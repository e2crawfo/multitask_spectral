12543 17
29 11 2 11 2 0 9 13 11 11 11 2 11 2 10 9 1 10 9 1 10 9 1 11 2 1 10 0 9 2
18 2 10 9 1 10 0 9 4 4 13 15 9 1 9 14 13 2 2
17 11 2 0 9 13 16 15 4 13 1 12 0 9 13 1 11 2
16 12 1 15 4 4 13 1 12 9 1 10 11 1 10 11 2
36 10 11 1 11 13 0 1 10 11 11 2 3 15 4 13 16 13 11 11 11 3 13 1 10 0 9 9 1 10 11 9 3 1 10 9 2
13 10 0 4 4 13 1 10 9 1 10 9 9 2
13 15 13 16 15 4 13 10 9 1 15 9 9 2
16 10 9 4 13 1 10 11 7 11 2 11 9 1 10 9 2
35 16 10 9 4 3 13 14 13 9 16 13 7 13 1 9 9 2 15 4 14 13 10 9 16 10 11 13 14 13 10 0 9 3 0 2
20 15 13 15 3 3 1 10 11 9 15 4 3 13 1 10 0 9 1 11 2
19 11 2 11 2 9 13 10 9 1 10 11 11 11 16 13 15 1 11 2
29 10 9 9 1 11 11 13 16 9 4 13 12 9 1 11 2 16 15 4 13 10 0 9 1 10 9 1 9 2
19 1 11 9 4 13 10 0 9 7 15 9 16 15 13 1 15 9 3 2
17 1 11 2 11 11 2 12 9 9 4 13 16 15 4 4 13 2
27 2 11 13 1 0 11 7 13 10 3 0 9 2 15 13 1 10 9 1 11 9 7 3 13 15 1 2
26 10 9 13 10 0 9 1 10 9 1 9 1 10 9 16 13 1 10 9 2 9 1 10 9 2 2
27 1 11 11 11 11 2 0 9 1 10 11 1 11 1 11 11 2 4 13 1 15 9 1 10 11 9 2
11 9 13 10 9 2 11 11 2 1 11 2
20 15 3 13 11 11 11 2 10 9 9 1 10 9 1 10 11 9 1 11 2
9 15 9 4 3 13 1 10 9 2
15 12 0 11 9 4 4 13 1 10 0 9 7 10 9 2
16 9 1 11 13 10 9 10 13 12 0 2 13 12 0 9 2
17 12 1 15 13 1 10 11 9 7 13 9 9 1 10 11 9 2
40 12 12 9 1 10 11 9 1 10 11 13 1 11 1 11 2 13 10 9 1 15 9 9 2 11 11 11 7 12 1 15 9 2 1 9 13 0 9 9 2
49 2 15 13 10 3 0 0 9 2 7 10 0 9 4 13 0 9 1 10 9 16 13 1 10 9 2 15 13 3 3 10 9 1 0 0 9 13 10 11 9 16 13 1 10 11 12 9 2 2
51 11 2 11 2 10 0 11 11 11 1 11 13 10 9 1 10 11 11 14 13 12 9 16 13 1 9 9 1 10 11 12 9 1 9 16 4 13 3 0 1 11 9 14 13 15 4 13 1 0 9 2
13 10 9 13 15 13 10 0 9 1 10 10 9 2
10 10 9 13 10 0 9 7 3 13 2
9 7 1 15 9 15 13 3 0 2
30 10 11 11 4 4 13 1 11 11 7 15 11 11 11 3 3 2 7 4 13 0 0 11 1 10 9 1 10 9 2
20 11 4 4 3 13 1 11 2 3 2 1 15 9 1 9 1 11 7 11 2
26 15 13 3 3 1 10 0 0 9 2 10 11 11 11 2 7 4 14 13 0 9 1 10 0 9 2
28 10 12 0 9 1 10 0 11 9 4 4 13 1 9 1 0 9 2 9 11 4 4 13 16 15 4 13 2
16 3 10 11 11 4 13 14 13 9 1 0 0 11 11 9 2
13 10 9 1 11 4 3 13 14 13 0 10 9 2
12 16 9 13 10 9 1 9 2 13 10 9 2
19 16 15 7 15 13 14 2 3 15 4 13 10 10 0 9 1 0 11 2
26 11 2 11 11 2 11 13 16 10 0 9 1 10 9 1 11 11 1 10 12 9 1 11 4 13 2
14 10 9 1 10 9 13 14 13 15 9 16 15 13 2
7 10 9 13 3 11 12 2
17 1 11 10 9 3 13 1 0 9 2 3 1 11 9 7 11 2
21 11 4 14 13 3 1 1 15 9 3 3 2 15 3 13 3 15 4 13 0 2
13 15 4 13 9 16 10 9 9 4 4 13 3 2
22 15 9 4 4 13 1 0 9 1 12 9 3 2 9 4 4 13 1 15 9 3 2
15 9 13 3 0 1 10 9 7 15 4 13 0 1 3 2
46 9 15 13 9 1 15 13 9 9 1 15 9 7 13 1 9 2 15 3 13 3 1 10 0 3 11 13 10 9 2 3 15 13 13 9 3 7 13 15 9 2 9 1 10 9 2
27 15 4 13 10 9 9 1 10 3 0 9 15 13 1 10 9 0 9 2 10 13 15 13 10 0 9 2
28 7 15 13 9 15 4 13 1 15 3 2 9 15 4 13 16 15 13 3 7 13 15 4 13 1 9 9 2
60 3 10 11 7 11 4 13 10 9 2 7 15 13 0 7 0 2 3 4 14 13 0 9 14 13 9 16 14 13 3 7 13 10 9 7 10 9 4 14 13 15 2 7 3 3 4 0 9 13 14 13 10 0 7 0 9 1 10 9 2
20 9 13 0 2 15 13 10 9 16 11 9 7 9 4 13 14 13 0 9 2
34 0 9 4 14 13 1 9 10 0 0 9 2 16 15 13 16 10 9 1 11 13 2 0 2 2 16 15 4 13 15 9 13 2 2
66 15 13 9 1 9 1 9 9 1 10 9 9 1 9 2 0 7 0 9 0 1 10 9 10 13 9 0 11 2 7 15 4 3 13 9 1 15 9 13 1 15 7 13 9 16 2 10 9 15 4 13 10 0 14 13 2 15 4 14 13 9 10 0 9 2 2
31 9 4 13 16 13 9 2 9 2 7 9 1 11 2 7 0 9 4 3 13 3 1 11 2 0 1 15 13 3 3 2
67 15 13 15 13 10 0 0 2 9 2 1 0 7 0 9 2 15 10 13 16 15 4 13 0 14 13 1 10 0 14 9 3 15 13 10 9 2 7 0 9 4 13 0 9 1 2 11 2 2 2 11 2 2 2 11 2 2 7 2 9 2 3 10 0 9 3 2
4 3 15 13 2
48 15 13 15 13 3 10 0 0 0 2 15 1 15 9 2 15 7 15 9 1 15 9 2 15 7 15 9 1 15 9 2 2 7 2 10 9 1 15 9 13 15 9 2 9 13 1 3 2
19 13 1 11 2 15 13 3 11 2 11 14 13 1 1 15 9 1 3 2
29 15 4 13 3 15 0 9 11 11 1 10 9 2 7 15 4 13 10 9 1 9 3 13 15 1 11 2 11 2
37 2 15 4 13 9 2 2 2 0 9 4 13 9 7 0 9 2 2 7 2 15 4 13 9 9 1 9 2 13 10 15 13 14 13 1 15 2
42 15 4 3 13 10 0 9 3 15 13 16 0 9 4 13 1 10 11 1 10 9 1 9 7 9 1 11 11 2 11 2 7 3 3 15 13 0 1 11 2 11 2
44 9 15 13 15 11 11 1 10 11 11 2 11 11 2 10 0 9 2 13 1 11 2 11 13 10 0 9 1 10 11 7 15 13 16 0 9 4 13 10 9 1 0 9 2
13 3 12 11 4 13 0 7 12 0 1 11 3 2
11 11 2 11 11 13 16 11 4 13 11 2
70 11 9 13 10 9 13 1 11 11 11 11 2 10 11 2 11 9 1 11 11 1 10 0 9 2 10 11 1 11 2 2 1 10 15 13 16 2 16 13 0 9 4 14 3 13 1 11 2 7 1 10 9 15 4 13 16 11 13 15 1 9 14 13 15 16 13 0 9 2 2
76 15 13 16 2 11 4 14 13 9 1 10 9 1 9 7 9 2 15 4 13 1 1 11 1 9 16 10 9 4 13 1 11 16 10 0 9 14 13 2 2 7 16 2 10 9 4 13 3 10 0 9 1 11 7 11 4 4 13 2 13 2 7 13 1 1 10 11 11 3 1 15 9 7 9 2 2
23 11 14 9 9 1 10 9 1 11 4 13 9 1 12 1 10 3 0 0 9 1 9 2
39 15 10 13 15 13 2 7 3 1 10 9 2 15 13 0 0 9 7 9 1 3 15 13 7 10 9 11 4 13 1 10 9 1 9 13 1 10 9 2
2 9 2
11 3 15 4 13 11 7 13 15 0 9 2
13 15 13 14 10 9 1 9 2 9 7 13 9 2
16 15 13 10 9 14 13 15 13 7 3 15 4 13 10 9 2
47 15 4 10 0 0 11 2 11 11 11 11 1 10 11 1 11 11 2 9 1 12 1 10 9 9 1 11 13 16 15 13 10 0 9 1 10 0 9 2 0 9 9 1 0 9 13 2
24 15 4 3 13 1 10 11 11 11 11 1 10 9 9 13 10 11 1 11 10 13 10 13 2
42 12 1 10 3 0 9 1 0 9 13 16 10 11 0 9 9 1 12 13 0 9 1 0 9 9 1 13 9 2 7 16 0 9 4 4 3 13 1 9 1 9 2
38 0 9 3 13 15 14 13 0 2 3 16 10 11 1 11 9 1 11 11 2 11 7 11 1 11 1 11 11 2 11 1 11 2 13 15 1 12 2
6 11 9 2 12 9 3
50 1 10 0 9 2 15 4 13 10 0 7 0 9 1 9 7 2 1 10 0 9 2 9 9 1 10 9 1 13 9 1 10 0 11 11 2 11 2 10 4 4 13 1 10 11 9 16 13 3 2
33 10 0 11 2 11 11 11 11 2 13 10 0 9 1 11 10 4 13 1 9 1 0 9 7 13 16 15 13 10 0 9 9 2
25 3 2 1 11 12 2 10 11 13 11 11 1 10 11 11 2 11 13 2 10 13 10 0 9 2
5 3 13 10 9 2
33 10 0 9 1 9 2 13 9 9 1 9 7 9 1 11 2 11 2 7 11 2 10 4 4 13 1 12 2 13 1 10 9 2
32 2 10 9 1 10 9 9 2 10 9 1 9 14 0 9 2 10 9 1 9 1 9 7 9 2 7 10 9 1 0 9 2
60 10 9 1 9 1 10 9 1 9 1 9 13 1 10 11 9 1 10 12 9 2 11 2 11 2 7 11 2 1 10 0 9 4 13 1 0 0 9 2 10 9 9 4 13 3 2 10 9 1 3 0 9 4 13 2 7 9 4 13 2
24 1 10 9 2 15 4 3 13 3 0 15 4 13 1 10 9 15 9 4 13 1 9 9 2
9 15 13 10 9 14 13 1 11 2
19 13 3 2 13 4 13 15 9 7 15 13 0 1 10 9 1 13 9 2
9 15 13 10 9 1 9 1 11 2
12 13 10 1 10 13 9 7 13 15 0 9 2
17 10 9 13 10 0 9 10 13 7 3 13 1 10 9 13 11 2
4 11 9 11 13
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
19 15 4 13 0 16 13 10 9 15 13 7 15 15 13 10 13 3 0 2
2 9 2
48 1 10 9 1 10 9 15 13 10 9 1 0 9 7 15 13 15 1 9 9 2 0 1 0 2 2 7 13 3 10 9 1 15 9 13 13 2 15 13 15 13 14 9 7 13 10 9 2
14 13 10 0 9 13 9 10 13 10 9 1 9 9 2
5 15 3 4 13 2
32 4 14 13 14 13 15 9 4 13 7 4 3 13 1 11 7 11 9 2 15 4 13 10 9 1 10 9 1 9 1 11 2
19 10 11 11 14 11 2 8 2 13 0 9 14 13 10 9 1 10 9 2
26 12 1 15 13 10 11 7 11 11 2 3 10 9 4 13 1 10 11 1 10 0 9 1 10 9 2
23 3 10 0 9 13 13 0 2 0 9 2 0 0 9 2 8 4 13 9 1 15 9 2
26 11 7 15 13 10 9 15 4 13 0 1 10 9 1 0 9 2 14 13 10 0 9 13 10 9 2
24 10 9 14 13 7 13 15 10 3 13 3 0 2 7 13 15 3 0 1 10 9 15 13 2
7 13 9 2 15 9 2 11
16 15 13 0 14 13 11 14 9 4 4 13 14 13 10 9 2
33 15 4 10 0 11 2 11 9 7 9 9 1 11 11 7 11 11 2 11 13 15 1 10 9 1 10 0 0 9 1 10 9 2
40 16 10 11 7 11 4 13 14 13 7 13 3 12 2 9 1 10 0 12 11 2 11 9 2 10 0 9 13 14 1 0 9 1 11 2 11 7 11 11 2
9 10 9 13 10 9 14 13 9 2
42 15 13 8 2 13 7 13 11 11 11 2 10 0 0 2 9 2 15 4 13 10 9 1 12 7 4 13 3 15 9 1 10 11 11 1 10 11 7 11 2 11 2
19 11 4 4 13 14 13 15 9 9 1 10 0 9 1 11 2 11 9 2
39 15 0 9 4 13 0 9 1 11 11 7 11 11 11 2 3 3 1 3 12 0 11 2 11 9 2 3 12 1 15 10 11 4 13 1 1 10 11 2
36 11 13 9 1 11 1 12 2 1 10 9 2 0 9 13 3 2 7 1 10 3 12 9 1 9 9 13 1 10 0 0 9 9 2 11 2
34 11 3 13 10 11 11 11 2 10 3 13 11 11 7 11 2 11 2 7 13 1 10 0 9 1 11 11 2 3 1 10 11 9 2
34 16 11 2 11 4 13 11 7 13 10 0 9 1 15 1 11 0 9 2 15 4 13 14 13 10 11 1 9 1 0 9 7 9 2
20 15 4 3 13 9 1 10 0 9 1 0 9 2 10 13 3 10 0 9 2
15 10 10 13 3 0 2 1 1 0 11 2 11 9 9 2
18 7 3 13 15 0 16 10 0 9 1 0 9 4 3 13 1 11 2
18 9 2 10 11 4 13 15 15 4 14 13 10 9 1 10 0 9 2
39 1 10 12 9 2 15 4 13 11 14 13 1 15 9 7 13 1 9 1 10 0 9 2 7 14 13 10 0 2 11 11 11 2 10 3 13 15 9 2
37 1 10 0 2 9 4 4 13 1 10 0 11 11 2 11 7 11 11 14 11 2 15 4 13 10 11 1 0 9 16 3 13 1 10 0 9 2
23 1 10 0 9 2 10 11 4 0 2 13 11 7 11 1 10 0 9 1 10 11 9 2
26 11 2 11 13 14 13 11 14 9 1 9 16 13 10 11 1 10 0 9 1 10 9 1 15 9 2
21 10 11 9 13 3 0 9 2 7 3 10 9 1 0 9 2 16 11 3 13 2
24 8 2 13 11 7 13 10 0 9 1 10 11 16 13 1 10 0 9 9 1 10 11 9 2
21 9 2 10 11 4 13 16 3 13 11 2 7 13 10 9 16 13 1 15 9 2
15 10 0 9 4 3 3 13 1 3 3 0 9 7 9 2
7 15 4 13 14 4 13 2
44 7 11 14 0 9 4 3 14 13 1 10 9 16 13 0 9 2 7 10 11 9 4 13 14 3 13 0 9 1 11 14 13 15 9 1 7 9 1 10 11 11 7 11 2
49 11 14 0 9 4 13 1 9 1 11 14 9 14 13 1 9 3 7 3 2 10 13 3 1 10 0 9 7 13 1 10 9 9 1 11 2 11 1 15 9 1 9 0 14 13 10 11 11 2
24 11 13 10 11 11 3 3 3 0 2 1 10 9 2 14 13 3 0 9 7 13 0 9 2
17 8 2 13 11 10 11 2 13 10 11 11 14 0 9 1 15 2
22 9 2 11 13 3 0 9 1 11 2 11 2 7 1 0 9 15 4 14 13 3 2
32 16 13 3 1 0 9 7 9 1 0 9 2 10 11 4 13 0 14 13 11 1 15 9 2 16 16 15 13 1 10 9 2
17 3 2 10 11 3 13 11 2 11 7 4 13 2 3 10 11 2
22 10 9 16 13 10 11 2 3 2 13 14 4 13 14 13 13 11 2 11 10 9 2
27 10 11 13 14 13 3 15 0 2 9 9 1 10 9 7 13 9 16 13 9 7 13 9 1 0 9 2
12 15 13 10 11 1 11 2 3 10 11 11 2
25 3 3 2 10 3 10 11 9 4 4 13 1 9 1 3 2 0 0 7 0 9 2 10 0 2
30 13 10 0 1 1 11 13 14 3 3 0 10 9 9 1 11 2 11 1 10 0 9 16 13 10 11 7 0 3 2
50 10 9 14 13 1 9 13 16 0 0 9 7 11 7 0 0 9 13 0 14 13 3 3 0 1 10 11 1 11 1 11 2 11 9 2 7 15 4 13 0 14 13 15 14 9 1 10 0 9 2
16 11 11 11 13 11 16 11 11 13 10 9 0 14 13 11 2
35 10 9 1 10 9 13 16 11 13 10 9 0 14 13 11 3 15 13 1 12 2 3 10 9 1 0 9 3 13 15 1 15 0 9 2
11 13 15 3 13 10 0 11 9 1 12 2
10 2 11 13 9 14 9 9 1 0 9
4 11 12 2 12
11 9 13 1 2 12 9 11 2 12 11 2
5 11 2 11 2 2
42 11 11 11 11 11 4 13 0 9 16 13 0 14 13 10 9 1 12 0 9 0 9 2 7 11 11 11 13 11 2 4 2 7 3 4 2 13 1 2 10 9 2
33 10 0 2 9 1 10 12 0 0 9 13 11 1 10 0 9 9 9 13 1 11 11 2 10 0 9 1 11 2 11 1 11 2
1 11
16 11 13 11 14 13 10 9 1 11 2 11 2 11 7 11 2
32 11 13 3 0 14 13 10 0 9 1 10 9 1 10 9 1 11 2 13 1 0 11 11 11 2 11 3 1 2 11 2 2
7 15 4 14 13 10 9 2
14 2 4 15 13 10 9 15 13 1 9 1 11 2 2
18 11 13 2 13 1 11 11 11 2 15 13 9 1 10 9 11 12 2
14 2 13 2 13 2 13 15 12 9 2 2 13 11 2
22 11 13 2 2 6 2 15 13 12 9 1 12 9 1 12 0 9 2 2 2 2 2
36 11 2 16 13 10 9 1 10 9 1 11 2 3 13 2 2 10 0 0 9 2 15 4 3 4 13 2 3 13 2 10 9 13 1 9 2
24 15 13 10 9 4 13 14 13 9 1 10 9 7 15 13 15 13 0 9 1 10 9 2 2
18 11 13 10 9 11 13 11 1 9 1 15 9 1 11 14 0 9 2
34 2 15 13 15 0 16 10 9 1 11 1 15 9 2 10 9 14 0 9 2 4 13 10 0 9 1 2 0 9 2 2 11 13 2
38 2 3 2 15 13 15 3 3 0 16 15 13 10 9 1 10 9 10 3 0 9 13 0 9 2 3 16 13 15 0 9 1 10 11 11 11 11 2
11 10 9 1 11 11 3 13 11 14 9 2
29 2 15 13 3 0 16 10 9 14 13 10 9 1 3 13 9 2 2 13 11 11 2 9 1 10 11 11 11 2
66 3 3 4 11 14 13 15 11 11 11 13 2 15 13 14 4 13 9 2 9 1 2 13 9 2 2 7 3 13 3 14 13 16 10 9 1 10 13 0 9 7 10 9 1 9 1 10 11 9 2 3 10 9 14 0 9 1 10 11 2 4 13 2 9 2 2
39 11 13 15 9 1 0 1 1 10 9 14 9 1 11 11 11 11 14 9 14 13 1 16 13 11 1 11 2 16 16 15 3 13 1 9 1 10 9 2
16 15 4 14 13 15 3 0 15 13 11 14 9 1 10 9 2
18 15 3 13 15 13 1 2 10 9 2 2 0 14 13 11 14 9 2
22 15 3 13 10 9 15 15 4 13 1 2 16 15 13 10 9 1 0 2 0 9 2
16 15 3 13 0 9 3 1 9 2 13 9 1 2 9 2 2
34 7 2 15 4 14 13 15 13 14 13 9 1 11 11 2 1 15 0 9 7 0 0 9 2 10 0 10 0 9 9 1 10 11 2
15 15 4 14 13 3 9 4 13 3 0 16 13 1 0 2
18 11 13 3 14 13 0 9 1 11 1 12 2 13 9 3 10 9 2
39 16 11 4 13 1 10 11 1 11 12 2 1 0 9 1 10 11 2 9 1 15 9 13 14 13 0 11 7 4 3 4 13 1 9 9 1 11 15 2
20 15 13 10 9 10 11 13 4 13 2 9 2 1 10 9 1 9 1 12 2
26 3 2 12 9 1 11 14 9 1 11 13 16 16 15 13 10 9 2 11 4 4 13 14 13 15 2
18 10 9 13 16 11 3 13 3 0 1 0 9 3 16 11 4 3 2
39 3 2 13 3 11 4 13 1 10 9 13 9 7 13 0 9 1 10 9 14 13 3 1 10 11 2 15 4 3 13 16 11 13 0 3 16 11 13 2
43 15 13 15 11 14 9 9 13 1 15 9 2 2 11 13 16 10 11 4 13 10 0 9 14 13 13 9 2 16 13 9 1 11 7 11 1 10 9 9 1 11 11 2
28 11 13 10 0 9 1 11 2 7 13 16 10 11 13 10 0 9 16 13 9 1 10 11 7 10 11 2 2
10 15 4 14 13 11 13 10 1 15 2
5 1 11 14 11 11
3 1 11 11
6 11 2 11 12 2 12
32 16 10 0 9 3 13 1 10 11 9 2 10 4 13 13 16 10 9 4 13 3 1 10 11 16 13 10 9 1 0 9 2
26 11 2 3 2 13 3 0 1 11 7 13 0 14 13 1 0 9 3 3 3 16 4 10 11 11 2
24 3 2 1 10 0 9 1 9 1 11 13 0 11 11 11 11 7 15 0 9 1 10 11 2
10 4 15 2 3 2 3 13 0 9 2
21 10 0 9 11 13 13 3 1 0 9 7 1 10 0 9 1 0 0 9 9 2
24 10 9 1 10 11 9 9 1 10 0 2 9 9 1 11 7 10 0 9 4 13 9 9 2
27 15 2 1 9 2 4 13 0 9 1 11 7 4 13 15 3 0 16 9 1 10 9 4 3 13 3 2
23 16 11 13 1 0 9 1 11 12 2 10 0 0 0 9 2 11 2 4 14 4 13 2
41 15 4 13 14 13 10 12 0 9 2 7 15 4 13 9 1 0 9 14 13 15 14 13 1 10 11 11 2 10 9 1 0 9 10 11 13 1 10 12 9 2
34 10 0 9 1 10 9 1 10 11 9 7 15 9 1 11 14 9 9 4 2 3 2 3 13 15 0 9 1 10 9 1 0 9 2
41 16 15 4 3 13 2 1 0 9 2 16 11 11 13 9 1 10 9 1 0 9 9 7 3 13 0 9 2 15 13 14 0 16 15 3 13 10 9 1 11 2
29 10 11 15 4 13 0 14 13 15 14 13 10 0 9 1 10 11 11 7 10 11 11 4 14 13 1 0 9 2
10 11 3 13 9 0 14 13 10 11 2
31 1 10 9 2 1 1 10 0 9 2 15 3 13 1 2 10 2 9 9 1 10 11 14 13 1 10 9 1 10 9 2
14 15 4 14 13 0 9 14 13 9 1 11 1 11 2
22 1 10 0 9 2 11 13 10 0 7 0 9 9 2 7 4 13 15 0 9 9 2
13 15 0 9 4 3 13 1 10 0 9 1 12 2
30 16 15 13 0 14 13 3 0 11 13 10 0 9 1 11 2 15 13 14 3 0 14 13 10 9 1 10 0 9 2
16 10 9 1 0 11 1 10 11 9 13 10 0 7 13 9 2
19 0 9 2 0 13 1 0 0 0 9 1 0 9 7 9 2 4 13 2
35 10 11 13 14 13 15 1 0 9 1 10 11 11 1 10 11 11 1 11 2 15 12 2 0 11 11 9 4 13 1 10 11 11 11 2
15 0 7 0 9 13 0 1 0 0 0 0 9 7 9 2
25 10 3 0 11 2 15 3 13 10 0 9 1 11 14 11 11 11 2 3 13 7 13 1 11 2
19 15 3 13 10 0 9 1 11 11 11 2 10 9 1 11 2 0 11 2
29 0 1 11 2 10 9 13 10 9 3 1 10 0 7 0 11 11 11 11 2 15 13 0 0 9 1 0 11 2
20 10 0 9 4 4 13 1 11 11 14 9 2 7 4 3 13 7 13 15 2
13 15 4 3 13 15 0 9 1 0 7 0 11 2
48 15 13 0 16 0 0 11 4 13 1 15 11 9 1 11 2 7 15 13 0 16 0 11 4 13 0 3 1 0 9 9 1 10 9 16 15 4 13 1 10 0 9 14 13 0 0 9 2
27 0 0 9 3 13 1 10 11 7 1 11 2 7 15 1 11 13 13 0 9 1 9 1 11 7 11 2
34 0 9 0 1 11 7 11 13 1 10 9 9 1 11 1 11 2 7 3 13 1 10 9 1 10 11 9 2 10 13 0 1 11 2
20 0 0 9 9 3 3 13 1 10 11 2 7 15 1 0 11 13 10 9 2
23 16 11 11 14 9 13 16 0 0 9 4 13 3 1 9 2 15 13 3 0 14 13 2
18 10 11 1 10 0 0 7 0 9 13 13 3 10 9 9 1 11 2
28 16 3 10 9 1 9 7 9 4 4 13 1 11 2 15 9 4 13 0 14 13 1 10 9 14 9 9 2
17 10 0 9 4 3 4 13 1 9 1 10 11 7 1 0 11 2
27 11 14 9 9 4 3 13 1 9 1 15 9 2 10 4 3 4 13 16 13 9 1 9 1 10 11 2
29 11 11 14 0 0 9 1 3 9 1 10 13 11 11 7 15 0 9 1 10 0 9 4 13 0 9 7 9 2
12 10 9 4 13 1 10 0 9 2 13 11 2
28 10 9 1 10 0 9 1 9 9 2 1 10 11 11 7 1 11 2 4 3 13 2 14 13 2 0 9 2
35 11 11 2 8 2 13 10 9 1 0 11 11 9 1 10 11 1 11 7 9 1 2 11 11 7 11 11 2 2 11 11 2 12 2 2
11 10 11 11 13 10 9 1 9 1 11 11
26 11 13 16 10 13 9 9 1 11 7 11 11 4 13 0 9 14 13 1 10 9 13 10 0 9 9
23 7 15 13 0 9 1 10 9 16 10 0 8 2 11 11 9 9 4 13 1 10 9 2
30 7 15 4 3 13 9 1 10 11 11 11 2 11 2 10 4 13 1 10 11 1 10 11 0 9 13 1 11 11 2
43 3 1 10 12 0 9 13 1 12 2 10 0 9 9 13 3 0 3 3 1 11 11 7 10 11 9 7 3 1 10 0 9 15 13 15 10 9 1 15 9 14 9 2
5 11 0 1 11 11
3 1 11 11
3 11 11 2
59 16 11 13 0 14 13 1 10 2 9 9 9 2 1 11 11 2 15 13 0 16 4 13 1 10 0 9 1 10 9 9 14 12 9 2 0 0 9 10 4 13 0 9 1 0 11 7 10 0 9 2 13 3 12 0 1 10 9 2
33 7 15 13 10 9 1 10 9 1 10 0 9 9 10 13 1 10 9 1 0 0 11 11 11 14 12 2 9 9 1 11 3 2
37 13 1 11 11 11 11 2 11 11 9 1 10 11 11 11 2 10 12 2 9 9 9 1 11 7 10 11 11 1 11 11 2 11 2 4 13 2
21 1 10 9 2 15 13 2 11 14 9 13 0 14 13 1 0 9 1 0 9 2
24 2 10 0 0 9 4 14 13 14 13 10 9 7 4 13 0 16 13 10 11 16 13 12 2
21 7 10 11 13 16 16 15 13 1 10 9 16 13 10 9 2 2 11 13 11 2
16 11 13 12 9 1 9 1 10 11 1 11 12 7 11 12 2
28 7 0 11 2 10 9 3 13 1 1 9 13 9 2 3 2 1 10 9 1 9 2 9 16 13 3 3 2
43 11 14 11 9 13 10 12 2 9 9 1 11 11 1 0 11 11 11 11 1 10 0 9 14 13 10 9 9 10 4 13 14 13 10 9 10 11 3 13 1 11 12 2
60 11 13 9 1 7 11 7 10 0 11 9 11 11 1 10 9 9 1 11 1 9 2 7 0 0 9 9 11 11 7 0 9 11 11 13 13 2 9 9 1 10 0 9 3 11 1 10 9 14 13 10 9 9 1 9 2 0 9 13 2
7 7 15 2 3 2 13 2
12 11 2 3 2 13 14 13 1 10 0 9 2
52 13 1 0 0 9 9 11 11 11 2 10 9 1 11 14 9 13 1 10 9 16 10 11 4 13 10 8 8 9 1 10 9 7 9 1 10 9 7 4 13 10 9 1 0 9 1 10 9 1 15 9 2
54 10 9 1 11 14 0 9 1 10 11 9 14 13 13 10 12 8 2 11 11 11 11 2 10 3 13 1 10 9 1 10 0 11 2 11 13 10 0 9 9 4 3 13 10 9 1 10 0 9 7 15 0 9 2
48 11 2 15 3 13 10 0 11 2 13 11 11 1 11 11 2 13 1 10 9 1 10 0 9 14 13 7 3 13 10 11 2 11 13 10 0 9 0 16 13 10 9 1 10 0 9 9 2
45 2 10 11 13 3 7 15 9 13 0 1 15 1 0 9 7 10 11 13 3 0 16 15 4 14 13 10 9 2 1 11 2 14 13 10 9 2 2 11 13 11 1 10 9 2
15 1 12 2 10 11 11 3 13 10 9 9 1 0 9 2
25 1 10 9 2 10 0 0 0 9 4 13 7 10 0 9 4 13 1 9 1 10 9 7 9 2
23 3 2 9 1 11 7 11 3 13 7 13 1 9 1 11 9 7 10 0 9 9 9 2
13 3 12 0 9 4 13 1 10 9 1 10 9 2
26 11 13 14 13 3 15 9 1 11 11 1 12 13 10 9 1 11 11 2 10 0 9 1 0 9 2
31 0 11 2 10 0 9 13 1 11 14 13 10 11 14 13 3 1 10 9 9 13 1 10 9 9 9 1 5 12 12 2
39 11 14 0 9 2 11 11 2 15 13 1 0 9 1 10 9 9 16 10 9 4 4 13 2 13 3 1 9 1 11 7 11 1 0 11 10 0 9 2
20 15 13 1 10 2 0 9 1 9 2 7 13 10 9 1 9 1 10 9 2
52 10 11 14 0 9 2 11 2 13 1 10 9 13 16 2 10 9 1 10 0 9 4 14 4 13 1 10 9 7 9 1 9 9 2 7 13 14 4 13 1 10 9 1 9 1 10 9 1 0 9 2 2
23 7 15 13 0 9 1 10 9 16 10 0 8 2 11 11 9 9 4 13 1 10 9 2
30 7 15 4 3 13 9 1 10 11 11 11 2 11 2 10 4 13 1 10 11 1 10 11 0 9 13 1 11 11 2
43 2 11 13 16 10 13 9 9 1 11 7 11 11 4 13 11 9 14 13 1 10 9 13 10 0 9 9 2 2 11 9 1 9 11 11 4 13 16 13 1 10 9 2
40 15 13 16 0 9 1 10 9 1 11 14 0 0 9 13 9 9 11 11 11 11 4 2 13 9 1 11 16 9 13 1 9 1 10 9 1 10 9 2 2
57 7 11 13 1 16 11 4 13 3 2 13 14 13 0 3 2 3 2 1 11 11 16 3 16 15 3 13 14 13 10 9 1 12 12 0 11 1 10 0 9 1 11 11 2 13 1 11 11 14 11 9 1 10 0 11 11 2
43 3 1 10 12 0 9 13 1 12 2 10 0 9 9 13 3 0 3 3 1 11 11 7 10 11 9 7 3 1 10 0 9 15 13 15 10 9 1 15 9 14 9 2
53 10 0 9 2 3 2 1 10 0 0 9 13 16 11 14 13 15 0 0 9 2 16 11 11 4 3 4 13 1 14 13 0 0 9 1 1 10 13 9 16 9 2 9 7 9 4 14 13 10 9 1 9 2
25 1 10 9 2 11 13 15 3 2 2 15 4 14 13 10 0 9 16 15 13 10 0 9 2 2
4 11 11 11 12
44 13 1 10 0 9 2 10 11 1 11 4 13 10 0 7 0 9 10 4 13 1 10 9 1 10 9 1 3 10 10 0 9 15 4 4 13 3 16 0 9 4 3 13 2
25 1 12 9 9 10 4 13 10 0 9 4 4 13 2 16 10 13 1 9 9 7 9 1 9 2
24 3 3 2 9 1 10 0 2 0 9 2 9 1 10 9 4 13 14 3 13 10 10 9 2
4 11 13 10 9
2 11 11
35 16 0 11 9 1 9 2 1 3 11 11 2 4 13 1 9 1 9 10 15 13 0 14 13 1 2 0 4 13 3 0 1 11 11 2
34 12 9 3 2 0 11 11 11 13 0 3 10 9 1 10 0 11 9 2 11 11 11 2 13 11 7 13 10 9 1 3 0 9 2
34 16 11 14 9 4 4 13 10 11 11 15 4 2 13 2 16 13 10 0 9 1 11 3 1 10 9 1 11 2 15 13 10 9 2
18 10 9 13 16 11 13 3 3 10 9 1 9 1 10 9 1 11 2
10 10 9 4 3 13 1 10 11 11 2
52 9 2 7 15 3 13 9 1 10 11 0 0 9 9 0 1 11 11 2 15 4 3 13 14 13 11 1 15 0 9 1 10 0 9 1 11 2 13 10 3 0 9 1 11 13 10 9 1 10 9 9 2
25 11 13 15 15 13 16 11 7 11 2 10 4 13 10 9 1 10 9 12 9 3 2 13 3 2
31 3 2 11 11 4 13 10 9 1 9 1 10 9 10 4 13 13 0 9 1 1 9 13 14 13 11 1 10 0 11 2
56 11 11 13 15 1 10 9 1 15 9 1 9 7 2 1 11 11 2 15 13 14 13 10 9 1 9 0 1 9 2 2 10 9 1 11 9 4 3 3 13 1 10 0 9 14 13 3 3 10 11 1 11 3 1 11 2
25 15 2 11 14 9 1 11 11 11 4 4 13 2 13 10 2 9 2 10 10 11 9 4 13 2
15 15 13 3 3 0 16 15 10 9 1 11 11 4 13 2
57 10 9 4 1 9 13 10 0 9 1 10 11 9 16 13 10 9 1 10 0 9 1 10 9 1 10 0 2 9 11 2 10 11 2 13 11 7 10 3 0 11 11 2 16 10 0 9 13 9 1 9 14 9 7 0 9 2
32 1 9 2 10 11 11 4 13 9 1 10 11 11 7 0 9 3 11 13 0 7 13 10 9 2 9 7 9 9 1 11 2
50 10 0 9 1 11 1 11 4 13 0 1 10 10 9 2 1 1 10 0 0 9 13 1 10 11 11 11 7 10 11 11 2 10 4 13 14 13 10 9 1 11 1 15 0 9 1 11 1 12 2
44 13 1 10 0 9 2 10 11 1 11 4 13 10 0 7 0 9 10 4 13 1 10 9 1 10 9 1 3 10 10 11 9 15 4 4 13 3 16 0 9 4 3 13 2
25 3 12 9 9 10 4 13 10 0 9 4 4 13 2 16 10 13 1 9 9 7 9 1 9 2
24 3 3 2 9 1 10 0 2 0 9 2 9 1 10 9 4 13 14 3 13 10 10 9 2
21 3 2 15 9 4 13 1 9 1 10 2 9 2 1 0 9 1 10 0 9 2
29 1 11 12 2 10 11 11 3 13 10 11 9 10 13 9 1 9 1 10 9 11 4 13 14 13 11 11 0 2
31 3 1 15 2 10 9 4 13 14 13 3 11 11 14 0 9 16 15 13 1 15 9 3 10 11 13 0 9 1 11 2
48 10 11 11 11 7 10 13 9 9 10 13 15 9 4 13 0 9 1 11 7 2 1 0 1 15 2 10 9 10 4 13 13 10 9 13 3 1 0 9 7 1 15 0 9 1 11 11 2
62 16 11 13 14 11 7 16 10 2 9 2 13 2 11 11 11 4 3 13 14 13 0 9 2 4 14 13 10 9 2 1 15 4 13 0 0 2 9 2 7 2 9 2 0 14 13 7 13 9 1 10 9 1 10 0 9 1 11 11 7 11 2
49 1 0 9 2 11 13 10 9 2 9 7 3 13 1 1 10 9 1 9 10 13 1 10 0 11 4 14 13 15 1 10 9 10 13 10 9 2 9 9 1 11 11 7 11 11 11 4 3 2
50 15 13 10 9 9 1 11 10 13 1 16 11 13 1 10 0 9 1 9 9 1 12 2 13 1 16 10 0 9 1 10 0 9 16 9 2 3 0 9 2 13 1 10 9 1 10 9 13 11 2
56 10 9 1 15 13 16 11 4 13 1 10 0 9 9 1 11 2 3 10 9 10 10 9 1 11 13 1 15 0 9 1 9 7 9 16 13 10 9 1 9 13 11 3 1 9 10 0 9 13 10 11 11 7 11 11 2
40 1 3 2 11 4 13 9 16 3 13 16 3 10 9 9 4 13 0 1 10 0 9 2 10 9 1 9 10 4 13 1 10 9 1 9 1 11 3 3 2
46 3 1 15 0 14 3 13 1 1 10 0 9 1 9 9 1 11 11 2 11 11 4 3 13 11 11 14 9 2 13 15 14 13 1 15 0 9 13 16 10 11 13 1 15 9 2
56 16 10 11 11 9 13 16 15 13 0 9 1 9 2 11 4 13 10 9 1 9 2 13 10 0 2 7 3 3 13 1 10 9 7 13 10 0 9 1 9 10 4 13 3 3 11 7 11 11 7 11 7 11 3 3 2
17 10 12 9 10 4 13 16 15 13 10 9 1 11 11 13 11 2
68 1 11 11 11 2 11 4 13 1 1 11 11 7 11 11 11 11 4 13 14 13 3 0 9 2 13 9 16 3 13 11 1 9 1 11 7 13 11 1 10 0 9 1 10 11 11 11 2 3 13 11 1 10 0 9 1 10 2 0 12 2 10 4 14 3 13 3 2
15 16 11 11 3 2 10 11 13 10 9 1 10 11 11 11
22 11 11 2 10 9 1 9 2 13 9 1 9 1 10 11 11 1 11 11 2 11 2
3 11 11 12
2 6 2
10 15 10 13 16 11 11 13 1 11 2
31 12 0 9 2 1 10 15 13 9 1 10 3 2 13 2 3 2 13 9 10 13 15 14 13 15 2 9 1 9 2 2
33 15 3 13 3 11 11 13 11 11 7 13 15 9 1 10 11 11 11 11 1 10 2 12 11 12 2 9 13 3 1 13 9 2
20 1 15 9 1 10 11 2 11 11 13 10 11 2 12 11 11 9 2 9 2
17 10 11 2 12 13 9 1 10 11 9 1 11 12 7 11 12 2
32 1 10 9 2 11 2 12 9 4 13 1 1 11 11 11 2 11 11 7 11 11 1 11 2 7 11 7 11 11 1 11 2
7 2 13 3 1 9 2 2
18 3 3 16 11 11 13 2 15 7 15 9 4 4 4 13 1 11 2
21 1 10 10 3 2 13 9 2 4 9 13 16 3 11 11 3 13 14 13 9 2
13 7 2 13 15 13 2 13 0 9 9 13 0 2
9 15 4 14 13 3 9 13 15 2
29 10 9 2 15 13 2 10 9 1 0 9 2 4 3 13 10 9 1 11 11 14 9 1 10 11 11 11 11 2
19 1 9 2 4 15 13 16 11 11 13 3 0 9 1 9 1 11 11 2
23 15 13 13 10 9 1 10 9 13 1 15 1 10 9 1 15 2 9 1 11 11 2 2
7 13 3 14 13 10 9 2
1 2
5 11 14 11 11 9
12 16 15 13 1 11 14 9 2 3 13 10 9
17 15 4 15 3 13 1 11 11 11 14 9 1 10 11 11 11 2
11 16 15 4 14 13 1 1 9 1 11 2
6 16 15 13 10 9 2
7 16 15 9 13 15 3 2
30 9 9 1 10 11 14 9 1 10 11 4 13 14 13 1 12 0 9 1 10 9 2 1 10 9 1 3 9 0 2
16 3 3 1 10 9 2 3 2 1 0 2 13 15 11 13 2
10 10 0 9 13 10 11 1 11 12 2
11 3 3 2 15 13 10 0 9 1 9 2
6 12 9 1 0 9 2
8 12 2 12 9 1 9 9 2
10 12 2 12 9 1 9 2 9 9 2
19 15 13 12 9 14 13 1 2 7 15 13 0 9 9 13 3 3 3 2
7 15 13 0 2 9 9 2
14 1 10 9 15 13 3 2 11 4 13 3 12 9 2
6 3 12 9 1 9 2
3 12 9 2
18 1 9 2 11 13 13 2 13 1 9 1 9 1 11 2 12 9 2
14 16 15 13 2 15 13 9 1 15 11 11 9 9 2
20 1 10 9 2 9 4 13 14 13 10 9 1 12 9 14 13 15 0 9 2
45 13 1 9 13 3 10 9 2 11 13 12 9 1 15 0 9 2 11 12 1 11 12 2 16 15 13 1 11 12 2 15 9 3 4 13 1 10 11 2 1 2 11 9 2 2
9 11 13 12 9 1 12 5 12 2
25 2 1 0 9 2 11 13 0 9 14 13 10 9 1 15 0 12 9 9 1 12 5 12 3 2
3 2 11 2
9 15 13 12 9 1 12 5 12 2
10 7 15 13 12 9 1 12 5 12 2
22 10 9 13 16 1 15 0 12 9 2 11 14 3 13 1 2 15 13 1 10 9 2
5 4 15 13 15 2
53 15 13 10 9 1 11 12 2 10 9 10 4 13 10 9 1 3 0 9 9 2 3 11 2 13 2 2 13 1 0 9 11 11 2 7 13 2 0 2 2 13 1 11 11 2 9 1 10 11 11 11 2 2
15 11 13 1 9 14 13 1 11 14 13 1 10 11 9 2
6 15 0 9 13 6 2
22 9 1 15 13 14 0 2 13 13 11 11 11 2 15 13 1 11 1 12 7 12 2
16 2 1 12 2 15 13 10 0 9 1 9 2 2 11 13 2
19 2 10 11 11 4 13 1 2 7 10 11 11 4 13 9 1 9 9 2
29 1 12 7 12 2 16 15 13 10 9 2 0 7 11 2 7 15 13 10 9 7 13 14 13 3 2 10 9 2
12 1 9 2 15 4 13 15 13 15 9 2 2
5 3 11 13 13 2
23 1 11 12 1 11 12 2 15 13 3 12 9 2 3 0 2 7 0 14 13 15 9 2
27 3 2 1 12 2 16 11 13 9 14 13 10 11 7 13 1 11 11 11 2 15 3 13 13 1 3 2
25 1 11 7 11 1 12 2 15 13 12 9 2 0 14 13 10 9 9 1 10 12 5 12 9 2
13 3 2 1 15 9 2 15 4 13 9 14 13 2
23 11 13 10 0 9 16 13 12 9 2 12 9 7 12 9 1 15 0 12 2 9 9 2
21 1 10 9 2 3 2 15 4 13 0 9 1 10 9 14 13 12 9 1 9 2
12 1 15 9 2 11 13 0 9 1 10 9 2
32 10 12 9 13 11 2 3 13 1 1 10 0 9 9 9 9 2 7 13 2 10 0 9 15 15 9 13 1 1 9 2 2
31 10 12 9 13 11 2 10 3 0 0 9 7 9 2 15 2 3 13 9 9 1 10 9 14 13 15 9 3 3 2 2
16 7 10 12 9 13 11 2 10 0 9 9 9 7 9 2 2
36 3 2 15 13 3 0 16 9 9 13 11 14 9 2 1 10 11 11 7 10 11 11 11 2 1 11 7 1 0 9 2 4 13 3 3 2
20 11 13 3 0 1 9 1 11 11 14 9 1 10 9 11 11 11 1 11 2
30 7 2 16 15 13 1 11 2 15 13 0 14 13 1 10 9 14 0 9 2 13 15 0 9 2 7 9 1 15 2
15 9 13 3 0 14 13 16 15 13 0 7 14 1 11 2
38 10 11 9 13 11 1 10 11 11 11 14 9 2 7 9 15 4 13 0 9 13 1 10 11 13 10 9 16 15 4 13 15 3 1 15 0 9 2
25 7 15 4 4 13 1 9 16 11 4 3 13 11 14 9 2 16 11 4 14 3 13 11 14 2
41 1 11 2 16 10 11 11 11 4 13 10 9 2 11 13 11 2 13 3 14 13 1 11 1 7 3 2 7 13 10 9 2 16 1 15 13 1 1 9 2 2
24 3 2 11 13 2 2 3 16 15 13 10 0 9 4 14 2 1 9 2 13 10 9 2 2
15 3 2 1 10 11 11 9 2 10 9 4 13 1 11 2
4 15 13 0 2
9 15 4 13 3 0 16 15 4 2
14 7 3 9 11 4 13 0 1 15 0 9 3 3 2
11 11 11 13 10 11 11 9 1 11 11 2
9 15 9 13 1 10 11 10 9 2
19 12 9 1 9 9 7 10 0 9 1 10 9 13 0 2 7 3 0 2
17 15 13 10 9 1 11 4 13 16 16 10 9 4 13 10 9 2
42 15 13 10 9 16 0 11 13 10 9 1 12 11 1 10 9 1 13 9 2 12 15 4 4 13 10 15 9 2 7 1 10 0 9 2 0 9 4 3 13 15 2
39 10 0 9 4 13 9 9 10 4 13 10 9 1 10 9 1 9 2 7 15 13 14 13 3 15 4 13 0 14 13 10 12 2 7 3 2 9 9 2
14 0 9 9 4 3 4 3 13 7 13 1 0 9 2
28 3 16 10 9 13 0 2 10 12 0 13 9 13 14 13 10 11 11 11 9 7 11 14 11 2 11 9 2
21 11 11 2 7 0 9 13 1 15 9 2 4 3 3 13 15 0 9 1 9 2
30 12 9 3 13 1 12 9 2 9 2 1 9 13 10 9 9 1 11 2 10 9 10 13 3 0 9 1 0 11 2
26 11 11 11 2 11 2 10 9 1 11 2 13 10 9 16 10 11 11 4 13 10 11 11 11 9 2
36 3 2 11 14 9 3 1 10 9 4 13 3 0 16 13 0 11 1 10 9 1 9 2 10 4 13 1 10 9 1 3 3 12 1 15 2
39 11 2 11 13 16 2 15 11 2 13 14 3 13 10 9 16 2 9 2 2 3 10 9 1 11 2 4 4 13 0 9 9 7 9 9 1 15 9 2
21 3 15 13 10 0 13 9 1 11 14 9 13 10 9 2 10 15 13 13 0 2
22 11 11 2 11 7 9 9 11 11 2 11 4 4 13 1 0 0 9 1 10 9 2
46 11 13 11 1 10 2 11 2 7 10 2 0 0 9 1 11 7 10 11 2 2 16 11 13 11 1 10 2 9 2 7 10 2 0 9 15 13 1 15 0 9 16 13 11 2 2
35 12 9 13 1 11 1 11 2 11 11 2 16 15 4 14 13 0 1 11 16 15 4 13 15 7 10 9 3 13 15 13 1 10 9 2
27 15 13 10 3 0 9 2 13 11 13 0 7 0 2 13 1 11 2 3 0 7 3 13 15 16 13 2
4 9 2 6 2
50 11 11 2 11 2 1 10 9 2 13 10 9 1 10 0 11 1 11 2 11 1 11 7 13 10 9 14 13 0 9 9 2 11 11 2 11 2 1 15 0 9 9 2 10 4 4 13 1 9 2
18 10 0 0 9 9 2 11 7 11 2 4 3 13 1 10 0 9 2
24 3 3 2 0 11 13 7 13 16 16 15 4 13 14 13 10 9 14 13 15 1 1 9 2
9 15 13 15 4 13 10 9 3 2
34 0 11 2 13 0 7 0 11 2 4 3 13 1 10 11 11 11 2 3 1 10 9 14 13 10 9 1 11 1 10 0 11 11 2
27 10 11 11 13 10 0 9 1 13 9 9 1 10 9 7 4 4 13 1 10 0 0 0 9 1 11 2
11 15 9 9 13 3 0 16 15 15 13 2
1 2
29 0 9 4 13 7 13 10 0 12 9 2 9 4 4 13 1 9 14 13 7 14 13 10 9 1 10 11 11 2
22 0 9 13 1 15 0 1 11 2 12 2 16 0 13 3 3 13 11 7 0 9 2
28 15 13 10 0 9 1 10 0 2 0 9 9 15 13 14 13 1 11 7 13 3 1 9 1 11 2 11 2
48 16 13 15 10 9 15 13 1 2 3 13 15 0 9 2 15 13 13 9 1 10 11 2 13 15 11 2 11 2 9 9 2 2 0 9 7 10 9 1 0 9 10 15 4 14 13 3 2
25 15 13 11 14 9 1 15 1 10 13 9 7 15 13 10 0 9 1 10 9 1 9 7 9 2
22 15 4 14 13 1 15 7 15 13 15 15 15 13 4 13 10 0 9 1 10 9 2
10 15 13 16 9 13 10 0 0 9 2
19 3 13 1 10 11 2 3 13 10 11 3 1 9 2 1 1 12 2 2
12 0 11 13 16 9 13 0 14 13 1 9 2
49 13 3 10 9 16 10 9 13 1 0 0 9 1 10 9 2 11 4 3 13 10 0 9 2 10 3 13 15 14 13 16 10 9 13 1 10 0 9 9 3 13 3 15 15 4 13 14 13 2
39 15 13 10 9 10 9 3 1 10 13 11 0 2 9 15 13 16 11 13 10 9 14 13 10 0 9 9 7 13 1 9 1 12 9 1 10 0 9 2
46 16 13 15 9 1 15 9 15 13 16 11 9 13 1 10 9 1 10 9 7 16 15 4 13 10 0 9 2 3 16 0 4 13 0 9 2 3 1 0 9 2 1 15 0 9 2
21 15 13 16 15 13 10 9 7 10 9 3 3 1 10 9 1 13 7 0 9 2
37 15 13 16 11 7 0 9 9 13 0 16 3 13 3 3 12 1 1 12 9 2 1 1 10 9 2 16 11 13 14 4 13 1 10 9 3 2
29 7 15 3 13 15 1 10 0 9 2 10 4 13 11 9 2 16 15 4 14 13 10 11 4 13 3 3 3 2
66 10 9 10 13 9 1 10 9 3 13 15 2 3 3 3 11 4 13 14 13 10 11 14 13 15 9 2 16 15 15 4 13 3 2 14 16 15 4 13 10 9 13 1 1 10 9 2 7 16 15 13 10 0 0 9 2 1 10 9 11 2 14 13 15 1 2
27 10 0 9 3 13 16 2 13 10 9 2 10 11 11 4 13 10 9 1 9 7 9 1 10 13 9 2
41 15 4 13 13 1 0 9 1 1 9 2 16 15 13 10 0 9 1 15 9 7 4 3 13 1 10 11 1 15 9 1 9 1 10 9 16 13 9 7 9 2
15 0 1 10 9 4 4 13 7 13 1 10 0 12 9 2
38 3 3 2 11 9 1 11 2 11 13 10 0 9 16 3 13 11 2 11 11 11 2 11 2 11 1 10 11 2 11 11 9 1 10 0 11 9 2
15 11 2 11 4 13 9 7 13 1 0 9 1 10 9 2
19 10 11 9 3 13 14 4 13 10 9 1 11 2 11 9 10 9 3 2
38 10 11 2 11 11 1 11 7 11 2 11 13 1 9 1 11 1 10 9 13 10 9 1 11 11 11 2 11 2 10 11 11 9 13 1 15 9 2
13 10 9 13 12 9 14 4 13 1 10 11 11 2
36 10 0 9 13 10 0 9 1 11 11 11 2 11 2 1 10 11 9 10 4 13 1 10 9 1 11 2 11 2 11 7 11 11 2 11 2
18 11 2 11 4 13 1 9 7 4 3 13 14 4 13 13 10 9 2
15 15 13 0 9 14 13 10 0 9 3 1 10 0 11 2
13 10 11 4 14 13 1 10 11 2 7 3 3 2
24 10 4 13 10 9 1 10 0 12 9 7 15 13 10 0 9 3 12 4 13 1 10 0 2
16 3 9 13 14 10 9 2 15 13 10 0 9 1 10 12 2
5 13 11 11 11 2
22 3 13 10 11 11 9 1 10 0 9 7 0 11 9 1 10 9 9 2 13 9 2
9 2 2 3 3 15 13 10 9 2
10 15 13 10 11 9 4 13 1 15 2
9 3 15 13 10 9 3 2 2 2
15 1 1 0 9 2 11 4 4 13 1 9 1 9 9 2
10 15 4 14 13 15 13 14 13 15 2
17 9 4 3 4 13 0 13 9 1 11 14 9 1 10 0 9 2
19 3 3 1 0 9 10 0 9 13 15 13 10 9 15 4 13 10 9 2
20 7 0 1 10 9 2 11 13 15 9 7 13 15 0 9 2 10 11 9 2
23 7 16 15 4 13 10 0 9 2 15 13 14 10 10 9 16 15 4 13 3 1 15 2
23 15 4 4 13 10 9 1 10 9 10 0 0 2 0 9 13 13 2 11 9 11 11 2
55 11 4 4 13 10 0 9 1 15 9 9 16 11 13 10 0 0 9 15 13 13 15 0 9 1 10 11 2 16 2 16 15 13 15 1 10 9 2 15 4 13 15 9 3 2 7 15 4 13 1 15 15 13 2 2
18 7 3 2 3 15 4 14 4 13 15 3 2 16 11 13 14 11 2
11 11 4 4 13 1 2 7 11 4 14 2
20 11 14 9 13 0 2 7 13 10 0 9 10 13 10 2 9 1 9 2 2
30 15 13 1 10 11 10 2 1 11 2 13 10 0 7 0 9 1 10 9 10 9 9 7 9 9 13 1 10 0 2
9 2 13 11 11 1 10 11 2 2
27 10 9 13 11 2 7 13 0 9 10 10 11 9 7 15 9 13 10 9 1 10 0 9 13 14 13 2
26 11 14 9 2 1 10 0 9 2 4 13 1 0 9 2 3 1 10 9 15 4 14 13 15 9 2
15 7 1 15 15 4 14 3 13 15 9 2 14 3 10 2
7 7 4 11 4 13 1 2
23 15 13 15 4 4 13 1 11 2 10 13 10 0 9 10 9 4 4 13 1 10 9 2
25 15 13 15 4 4 13 16 2 1 2 0 9 2 11 11 2 11 4 14 4 13 10 0 9 2
20 10 9 4 13 16 11 4 3 4 13 1 10 0 11 2 0 9 1 11 2
20 16 10 10 9 4 13 7 13 4 13 10 9 2 9 4 14 4 13 3 2
20 7 11 13 3 12 9 0 2 7 10 0 9 4 13 15 13 10 0 9 2
12 3 3 11 4 4 13 3 2 1 0 9 2
25 10 9 1 10 11 3 2 3 14 3 0 16 13 10 0 9 13 1 11 2 13 1 15 9 2
7 11 13 0 1 10 9 2
14 15 9 13 10 9 9 1 10 2 9 1 9 2 2
7 3 15 9 4 13 0 2
26 10 9 1 0 9 7 9 13 2 13 1 10 9 2 4 13 1 10 9 11 11 2 1 11 11 2
27 11 2 10 11 9 3 13 1 10 11 9 2 13 10 9 13 14 13 15 1 10 0 9 1 11 11 2
11 15 13 14 13 10 9 13 14 13 9 2
1 8
74 15 4 13 10 9 2 15 13 10 0 9 9 1 10 9 1 9 2 3 16 3 0 1 10 0 9 4 13 10 9 1 11 9 9 10 13 16 11 13 10 9 1 9 1 10 11 9 9 10 13 9 1 10 11 9 2 13 1 0 9 9 13 11 11 2 11 11 2 11 11 7 11 11 2
21 11 11 11 13 10 9 16 3 11 14 9 4 13 1 15 1 15 9 11 11 2
7 2 0 0 2 0 0 2
34 1 16 10 9 1 10 12 9 13 16 10 11 9 4 14 13 13 10 9 2 3 13 15 1 9 1 11 2 10 9 13 10 9 2
23 15 13 9 10 4 13 10 9 15 4 13 0 14 13 10 0 9 1 11 9 1 11 2
21 11 4 13 16 15 4 4 13 1 10 11 3 15 13 10 9 2 12 1 11 2
26 10 9 4 13 15 13 10 9 13 15 9 1 0 9 1 7 11 7 10 2 11 1 11 11 2 2
34 11 4 13 0 14 13 16 15 4 13 0 1 12 2 0 9 2 1 10 11 1 15 9 1 12 2 13 10 9 14 9 1 9 2
9 3 11 11 11 13 1 10 9 2
65 3 13 11 9 2 11 13 10 9 1 11 9 2 12 2 16 1 11 9 2 12 2 15 4 13 10 9 1 11 9 2 1 10 0 10 1 10 9 13 1 11 11 11 2 7 10 0 9 13 15 9 1 11 9 2 12 2 3 15 13 1 10 11 2 2
26 10 11 11 13 16 1 12 9 1 12 2 11 4 14 13 2 3 7 3 2 1 10 11 16 13 2
1 8
23 0 9 2 11 11 11 11 11 1 11 2 11 2 13 1 11 14 12 2 9 0 9 2
23 11 11 13 2 2 9 3 13 0 9 1 15 2 2 13 2 9 13 3 1 9 2 2
1 8
1 8
11 13 16 15 4 13 15 9 3 1 11 2
10 0 9 2 9 13 1 9 9 9 9
4 11 2 11 2
34 9 14 9 1 11 13 10 0 9 11 1 10 0 9 1 10 9 13 9 1 0 9 1 9 7 9 1 10 11 2 11 2 9 2
24 11 11 11 11 2 12 2 4 13 1 10 9 1 13 9 1 10 9 1 10 9 1 12 2
35 9 13 11 13 1 9 16 15 13 9 1 10 0 9 1 11 12 7 13 16 13 1 0 9 13 9 7 10 9 10 13 1 11 11 2
28 11 11 9 14 9 11 11 11 2 12 2 4 13 11 1 12 9 1 13 9 7 12 9 1 9 1 9 2
60 1 11 2 11 11 2 12 2 10 0 9 1 11 11 2 4 13 1 12 9 1 13 9 7 12 9 1 9 1 9 16 15 13 1 1 10 11 11 11 14 11 7 13 15 4 13 9 1 10 9 1 10 9 10 3 13 12 9 3 2
25 15 13 10 0 9 13 3 3 1 10 9 1 10 9 1 10 9 7 0 9 13 1 10 9 2
16 16 15 13 11 15 4 13 11 1 11 14 13 9 1 3 2
6 6 2 2 9 2 2
22 9 9 2 10 11 9 4 13 1 10 0 9 9 9 1 11 2 11 2 11 2 2
15 10 3 13 9 2 13 15 0 1 10 9 9 2 4 13
1 11
10 3 15 13 10 9 15 4 13 1 2
12 15 3 13 15 13 2 15 13 13 10 9 2
21 15 4 14 13 3 9 13 2 7 15 4 3 13 1 9 1 11 1 10 9 2
14 10 0 0 11 1 11 13 14 15 15 13 14 13 2
5 15 13 15 9 2
11 6 13 1 15 15 13 10 9 1 9 2
17 6 15 13 10 0 9 2 15 3 13 10 9 1 11 11 0 9
10 15 4 13 15 1 2 11 11 0 9
6 15 13 10 0 9 2
4 13 15 13 2
15 15 4 13 1 9 1 15 15 13 10 0 0 9 9 2
7 15 3 3 13 9 9 2
8 15 4 13 0 14 13 3 2
7 6 15 3 13 15 9 2
10 15 3 13 10 9 9 9 5 9 2
6 15 3 13 1 9 9
12 6 13 7 13 15 1 16 15 13 10 9 2
12 15 4 13 1 9 9 9 7 13 10 9 2
4 15 13 3 2
1 11
31 3 4 15 13 14 13 3 15 4 13 1 10 0 0 9 10 4 9 2 13 1 15 9 2 7 1 10 9 1 15 2
5 15 4 13 15 2
13 7 15 13 14 0 14 13 2 16 15 13 3 2
14 4 14 13 15 13 15 3 16 3 3 13 10 9 2
28 10 0 9 13 16 15 13 14 13 10 9 1 5 12 2 7 2 15 13 14 13 10 0 9 13 1 15 2
1 8
20 5 16 10 9 1 10 11 11 9 13 3 2 0 9 4 3 13 1 9 2
10 1 0 9 2 15 9 4 13 0 2
60 10 9 14 13 1 9 10 9 9 1 10 0 0 9 7 0 0 0 9 11 11 11 0 11 12 1 10 0 9 1 11 2 7 10 0 2 9 2 1 0 11 11 13 15 9 7 13 10 0 0 9 2 13 0 9 1 9 9 2 5
5 9 1 11 14 9
2 11 11
30 1 0 11 2 11 13 12 0 9 1 11 16 13 1 10 11 11 2 9 1 10 11 11 9 2 13 9 9 2 2
26 10 0 9 1 10 11 11 2 10 0 9 1 10 11 11 11 1 11 2 4 4 13 1 0 9 2
16 15 13 0 2 7 3 0 2 16 15 4 4 13 1 11 2
31 7 10 9 1 10 0 9 13 3 10 9 1 10 9 3 15 13 1 13 9 1 11 11 1 10 9 1 10 11 11 2
19 9 4 13 1 10 9 9 16 10 11 11 13 14 3 0 1 11 9 2
27 15 4 3 13 10 9 9 1 10 11 11 1 11 11 2 11 2 2 15 13 3 3 1 10 11 11 2
23 9 13 1 10 9 13 1 9 1 10 11 12 9 2 10 13 10 0 9 1 10 11 2
42 9 15 13 3 14 13 10 9 13 15 3 13 10 9 2 10 0 9 9 13 10 0 9 14 11 11 11 11 2 3 4 13 1 1 11 14 2 0 9 9 2 2
2 13 9
50 9 9 1 10 11 11 13 14 0 2 7 15 4 13 1 10 0 0 9 2 1 9 1 10 9 1 10 9 9 1 11 2 11 7 11 2 7 3 1 10 0 0 9 1 11 2 11 7 11 2
68 16 10 0 9 4 13 9 2 0 1 10 0 9 2 7 4 13 10 9 16 13 10 0 9 1 10 9 2 15 4 13 3 0 1 15 0 9 2 3 15 9 13 14 10 0 9 7 10 9 1 0 2 0 7 9 2 13 9 13 1 11 11 7 0 11 1 11 2
31 10 11 11 13 10 0 9 1 10 9 2 7 10 12 0 7 0 9 10 13 10 11 7 11 9 13 10 0 9 9 2
9 10 9 7 9 13 1 10 9 2
53 16 10 2 11 11 2 1 10 11 2 3 13 1 10 11 11 2 13 10 9 15 13 10 11 11 2 15 13 10 9 7 9 1 15 0 9 7 3 14 13 1 9 1 11 7 3 1 10 0 9 1 11 2
17 15 13 0 9 16 10 11 11 4 13 10 0 9 1 11 11 2
8 15 13 14 0 1 11 11 2
62 10 0 9 1 10 9 1 11 11 2 1 10 11 2 13 10 0 9 13 16 9 1 11 2 11 7 11 11 4 3 13 1 10 9 2 13 0 0 9 9 2 16 9 1 11 2 11 2 11 7 11 4 13 3 14 13 10 0 9 7 13 2
30 2 11 11 2 11 11 2 11 2 11 11 2 11 14 11 2 11 11 7 11 4 3 13 1 9 2 2 15 13 2
27 10 0 9 13 1 12 13 15 13 12 2 9 2 1 10 11 11 2 7 0 9 13 3 0 1 15 2
24 10 0 9 1 15 13 11 2 15 1 9 1 15 9 4 13 15 3 13 9 14 13 3 2
30 16 0 1 15 13 0 0 9 2 7 10 11 13 0 9 1 15 1 10 9 2 15 13 1 9 7 0 0 9 2
21 10 9 1 10 11 11 1 10 9 1 9 2 9 7 9 13 10 9 3 0 2
39 9 1 11 11 13 15 0 16 11 11 13 0 1 2 10 2 9 9 2 7 10 0 11 11 13 3 0 14 13 1 10 9 1 0 9 1 10 9 2
21 12 0 0 9 4 13 13 2 2 9 9 13 10 3 0 9 1 10 9 2 2
18 13 10 9 14 0 0 9 2 15 13 0 3 0 11 11 4 13 2
35 10 9 13 1 10 0 9 9 1 10 11 1 11 2 1 10 12 9 7 9 9 13 3 2 13 3 9 1 10 11 11 7 11 11 2
2 9 9
19 16 10 9 1 10 11 11 9 13 3 2 0 9 4 3 13 1 9 2
10 1 0 9 2 15 9 4 13 0 2
59 10 9 14 13 1 9 10 9 9 1 10 0 0 9 7 0 0 0 9 11 11 11 0 11 12 1 10 0 9 1 11 2 7 10 0 2 9 2 1 0 11 11 13 15 9 7 13 10 0 0 9 2 13 0 9 1 9 9 2
23 1 13 0 7 0 9 2 11 4 13 0 1 0 9 1 10 9 3 14 13 0 9 2
36 16 11 11 13 3 16 13 9 1 15 0 9 1 9 2 9 2 9 9 7 9 9 2 15 4 14 13 0 9 1 10 9 1 13 9 2
40 1 9 2 15 4 13 14 13 3 0 0 9 2 0 1 10 0 8 11 11 2 11 2 7 3 2 13 11 2 14 13 10 9 7 13 11 14 0 9 2
13 0 9 14 0 9 16 13 1 10 11 13 0 2
32 10 0 9 2 10 13 10 0 9 10 0 9 1 10 9 2 4 4 13 1 0 11 7 1 10 11 11 1 10 0 9 2
36 1 12 2 13 1 0 9 9 2 9 9 13 10 3 2 13 9 1 10 12 2 10 13 9 13 11 7 11 2 7 13 0 9 1 9 2
16 10 9 4 13 14 13 1 10 11 7 2 0 9 9 2 2
20 10 13 2 7 2 13 9 4 13 1 1 10 0 9 1 13 9 1 11 2
16 1 9 2 11 9 1 10 11 11 13 3 0 1 0 9 2
16 10 0 11 0 9 4 13 1 10 3 2 0 11 1 12 2
41 10 9 1 9 2 9 7 9 2 13 14 4 4 13 1 11 7 0 0 12 9 2 13 10 9 1 11 1 11 1 0 11 12 1 10 9 11 2 11 12 2
16 16 13 11 0 9 2 10 9 13 15 9 1 9 1 11 2
43 1 15 9 1 10 11 1 11 10 9 4 13 1 10 0 9 7 11 2 13 9 9 1 11 14 11 11 11 2 15 4 13 1 0 0 9 1 11 11 14 0 9 2
4 11 9 2 9
36 1 12 2 10 0 9 13 10 9 1 10 12 2 9 9 1 10 9 1 10 0 9 1 11 2 7 10 9 1 12 9 1 9 7 9 2
30 1 10 9 13 13 12 9 2 13 2 9 9 2 12 9 9 2 9 2 12 9 9 7 0 1 12 9 1 9 2
15 12 9 4 13 2 3 13 1 10 11 11 11 14 11 2
11 12 9 9 13 1 10 11 9 1 11 2
11 10 9 4 13 1 11 14 11 1 11 2
24 1 12 10 11 13 10 9 1 11 2 10 9 1 10 9 1 11 2 3 1 10 11 9 2
11 3 2 11 13 10 11 14 0 9 9 2
24 10 11 11 2 13 11 1 10 0 9 4 13 1 0 9 1 12 1 15 9 1 10 11 2
34 1 10 9 1 15 9 2 10 9 13 3 0 16 13 10 2 9 2 1 10 9 1 10 9 1 11 1 11 1 10 11 11 9 2
2 0 9
32 10 0 9 1 10 11 9 13 10 0 9 2 9 1 9 7 9 10 13 10 11 11 7 10 9 1 3 2 0 0 9 2
15 1 10 0 9 2 11 4 3 13 1 10 9 1 9 2
27 10 9 1 9 9 2 1 10 9 1 10 11 9 2 4 13 0 1 9 9 2 9 9 7 0 9 2
55 15 4 3 13 16 10 0 11 4 13 10 9 1 9 11 9 2 0 1 10 11 2 11 2 11 2 11 2 11 2 1 10 9 9 1 11 2 7 13 10 9 1 9 9 1 11 14 9 1 9 1 10 9 9 2
28 1 10 9 2 3 1 10 11 11 2 0 9 9 4 13 10 9 1 9 0 1 10 9 1 9 7 9 2
34 10 9 1 9 7 9 13 16 9 4 13 1 10 11 1 11 2 11 7 11 1 11 2 1 3 15 4 13 3 1 9 1 11 2
24 10 9 1 11 1 11 1 11 14 11 13 1 0 11 2 11 7 11 2 7 3 1 11 2
1 9
24 11 14 11 7 11 11 13 0 1 12 9 13 12 9 3 1 11 11 1 10 11 1 11 2
22 13 12 9 1 9 1 9 2 15 13 1 1 10 9 1 11 3 1 11 1 11 2
30 10 11 11 11 13 10 11 2 10 13 10 0 7 3 3 13 0 9 2 1 10 12 7 3 11 11 1 10 9 2
28 1 11 11 2 10 3 3 13 9 2 13 11 11 2 10 13 10 9 7 10 3 0 9 1 10 0 9 2
24 9 1 10 11 11 13 0 1 11 2 7 15 4 3 14 13 1 10 9 1 11 11 11 2
30 11 11 13 1 10 9 1 0 9 7 13 10 0 9 1 10 11 2 13 11 7 10 11 11 2 13 11 11 11 2
14 15 3 13 1 11 2 11 14 9 2 13 0 9 2
18 2 11 3 13 14 13 1 10 13 1 9 1 11 7 11 1 11 2
23 11 13 11 11 16 13 15 9 1 11 7 11 14 13 0 9 15 13 0 1 0 11 2
20 0 9 13 15 13 3 0 1 12 11 9 13 1 11 7 10 12 1 11 2
19 2 15 13 10 9 13 3 16 15 4 13 11 2 2 13 10 0 9 2
8 7 11 7 11 13 10 9 2
40 2 4 11 13 15 10 9 1 10 0 9 13 0 9 14 13 1 15 9 15 4 13 15 3 3 2 2 13 11 11 10 9 1 11 14 11 11 11 2 2
6 11 2 11 0 0 9
2 11 2
33 1 10 0 12 9 0 11 4 13 1 0 9 1 15 9 2 11 2 11 7 10 0 0 9 2 7 0 9 2 11 7 11 2
26 10 9 4 3 13 2 7 15 13 9 16 1 16 13 11 14 9 15 4 3 4 13 14 13 15 2
24 2 10 9 4 13 10 9 1 10 15 9 16 10 0 11 2 10 0 11 13 0 1 10 2
20 9 4 13 10 9 1 11 2 2 11 11 11 13 11 14 11 9 10 11 2
30 2 10 0 9 4 3 13 10 11 9 7 13 10 0 9 2 7 0 9 13 16 15 10 13 15 0 9 1 11 2
55 1 11 12 2 11 4 4 3 13 1 0 7 0 9 16 13 11 9 15 4 13 14 13 10 9 2 7 1 10 0 9 10 11 4 13 13 11 11 11 1 10 9 16 15 4 13 10 11 13 11 11 9 1 11 2
31 15 13 1 11 12 3 11 11 11 11 2 11 7 11 13 10 12 9 9 1 11 11 1 10 9 1 10 11 11 11 2
33 10 9 4 13 3 1 10 11 7 10 11 11 11 15 13 3 0 14 13 10 0 9 1 11 7 10 9 1 0 0 13 11 2
28 0 7 0 9 3 0 1 10 9 2 13 11 13 11 3 16 13 1 10 11 16 10 9 4 13 9 3 2
13 2 3 13 11 11 2 11 11 7 11 11 2 2
10 11 4 13 14 4 13 10 0 11 2
16 10 12 13 9 11 7 15 9 7 13 14 4 13 1 11 2
40 2 11 11 13 9 1 10 11 2 11 13 10 0 9 9 1 11 1 10 11 9 7 3 10 9 1 11 9 16 11 13 10 9 11 2 11 2 11 2 2
28 2 15 13 10 0 9 3 11 3 13 1 10 11 9 1 1 11 11 1 10 11 2 2 13 10 0 9 2
15 2 11 4 3 3 13 1 10 9 2 2 10 9 13 2
28 10 0 9 1 10 9 13 2 2 10 11 3 13 16 10 11 13 10 0 9 1 15 9 1 11 11 2 2
8 11 13 3 0 1 10 9 2
23 2 11 11 13 14 13 15 7 13 1 15 16 13 0 9 1 10 11 2 2 13 11 2
25 10 0 9 10 0 11 3 13 16 11 4 14 13 0 9 1 11 2 10 0 9 1 10 11 2
11 1 3 15 4 13 11 14 9 13 0 2
14 3 0 9 13 16 10 9 13 0 1 10 0 9 2
38 11 7 11 0 9 1 11 13 15 13 3 0 14 13 16 11 14 0 9 13 0 16 13 11 7 10 11 14 13 10 11 14 13 16 13 10 9 2
13 3 15 13 0 9 1 10 9 1 10 11 9 2
23 2 11 3 13 10 0 9 13 1 11 10 13 14 3 3 2 2 13 11 11 11 11 2
32 2 15 13 3 0 0 9 1 15 9 1 10 9 1 10 9 2 7 10 9 1 11 3 13 1 10 9 2 2 15 13 2
28 3 0 9 1 10 9 11 13 10 9 9 9 1 11 1 11 10 13 10 0 9 9 1 10 11 1 11 2
38 3 11 0 9 13 0 9 9 2 0 1 15 0 2 13 9 1 10 11 11 15 13 1 10 9 13 3 0 1 10 11 7 10 9 1 10 11 2
26 1 10 0 9 10 11 13 0 1 10 0 9 7 0 9 10 10 9 4 13 1 15 9 1 11 2
42 3 3 4 10 9 13 0 0 9 2 13 9 7 0 9 1 10 0 9 7 15 4 3 13 0 9 2 1 12 5 12 0 9 4 4 13 1 10 9 1 11 2
19 11 4 3 13 16 10 11 4 3 13 0 9 1 11 9 13 1 11 2
5 15 3 4 13 2
21 11 7 0 9 4 3 4 13 10 11 1 10 9 1 11 9 7 15 13 9 2
37 3 15 13 3 0 0 9 1 9 14 13 7 13 3 1 11 13 11 9 2 15 4 4 13 3 1 11 7 4 13 10 9 1 10 11 9 2
26 1 10 11 9 14 13 10 0 9 2 10 9 13 3 3 0 1 10 0 11 15 13 14 13 3 2
29 1 3 11 4 14 13 10 10 9 7 3 15 4 14 13 16 15 13 7 10 9 1 11 7 10 9 1 11 2
48 1 11 11 0 14 13 10 9 7 10 9 1 0 0 11 11 9 0 1 11 11 7 9 11 11 2 15 13 3 0 9 16 0 11 9 14 13 9 1 0 11 11 9 16 15 13 3 2
17 15 9 4 3 13 13 9 16 11 14 13 10 9 1 0 11 2
19 0 9 13 10 9 1 11 12 1 11 11 11 11 1 10 0 11 9 2
36 11 4 3 13 7 13 1 11 16 1 10 0 9 15 13 10 0 9 1 10 0 0 9 1 10 0 7 11 9 1 9 0 1 9 9 2
17 11 3 13 14 13 1 10 13 1 9 1 11 7 11 1 11 2
23 11 13 11 11 16 13 15 9 1 11 7 11 14 13 0 9 15 13 0 1 0 11 2
20 0 9 13 15 13 3 0 1 12 11 9 13 1 11 7 10 12 1 11 2
19 2 15 13 10 9 13 3 16 15 4 13 11 2 2 13 10 0 9 2
8 7 11 7 11 13 10 9 2
39 2 4 11 13 15 10 9 1 10 0 9 13 0 9 14 13 1 15 9 15 4 13 15 3 3 2 2 13 11 11 10 9 1 11 14 11 11 11 2
27 11 3 13 16 15 4 13 11 3 16 10 0 9 1 11 13 1 0 9 1 11 4 4 13 1 3 2
11 0 11 9 7 0 9 4 13 11 3 2
52 1 10 0 0 9 13 10 3 13 9 1 11 2 11 2 11 7 11 10 4 3 13 10 11 13 0 11 11 13 0 9 14 13 0 9 11 11 14 13 10 9 1 11 1 10 9 7 14 14 13 11 2
17 11 1 0 13 16 11 4 13 7 3 4 3 13 1 10 9 2
19 11 13 14 13 10 0 9 16 15 0 0 11 13 15 14 13 1 11 2
33 3 1 10 9 0 9 4 13 0 16 13 10 11 11 9 11 11 14 13 10 9 1 10 9 7 3 13 11 14 13 10 0 2
37 16 10 11 0 9 13 10 9 1 15 9 1 7 11 7 11 2 11 14 0 9 13 0 14 13 13 11 16 16 10 11 9 1 11 4 13 2
26 3 0 9 1 11 4 4 13 14 13 10 9 7 10 0 9 13 0 14 13 10 9 1 10 9 2
26 0 9 13 3 0 1 10 11 9 1 11 2 10 0 11 2 9 9 3 12 9 1 11 14 9 2
37 10 13 11 9 1 0 11 4 3 13 0 1 10 9 1 11 11 2 10 9 7 11 1 11 9 0 9 2 15 13 10 0 9 1 0 9 2
22 0 9 13 15 13 10 9 1 11 14 9 16 15 13 14 13 11 14 9 1 9 2
61 1 10 9 1 13 9 1 11 7 11 1 11 14 0 9 9 7 9 1 9 1 11 16 10 0 11 9 4 13 1 11 3 2 10 11 13 16 11 4 4 13 1 10 9 9 2 9 9 7 3 10 9 9 1 10 0 11 9 1 11 2
16 0 9 13 10 11 4 13 3 12 0 9 7 9 1 11 2
13 3 11 11 13 10 11 9 13 10 9 1 11 2
20 2 15 13 10 3 0 9 1 9 1 11 1 10 0 9 2 2 13 11 2
24 3 15 13 11 1 10 0 7 0 9 16 15 13 14 13 0 9 1 7 10 11 7 11 2
15 2 11 4 13 10 9 1 9 1 7 10 11 7 11 2
27 3 3 15 15 4 13 3 4 13 0 1 15 7 15 13 3 15 4 13 14 13 15 2 2 13 11 2
31 9 4 13 16 10 9 1 11 14 9 13 3 2 7 10 9 4 13 0 14 13 11 7 13 3 3 1 9 14 9 2
27 1 10 8 0 9 15 4 13 3 0 16 10 11 4 14 13 10 9 1 10 0 9 7 10 0 11 2
33 1 10 3 0 9 0 0 9 1 10 11 9 13 10 11 1 11 7 11 16 16 15 13 7 13 10 9 2 15 4 4 13 2
10 0 11 13 1 11 13 1 11 11 2
46 15 13 3 3 0 16 1 10 3 13 9 1 11 2 10 9 1 0 11 11 9 7 10 0 0 9 1 11 2 11 4 13 15 9 16 13 0 9 1 11 9 13 1 0 9 2
3 11 11 12
28 10 9 10 10 9 1 11 9 0 1 10 11 9 4 3 13 1 11 11 14 9 9 13 0 1 10 9 2
27 10 9 10 15 4 13 10 9 1 16 13 1 11 13 0 7 4 4 13 1 10 0 9 14 13 0 2
15 0 1 15 13 10 9 4 3 13 2 13 2 13 15 2
10 7 15 13 14 9 7 4 3 13 2
17 7 14 13 10 9 1 10 0 9 13 14 13 13 1 15 9 2
30 10 0 9 1 10 0 9 4 3 13 3 15 13 16 11 11 11 3 13 10 9 3 3 1 10 9 1 15 9 2
9 15 4 3 13 1 10 9 9 2
15 16 10 1 11 11 14 9 13 0 2 11 13 10 9 2
50 2 7 2 10 9 1 9 1 10 9 10 13 3 10 0 9 4 4 13 4 15 13 10 9 7 13 1 10 9 2 10 9 13 1 15 9 13 15 13 1 0 9 7 4 14 13 15 1 15 2
9 15 13 10 9 1 10 9 2 2
10 11 13 10 9 14 9 16 1 9 2
6 11 13 10 0 9 2
8 15 4 11 13 1 15 9 2
4 15 4 13 2
15 15 4 13 1 10 9 2 10 9 2 1 10 0 9 2
3 1 9 2
18 15 13 10 9 1 9 2 13 9 2 7 4 14 3 13 1 3 2
41 10 9 1 9 7 3 0 9 9 13 10 0 9 16 15 3 3 13 1 11 14 9 1 10 0 9 2 7 4 13 15 9 1 15 0 7 0 9 1 9 2
41 15 0 9 3 13 10 0 9 1 11 0 9 2 13 12 11 2 0 1 15 9 7 9 2 1 9 1 10 9 1 12 0 9 2 12 1 15 10 11 11 2
16 2 11 13 16 11 13 15 9 2 2 13 9 13 2 2 2
7 10 9 13 3 12 9 2
6 11 13 10 0 9 2
10 15 3 13 2 1 9 2 13 9 2
33 15 9 16 13 9 13 10 9 9 1 12 3 15 13 2 1 12 9 2 14 13 10 9 16 13 0 2 9 10 0 3 3 2
15 15 4 3 13 1 13 13 9 1 10 0 9 1 11 2
16 9 9 4 13 10 9 1 10 9 14 13 0 9 1 9 2
18 12 9 16 13 15 0 9 1 0 3 0 9 4 13 11 13 9 2
31 3 1 15 15 3 13 2 2 0 2 0 9 2 9 2 9 9 2 7 0 2 9 9 2 13 10 0 14 13 2 2
23 16 15 13 14 13 1 10 9 2 16 1 10 9 9 2 15 13 3 3 2 13 0 2
31 7 15 13 10 0 9 1 10 9 2 7 15 4 3 13 1 1 15 3 2 16 15 13 10 3 0 9 1 10 9 2
37 15 10 13 1 3 16 11 4 14 3 13 15 0 9 1 10 11 11 11 11 2 13 15 14 13 1 10 11 9 9 1 11 2 11 2 11 2
11 16 15 13 3 0 1 10 9 13 0 2
26 7 15 13 0 16 14 3 4 11 13 1 1 15 11 11 9 2 7 15 13 1 1 15 9 9 2
48 10 3 2 13 9 1 11 14 9 11 11 2 10 13 1 11 11 11 14 2 10 11 13 1 11 12 2 12 2 13 10 0 9 16 15 15 13 1 14 13 14 13 1 11 1 10 9 2
16 2 10 11 13 2 12 9 11 2 2 11 11 12 2 12 11
29 10 9 9 2 15 4 13 9 16 16 11 11 11 13 15 9 1 10 11 11 1 10 0 9 1 10 0 9 2
31 1 9 2 9 13 11 1 9 1 9 7 9 15 4 4 13 13 11 11 1 10 9 15 4 13 1 10 11 11 3 2
29 15 13 12 9 1 11 3 11 11 13 0 3 3 9 2 10 9 1 11 1 11 11 9 11 2 11 2 11 2
21 11 11 4 3 13 16 13 1 11 13 10 9 15 13 1 10 11 11 11 11 2
16 11 14 11 11 13 10 9 1 11 11 14 9 1 10 9 2
4 11 11 13 2
25 1 12 2 11 11 13 10 0 2 0 0 9 3 2 3 1 10 9 1 10 0 11 11 9 2
22 11 13 11 11 11 14 9 2 7 1 10 9 2 15 13 10 9 1 10 9 9 2
22 13 15 1 10 0 0 9 1 11 2 7 15 13 15 12 9 3 16 15 13 9 2
9 11 11 11 2 0 9 9 2 2
10 15 4 13 9 9 7 10 0 9 2
11 15 13 3 0 14 13 3 1 10 9 2
10 1 10 9 2 15 4 13 15 9 2
6 15 13 10 11 9 2
7 7 15 3 13 1 9 2
23 11 2 10 9 11 11 4 13 1 2 11 11 2 4 13 0 1 11 1 10 9 9 2
13 0 0 11 13 9 1 10 0 9 1 10 9 2
17 11 14 9 1 10 9 13 15 14 4 13 11 11 14 11 11 2
19 1 11 2 11 13 9 7 9 9 1 11 11 14 9 2 3 11 11 2
22 15 13 3 12 2 9 2 0 11 11 13 1 11 2 1 15 9 14 9 2 2 2
18 15 13 11 11 14 9 14 13 10 0 9 9 1 10 12 11 9 2
24 3 1 12 1 10 0 9 2 0 0 9 4 14 13 0 1 10 9 1 0 11 11 9 2
16 7 1 11 2 15 13 11 7 11 15 13 14 13 11 11 2
28 15 13 10 0 11 14 9 14 13 1 15 10 9 9 13 1 10 9 1 9 9 7 13 10 9 1 15 2
20 11 13 10 9 13 11 11 13 3 3 1 10 0 11 9 2 9 13 0 2
32 2 2 2 11 11 13 11 11 14 9 1 9 2 7 1 12 2 15 4 13 1 10 12 2 9 9 1 11 1 10 9 2
19 11 13 16 1 10 9 0 1 0 9 2 11 11 13 14 12 1 15 2
25 11 11 11 2 9 1 11 11 2 2 6 2 15 4 13 3 3 1 10 9 7 13 1 9 2
21 3 2 11 4 13 3 3 9 2 15 4 3 13 3 12 7 12 1 10 9 2
47 11 2 11 13 16 12 9 1 10 9 2 1 11 1 12 2 11 11 14 9 9 13 1 15 7 13 16 15 3 13 1 11 11 14 9 16 10 9 9 4 14 13 3 1 10 9 2
24 11 11 2 11 3 4 14 13 14 13 10 9 16 15 13 1 10 9 1 10 9 9 3 2
26 15 0 9 13 16 15 4 14 13 3 0 1 10 9 1 10 0 9 15 4 13 1 10 9 9 2
24 11 2 11 11 13 16 3 3 2 15 4 14 13 16 11 11 4 13 1 10 11 11 11 2
18 16 15 13 1 1 9 0 2 11 13 14 13 1 11 11 1 15 2
23 10 11 13 10 9 7 11 4 13 10 9 2 3 2 15 13 15 13 9 14 13 1 2
17 11 11 2 11 4 14 13 10 9 3 3 16 13 1 10 9 2
17 1 9 2 3 15 13 10 9 1 15 2 15 3 13 10 9 2
20 15 13 14 0 1 15 2 7 15 3 13 10 9 7 4 14 13 1 15 2
16 11 2 3 1 11 7 11 2 11 2 11 11 13 15 9 2
11 15 13 10 0 0 9 13 1 10 9 2
12 15 13 3 1 10 9 7 13 10 0 9 2
38 1 9 2 15 13 10 9 15 13 1 0 9 2 1 9 1 10 9 7 10 9 13 2 16 10 11 9 15 13 15 3 13 1 10 0 9 9 2
36 11 13 11 11 4 13 1 10 9 7 2 1 10 0 9 2 13 1 9 1 10 9 15 4 13 10 9 3 2 3 3 1 10 9 9 2
15 11 11 2 9 13 0 9 16 13 10 9 1 10 9 2
26 15 4 13 14 13 1 15 9 2 15 4 13 14 13 1 9 2 15 4 13 14 13 1 10 9 2
24 7 15 13 3 15 13 9 2 15 4 13 13 16 16 15 4 13 3 3 10 9 3 13 2
20 11 2 11 13 10 9 1 10 11 11 13 10 9 13 3 2 0 1 15 2
22 11 11 2 15 13 2 1 10 9 2 15 13 12 2 11 4 4 13 12 7 12 2
39 7 15 13 15 13 3 0 16 9 1 15 9 4 13 9 2 3 1 10 9 1 9 3 3 1 10 11 0 9 2 16 13 1 15 9 10 9 3 2
10 15 13 15 0 7 2 3 2 0 2
51 11 2 13 1 11 2 11 11 4 3 3 13 9 1 15 9 1 11 1 11 11 2 7 3 3 15 4 13 3 1 0 9 2 15 4 13 13 16 10 9 13 15 13 10 9 1 10 11 11 11 2
27 11 2 10 0 2 9 11 9 2 15 2 1 10 9 2 13 3 10 13 11 2 4 14 13 10 9 2
34 11 11 2 15 13 15 3 15 4 13 2 3 3 16 10 9 9 13 1 16 15 13 10 9 1 11 11 2 15 4 13 15 13 2
9 7 15 4 3 13 1 15 2 2
14 11 3 13 16 11 11 4 14 13 11 13 0 9 2
22 7 15 13 9 2 16 15 13 14 10 9 1 9 9 1 11 13 10 2 9 2 2
11 15 4 13 14 13 1 11 7 13 15 2
15 3 2 9 1 10 9 1 9 4 14 13 10 9 0 2
12 15 9 13 1 9 7 15 9 13 1 9 2
18 15 4 14 4 13 1 10 9 1 10 9 15 13 15 9 1 15 2
12 3 10 9 13 1 9 1 10 13 9 1 9
8 3 13 16 9 13 14 10 9
12 7 15 13 1 0 14 13 3 12 9 13 9
11 3 13 16 9 13 14 10 9 2 11 11
17 0 15 4 14 13 9 9 14 13 15 2 7 10 9 13 9 2
20 1 11 14 11 10 9 2 2 4 12 9 13 1 10 9 1 11 9 2 2
12 2 3 13 10 9 1 10 11 9 9 2 2
22 10 12 9 10 11 13 1 0 9 9 4 4 4 13 1 9 2 15 4 13 9 2
21 10 12 2 9 9 1 9 13 14 4 4 3 13 3 1 10 11 9 1 11 2
9 7 10 12 9 1 9 4 13 2
16 9 16 10 9 14 13 3 4 13 1 10 11 11 1 11 2
15 7 10 9 4 13 1 1 10 0 9 1 0 9 9 2
29 7 10 0 9 13 14 13 10 9 4 13 1 10 11 1 12 16 13 9 1 11 2 0 9 9 11 4 13 2
24 15 13 10 0 9 13 16 9 1 9 13 1 11 14 9 7 9 3 13 1 11 2 11 2
21 11 0 9 11 11 13 2 2 15 13 0 16 10 9 4 13 1 12 9 9 2
13 16 10 9 4 13 0 15 13 10 0 9 2 2
21 0 9 9 13 10 11 9 14 13 10 9 2 1 10 9 0 9 2 1 11 2
24 7 9 9 9 1 11 13 10 9 1 10 9 2 10 3 13 1 1 11 12 7 11 12 2
31 10 9 9 9 13 15 4 14 13 2 10 9 1 11 2 7 13 15 13 2 14 0 1 10 9 1 11 1 11 2 2
27 11 7 11 9 4 3 13 9 16 0 9 2 13 1 11 2 0 7 0 9 2 4 4 13 1 9 2
22 10 11 9 13 2 2 15 13 10 9 9 14 13 15 4 14 13 1 10 0 9 2
12 15 13 9 16 10 4 4 4 13 1 2 2
28 10 9 10 9 13 12 11 9 13 0 1 10 9 1 10 9 1 9 1 0 9 4 13 1 11 2 11 2
17 10 0 9 13 11 2 7 6 2 15 13 12 1 11 11 14 2
37 15 13 3 10 13 2 15 2 9 2 1 2 10 2 9 9 2 13 3 10 9 10 9 9 13 2 3 1 10 1 10 9 14 0 0 9 2
51 7 3 2 3 14 13 1 10 2 9 2 4 13 9 1 10 9 2 13 3 0 0 9 13 1 10 11 11 10 9 2 7 3 0 1 2 0 9 2 4 4 13 1 10 0 9 1 9 7 9 2
43 1 10 9 1 9 1 9 10 4 4 2 13 2 1 11 2 9 1 9 4 14 3 2 13 2 2 3 3 10 11 13 10 9 1 10 0 9 1 11 14 0 9 2
31 7 11 14 9 13 14 0 14 4 13 16 10 9 10 9 13 2 16 15 13 1 3 0 9 1 10 9 14 13 9 2
16 3 2 10 9 4 4 13 1 10 9 1 11 9 11 11 2
5 7 15 13 9 2
33 10 11 11 11 13 0 2 0 16 10 9 14 9 9 4 13 2 7 15 13 3 7 13 1 15 9 16 4 13 3 1 9 2
1 5
21 10 9 13 1 10 9 13 10 9 9 1 0 9 1 10 11 1 11 1 12 2
38 9 13 10 9 2 11 11 11 2 12 2 4 13 7 3 13 2 16 12 9 1 15 9 13 10 9 1 10 13 9 2 10 3 2 13 0 9 2
23 10 9 9 4 13 1 15 3 2 0 9 2 10 4 13 16 16 15 4 4 3 13 2
21 2 15 13 16 3 15 4 13 15 10 3 2 2 9 11 11 13 1 13 9 2
16 2 15 13 10 9 16 9 14 13 2 3 1 11 15 2 2
52 1 10 9 12 1 11 14 0 9 2 13 1 11 11 2 10 0 9 1 10 11 11 1 15 13 1 11 2 11 2 2 15 4 13 13 10 9 2 7 13 15 2 2 15 13 15 13 1 9 2 2 2
9 1 11 14 9 1 10 11 9 2
30 3 1 3 2 9 7 9 13 10 9 7 10 9 14 13 1 0 9 2 3 3 10 9 13 3 0 9 7 9 2
10 3 9 7 9 13 0 2 9 13 2
25 3 9 7 9 13 1 2 3 3 3 10 9 4 13 2 10 9 4 13 2 7 9 4 13 2
9 10 9 9 2 11 14 9 9 2
22 3 2 1 10 9 2 10 9 2 9 1 10 9 1 10 9 1 10 11 9 9 2
21 11 11 11 11 11 11 2 10 9 15 13 10 9 0 9 2 4 3 13 3 2
42 7 1 10 10 9 15 10 9 4 13 14 13 10 9 2 13 9 0 1 11 11 2 10 0 9 1 10 11 11 2 15 13 1 9 1 10 9 7 10 0 9 2
6 11 13 0 1 0 2
7 9 7 9 13 10 9 2
6 10 9 13 10 9 2
5 10 4 2 3 2
3 7 3 2
11 15 13 3 10 9 1 15 15 13 14 2
20 9 1 0 9 3 3 9 11 2 13 11 7 10 0 0 9 1 10 9 2
8 4 15 13 15 1 11 3 2
9 13 16 9 9 3 13 10 9 2
4 9 1 9 9
40 0 0 9 4 13 1 10 0 11 1 10 0 7 3 0 9 1 9 3 16 10 9 13 1 10 11 11 11 11 2 11 2 13 15 1 0 11 1 12 2
1 5
73 3 2 11 9 11 11 4 4 13 1 10 11 14 9 1 2 12 3 13 9 2 2 10 9 10 13 9 9 14 0 9 1 9 1 10 0 9 1 0 9 2 2 1 1 2 10 9 10 10 9 14 9 2 9 9 9 13 2 4 13 1 10 3 0 1 10 9 2 3 9 7 9 2
95 3 10 11 1 11 11 2 7 15 9 1 15 2 13 1 10 12 9 1 0 0 9 1 13 9 1 5 12 12 2 3 15 13 0 16 9 9 2 9 9 2 7 9 1 10 9 4 13 0 1 10 9 2 3 9 3 13 9 7 0 9 9 2 3 13 0 9 13 14 13 0 9 2 2 7 3 10 9 13 14 13 0 9 2 9 7 0 9 13 14 13 3 3 3 2
1 5
28 3 2 11 4 13 1 11 7 11 1 0 9 1 0 9 7 16 13 2 0 2 9 1 9 7 0 9 2
32 1 9 9 9 1 11 11 11 7 11 2 11 7 9 9 13 11 2 4 13 0 7 0 7 4 4 13 1 0 9 2 2
23 1 10 9 2 15 4 13 1 0 9 1 10 0 9 1 10 9 2 13 1 0 9 2
1 5
28 1 1 11 11 7 0 9 2 0 9 13 1 10 11 11 7 10 0 11 11 2 11 4 13 9 3 3 2
40 2 10 0 9 13 10 9 1 10 10 9 4 3 13 0 14 13 9 1 10 9 2 2 11 4 13 16 13 1 10 11 11 11 11 14 2 9 9 2 2
71 10 9 1 10 9 2 13 11 11 11 1 11 11 11 3 10 9 13 16 2 10 9 14 9 2 10 0 9 1 0 9 2 7 10 9 14 13 1 10 9 14 9 1 10 0 9 4 3 3 13 1 10 9 2 9 9 9 7 9 2 9 9 4 13 3 13 1 0 9 2 2
1 8
20 3 15 4 13 9 3 2 7 3 2 3 2 4 15 2 13 2 12 9 2
10 2 15 13 10 9 9 1 9 2 2
3 6 6 2
5 10 9 14 13 2
13 15 13 0 10 9 1 9 13 3 10 10 9 2
10 15 3 13 15 1 15 3 13 9 2
8 3 13 3 2 15 13 3 0
3 10 11 11
7 15 13 6 12 0 9 2
20 3 2 3 3 2 15 13 10 9 10 9 4 14 13 1 1 10 11 9 2
13 0 3 10 9 4 13 3 1 3 2 13 9 2
16 3 16 15 13 1 10 0 9 5 9 1 9 5 0 9 2
28 15 13 1 10 9 14 3 3 3 10 9 4 13 14 13 10 0 9 13 1 10 9 16 3 13 9 9 2
18 3 3 9 9 4 13 15 9 3 9 4 13 9 1 10 9 15 2
22 3 15 4 14 13 10 9 15 9 13 1 12 10 3 3 16 15 13 10 9 13 2
18 15 13 10 9 9 1 0 9 1 0 9 3 0 9 10 13 15 2
22 3 10 9 13 9 7 10 9 7 9 13 1 9 16 10 9 4 13 10 0 9 2
20 1 10 11 11 9 15 13 9 16 10 9 13 15 7 14 13 10 0 9 2
11 9 13 9 7 9 9 1 10 0 9 2
19 10 0 9 1 9 4 13 3 1 10 9 3 1 3 3 1 10 9 2
25 15 13 0 7 10 9 13 14 13 10 9 1 10 9 14 13 1 10 9 3 1 10 13 9 2
18 10 9 13 15 14 13 13 7 15 13 15 13 14 13 10 9 0 2
8 13 1 9 9 1 0 9 2
7 3 13 1 10 11 9 2
26 12 9 3 4 13 16 13 15 9 9 0 3 15 13 3 1 2 9 2 1 15 9 14 0 9 2
12 10 9 4 13 1 13 9 2 3 10 9 2
8 3 15 2 13 2 10 9 2
7 15 13 10 0 9 3 2
16 15 4 14 13 10 9 14 13 1 1 9 14 13 1 15 2
14 3 10 9 4 13 7 10 10 0 9 4 3 13 2
21 15 13 10 0 0 9 1 9 16 13 10 10 9 9 0 1 10 10 9 9 2
13 15 3 4 13 10 9 9 3 2 13 14 15 2
9 3 10 0 11 9 9 2 6 2
26 6 2 15 4 13 11 4 13 10 9 0 16 10 9 13 15 16 15 4 13 1 9 1 0 9 2
18 15 13 16 15 13 3 0 1 10 11 16 15 4 13 1 0 9 2
14 11 13 0 9 2 9 1 11 9 9 2 9 9 13
39 10 11 4 13 0 11 9 9 7 13 1 10 0 7 0 9 1 9 1 9 14 13 9 1 11 1 9 1 10 0 9 2 0 7 0 9 9 13 2
1 8
11 10 9 13 10 9 15 13 2 15 9 2
20 7 11 2 10 0 2 3 0 2 9 9 1 9 2 13 3 3 10 9 2
14 16 10 9 13 14 13 2 10 11 13 10 9 9 2
17 2 2 15 13 12 9 1 9 2 9 2 9 2 9 2 2 2
24 0 1 10 9 15 4 13 4 13 3 1 11 9 1 11 2 3 15 13 13 1 15 9 2
10 9 9 4 13 1 11 9 7 11 2
46 3 11 13 11 2 0 1 10 9 4 13 1 11 7 3 13 1 0 9 2 11 2 11 2 11 2 11 2 11 2 10 11 11 2 3 15 4 13 1 9 15 13 3 11 9 2
26 3 15 13 12 7 12 2 0 1 15 13 14 13 3 1 11 7 13 10 9 1 10 0 11 9 2
37 16 2 9 2 13 3 14 10 0 9 2 16 1 10 9 15 4 13 2 10 9 7 9 4 14 13 14 13 1 15 7 14 3 13 15 9 2
50 2 10 9 7 9 2 10 9 2 13 3 3 1 12 7 12 2 13 14 13 1 10 9 1 11 7 11 2 13 15 7 13 9 1 15 2 2 11 11 2 10 0 11 0 2 9 2 13 15 2
39 11 2 15 4 13 1 11 7 13 0 16 13 11 9 1 10 11 11 2 13 16 3 10 0 9 13 14 13 11 9 1 15 9 9 2 10 11 13 2
14 0 1 10 9 4 13 1 11 9 2 3 1 11 2
20 10 11 2 11 13 3 14 13 2 2 13 10 9 1 10 0 9 14 9 2
10 15 13 14 13 15 7 13 15 2 2
33 10 4 13 10 9 1 15 9 2 10 9 1 9 2 9 7 10 9 1 9 2 9 13 1 10 9 7 9 1 11 7 11 2
1 9
37 15 13 14 13 16 10 0 9 1 15 9 7 9 15 13 1 10 9 1 10 9 4 14 13 15 15 13 2 4 14 13 2 7 13 3 3 2
2 11 2
12 11 13 15 1 10 9 1 10 9 9 2 8
2 6 2
2 9 9
14 11 11 2 11 13 10 9 9 9 9 1 0 9 2
15 15 13 10 15 13 2 15 4 13 9 14 13 1 15 2
9 11 3 13 11 13 0 1 9 2
5 7 9 1 15 2
1 8
23 2 10 9 1 0 9 4 13 1 2 7 2 6 2 15 13 14 3 1 9 7 9 2
10 6 2 15 13 3 1 9 7 9 2
8 7 15 4 13 3 1 15 2
26 7 3 7 3 2 16 9 13 1 10 0 0 9 10 13 1 9 2 15 4 13 14 13 9 0 2
15 15 4 13 10 9 1 9 2 14 9 9 2 0 9 2
36 9 13 2 13 10 9 1 0 9 1 9 2 9 2 0 9 7 9 2 10 9 16 13 15 9 1 10 9 1 9 4 13 1 2 11 2
2 6 2
21 10 9 15 13 1 10 0 9 5 9 5 9 9 9 13 9 13 9 13 9 2
17 10 0 9 13 11 2 7 6 2 15 13 12 1 11 11 14 2
20 10 11 9 1 11 13 3 10 9 2 13 1 9 14 13 10 9 1 15 2
1 8
8 3 2 13 10 9 1 3 2
9 15 13 2 9 13 10 9 2 5
2 11 2
5 15 13 2 6 2
10 3 13 9 1 9 7 9 2 9 2
15 15 1 11 14 9 13 10 9 2 2 13 15 9 2 2
19 7 4 10 11 9 13 1 10 2 0 9 2 3 15 3 13 15 9 2
18 15 13 9 9 13 9 2 3 13 10 9 9 9 2 6 2 9 2
28 2 14 9 9 2 6 15 13 0 2 13 15 9 2 6 6 2 13 15 9 2 3 15 13 0 9 2 2
5 3 2 6 3 2
13 15 13 10 13 9 1 10 13 9 1 10 9 2
9 10 0 9 1 9 2 1 11 2
21 15 13 10 9 13 3 3 16 3 15 13 10 9 3 1 9 1 10 11 9 2
62 3 15 4 13 1 10 9 9 9 3 1 10 9 1 9 1 1 10 0 9 1 10 8 9 1 10 0 9 1 10 2 9 2 9 2 9 2 10 13 10 9 1 9 9 16 13 15 9 2 7 4 14 13 10 9 3 3 1 15 0 9 2
33 10 0 15 13 2 10 11 13 10 0 9 14 13 14 13 1 1 10 9 7 9 13 1 1 9 2 13 2 16 0 2 11 2
8 9 13 0 2 3 13 9 2
4 15 13 15 2
6 15 4 13 15 9 2
14 6 2 15 13 14 3 0 7 0 0 1 10 10 2
24 15 4 13 1 10 0 7 3 3 0 0 2 0 9 3 10 4 13 0 9 7 0 9 2
20 10 11 11 9 13 1 10 0 9 4 13 1 10 0 9 9 1 0 9 2
9 10 13 9 13 1 10 11 9 2
18 0 9 13 0 7 0 2 0 9 13 0 2 0 2 0 2 0 2
15 0 9 13 0 2 0 9 13 3 0 2 0 2 0 2
3 2 11 11
2 11 2
7 15 4 14 13 3 3 2
22 10 9 13 3 9 2 10 1 10 0 2 1 16 15 13 10 0 9 15 13 1 2
13 7 1 15 2 1 9 2 15 3 13 3 3 2
32 3 13 10 9 2 3 10 3 3 0 13 9 10 13 0 7 0 2 15 13 10 3 0 9 16 15 13 0 7 0 9 2
21 15 13 15 7 15 14 4 13 1 15 9 2 16 15 2 13 16 15 4 2 2
1 8
5 16 3 13 10 9
13 7 3 15 13 13 16 15 3 4 4 13 0 2
28 16 10 9 13 3 1 2 9 9 2 15 13 10 9 13 10 0 9 7 15 3 13 3 0 9 1 9 2
1 8
40 12 9 14 0 9 1 15 0 9 13 15 14 13 12 1 10 3 0 9 1 0 11 2 10 9 1 11 7 9 10 4 13 10 9 1 0 1 10 9 2
15 1 11 12 11 11 7 11 11 2 3 3 12 2 13 2
27 15 4 4 13 1 10 9 13 10 11 2 10 9 1 10 0 9 9 1 11 2 7 15 3 13 3 2
15 10 9 7 0 1 15 9 3 13 15 4 13 3 3 2
8 7 15 9 13 14 13 15 2
26 11 11 2 11 14 9 2 13 14 13 9 9 7 9 1 11 2 13 1 9 7 13 11 14 9 2
42 11 7 15 9 13 1 10 3 0 9 1 0 9 9 2 9 9 7 0 9 2 9 0 1 9 1 9 7 11 2 7 10 9 1 10 9 13 0 1 10 9 2
16 10 9 4 13 15 3 15 13 16 0 9 7 11 4 3 13
2 11 11
24 15 13 16 11 2 10 9 15 13 1 11 2 13 10 9 1 0 9 7 9 1 15 9 2
20 1 10 9 2 11 11 13 0 16 11 13 9 14 13 1 15 9 14 9 2
18 2 10 9 4 13 15 3 15 13 16 0 9 7 11 4 3 13 2
8 15 13 0 2 2 15 13 2
25 6 2 15 13 11 13 1 12 1 15 9 3 1 10 0 0 9 2 2 1 9 1 9 2 2
20 15 3 13 2 7 4 13 10 9 14 13 2 2 1 9 1 9 9 2 2
20 10 0 9 3 13 16 10 9 4 3 13 10 0 0 9 2 2 2 2 2
16 13 1 10 13 2 15 2 9 2 1 2 10 2 9 9 2
15 7 1 2 11 2 3 2 13 1 10 9 9 4 13 2
6 15 4 13 15 3 2
20 4 15 3 13 11 2 7 9 1 0 13 0 1 0 9 1 11 1 11 2
28 2 15 13 2 0 9 2 3 3 13 15 2 7 10 0 9 2 11 2 2 3 16 15 15 13 10 9 2
5 15 13 3 9 2
12 9 15 13 13 10 9 2 7 15 1 10 2
7 3 3 3 13 15 9 2
6 15 3 13 15 9 2
50 15 13 14 4 13 1 2 11 2 2 7 15 3 13 16 1 10 1 15 2 10 9 1 15 9 13 0 1 0 0 9 2 7 13 10 9 0 14 13 1 10 0 9 14 9 1 10 9 9 2
15 15 13 14 13 3 2 0 2 16 3 15 13 10 9 2
14 13 15 16 15 13 2 7 16 15 15 13 14 13 2
37 2 10 3 0 9 1 0 9 9 2 9 9 7 0 9 2 9 0 1 9 1 9 7 11 2 7 10 9 1 10 9 13 0 1 10 9 2
29 3 10 1 10 9 9 9 9 1 10 0 0 9 2 1 1 0 9 2 4 13 2 0 2 1 10 11 11 2
28 11 11 3 13 10 9 1 2 0 9 2 1 12 2 16 13 10 0 9 1 2 0 2 9 1 10 9 2
10 10 0 9 9 4 13 1 10 9 2
17 3 13 10 0 9 1 10 11 11 2 11 11 2 9 1 12 2
1 8
48 3 2 7 3 14 2 2 10 9 1 10 2 9 2 7 2 0 9 2 4 13 1 10 11 7 15 9 4 4 13 3 1 0 2 9 2 11 11 7 10 12 9 15 13 13 11 2 2
12 11 13 3 10 8 9 1 10 11 11 11 2
27 3 10 3 3 0 13 9 10 13 0 7 0 2 15 13 10 3 0 9 16 15 13 0 7 0 9 2
21 15 13 15 7 15 14 4 13 1 15 9 2 16 15 2 13 16 15 4 2 2
3 10 9 2
25 4 10 9 1 2 0 11 2 7 9 1 0 9 13 7 13 1 10 9 14 13 2 9 2 2
12 4 10 9 13 1 7 13 1 10 0 9 2
31 13 16 16 15 13 10 0 9 4 13 1 10 2 0 2 11 1 11 7 10 3 11 1 11 2 10 13 10 0 9 2
7 13 10 9 0 7 0 2
6 4 10 9 3 13 2
15 15 13 3 10 8 2 0 9 1 10 9 13 1 9 2
2 0 2
2 6 2
9 3 2 11 2 15 13 15 9 2
7 3 4 14 15 13 15 2
18 15 9 13 16 15 13 3 3 9 7 15 13 0 1 1 10 9 2
6 3 13 10 0 9 2
5 11 11 1 11 2
25 2 4 14 13 14 13 11 3 2 15 13 3 0 16 13 9 13 1 0 0 7 0 9 2 2
1 8
1 8
10 11 13 1 12 1 10 2 9 2 2
37 15 13 9 9 0 1 11 2 11 2 11 2 11 2 11 7 11 7 13 11 14 0 9 1 10 0 9 13 14 13 10 3 0 9 1 9 2
10 14 12 9 2 10 9 4 14 13 2
16 12 9 1 9 2 12 9 13 12 9 2 0 1 12 9 2
13 16 10 9 13 12 9 3 13 3 0 1 12 2
2 11 2
19 3 16 15 13 15 9 10 0 3 3 15 4 13 15 16 13 10 9 2
9 2 15 13 2 3 15 13 2 5
13 13 1 10 9 3 11 11 14 9 4 13 1 2
17 15 13 1 10 9 0 9 14 13 10 9 14 9 7 9 9 2
12 6 7 6 2 10 11 13 3 1 10 9 2
11 12 0 9 13 9 1 10 0 9 9 2
20 3 13 15 9 7 5 7 9 9 1 10 9 7 15 4 13 1 15 9 2
9 15 4 13 1 10 9 15 13 2
12 0 0 9 2 7 3 13 7 9 2 0 2
15 15 13 13 10 9 10 4 4 13 10 1 15 14 13 2
9 15 4 4 13 3 0 14 13 2
12 4 9 13 10 9 3 1 11 1 11 11 2
1 8
10 15 4 14 13 16 15 4 4 13 2
21 7 3 13 9 1 0 9 2 10 9 1 10 9 13 1 15 0 9 2 3 2
34 15 13 14 13 10 9 9 13 1 1 11 14 9 16 15 13 14 3 13 10 9 2 7 15 13 0 14 13 15 3 13 10 9 2
37 16 15 13 10 9 2 15 13 10 0 9 1 9 7 9 1 15 13 15 2 7 15 1 10 9 1 10 9 15 3 13 2 13 15 1 2 2
11 11 2 15 9 13 0 2 0 7 0 2
33 1 10 9 9 9 2 11 4 3 13 9 2 9 1 2 11 11 2 2 2 11 11 2 9 1 15 0 9 2 11 11 11 2
14 0 11 11 1 11 14 9 1 10 13 9 1 9 2
1 8
4 5 0 9 2
5 3 0 2 3 0
22 15 4 4 13 1 9 2 7 3 13 10 11 14 13 10 9 3 15 13 1 15 2
13 7 15 4 13 10 9 1 15 2 6 13 10 9
10 5 3 4 11 13 11 11 12 9 2
2 1 11
9 11 11 12 2 12 1 12 9 11
14 16 13 10 11 9 9 2 15 13 10 13 0 9 2
27 0 9 2 9 1 0 9 12 2 12 2 12 2 12 2 7 12 2 7 2 9 2 1 0 9 12 2
14 15 4 14 13 15 13 10 0 9 9 15 13 11 2
18 15 13 0 16 13 1 10 9 1 9 2 15 13 1 3 0 2 5
22 15 13 10 0 9 7 1 10 9 11 4 14 13 15 1 9 2 7 13 15 11 2
2 11 2
33 3 2 10 9 13 10 0 2 0 2 9 2 9 2 7 3 2 0 2 3 3 2 16 15 13 1 10 9 1 9 7 9 2
14 1 9 2 13 10 9 1 0 11 10 13 0 9 2
13 7 4 15 13 14 3 13 10 9 1 0 9 2
18 3 2 13 13 0 0 9 7 9 10 9 1 10 0 7 0 9 2
20 1 15 9 2 9 4 3 3 13 14 13 1 7 13 0 0 7 0 9 2
21 10 2 0 9 2 7 3 0 0 2 9 2 4 3 13 7 13 1 10 9 2
29 1 9 1 9 9 2 10 9 13 2 3 3 2 10 9 1 9 2 9 7 10 0 9 1 9 1 0 9 2
12 4 15 13 10 9 1 9 9 11 3 3 2
13 11 13 3 12 1 10 0 2 9 9 2 9 2
10 11 2 16 15 4 3 13 10 9 2
19 10 9 1 10 9 2 9 9 1 15 3 2 7 15 13 1 15 9 2
12 15 0 9 13 1 9 9 2 1 10 9 2
6 0 9 13 0 9 2
21 15 3 13 0 0 1 2 11 2 2 16 15 13 10 0 9 3 15 13 1 2
54 3 2 15 13 3 0 1 10 9 16 15 1 9 3 2 7 2 1 0 2 3 9 1 10 9 1 10 0 9 9 2 13 14 13 10 0 9 1 10 9 14 13 15 0 9 7 1 10 9 14 13 10 9 2
27 15 13 10 9 16 9 4 13 1 9 9 11 14 9 14 13 10 11 2 7 0 13 14 13 3 10 2
16 15 13 14 13 9 1 2 1 15 9 4 15 13 15 2 2
27 15 4 13 15 9 3 10 9 3 9 13 3 10 0 2 9 2 7 2 9 13 15 13 15 2 9 2
50 16 15 4 14 13 1 10 9 16 10 9 15 13 7 13 1 13 10 9 1 15 9 2 10 15 13 13 3 0 2 2 15 4 13 15 3 9 13 1 10 0 9 1 9 14 13 10 9 1 2
14 9 2 16 10 9 13 2 4 14 13 1 10 9 2
29 3 2 15 13 10 9 13 9 15 13 3 3 1 15 0 9 2 7 13 14 13 15 0 9 10 9 3 3 2
25 10 9 13 0 16 15 4 9 2 13 1 2 11 11 2 7 13 3 1 2 3 11 11 2 2
14 2 10 9 1 9 7 9 13 10 0 0 9 2 2
41 15 13 9 1 9 1 9 15 13 1 9 2 9 2 7 9 2 7 15 13 0 14 13 16 11 2 7 2 11 2 2 4 14 13 10 9 1 10 0 9 2
2 9 2
41 10 9 16 10 11 9 7 9 4 13 10 9 9 16 11 13 14 13 9 2 7 3 12 1 10 9 11 13 14 13 13 0 1 15 9 1 11 13 3 0 2
39 15 13 10 9 4 4 13 3 1 11 7 13 1 9 3 1 12 1 10 11 14 0 9 7 15 3 13 10 9 14 13 10 9 1 10 9 7 12 2
14 9 3 1 15 9 11 11 16 13 15 3 1 9 2
22 15 13 10 9 1 10 9 13 1 10 0 9 1 10 0 9 1 10 0 0 9 2
9 15 13 10 0 7 3 0 9 2
10 2 10 11 1 10 11 1 10 11 2
23 9 13 1 11 11 1 10 9 1 10 11 11 11 1 10 0 0 9 2 11 2 12 2
48 2 16 15 13 2 15 3 13 10 0 7 0 2 9 2 1 15 9 2 7 2 1 10 9 2 15 11 13 16 15 13 15 0 0 9 1 9 1 10 9 1 10 9 1 10 15 13 2
19 15 4 3 13 7 15 4 3 13 10 9 9 7 15 13 10 0 9 2
31 15 9 4 3 13 16 15 15 13 2 16 15 15 13 7 1 10 9 16 15 9 4 13 1 10 9 1 3 12 9 2
26 15 4 13 15 9 1 15 1 10 0 9 9 2 10 15 4 13 14 13 2 3 15 13 10 9 2
20 15 4 4 13 1 15 10 0 9 7 10 0 9 1 10 0 2 0 9 2
11 3 2 15 4 13 1 15 3 1 9 2
22 15 13 14 13 0 1 15 9 1 10 0 9 1 10 9 7 15 9 1 9 9 2
29 15 13 1 10 0 9 1 11 7 11 2 10 13 3 0 2 3 0 2 7 13 0 0 7 3 0 0 9 2
12 3 4 15 13 1 11 7 15 0 0 9 2
43 16 11 7 10 9 0 1 15 2 1 9 16 15 15 4 13 7 13 1 10 9 9 2 13 14 10 0 9 2 7 4 3 13 10 0 9 1 10 9 1 10 9 2
24 6 2 15 13 10 12 9 2 0 0 2 0 9 2 7 15 13 14 3 10 0 9 13 2
17 10 9 15 13 1 10 11 2 11 9 13 9 14 13 1 11 2
28 10 0 9 13 3 3 1 11 2 3 10 0 0 9 4 13 15 0 0 9 2 13 9 14 13 1 11 2
27 10 0 9 1 11 1 10 9 1 9 1 9 1 12 9 7 10 1 0 11 13 9 14 13 1 11 2
19 11 11 4 14 13 11 2 13 11 11 7 13 15 0 9 1 1 11 2
15 11 4 14 13 0 9 1 11 1 10 9 1 1 11 2
25 11 10 11 4 14 13 9 1 9 1 15 0 9 1 12 9 1 11 11 1 11 1 1 11 2
17 10 11 9 1 11 7 10 0 9 3 13 9 14 13 1 11 2
27 10 0 9 9 1 10 11 2 11 9 13 9 14 13 1 11 2 7 15 4 13 3 7 3 7 3 2
45 10 9 1 10 9 13 16 10 9 0 9 13 3 0 2 1 10 9 1 10 9 2 7 4 4 13 3 3 16 11 4 13 10 11 11 7 10 0 11 4 13 1 12 9 2
39 10 12 9 9 1 10 11 11 2 1 11 1 10 11 11 2 13 10 0 9 1 12 9 2 0 1 10 11 7 3 3 0 1 10 11 1 15 9 2
15 15 13 10 9 9 0 1 7 10 11 7 10 1 11 2
34 10 12 9 2 1 10 15 9 7 0 9 2 13 10 13 11 0 1 15 1 11 7 11 7 0 1 9 1 10 11 1 11 3 2
35 1 10 0 11 2 10 9 1 0 7 0 13 1 9 7 3 0 1 10 0 13 15 9 3 16 13 1 9 2 7 16 13 0 9 2
19 10 0 9 1 9 13 3 16 15 15 13 1 10 11 11 12 9 3 2
26 0 9 13 1 10 0 9 2 1 9 1 10 0 9 16 11 4 13 9 1 10 11 11 11 9 2
40 13 1 10 9 13 1 10 9 1 0 9 7 13 1 10 9 1 10 11 2 10 9 1 9 13 1 10 0 0 9 13 3 0 16 15 0 11 3 13 2
19 10 0 9 1 0 9 1 12 12 11 13 0 1 15 1 12 12 11 2
21 9 9 1 10 9 13 3 0 2 13 10 9 2 10 0 9 7 10 0 9 2
53 7 10 1 15 4 13 1 10 9 2 10 3 12 9 3 2 4 13 14 13 10 0 0 9 1 10 9 2 7 1 10 0 9 2 10 13 2 1 10 9 1 9 2 12 1 10 3 0 9 1 10 9 2
29 15 13 0 14 13 16 15 13 10 0 9 9 1 0 9 2 9 9 2 9 2 9 2 9 9 7 0 9 2
39 15 13 3 10 9 16 3 9 1 10 9 13 10 9 1 10 11 11 2 1 11 2 1 0 9 2 1 11 7 11 2 1 9 7 9 2 1 15 2
57 10 9 1 10 9 1 0 2 0 2 0 9 15 13 7 0 11 7 13 14 3 0 7 13 1 1 0 9 2 15 13 0 9 1 10 0 9 2 10 3 13 9 2 7 1 15 0 9 10 13 15 9 16 13 3 0 2
31 10 9 13 16 10 0 0 9 1 10 11 13 14 9 1 10 9 7 10 9 2 7 15 3 4 14 13 1 1 15 2
22 15 13 9 2 1 9 2 7 15 13 1 0 9 2 9 2 9 9 7 0 9 2
18 0 1 15 4 3 13 9 1 9 2 7 13 0 14 13 15 9 2
32 10 9 1 10 0 0 9 4 13 12 9 2 10 4 3 13 2 7 4 3 13 3 0 1 1 10 0 9 1 10 9 2
24 10 0 0 9 4 13 16 9 13 16 15 13 10 11 11 2 7 15 13 3 3 1 15 2
29 15 13 10 12 0 9 1 10 0 9 9 2 7 3 15 4 3 13 1 15 1 2 10 0 11 11 11 2 2
12 2 8 2 10 0 9 13 10 9 9 2 2
24 9 9 13 14 10 0 9 7 15 4 4 13 0 2 16 15 4 13 10 9 2 3 3 2
20 3 1 11 12 2 15 13 16 0 1 10 11 11 4 14 3 13 10 9 2
8 15 13 10 3 0 0 9 2
8 15 0 0 9 13 3 0 2
27 10 0 9 1 9 1 9 1 9 9 1 11 1 10 0 12 9 13 3 0 1 15 1 1 9 9 2
10 11 12 13 3 3 3 0 1 0 9
31 0 9 13 1 9 1 12 9 1 11 1 10 10 11 15 13 1 10 9 1 11 2 13 0 9 9 16 10 9 13 2
21 11 13 0 9 0 9 1 10 10 15 13 1 9 9 1 10 11 9 1 11 2
10 3 15 13 10 10 9 1 9 9 2
4 15 13 9 2
4 15 13 0 2
4 15 13 0 2
20 15 13 10 3 0 9 1 9 13 7 0 0 0 9 1 0 1 10 0 2
10 15 4 3 13 1 9 1 0 9 2
34 12 0 9 2 1 10 9 1 0 9 9 2 4 13 10 9 9 1 10 9 1 10 10 9 2 16 15 4 1 11 7 1 11 2
24 7 10 0 9 13 1 10 0 9 16 10 9 7 10 0 9 4 13 1 10 0 9 9 2
12 15 4 14 3 13 10 9 1 10 11 11 2
19 10 11 7 11 4 3 13 15 9 1 10 0 9 2 3 10 0 12 2
12 15 4 13 1 10 0 9 9 1 10 9 2
27 7 16 15 13 14 13 1 9 2 15 4 14 13 14 13 10 9 1 9 14 13 15 7 13 0 9 2
23 15 4 13 10 9 9 1 10 9 1 10 0 9 13 14 4 13 1 10 9 9 9 2
16 3 1 10 9 1 10 13 2 1 9 1 10 0 9 9 2
20 13 10 9 9 1 9 1 10 9 9 1 11 7 10 9 4 13 10 9 2
23 13 10 9 7 15 4 13 1 9 9 2 9 9 2 9 2 9 9 2 9 7 9 2
40 13 9 1 9 1 10 9 9 7 15 4 3 13 10 9 1 9 14 4 13 1 10 9 7 10 9 4 13 10 9 2 3 14 13 16 13 10 9 15 2
31 15 4 3 13 15 9 1 0 7 0 9 7 1 0 9 9 7 14 13 15 7 3 14 13 10 9 1 10 0 9 2
6 7 15 13 10 9 2
7 15 13 1 10 9 9 2
16 9 13 2 9 7 9 7 0 2 0 0 9 2 9 0 2
11 15 13 9 14 13 1 0 0 0 9 2
9 10 0 9 4 3 13 15 1 2
15 10 9 1 10 0 9 7 0 9 4 3 13 15 1 2
9 10 9 1 9 0 4 13 15 2
34 4 14 15 13 9 1 10 0 9 14 13 15 15 2 7 14 13 15 9 16 13 15 2 16 15 13 3 10 0 9 1 0 9 2
12 13 14 15 0 1 10 9 16 13 1 11 2
17 3 2 15 13 0 9 2 0 9 2 0 9 7 0 13 9 2
32 15 13 15 10 9 2 3 0 2 1 10 0 9 2 7 13 15 9 3 16 10 0 9 4 13 7 0 0 9 13 0 2
12 9 9 3 13 9 14 13 1 9 7 9 2
13 10 0 9 1 10 9 2 1 3 2 13 11 2
5 15 3 13 3 2
17 15 13 0 0 9 1 10 9 2 1 0 9 2 9 7 9 2
12 9 4 14 13 9 1 9 2 9 7 9 2
22 15 13 3 0 9 1 11 14 11 1 1 11 11 14 11 2 7 10 9 13 15 2
55 10 9 9 13 3 10 0 2 0 9 1 0 2 0 2 0 2 3 2 13 9 2 1 10 9 1 0 9 2 13 10 9 1 15 0 9 2 7 1 3 0 9 1 15 0 0 3 2 9 7 15 9 1 9 2
34 10 0 9 14 13 10 0 2 0 2 9 13 0 1 10 0 9 1 10 15 13 0 9 7 9 1 10 0 9 2 10 0 9 2
32 1 1 10 9 1 0 9 2 15 13 0 16 10 9 1 10 9 13 0 7 15 13 0 14 13 10 9 1 10 9 9 2
17 15 4 14 13 0 9 16 13 10 0 9 9 1 10 9 9 2
12 15 4 13 1 10 9 1 10 2 9 2 2
41 16 9 1 10 9 13 15 2 9 13 15 2 0 13 0 1 15 7 10 13 14 13 15 3 1 9 7 1 10 0 9 2 0 9 4 13 7 3 4 9 2
11 10 11 11 13 15 3 2 1 11 12 2
7 11 4 13 14 13 15 2
5 11 13 15 3 2
15 15 13 3 3 0 16 0 1 11 3 4 14 13 15 2
21 3 2 15 13 16 11 4 13 15 3 16 9 9 13 1 11 1 10 0 9 2
10 1 15 0 9 2 15 4 3 13 2
12 10 0 9 7 10 11 9 13 3 10 9 2
14 10 9 1 10 0 9 16 13 10 9 13 3 0 2
12 16 11 13 1 2 10 9 4 14 4 13 2
14 2 8 2 10 0 9 13 9 2 3 3 9 2 2
5 9 4 13 0 2
4 15 13 9 2
26 15 4 3 13 16 9 2 9 7 3 3 9 7 9 9 4 3 13 2 1 9 1 15 0 9 2
36 7 10 9 1 9 7 9 13 0 2 1 9 1 10 9 1 9 7 0 0 0 9 2 10 4 13 0 9 1 10 9 15 4 13 1 2
30 10 0 9 1 9 1 10 0 9 13 16 11 12 3 13 2 7 13 10 0 9 7 2 3 3 2 10 0 9 2
28 15 10 13 10 0 11 1 11 2 11 11 11 11 2 11 7 15 9 9 3 10 11 9 13 3 1 11 2
10 9 1 9 1 9 13 10 13 9 2
38 7 14 13 2 9 1 9 2 7 14 13 0 0 9 2 0 1 9 14 13 9 2 16 3 4 13 1 15 0 9 2 4 3 13 1 10 9 2
27 11 11 3 13 10 0 9 1 10 9 9 2 7 15 4 14 13 10 3 0 9 16 13 15 0 9 2
22 15 3 4 14 13 10 0 9 16 13 9 2 10 9 2 3 3 2 1 0 9 2
19 3 3 2 16 15 13 14 13 10 9 2 15 13 0 9 16 13 15 2
22 15 4 14 13 14 13 16 10 11 3 13 2 7 16 10 0 9 1 11 3 13 2
15 7 9 1 11 4 13 1 15 9 16 15 13 10 9 2
20 3 10 0 9 13 0 9 2 10 0 9 13 15 16 16 15 4 13 0 2
42 15 13 10 0 9 16 10 0 9 15 13 2 13 7 13 9 9 2 13 10 9 1 11 1 9 1 0 9 9 2 13 1 10 9 9 2 10 3 3 13 15 2
28 15 13 10 0 9 14 13 10 0 9 13 0 9 1 11 1 15 9 7 1 11 1 10 9 1 10 9 2
30 9 1 0 9 2 13 1 9 9 1 13 9 2 4 13 10 0 9 1 15 15 13 2 13 7 13 14 13 9 2
39 0 9 4 13 1 0 9 7 1 9 1 3 2 13 9 2 7 10 0 9 4 14 13 15 16 15 0 9 9 4 3 13 1 9 9 7 9 9 2
25 15 13 1 15 2 3 16 0 1 15 4 14 13 11 2 14 13 11 11 2 1 9 1 9 2
8 15 4 14 13 15 0 9 2
11 7 9 3 13 1 0 9 2 3 0 2
39 10 9 1 11 2 13 9 13 11 14 9 7 13 12 2 9 0 9 13 1 9 9 2 4 13 1 10 9 7 1 0 9 1 10 2 9 9 2 2
30 15 4 13 7 13 10 11 9 2 7 14 13 1 9 1 11 2 11 7 11 11 1 9 9 13 10 9 3 0 2
31 10 9 13 1 10 0 9 1 9 2 13 2 13 9 1 0 9 7 9 13 15 9 1 10 0 9 7 13 10 9 2
24 15 3 13 15 1 2 13 12 9 2 13 0 9 2 16 9 7 9 13 3 1 10 9 2
19 15 4 13 2 9 2 1 0 0 9 7 2 9 2 1 10 0 9 2
14 9 13 10 9 7 13 15 0 9 7 10 9 13 2
52 15 13 10 0 9 1 9 2 10 0 9 4 13 2 10 0 9 2 2 10 9 15 13 15 2 13 15 7 13 15 4 3 13 2 10 0 9 2 7 10 9 1 10 9 4 13 10 2 0 9 2 2
24 15 13 0 0 9 1 0 0 9 2 13 10 9 3 3 1 9 9 7 3 1 0 9 2
11 10 9 13 3 3 0 16 0 9 13 2
8 15 13 10 0 9 1 9 2
20 15 13 11 11 15 13 16 16 15 13 10 9 3 3 2 9 4 13 15 2
9 15 4 3 4 13 1 15 9 2
10 2 8 2 10 0 9 13 9 2 2
31 0 9 1 9 2 10 4 4 13 0 0 9 1 10 0 9 1 10 9 2 4 13 1 12 0 9 13 9 7 9 2
9 1 10 0 9 13 10 9 15 2
17 10 9 13 15 9 2 9 2 9 7 0 9 1 0 0 9 2
31 10 0 9 4 3 13 1 9 9 1 11 7 11 2 1 3 3 1 11 7 11 7 3 3 1 10 1 10 0 9 2
20 10 9 2 3 3 1 10 11 11 2 13 10 0 9 1 10 0 9 9 2
37 15 4 13 1 10 0 0 9 1 0 9 2 9 2 9 2 9 2 10 1 15 13 10 9 2 3 10 3 0 9 2 16 13 1 9 9 2
44 3 2 15 13 10 0 9 1 3 2 13 0 2 0 7 9 9 2 10 3 13 10 9 2 13 10 0 7 13 10 9 2 7 13 10 0 9 1 9 2 9 7 9 2
21 10 9 13 3 1 9 2 9 7 0 0 9 7 3 1 13 0 7 13 9 2
26 15 13 10 9 10 13 0 16 9 13 0 2 16 9 13 0 7 16 9 1 10 0 9 13 0 2
24 15 13 3 10 9 10 13 10 9 16 13 9 1 10 0 9 2 1 10 9 1 10 9 2
65 10 0 9 4 3 13 1 11 11 2 7 3 1 9 1 0 0 9 1 10 11 11 7 11 7 2 1 10 0 9 2 1 9 1 0 9 1 0 9 7 1 0 11 11 9 2 15 9 4 13 0 2 7 15 4 13 7 13 1 9 1 10 0 9 2
27 10 0 9 2 3 3 2 4 13 10 0 9 1 0 9 2 3 10 0 9 4 13 1 10 0 9 2
25 10 11 4 13 14 13 15 2 7 15 13 10 0 9 2 16 3 13 10 9 1 10 0 9 2
36 3 13 2 10 0 9 13 10 9 2 10 13 0 16 10 9 13 7 13 3 1 10 0 9 1 9 7 9 2 3 1 1 10 9 0 2
24 10 9 1 10 0 0 9 3 13 1 10 9 1 9 1 2 7 9 1 2 10 0 9 2
10 10 0 13 9 13 10 0 9 9 2
30 9 1 10 9 1 10 0 9 13 1 10 9 1 12 2 10 3 0 9 1 9 2 13 12 0 9 1 0 9 2
15 10 1 10 9 1 10 0 9 13 3 3 1 15 9 2
21 15 13 15 9 1 10 0 0 9 1 11 2 3 1 10 9 9 1 9 9 2
24 10 9 2 9 2 13 13 9 9 1 11 7 0 9 2 16 10 1 15 9 13 1 11 2
62 11 11 2 15 13 1 11 1 15 9 2 13 9 1 9 1 9 1 9 1 10 13 0 11 11 2 16 10 0 0 9 1 10 11 2 11 9 2 13 1 11 2 13 3 10 9 9 1 10 9 1 12 9 2 16 13 9 1 10 9 9 2
20 2 8 2 10 0 9 1 10 0 9 9 13 10 0 9 1 10 9 2 2
29 10 0 9 13 1 9 2 10 9 1 9 2 13 0 9 2 0 9 2 0 9 7 0 9 2 1 0 9 2
42 15 13 0 0 2 0 9 0 16 13 0 9 7 9 2 14 13 9 7 9 1 9 1 9 2 13 10 9 1 0 9 7 14 13 9 1 0 9 7 0 9 2
26 3 1 9 2 14 3 1 10 11 9 2 13 15 0 0 9 1 10 1 10 0 16 15 13 3 2
21 10 9 1 0 9 13 3 15 13 10 0 9 16 13 10 0 9 7 13 9 2
11 0 9 1 10 0 9 4 3 13 9 2
12 4 10 9 13 9 1 9 13 14 13 15 2
13 4 10 9 13 1 9 9 1 9 7 9 9 2
16 4 0 9 13 15 3 15 13 2 9 2 1 10 0 9 2
11 4 15 13 9 9 2 1 0 0 9 2
8 15 13 10 0 2 0 9 2
9 7 3 15 13 10 0 0 9 2
14 4 15 13 10 9 2 10 13 1 10 0 9 9 2
13 4 15 13 9 2 16 15 4 13 1 10 9 2
15 4 15 13 10 9 13 1 1 9 15 13 10 9 9 2
17 4 15 13 10 9 16 10 0 9 9 13 9 14 13 15 9 2
20 4 15 13 10 9 16 12 13 14 13 0 7 13 10 9 9 1 15 9 2
19 4 15 13 3 1 9 13 14 13 15 2 13 3 1 10 9 1 9 2
12 4 15 13 0 9 2 13 1 10 0 9 2
19 4 15 13 10 9 15 3 13 1 12 9 1 10 2 3 13 1 9 2
13 10 1 15 13 3 1 11 7 1 10 0 9 2
5 15 4 15 13 2
11 6 2 15 4 14 13 14 13 10 9 2
7 7 15 4 14 4 13 2
97 13 2 1 10 9 1 9 2 16 9 4 3 13 1 10 3 2 0 9 1 11 2 13 1 10 0 9 7 13 1 15 2 13 12 9 1 10 1 11 7 1 11 2 13 9 1 0 9 2 13 9 1 10 9 2 13 1 0 9 9 14 13 0 1 10 0 2 16 10 9 1 11 13 0 9 1 15 9 7 13 14 13 15 2 13 15 1 0 9 7 13 15 1 10 0 9 2
23 15 13 15 1 15 1 9 14 13 1 15 11 7 11 4 4 13 2 1 10 10 9 2
22 10 9 13 16 10 0 9 4 3 13 9 1 10 9 1 9 1 10 3 0 9 2
29 15 4 13 14 13 9 9 16 13 10 9 9 2 9 1 10 9 7 14 13 1 10 9 9 1 10 9 9 2
47 1 10 0 9 3 10 9 13 10 9 16 9 13 15 0 9 2 16 10 10 9 13 0 2 0 9 4 14 13 9 13 1 9 2 9 7 9 2 16 4 13 1 15 9 7 9 2
36 0 9 4 14 13 3 14 13 9 15 13 9 14 13 9 2 13 1 15 7 13 1 9 7 4 14 4 13 16 15 4 13 1 10 9 2
40 0 9 4 14 13 3 14 13 1 10 9 1 9 15 4 3 7 3 13 1 10 9 2 10 13 14 13 15 9 7 3 13 14 13 3 0 14 13 15 2
36 10 0 9 13 16 10 1 10 9 13 9 1 0 9 2 7 13 10 10 15 13 15 1 2 9 9 2 2 16 10 0 9 13 10 9 2
24 10 0 9 13 16 10 1 15 13 0 2 16 10 9 1 0 9 4 3 13 15 1 9 2
20 10 9 1 9 9 4 13 9 7 9 1 10 9 2 14 3 7 14 3 2
23 1 10 9 9 2 10 9 1 0 9 4 13 2 7 10 0 4 13 1 10 0 9 2
14 7 1 10 9 9 2 10 9 1 9 4 4 13 2
9 10 9 15 13 3 13 14 0 2
7 15 4 15 13 1 15 2
10 1 10 0 9 2 3 13 7 13 2
17 1 10 0 9 2 3 13 10 0 9 7 13 15 1 10 9 2
11 10 0 9 4 7 4 4 13 1 9 2
10 10 0 9 4 14 4 13 1 9 2
35 3 15 13 0 9 1 10 13 0 2 0 9 1 9 2 0 9 2 9 2 9 3 0 7 9 1 0 9 2 9 7 10 0 9 2
22 1 10 2 15 13 10 0 0 9 7 9 1 10 0 9 1 10 12 9 1 9 2
22 13 15 2 1 10 9 2 14 13 1 15 0 9 1 10 9 9 7 13 1 9 2
15 3 15 13 10 0 9 2 15 4 13 10 9 15 3 2
30 15 4 3 13 15 16 13 0 9 16 13 15 1 0 9 1 10 9 2 3 13 0 2 9 2 16 13 10 9 2
14 16 15 13 14 13 0 2 15 13 0 14 13 10 2
33 7 16 15 13 7 13 2 1 9 7 3 2 15 13 14 13 16 15 13 1 10 9 2 7 15 4 13 11 10 0 0 9 2
32 1 9 14 13 2 15 13 0 14 3 13 10 0 9 2 16 16 10 9 1 10 9 4 13 1 10 0 9 1 10 9 2
46 15 4 14 13 14 13 3 16 16 10 0 2 13 9 1 11 13 0 1 10 9 1 9 1 9 1 0 9 7 10 0 0 9 2 7 15 4 13 1 10 0 9 1 0 11 2
31 3 16 11 2 11 7 11 13 3 2 12 7 10 9 0 9 13 2 11 2 11 7 11 2 10 0 13 10 0 9 2
9 3 11 4 4 13 1 10 9 2
25 1 10 9 1 10 9 1 11 7 11 2 7 11 7 11 4 3 3 13 1 9 0 1 15 2
22 11 4 13 1 11 2 1 10 11 11 2 11 7 10 0 9 1 10 0 11 11 2
12 11 4 13 1 11 2 11 2 11 7 11 2
16 15 13 10 0 0 9 7 15 13 0 9 1 10 0 9 2
19 15 13 14 0 16 11 13 3 0 16 13 14 13 10 0 9 1 11 2
24 15 4 14 13 16 10 0 9 13 3 14 13 7 11 7 11 2 7 15 13 10 13 9 2
19 1 15 0 9 2 10 9 12 9 1 10 9 9 13 11 7 15 9 2
15 15 3 13 9 14 13 0 9 7 14 13 1 10 9 2
11 15 13 10 9 10 13 9 1 0 9 2
4 15 13 0 2
20 15 4 13 16 15 4 13 0 0 9 16 13 3 0 9 2 13 0 11 2
9 15 4 3 13 14 13 0 9 2
25 15 3 2 13 9 7 9 13 15 0 9 9 1 10 2 0 2 9 1 0 2 9 2 9 2
81 11 13 0 9 2 15 13 3 1 0 1 10 9 1 11 2 15 4 3 13 10 11 7 2 1 15 2 10 0 11 7 11 11 2 15 13 9 1 9 3 3 1 11 7 1 11 11 7 3 3 1 11 7 11 11 7 15 3 13 10 0 9 9 2 10 13 2 1 0 9 2 11 2 11 7 0 0 9 1 11 2
22 3 2 0 0 9 3 13 1 11 2 13 14 13 15 7 13 14 13 10 0 9 2
20 1 9 14 13 10 9 15 13 3 0 14 13 10 0 9 1 10 9 9 2
34 15 13 0 14 13 14 13 10 0 9 1 10 0 9 1 11 11 7 11 7 10 0 9 1 11 2 11 7 0 0 2 13 9 2
13 3 15 13 15 9 9 2 10 1 15 13 3 2
24 15 13 0 14 13 0 7 0 0 9 1 10 0 9 2 10 13 10 0 9 9 1 9 2
46 15 13 0 14 13 10 9 1 10 0 9 1 0 9 2 14 13 10 9 1 0 9 9 7 14 13 1 0 0 9 1 10 0 9 1 0 9 1 10 1 10 12 9 1 9 2
33 15 13 3 0 14 13 3 1 10 9 1 9 7 9 7 14 13 10 0 9 15 13 1 15 1 1 9 2 0 9 7 9 2
8 1 10 2 3 13 1 9 2
29 10 9 4 3 13 16 10 0 9 1 11 4 4 13 10 0 9 2 16 3 1 10 9 9 10 0 9 3 2
7 7 15 3 4 14 13 2
23 15 13 13 16 10 9 13 16 15 13 10 9 7 16 15 13 16 13 11 1 1 11 2
36 10 0 9 4 3 13 1 13 3 0 1 0 0 9 2 13 11 2 15 4 3 13 13 9 7 13 9 7 13 9 15 13 9 1 11 2
12 1 10 0 9 2 11 15 4 13 3 0 2
8 13 10 9 10 0 0 9 2
68 16 1 9 15 13 0 9 7 3 0 9 2 0 9 2 10 13 0 9 2 0 9 2 9 1 9 2 0 0 9 2 9 1 0 9 7 9 2 9 1 0 9 7 1 9 2 7 9 1 0 9 13 9 2 9 1 9 7 9 2 3 6 2 9 13 10 9 2
30 16 9 13 3 0 9 2 15 13 0 16 10 3 0 9 4 4 13 2 10 9 15 9 7 9 13 10 3 0 2
17 15 4 13 15 3 1 11 7 2 1 10 0 9 2 1 11 2
14 15 4 13 3 2 16 10 9 4 14 13 3 3 2
52 1 10 0 9 2 10 0 9 9 2 1 1 11 2 4 13 10 0 0 9 2 13 10 9 1 10 0 9 2 3 1 10 0 9 3 10 0 0 9 4 14 13 1 11 7 4 14 4 13 1 11 2
11 15 13 10 9 16 10 0 9 4 13 2
25 7 10 3 15 13 15 14 13 10 0 9 1 10 9 2 10 3 0 7 0 10 9 4 13 2
12 11 2 3 1 10 0 9 2 13 10 9 2
29 15 0 9 1 9 2 13 10 9 1 11 11 11 2 4 13 9 1 0 0 9 2 16 10 9 4 13 2 2
18 11 4 13 1 10 9 1 10 11 11 11 13 1 10 11 1 11 2
26 11 7 10 11 1 11 4 13 14 13 11 14 9 1 11 1 10 0 9 1 0 9 1 0 9 2
31 1 12 2 11 4 13 16 10 11 11 11 4 13 1 15 9 1 10 11 11 7 13 1 1 0 9 1 10 0 9 2
22 10 0 9 13 3 15 13 10 9 9 3 13 1 10 11 11 11 11 11 1 12 2
39 13 1 0 8 9 9 2 7 3 7 3 2 1 10 9 1 10 0 9 13 9 15 13 1 9 7 13 0 14 13 3 10 9 1 10 9 13 15 2
15 11 11 2 11 7 11 2 9 2 9 2 9 9 7 9
2 9 9
44 1 0 11 12 2 10 11 11 11 2 2 11 2 2 9 3 13 16 10 9 1 11 11 14 7 11 11 14 9 1 9 13 1 10 13 9 16 13 0 9 0 1 9 2
52 10 0 11 12 11 9 13 10 9 1 10 11 9 16 1 10 9 1 11 12 11 11 4 13 10 2 0 2 0 9 2 10 9 1 10 4 13 10 9 1 10 9 1 11 11 11 2 2 11 2 2 2
12 15 4 4 13 10 0 9 1 11 2 11 2
32 1 11 12 2 10 9 1 10 11 9 1 9 13 16 11 11 13 0 14 13 0 7 0 9 7 4 13 3 1 0 9 2
39 1 10 9 13 11 12 2 12 2 10 11 11 9 13 16 2 11 11 13 10 0 0 9 9 7 4 13 9 1 15 9 14 13 9 0 1 11 12 2
34 13 1 11 1 11 11 11 11 2 11 11 14 9 14 13 10 9 9 13 12 1 10 3 0 9 10 11 11 13 0 14 13 2 2
48 1 11 12 2 12 2 15 4 13 16 1 10 9 1 12 2 10 9 13 11 2 11 2 3 13 1 11 10 11 2 15 13 9 1 10 2 0 9 2 2 4 4 13 11 11 11 9 2
21 9 1 10 13 9 9 13 10 9 7 10 9 1 10 9 1 10 9 7 9 2
23 1 10 9 2 10 11 13 16 10 9 4 13 1 10 9 14 13 10 0 7 0 9 2
18 10 11 3 4 4 3 13 10 9 16 10 9 9 13 10 0 9 2
5 15 13 0 9 2
24 15 13 3 3 3 3 0 14 3 13 10 11 14 2 0 2 9 1 10 0 2 0 9 2
35 0 9 4 13 16 10 11 2 13 11 11 9 13 1 10 0 9 12 9 9 1 10 11 2 7 16 10 9 13 1 10 9 7 9 2
39 11 9 9 11 11 4 13 16 16 9 4 13 16 16 13 9 4 13 1 10 9 1 9 2 9 1 11 13 16 9 4 4 13 16 0 9 4 13 2
76 2 10 11 14 9 2 2 13 11 11 2 10 11 2 11 9 15 3 13 1 10 11 7 3 13 15 11 11 9 2 2 13 3 2 16 15 13 9 2 13 15 3 3 2 2 10 9 9 13 10 9 1 9 15 13 1 11 12 1 9 9 1 11 2 11 7 11 11 11 2 3 3 1 0 9 2
29 10 9 9 4 13 1 9 1 10 9 1 10 0 9 11 11 7 15 0 1 10 0 11 11 11 9 1 12 2
38 0 9 7 9 1 10 9 13 1 10 9 1 11 2 11 11 14 9 12 2 13 10 0 9 9 9 13 10 9 9 7 13 10 9 1 0 9 2
35 15 15 9 9 4 14 13 15 2 3 2 13 16 10 11 13 10 0 9 1 11 11 14 0 2 9 2 11 11 11 2 12 9 3 2
23 10 9 9 4 13 1 15 1 15 9 1 10 11 1 11 7 13 1 1 10 0 9 2
15 11 2 1 10 9 2 13 10 9 1 11 14 0 9 2
25 15 13 10 9 16 9 13 10 9 10 11 11 4 13 14 13 9 1 0 9 7 9 7 9 2
31 10 4 3 13 16 3 1 10 0 9 1 10 12 9 2 11 11 4 13 14 13 10 0 9 1 10 11 7 11 11 2
22 9 13 16 15 13 14 13 9 1 10 0 9 1 9 13 1 9 1 10 0 9 2
33 15 4 10 9 1 11 2 3 2 13 11 12 2 12 13 16 15 13 14 13 10 9 9 9 10 13 14 13 1 1 12 9 2
29 1 11 12 2 11 3 13 16 11 4 14 13 14 13 9 1 12 7 13 14 13 9 1 10 2 0 9 2 2
36 16 11 11 13 15 5 12 1 11 2 13 11 12 9 11 11 13 15 9 9 16 15 13 10 11 11 9 10 4 4 13 1 10 9 9 2
33 11 13 16 11 14 9 1 9 9 4 4 13 0 1 10 9 9 4 13 1 11 2 13 9 7 11 11 9 2 0 11 11 2
40 11 11 2 3 10 0 9 1 10 9 7 13 1 15 9 14 13 0 2 4 13 10 9 1 15 9 1 10 9 16 15 13 2 9 1 11 9 3 2 2
24 11 11 14 0 9 2 11 2 15 13 1 10 0 11 12 9 7 13 11 2 4 4 13 2
8 11 3 4 13 1 10 9 2
28 11 7 11 13 11 2 11 2 11 2 11 2 2 1 1 11 10 11 2 14 13 11 9 1 10 0 9 2
22 15 13 1 9 1 10 9 1 0 12 3 11 10 11 13 9 9 1 10 11 9 2
23 11 2 13 1 7 11 7 11 2 4 14 13 10 0 11 11 11 9 10 4 4 13 2
11 15 4 13 9 15 13 9 1 10 9 2
42 7 16 9 13 10 9 2 9 4 13 1 10 9 1 11 11 11 14 9 2 0 9 14 13 7 13 9 1 11 9 10 4 13 1 12 9 1 10 0 9 9 2
17 10 9 4 4 13 1 0 9 7 4 13 11 3 1 0 9 2
23 9 1 11 1 11 1 10 9 1 12 13 16 11 13 10 0 9 1 10 11 9 9 2
18 15 13 16 10 11 13 16 10 9 4 13 10 9 13 1 10 9 2
37 2 15 15 13 13 16 15 4 3 13 15 13 10 0 9 14 13 10 0 9 1 15 9 2 2 0 11 11 9 8 9 9 11 11 4 13 2
61 10 11 11 11 13 16 10 9 13 1 11 13 10 11 12 9 10 2 13 10 9 4 13 9 7 9 1 0 9 2 10 15 13 13 2 3 0 1 15 7 13 0 9 1 9 2 10 4 3 13 15 1 10 0 9 2 11 0 2 2 2
18 11 4 13 1 10 9 1 10 11 11 11 13 1 10 11 1 11 2
26 11 7 10 11 1 11 4 13 14 13 11 14 9 1 11 1 10 0 9 1 0 9 1 0 9 2
31 1 12 2 11 4 13 16 10 11 11 11 4 13 1 15 9 1 10 11 11 7 13 1 1 0 9 1 10 0 9 2
22 10 0 9 13 3 15 13 10 9 9 3 13 1 10 11 11 11 11 11 1 12 2
39 13 1 0 8 9 9 2 7 3 7 3 2 1 10 9 1 10 0 9 13 9 15 13 1 9 7 13 0 14 13 3 10 9 1 10 9 13 15 2
36 10 0 9 1 11 12 2 1 10 13 9 9 1 11 1 9 2 14 13 1 10 11 9 2 10 9 9 4 13 1 0 7 2 0 2 2
19 16 10 9 9 4 3 3 13 1 0 2 11 1 0 11 13 10 9 2
22 15 13 10 11 16 9 7 9 4 4 13 1 10 9 1 9 13 9 7 13 9 2
13 11 13 16 10 11 4 13 10 12 1 11 9 2
21 13 1 10 9 2 11 4 13 1 9 14 13 3 1 10 9 1 11 7 11 2
13 1 12 9 2 10 13 15 4 4 13 1 11 2
21 3 15 13 2 9 13 14 13 1 10 0 9 1 15 7 15 15 7 11 13 2
33 1 11 12 2 4 10 11 9 13 1 10 9 9 11 11 13 1 10 13 9 2 1 12 2 10 4 13 2 11 11 11 2 2
15 10 9 13 14 13 0 9 16 10 0 9 4 14 13 2
16 2 11 11 14 9 13 3 1 11 2 16 13 11 14 2 2
21 9 1 0 9 1 9 7 13 9 1 0 9 13 10 0 9 1 10 11 9 2
28 1 11 12 2 11 11 2 11 11 2 0 2 2 11 11 1 11 11 2 11 11 11 13 1 10 11 11 2
25 15 13 16 9 7 0 9 13 16 11 11 13 14 13 10 11 1 10 0 9 2 3 3 9 2
41 10 0 9 2 10 11 9 13 16 16 15 4 14 13 10 9 1 10 9 1 9 2 15 4 13 9 14 13 1 10 9 13 9 13 1 9 10 4 4 13 2
44 11 11 4 13 9 2 10 0 9 9 1 15 0 9 2 1 3 3 12 2 3 15 4 13 1 11 11 1 10 11 11 11 11 2 2 11 11 2 7 2 11 2 2 2
17 11 2 11 11 14 9 12 2 13 9 1 11 11 14 0 9 2
16 10 11 4 13 1 11 14 9 14 13 9 1 10 0 9 2
27 10 9 7 0 2 9 9 1 11 11 11 13 16 11 13 16 13 9 7 13 14 13 15 1 11 9 2
35 10 0 11 11 9 2 10 9 7 9 2 13 9 9 3 3 2 4 13 1 10 0 9 9 7 15 13 10 9 1 10 13 0 9 2
34 3 11 14 9 1 12 13 16 11 11 7 11 13 0 14 13 1 10 0 7 0 9 15 13 13 10 9 9 0 11 11 9 13 2
39 10 3 13 9 15 4 13 10 0 9 1 11 13 16 11 13 10 9 7 4 13 12 0 9 14 13 10 0 9 14 13 9 1 11 7 10 11 11 2
29 10 11 11 9 4 14 13 2 7 13 10 0 11 9 1 9 13 4 14 13 10 9 13 15 1 10 9 9 2
34 15 13 0 9 1 10 9 1 10 11 9 10 4 13 2 3 1 9 1 10 9 16 9 4 14 3 13 14 4 13 0 1 12 2
39 3 2 10 0 15 13 15 3 10 0 9 3 2 3 0 2 2 16 4 13 2 4 14 3 13 16 15 3 13 10 0 9 1 10 9 1 11 11 2
25 11 11 11 1 10 0 9 1 10 9 1 12 13 16 10 11 4 13 10 11 9 1 12 9 2
47 1 9 12 2 11 2 13 1 10 0 11 9 2 13 16 10 11 4 13 10 9 1 9 13 14 4 13 11 10 13 10 9 1 12 1 12 7 4 14 13 1 16 15 4 13 3 2
25 11 11 14 9 9 9 1 11 11 14 9 4 14 13 9 1 0 9 1 10 3 0 0 9 2
27 3 3 13 1 10 0 9 1 9 9 11 11 7 11 11 2 1 10 0 9 2 15 13 10 0 9 2
17 1 10 9 1 10 9 13 1 10 9 2 15 13 10 0 9 2
25 16 3 13 10 9 1 0 9 7 10 12 9 9 2 15 13 9 3 0 1 12 5 12 9 2
14 2 9 4 13 3 0 1 12 9 14 13 0 2 2
10 0 13 1 10 12 9 9 1 0 2
31 15 13 3 0 2 3 2 14 13 10 12 9 9 1 10 9 1 10 0 9 1 1 0 9 0 1 10 9 13 9 2
27 10 2 12 9 2 9 13 1 10 9 1 10 9 1 0 9 1 10 9 13 16 9 9 4 3 13 2
41 10 13 9 1 11 13 10 9 1 7 10 2 13 11 2 9 7 10 9 0 1 11 11 11 15 13 1 11 9 9 16 15 13 15 16 13 0 1 0 9 2
23 11 9 11 11 3 13 15 2 1 0 9 2 1 11 14 9 16 13 7 13 10 9 2
24 11 11 3 13 9 16 11 11 14 9 1 9 9 4 4 13 1 11 11 14 9 9 9 2
37 16 10 9 1 10 9 1 11 14 9 4 2 7 4 14 2 13 1 0 9 1 0 9 2 15 13 3 0 1 10 9 13 1 10 9 9 2
9 11 11 13 7 10 9 7 9 2
18 11 2 13 0 9 11 11 13 1 12 9 7 12 9 1 11 12 2
19 11 13 10 9 1 11 11 7 10 9 1 11 11 2 2 11 2 2 2
8 11 13 9 1 10 11 11 2
16 11 13 15 9 13 11 11 11 14 13 9 0 1 11 11 2
14 2 9 13 2 11 2 7 11 11 14 0 9 2 2
33 11 11 2 15 13 10 9 9 9 3 15 4 13 2 13 1 11 14 9 1 12 3 15 4 13 14 13 1 9 9 1 11 2
24 11 11 13 11 1 10 9 13 16 15 13 10 9 9 1 11 11 7 3 13 15 5 12 2
14 10 9 9 13 14 13 9 1 10 2 0 9 2 2
25 1 12 2 11 11 13 1 11 7 11 14 13 1 10 11 11 11 7 14 13 15 9 1 9 2
36 16 13 1 11 11 2 10 0 9 1 10 11 11 3 4 4 13 11 2 16 13 15 2 16 13 1 11 1 11 12 2 13 15 1 0 2
16 10 9 4 13 9 1 11 7 13 1 15 9 14 13 9 2
12 11 4 13 1 11 12 1 15 9 1 11 2
30 11 13 16 10 2 0 9 2 13 0 9 4 4 13 1 10 9 1 11 11 9 15 4 4 13 14 13 0 9 2
38 0 9 2 7 0 7 0 2 4 13 1 11 11 9 7 9 2 14 13 10 9 11 11 11 2 10 9 1 11 7 11 11 2 9 2 1 11 2
18 9 11 11 11 4 13 1 1 15 9 2 11 2 16 13 10 9 2
25 1 1 11 12 2 12 2 15 13 1 10 9 1 10 0 9 7 4 4 13 2 0 9 2 2
36 7 10 15 13 1 1 10 9 13 10 9 1 10 9 11 11 11 2 15 13 10 9 1 10 11 16 13 3 0 2 9 1 1 9 9 2
20 15 13 11 11 15 13 9 1 11 11 2 15 13 10 9 1 11 1 9 2
24 10 0 9 13 16 15 4 13 1 11 16 4 13 1 10 9 1 0 11 7 0 11 12 2
11 16 0 2 3 4 10 9 3 13 1 2
8 3 2 11 13 10 0 9 2
16 10 11 11 7 11 3 13 9 9 1 9 1 10 0 9 2
18 10 11 4 14 3 13 10 11 9 1 11 1 12 9 1 15 9 2
30 16 9 11 11 2 3 9 1 10 11 9 13 2 10 9 13 1 11 11 13 0 16 10 9 13 3 0 0 9 2
26 16 15 13 14 0 14 13 9 1 9 2 11 11 11 7 11 11 4 3 13 11 4 3 4 13 2
4 15 4 13 2
21 15 9 11 3 13 11 7 15 9 16 15 13 1 10 9 1 10 9 1 11 2
18 11 13 1 15 9 1 15 9 14 13 10 9 7 10 9 1 11 2
29 13 1 10 11 9 2 11 11 4 13 16 4 13 1 11 11 11 2 16 15 4 13 1 10 9 14 9 2 2
8 2 11 13 1 10 9 2 2
21 10 9 13 15 4 13 16 4 13 10 9 1 11 11 14 2 11 11 11 2 2
31 10 9 14 9 13 15 16 11 4 14 13 0 9 14 13 1 9 9 1 15 7 10 9 7 13 11 1 10 9 9 2
9 15 13 10 0 11 13 1 15 2
8 11 3 13 10 9 14 9 2
27 3 9 13 0 1 10 9 2 7 10 9 2 11 11 11 2 4 13 1 10 10 11 11 7 11 9 2
25 10 9 14 9 13 15 16 11 13 10 9 1 9 2 7 15 4 14 13 14 13 15 9 2 2
31 15 3 13 10 3 0 9 1 10 2 11 2 9 2 11 2 11 11 11 2 15 11 4 13 14 4 13 7 4 13 2
9 15 9 13 2 11 10 11 2 2
14 10 0 11 9 13 16 11 13 9 1 10 0 9 2
18 15 4 13 1 12 11 9 14 13 2 3 2 3 2 3 2 0 2
23 15 3 13 1 12 7 0 9 1 10 9 1 12 1 11 1 10 11 7 11 13 0 2
25 15 4 4 4 13 1 11 2 11 2 1 1 11 11 2 11 2 15 3 3 4 13 9 9 2
17 10 11 11 3 3 3 13 9 1 0 9 7 3 2 13 9 2
37 1 0 11 12 2 10 11 9 13 16 10 9 1 11 14 7 11 11 14 9 1 9 13 1 9 1 10 13 9 16 13 0 9 0 1 9 2
28 15 4 3 4 13 11 11 11 13 0 16 13 9 14 13 0 9 2 1 10 9 1 9 9 11 11 2 2
13 10 9 11 11 13 14 4 13 0 9 1 11 2
26 15 13 0 14 13 15 9 16 15 13 10 9 16 13 1 10 9 15 4 13 1 10 9 1 11 2
15 10 9 13 0 9 1 11 11 14 9 9 9 1 11 2
26 10 0 9 13 1 11 14 0 9 1 11 4 14 13 10 9 16 11 11 13 10 11 9 1 11 2
12 11 2 3 2 13 10 0 9 1 10 11 2
22 0 0 9 11 11 4 13 16 10 0 0 9 13 11 7 16 11 13 10 11 9 2
38 2 15 9 4 4 13 13 1 10 0 0 9 9 13 1 10 11 1 10 11 9 2 11 2 2 10 11 13 14 13 0 1 0 0 9 9 2 2
20 11 4 13 1 11 1 12 1 10 9 14 13 10 9 9 1 11 14 9 2
34 10 9 13 1 9 1 10 11 2 11 14 0 9 2 13 16 10 9 1 11 11 9 4 13 1 10 0 9 1 11 12 1 11 2
26 13 1 3 3 10 9 2 11 11 13 10 9 1 10 0 9 2 13 14 13 15 0 9 1 9 2
44 12 0 0 9 2 9 13 11 7 11 2 4 13 10 9 14 13 0 1 11 14 9 9 2 13 1 11 11 11 2 9 1 10 11 9 9 1 9 1 10 9 1 11 2
20 15 4 13 16 10 11 13 0 9 1 10 9 7 9 9 13 14 13 9 2
34 10 9 9 4 13 3 0 1 10 9 1 9 7 10 9 11 11 7 11 4 4 4 13 2 13 14 3 13 15 1 2 9 2 2
37 11 3 13 11 11 7 11 14 13 9 9 2 1 9 1 0 9 9 2 1 1 10 9 13 3 1 10 2 11 11 2 1 0 7 9 9 2
12 10 9 4 13 10 0 9 16 13 15 9 2
34 11 11 9 7 9 13 16 10 11 14 9 1 9 1 11 2 11 11 2 11 2 11 2 7 10 11 13 1 10 9 1 10 9 2
36 13 1 10 9 15 13 1 10 9 2 11 11 13 10 0 9 1 9 1 11 9 13 1 9 1 10 9 1 11 12 9 11 11 1 11 2
24 11 11 13 9 1 7 10 11 11 13 10 11 7 11 11 1 9 1 0 9 1 10 9 2
36 1 0 11 12 2 15 4 13 16 10 11 4 13 10 9 9 10 4 13 10 9 1 9 1 0 7 9 9 1 9 16 13 10 0 9 2
31 10 9 7 9 1 11 11 9 2 1 1 11 9 1 11 7 10 11 9 1 11 2 13 0 1 10 9 1 11 11 2
35 1 10 9 1 10 9 1 15 0 9 9 2 15 9 4 13 3 1 10 9 9 1 10 2 0 9 2 9 2 3 15 13 9 2 2
31 15 13 0 14 13 1 1 10 9 1 12 9 9 2 9 9 2 7 9 9 1 9 1 11 7 11 7 3 3 11 2
20 10 9 13 1 9 1 10 0 9 1 9 1 9 13 1 10 9 1 11 2
8 11 11 13 10 9 1 9 2
55 1 15 9 12 9 13 11 1 10 11 1 10 11 2 11 13 16 10 0 9 4 13 2 9 2 1 10 0 9 2 14 13 10 9 16 10 0 9 13 3 10 9 1 10 11 11 1 9 16 13 10 11 1 11 2
32 11 13 3 16 15 4 13 0 1 10 9 1 11 11 1 11 1 1 10 11 11 11 7 10 13 9 9 1 11 7 11 2
32 10 9 9 4 13 1 10 9 1 10 11 11 11 7 3 10 9 11 11 4 13 16 16 14 13 10 9 1 9 13 9 2
38 0 1 10 2 13 9 2 1 9 2 3 2 13 3 16 11 7 11 13 0 9 7 4 14 13 9 1 11 11 16 15 15 13 1 10 11 9 2
15 10 11 14 9 13 10 11 2 13 9 1 10 0 9 2
16 11 11 11 13 16 10 2 7 2 7 2 9 13 14 0 2
35 10 9 4 13 14 13 10 9 16 3 10 11 13 10 9 2 9 2 10 9 13 10 11 2 13 2 3 2 0 9 1 10 0 9 2
39 15 13 10 13 9 16 9 4 13 1 10 9 1 11 2 10 9 1 10 11 11 2 1 10 0 9 9 1 11 11 13 10 11 1 11 7 13 9 2
41 10 9 1 10 11 1 11 11 1 9 1 11 9 2 3 3 1 0 9 1 9 11 11 2 13 10 9 16 15 13 3 12 2 7 12 2 0 9 13 9 2
21 2 10 9 13 1 0 11 9 2 12 1 10 11 11 7 10 1 10 11 2 2
20 2 9 9 11 11 13 10 9 13 10 9 14 4 4 13 1 10 11 2 2
23 10 9 1 9 13 14 3 10 9 9 1 10 0 9 13 1 11 2 15 13 15 9 2
20 10 9 13 9 9 1 11 12 1 9 9 1 11 11 11 7 11 2 11 2
26 15 4 13 1 9 1 10 0 9 1 10 11 11 11 7 10 9 1 10 0 9 2 11 11 11 2
29 10 0 9 1 10 0 11 2 11 11 2 11 2 2 11 11 2 2 2 15 13 3 10 0 9 1 11 11 2
27 10 9 9 4 13 1 9 1 10 9 1 10 0 9 13 1 10 0 9 1 10 11 7 10 0 9 2
19 10 9 1 10 9 9 2 10 13 1 0 9 2 13 14 13 10 9 2
30 2 15 3 13 10 0 5 12 12 9 2 1 10 9 1 9 9 2 10 9 3 13 3 1 5 12 12 2 2 2
7 15 13 10 9 1 9 2
5 15 13 10 9 2
20 16 12 4 4 13 2 10 0 9 2 13 1 12 0 9 2 4 3 13 2
3 13 0 2
24 12 9 4 3 13 1 11 2 3 10 0 11 12 9 4 13 2 13 1 2 9 9 2 2
8 2 10 9 4 14 13 2 2
14 11 11 14 9 4 13 1 11 2 11 1 9 12 2
19 10 9 1 9 13 1 10 0 9 1 11 11 2 11 11 14 9 12 2
16 11 3 4 13 1 10 9 1 10 0 9 11 11 11 11 2
18 1 1 11 2 11 11 7 15 12 9 4 13 0 9 1 11 11 2
7 15 3 13 15 1 9 2
43 16 16 1 9 1 10 0 9 2 11 13 0 9 16 13 10 0 9 14 9 14 13 10 9 1 10 0 11 11 7 10 0 11 11 2 11 7 11 13 11 14 9 2
11 10 13 11 12 9 11 13 11 14 9 2
32 3 2 10 9 1 9 1 11 11 14 9 9 9 13 10 0 9 1 15 13 1 9 1 10 0 9 1 10 11 11 11 2
46 13 1 10 0 2 11 9 2 2 10 13 13 9 13 10 0 5 11 11 9 2 11 11 11 4 13 0 9 1 0 9 16 13 9 9 10 0 9 16 10 11 11 9 4 13 2
28 3 16 11 11 13 15 9 9 7 10 0 14 13 0 4 14 13 15 4 14 13 10 9 1 10 0 9 2
12 16 11 11 3 13 2 2 9 13 9 2 2
28 10 9 13 14 13 0 13 9 1 7 0 12 7 0 12 1 11 11 7 9 1 9 9 1 11 1 12 2
16 15 13 3 10 9 13 2 11 11 2 1 10 11 11 9 2
17 10 2 0 9 2 9 13 1 10 9 9 13 10 9 2 9 2
22 15 4 3 13 1 10 0 9 16 9 13 1 9 2 1 10 9 1 0 9 2 2
50 1 10 0 9 1 10 15 13 12 2 7 13 10 9 13 1 10 12 9 1 10 9 2 10 9 13 1 10 11 9 2 10 9 16 13 10 9 12 2 7 13 10 9 1 10 2 0 9 2 2
16 11 11 11 3 13 10 9 1 15 9 2 10 11 11 2 2
23 10 9 1 10 11 11 9 13 16 2 1 10 9 1 0 9 2 13 16 15 13 3 2
23 10 9 14 9 1 2 11 11 2 1 10 9 9 1 10 9 1 10 9 13 3 0 2
33 10 11 12 9 10 11 13 1 0 11 11 9 3 13 16 11 13 2 9 2 1 10 9 9 1 10 0 0 9 1 15 9 2
11 9 13 11 7 13 10 11 11 14 9 2
26 1 11 11 2 10 9 9 4 13 0 2 3 16 11 11 4 13 0 16 13 15 9 11 11 11 2
9 2 9 2 13 2 9 9 2 2
20 11 3 13 1 0 9 9 2 8 2 11 14 0 11 11 7 10 11 11 2
44 10 9 3 4 13 16 15 13 1 7 0 11 11 2 0 11 11 7 11 2 11 11 2 10 13 3 10 0 9 1 10 9 1 10 9 1 10 0 11 11 7 11 11 2
22 1 10 11 9 3 9 13 2 9 4 13 0 9 2 1 1 11 3 15 4 13 2
30 1 10 11 10 11 1 11 13 16 10 9 1 10 9 13 1 10 9 1 0 9 10 13 3 15 13 1 10 9 2
37 1 1 9 2 16 3 13 2 15 13 10 9 1 2 0 9 2 9 1 0 11 11 7 0 11 11 7 0 11 11 1 10 11 11 7 11 2
23 10 0 9 3 13 1 10 13 9 15 4 4 13 7 15 13 1 0 7 4 4 13 2
22 11 14 9 1 10 11 11 1 12 13 14 13 9 1 9 2 3 9 1 0 9 2
18 15 13 1 10 9 7 4 13 1 10 0 11 11 9 13 11 11 2
12 10 9 3 4 15 13 7 15 4 15 13 2
13 10 15 0 9 2 10 11 7 11 13 15 9 2
10 15 13 2 3 3 2 1 15 3 2
29 3 2 10 9 1 10 10 9 13 16 15 13 0 9 14 3 2 13 2 7 3 13 2 15 10 11 4 13 2
16 9 9 13 10 0 9 1 9 1 1 10 9 1 0 9 2
8 3 2 9 13 12 2 12 2
38 3 2 16 10 2 0 9 2 11 11 2 11 1 9 1 10 9 2 15 13 14 0 15 4 13 3 16 13 10 0 9 1 0 9 7 0 9 2
19 3 2 10 2 11 9 2 13 14 4 4 13 7 3 3 13 0 9 2
14 10 2 11 9 2 13 11 11 11 13 3 3 0 2
21 10 9 4 13 1 0 0 9 2 7 15 13 10 0 3 13 9 13 15 9 2
31 10 11 14 9 1 11 2 3 3 16 13 1 10 9 2 4 4 13 1 10 9 1 12 9 16 9 13 1 10 9 2
26 11 14 9 1 9 3 13 1 10 0 9 16 10 0 2 9 13 0 16 12 0 9 4 4 13 2
34 10 11 9 2 14 13 0 9 7 0 12 2 12 9 1 12 9 9 2 13 3 10 9 1 0 0 9 7 9 9 1 0 9 2
18 10 9 1 10 11 11 11 7 9 11 11 4 13 1 0 11 12 2
18 10 9 4 13 14 13 10 0 9 9 1 9 1 3 3 11 12 2
45 10 9 2 13 1 10 0 9 1 9 2 13 16 10 9 13 10 13 9 10 4 13 10 0 9 14 13 2 7 10 9 4 13 16 10 9 14 13 10 9 1 10 9 2 2
25 10 11 9 3 4 3 4 13 1 10 11 11 9 2 1 10 0 0 9 13 1 10 0 9 2
43 13 10 0 9 16 15 13 1 9 2 15 13 3 0 16 10 11 13 1 0 9 10 9 16 11 11 4 3 4 13 1 10 9 16 7 3 15 13 14 13 10 9 2
22 10 9 1 11 11 11 14 9 3 4 13 3 3 10 0 9 1 10 9 9 9 2
26 0 9 4 4 13 1 10 9 16 13 16 10 9 13 1 10 9 16 13 15 3 3 16 13 15 2
2 11 2
30 11 4 13 14 13 1 10 9 1 9 13 1 10 0 9 2 11 9 9 2 12 0 9 16 15 13 15 1 15 2
43 15 4 13 0 16 15 4 14 13 9 7 9 2 9 2 9 2 8 2 9 3 3 12 1 10 9 4 3 4 13 1 10 9 9 7 14 13 10 9 9 4 13 2
20 3 2 15 13 7 9 7 9 1 15 2 7 10 9 4 14 3 4 13 2
16 15 13 16 15 4 13 15 10 9 9 16 13 10 0 9 2
23 1 3 2 15 13 10 9 1 9 1 10 15 4 3 13 10 9 7 2 7 9 9 2
10 15 4 13 10 9 1 11 3 9 2
1 11
1 11
1 11
1 11
1 11
1 11
1 11
14 11 11 9 3 2 15 13 0 9 9 2 3 3 2
1 11
6 11 15 13 0 9 3
6 11 15 13 0 9 3
3 11 9 3
29 15 13 14 0 1 10 9 1 10 11 9 2 9 9 7 4 13 10 9 1 15 16 15 4 14 13 3 3 2
2 9 2
1 11
4 11 7 11 2
23 6 13 15 10 9 1 10 9 10 15 4 13 14 13 15 0 9 1 10 11 9 9 2
2 9 2
1 11
2 11 2
9 15 13 14 13 10 9 1 9 2
8 15 13 3 0 9 3 3 2
2 11 11
2 0 11
41 3 10 0 9 14 13 1 1 10 9 10 15 13 15 3 13 15 14 13 1 15 0 9 2 11 12 11 2 10 4 13 9 1 11 1 12 7 12 11 12 2
11 4 15 13 10 9 14 13 10 9 3 2
35 15 4 13 14 13 10 9 13 0 9 2 3 15 4 3 13 14 13 3 3 16 0 16 15 4 13 0 14 13 1 10 9 14 9 2
32 15 4 13 1 15 11 11 9 1 10 9 3 2 9 2 12 12 12 2 2 7 15 4 4 13 1 9 3 7 1 9 2
3 0 9 2
1 11
16 11 11 9 9 11 11 11 12 12 12 12 12 12 12 12 8
22 11 4 13 15 9 1 10 0 9 11 9 2 12 2 1 11 14 11 11 1 12 2
9 13 15 10 3 2 15 13 3 0
1 11
2 11 2
4 9 10 9 2
7 4 15 13 1 10 9 2
1 11
22 11 4 13 15 9 1 10 11 11 11 9 2 12 2 1 11 14 11 11 1 12 2
9 13 15 10 3 2 15 13 3 0
1 11
1 3
1 11
9 11 2 11 4 13 15 13 11 2
2 11 2
27 16 15 13 1 15 9 9 2 11 11 13 14 13 11 11 2 10 0 9 9 1 11 2 1 15 9 2
16 3 2 3 15 4 13 1 10 9 2 11 13 11 1 11 2
28 11 14 9 13 0 9 2 7 15 13 16 11 4 14 13 10 9 2 7 3 4 14 13 16 11 4 3 2
7 0 9 13 3 0 9 2
45 15 13 16 15 13 11 7 11 14 9 2 9 1 0 0 9 1 15 9 0 1 11 11 7 11 14 13 16 15 13 0 2 7 16 15 9 1 9 7 9 13 14 3 0 2
30 16 10 0 13 10 9 2 15 4 13 7 11 7 11 1 10 9 9 9 2 10 9 9 13 12 5 12 12 2 2
3 6 13 2
2 9 2
1 11
2 11 2
4 9 10 9 2
6 15 13 10 15 9 2
1 11
2 11 2
3 0 9 2
22 11 14 9 4 13 3 2 15 4 13 9 13 1 15 7 13 15 10 9 1 11 2
10 15 13 2 10 2 0 9 1 11 2
33 15 13 5 12 1 0 9 10 9 2 10 9 9 11 4 13 11 1 15 0 9 2 13 10 9 10 4 14 4 13 1 9 2
6 15 13 0 1 15 2
1 11
2 11 2
2 9 2
11 11 2 6 2 13 10 9 1 11 14 9
1 11
2 11 2
7 9 16 13 10 9 3 2
22 15 4 13 9 1 9 16 15 4 13 0 9 9 10 15 4 14 13 9 1 3 2
47 0 1 15 9 1 0 9 1 10 9 4 13 16 15 13 10 0 9 2 13 15 14 13 1 11 11 2 11 2 7 11 2 7 13 14 13 1 15 9 14 0 9 9 1 9 0 2
10 10 0 9 13 10 9 1 15 3 2
33 16 15 4 13 9 0 1 9 1 0 9 7 9 9 2 7 0 9 1 0 9 9 7 0 9 1 10 9 2 15 4 13 2
1 11
2 11 2
14 15 4 13 10 9 3 7 13 1 15 1 0 9 2
29 1 10 9 2 15 4 13 14 13 1 10 9 9 1 0 9 2 3 1 9 7 10 0 9 16 10 9 13 2
20 11 11 9 9 9 11 11 11 11 2 11 12 12 9 9 2 12 9 2 12
2 11 2
4 13 10 9 2
18 3 2 1 15 0 9 2 15 4 14 13 14 3 13 1 10 9 2
30 15 13 11 4 13 14 13 9 0 2 7 16 9 15 13 14 2 15 4 14 13 14 13 12 5 1 15 9 9 2
24 15 4 9 9 16 3 15 4 13 14 13 1 9 1 11 7 4 13 9 14 13 10 9 2
15 1 10 9 2 15 13 15 4 14 13 14 13 0 9 2
18 15 4 13 10 9 1 9 14 13 10 9 15 13 1 0 0 9 2
7 6 13 1 15 1 15 2
2 11 2
2 11 2
24 15 4 13 1 10 0 9 1 11 7 13 15 4 13 10 9 14 13 1 10 9 15 13 2
21 3 3 2 15 4 3 13 1 10 9 14 13 9 3 16 10 9 13 10 9 2
17 15 13 14 0 16 11 1 12 13 10 9 2 7 3 1 12 2
7 13 15 16 15 13 0 2
20 11 11 9 9 9 11 11 11 11 2 11 12 12 9 9 2 12 9 2 12
27 9 13 9 1 9 7 9 2 6 4 14 13 9 7 2 7 9 13 15 11 9 2 8 2 1 9 2
30 9 7 2 7 9 13 1 9 4 14 4 13 1 11 7 11 4 14 13 0 16 13 1 0 9 7 2 7 9 2
29 9 13 9 7 9 2 11 13 10 9 14 13 7 13 10 9 1 10 9 9 13 7 2 7 13 1 15 9 2
27 9 13 9 1 9 7 9 2 6 4 14 13 9 7 2 7 9 13 15 11 9 2 8 2 1 9 2
30 9 7 2 7 9 13 1 9 4 14 4 13 1 11 7 11 4 14 13 0 16 13 1 0 9 7 2 7 9 2
29 11 13 9 7 9 2 11 13 10 9 14 13 7 13 10 9 1 10 9 9 13 7 2 7 13 1 15 9 2
27 9 13 9 1 9 7 9 2 6 4 14 13 9 7 2 7 9 13 15 11 9 2 8 2 1 9 2
30 9 7 2 7 9 13 1 9 4 14 4 13 1 11 7 11 4 14 13 0 16 13 1 0 9 7 2 7 9 2
29 9 13 9 7 9 2 11 13 10 9 14 13 7 13 10 9 1 10 9 9 13 7 2 7 13 1 15 9 2
3 15 13 2
12 6 13 16 0 3 15 9 9 4 13 1 8
6 15 3 13 1 11 2
8 3 1 9 1 11 1 15 2
6 15 9 11 13 15 2
11 3 1 0 1 15 7 1 15 1 11 2
3 14 3 2
6 3 13 9 1 11 2
11 4 15 13 1 10 11 9 9 9 11 2
7 6 11 13 15 10 9 2
6 4 9 11 13 3 2
3 14 3 2
6 3 13 9 1 11 2
11 4 15 13 1 10 11 9 9 9 11 2
7 6 11 13 15 10 9 2
7 11 4 14 13 1 15 2
8 3 1 11 1 12 11 9 2
4 15 3 13 2
38 15 4 13 14 13 10 9 3 10 9 1 12 5 12 9 1 10 12 1 15 3 14 13 0 15 4 13 3 7 14 13 10 9 7 9 7 9 2
15 15 0 9 13 16 15 13 10 9 3 1 15 0 9 2
6 15 4 15 9 13 2
1 11
2 6 2
11 15 4 13 14 13 15 0 9 1 11 2
7 11 13 0 9 1 12 2
7 11 4 14 13 1 15 2
8 3 1 11 1 12 11 9 2
4 15 3 13 2
38 15 4 13 14 13 10 9 3 10 9 1 12 5 12 9 1 10 12 1 15 3 14 13 0 15 4 13 3 7 14 13 10 9 7 9 7 9 2
15 15 0 9 13 16 15 13 10 9 3 1 15 0 9 2
6 15 4 15 9 13 2
1 11
3 14 3 2
9 4 15 13 14 13 15 9 9 2
6 6 13 1 9 3 2
2 9 2
8 11 11 4 13 10 13 9 2
16 15 13 0 1 10 9 1 9 2 1 0 2 11 11 11 2
28 16 15 4 2 6 13 10 0 9 7 13 15 13 16 15 13 1 9 1 10 9 1 9 9 2 16 0 2
10 15 13 1 9 16 15 13 10 9 2
2 9 2
45 15 13 10 1 10 9 2 3 2 10 9 13 16 15 13 11 2 10 15 4 16 15 4 14 13 12 12 5 12 12 2 2 15 4 13 1 13 10 9 1 12 5 12 9 2
8 15 13 3 0 9 1 15 2
20 15 13 15 13 1 10 9 2 7 10 9 1 0 9 13 3 0 3 3 2
9 15 4 13 14 13 15 13 3 2
2 9 2
15 15 4 13 10 9 1 10 9 9 9 1 11 11 11 2
21 11 13 10 9 1 15 7 3 13 10 9 4 13 14 13 15 14 13 10 13 2
5 0 9 2 5 12
4 9 9 2 9
5 9 9 9 2 0
3 9 9 2
4 9 9 12 9
3 12 9 9
3 5 12 9
3 13 9 2
5 9 9 2 12 12
3 12 9 9
3 5 12 9
41 9 9 2 16 15 13 0 12 12 7 12 12 15 4 3 13 10 1 10 5 12 9 2 3 12 5 2 7 13 1 9 15 4 13 1 0 1 10 0 9 2
15 3 2 10 9 1 10 0 9 1 10 9 13 12 9 2
19 15 4 3 13 15 9 14 13 1 10 0 9 9 4 15 14 4 13 2
36 3 2 15 4 3 8 13 9 10 15 13 1 10 0 9 9 10 13 0 7 0 9 3 8 11 11 2 11 11 2 11 11 7 11 11 2
6 11 11 1 11 11 2
5 11 11 0 5 12
5 11 11 0 5 12
5 11 11 0 5 12
5 11 11 0 5 12
5 11 11 0 5 12
14 13 15 13 15 9 2 3 15 4 13 15 1 11 2
6 4 15 13 14 13 2
17 9 9 7 11 1 11 11 11 12 5 12 2 12 2 11 2 11
1 9
39 10 9 4 13 10 9 7 0 9 1 11 0 9 1 9 16 3 13 9 9 14 13 0 9 1 10 0 7 0 0 0 9 13 1 11 14 11 9 2
15 10 9 4 13 10 9 1 10 9 7 0 9 1 15 2
13 15 4 13 9 9 7 0 9 9 1 9 9 2
25 15 4 13 13 9 1 0 9 9 7 9 2 13 9 2 13 9 9 1 11 14 0 9 9 2
34 10 9 4 3 13 15 15 4 13 1 0 9 7 0 9 14 13 10 0 9 16 13 16 10 9 13 10 0 9 7 0 9 9 2
24 10 9 1 10 11 7 0 11 4 4 13 16 13 1 10 9 3 2 2 8 2 2 8 2
14 9 11 11 11 11 12 5 12 2 12 2 11 2 11
12 15 13 14 13 9 1 12 14 12 9 9 2
10 15 13 10 12 9 9 9 1 12 2
1 11
2 11 11
3 12 12 9
9 2 13 9 2 9 0 9 2 2
17 15 13 16 15 13 1 15 16 15 4 14 13 10 1 10 9 2
3 15 2 11
7 15 2 0 9 1 11 11
6 3 2 9 1 12 9
12 3 2 10 11 11 12 11 11 2 12 2 12
11 3 2 9 13 11 14 0 9 1 11 2
9 15 13 14 10 11 2 13 9 2
10 3 4 15 13 16 13 1 10 9 2
16 11 7 11 4 13 13 9 12 1 15 9 2 13 3 2 2
4 4 15 13 2
7 6 13 15 13 11 9 2
2 9 2
1 11
16 16 15 4 14 3 13 10 9 2 11 14 9 4 13 0 2
7 11 11 0 9 9 11 12
8 6 13 15 9 1 0 3 2
1 11
2 11 2
13 4 15 13 3 10 9 10 13 1 10 0 9 2
17 16 0 2 4 15 3 13 10 9 1 10 9 2 12 1 12 2
2 9 2
1 11
18 15 13 10 0 9 10 4 13 14 13 9 7 4 13 1 10 9 2
6 9 2 11 11 11 11
12 10 9 13 14 1 11 2 11 2 7 11 2
13 10 12 9 9 13 10 9 2 9 2 7 9 2
23 15 13 10 0 9 9 1 10 9 2 7 10 9 13 14 4 13 0 1 15 13 9 2
6 9 2 11 11 11 11
13 1 10 9 2 10 9 13 14 13 10 11 9 2
24 1 11 9 2 10 9 13 3 5 12 12 1 11 7 3 5 12 12 1 9 2 9 0 2
20 10 0 12 9 13 15 9 16 1 11 2 7 4 14 4 13 1 10 9 2
8 9 2 11 11 11 2 11 2
30 10 9 4 13 1 12 1 10 9 1 11 11 2 3 11 11 11 2 11 9 2 2 7 3 13 1 9 1 9 2
17 9 13 3 1 10 0 9 1 9 7 9 2 7 10 9 9 2
5 9 13 15 9 2
9 15 13 10 9 4 13 1 9 2
9 3 15 13 15 4 13 1 11 2
7 15 4 13 12 2 0 2
9 12 2 11 11 11 9 1 9 2
12 10 9 4 3 4 13 1 9 7 9 9 2
8 14 3 1 15 9 1 9 2
24 15 13 15 4 13 1 10 9 2 0 9 2 0 1 9 2 7 9 7 9 2 11 2 2
4 12 2 0 2
6 12 2 11 2 11 11
10 13 1 0 9 14 13 9 9 9 2
7 13 1 10 9 1 12 2
30 10 0 9 2 12 2 4 13 1 9 7 9 2 11 11 7 11 11 2 3 10 9 4 4 13 1 15 3 3 2
4 12 2 0 2
7 12 2 11 2 11 2 11
10 13 1 1 11 11 11 2 10 9 2
16 11 11 11 4 13 1 11 11 2 11 11 7 11 11 2 2
23 3 10 9 4 3 13 1 15 16 10 0 9 10 4 13 14 4 13 4 13 0 9 2
4 12 2 0 2
8 12 2 11 2 11 11 2 11
10 13 1 0 9 14 13 9 9 9 2
7 13 1 10 9 1 12 2
4 0 1 12 2
15 15 4 4 13 1 11 11 2 11 11 7 11 11 2 2
4 12 2 0 2
9 13 15 13 16 15 13 10 9 2
14 11 11 0 9 9 9 7 9 2 12 2 12 9 8
7 10 9 16 13 9 12 3
15 15 13 16 15 13 10 12 2 3 15 4 13 10 9 2
10 3 4 15 13 16 13 1 10 9 2
16 11 7 11 4 13 13 9 12 1 15 9 2 13 3 2 2
4 4 15 13 2
7 6 13 15 13 11 9 2
2 9 2
1 11
16 16 15 4 14 3 13 10 9 2 11 14 9 4 13 0 2
7 11 11 0 9 9 11 12
8 6 13 15 9 1 0 3 2
1 11
2 11 2
13 4 15 13 3 10 9 10 13 1 10 0 9 2
17 16 0 2 4 15 3 13 10 9 1 10 9 2 12 1 12 2
2 9 2
1 11
2 11 2
2 6 2
13 15 4 3 13 16 13 10 11 7 11 0 9 2
15 15 13 15 7 13 10 1 10 9 1 11 2 11 11 2
7 15 4 4 13 10 9 2
12 15 13 0 7 4 13 10 9 1 15 9 2
19 1 10 9 10 11 13 3 7 13 1 15 0 9 9 7 15 13 0 2
11 15 4 3 13 10 11 1 10 0 9 2
7 15 13 0 1 0 9 2
5 3 2 10 9 2
12 15 4 4 13 1 12 7 0 1 10 13 2
31 15 9 13 16 1 9 15 4 13 14 13 12 1 10 10 13 9 7 15 4 3 13 3 15 13 9 10 15 3 13 2
17 15 13 10 1 15 2 3 15 1 15 9 14 9 7 9 2 2
24 15 13 3 3 1 9 9 7 16 15 13 16 15 13 10 9 10 15 13 15 4 13 15 2
6 15 13 13 7 13 2
21 15 13 16 10 4 14 13 1 10 9 7 15 13 10 0 9 1 15 9 9 2
19 15 3 13 16 10 4 14 4 13 10 9 1 9 7 15 13 3 0 2
18 1 9 2 15 4 13 14 13 16 11 7 11 13 10 9 1 9 2
10 3 3 15 13 15 15 4 13 3 2
5 11 2 0 3 2
1 11
8 11 2 10 9 1 9 2 2
9 15 4 14 13 16 15 13 10 2
6 0 0 7 8 0 9
1 11
1 11
1 11
1 11
1 11
1 11
1 11
1 11
28 1 10 9 2 15 13 0 16 13 1 10 11 2 16 15 13 12 2 10 15 9 13 10 9 1 9 3 2
31 15 13 10 0 9 1 10 9 7 15 13 15 13 10 9 10 2 9 9 2 2 9 1 10 9 1 10 0 9 2 2
17 15 13 1 9 1 10 9 1 9 1 11 7 13 3 5 12 2
5 13 15 12 0 2
42 3 15 4 3 13 1 10 11 15 13 3 7 16 15 4 13 2 15 13 10 9 1 0 9 15 13 0 1 7 15 4 13 1 10 0 9 16 15 3 13 12 2
2 9 2
1 11
5 11 13 1 11 2
3 8 8 8
3 12 12 9
6 11 13 2 11 13 2
2 8 8
3 12 12 9
5 9 1 10 9 2
3 11 13 2
9 15 4 13 9 3 9 13 1 2
1 11
3 8 8 8
3 12 12 9
1 11
11 15 13 16 15 4 13 14 13 9 9 2
16 15 4 13 14 13 3 2 15 4 13 15 13 3 10 9 2
29 15 13 3 10 9 7 15 13 14 13 10 0 9 1 10 9 9 3 1 11 9 3 15 4 4 13 1 9 2
30 3 2 15 13 15 13 1 3 0 9 3 15 4 3 4 13 9 7 3 4 14 13 3 0 16 15 13 14 13 2
1 11
52 9 15 9 13 15 15 13 1 12 9 9 2 3 15 13 1 16 12 1 15 13 10 8 9 7 10 9 1 11 2 15 4 14 13 10 9 1 15 2 15 13 15 13 10 3 2 3 0 9 9 9 2
8 11 2 3 13 10 0 9 2
17 6 13 1 10 11 9 7 13 10 9 7 9 10 15 13 0 2
14 15 4 14 3 13 10 9 16 15 3 13 15 3 2
1 11
12 11 2 15 13 15 4 13 10 9 1 15 2
1 11
3 8 8 8
3 12 12 9
1 11
11 15 13 16 15 4 13 14 13 9 9 2
16 15 4 13 14 13 3 2 15 4 13 15 13 3 10 9 2
29 15 13 3 10 9 7 15 13 14 13 10 0 9 1 10 9 9 3 1 11 9 3 15 4 4 13 1 9 2
30 3 2 15 13 15 13 1 3 0 9 3 15 4 3 4 13 9 7 3 4 14 13 3 0 16 15 13 14 13 2
1 11
52 9 15 9 13 15 15 13 1 12 9 9 2 3 15 13 1 16 12 1 15 13 10 8 9 7 10 9 1 11 2 15 4 14 13 10 9 1 15 2 15 13 15 13 10 3 2 3 0 9 9 9 2
8 15 4 13 15 1 15 9 2
15 3 0 15 4 14 13 10 11 9 2 7 3 0 9 2
13 11 11 2 6 10 10 9 9 1 10 0 9 2
10 15 4 13 10 0 9 1 9 3 2
17 15 4 13 10 0 9 16 15 13 11 3 0 9 1 15 9 2
11 15 13 1 10 11 7 13 10 0 9 2
2 8 8
3 12 12 9
26 10 11 2 11 13 1 10 9 1 11 11 2 10 4 13 15 0 9 2 3 3 2 3 0 2 2
6 15 4 13 3 3 12
26 0 11 15 4 13 14 13 14 13 11 3 16 15 13 3 3 3 2 10 13 13 1 12 7 3 2
9 11 12 2 11 9 1 10 9 2
25 11 12 2 12 2 11 13 1 1 9 2 3 15 13 14 13 11 3 1 9 2 13 1 12 2
11 11 12 2 12 2 13 14 13 9 9 2
26 11 13 10 9 1 11 11 2 3 15 13 1 11 2 11 11 2 11 2 14 3 0 10 9 2 2
14 15 13 10 9 14 9 1 11 2 7 9 4 13 2
13 15 13 15 4 14 13 1 9 1 10 11 9 2
5 13 2 3 3 2
4 9 16 13 2
11 15 4 13 1 10 0 9 9 2 3 2
5 3 2 9 2 9
14 15 13 10 9 1 9 16 15 4 13 1 10 9 2
9 15 13 1 13 9 9 9 9 2
16 4 15 13 14 13 10 0 9 2 7 4 15 13 3 0 2
31 4 15 13 14 13 10 9 1 10 9 9 2 7 13 10 0 9 16 13 1 9 3 10 0 16 15 13 1 10 9 2
19 15 13 10 9 16 10 11 9 9 4 13 15 1 10 9 1 10 9 2
12 4 15 13 14 13 12 9 9 2 7 0 2
23 15 4 13 1 10 9 9 2 10 4 13 1 11 14 9 2 4 14 13 3 3 2 2
14 16 9 13 15 0 2 15 4 13 9 1 1 15 2
2 9 2
1 11
8 13 10 12 7 0 9 9 2
12 15 13 15 13 14 13 0 9 1 10 9 2
14 15 13 10 9 1 9 16 15 4 13 1 10 9 2
9 15 13 1 13 9 9 9 9 2
16 4 15 13 14 13 10 0 9 2 7 4 15 13 3 0 2
31 4 15 13 14 13 10 9 1 10 9 9 2 7 13 10 0 9 16 13 1 9 3 10 0 16 15 13 1 10 9 2
19 15 13 10 9 16 10 11 9 9 4 13 15 1 10 9 1 10 9 2
12 4 15 13 14 13 12 9 9 2 7 0 2
23 15 4 13 1 10 9 9 2 10 4 13 1 11 14 9 2 4 14 13 3 3 2 2
14 16 9 13 15 0 2 15 4 13 9 1 1 15 2
2 9 2
1 11
24 1 10 9 1 10 9 2 10 9 13 16 10 5 12 12 4 13 3 10 9 9 4 13 2
21 4 15 13 16 10 9 0 1 10 9 4 4 13 16 10 0 9 9 4 13 2
2 9 2
1 11
35 8 2 10 9 10 15 4 13 11 13 0 1 11 11 7 4 14 13 0 16 13 10 9 2 8 2 11 4 13 10 9 0 9 2 2
12 3 2 15 13 16 15 13 14 13 10 9 2
13 8 2 10 9 1 10 9 9 13 10 11 9 2
22 1 9 14 13 10 12 9 2 15 4 13 14 13 11 14 13 10 9 9 1 12 2
23 1 15 9 2 15 4 13 11 10 9 1 10 9 1 10 9 16 10 9 9 4 13 2
16 15 4 3 13 15 10 9 9 9 10 9 9 1 10 9 2
23 13 16 3 11 13 2 15 4 13 10 0 9 16 10 9 13 14 4 13 1 10 9 2
12 8 2 15 13 3 3 12 9 9 1 9 2
18 15 4 14 13 14 13 10 9 1 12 9 1 10 9 1 10 9 2
21 9 9 4 7 4 13 1 10 9 9 7 10 9 1 9 9 1 10 13 9 2
4 3 0 9 2
5 13 1 2 8 8
5 3 2 13 3 2
6 11 14 9 13 9 2
8 15 4 15 13 14 13 15 2
1 11
6 15 13 10 0 9 2
9 15 13 15 4 13 15 9 3 2
8 13 3 16 13 10 0 9 2
1 11
9 11 11 2 8 2 1 12 12 9
6 15 9 13 3 0 2
17 15 9 13 3 0 2 3 15 13 9 15 13 14 13 12 9 2
9 3 15 13 15 13 10 9 13 2
18 3 15 4 13 1 10 9 13 9 10 9 13 15 12 9 14 13 2
12 15 13 9 1 9 2 2 5 3 10 9 2
8 15 9 9 13 1 10 9 2
12 3 15 13 1 10 9 10 9 13 15 9 2
10 15 0 9 9 9 13 10 0 9 2
13 15 9 14 9 13 2 9 13 1 0 9 2 2
10 15 13 14 13 15 9 1 10 9 2
13 10 9 1 15 9 13 1 10 9 1 0 9 2
49 15 9 13 3 0 2 10 10 9 1 9 13 9 10 13 2 2 0 9 2 12 9 7 15 9 2 15 9 13 3 0 2 3 15 13 3 2 15 13 14 13 10 12 9 1 10 9 9 2
17 15 9 13 3 0 2 3 1 11 12 9 2 15 13 11 9 2
19 15 9 13 3 0 2 3 15 13 1 10 9 2 15 13 14 13 3 2
17 15 9 13 3 0 2 15 4 13 1 10 9 9 1 15 9 2
16 15 9 13 3 0 2 15 4 13 0 0 9 13 1 15 2
11 15 9 13 3 0 2 15 4 13 9 2
8 15 4 13 14 13 7 13 5
2 0 2
7 13 10 9 1 11 9 2
1 11
7 15 13 10 0 9 9 2
4 13 15 9 2
1 11
27 15 13 11 16 15 13 15 9 3 3 16 15 4 14 13 14 13 15 9 16 15 13 9 13 1 9 2
20 15 13 15 15 13 15 14 13 15 1 7 3 3 13 15 15 13 14 13 2
20 15 13 15 4 13 1 9 7 13 16 15 15 13 15 10 9 13 10 9 2
1 11
10 13 10 9 10 15 13 11 3 0 2
22 10 10 9 1 9 4 13 15 4 14 13 13 15 13 15 4 3 13 10 0 9 2
1 11
3 11 11 12
8 15 4 14 13 1 10 5 2
24 4 15 13 14 9 13 10 9 1 15 9 1 10 9 1 10 9 7 4 15 3 13 15 2
1 11
2 11 2
12 4 14 13 10 9 1 16 15 13 1 15 2
27 15 13 15 13 15 7 15 13 14 13 15 1 10 0 9 9 2 15 3 13 15 1 15 0 9 2 2
2 9 2
1 11
10 3 10 9 14 13 15 10 9 9 2
2 9 2
1 11
5 11 13 15 9 2
16 15 4 13 1 11 1 10 9 1 9 7 4 13 15 3 2
1 11
5 15 4 13 3 2
8 4 14 13 11 7 11 13 2
1 11
12 15 4 14 13 10 9 14 13 1 11 9 2
6 13 15 10 9 9 2
1 11
13 4 15 6 13 10 11 9 2 9 1 15 9 2
1 11
8 3 16 13 1 12 7 12 2
11 15 13 1 10 9 3 13 15 10 9 2
2 11 12
5 10 9 13 0 2
1 11
7 13 13 9 7 9 9 2
8 3 15 4 14 13 9 3 2
9 11 13 3 0 7 10 0 9 2
9 15 13 15 4 13 10 0 9 2
18 13 15 10 9 11 9 14 13 2 13 1 11 13 1 10 9 2 2
2 9 2
1 11
11 15 4 14 13 10 9 14 13 15 3 2
19 11 13 1 1 10 9 9 3 15 4 14 13 10 9 14 13 1 15 2
15 15 4 13 15 3 3 16 15 13 16 15 4 7 14 2
1 11
9 4 15 9 3 13 1 10 9 2
11 4 15 13 10 9 1 11 7 15 3 2
16 11 11 11 11 9 12 2 12 11 11 11 2 11 9 9 12
5 11 11 2 9 12
5 11 11 2 9 12
19 13 4 10 9 1 10 9 1 10 9 1 10 9 2 9 7 9 2 2
20 15 4 13 14 13 10 9 9 1 10 0 9 14 13 3 3 16 15 4 2
1 11
4 13 15 3 2
1 11
3 9 9 2
5 11 11 13 6 2
1 11
7 15 4 13 0 14 13 2
1 11
2 11 11
2 12 12
3 11 2 11
32 3 7 3 2 1 11 11 14 9 2 15 4 13 3 10 12 9 9 9 1 15 0 9 9 2 15 10 12 9 9 2 2
32 15 13 1 10 0 9 1 10 9 2 3 15 13 10 9 9 1 11 10 4 13 15 1 9 1 11 2 10 11 11 9 2
10 13 15 10 9 1 9 7 9 9 2
1 11
5 0 11 13 0 2
43 11 4 13 10 9 1 0 9 1 10 9 1 11 2 11 11 11 11 11 2 0 9 10 15 7 15 13 0 14 13 1 2 2 10 11 11 7 10 9 9 1 11 2
18 15 13 16 15 13 12 9 1 10 9 2 11 12 2 12 7 9 2
22 3 10 0 9 1 11 4 13 3 2 7 15 4 13 10 9 1 0 9 2 2 2
6 4 15 13 1 15 2
13 7 4 15 13 14 13 15 1 10 11 7 11 2
22 11 3 13 3 1 15 2 3 16 16 15 13 3 1 11 7 13 9 1 11 9 2
2 6 2
10 13 1 10 0 9 2 9 2 9 2
8 15 13 10 9 4 13 0 2
7 15 13 10 0 9 11 2
8 3 4 0 11 13 1 15 2
7 4 15 13 10 9 3 2
6 4 15 13 1 9 2
1 11
38 15 13 16 15 13 10 0 9 14 13 10 9 13 15 0 9 9 2 7 15 13 1 10 3 0 9 2 0 1 10 0 9 7 10 9 1 9 2
22 1 10 9 1 9 2 15 13 14 0 1 15 9 16 7 3 15 3 13 10 9 2
36 13 15 10 9 14 4 13 1 10 11 9 7 1 9 10 9 14 4 13 1 11 14 9 2 16 3 2 1 15 4 10 9 4 13 2 2
19 7 13 10 9 1 11 10 9 14 4 13 1 10 9 9 1 10 9 2
44 1 9 1 10 0 9 2 15 13 16 12 1 10 0 9 1 0 9 9 13 16 15 4 13 14 13 0 1 9 2 13 1 10 9 7 10 9 3 15 13 1 9 9 2
37 16 10 9 9 13 3 2 15 4 13 1 9 9 16 9 4 4 13 7 15 4 13 0 14 13 11 9 9 16 15 13 9 1 9 9 3 2
25 10 0 9 3 4 13 11 14 13 15 9 9 3 3 2 1 3 13 9 1 9 1 9 9 2
19 15 13 14 0 1 10 9 16 13 16 10 0 9 1 10 9 13 3 2
7 3 2 10 9 13 9 2
42 10 0 15 13 16 15 7 11 13 10 9 9 1 0 9 9 13 16 15 4 4 13 2 11 13 15 14 13 1 11 14 9 1 11 2 1 9 1 10 9 9 2
30 15 4 14 13 16 15 13 3 1 10 9 3 15 4 13 16 10 9 9 3 4 13 2 13 7 4 13 10 9 2
36 7 3 14 13 10 9 16 13 10 9 2 10 0 9 2 7 10 0 9 1 15 2 4 13 10 0 9 9 1 10 0 9 1 10 9 2
22 15 9 1 11 11 13 16 15 4 13 10 0 9 1 9 1 10 9 1 10 9 2
32 15 13 0 9 14 13 16 13 10 9 7 9 1 10 9 7 3 0 9 14 13 14 13 0 9 1 9 16 13 10 9 2
23 11 4 13 11 11 14 13 1 15 2 7 15 13 16 11 4 3 4 13 1 11 11 2
22 3 15 13 16 7 3 15 13 14 13 9 1 0 9 10 15 4 14 3 13 1 2
40 4 10 3 0 9 13 1 10 11 11 11 9 1 11 3 15 4 13 0 9 2 9 7 9 1 10 9 7 2 3 2 15 0 9 1 10 0 9 9 2
8 0 16 10 9 13 3 0 2
17 15 4 4 13 12 9 16 13 2 3 15 13 16 15 13 9 2
7 9 16 13 15 1 15 2
19 16 15 13 1 9 2 15 13 16 15 4 14 13 16 15 13 15 10 2
2 2 11
3 8 8 8
3 12 12 9
31 11 2 15 13 16 15 9 1 12 1 12 4 13 3 1 12 5 9 1 9 2 8 2 5 12 12 1 5 12 12 2
32 15 4 13 0 14 13 11 14 0 9 9 0 9 1 9 2 15 4 13 3 14 13 10 0 9 0 9 1 9 3 3 2
16 4 15 13 10 9 16 3 15 4 13 0 14 13 10 9 2
1 9
1 11
14 4 14 13 1 15 2 0 16 13 15 3 1 9 2
15 15 3 13 11 14 13 2 15 13 9 9 3 3 2 2
8 9 1 10 9 1 10 9 2
28 1 10 9 15 4 14 13 10 0 9 4 4 13 3 3 2 9 13 11 16 13 2 16 1 0 9 2 2
9 10 0 9 9 4 3 13 0 2
17 11 11 4 13 10 9 2 9 14 0 14 13 15 16 15 13 2
2 11 11
5 13 1 2 11 11
3 12 12 9
7 15 13 16 15 13 9 2
20 6 13 15 13 16 15 4 3 13 10 9 1 10 0 2 13 9 1 11 2
8 9 16 13 10 9 1 15 2
17 15 13 10 0 9 1 10 9 2 15 13 3 3 16 15 13 2
2 0 2
1 11
22 4 15 13 10 9 16 13 12 2 1 2 12 7 4 15 3 13 1 10 0 9 2
21 15 13 0 16 16 15 4 3 13 10 9 1 9 1 9 15 4 13 15 9 2
2 11 11
5 13 1 2 11 11
3 12 12 9
50 13 10 0 9 2 15 4 3 13 14 13 1 10 9 1 11 2 7 4 13 10 0 9 13 16 2 1 0 2 15 13 14 13 3 1 10 9 7 13 14 13 11 13 10 9 10 13 1 9 2
2 6 2
3 13 3 2
10 4 15 13 10 9 1 10 11 9 2
2 11 11
3 12 12 9
2 11 2
23 1 10 9 2 15 9 9 4 13 10 9 7 13 15 4 13 10 9 7 9 9 9 2
9 15 13 3 12 0 9 2 3 2
11 9 3 4 14 13 16 13 9 1 9 2
25 15 13 16 9 13 1 11 7 13 1 10 0 11 9 4 14 13 10 9 9 1 10 11 9 2
27 10 9 4 13 10 11 9 16 11 13 3 14 13 15 0 9 9 9 2 11 2 7 4 13 11 3 2
15 11 4 13 1 11 2 16 15 4 13 1 10 0 9 2
25 9 2 13 14 13 10 0 9 1 10 9 2 4 14 13 11 16 9 9 4 14 4 13 0 2
14 9 4 3 13 10 9 13 11 10 4 13 0 9 2
33 9 4 14 4 13 3 1 10 9 1 10 0 9 2 7 4 15 4 13 1 12 1 12 9 16 15 4 13 1 10 9 9 2
40 10 9 14 13 13 16 10 9 4 13 0 14 13 7 13 1 10 13 9 1 9 2 13 9 4 14 13 15 7 13 15 3 2 16 15 4 1 9 2 2
32 15 13 16 15 4 13 3 1 10 9 1 0 9 7 13 10 9 3 2 16 15 4 4 13 7 13 1 10 9 15 13 2
21 10 0 9 13 16 10 0 9 1 9 4 13 10 9 2 7 15 13 0 9 2
27 15 4 13 11 4 13 10 9 1 10 9 10 4 13 15 14 3 13 10 9 16 13 15 9 2 3 2
10 6 13 15 13 16 15 13 0 9 2
2 2 11
3 11 11 11
3 12 12 9
22 4 15 13 10 9 1 3 0 15 4 13 2 3 0 15 4 14 7 3 15 13 2
18 13 0 9 2 8 11 2 0 7 13 15 3 10 15 13 9 9 2
2 11 11
3 12 12 9
4 11 7 11 2
20 11 11 7 15 4 13 14 13 1 15 14 13 10 9 13 11 16 15 13 2
14 16 15 4 13 1 10 9 9 2 15 13 3 0 2
2 9 2
1 11
1 9
2 8 8
5 13 1 2 8 8
3 12 12 9
23 11 11 4 13 15 14 13 10 9 9 14 13 10 11 9 10 4 13 11 2 11 9 2
12 6 4 13 16 15 4 13 10 9 16 13 2
6 9 2 11 2 11 9
12 9 2 12 9 2 12 9 11 2 12 9 11
5 13 1 9 2 12
4 9 9 2 12
8 9 9 1 11 11 3 2 12
10 16 15 13 10 9 2 6 13 12 2
6 11 11 9 1 11 11
4 15 13 3 9
12 15 13 4 15 13 15 9 1 9 0 9 2
13 10 9 9 13 12 2 3 4 14 15 13 15 2
18 4 15 13 10 9 1 11 11 11 13 12 9 1 11 9 1 12 2
15 15 4 13 1 15 7 15 4 14 13 10 9 1 15 2
9 4 15 13 15 10 11 9 9 2
1 9
1 11
11 0 14 13 1 15 7 15 9 2 11 2
10 15 4 13 10 0 0 11 11 9 2
8 0 9 1 9 9 1 12 2
10 16 15 13 10 0 9 2 6 13 2
12 3 2 15 4 13 15 4 13 10 12 9 2
3 13 15 2
18 3 2 1 0 9 10 9 9 13 12 2 3 4 14 15 13 15 2
18 4 15 13 10 9 1 11 11 11 13 12 9 1 11 9 1 12 2
15 15 4 13 1 15 7 15 4 14 13 10 9 1 15 2
9 4 15 13 15 10 11 9 9 2
1 9
1 11
4 4 13 8 9
19 11 2 1 9 12 1 11 12 9 1 11 11 2 15 13 10 9 9 2
19 15 9 13 9 9 9 7 11 4 13 14 13 15 13 1 9 9 9 2
17 4 15 6 13 10 9 13 0 7 13 10 9 1 11 16 0 2
1 9
23 11 11 11 11 11 11 9 9 9 2 2 12 2 12 9 2 2 12 2 12 9 2 8
5 0 1 10 9 2
8 13 15 7 15 9 13 3 2
10 13 4 10 9 9 7 9 1 11 2
10 10 0 9 15 13 13 1 9 9 2
15 11 11 13 16 3 16 9 9 13 2 10 9 13 9 2
5 13 10 0 9 2
1 11
7 2 9 2 9 2 9 2
7 2 9 2 9 2 9 2
30 3 2 1 9 13 1 1 13 2 10 13 9 9 12 9 13 0 9 2 1 11 2 9 9 12 2 9 13 9 9
19 11 2 1 9 12 1 11 12 9 1 11 11 2 15 13 10 9 9 2
19 15 9 13 9 9 9 7 11 4 13 14 13 15 13 1 9 9 9 2
17 4 15 6 13 10 9 13 0 7 13 10 9 1 11 16 0 2
1 9
23 11 11 11 11 11 11 9 9 9 2 2 12 2 12 9 2 2 12 2 12 9 2 8
5 0 1 10 9 2
8 13 15 7 15 9 13 3 2
10 13 4 10 9 9 7 9 1 11 2
10 10 0 9 15 13 13 1 9 9 2
15 11 11 13 16 3 16 9 9 13 2 10 9 13 9 2
5 13 10 0 9 2
1 11
7 2 9 2 9 2 9 2
7 2 9 2 9 2 9 2
12 15 13 1 11 1 11 11 2 3 13 15 9
16 11 2 4 15 6 13 1 11 10 9 1 10 9 1 9 2
16 15 9 4 13 15 9 1 9 9 9 3 1 9 9 9 2
1 9
23 11 11 11 11 11 11 9 9 9 2 2 12 2 12 9 2 2 12 2 12 9 2 8
30 3 2 1 9 13 1 1 13 2 10 13 9 9 12 9 13 9 9 2 1 11 2 9 9 12 2 9 13 9 9
19 11 2 1 9 12 1 11 12 9 1 11 11 2 15 13 10 9 9 2
19 15 9 13 9 9 9 7 11 4 13 14 13 15 13 1 9 9 9 2
17 4 15 6 13 10 9 13 0 7 13 10 9 1 11 16 0 2
1 9
23 11 11 11 11 11 11 9 9 9 2 2 12 2 12 9 2 2 12 2 12 9 2 8
5 0 1 10 9 2
8 13 15 7 15 9 13 3 2
10 13 4 10 9 9 7 9 1 11 2
10 10 0 9 15 13 13 1 9 9 2
15 11 11 13 16 3 16 9 9 13 2 10 9 13 9 2
5 13 10 0 9 2
1 11
7 2 9 2 9 2 9 2
7 2 9 2 9 2 9 2
15 6 13 13 11 14 9 1 9 1 11 11 9 0 12 2
4 13 13 9 2
9 6 13 10 9 1 10 13 9 2
11 16 15 13 10 9 7 9 2 6 13 2
24 15 4 14 13 10 9 14 13 15 13 2 15 4 13 15 10 9 7 15 4 13 1 15 2
8 3 13 15 9 1 11 11 2
9 4 10 9 1 11 13 15 9 2
3 6 11 2
9 3 4 15 13 14 13 11 13 2
6 3 13 11 14 9 2
9 4 15 3 13 1 10 0 9 2
6 2 11 2 11 11 2
11 6 15 4 13 0 3 12 9 10 9 2
7 15 13 15 4 13 0 2
17 15 4 14 13 15 1 10 9 1 9 7 4 3 13 1 15 2
30 15 4 3 4 13 15 0 9 2 10 9 13 15 14 13 3 0 1 0 9 3 15 4 13 15 9 1 10 9 2
25 11 3 13 15 15 13 10 9 1 9 1 15 9 7 15 13 15 13 0 14 13 3 0 3 2
4 0 1 15 2
17 11 2 11 7 15 4 13 14 13 3 10 10 11 9 9 9 2
16 16 10 9 13 2 15 4 13 10 0 9 1 11 13 9 2
8 6 9 2 15 13 9 3 2
7 15 13 3 3 3 3 2
2 11 2
10 15 4 14 13 16 15 9 13 11 2
5 4 15 13 15 2
13 11 11 9 9 9 2 12 9 2 12 9 2 12
1 2
31 10 9 7 10 9 13 1 15 1 10 11 11 13 0 7 13 3 1 10 9 1 10 9 7 9 1 15 15 4 13 2
13 16 15 4 13 10 9 1 9 6 13 10 9 2
1 2
17 11 2 11 7 15 4 13 14 13 3 10 10 11 9 9 9 2
16 16 10 9 13 2 15 4 13 10 0 9 1 11 13 9 2
17 6 2 15 3 13 14 13 1 11 16 15 13 3 1 10 9 2
12 7 15 13 15 13 1 10 9 1 11 3 2
25 4 15 10 13 3 7 13 10 9 9 1 11 16 15 4 3 7 4 15 3 13 11 11 15 2
18 15 0 9 13 11 11 2 11 11 2 9 2 2 2 7 11 11 2
6 4 14 13 1 15 2
20 15 4 3 13 14 13 1 15 15 4 13 14 13 9 9 7 9 9 9 2
10 10 9 1 10 9 2 3 10 9 2
21 3 2 15 4 13 3 0 16 15 9 14 13 16 0 1 10 9 4 13 0 2
9 11 2 9 13 0 1 12 9 2
16 10 9 9 1 11 4 13 7 9 2 12 7 9 2 12 2
8 15 4 14 13 1 1 11 2
27 15 13 7 13 15 2 13 15 1 15 9 2 7 15 4 13 3 7 13 10 9 1 15 9 1 11 2
11 3 15 4 13 15 1 11 1 15 9 2
19 1 10 9 2 11 7 11 4 13 9 16 15 15 4 13 1 11 11 2
2 11 2
15 1 15 9 10 0 9 3 2 13 6 13 10 13 9 2
26 10 9 4 4 13 1 10 9 10 13 1 10 9 2 9 15 13 1 11 11 3 10 0 9 3 2
21 15 3 13 2 0 1 9 2 13 1 15 9 2 13 15 13 9 1 10 9 2
12 15 13 15 16 15 4 13 15 1 15 9 2
28 3 2 16 15 13 1 15 2 15 4 13 15 9 2 9 1 11 11 1 11 11 1 11 14 13 15 0 2
15 2 15 9 9 13 15 13 1 1 10 9 1 11 2 2
8 9 1 10 15 9 1 15 2
24 11 11 11 11 7 11 11 12 11 11 11 2 11 11 12 9 2 12 9 2 12 9 2 8
1 5
28 10 9 4 13 9 10 13 0 2 0 7 2 7 9 9 9 1 10 0 9 1 10 13 9 2 8 2 2
17 10 9 2 9 7 9 1 9 7 9 1 0 9 4 3 13 2
17 16 15 13 14 10 13 9 2 6 13 10 9 7 13 10 9 2
11 2 8 8 8 8 8 8 8 8 9 2
9 2 8 8 8 8 8 8 9 2
18 2 8 8 8 8 8 8 8 8 9 2 8 8 8 8 8 8 9
15 10 0 9 1 10 9 1 9 16 13 9 1 10 9 2
17 11 11 13 10 9 1 9 9 1 11 0 9 1 10 11 11 2
14 15 13 3 16 9 3 13 3 12 9 1 15 9 2
18 15 13 1 11 3 7 13 16 10 9 3 13 0 9 1 15 9 2
15 11 11 13 12 1 10 9 7 13 2 2 15 13 0 2
19 4 15 13 10 0 9 3 15 13 9 3 14 13 10 9 1 9 2 2
10 2 9 9 2 2 13 10 0 9 2
30 11 7 11 2 9 1 11 11 11 2 13 10 1 15 9 1 10 9 14 13 10 11 7 11 9 3 1 11 11 2
29 15 3 13 12 0 9 2 15 4 13 1 10 2 0 1 9 2 9 1 10 9 1 9 12 1 9 9 12 2
10 15 4 4 13 10 13 9 1 15 2
10 15 4 13 15 1 15 1 15 9 2
7 3 15 4 13 13 3 2
5 15 4 13 0 2
12 15 4 13 1 15 9 1 12 7 12 9 2
8 15 3 4 14 13 14 13 2
15 15 13 15 13 10 9 13 1 1 15 7 10 0 9 2
6 15 4 13 10 9 2
15 13 14 13 15 3 1 10 9 2 7 15 13 14 0 2
10 15 13 10 9 1 15 9 2 9 2
5 8 1 12 12 9
2 0 2
2 6 2
25 15 4 14 13 0 1 10 9 9 2 15 13 3 15 13 0 2 4 13 1 12 1 9 6 2
11 15 4 13 0 16 15 13 10 10 9 2
16 3 15 4 13 1 15 2 15 13 1 10 9 7 10 9 2
2 9 2
11 11 11 13 10 9 1 11 2 7 11 2
2 11 11
3 10 11 9
15 15 3 13 15 14 13 10 11 2 9 9 2 1 15 2
13 10 9 13 0 7 2 1 10 9 2 3 0 2
13 15 0 9 13 1 9 1 11 11 1 11 11 2
18 1 10 2 15 13 9 1 12 9 3 1 11 14 13 10 11 9 2
24 15 13 15 4 13 14 13 15 15 9 13 0 2 3 15 4 13 10 9 1 10 9 3 2
9 3 13 10 0 12 3 13 9 2
9 8 2 11 11 2 9 2 11 11
9 8 2 11 11 2 9 2 11 11
5 8 2 0 11 9
14 8 2 11 11 2 9 2 10 11 11 1 3 11 11
7 8 2 11 11 2 9 9
16 8 2 11 11 11 2 0 11 2 11 11 1 11 2 11 2
12 8 2 11 11 2 11 2 11 11 2 11 2
7 8 2 0 11 11 11 11
8 8 2 11 11 2 9 2 11
7 8 2 11 11 11 11 11
24 16 15 4 14 13 10 9 2 15 4 13 15 0 14 13 3 3 3 10 1 10 0 9 2
24 16 15 13 10 9 15 4 13 15 13 1 9 1 10 9 9 2 6 13 15 13 1 8 2
12 9 13 10 0 9 3 7 3 2 3 11 2
11 15 13 9 1 0 9 13 2 3 3 2
23 10 9 4 13 3 0 14 13 2 16 13 9 1 10 1 15 9 4 13 10 10 9 2
7 13 15 10 1 15 9 2
2 11 2
2 13 2
1 11
2 11 2
10 12 9 1 11 11 11 4 13 0 2
11 15 4 13 15 1 10 9 1 12 9 2
3 0 9 2
1 11
2 11 2
13 11 13 10 0 9 2 9 9 9 10 9 2 2
12 15 1 12 1 10 9 7 9 9 1 12 2
12 15 4 13 1 11 11 11 2 11 11 2 2
1 11
2 11 2
15 4 15 13 3 11 9 3 12 1 12 9 1 15 9 2
8 15 4 13 3 0 1 15 2
14 15 4 13 14 13 9 1 3 12 14 13 10 9 2
15 15 4 13 16 15 4 14 13 1 3 0 1 15 9 2
14 9 1 15 9 3 2 7 9 16 13 0 1 15 2
2 11 11
1 3
3 11 13 2
6 15 4 13 10 9 2
2 11 2
5 11 13 1 15 2
6 15 1 12 15 9 2
1 11
6 6 13 1 2 8 2
7 3 1 11 2 11 12 2
2 11 2
3 10 9 2
18 15 4 13 10 0 9 1 9 2 9 9 2 1 11 2 11 12 2
6 4 15 13 1 10 9
1 11
6 6 13 1 2 8 2
16 15 4 3 13 3 1 11 3 15 4 13 15 1 10 9 2
2 6 2
2 11 2
17 4 15 13 1 11 1 10 9 7 15 4 13 15 1 10 9 2
1 11
6 6 13 1 2 8 2
2 11 2
17 3 1 10 0 9 9 9 1 11 2 11 12 1 12 9 11 2
1 11
2 11 2
7 11 12 2 12 15 13 2
8 15 4 13 10 0 9 9 2
6 3 4 15 13 15 2
1 11
6 6 13 1 2 8 2
2 11 2
10 15 13 3 0 1 12 1 11 12 2
17 3 1 10 0 9 9 9 1 11 2 11 12 1 12 9 11 2
1 11
2 11 2
11 11 2 11 12 2 12 4 13 1 15 2
11 15 4 13 0 14 13 15 9 2 8 2
16 15 4 13 10 9 15 13 1 9 1 15 9 14 13 15 2
1 11
6 6 13 1 2 8 2
2 11 2
13 0 14 13 1 15 7 15 13 0 15 13 0 2
6 3 13 11 1 12 2
14 15 4 13 1 9 7 13 14 0 14 13 15 9 2
21 15 13 0 14 13 0 1 15 1 15 9 9 9 7 9 9 1 1 9 9 2
6 3 4 10 9 13 2
33 15 4 13 1 10 9 1 9 9 7 13 0 14 13 16 11 2 11 2 11 7 11 4 13 14 13 10 9 14 13 1 15 2
6 13 1 10 9 9 2
17 16 15 13 9 0 9 2 15 4 13 15 1 15 9 2 8 2
10 15 13 3 0 16 15 15 4 13 2
26 15 4 14 13 1 10 9 3 7 4 13 0 14 13 1 10 9 1 15 1 10 9 13 15 9 2
39 15 13 10 3 0 9 2 16 9 2 1 2 10 2 9 9 9 2 0 2 12 5 12 2 7 9 1 9 2 13 10 0 9 9 1 11 7 11 2
27 11 13 9 7 9 9 9 9 2 9 9 2 7 2 9 2 9 14 13 9 9 9 1 0 9 9 2
34 1 12 9 14 0 2 9 9 2 15 13 0 1 10 9 2 8 2 15 13 11 3 14 13 5 12 7 15 13 1 5 12 2 2
5 13 10 0 9 2
1 11
2 11 2
8 15 4 13 0 1 10 9 2
12 15 1 11 2 11 12 2 1 12 7 12 2
12 6 2 13 15 13 10 9 4 13 1 15 2
9 15 4 13 0 14 13 15 3 2
1 11
18 9 1 10 9 2 4 15 13 10 9 14 13 10 9 1 10 9 2
4 6 13 1 8
2 8 8
3 12 12 9
5 15 4 15 13 2
5 8 1 12 12 9
11 3 11 7 11 13 10 12 12 9 9 2
24 16 0 2 15 13 10 0 9 14 13 10 9 4 13 14 13 10 9 1 10 0 9 9 2
22 15 4 3 13 1 10 9 9 7 4 13 1 10 3 0 9 9 9 1 10 9 2
16 15 4 3 13 10 12 9 13 1 9 9 1 10 9 9 2
16 10 9 1 10 9 13 10 0 7 0 9 1 10 0 9 2
7 10 12 12 13 0 9 2
12 13 15 13 16 15 13 15 13 0 7 0 2
23 15 3 2 13 0 1 9 16 10 11 7 11 9 13 3 0 7 10 0 9 1 15 2
1 9
1 11
2 11 2
10 10 0 9 13 10 9 2 11 9 2
20 15 4 13 14 13 1 3 0 9 15 3 13 0 2 15 3 3 13 15 2
30 15 4 13 10 9 1 11 10 4 13 10 9 1 0 11 9 13 10 9 2 13 15 1 10 9 2 16 15 13 2
11 15 4 13 10 9 1 10 9 1 15 2
13 15 4 14 13 1 11 14 9 1 10 11 9 2
9 15 13 15 4 13 15 0 9 2
16 6 13 15 13 2 15 13 0 14 13 13 1 11 7 15 2
2 9 2
1 11
2 11 2
10 13 15 13 16 15 13 14 13 9 2
12 15 13 0 16 15 13 0 14 13 9 9 2
2 9 2
2 11 11
2 11 11
3 12 12 9
2 11 2
27 13 1 15 9 4 10 13 9 1 10 2 2 8 2 9 7 2 8 2 9 12 1 10 9 9 9 2
47 15 4 4 13 1 10 9 13 12 2 7 13 11 14 13 9 1 15 2 8 2 13 9 13 1 11 1 11 12 2 12 2 7 2 8 2 9 9 13 1 11 1 11 9 2 12 2
7 15 13 3 1 15 9 2
2 3 2
3 11 11 11
9 15 4 14 13 9 1 10 9 2
2 11 11
3 8 8 8
3 12 12 9
4 0 9 11 2
30 15 13 14 13 1 1 15 13 10 9 7 9 1 9 9 1 10 13 9 9 10 15 13 11 4 13 1 15 3 2
15 8 2 11 11 2 9 1 11 11 11 2 12 1 0 2
14 8 2 9 2 9 1 11 11 11 2 12 1 0 2
3 6 13 2
2 9 2
1 11
28 2 9 1 13 9 2 10 13 9 0 1 2 11 2 1 10 9 9 4 4 13 1 10 9 9 16 13 2
19 13 9 5 2 0 9 1 9 9 1 13 9 2 2 9 2 12 2 2
2 11 11
56 2 0 9 2 1 10 9 9 2 2 11 2 4 13 2 10 9 1 2 2 10 9 0 1 2 9 2 12 2 2 2 10 13 4 13 0 1 10 9 9 1 10 2 9 9 2 3 4 15 13 1 10 9 2 2 2
2 11 11
2 11 11
3 12 12 9
28 2 9 1 13 9 2 10 13 9 0 1 2 11 2 1 10 9 9 4 4 13 1 10 9 9 16 13 2
19 13 9 5 2 0 9 1 9 9 5 13 9 2 2 9 2 12 2 2
2 11 11
17 10 9 2 8 2 1 11 13 9 1 10 0 7 11 0 9 2
38 1 10 9 1 10 3 3 0 9 2 10 11 7 11 9 9 13 14 13 1 9 16 10 13 10 2 9 2 1 9 9 1 10 9 7 9 9 2
8 15 13 3 16 13 1 15 2
2 9 2
1 11
6 9 9 1 15 9 2
18 15 4 14 13 10 9 14 13 1 15 1 10 9 14 13 15 9 2
8 13 15 13 15 9 1 11 2
2 13 0
2 11 11
2 8 8
3 12 12 9
2 11 2
12 15 13 14 13 10 9 9 1 10 9 9 2
31 10 9 13 3 1 10 9 9 9 2 10 3 1 2 2 12 9 9 1 10 9 1 10 9 2 2 4 13 1 13 2
13 1 11 11 11 2 11 2 12 11 12 9 2 9
91 10 9 9 1 11 11 11 7 11 11 2 2 11 2 2 1 9 1 11 11 7 11 11 1 10 7 2 8 2 1 10 9 1 10 9 13 10 9 14 13 1 11 2 9 4 13 10 9 9 9 7 4 13 10 0 9 9 2 7 2 8 2 1 10 9 1 10 9 13 10 9 14 13 1 11 2 9 4 13 10 9 9 9 7 4 13 10 0 9 9 2
16 10 9 9 9 4 13 10 9 13 1 10 9 1 10 9 2
49 10 0 9 9 4 13 10 9 9 9 2 13 1 10 0 11 11 11 2 11 2 9 9 16 13 1 11 1 9 9 1 10 9 1 10 9 2 13 1 10 9 13 1 10 9 1 10 9 2
23 10 9 1 10 9 4 13 1 10 9 2 8 2 13 3 1 10 9 9 1 10 9 2
20 10 9 9 4 13 10 9 2 8 2 13 3 1 10 9 9 1 10 9 2
24 10 9 4 13 1 9 2 10 2 0 9 2 2 1 11 9 2 10 2 9 9 2 2 2
15 10 9 1 9 1 10 10 9 4 13 4 13 11 9 2
12 6 13 15 13 15 9 16 15 13 10 9 2
1 9
1 11
20 15 13 14 13 10 9 13 1 10 13 15 4 14 13 9 9 9 1 11 2
14 4 15 13 1 15 15 13 14 13 15 1 1 9 2
2 9 2
1 11
16 15 9 3 13 7 13 15 9 14 9 4 13 1 12 9 2
5 11 2 11 9 2
34 15 4 13 3 1 9 1 10 9 2 7 10 9 4 13 12 9 7 3 15 4 13 15 1 12 0 9 16 15 13 15 1 9 2
13 15 4 13 15 4 3 13 1 10 9 12 9 2
1 11
9 9 9 1 9 9 2 16 13 2
9 15 13 10 9 1 9 0 9 2
19 15 9 4 13 9 1 11 11 2 3 15 4 4 13 10 9 1 11 2
27 15 4 13 14 13 1 9 3 2 7 15 4 13 10 9 9 1 11 11 10 15 4 14 4 13 3 2
7 15 4 13 9 9 3 2
1 11
15 15 13 15 4 14 13 15 9 16 13 1 10 9 11 2
18 15 13 16 13 11 1 10 0 11 11 9 1 10 11 1 11 11 2
15 15 13 10 9 1 9 2 7 15 4 3 13 1 15 2
4 5 9 9 5
13 10 9 1 10 9 4 13 0 7 2 7 0 2
16 10 9 4 13 14 4 13 1 3 10 9 7 9 13 3 2
45 16 15 13 14 10 13 9 7 10 13 9 1 10 13 9 2 15 4 3 13 16 10 9 2 9 7 9 1 10 9 7 15 9 2 16 10 2 7 10 9 13 3 4 13 2
25 16 15 4 13 10 9 1 9 2 6 3 13 10 9 1 9 9 7 13 10 9 1 15 9 2
2 13 15
2 11 11
3 12 12 9
9 15 13 10 9 1 9 0 9 2
19 15 9 4 13 9 1 11 11 2 3 15 4 4 13 10 9 1 11 2
27 15 4 13 14 13 1 9 3 2 7 15 4 13 10 9 9 1 11 11 10 15 4 14 4 13 3 2
7 15 4 13 9 9 3 2
1 11
13 15 4 14 13 14 13 0 16 15 13 15 9 2
6 13 15 0 1 15 2
4 8 8 8 8
3 12 12 9
8 11 11 4 4 13 10 9 2
9 10 9 2 11 2 11 9 2 12
4 10 9 2 12
4 10 9 2 12
9 10 9 2 12 9 5 12 9 11
5 10 9 2 11 9
10 10 9 2 9 12 7 9 12 9 9
17 16 15 13 10 9 7 9 2 6 13 0 14 13 15 1 12 2
3 13 15 2
2 11 11
20 6 2 7 10 9 15 13 15 9 9 2 10 9 10 13 9 1 10 9 2
6 0 9 9 1 9 2
9 15 13 15 9 14 9 13 3 2
16 13 15 0 1 10 9 15 4 13 13 3 2 0 2 2 2
1 11
2 11 11
3 12 12 9
2 11 11
3 12 12 9
9 15 13 10 9 1 9 0 9 2
19 15 9 4 13 9 1 11 11 2 3 15 4 4 13 10 9 1 11 2
27 15 4 13 14 13 1 9 3 2 7 15 4 13 10 9 9 1 11 11 10 15 4 14 4 13 3 2
7 15 4 13 9 9 3 2
1 11
30 1 0 7 0 2 10 10 9 1 10 9 2 9 2 7 2 9 2 13 15 2 16 11 13 10 0 9 1 9 2
1 11
16 3 2 13 9 12 5 12 2 9 9 5 9 1 15 9 2
1 11
4 8 8 8 8
3 12 12 9
22 15 13 10 9 1 9 7 15 13 15 13 13 9 13 10 1 10 9 1 0 9 2
13 6 13 16 10 9 13 0 1 9 1 15 9 2
11 10 9 10 15 13 9 1 13 1 0 2
2 9 2
2 11 2
15 15 13 10 9 16 16 15 4 13 1 12 0 9 9 2
14 6 13 10 0 9 1 13 1 10 9 15 13 3 2
16 6 13 10 13 9 9 1 11 7 13 10 9 1 9 9 2
32 15 13 0 16 10 1 10 9 1 10 13 9 13 0 2 13 9 2 16 10 9 4 4 13 3 1 11 11 7 11 11 2
2 9 2
2 11 2
7 3 13 10 9 13 9 2
2 11 2
8 15 3 13 15 14 13 3 2
4 3 15 13 2
14 3 13 4 10 9 9 9 2 3 12 0 9 2 2
2 2 9
2 2 9
4 8 8 8 8
3 12 12 9
8 11 11 4 4 13 10 9 2
9 10 9 2 11 2 11 9 2 12
4 10 9 2 12
4 10 9 2 12
9 10 9 2 12 9 5 12 9 11
5 10 9 2 11 9
10 10 9 2 9 12 7 9 12 9 9
17 16 15 13 10 9 7 9 2 6 13 0 14 13 15 1 12 2
3 13 15 2
3 11 11 12
2 11 11
3 12 12 9
3 0 9 2
17 15 4 13 10 13 9 9 9 9 2 13 9 1 15 0 9 2
8 15 13 3 16 13 15 3 2
2 9 2
1 11
10 11 11 13 10 11 9 15 13 11 2
2 8 8
3 12 12 9
12 15 4 14 13 10 0 9 13 3 1 11 2
9 13 10 1 15 0 1 10 9 2
26 15 4 13 10 9 1 10 11 2 11 11 0 7 0 9 7 15 4 14 13 14 13 10 9 9 2
32 15 9 9 2 11 11 2 7 9 2 11 11 2 13 14 13 10 9 9 14 13 9 9 1 10 9 14 13 10 11 9 2
24 15 3 13 16 9 1 11 2 11 11 2 11 11 4 13 10 9 9 1 11 1 10 9 2
17 15 13 14 1 10 9 9 2 3 6 13 11 11 1 15 9 2
1 11
3 6 11 2
14 15 13 15 0 9 7 13 0 14 13 1 15 9 2
10 15 13 16 16 15 9 4 13 3 2
6 15 13 3 0 9 2
26 16 15 13 15 9 7 9 14 9 13 7 3 13 15 13 2 15 13 10 3 0 9 1 15 9 2
26 7 15 4 13 3 0 14 13 0 0 9 7 14 4 13 10 9 14 4 4 13 1 0 0 9 2
11 13 16 16 11 4 13 3 3 1 11 2
7 15 4 13 10 0 9 2
17 15 13 3 0 14 13 16 15 4 13 15 9 13 1 10 9 2
31 16 15 4 13 1 10 9 3 0 9 13 3 0 2 15 13 0 16 10 0 9 14 13 10 3 0 0 9 15 4 2
26 1 1 15 9 2 1 10 0 12 9 15 0 9 11 4 13 1 10 0 9 1 11 11 2 11 2
16 15 13 16 15 4 3 13 1 10 9 1 9 1 11 11 2
21 15 13 3 1 15 9 7 3 16 13 4 4 13 1 11 11 1 11 2 11 2
10 10 0 11 9 15 0 9 4 13 2
12 15 4 13 1 15 9 11 7 15 9 11 2
14 15 13 10 12 9 2 12 9 2 12 9 0 9 2
23 3 15 3 13 12 9 7 12 9 13 1 3 12 9 5 12 9 3 1 10 0 9 2
8 15 13 10 0 9 1 9 2
6 15 4 13 3 3 2
17 15 4 13 3 16 13 11 2 11 2 11 3 15 13 1 11 2
21 15 4 13 0 14 13 9 1 15 7 15 9 4 15 3 13 9 14 13 11 2
8 15 13 15 13 10 0 9 2
15 13 15 1 15 0 9 16 11 11 14 13 1 15 9 2
16 3 2 1 1 11 11 14 9 15 4 14 13 0 14 13 2
4 13 15 3 2
5 11 11 11 0 9
2 6 2
14 3 14 13 15 13 16 15 13 16 12 9 4 13 2
10 15 13 14 13 1 11 11 16 13 2
2 9 2
1 11
3 0 11 2
19 16 15 13 2 15 0 9 13 1 11 2 11 12 1 12 5 12 9 2
43 1 10 0 9 7 3 2 15 4 4 13 3 10 9 9 10 15 13 13 10 9 2 7 15 4 13 14 13 1 3 0 1 15 16 0 1 10 9 14 13 1 15 2
37 3 2 11 11 4 13 14 13 1 15 1 11 14 13 1 10 9 15 4 13 7 3 14 13 15 10 9 1 10 1 10 9 16 15 13 15 2
44 15 13 12 0 9 1 10 9 2 10 15 13 13 1 12 9 2 3 2 10 9 1 10 9 3 1 12 5 12 9 2 7 3 10 9 1 9 11 1 12 5 12 9 2
5 3 13 10 9 2
15 4 15 6 13 15 13 10 1 15 4 13 0 1 15 2
9 5 11 2 11 12 12 5 12 9
9 5 11 2 11 12 12 5 12 9
9 5 11 2 11 12 12 5 12 9
3 0 9 2
2 11 11
5 0 9 2 11 2
23 11 11 4 13 14 13 10 11 11 9 2 2 10 0 8 0 9 13 1 10 9 2 2
16 11 13 14 13 3 7 13 15 16 15 15 13 15 4 13 2
12 6 13 15 13 3 15 4 13 14 13 15 2
4 9 2 11 2
1 11
22 3 13 10 9 1 10 0 0 9 1 10 9 2 15 4 13 1 1 10 9 9 2
18 10 11 9 13 10 0 7 10 9 13 10 10 1 12 7 3 0 2
1 8
5 2 8 8 9 2
4 2 8 8 9
26 3 2 11 11 4 13 1 11 11 2 11 13 1 10 9 2 3 15 13 10 9 2 1 11 12 2
2 11 11
3 1 2 5
3 11 12 9
32 3 11 11 7 11 11 13 15 10 9 1 10 9 10 15 4 13 1 11 12 1 12 9 14 4 13 1 10 11 11 11 2
12 15 13 16 15 4 13 0 14 13 10 9 2
22 1 10 9 1 11 11 7 9 15 4 13 0 9 1 9 1 11 1 10 0 9 2
20 3 15 13 9 14 13 10 0 9 7 13 3 0 9 1 15 0 9 9 2
29 10 11 11 11 11 4 13 1 1 9 9 2 9 2 7 13 9 0 16 13 0 9 9 16 13 9 1 11 2
13 15 4 13 10 9 14 13 1 15 1 10 9 2
2 11 11
4 11 11 11 12
1 2
26 15 13 0 1 11 11 2 7 15 4 13 1 10 3 0 9 2 3 4 3 13 0 14 13 8 2
17 15 13 10 2 9 9 9 2 1 10 11 11 11 1 11 11 2
28 1 9 9 2 6 13 16 15 13 10 9 7 13 15 13 16 15 13 10 9 9 10 15 13 15 14 13 2
3 13 15 2
8 11 11 0 9 1 11 11 12
1 5
15 9 2 10 9 1 10 9 13 0 7 4 13 3 0 2
19 16 15 13 14 10 13 9 2 15 4 14 13 2 13 7 13 10 9 2
71 16 10 9 7 10 9 4 13 14 13 0 1 10 9 7 0 9 10 4 13 10 9 9 1 10 15 4 13 7 13 2 15 13 10 9 1 10 9 14 13 16 15 13 9 0 7 10 9 4 13 1 11 11 7 10 1 15 9 1 10 9 7 9 13 1 10 9 1 15 9 2
1 5
12 11 11 4 13 10 13 9 9 1 11 11 2
4 6 11 11 2
28 15 13 9 13 1 15 9 2 7 11 11 13 15 14 13 15 13 16 10 9 4 14 13 1 15 2 3 2
2 0 2
1 11
19 13 15 13 16 15 13 10 9 1 10 11 2 11 11 9 1 10 9 2
18 15 4 13 11 9 1 9 7 13 11 7 11 1 9 2 5 12 2
13 15 4 14 13 16 15 9 4 13 15 7 14 2
11 4 15 13 15 10 9 9 15 4 13 2
10 6 13 11 9 12 1 10 9 9 2
7 11 4 14 13 10 9 2
2 9 2
1 11
2 11 2
5 5 12 1 9 2
13 11 11 11 2 11 9 9 12 11 11 2 11 12
8 3 15 13 14 10 0 9 2
19 13 12 9 2 11 12 12 2 12 9 2 12 5 12 2 12 11 9 2
23 9 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 9 2 12 9 9 2
18 6 2 15 4 13 1 1 12 0 9 1 11 11 14 13 10 9 2
6 13 15 13 14 13 2
11 15 13 10 9 9 4 13 0 3 3 2
6 3 2 11 13 15 2
7 15 13 5 12 7 9 2
17 15 13 3 0 7 13 9 2 9 7 9 1 10 9 1 9 2
3 3 0 2
12 15 13 14 13 1 0 9 3 1 11 14 2
18 11 13 2 15 4 13 14 13 0 1 15 14 13 15 0 11 9 2
17 15 13 6 2 13 10 9 3 16 15 4 13 0 1 15 9 2
9 15 3 13 14 13 9 16 13 2
17 15 4 13 9 9 7 13 14 13 11 11 9 1 11 1 9 2
15 12 9 13 1 0 2 10 9 4 14 13 1 15 9 2
9 11 9 13 3 1 1 5 12 2
4 6 2 6 2
13 13 14 13 1 5 12 7 3 15 4 13 0 2
19 15 13 1 11 7 15 13 15 13 10 9 1 9 13 1 11 14 9 2
14 15 13 14 13 10 9 7 13 13 9 1 10 9 2
12 15 4 13 14 13 10 9 7 9 3 3 2
11 15 4 13 3 3 7 13 10 9 13 2
8 11 13 15 4 13 15 3 2
14 15 3 3 13 10 9 16 15 4 13 1 1 15 2
6 3 13 2 3 13 2
5 3 13 10 9 2
6 15 4 13 1 12 2
18 13 0 14 13 15 9 3 1 10 9 9 7 13 1 10 0 9 2
9 15 13 3 0 13 3 0 9 2
20 15 13 14 13 3 7 13 1 10 9 1 10 9 7 13 1 10 9 9 2
25 15 13 10 9 1 9 1 15 9 10 9 3 7 10 9 10 13 14 13 16 15 13 9 9 2
3 3 0 2
19 15 9 4 13 0 9 7 4 13 15 15 4 13 1 10 12 9 9 2
18 15 3 13 10 9 1 9 7 15 13 14 1 0 3 0 15 13 2
12 15 4 13 14 13 10 9 2 9 9 9 2
14 15 13 15 3 13 14 13 0 14 13 9 9 9 2
7 15 4 13 12 1 12 2
7 15 13 3 0 1 15 2
9 11 13 11 4 13 1 3 3 2
7 15 4 8 13 15 3 2
11 15 13 0 15 4 13 14 13 1 15 2
2 8 2
10 1 10 9 2 13 0 7 13 0 2
25 15 4 4 13 1 9 2 3 3 16 15 13 15 9 0 7 15 9 0 2 15 4 13 0 2
13 6 2 13 9 1 15 12 13 0 9 1 15 2
10 6 2 11 11 13 10 0 9 3 2
4 13 1 11 2
12 15 13 10 3 0 9 3 1 12 2 12 2
9 15 4 13 12 9 1 10 9 2
17 15 13 8 3 1 10 0 7 15 4 13 15 3 15 13 3 2
8 15 3 13 15 9 1 9 2
9 15 9 13 3 0 14 13 1 2
10 1 10 13 11 9 15 13 12 9 2
5 13 15 9 0 2
2 6 2
1 9
1 11
34 11 11 11 2 11 12 11 11 11 11 12 2 9 9 11 2 11 12 9 12 12 12 12 2 12 2 9 12 12 12 9 12 12 12
4 15 4 13 2
9 15 13 15 13 10 3 0 9 2
6 4 13 0 13 9 2
7 15 13 12 9 1 15 2
22 8 2 15 13 10 9 1 10 12 9 7 15 4 13 14 13 15 1 1 15 9 2
5 15 4 15 13 2
24 16 15 13 0 2 3 4 15 13 15 9 14 13 1 1 10 9 7 10 9 4 15 13 2
13 8 2 15 4 13 0 14 13 1 10 11 9 2
10 3 0 1 9 14 9 4 15 13 2
15 0 9 2 13 15 10 12 9 2 15 13 0 16 13 2
16 15 13 15 3 13 9 2 3 3 12 9 2 1 10 11 2
5 15 4 14 13 2
24 15 4 13 16 0 1 10 9 10 9 4 14 13 16 15 4 1 11 7 11 1 10 9 2
12 15 13 15 3 13 10 9 7 13 1 11 2
3 6 9 2
14 4 15 6 13 10 11 9 1 11 12 5 11 12 2
14 4 15 13 14 13 10 9 13 1 11 1 10 9 2
8 11 8 13 15 9 10 9 2
17 15 13 16 11 13 15 10 0 13 1 10 9 10 4 14 13 2
1 9
1 11
9 15 4 14 13 3 1 10 9 2
4 6 13 15 12
3 6 11 2
6 15 4 13 15 9 2
12 15 13 15 13 15 9 7 4 14 13 15 2
3 6 11 2
8 15 13 15 1 11 0 9 2
14 15 4 13 3 16 1 10 9 15 3 13 3 3 2
6 15 13 10 9 3 2
5 4 15 13 1 2
2 9 2
2 11 11
3 12 12 9
5 13 1 2 11 11
3 6 11 2
6 15 13 15 9 3 2
11 15 13 9 1 11 2 11 2 7 11 2
2 9 2
5 8 1 12 12 9
4 6 13 1 8
2 9 2
8 9 2 1 2 11 11 11 11
8 11 12 11 12 11 12 11 12
5 8 1 12 12 9
3 6 11 2
21 6 13 15 10 9 7 13 15 10 9 9 1 11 2 11 2 11 7 11 12 2
2 9 2
2 11 11
3 12 12 9
2 11 2
20 4 15 6 13 10 0 9 1 10 9 9 9 2 7 13 1 11 11 2 2
24 1 9 1 10 9 13 9 2 15 13 3 0 1 10 9 9 3 13 9 0 9 1 9 2
26 15 13 16 15 13 9 9 1 10 9 9 3 15 4 14 13 3 16 15 13 10 9 15 3 13 2
7 13 15 13 15 15 13 2
2 9 2
1 11
1 8
3 12 12 9
9 13 6 13 10 0 9 9 9 2
17 15 9 7 0 9 9 4 13 12 9 9 13 9 12 9 9 2
6 11 2 8 8 9 2
4 2 8 8 9
6 15 13 3 1 9 2
6 15 4 13 3 9 2
14 15 13 10 9 9 1 9 2 3 2 16 15 13 2
26 3 2 15 4 13 15 15 4 13 1 1 10 9 2 7 15 4 13 11 13 7 15 4 13 3 2
5 10 4 15 13 2
1 11
11 13 15 1 10 9 14 13 9 9 9 2
10 16 14 2 13 15 9 0 10 4 2
8 15 13 16 11 13 1 11 2
1 11
2 11 11
3 12 12 9
9 16 11 13 0 2 15 13 0 2
1 11
2 6 2
16 15 13 1 11 11 9 13 10 0 9 1 9 13 9 9 2
22 15 0 9 13 16 15 9 13 3 0 7 1 9 1 10 9 1 10 3 13 9 2
15 3 2 15 4 13 10 9 0 9 14 13 11 14 9 2
28 8 2 13 16 9 4 3 4 13 10 13 0 1 9 7 8 2 16 10 13 9 4 13 10 0 9 9 2
10 10 9 4 4 13 1 10 13 9 2
18 15 9 2 3 0 2 13 14 13 10 9 9 1 10 9 1 9 2
17 9 4 13 1 3 7 10 0 9 4 13 3 0 10 13 9 2
18 3 2 15 13 14 13 3 16 15 13 10 9 1 10 9 16 13 2
17 3 2 15 4 4 13 15 1 9 1 15 0 9 1 8 9 2
8 9 1 15 0 9 1 15 2
2 9 2
1 11
2 11 11
3 12 12 9
2 11 2
20 4 15 6 13 10 0 9 1 10 9 9 9 2 7 13 1 11 11 2 2
24 1 9 1 10 9 13 9 2 15 13 3 0 1 10 9 9 3 13 9 0 9 1 9 2
26 15 13 16 15 13 9 9 1 10 9 9 3 15 4 14 13 3 16 15 13 10 9 15 3 13 2
7 13 15 13 15 15 13 2
2 9 2
1 11
1 8
3 12 12 9
9 13 6 13 10 0 9 9 9 2
17 15 9 7 0 9 9 4 13 12 9 9 13 9 12 9 9 2
1 11
5 2 8 8 9 2
4 2 8 8 9
29 15 13 3 0 16 15 14 13 7 13 16 14 13 1 9 15 4 14 13 9 1 15 7 13 15 14 13 15 2
17 15 4 13 15 3 2 13 15 2 7 13 15 16 15 15 13 2
30 7 2 15 13 1 11 10 9 3 15 4 13 10 9 1 15 2 3 16 13 10 9 15 4 14 13 1 13 15 2
14 15 13 3 0 1 15 15 13 2 7 15 13 15 2
9 13 10 13 9 10 0 0 9 2
10 3 7 1 15 4 15 13 15 13 2
2 9 2
1 11
21 16 15 4 13 11 13 2 15 4 3 13 0 14 13 10 9 1 10 9 3 2
8 7 9 7 9 0 13 3 2
11 13 15 13 10 13 0 7 15 4 13 2
1 11
2 11 11
3 12 12 9
6 15 13 3 1 9 2
6 15 4 13 3 9 2
14 15 13 10 9 9 1 9 2 3 2 16 15 13 2
26 3 2 15 4 13 15 15 4 13 1 1 10 9 2 7 15 4 13 11 13 7 15 4 13 3 2
5 10 4 15 13 2
1 11
11 13 15 1 10 9 14 13 9 9 9 2
10 16 14 2 13 15 9 0 10 4 2
8 15 13 16 11 13 1 11 2
1 11
2 11 11
3 12 12 9
9 16 11 13 0 2 15 13 0 2
1 11
2 6 2
16 15 13 1 11 11 9 13 10 0 9 1 9 13 9 9 2
22 15 0 9 13 16 15 9 13 3 0 7 1 9 1 10 9 1 10 3 13 9 2
15 3 2 15 4 13 10 9 0 9 14 13 11 14 9 2
28 8 2 13 16 9 4 3 4 13 10 13 0 1 9 7 8 2 16 10 13 9 4 13 10 0 9 9 2
10 10 9 4 4 13 1 10 13 9 2
18 15 9 2 3 0 2 13 14 13 10 9 9 1 10 9 1 9 2
17 9 4 13 1 3 7 10 0 9 4 13 3 0 10 13 9 2
18 3 2 15 13 14 13 3 16 15 13 10 9 1 10 9 16 13 2
17 3 2 15 4 4 13 15 1 9 1 15 0 9 1 8 9 2
8 9 1 15 0 9 1 15 2
2 9 2
1 11
2 11 11
3 12 12 9
2 11 2
20 4 15 6 13 10 0 9 1 10 9 9 9 2 7 13 1 11 11 2 2
24 1 9 1 10 9 13 9 2 15 13 3 0 1 10 9 9 3 13 9 0 9 1 9 2
26 15 13 16 15 13 9 9 1 10 9 9 3 15 4 14 13 3 16 15 13 10 9 15 3 13 2
7 13 15 13 15 15 13 2
2 9 2
1 11
1 8
3 12 12 9
9 13 6 13 10 0 9 9 9 2
17 15 9 7 0 9 9 4 13 12 9 9 13 9 12 9 9 2
1 11
5 2 8 8 9 2
4 2 8 8 9
7 15 4 13 1 15 3 2
17 3 15 2 11 2 4 13 15 9 9 2 3 13 15 1 11 2
6 15 4 13 3 12 2
15 10 9 2 15 4 13 15 1 15 1 9 1 9 9 2
4 4 15 13 2
1 11
8 15 13 0 14 13 1 15 2
8 15 13 10 0 11 3 3 2
55 15 13 0 2 16 3 15 13 3 15 2 9 2 11 7 11 2 7 11 4 14 3 13 13 9 7 0 9 2 14 16 15 4 13 15 1 15 2 2 2 3 15 13 14 3 10 0 9 1 9 15 4 13 3 2
8 15 13 0 13 10 9 3 2
24 15 13 10 0 9 1 11 13 2 0 11 2 10 13 0 2 0 7 1 9 2 3 0 2
7 15 13 14 1 10 0 2
10 15 13 0 10 10 0 9 11 13 2
29 15 13 15 9 13 3 3 1 9 0 14 2 3 15 13 15 4 13 3 15 4 13 9 0 14 9 2 2 2
16 15 13 11 4 14 13 9 14 13 15 9 16 15 13 0 2
14 15 13 13 1 15 9 2 15 13 0 1 15 9 2
29 3 2 3 2 15 4 13 3 0 9 1 3 3 3 2 16 15 4 14 13 3 15 4 13 14 13 9 9 2
28 15 4 3 13 15 10 12 9 9 3 15 13 15 9 0 9 16 15 4 14 13 12 9 1 10 0 9 2
13 3 15 4 13 14 13 14 13 13 1 10 9 2
19 7 15 9 13 3 0 1 1 15 13 0 9 4 4 13 1 10 9 2
20 15 13 9 4 13 14 13 3 3 3 1 11 7 11 14 13 10 0 9 2
13 15 4 13 14 13 13 14 13 1 15 0 9 2
10 10 0 2 9 9 2 13 3 0 2
14 15 4 13 15 0 9 7 9 2 7 13 3 0 2
26 3 3 16 10 9 1 9 11 13 2 16 15 13 0 14 13 1 15 15 4 14 13 1 15 9 2
11 15 13 10 3 0 9 1 10 1 15 2
10 7 2 15 13 2 15 13 10 9 2
8 15 4 3 13 15 11 9 2
27 15 13 10 9 1 10 9 2 15 9 13 3 1 12 9 2 7 13 10 9 1 10 9 1 12 9 2
7 15 13 0 13 1 15 2
4 13 1 9 2
1 8
3 12 12 9
2 11 2
17 15 4 14 13 2 15 4 15 13 16 2 13 1 10 9 2 2
20 3 2 15 13 15 9 2 7 15 13 10 11 11 9 2 16 15 4 3 13
45 11 7 11 13 10 0 9 1 11 2 15 4 13 16 15 13 12 1 10 0 11 9 15 4 3 13 2 15 3 13 14 13 15 15 2 15 4 14 13 15 13 0 9 2 2
24 9 13 15 13 10 0 9 1 11 2 15 13 0 14 13 15 2 3 3 1 11 7 11 2
11 15 13 15 13 15 0 9 1 15 9 2
28 15 4 13 14 13 10 0 14 13 10 0 9 2 4 14 15 13 0 16 10 9 4 13 1 11 9 2 2
9 3 4 14 11 13 9 15 9 2
18 15 4 15 13 1 15 9 9 1 9 11 2 15 13 3 0 2 2
6 4 15 13 1 11 2
6 13 14 13 1 3 2
3 13 15 2
1 11
1 5
8 2 11 2 11 11 0 9 9
1 5
38 11 12 11 1 10 11 0 9 11 11 2 11 12 11 9 2 12 2 12 2 12 9 2 12 2 12 2 12 9 2 12 2 12 2 12 9 2 8
1 5
7 13 15 9 9 1 2 8
1 5
25 5 5 5 8 5 5 5 8 5 5 5 5 5 5 12 5 5 5 12 9 5 5 5 5 5
4 5 5 5 5
16 6 2 11 11 2 15 4 14 13 10 9 1 1 15 9 2
1 8
2 9 9
24 15 11 11 1 9 9 2 4 13 11 11 2 11 2 11 2 11 1 2 1 2 12 9 9
12 15 4 13 15 9 11 11 1 10 9 3 2
2 9 2
2 8 8
3 12 12 9
17 13 4 10 9 9 1 9 9 1 12 16 9 9 13 1 9 2
2 11 11
2 8 8
3 12 12 9
2 9 2
1 11
6 13 4 10 13 9 2
12 13 15 13 16 10 9 9 13 0 1 15 2
21 16 3 2 15 4 13 15 13 1 11 11 9 2 3 13 15 1 15 1 9 2
9 13 1 15 2 15 13 15 9 2
15 15 13 14 0 15 13 10 9 14 13 9 1 0 9 2
8 6 2 15 4 14 13 15 2
28 13 10 10 11 2 13 9 2 4 3 13 10 9 1 10 0 9 1 10 0 11 9 10 9 1 10 9 2
29 15 9 13 16 15 4 14 13 10 9 0 9 14 3 13 10 9 1 10 9 9 10 13 10 9 1 10 9 2
2 11 11
3 12 12 9
26 16 15 4 13 10 10 9 2 4 15 13 16 15 4 14 13 14 13 1 9 10 0 9 1 11 2
68 1 9 1 11 11 2 2 11 2 2 2 15 13 12 9 9 13 2 11 4 13 15 14 13 10 10 11 9 9 11 13 1 1 13 9 1 10 9 9 9 7 15 13 3 0 14 13 3 2 16 15 4 3 13 1 9 1 13 9 9 1 10 9 1 10 9 9 2
20 11 7 11 11 1 9 4 13 14 13 1 10 11 9 9 1 10 13 9 2
38 1 9 1 11 11 11 11 2 10 9 15 4 13 1 13 3 0 16 15 13 14 13 1 15 0 9 1 9 10 4 13 1 15 1 12 1 9 2
15 11 4 13 1 15 1 11 11 2 10 9 1 15 9 2
2 11 11
3 12 12 9
2 11 2
33 4 15 6 13 15 10 9 16 3 15 13 1 10 9 1 10 9 1 10 13 9 7 13 10 11 9 15 4 13 1 9 1 2
2 9 2
1 11
4 11 11 11 11
3 11 11 11
49 15 13 1 11 11 1 15 9 9 2 7 15 13 16 15 4 14 13 10 9 14 13 9 1 15 0 2 7 3 3 16 15 4 3 13 9 13 1 10 13 9 1 10 9 9 15 13 0 2
4 11 2 11 2
32 10 13 9 9 4 13 1 10 2 0 9 2 2 4 15 6 13 15 13 10 9 15 13 16 15 4 3 13 10 9 9 2
3 13 15 2
1 11
4 6 3 15 2
16 0 15 4 14 13 15 9 1 10 9 14 13 15 3 13 2
26 15 4 3 13 1 9 1 11 7 4 14 13 15 4 13 14 13 1 3 10 0 9 1 15 9 2
24 3 0 9 16 15 13 2 15 13 15 4 3 13 10 0 9 16 15 15 4 13 1 15 2
28 1 1 11 2 9 4 3 13 3 16 15 4 14 13 15 3 3 10 9 2 15 13 12 3 0 9 2 2
31 7 2 15 13 10 0 0 0 9 0 11 7 15 13 4 13 10 0 9 2 15 13 2 14 3 3 0 1 9 8 2
18 1 12 9 15 13 0 2 7 15 3 13 9 10 9 0 14 13 2
25 3 2 15 13 0 15 9 13 15 9 7 11 7 11 13 14 13 15 7 15 13 15 13 3 2
23 3 2 16 15 4 3 13 13 11 2 15 7 11 4 13 15 3 15 13 3 14 13 2
57 15 4 13 16 13 15 1 3 3 12 1 10 11 9 2 15 3 13 14 13 1 3 15 13 14 13 2 3 3 1 3 13 15 1 10 11 2 11 2 11 2 11 11 9 7 10 0 2 9 9 10 13 10 11 9 2 2
9 9 1 11 13 0 7 3 0 2
21 15 13 1 11 7 15 9 0 9 14 13 10 9 2 11 2 7 15 13 0 2
21 3 2 15 4 13 3 1 11 11 1 10 11 11 9 14 13 11 14 9 11 2
8 0 14 13 15 13 3 0 2
6 13 1 15 9 3 2
1 11
3 6 9 2
5 3 4 15 13 2
9 4 14 13 1 15 1 10 9 2
14 10 0 9 13 15 16 15 4 13 1 9 1 11 2
4 13 15 3 2
9 4 15 13 1 15 9 7 3 2
33 1 10 9 2 15 4 13 10 0 9 14 13 10 9 2 7 9 2 2 3 15 13 10 0 9 16 15 14 13 16 15 13 2
43 15 13 16 15 4 13 1 11 3 15 9 13 7 13 10 0 9 9 2 10 4 13 3 10 0 9 2 3 2 2 7 4 13 13 1 11 7 3 1 9 1 11 2
13 15 4 13 15 15 13 13 16 15 3 4 13 2
17 13 15 13 10 0 1 11 7 3 16 15 4 13 1 1 11 2
3 13 9 2
1 11
1 5
4 4 15 13 2
11 13 0 9 7 13 9 9 1 11 11 2
1 8
26 6 11 2 1 2 10 0 2 7 0 2 9 2 9 1 10 11 11 7 1 10 9 10 11 11 2
11 10 9 13 3 0 7 15 13 3 13 2
22 15 4 13 3 13 3 15 13 1 10 1 10 9 10 0 9 15 13 15 1 11 2
31 10 9 9 3 13 14 13 3 0 9 14 13 1 10 9 1 10 3 0 9 2 15 13 15 4 13 15 0 9 2 2
35 15 13 10 0 9 1 11 14 11 9 0 9 3 1 10 9 2 6 2 15 13 14 13 3 1 10 9 2 15 13 15 9 2 2 2
19 3 2 15 13 0 15 4 13 15 3 7 6 15 13 10 3 0 9 2
43 1 10 9 1 15 2 15 4 13 1 0 9 1 10 9 14 13 1 15 9 16 13 11 11 7 13 11 16 3 13 15 2 10 9 3 13 15 0 9 1 9 2 2
26 11 13 15 15 13 15 0 9 1 9 9 7 13 15 16 15 13 14 13 3 10 0 9 15 13 2
34 15 4 13 15 13 3 16 15 13 3 0 10 9 16 15 4 14 13 15 9 0 1 10 9 2 15 13 15 13 10 10 0 9 2
21 3 13 11 3 0 9 14 13 15 7 4 15 3 13 15 4 13 10 0 9 2
7 15 13 10 3 0 9 2
18 13 15 9 4 13 3 7 16 10 9 1 12 13 1 1 10 9 2
11 0 9 1 10 1 10 2 0 2 9 2
1 11
22 2 1 1 10 9 1 9 9 2 15 4 13 14 13 1 15 9 1 10 9 9 2
14 15 4 13 14 13 16 15 4 14 13 3 1 15 2
2 11 11
3 12 12 9
5 3 13 10 9 2
29 15 13 14 13 15 16 15 13 15 9 1 10 9 11 10 0 9 7 15 3 13 15 7 15 13 3 1 12 2
3 0 9 2
20 15 13 1 11 0 9 1 11 14 7 15 4 13 15 13 10 9 1 11 2
8 3 2 9 1 0 9 9 2
7 15 4 13 1 15 3 2
13 3 15 4 13 10 9 1 10 9 15 13 3 2
11 15 13 15 4 4 13 1 15 3 3 2
20 1 10 9 15 4 13 14 13 13 9 1 15 9 14 13 15 14 13 9 2
24 3 2 4 13 1 15 1 0 9 15 13 0 15 4 13 0 14 13 10 9 1 13 9 2
34 13 1 9 3 16 16 15 13 1 13 15 4 14 13 15 13 15 2 7 2 16 15 4 13 2 15 13 10 9 1 10 9 2 2
19 15 4 13 9 1 15 1 10 9 7 3 13 16 9 13 0 1 12 2
10 3 3 1 15 13 3 0 2 15 2
40 13 15 4 13 14 13 16 10 11 11 4 13 3 1 11 11 12 7 4 13 3 1 10 9 1 15 1 10 11 11 2 15 13 3 1 15 7 15 9 2
2 11 11
3 12 12 9
2 6 2
21 15 3 13 1 16 15 13 14 13 10 11 9 14 9 7 13 7 1 10 9 2
16 15 13 10 12 9 9 7 3 16 15 13 15 11 9 13 2
10 15 13 15 13 10 1 15 0 9 2
26 15 4 13 14 13 3 7 13 10 9 10 9 16 15 4 13 1 12 2 15 3 3 13 15 2 2
20 3 13 9 1 12 9 2 6 15 13 0 1 15 13 15 13 3 1 15 2
23 15 13 10 9 16 13 9 14 13 2 10 9 13 16 13 9 14 13 7 14 13 15 2
3 2 11 11
2 11 11
3 12 12 9
17 13 16 10 10 2 9 2 9 13 15 14 13 10 9 1 11 2
1 8
3 12 12 9
19 16 15 13 2 10 13 13 13 9 13 0 9 14 13 1 10 9 9 2
34 11 4 13 9 2 1 9 2 16 13 1 10 9 1 2 9 2 9 7 0 9 1 0 9 1 11 2 1 10 9 1 9 9 2
19 0 9 9 4 13 9 14 13 11 3 3 16 13 3 0 1 9 9 2
8 6 13 16 15 13 14 13 2
5 13 10 0 9 2
18 10 9 4 13 1 10 9 9 7 13 9 10 4 13 0 7 0 2
17 16 15 13 14 10 13 9 2 6 13 10 9 7 13 15 3 2
11 10 0 15 4 13 13 13 10 9 3 2
8 13 15 9 0 15 4 13 2
5 11 11 2 8 2
3 12 12 9
11 3 2 15 13 16 11 13 1 0 9 2
2 9 2
1 11
19 15 13 15 4 13 15 10 9 16 15 13 1 1 9 7 1 10 9 2
21 3 15 13 3 0 14 13 11 11 14 13 1 10 9 9 2 10 9 13 3 2
11 15 4 14 13 16 15 4 13 9 3 2
2 11 2
6 9 1 10 9 9 2
9 4 15 13 10 9 14 13 9 2
9 4 15 13 16 11 4 13 9 2
10 10 1 10 9 3 4 13 14 13 2
2 9 2
1 11
7 13 15 4 13 14 13 2
18 11 11 11 11 9 9 2 12 9 2 12 8 2 8 2 8 2 2
20 11 2 13 10 9 7 13 15 14 13 10 9 1 10 9 2 13 11 11 2
27 11 13 10 9 1 10 9 9 2 16 13 10 9 2 15 7 0 9 1 15 9 4 13 1 10 9 2
15 15 13 12 9 1 10 13 9 7 10 9 1 0 9 2
9 11 13 12 1 15 1 0 9 2
12 15 13 3 1 10 9 9 1 11 11 11 2
19 11 11 11 4 13 1 12 11 11 2 11 2 11 2 9 9 2 12 2
21 15 4 14 13 9 2 9 7 9 1 10 9 2 16 15 13 1 10 9 9 2
13 10 9 4 4 13 2 3 3 16 12 13 0 2
13 13 11 2 15 9 9 7 15 9 1 15 9 2
18 11 11 0 9 11 11 2 12 2 12 12 8 2 8 2 8 2 2
60 15 13 15 13 10 0 9 16 10 0 9 13 1 9 2 11 13 10 0 9 15 4 13 9 1 10 9 9 3 15 4 13 0 9 1 3 10 9 4 4 13 7 0 9 7 9 2 15 4 13 1 10 9 9 7 3 0 9 2 2
2 8 8
3 12 12 9
2 11 2
19 15 4 13 16 13 10 9 9 9 1 0 11 9 2 1 10 9 2 2
9 4 15 13 9 2 9 2 9 2
1 11
18 4 15 13 9 16 15 14 13 1 10 9 16 15 13 1 11 11 2
38 15 13 14 0 15 13 0 14 13 15 1 10 9 2 3 2 15 13 0 15 4 14 13 9 0 14 13 7 16 15 13 15 4 13 0 1 15 2
2 8 8
3 12 12 9
17 11 7 15 4 13 14 13 1 11 1 11 7 11 1 10 9 2
13 15 13 14 13 3 0 9 16 0 13 9 9 2
11 15 4 13 11 11 7 15 9 1 9 2
15 15 4 13 14 13 10 9 1 15 1 10 9 7 3 2
24 6 13 15 13 1 15 9 7 16 15 13 0 14 13 1 0 1 12 1 15 1 12 9 2
2 13 15
1 3
2 8 8
3 12 12 9
3 0 9 2
14 11 13 14 13 3 3 13 10 9 1 9 2 8 2
20 15 13 14 13 1 11 12 2 13 15 4 13 14 4 13 9 3 1 11 2
1 11
2 11 11
3 12 12 9
2 11 2
15 3 13 14 13 3 15 13 1 10 9 7 9 1 11 2
5 9 1 15 9 2
4 11 11 9 12
41 16 15 13 0 2 15 13 10 9 1 10 9 9 1 10 0 9 16 13 9 9 2 15 13 1 15 1 11 2 10 15 13 4 13 3 0 1 10 9 9 2
30 15 4 14 13 3 15 13 3 2 15 4 14 13 10 9 1 11 2 7 15 4 13 1 1 11 11 16 15 13 2
3 11 11 11
3 12 12 9
22 15 4 13 11 9 9 2 11 9 1 9 7 10 9 1 9 9 9 1 11 11 2
18 15 4 3 13 10 0 9 1 0 9 7 10 11 0 9 9 9 2
9 15 4 13 12 9 1 10 0 2
6 13 15 15 15 13 2
1 11
3 0 9 2
28 9 3 2 11 12 1 11 12 2 13 15 13 1 10 9 15 13 7 13 3 1 9 10 9 16 15 13 2
3 12 9 9
9 11 11 12 2 13 11 3 12 9
14 11 11 12 2 13 11 0 9 2 13 1 9 1 11
6 2 13 11 1 9 2
16 13 9 7 13 1 0 9 2 0 1 12 9 3 2 2 13
14 11 11 12 2 13 1 0 9 2 13 11 2 11 2
23 11 11 12 2 13 1 11 11 2 1 11 2 11 7 0 0 9 2 13 2 1 8 9
6 11 11 12 2 11 11
6 11 11 12 2 11 11
14 11 11 12 2 13 1 11 2 13 9 2 13 1 11
5 11 11 12 2 11
15 11 11 12 2 11 2 9 7 11 2 0 9 9 9 2
19 11 11 12 2 11 2 11 2 11 14 9 2 12 2 12 9 9 9 2
5 11 11 12 2 11
21 11 11 12 2 11 1 11 1 9 2 3 1 11 9 2 2 13 11 0 9 2
10 11 11 12 2 11 2 9 1 11 2
18 11 11 12 2 13 11 1 11 2 13 1 9 2 13 1 12 9 2
13 14 13 9 3 3 0 2 15 13 12 11 11 2
21 15 13 10 9 15 13 1 15 13 1 10 11 11 1 11 2 13 1 11 2 2
23 3 2 15 4 14 3 15 9 1 15 3 2 15 13 14 13 10 9 1 10 9 2 2
19 16 15 3 13 15 2 4 15 13 15 1 15 1 2 11 11 11 2 2
7 15 4 13 9 1 15 2
5 9 1 10 9 2
2 9 2
8 13 4 10 9 1 11 11 2
16 11 13 10 0 9 10 13 10 9 1 15 9 1 10 11 2
19 13 16 10 9 9 13 1 11 9 2 7 10 9 4 13 1 0 9 2
15 6 13 10 9 1 11 11 7 15 4 13 1 10 9 2
9 6 13 10 9 1 15 3 3 2
5 13 10 0 9 2
1 11
5 2 9 2 9 2
2 11 2
9 15 13 15 10 9 9 1 11 2
42 15 13 1 10 11 9 7 13 10 9 2 0 1 15 9 13 0 2 10 9 9 9 1 15 4 13 11 9 7 3 9 2 7 15 13 10 0 0 9 15 13 2
1 11
2 6 2
11 13 4 11 14 0 9 1 10 9 9 2
15 11 11 4 13 11 14 0 9 1 2 9 1 10 9 2
20 4 15 6 13 10 0 9 1 10 9 1 11 2 11 2 11 7 15 9 2
23 16 15 13 0 1 15 2 15 4 13 14 13 15 3 3 16 0 16 15 13 10 9 2
1 9
1 11
2 11 2
8 6 13 13 10 11 9 9 2
11 15 4 13 10 9 9 1 11 16 13 2
19 15 4 3 13 10 9 1 10 9 9 9 1 12 9 3 1 12 9 2
7 2 9 12 7 12 2 2
10 15 4 13 10 9 1 9 1 9 2
16 16 10 9 13 0 1 15 4 15 6 13 7 13 1 9 2
15 16 15 13 10 9 6 4 14 13 14 13 15 10 9 2
2 9 2
30 11 11 0 9 11 11 12 11 11 11 2 11 12 2 9 2 12 2 12 12 9 2 12 2 12 12 9 12 12 12
9 2 8 8 8 8 8 8 9 2
7 13 1 15 9 10 9 2
2 9 2
15 9 9 1 11 1 12 9 1 11 14 9 2 11 9 2
2 11 2
20 13 1 15 0 9 4 10 9 9 11 11 1 11 7 11 11 11 11 11 2
10 6 13 16 10 0 9 4 4 13 2
14 6 13 15 13 16 15 13 10 9 7 13 9 0 2
2 11 9
2 11 2
7 3 13 9 1 10 11 2
1 11
2 9 2
18 15 4 4 13 9 16 9 4 13 16 10 2 11 11 2 4 13 2
21 0 14 13 16 15 13 3 0 7 13 10 0 9 2 7 16 9 4 13 3 2
10 13 3 16 13 9 1 10 0 9 2
14 15 13 15 10 4 13 14 13 3 0 9 1 15 2
22 13 15 4 4 13 1 9 2 16 15 13 16 15 4 14 4 13 0 1 10 9 2
4 3 2 9 2
28 10 12 0 9 4 14 13 3 0 15 13 14 13 10 10 0 9 2 7 15 13 0 15 4 13 1 3 2
2 13 9
1 11
4 9 7 9 2
24 15 13 3 14 13 15 13 16 11 13 9 1 9 12 1 11 2 9 11 2 1 15 9 2
11 11 11 2 1 12 9 2 12 9 12 9
8 11 11 2 12 9 2 12 9
11 11 11 2 12 9 2 12 9 12 9 2
48 16 0 2 15 13 3 2 3 0 2 7 3 0 2 15 13 1 10 0 9 1 0 9 2 7 15 4 3 13 1 3 1 10 12 1 12 9 2 16 15 4 13 3 7 13 15 9 2
9 11 13 0 2 3 2 3 0 2
6 10 10 0 7 0 9
1 11
2 6 2
20 13 4 10 9 9 9 1 10 1 10 11 7 11 11 11 15 3 13 15 2
1 11
2 11 2
19 15 4 13 10 0 7 13 9 1 10 13 9 13 10 9 1 9 9 2
11 15 4 13 14 13 15 14 13 15 0 2
29 3 11 11 4 13 16 13 15 16 15 13 0 15 13 3 0 1 10 9 11 11 13 15 9 13 16 15 13 2
13 13 15 13 16 15 13 10 9 7 13 9 0 2
2 11 9
7 13 1 15 9 10 9 2
4 6 2 11 2
2 9 2
1 11
5 11 11 0 0 9
3 11 11 2
24 15 4 13 1 13 10 9 1 15 9 1 10 9 1 9 1 11 10 15 13 1 11 11 2
19 6 4 14 13 14 13 7 11 11 2 11 7 15 1 10 9 7 9 2
8 15 13 3 16 13 15 9 2
5 11 11 0 0 9
3 11 11 2
18 13 4 10 0 7 13 9 1 15 9 1 9 2 10 13 15 9 2
27 6 4 14 13 14 13 7 11 11 2 11 2 0 9 2 12 2 8 2 7 15 1 10 9 7 9 2
6 13 15 1 15 9 2
5 11 11 0 0 9
2 11 2
14 15 13 10 9 1 11 11 11 2 11 1 15 9 2
9 4 15 13 3 1 10 0 9 2
2 9 2
1 11
2 11 2
22 1 15 9 9 9 2 13 4 13 9 1 10 9 7 10 9 12 3 1 10 9 2
54 4 13 1 11 11 2 15 4 13 16 15 13 3 12 9 1 9 1 10 9 1 5 12 12 10 2 12 1 11 11 11 11 1 2 9 2 1 11 2 7 12 1 11 11 1 2 9 2 1 11 11 11 11 2
36 15 4 13 16 15 0 9 9 13 14 13 10 9 9 1 5 12 12 1 10 9 2 7 1 9 16 15 4 13 14 13 10 13 9 3 2
12 13 15 13 16 15 13 15 9 2 3 3 2
28 16 15 4 13 10 9 14 13 10 13 2 6 13 15 10 13 2 1 9 7 15 4 13 15 9 1 3 2
12 4 15 13 10 9 2 13 0 14 13 15 2
7 15 4 4 13 1 12 2
17 10 9 9 4 4 13 1 11 11 2 15 4 4 13 1 12 2
8 15 13 3 16 13 1 15 2
2 11 11
26 2 13 13 9 2 8 8 8 8 8 8 9 2 2 13 13 9 2 8 8 8 8 8 8 9 2
8 2 8 8 8 8 8 8 9
8 2 8 8 8 8 8 8 9
2 6 11
18 4 15 13 10 9 14 13 10 9 1 9 10 15 4 13 10 9 2
8 9 2 15 13 15 13 0 2
1 11
2 11 2
22 13 13 10 9 9 1 10 11 9 9 2 3 1 9 12 1 10 11 9 9 9 2
20 15 4 13 10 9 9 1 10 9 9 1 15 3 3 16 15 13 10 9 2
13 13 15 13 16 15 13 10 9 7 13 9 0 2
2 11 9
3 6 9 2
62 15 3 13 1 10 9 1 11 7 15 13 15 3 14 13 10 9 1 10 9 1 9 9 1 9 1 0 9 7 15 3 13 15 13 3 14 13 10 0 9 9 0 2 16 9 4 13 10 9 9 9 4 3 3 13 1 16 9 4 4 13 2
39 4 15 13 16 1 11 7 1 10 0 9 1 11 15 4 14 13 9 7 3 13 9 1 10 13 3 9 2 7 13 9 4 13 1 1 9 9 2 2
42 16 15 13 10 9 15 4 13 9 14 13 15 1 11 14 13 16 10 9 4 3 13 15 1 16 15 13 10 0 9 1 0 9 1 11 12 10 4 14 13 1 2
13 13 15 13 16 12 1 15 4 13 15 13 15 2
2 11 2
19 3 2 15 10 9 10 11 11 4 13 0 1 1 10 9 1 9 3 2
22 15 13 10 9 13 1 10 9 1 10 9 9 7 15 4 3 13 1 10 9 9 2
1 11
4 11 2 11 2
11 15 4 3 13 3 1 10 9 9 9 2
20 15 13 16 15 4 13 10 9 2 9 9 1 9 10 4 13 10 0 9 2
6 15 4 13 15 0 2
12 11 2 15 13 3 10 9 1 15 0 9 2
18 15 4 13 3 1 15 3 3 16 15 13 0 9 2 3 3 9 2
16 11 11 11 0 9 9 11 11 2 11 2 11 2 12 2 12
12 10 9 9 15 4 13 1 1 11 13 12 2
30 15 4 13 1 10 9 9 9 7 10 1 10 5 12 9 13 1 10 9 7 10 5 12 9 13 3 1 10 9 2
24 4 14 10 10 9 9 1 10 9 1 10 9 13 10 9 2 13 0 9 2 1 10 9 2
9 10 9 9 1 10 9 13 0 2
1 11
2 11 2
38 15 4 14 13 14 13 1 9 9 2 13 15 13 10 9 3 7 1 10 11 12 0 9 2 13 15 13 10 9 1 11 16 15 13 1 11 9 2
3 6 9 2
62 15 3 13 1 10 9 1 11 7 15 13 15 3 14 13 10 9 1 10 9 1 9 9 1 9 1 0 9 7 15 3 13 15 13 3 14 13 10 0 9 9 0 2 16 9 4 13 10 9 9 9 4 3 3 13 1 16 9 4 4 13 2
39 4 15 13 16 1 11 7 1 10 0 9 1 11 15 4 14 13 9 7 3 13 9 1 10 13 3 9 2 7 13 9 4 13 1 1 9 9 2 2
42 16 15 13 10 9 15 4 13 9 14 13 15 1 11 14 13 16 10 9 4 3 13 15 1 16 15 13 10 0 9 1 0 9 1 11 12 10 4 14 13 1 2
13 13 15 13 16 12 1 15 4 13 15 13 15 2
2 11 2
19 3 2 15 10 9 10 11 11 4 13 0 1 1 10 9 1 9 3 2
22 15 13 10 9 13 1 10 9 1 10 9 9 7 15 4 3 13 1 10 9 9 2
1 11
4 11 2 11 2
11 15 4 3 13 3 1 10 9 9 9 2
20 15 13 16 15 4 13 10 9 2 9 9 1 9 10 4 13 10 0 9 2
6 15 4 13 15 0 2
12 11 2 15 13 3 10 9 1 15 0 9 2
18 15 4 13 3 1 15 3 3 16 15 13 0 9 2 3 3 9 2
16 11 11 11 0 9 9 11 11 2 11 2 11 2 12 2 12
12 10 9 9 15 4 13 1 1 11 13 12 2
30 15 4 13 1 10 9 9 9 7 10 1 10 5 12 9 13 1 10 9 7 10 5 12 9 13 3 1 10 9 2
24 4 14 10 10 9 9 1 10 9 1 10 9 13 10 9 2 13 0 9 2 1 10 9 2
9 10 9 9 1 10 9 13 0 2
1 11
21 0 14 13 1 10 9 1 1 10 0 9 2 15 4 13 1 15 3 3 10 9
17 6 2 3 16 15 4 13 15 9 2 15 3 4 13 0 9 2
33 15 4 13 14 3 13 3 1 15 1 11 2 11 12 1 12 9 5 12 9 2 9 2 14 13 1 15 9 9 1 11 11 2
32 15 4 13 1 1 15 12 2 12 9 9 7 15 13 15 9 4 13 15 13 15 13 3 7 15 4 4 13 1 15 9 2
21 1 15 1 15 1 11 2 15 13 16 3 13 0 14 13 15 1 15 9 9 2
21 3 2 16 15 4 13 1 12 9 14 13 2 13 3 7 13 9 7 13 15 2
9 15 4 13 15 9 1 1 9 2
8 15 4 13 9 9 9 12 2
17 6 13 15 13 16 7 3 15 4 13 16 15 4 13 0 9 2
2 9 2
3 4 13 0
28 3 13 15 9 14 13 10 9 7 9 9 9 13 1 11 2 11 9 1 12 9 2 12 9 11 9 2 2
10 10 9 4 14 13 0 1 12 9 2
9 10 11 9 4 4 9 13 3 2
2 9 2
1 11
15 13 15 13 1 11 2 16 15 4 13 14 13 10 9 3
18 13 4 10 13 9 9 10 13 15 9 9 1 11 11 3 10 9 2
31 15 13 15 13 10 9 9 1 11 11 1 11 11 12 1 12 9 11 9 14 13 10 9 1 9 2 9 15 4 13 2
38 3 2 4 15 1 15 15 4 14 13 1 15 1 9 13 15 9 1 10 9 1 10 15 12 9 4 13 14 13 9 9 1 10 9 13 1 15 2
16 13 4 10 9 15 3 13 1 15 1 11 12 1 10 9 2
10 2 9 2 8 8 8 8 8 9 2
2 9 2
1 11
2 11 2
14 10 9 13 10 9 15 13 1 15 9 10 0 9 2
10 15 4 3 13 10 13 9 13 9 2
2 9 2
1 11
9 2 8 8 8 8 8 8 9 2
10 2 8 8 8 8 8 8 8 9 2
19 2 8 8 8 8 8 8 9 2 9 2 8 8 8 8 8 8 9 2
21 2 8 8 8 8 8 8 8 9 2 9 2 8 8 8 8 8 8 8 9 2
1 6
3 6 11 2
27 1 9 1 9 12 2 9 12 2 9 2 2 4 15 13 14 13 10 0 13 9 1 9 1 0 9 2
2 9 2
1 11
7 2 11 11 2 2 8 2
3 12 12 9
4 6 13 1 11
2 9 2
27 11 4 4 13 10 9 1 11 11 11 11 1 11 2 11 12 2 12 1 10 0 11 11 11 1 11 2
38 15 4 4 13 14 13 3 3 5 12 3 9 9 4 13 1 5 12 5 5 12 1 9 2 5 12 12 9 1 9 2 13 1 10 9 1 9 2
10 15 4 3 13 0 9 1 12 9 2
14 16 15 13 0 16 13 6 13 15 3 3 16 0 2
10 10 0 9 4 13 1 15 15 13 2
18 15 13 9 7 9 1 3 3 1 9 1 11 2 11 12 2 12 2
7 6 13 15 1 10 9 2
3 13 15 2
10 11 11 9 1 9 11 2 12 2 12
2 9 2
9 9 13 3 0 16 15 4 13 2
12 0 1 9 7 3 3 13 3 16 13 3 2
2 0 2
1 11
9 15 4 13 15 3 15 13 15 2
19 13 1 10 0 9 14 13 10 9 1 11 7 11 3 1 1 11 12 2
2 9 2
42 15 13 0 15 13 14 13 2 1 1 11 2 15 4 4 13 15 2 7 15 4 13 10 9 2 9 3 3 13 1 9 15 13 1 10 9 1 11 1 9 3 2
6 13 15 13 1 11 2
10 15 4 13 1 11 7 4 13 15 2
2 0 2
1 11
5 11 11 2 8 2
3 12 12 9
2 11 2
20 3 2 15 13 10 0 9 1 10 9 9 1 11 1 11 7 11 8 8 2
15 15 13 15 4 13 11 14 9 9 1 9 1 10 9 2
33 15 4 13 1 1 11 7 11 1 10 9 0 9 2 9 9 7 11 9 2 9 9 2 7 13 15 13 16 15 13 0 9 2
16 15 13 9 1 10 0 9 9 7 4 3 13 1 10 11 2
9 13 15 13 10 9 13 1 15 2
30 3 2 4 15 13 10 0 9 2 9 9 2 9 1 10 0 9 1 11 14 9 2 11 11 2 11 2 11 11 2
2 9 2
5 11 11 11 7 11
23 13 1 15 9 4 9 9 9 1 10 11 11 11 9 15 4 13 1 1 11 1 11 2
9 10 9 2 9 2 8 4 13 2
2 9 2
8 6 2 15 4 13 14 13 2
2 9 2
4 9 10 12 2
5 13 1 15 3 2
3 8 8 8
3 12 12 9
10 3 13 10 9 16 13 3 2 9 2
1 11
2 11 11
3 12 12 9
17 10 13 2 3 9 7 9 1 10 12 12 9 9 13 16 13 2
9 9 4 13 10 9 0 9 12 2
17 10 10 0 9 4 4 13 14 13 15 9 9 2 10 13 12 2
19 11 2 15 9 9 2 9 12 2 16 13 10 9 0 9 4 13 12 2
29 15 4 13 1 12 0 9 7 4 9 0 13 14 13 3 2 15 4 13 3 1 10 9 9 7 1 9 9 2
9 10 9 1 10 9 13 12 9 2
10 10 9 4 13 16 9 4 13 1 2
12 6 13 15 13 16 10 1 15 13 0 9 2
2 9 2
6 11 11 11 2 11 9
59 13 1 15 9 4 9 1 10 9 9 10 4 13 9 1 10 11 11 11 2 11 11 11 9 2 13 10 9 1 9 1 10 0 9 10 4 13 1 12 9 1 10 0 9 2 10 0 9 9 15 2 7 10 0 9 1 10 9 2
24 16 10 9 1 10 9 7 9 9 13 14 3 0 3 2 15 4 14 4 13 1 10 9 2
29 0 9 1 10 0 9 2 13 10 9 7 9 9 2 4 4 13 9 1 11 9 1 10 9 1 10 9 9 2
33 0 13 9 4 13 0 1 10 0 9 7 3 7 15 4 13 15 0 1 10 1 15 2 3 13 15 13 3 0 9 15 13 2
16 15 4 13 14 13 10 1 10 9 15 13 1 10 9 9 2
21 15 4 3 13 0 9 2 9 7 9 1 10 9 1 10 9 2 7 15 13 2
54 15 3 13 10 9 1 10 9 10 13 9 9 2 0 7 0 9 2 0 9 2 9 2 9 2 0 9 9 2 9 9 2 9 2 9 2 9 2 9 9 2 0 9 2 9 2 7 9 0 9 2 1 9 2
26 16 15 4 13 0 1 15 9 2 15 3 4 13 1 10 9 16 13 15 9 0 1 11 12 9 2
20 9 4 3 4 13 7 15 4 13 10 9 9 3 10 9 14 13 0 9 2
8 3 3 16 13 1 15 9 2
11 3 3 2 13 15 10 1 10 0 9 2
37 2 9 2 2 9 2 2 2 9 2 2 9 2 2 9 2 2 9 2 2 9 2 2 9 2 2 8 8 8 9 2 2 9 2 2 9 2
2 2 9
2 2 9
2 2 9
2 2 9
2 2 9
2 2 9
2 2 9
2 2 9
5 2 8 8 8 9
2 2 9
2 2 9
2 11 11
50 11 11 9 1 9 9 7 9 9 9 11 11 1 11 11 11 11 11 1 11 12 11 11 11 2 11 12 11 2 11 12 2 9 2 12 2 9 2 12 2 9 2 12 8 9 2 8 9 2 8
26 13 4 10 0 9 1 15 9 9 1 10 9 15 4 13 1 1 10 11 9 1 11 1 11 9 2
21 4 13 1 0 9 9 2 7 11 2 1 9 7 13 15 4 13 10 2 3 2
9 9 1 9 2 2 9 9 2 2
54 9 13 14 2 3 2 2 13 11 11 14 7 11 11 14 13 9 16 8 2 11 14 9 14 13 4 13 3 1 9 1 10 9 1 9 7 8 2 10 9 13 14 13 1 10 9 1 13 2 7 2 13 9 2
12 10 11 9 9 13 0 14 13 10 9 3 2
5 9 4 3 13 2
2 0 2
1 11
2 11 2
22 16 15 13 9 2 11 7 15 13 7 15 13 16 10 9 13 0 14 13 1 11 2
17 15 4 13 14 13 10 9 1 10 9 15 13 1 11 0 9 2
13 15 4 13 16 15 4 13 14 13 10 13 9 2
5 15 3 13 15 2
23 13 15 13 7 15 4 13 15 2 7 13 10 0 9 15 4 13 14 13 1 10 9 2
11 15 9 13 1 11 1 1 12 1 11 2
2 0 2
1 11
16 11 13 15 4 3 13 1 12 9 7 15 13 0 2 13 2
2 11 11
3 12 12 9
1 3
2 0 11
8 11 13 15 14 13 1 15 2
17 16 15 13 2 10 9 9 13 3 0 7 3 13 1 0 9 2
35 3 2 10 9 9 9 10 13 10 9 9 1 10 9 1 10 9 3 15 13 15 4 14 13 15 9 14 13 9 16 13 10 9 9 2
47 13 10 0 2 16 15 13 0 9 1 10 9 11 2 10 13 10 9 10 15 13 1 2 9 3 3 1 15 0 9 2 2 15 4 13 16 10 9 1 10 9 11 11 13 3 0 2
20 3 2 16 15 13 10 0 9 1 10 1 2 9 9 2 15 4 4 13 2
7 15 13 10 0 13 0 2
2 11 11
2 11 2
11 16 15 4 13 1 15 1 10 9 2 9
1 11
2 11 11
2 12 12
12 4 12 1 15 13 15 10 0 9 14 13 2
5 15 13 1 9 2
2 9 2
30 15 13 15 4 1 10 9 3 13 1 2 11 2 13 1 9 2 7 11 2 9 2 2 8 3 13 15 0 9 2
15 15 13 15 13 0 16 3 11 14 13 2 11 2 9 2
2 11 11
2 12 12
2 11 2
11 4 15 6 13 15 10 9 14 13 9 2
14 8 4 15 13 16 15 13 10 9 1 2 11 2 2
4 8 2 11 2
13 16 15 4 13 2 3 13 15 0 14 13 11 2
2 9 2
1 11
1 5
5 10 9 13 0 2
17 15 4 3 13 0 7 3 13 1 9 9 9 7 0 0 9 2
34 16 15 4 13 15 1 9 6 13 15 13 1 9 7 3 13 15 1 15 9 2 15 4 14 13 10 9 7 13 15 9 1 9 2
1 5
41 1 15 9 1 11 10 9 2 15 4 13 10 13 9 1 10 0 9 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 11 2 7 11 2
12 3 13 10 9 2 3 13 14 13 10 9 2
27 9 10 13 4 13 14 13 9 9 2 11 2 11 2 11 2 11 2 11 2 10 11 2 7 10 11 2
50 9 10 4 14 13 14 13 9 9 13 2 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 7 10 11 2
33 1 9 13 1 10 0 9 2 15 4 13 0 16 15 14 13 1 1 10 9 13 1 10 13 9 2 8 11 7 11 9 2 2
13 15 4 13 14 4 13 1 10 9 1 9 9 2
13 6 13 15 13 16 15 13 10 9 1 10 9 2
5 13 1 2 11 11
39 6 2 15 4 13 9 1 9 9 7 2 7 9 9 7 0 9 9 1 10 11 11 2 11 2 2 11 11 2 11 11 2 7 11 11 2 11 2 2
2 9 2
1 11
35 1 9 1 15 0 9 1 10 9 1 9 15 13 14 13 1 2 4 15 14 13 14 13 10 0 9 0 2 0 9 9 2 9 9 2
2 11 11
3 12 12 9
10 6 13 13 9 14 9 9 1 12 2
1 9
1 11
5 15 13 10 0 2
10 3 4 15 3 13 14 13 15 9 2
25 15 4 13 10 0 9 1 10 11 9 9 1 11 12 1 12 1 11 1 10 11 1 12 11 2
16 10 9 1 10 9 13 10 0 9 1 10 0 9 9 9 2
12 15 4 13 0 16 11 7 11 11 4 13 2
9 3 15 4 13 15 10 0 9 2
36 15 4 13 10 9 1 10 11 11 11 9 13 1 11 11 2 10 13 10 0 9 9 2 16 15 4 14 13 14 13 10 9 1 10 9 2
19 11 11 4 14 13 10 9 16 10 9 3 2 7 15 4 13 0 9 2
26 15 4 13 14 13 15 1 13 2 16 11 11 4 13 2 7 15 3 13 15 14 4 13 1 11 2
11 4 15 13 15 13 3 7 3 1 15 2
3 0 9 2
20 15 4 13 10 13 9 1 10 9 9 1 11 2 11 13 11 12 2 12 2
21 10 9 13 10 9 9 13 1 9 2 9 2 1 10 9 9 1 10 9 9 2
5 9 4 4 13 2
22 13 10 0 9 16 11 11 2 10 9 2 4 14 13 15 14 13 9 7 9 9 2
29 15 13 15 13 10 9 1 10 13 9 16 11 13 10 9 9 9 3 2 7 15 3 4 14 13 15 3 3 2
16 15 4 14 3 16 15 13 1 10 9 9 7 15 13 1 2
26 3 15 13 10 9 2 15 4 13 15 10 9 7 15 4 13 3 7 13 15 3 14 13 10 9 2
43 15 13 1 11 14 13 10 9 16 15 15 4 13 14 4 13 1 10 9 1 9 9 2 7 15 13 16 15 0 9 13 16 10 1 10 9 4 4 13 1 1 11 2
7 15 13 15 1 11 11 2
20 15 3 13 16 11 4 13 14 4 13 12 9 14 13 1 10 9 9 9 2
2 6 2
9 11 2 4 15 13 15 7 11 2
2 11 11
3 12 12 9
3 6 11 2
23 15 13 10 9 9 1 10 0 9 7 12 1 15 9 13 10 9 1 15 0 9 9 2
15 10 9 13 11 11 2 7 15 9 13 1 10 13 9 2
13 4 15 13 10 9 1 15 7 13 15 10 9 2
2 9 2
18 11 2 16 13 15 4 13 11 14 13 9 1 10 11 0 9 9 2
20 15 13 3 16 13 1 10 3 0 9 1 10 0 7 0 9 1 9 9 2
1 11
7 2 13 13 9 2 9 2
2 2 9
19 15 4 13 10 13 0 9 1 9 9 9 13 1 1 11 12 2 12 2
13 10 9 13 10 11 11 11 11 9 1 10 9 2
5 9 4 4 13 2
14 9 9 2 15 4 13 13 10 9 1 10 9 3 2
2 11 11
3 12 12 9
10 6 13 13 9 14 9 9 1 12 2
2 9 2
1 11
9 3 13 10 9 1 10 0 9 2
2 11 11
3 12 12 9
10 6 13 13 9 14 9 9 1 12 2
1 9
1 11
2 6 2
2 3 2
32 15 3 13 10 9 1 11 7 11 7 15 13 15 15 13 10 0 9 10 9 14 13 10 0 9 9 14 13 0 0 9 2
11 15 4 13 14 13 1 15 1 10 11 2
7 6 9 2 13 11 3 2
2 11 11
3 12 12 9
10 6 13 9 13 10 9 9 1 12 2
1 9
1 11
2 11 11
3 12 12 9
11 6 13 13 10 3 0 9 1 11 11 2
14 1 9 10 13 9 9 7 0 9 9 13 1 9 2
24 0 9 4 4 13 7 10 9 4 4 3 13 2 7 1 9 9 9 7 8 0 9 2 2
9 6 13 15 16 15 13 10 0 9
1 11
2 11 11
2 12 12
60 10 9 1 10 9 7 9 13 1 15 0 9 2 13 13 9 2 13 14 13 10 0 9 9 9 1 0 9 9 2 9 7 9 7 9 10 0 9 1 9 1 9 9 0 9 9 7 9 9 9 0 9 7 10 9 1 10 11 0 9
77 1 10 0 9 1 9 2 13 9 1 10 9 9 2 10 0 9 1 10 9 1 9 9 9 2 7 9 1 10 9 1 10 0 9 9 9 13 0 16 15 13 3 14 0 16 13 0 0 9 1 9 14 13 15 9 9 2 10 1 10 0 9 13 10 0 9 9 1 9 7 0 9 1 0 9 9 2
19 3 15 13 14 13 15 1 2 7 2 7 13 15 9 1 2 10 13 2
7 15 4 13 1 9 10 13
27 16 9 9 1 10 13 9 9 4 4 13 1 1 9 9 2 1 7 1 13 9 1 9 1 9 9 2
41 16 15 13 9 9 1 9 9 9 2 9 1 9 9 7 10 0 0 9 9 2 10 9 4 1 0 14 13 7 4 13 14 4 13 1 9 1 10 9 9 2
26 10 9 1 10 0 9 9 9 9 13 1 15 0 9 10 4 3 4 13 7 13 2 13 9 9 2
31 10 9 1 10 9 9 9 2 3 1 0 0 9 2 1 0 11 9 15 13 14 13 3 0 9 14 13 10 3 13 9
25 10 9 1 0 0 2 11 2 9 15 4 2 13 2 0 0 9 9 9 3 13 10 13 11 9
23 10 9 9 1 5 12 12 13 1 10 13 9 7 10 0 9 9 16 13 1 10 9 2
29 15 4 13 14 13 0 9 1 10 9 9 2 1 10 9 1 9 7 9 9 9 2 1 10 9 9 9 9 2
23 3 2 10 9 4 13 14 4 13 16 13 10 0 9 7 9 1 9 9 9 1 9 2
34 10 9 1 10 9 9 1 0 11 7 9 1 9 9 2 13 3 3 0 2 16 9 4 3 13 7 0 0 9 9 4 4 13 2
8 11 11 9 4 13 13 16 13
55 10 9 9 13 1 9 1 9 9 2 1 0 9 1 9 1 0 9 9 1 9 2 9 10 9 1 10 9 7 0 9 9 1 10 9 2 13 13 9 9 1 1 9 9 2 2 13 0 9 1 9 9 1 0 9
14 9 1 9 9 1 9 7 9 9 9 1 9 0 9
14 0 9 9 1 10 9 9 10 4 4 13 1 11 9
13 9 9 1 9 9 9 13 10 0 3 13 9 9
15 10 9 1 11 0 9 7 9 1 15 9 9 7 9 9
12 10 9 2 9 0 9 13 1 9 1 9 9
11 15 4 13 1 9 3 1 10 9 13 9
1 9
1 11
2 11 11
2 12 12
20 0 0 9 4 13 1 10 9 1 10 9 1 9 9 1 10 11 11 9 2
24 9 13 10 9 1 10 1 9 9 9 2 2 9 2 2 10 13 12 9 1 10 9 9 2
20 10 9 13 1 10 9 1 9 14 9 1 10 9 3 1 10 9 9 9 2
34 10 9 1 10 9 1 2 9 2 1 10 9 11 9 2 13 1 10 9 1 9 13 9 2 10 13 10 0 9 16 13 10 9 2
28 10 9 14 13 10 0 9 7 9 9 9 1 10 9 1 10 0 9 1 10 9 1 11 2 7 9 2 2
15 10 0 9 9 1 11 4 13 7 4 13 1 9 9 2
20 10 0 9 14 13 9 9 9 1 10 11 9 3 1 10 0 0 9 9 2
38 0 9 9 4 13 7 4 13 13 14 13 9 2 13 9 1 9 9 7 14 13 9 1 0 9 1 1 10 9 1 10 9 9 7 9 9 9 2
38 10 9 1 9 1 10 11 9 4 4 13 7 3 13 1 10 0 9 2 0 9 2 9 9 2 9 13 14 13 0 9 1 9 1 9 11 9 2
25 10 9 2 9 9 9 9 9 1 10 9 4 13 16 16 14 13 10 0 9 1 1 9 9 2
26 11 11 4 13 10 0 0 9 9 9 9 13 9 9 2 9 9 1 9 9 9 1 10 11 9 2
26 10 13 9 9 9 4 4 13 0 1 9 9 13 0 9 2 9 9 7 13 9 1 9 7 9 2
33 10 0 9 9 4 13 0 1 10 9 2 3 9 4 4 13 14 13 0 11 2 11 9 1 1 10 9 7 13 9 9 9 2
40 9 9 1 0 9 9 7 9 4 4 3 13 7 10 9 9 4 13 0 1 10 9 1 9 13 10 9 1 12 9 13 1 0 9 1 10 9 1 9 2
26 10 9 1 10 0 9 9 4 4 13 1 10 9 9 9 13 10 0 9 9 1 9 9 7 9 9
16 10 0 0 9 9 9 4 4 13 1 10 9 9 9 10 13
14 10 0 9 1 9 9 2 7 9 1 9 9 1 11
30 9 1 0 1 10 0 9 9 2 1 0 9 9 2 3 15 13 10 9 16 9 9 4 14 4 13 1 10 0 9
28 0 9 3 1 9 9 9 1 10 0 0 7 0 9 9 2 9 13 10 0 9 9 13 1 1 10 9 2
9 0 9 7 9 1 9 9 9 9
28 0 9 1 9 1 10 9 1 11 9 2 3 13 9 1 9 10 15 13 9 14 13 2 7 1 9 11 9
22 10 9 13 9 9 2 13 1 9 9 2 3 0 2 7 10 0 8 0 9 9 9
21 10 0 9 1 9 1 0 2 9 9 2 7 0 9 2 9 2 9 1 9 2
6 10 0 9 1 0 9
9 10 0 0 9 1 9 7 9 9
15 15 13 14 13 0 9 1 10 9 1 10 0 9 1 11
10 16 15 13 10 9 6 13 15 1 9
1 9
1 11
3 11 11 2
17 15 4 13 14 13 15 16 3 13 10 9 14 3 13 15 9 2
22 16 15 13 0 1 10 9 15 13 3 0 14 13 10 11 11 11 1 11 0 9 2
34 15 13 3 0 10 9 4 13 2 7 15 13 16 1 15 9 9 2 9 2 9 2 0 9 2 8 16 15 4 13 1 15 9 2
31 16 13 1 11 11 2 11 2 11 7 11 2 15 13 0 16 10 9 13 10 0 9 14 13 10 9 15 4 13 1 2
41 15 13 3 0 16 10 9 13 10 0 9 16 13 10 0 9 2 9 9 2 3 15 13 15 14 13 16 15 4 13 14 13 15 15 13 14 13 3 0 9 2
35 15 13 16 13 12 7 12 9 9 9 9 1 10 11 1 11 10 9 7 9 14 13 1 10 9 9 16 15 4 13 1 10 9 9 2
9 15 3 13 16 13 10 11 9 2
34 1 1 15 9 2 15 4 13 10 0 9 2 7 15 13 0 14 13 1 10 9 16 15 4 13 0 1 10 11 11 11 1 11 2
26 15 4 13 14 13 3 1 11 10 9 14 13 1 15 14 3 13 15 9 9 7 14 3 13 15 2
24 16 15 13 1 9 0 15 4 13 14 13 15 0 9 9 1 0 9 2 6 13 15 13 2
10 13 9 7 13 14 13 1 15 3 2
2 3 2
2 11 11
3 11 11 2
18 15 4 13 14 13 15 16 13 10 9 14 13 15 1 10 9 9 2
10 1 10 9 2 10 9 13 14 0 2
38 15 13 16 15 13 10 0 9 2 7 15 13 16 1 15 9 9 2 9 2 0 9 2 8 2 16 15 4 13 15 9 7 3 13 1 15 9 2
29 16 13 1 15 7 11 11 2 11 7 11 2 15 13 0 16 11 13 10 0 9 14 13 13 1 9 2 9 2
39 15 13 3 0 16 11 13 10 9 16 13 10 0 9 2 9 9 2 3 15 13 15 14 13 16 15 4 13 14 13 15 15 13 14 13 3 0 9 2
34 15 13 16 13 12 7 12 9 9 9 9 1 10 11 1 11 10 9 7 9 14 13 1 10 9 9 16 15 4 13 1 10 9 2
11 15 3 13 16 13 14 13 10 11 9 2
38 1 1 15 9 2 15 4 13 10 0 9 2 7 15 13 0 14 13 1 10 9 9 16 15 4 13 1 10 9 1 10 11 11 11 11 1 11 2
13 9 3 16 13 10 9 14 13 7 13 1 15 2
23 15 4 13 10 9 13 15 7 15 13 15 4 13 14 13 1 9 7 9 1 10 9 2
27 3 2 16 15 4 13 1 9 0 15 4 13 14 13 15 0 9 9 1 0 9 2 6 13 15 13 2
10 13 9 7 13 14 13 1 15 3 2
2 3 2
2 11 11
3 11 11 2
18 15 4 13 14 13 15 16 13 10 9 14 13 15 1 10 9 9 2
10 1 10 9 2 10 9 13 14 0 2
37 15 13 16 15 13 10 0 9 2 7 15 13 16 1 15 9 9 2 9 2 0 9 2 8 2 16 15 4 13 15 9 7 3 13 15 9 2
29 16 13 1 15 7 11 11 2 11 7 11 2 15 13 0 16 11 13 10 0 9 14 13 13 1 9 2 9 2
40 15 13 3 0 16 11 13 10 9 16 13 10 0 9 2 9 9 2 3 15 13 15 14 13 16 15 4 13 14 13 8 15 15 13 14 13 3 0 9 2
34 15 13 16 13 10 9 1 9 9 9 9 1 10 11 1 11 10 9 7 9 14 13 1 10 9 9 16 15 4 13 1 10 9 2
11 15 3 13 16 13 14 13 10 9 9 2
37 1 1 15 9 2 15 4 13 10 0 9 2 7 15 13 0 14 13 1 10 9 9 16 15 4 13 10 9 1 10 11 11 11 11 1 11 2
21 3 2 15 4 13 14 13 15 9 13 13 10 9 2 9 0 9 9 1 11 2
22 15 13 16 1 15 9 2 0 7 9 9 9 16 15 4 13 13 9 1 10 9 2
18 15 13 3 0 1 9 2 9 7 13 16 15 9 13 10 3 0 2
13 9 3 16 13 10 9 14 13 7 13 1 15 2
25 15 4 13 10 9 14 13 1 15 7 15 13 15 4 13 14 13 1 9 7 9 1 10 9 2
26 3 2 16 15 13 1 9 0 15 4 13 14 13 15 0 9 9 1 0 9 2 6 13 15 13 2
10 13 9 7 13 14 13 1 15 3 2
2 3 2
2 11 11
9 13 15 13 16 15 13 10 9 2
1 9
1 11
13 0 1 15 2 15 4 13 1 10 11 11 9 2
1 9
1 11
21 6 13 15 10 11 9 10 13 10 9 10 15 13 13 1 10 9 9 9 9 2
23 15 13 14 13 0 16 15 13 3 3 15 13 13 10 9 7 3 10 9 4 4 13 2
9 1 0 2 6 13 10 13 9 2
20 4 15 4 13 2 13 10 9 1 0 9 9 7 10 9 1 0 9 9 2
16 10 9 9 4 15 13 10 9 1 2 11 11 7 11 11 2
20 6 13 15 10 0 9 9 10 15 4 13 1 5 5 9 14 13 10 9 2
38 10 9 4 15 13 14 13 10 9 2 0 9 7 0 9 7 10 9 1 10 12 2 16 13 6 13 15 10 9 15 13 14 13 10 12 9 2 2
25 10 9 9 4 15 13 2 8 2 1 0 9 9 10 9 1 10 0 9 2 7 1 0 9 2
13 10 9 4 15 13 2 12 5 0 1 12 9 2
13 4 15 13 10 9 9 1 10 9 1 10 9 2
15 4 15 13 10 2 9 2 0 9 9 14 13 10 9 2
14 4 15 13 10 5 5 9 9 9 9 1 15 9 2
8 4 11 13 10 13 9 9 2
12 10 9 4 4 13 7 9 7 3 3 9 2
23 11 2 7 11 2 6 13 9 1 10 9 1 13 9 16 16 15 13 0 9 1 9 2
13 13 15 10 3 3 1 15 9 7 9 3 3 2
58 3 2 15 4 13 14 13 16 9 14 9 2 0 16 13 10 9 9 2 13 14 13 12 5 0 16 2 2 8 2 10 9 10 4 4 13 13 0 1 10 0 9 2 7 2 8 2 10 0 9 1 10 9 9 9 9 13 2
19 15 13 9 14 13 10 13 9 1 10 9 1 10 9 7 3 7 3 2
2 9 2
1 11
14 11 2 15 13 10 9 15 13 15 10 9 9 1 2
50 9 12 1 10 11 11 11 9 2 10 15 4 13 1 15 3 2 1 11 13 11 14 2 13 1 0 9 1 11 2 14 13 10 0 9 10 4 3 4 13 15 1 9 9 9 1 11 14 9 2
76 15 13 10 3 0 9 3 15 13 10 9 16 11 4 14 13 0 14 13 15 1 10 9 9 9 2 3 15 13 10 13 3 9 1 10 11 4 13 14 2 13 2 11 2 16 13 10 0 9 14 13 10 0 9 7 4 13 0 7 13 2 11 2 0 1 10 9 7 9 2 13 1 10 0 9 2
30 15 4 13 1 15 16 15 13 10 5 12 12 10 11 13 3 13 1 15 9 14 2 13 2 15 16 13 10 9 2
29 1 10 9 9 2 15 13 14 13 0 16 15 4 13 9 15 4 14 13 10 9 1 10 9 14 13 0 9 2
11 4 15 13 9 15 4 13 15 3 3 2
33 15 4 13 3 3 3 1 11 16 15 4 14 13 3 0 9 14 13 10 9 16 15 13 2 7 13 15 13 15 15 4 13 2
42 11 4 13 16 12 9 9 13 10 9 1 10 9 9 2 15 13 1 11 7 11 2 10 4 13 11 14 13 1 15 10 9 16 3 14 13 10 0 9 1 11 2
29 15 13 1 10 9 9 1 11 2 7 16 15 13 15 15 4 13 2 13 15 13 7 15 4 13 1 10 9 2
2 9 2
1 11
2 11 11
3 12 12 9
21 4 15 6 13 11 11 7 13 10 11 11 11 11 1 9 1 10 9 9 9 2
36 15 9 13 16 11 13 14 13 10 9 14 13 11 14 0 9 1 9 16 15 14 13 10 9 14 13 13 10 9 1 11 14 9 9 9 2
28 15 4 14 13 9 1 10 9 10 4 13 3 3 1 0 0 9 1 5 12 1 10 9 1 11 1 11 2
22 0 9 4 4 13 1 10 9 1 10 9 2 10 15 4 14 13 0 14 13 3 2
23 10 9 4 13 5 12 1 9 16 15 13 14 13 10 9 16 15 4 1 11 7 11 2
25 0 9 2 7 15 13 0 15 4 13 16 15 9 4 3 13 1 10 9 1 9 7 0 9 2
44 15 4 13 14 13 1 9 16 15 13 0 9 9 2 15 13 1 10 9 2 7 16 15 13 14 13 10 9 10 13 10 0 9 1 9 7 9 2 15 4 4 13 3 2
15 9 1 15 13 2 7 3 3 2 10 13 9 13 14 2
22 15 9 9 3 13 16 15 4 13 10 0 13 9 16 10 9 13 1 9 7 9 2
18 15 13 1 15 9 15 13 0 1 15 7 15 4 13 15 13 3 2
1 11
43 15 3 4 13 13 1 10 0 9 9 16 13 3 1 10 8 8 9 9 1 10 9 7 15 3 13 16 10 0 9 4 13 16 10 9 7 13 9 4 4 13 1 2
46 15 9 16 13 10 9 3 13 2 4 15 4 13 16 3 9 13 10 9 4 7 4 13 1 10 9 2 16 15 3 13 11 7 11 7 16 15 13 15 4 4 13 10 0 9 2
2 11 11
3 12 12 9
31 1 9 1 10 0 9 15 13 16 10 0 9 4 13 1 10 13 11 9 7 1 10 12 0 13 9 9 15 4 13 2
14 16 15 13 10 9 15 13 14 13 3 1 15 3 2
3 6 13 2
1 11
23 1 9 1 11 2 15 13 15 4 13 0 14 13 15 3 1 10 9 1 9 7 9 2
27 3 2 16 15 4 13 2 10 9 15 13 1 13 3 0 2 7 15 13 15 13 9 1 10 1 15 2
26 12 9 13 14 13 3 10 9 1 10 9 9 7 3 13 3 1 10 0 12 9 16 15 4 13 2
7 6 13 15 15 9 3 2
1 11
2 6 2
4 3 15 13 2
2 9 2
1 11
5 3 13 10 9 2
10 13 4 15 9 1 10 9 1 9 2
12 15 13 11 11 14 7 11 11 14 0 9 2
28 6 13 15 7 13 15 13 16 15 13 10 9 1 7 1 11 9 2 15 4 13 1 1 10 9 11 2 2
3 13 15 2
2 6 2
1 11
2 11 11
3 12 12 9
18 6 13 11 14 13 9 9 7 13 1 9 1 10 9 2 1 15 2
2 9 2
5 13 14 13 15 2
1 11
2 11 11
3 12 12 9
2 6 2
1 11
2 11 11
3 12 12 9
18 6 13 11 14 13 9 9 7 13 1 9 1 10 9 2 1 15 2
2 9 2
14 11 2 4 15 13 10 9 1 9 1 9 1 15 2
23 11 11 13 10 0 9 0 9 7 15 13 15 10 9 2 15 3 13 12 2 3 2 2
5 11 2 10 9 2
2 11 11
3 12 12 9
21 11 11 4 13 9 14 13 10 11 9 1 10 1 15 9 2 1 12 7 12 2
15 10 0 9 4 13 14 13 1 9 9 2 10 15 13 2
27 0 9 1 11 3 13 10 9 1 9 2 7 15 3 2 16 3 2 13 10 9 16 15 13 3 0 2
10 10 9 13 5 12 1 9 7 9 2
7 6 13 10 9 1 12 2
2 9 2
10 6 2 15 13 11 1 1 10 9 2
2 11 11
3 12 12 9
14 11 2 4 15 13 10 9 1 9 1 9 1 15 2
23 11 11 13 10 0 9 0 9 7 15 13 15 10 9 2 15 3 13 12 2 3 2 2
5 11 2 10 9 2
2 11 11
3 12 12 9
21 11 11 4 13 9 14 13 10 11 9 1 10 1 15 9 2 1 12 7 12 2
15 10 0 9 4 13 14 13 1 9 9 2 10 15 13 2
27 0 9 1 11 3 13 10 9 1 9 2 7 15 3 2 16 3 2 13 10 9 16 15 13 3 0 2
10 10 9 13 5 12 1 9 7 9 2
7 6 13 10 9 1 12 2
2 9 2
22 15 13 15 13 10 9 1 10 11 11 9 1 9 13 11 12 10 11 14 9 13 2
13 15 13 10 11 9 1 11 7 13 15 1 15 2
45 11 7 15 13 15 9 16 13 10 13 9 1 11 7 11 13 1 11 14 9 2 7 16 9 13 2 11 7 15 13 3 14 13 15 1 11 7 13 15 14 13 10 13 9 2
29 16 15 13 2 11 7 15 4 3 13 15 1 1 11 1 11 11 7 3 13 10 9 1 13 9 1 10 9 2
30 11 4 3 13 10 9 1 3 0 9 15 13 1 10 9 1 11 7 11 1 10 9 16 3 3 14 13 10 9 2
7 6 2 15 13 0 9 2
4 10 10 9 2
16 4 14 13 15 10 9 7 12 13 15 0 1 15 0 9 2
1 11
2 11 2
13 15 13 0 16 13 10 9 16 13 10 0 9 2
11 13 15 9 1 15 9 7 9 1 9 2
24 15 4 13 10 9 16 13 9 13 3 7 15 13 14 13 0 16 15 13 15 13 1 9 2
1 11
6 4 15 13 14 13 2
1 11
28 10 0 9 1 10 11 9 1 9 4 4 13 1 11 2 11 12 2 1 10 11 11 11 1 11 2 11 2
19 10 9 4 4 13 1 9 1 10 0 9 1 15 11 1 10 11 11 2
17 2 6 13 15 3 13 9 8 1 0 9 1 10 11 11 2 2
31 13 10 9 9 1 11 2 15 4 13 14 13 1 9 1 10 11 11 1 10 11 9 9 7 9 2 13 10 9 9 2
21 9 9 4 3 13 14 13 1 10 0 9 1 10 11 11 1 11 2 11 12 2
25 1 1 10 0 0 9 0 1 11 1 10 0 9 1 15 9 2 10 11 11 3 4 3 13 2
15 3 2 15 4 13 10 9 1 9 1 10 0 11 11 2
22 14 13 12 1 10 9 2 15 4 13 10 11 9 16 15 13 9 1 10 11 9 2
26 16 15 4 13 14 13 9 1 10 0 9 2 6 13 3 3 16 15 13 0 9 1 10 13 9 2
18 15 4 4 13 10 11 9 0 1 9 1 10 11 11 1 11 12 2
24 16 15 13 10 9 7 13 10 9 3 3 2 6 13 11 11 1 12 7 11 11 1 12 2
11 15 4 13 3 16 13 15 1 11 12 2
3 9 9 2
21 11 11 11 12 11 11 11 11 11 12 9 2 12 7 12 9 2 12 9 2 8
22 11 11 11 12 11 11 11 11 2 11 12 9 2 12 7 12 9 2 12 9 2 8
2 0 2
4 13 15 0 2
8 16 3 2 15 4 13 15 2
3 9 11 2
2 8 8
3 12 12 9
3 0 11 2
17 15 4 13 9 1 11 11 11 1 9 1 10 0 11 9 9 2
16 11 11 13 15 4 4 13 1 11 11 14 9 9 2 8 2
11 4 15 13 15 14 13 10 9 1 15 2
4 13 15 13 2
3 0 9 2
1 11
26 11 11 0 9 9 9 11 12 11 11 2 11 9 12 11 2 11 12 12 12 2 9 2 9 2 8
9 2 13 9 2 9 0 9 2 2
6 15 13 3 10 9 2
1 11
18 4 15 13 16 15 13 3 1 11 1 10 11 9 3 15 13 1 2
6 11 11 2 11 11 2
15 10 13 9 1 10 9 9 1 9 7 9 4 13 3 2
28 6 13 7 13 10 9 15 13 1 11 12 2 3 3 1 10 0 9 13 1 10 9 9 0 1 10 9 2
10 6 13 10 13 1 9 7 9 9 2
13 10 9 1 9 7 9 4 4 13 13 10 9 2
13 2 11 2 8 9 2 9 2 11 2 8 9 2
4 11 7 11 2
17 4 15 13 10 9 10 9 2 3 11 1 12 2 14 13 15 2
1 11
7 15 4 13 10 0 9 2
17 15 4 4 13 3 3 14 13 10 9 16 15 13 7 13 9 2
12 11 4 4 13 15 1 10 0 0 9 9 2
18 15 4 13 0 16 13 10 9 1 10 0 9 7 11 7 13 9 2
23 10 9 13 3 3 0 1 9 9 10 4 13 10 9 2 13 0 9 7 13 10 9 2
6 0 2 9 4 13 2
16 15 15 13 1 1 9 7 4 14 13 1 9 4 3 13 2
29 15 15 13 1 7 13 2 7 4 14 13 1 10 13 9 7 10 0 11 9 9 2 9 9 2 8 4 13 2
15 11 7 15 13 1 10 9 1 11 7 4 13 0 9 2
8 11 7 15 3 13 1 15 2
19 11 11 13 10 9 9 1 11 11 7 13 15 14 13 10 11 9 13 2
35 2 3 16 15 13 0 9 14 13 1 11 2 15 13 15 9 7 15 13 16 16 9 4 14 13 1 11 2 10 9 4 13 0 2 2
18 11 11 7 11 11 2 1 10 11 9 2 4 3 13 1 9 9 2
15 15 4 4 13 1 10 9 9 0 9 7 13 15 13 2
14 15 13 10 0 9 9 9 13 1 11 9 7 9 2
10 10 9 4 13 14 13 13 9 3 2
17 15 3 13 1 9 13 11 9 7 11 14 11 11 7 11 11 2
26 10 9 4 13 1 10 9 7 15 13 10 9 14 13 10 0 9 1 11 14 13 1 11 7 11 2
24 3 16 11 13 14 10 9 1 11 11 2 15 13 0 9 14 13 1 7 13 10 0 9 2
13 11 13 1 11 1 11 2 7 13 0 1 9 2
12 15 4 13 1 10 9 1 11 1 12 9 2
12 4 15 13 10 9 10 13 1 15 14 13 2
13 11 13 1 10 11 9 9 11 1 12 1 12 2
15 15 13 0 1 11 14 11 9 9 2 13 15 0 3 2
18 15 13 0 2 15 4 13 10 0 9 2 11 4 13 10 0 9 2
3 9 2 11
4 11 7 11 2
33 13 1 0 9 2 11 11 13 16 15 13 9 4 13 1 11 1 10 0 9 9 7 9 1 0 9 13 14 0 1 13 9 2
29 11 13 14 13 10 9 14 3 13 15 9 3 1 10 11 7 11 9 16 15 4 13 10 9 7 15 13 9 2
32 16 11 13 10 9 1 11 2 7 1 1 9 9 7 0 9 9 9 2 15 4 13 10 0 9 1 9 7 1 11 11 2
17 3 0 2 10 0 11 9 13 10 9 3 3 16 13 10 9 2
15 13 15 13 15 14 13 0 9 10 4 13 10 0 9 2
28 11 7 11 2 15 13 16 15 13 10 0 9 16 15 14 13 1 10 0 12 5 12 9 14 13 10 9 2
12 15 4 13 14 13 15 1 15 1 11 9 2
14 15 13 0 1 12 9 1 11 1 11 14 9 9 2
1 11
2 3 2
8 15 4 13 14 13 1 11 2
1 11
64 1 10 9 1 10 9 11 7 15 13 1 11 7 11 10 9 1 9 3 2 15 4 13 9 14 13 10 0 9 10 4 13 15 14 13 0 9 1 9 9 9 2 7 3 9 9 2 1 10 9 10 4 4 13 1 10 11 9 9 13 1 10 9 2
37 15 13 10 9 10 4 13 10 0 9 7 9 1 10 9 2 9 2 8 1 10 9 1 10 9 9 3 3 1 15 15 4 13 3 0 9 2
14 15 4 13 10 9 9 15 7 15 9 4 3 13 2
15 0 9 13 14 4 13 1 2 7 15 4 13 15 13 2
21 1 10 9 2 4 15 6 13 10 9 1 15 9 1 15 15 4 13 0 9 2
7 15 4 15 13 14 13 2
1 11
3 8 8 8
3 12 12 9
27 15 4 13 1 15 9 10 9 1 11 11 15 13 10 0 9 16 13 0 9 1 0 9 1 9 9 2
8 11 4 13 3 1 10 9 2
23 15 13 15 0 9 1 10 9 1 10 11 7 11 11 1 11 9 1 10 11 1 11 2
30 10 9 1 0 9 1 9 9 7 0 9 4 13 11 14 13 0 9 1 15 9 9 7 13 10 9 1 9 9 2
17 6 2 13 15 13 16 15 0 16 13 11 1 9 1 15 9 2
11 15 4 13 0 14 13 9 1 10 9 2
2 11 11
9 11 11 2 8 2 1 12 12 9
18 15 13 15 9 2 7 13 15 3 3 2 1 10 11 9 0 11 2
29 15 13 0 9 1 10 0 9 1 10 9 7 9 1 9 7 9 9 9 2 3 1 10 9 7 9 9 9 2
16 15 4 13 1 10 9 10 4 13 15 9 9 7 0 9 2
16 13 1 1 10 0 9 1 10 9 9 9 4 13 10 9 2
10 6 13 16 15 4 13 1 15 9 2
17 15 9 1 10 9 13 16 15 13 0 1 10 9 15 13 1 2
33 3 2 6 13 15 13 2 1 9 2 10 9 7 9 9 1 0 9 1 11 15 4 13 16 13 9 1 15 9 1 15 9 2
13 13 4 15 9 7 10 9 13 0 7 9 9 2
6 9 13 0 1 9 2
16 15 4 13 15 1 10 9 1 9 14 13 1 1 10 9 2
6 13 15 1 15 9 2
17 11 11 12 11 11 8 11 2 11 12 2 12 2 12 9 7 9
5 2 8 8 8 9
7 2 8 8 8 8 8 9
11 0 15 13 15 4 14 13 15 3 3 2
6 15 13 0 1 15 2
2 6 2
8 13 11 11 14 13 10 9 2
3 8 8 8
3 12 12 9
2 11 2
16 15 4 4 13 15 9 1 9 1 11 1 11 1 10 9 2
19 15 4 13 1 10 9 1 9 13 9 1 10 0 9 3 1 11 9 2
16 13 16 15 4 13 1 11 2 13 1 15 9 1 0 9 2
1 11
2 8 8
3 12 12 9
11 15 13 10 9 9 15 13 14 13 1 2
3 8 8 8
3 12 12 9
2 11 2
21 15 4 13 1 11 1 11 9 7 4 13 14 13 1 15 1 0 9 16 0 2
11 6 13 15 13 10 9 4 13 1 15 2
2 9 2
2 11 11
10 15 13 10 9 13 1 12 1 15 2
8 6 13 10 9 1 11 11 2
5 8 1 12 12 9
4 0 11 11 2
22 15 4 3 4 13 0 1 10 9 9 9 9 9 12 10 4 13 0 1 15 9 2
33 15 4 3 13 1 10 9 9 2 9 9 2 1 11 7 4 13 14 13 15 0 9 7 9 14 13 15 9 1 10 9 9 2
18 15 4 13 3 16 15 4 13 15 10 9 7 9 1 9 9 9 2
13 9 15 4 13 14 13 13 15 9 4 4 13 2
2 3 2
4 11 11 12 8
13 15 4 13 10 0 9 1 15 9 1 10 9 2
5 8 1 12 12 9
4 0 11 11 2
22 15 4 3 4 13 0 1 10 9 9 9 9 9 12 10 4 13 0 1 15 9 2
33 15 4 3 13 1 10 9 9 2 9 9 2 1 11 7 4 13 14 13 15 0 9 7 9 14 13 15 9 1 10 9 9 2
18 15 4 13 3 16 15 4 13 15 10 9 7 9 1 9 9 9 2
13 9 15 4 13 14 13 13 15 9 4 4 13 2
2 3 2
4 11 11 12 8
6 15 13 0 1 15 2
7 11 13 1 10 0 9 2
3 8 8 8
3 12 12 9
3 0 9 2
23 15 4 13 14 13 10 9 1 11 11 0 1 10 0 0 9 9 1 11 12 2 12 2
11 6 13 15 9 7 9 3 3 16 0 2
11 15 4 13 13 10 9 9 7 15 9 2
2 9 2
5 11 11 7 11 11
27 15 13 14 13 15 16 15 13 0 2 1 15 9 7 0 9 2 11 14 12 2 12 2 11 11 9 2
15 10 9 13 1 9 12 2 9 9 2 9 12 5 12 2
6 15 9 4 13 3 2
14 6 13 15 13 16 15 13 0 1 10 1 10 9 2
14 15 4 4 13 1 10 9 9 3 2 3 0 9 2
14 9 9 9 2 11 2 11 12 1 12 9 1 11 11
14 9 9 9 2 11 2 11 12 1 12 9 1 11 11
14 9 12 2 11 2 11 12 1 12 9 1 11 11 11
14 9 12 2 11 2 11 12 1 12 9 1 11 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
14 9 12 2 11 2 11 12 1 12 9 1 11 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
13 9 12 2 11 2 11 12 1 12 9 1 11 11
16 6 13 16 9 7 9 13 0 1 9 2 6 13 0 9 2
2 9 2
2 11 12
8 13 15 1 10 9 13 0 2
8 15 4 13 15 10 9 9 2
2 9 2
5 8 1 12 12 9
6 3 0 1 15 9 2
33 13 15 10 0 3 14 13 7 13 11 14 0 9 16 15 4 13 2 15 13 10 9 13 1 3 2 16 15 4 13 3 2 2
11 15 13 14 13 15 3 1 15 3 9 2
22 16 11 13 10 9 3 2 15 13 15 4 3 13 15 1 15 9 16 15 13 3 2
1 11
3 0 9 2
5 9 7 0 9 2
4 6 2 11 2
6 11 4 13 1 9 2
1 11
2 8 8
3 12 12 9
4 0 9 0 9
6 9 2 11 2 11 9
7 9 2 12 9 2 11 2
5 9 2 0 9 9
12 9 2 9 4 4 13 1 0 9 1 9 2
9 9 9 2 11 9 4 4 13 2
23 6 13 11 11 2 12 2 7 11 11 2 12 2 1 10 0 13 2 1 9 7 9 2
17 6 13 3 16 7 3 15 13 14 13 10 9 7 1 10 9 2
8 6 2 15 4 13 1 9 5
5 1 9 9 1 5
4 1 9 9 5
7 6 2 15 4 14 13 5
1 2
17 6 13 10 9 1 15 1 15 9 1 12 9 2 11 2 11 9
3 13 15 2
3 11 11 2
6 13 15 1 10 9 2
15 3 11 7 15 4 14 13 0 14 13 1 1 0 9 2
2 11 2
6 6 13 10 9 3 2
21 1 9 2 11 4 13 10 0 9 9 1 10 9 13 10 9 16 15 13 3 2
23 3 10 9 4 13 1 1 10 11 9 15 13 10 9 1 10 9 7 13 10 9 9 2
24 11 2 6 13 2 11 11 3 13 10 9 14 13 9 1 10 9 7 9 1 15 0 9 2
16 13 15 13 16 15 13 10 0 9 10 15 4 13 14 13 2
2 9 2
1 11
4 11 7 11 2
5 1 2 11 11 11
23 15 13 15 9 1 10 11 9 16 10 9 4 13 10 0 13 9 1 9 1 10 9 2
48 11 2 15 15 9 13 14 13 15 9 9 3 7 13 15 14 13 15 14 13 9 1 2 11 11 11 2 10 9 1 11 2 11 2 7 2 11 2 11 13 1 15 11 11 11 9 2 2
2 11 11
3 12 12 9
9 10 9 9 4 4 13 1 0 2
3 9 11 2
11 15 13 10 0 11 9 13 1 10 11 2
3 6 13 2
3 0 9 2
3 11 9 11
4 6 13 13 2
2 11 2
10 13 15 10 0 9 14 13 1 15 2
3 11 11 11
3 12 12 9
12 6 13 10 13 9 9 1 11 1 12 9 2
7 13 10 9 1 9 3 2
6 11 9 0 13 9 9
12 9 0 9 1 9 9 2 11 9 9 9 9
3 9 9 2
3 9 9 2
26 10 9 1 10 9 4 13 1 10 0 9 2 7 9 9 2 1 10 9 9 2 7 9 9 2 2
13 10 0 9 2 7 9 9 2 13 12 11 12 2
13 10 9 9 2 7 9 9 2 13 12 11 12 2
7 9 0 9 2 9 2 2
20 10 9 13 1 0 13 9 1 10 9 1 12 9 7 10 9 1 12 9 2
14 10 9 13 11 11 11 11 1 11 2 11 0 9 2
36 11 13 1 10 13 9 2 9 13 0 1 9 2 9 7 9 1 1 7 13 9 1 9 2 9 13 0 1 9 2 9 7 9 1 9 2
24 10 9 9 4 13 9 13 1 9 1 11 2 12 5 0 7 0 9 1 9 14 9 2 2
15 10 9 9 1 10 9 1 10 9 4 13 10 9 9 2
24 11 4 13 9 1 10 9 1 10 13 9 9 7 13 9 1 10 9 1 10 13 9 9 2
45 9 4 4 13 2 1 10 9 1 10 13 9 13 1 10 0 9 7 9 2 1 10 0 9 1 0 9 3 3 1 12 9 9 1 10 9 1 10 10 9 4 13 1 9 2
2 9 2
19 10 9 4 13 1 11 9 1 9 1 9 2 10 4 13 10 0 9 2
4 9 1 9 2
30 10 9 1 9 1 10 10 9 4 13 4 13 0 9 2 12 9 2 7 10 9 13 4 13 1 0 9 1 9 2
4 9 1 9 2
4 13 10 9 9
2 13 9
3 13 9 9
6 13 11 9 2 9 2
6 13 1 0 9 2 9
10 13 10 11 11 9 9 2 9 2 9
9 13 11 2 15 13 10 11 9 2
6 13 1 11 9 2 9
8 13 1 10 2 5 2 1 11
9 13 1 10 2 5 2 1 9 9
18 13 1 10 2 5 2 1 2 13 9 2 2 7 2 3 13 2 2
10 13 10 9 13 9 16 13 1 9 3
15 0 2 9 2 13 1 2 9 2 14 13 9 9 2 9
10 14 13 2 0 9 13 1 2 9 2
7 9 11 2 13 15 9 2
3 11 11 11
3 12 12 9
22 15 13 11 16 15 13 10 9 1 0 9 14 13 2 2 10 9 1 11 11 2 2
21 15 4 13 1 10 0 9 14 13 10 9 13 9 7 9 9 9 1 0 9 2
1 11
2 11 2
23 16 11 14 9 3 1 10 9 9 13 0 2 15 13 1 15 16 9 13 14 4 13 2
19 10 9 13 1 10 9 16 10 9 9 13 10 9 14 9 1 0 9 2
21 16 9 1 9 13 14 0 9 15 4 14 13 10 9 14 13 1 15 0 9 2
28 16 10 0 0 9 13 14 1 0 9 2 10 9 13 3 1 10 0 0 9 1 15 3 13 10 9 15 2
18 15 13 10 9 1 11 14 9 13 10 0 9 1 9 1 10 9 2
40 15 9 13 16 0 9 13 10 0 9 10 10 9 4 13 1 10 11 9 9 2 15 9 13 16 10 11 9 13 0 9 1 10 9 16 15 4 3 13 2
32 1 10 0 9 16 10 9 4 3 14 13 14 13 1 11 3 10 9 16 13 3 15 9 15 13 3 0 7 4 3 13 2
30 15 4 13 15 16 15 4 13 10 9 13 9 7 2 16 15 13 10 9 16 13 10 9 9 2 6 13 15 13 2
1 11
2 11 11
3 12 12 9
2 11 11
3 12 12 9
2 3 2
20 11 11 11 4 13 1 3 1 10 0 9 9 1 10 9 1 11 2 11 2
33 11 11 11 13 10 0 9 1 10 9 7 13 1 1 0 1 9 1 10 9 2 1 2 0 9 1 11 2 11 1 9 9 2
26 3 2 10 0 9 9 2 11 11 2 4 13 0 9 9 9 1 10 9 1 9 14 13 10 9 2
3 0 9 2
12 11 9 2 9 2 11 11 11 5 0 9 9
13 10 9 16 13 10 0 0 9 1 10 9 9 2
2 6 2
20 6 2 9 13 10 9 14 13 10 9 1 10 9 7 9 1 15 0 9 2
23 9 9 13 14 13 9 9 10 13 7 10 9 2 9 9 7 9 9 2 3 10 3 2
15 2 16 2 15 4 13 10 9 1 0 1 10 9 2 2
9 15 13 10 9 16 13 10 9 2
3 0 9 2
1 11
2 11 2
6 6 13 10 9 3 2
21 1 9 2 11 4 13 10 0 9 9 1 10 9 13 10 9 16 15 13 3 2
23 3 10 9 4 13 1 1 10 11 9 15 13 10 9 1 10 9 7 13 10 9 9 2
24 11 2 6 13 2 0 9 3 13 10 9 14 13 9 1 10 9 7 9 1 15 0 9 2
16 13 15 13 16 15 13 10 0 9 10 15 4 13 14 13 2
2 9 2
1 11
4 11 7 11 2
5 1 2 11 11 11
23 15 13 15 9 1 10 11 9 16 10 9 4 13 10 0 13 9 1 9 1 10 9 2
48 11 2 15 15 9 13 14 13 15 9 9 3 7 13 15 14 13 15 14 13 9 1 2 11 11 11 2 10 9 1 11 2 11 2 7 2 11 2 11 13 1 15 11 11 11 9 2 2
2 11 11
3 12 12 9
9 10 9 9 4 4 13 1 0 2
3 9 11 2
11 15 13 10 0 11 9 13 1 10 11 2
3 6 13 2
3 0 9 2
3 11 9 11
4 6 13 13 2
2 11 2
9 15 4 13 1 9 1 11 9 2
11 10 9 15 4 13 3 1 9 11 9 2
1 11
14 15 4 13 10 9 2 15 13 16 11 13 10 9 2
1 11
7 4 15 13 1 15 9 2
5 15 13 1 9 2
19 15 13 10 9 1 11 11 2 3 3 2 3 14 13 0 15 4 13 2
7 15 9 13 10 9 9 2
7 4 15 13 12 9 9 2
11 16 3 2 15 4 13 14 13 7 13 2
4 9 10 9 2
9 15 4 13 15 0 9 1 11 2
2 9 2
1 11
19 11 11 11 11 11 2 0 11 12 2 12 2 12 9 2 12 2 12 9
4 15 13 15 2
8 15 13 15 13 12 11 11 2
28 3 2 11 2 11 12 2 12 12 9 5 12 9 2 11 5 12 2 11 11 2 11 7 11 2 2 11 2
4 3 2 9 9
1 5
4 12 5 12 11
6 13 2 3 9 2 12
3 9 2 12
11 3 13 10 9 1 11 11 14 9 9 2
5 15 4 15 13 2
1 11
5 11 2 6 13 2
20 6 13 15 10 9 9 16 16 15 7 11 11 13 0 16 15 15 4 13 2
8 1 15 2 15 4 15 13 2
1 11
19 1 10 9 1 11 11 15 3 6 13 1 9 15 9 1 9 1 11 2
5 6 13 13 11 9
2 0 9
2 11 11
5 6 13 10 13 2
1 11
27 6 13 11 11 9 1 15 0 0 9 9 7 10 0 9 9 2 13 11 9 2 1 7 1 9 2 2
1 11
17 15 4 13 12 10 9 2 7 15 4 13 15 3 15 13 0 2
1 11
4 9 3 3 2
10 4 15 3 13 10 9 15 4 13 2
1 11
23 2 9 2 8 8 8 8 8 8 8 9 2 2 9 2 8 8 8 8 8 8 9 2
6 3 13 10 9 9 2
10 6 13 15 13 16 15 13 9 0 2
2 9 2
4 11 11 0 9
16 15 13 3 2 7 15 4 14 13 10 10 9 7 9 0 2
11 4 15 13 10 2 6 2 9 1 15 2
8 4 15 6 13 1 10 9 2
9 15 13 16 15 10 9 13 3 2
17 15 13 9 9 2 7 9 2 0 9 2 3 1 9 9 2 2
12 15 13 15 4 13 14 13 1 12 1 15 2
16 6 13 15 13 10 9 1 9 15 4 13 3 1 10 9 2
2 9 2
2 11 2
11 1 15 9 9 2 6 13 10 9 3 2
14 15 4 13 14 13 1 15 1 10 9 1 10 9 2
2 9 2
1 11
10 11 11 9 9 9 9 7 9 9 8
11 2 9 9 2 9 2 9 0 9 2 2
3 8 8 8
3 12 12 9
6 16 15 15 4 13 2
17 1 9 7 9 2 15 13 3 1 9 9 13 13 0 9 9 2
8 15 13 3 0 1 10 9 2
9 15 13 10 13 9 1 15 9 2
33 16 11 14 9 4 13 10 9 9 9 2 9 9 2 7 10 9 9 2 4 11 1 10 9 13 10 9 3 1 10 9 9 2
8 15 4 13 0 1 10 9 2
23 1 9 2 15 13 0 3 15 13 10 0 9 9 7 15 13 14 13 1 15 9 9 2
33 15 4 14 13 0 3 3 14 13 15 9 1 3 0 9 1 11 2 3 3 10 9 13 1 0 2 9 2 9 2 9 2 2
12 15 4 13 15 9 9 3 3 1 15 9 2
22 6 13 15 13 3 15 9 4 13 10 11 9 13 0 1 10 9 1 15 9 9 2
11 6 13 7 13 1 15 9 1 10 9 2
2 9 2
1 11
2 10 2
14 10 9 16 10 9 9 9 9 4 13 9 1 3 2
14 11 2 9 11 12 9 5 12 9 2 11 12 2 2
11 10 9 15 13 0 1 9 13 16 13 2
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
3 11 11 11
2 11 11
10 9 9 4 3 4 13 1 10 0 2
20 1 9 2 15 4 13 1 10 1 15 10 9 1 10 9 1 15 0 9 2
17 1 9 15 4 4 13 15 14 13 15 9 1 9 1 15 9 2
32 15 15 4 14 13 10 9 4 3 13 9 2 10 9 1 12 2 1 10 9 13 1 9 1 15 9 1 10 0 9 9 2
13 16 9 13 10 9 1 10 0 6 13 15 13 2
3 0 9 2
3 11 2 9
10 11 2 15 13 1 11 9 1 15 2
5 13 15 13 9 2
2 9 2
1 11
10 15 13 10 9 1 15 9 1 11 2
14 15 13 10 9 1 10 9 15 4 13 1 15 9 2
7 9 16 13 1 1 15 2
1 11
2 11 2
11 15 4 14 13 3 1 11 7 11 11 2
13 4 15 6 13 11 14 13 10 9 1 11 9 2
22 11 2 11 7 15 13 10 0 9 9 7 15 13 3 0 16 15 4 13 10 9 2
35 15 13 9 1 10 9 7 11 13 1 1 9 7 15 4 13 14 13 0 16 15 13 1 1 15 7 10 9 2 0 9 10 4 13 2
2 13 15
1 11
13 13 15 13 3 15 4 13 3 2 9 2 8 2
2 9 2
1 11
3 6 15 2
15 15 13 14 13 15 13 1 15 16 15 13 1 15 9 2
9 13 15 13 16 15 13 10 9 2
2 9 2
1 11
40 11 11 13 16 15 13 15 1 10 9 14 13 9 1 2 11 14 0 9 9 7 9 2 3 3 1 0 9 1 9 2 9 2 9 2 0 9 2 9 2
26 11 11 4 13 14 13 1 11 11 11 2 11 2 1 10 12 2 9 9 9 13 2 11 11 2 2
34 11 4 13 11 7 10 9 1 0 9 1 10 0 12 9 14 13 3 15 13 1 9 9 7 14 13 3 15 13 1 10 9 9 2
14 6 13 15 13 1 15 0 9 16 15 4 13 15 2
2 9 2
1 11
7 6 13 10 10 1 15 2
2 9 2
1 11
2 11 2
3 13 15 2
2 11 11
7 3 1 2 11 9 9 2
1 11
2 11 2
5 12 1 12 9 2
20 15 13 16 10 9 9 4 3 13 14 13 10 11 11 2 11 9 3 3 2
23 15 9 9 13 14 13 10 9 7 9 1 10 9 4 15 13 1 10 9 1 10 9 2
24 1 10 9 2 15 13 14 13 1 11 11 7 11 14 13 7 13 10 9 1 10 9 9 2
19 15 13 10 0 9 13 10 9 1 15 2 15 2 11 11 7 11 11 2
19 7 3 10 9 1 10 9 7 10 9 1 10 9 14 13 1 10 9 2
16 11 2 6 13 10 9 1 11 2 11 2 11 11 7 15 2
2 9 2
2 11 2
46 15 4 4 13 1 15 9 9 2 11 11 11 16 16 15 4 13 10 11 1 11 11 11 11 7 11 11 13 15 9 9 15 13 16 10 9 4 13 1 9 9 14 13 15 9 2
11 3 10 9 13 15 16 10 9 4 13 2
18 15 4 13 16 10 9 4 13 10 9 9 1 10 11 11 9 9 2
13 15 4 13 0 0 9 14 13 15 1 10 9 2
20 11 11 2 15 13 16 11 11 11 14 9 9 1 11 13 11 12 2 12 2
13 6 13 1 1 15 15 9 13 7 15 9 9 2
2 9 2
37 11 11 11 9 9 11 11 11 11 2 11 2 12 11 11 11 11 11 2 11 12 11 9 2 12 9 2 12 9 2 12 9 2 2 8 2 8
2 8 8
3 12 12 9
8 11 2 9 13 3 14 0 2
10 13 15 1 10 9 1 10 9 9 2
10 15 4 13 7 11 7 15 14 13 2
8 15 13 15 4 13 3 11 2
6 4 15 13 15 3 2
1 9
1 11
16 2 4 15 13 15 14 13 3 1 10 11 9 1 15 9 2
1 4
2 8 8
3 12 12 9
15 4 15 13 15 4 4 13 9 2 3 1 10 12 9 2
35 15 13 10 9 9 10 9 1 12 9 2 11 9 2 1 11 11 11 11 11 1 10 11 9 13 0 9 1 0 9 16 13 1 11 2
14 13 4 10 9 1 9 7 10 0 11 9 13 9 2
17 16 15 4 13 14 13 1 9 7 1 9 2 6 13 15 13 2
20 15 4 13 1 11 11 1 11 12 5 12 7 11 11 1 11 12 5 12 2
12 1 11 2 15 4 4 13 3 1 11 9 2
11 1 11 2 15 4 4 13 1 11 9 2
13 13 15 13 16 15 4 13 14 13 1 10 9 2
1 11
5 6 13 14 13 2
2 9 2
1 11
2 11 11
3 12 12 9
24 3 1 11 2 11 12 2 1 12 9 2 11 9 2 10 13 12 9 2 11 11 2 9 2
3 6 13 2
1 11
1 5
1 9
7 9 2 10 9 13 0 2
34 16 15 4 13 15 1 9 6 13 15 13 1 9 7 3 13 15 1 15 9 2 15 4 14 13 10 9 7 13 15 9 1 9 2
3 13 15 2
2 2 9
5 10 9 4 13 2
12 15 4 13 14 13 1 10 0 9 11 9 2
1 11
2 8 8
3 12 12 9
2 6 2
16 16 9 13 3 15 13 3 0 14 13 15 4 13 15 13 2
2 9 2
2 8 8
3 12 12 9
22 10 9 4 4 13 1 12 9 2 11 9 2 10 13 12 9 2 11 11 9 2 2
15 6 13 15 13 16 15 4 13 16 15 14 13 15 3 2
1 11
10 10 9 15 13 4 4 13 1 11 2
12 16 15 4 13 15 13 2 6 13 15 13 2
1 11
3 8 8 8
3 12 12 9
2 11 2
3 13 0 2
1 11
2 8 8
3 12 12 9
10 11 2 6 13 16 10 13 9 13 2
5 15 9 13 12 2
1 11
23 1 10 9 1 15 9 1 10 9 9 9 2 4 9 13 10 0 9 13 10 9 9 2
18 16 15 13 10 0 0 9 4 4 13 2 6 13 0 14 13 15 2
2 9 2
1 11
13 15 13 15 9 3 10 9 7 4 13 10 9 2
26 4 15 13 10 9 9 1 12 9 2 11 2 10 13 12 9 2 11 11 2 1 11 2 11 12 2
3 6 13 2
1 11
26 10 9 9 4 4 13 1 11 2 11 12 1 12 9 2 11 2 10 13 12 9 2 11 11 2 2
6 15 4 13 10 9 2
18 16 9 4 13 14 4 13 3 7 13 1 9 2 6 13 15 13 2
2 9 2
1 11
12 15 4 13 1 15 9 13 1 0 9 9 2
7 15 13 10 0 9 9 2
17 15 4 3 13 1 9 1 11 10 4 13 7 0 7 0 9 2
17 0 2 9 2 13 1 0 9 1 10 0 9 1 11 7 11 2
6 15 4 13 1 11 2
13 15 13 14 3 0 1 16 15 15 4 13 1 2
31 3 10 0 9 13 9 10 4 14 13 1 10 11 2 16 11 13 3 3 0 16 15 4 13 1 10 0 9 9 2 2
16 12 9 10 4 14 13 1 1 10 9 13 10 9 9 9 2
9 13 15 13 3 15 4 13 3 2
1 11
2 11 11
3 12 12 9
14 3 15 13 2 15 13 15 12 2 0 7 13 15 2
9 11 4 13 15 10 0 9 9 2
4 9 9 3 2
3 13 3 2
13 15 13 16 10 12 2 9 9 9 13 10 9 2
6 15 4 13 15 3 2
29 11 11 1 11 13 15 0 9 14 13 15 4 3 13 10 9 9 9 16 10 13 9 13 1 7 13 1 9 2
13 15 13 15 1 15 7 4 13 10 0 13 3 2
10 13 15 4 13 9 14 13 15 9 2
11 9 4 3 13 1 10 9 7 9 9 2
14 15 4 14 13 9 1 15 1 9 13 10 13 9 2
59 11 13 16 15 13 10 13 9 9 10 4 4 13 2 15 13 15 13 15 13 14 13 10 9 9 1 12 9 3 1 12 2 7 10 0 9 9 2 13 10 12 9 9 14 13 10 9 1 10 0 9 16 10 0 13 14 13 2 2
42 15 13 15 13 1 10 9 3 2 7 11 14 9 13 14 13 9 13 1 9 3 16 0 9 4 4 13 1 9 2 3 16 15 13 10 9 13 10 9 7 9 2
2 9 2
14 13 16 15 13 9 7 16 15 4 13 1 10 9 2
15 15 13 10 0 9 15 4 13 9 0 14 13 10 9 2
4 1 0 9 2
1 11
3 6 3 2
6 7 0 11 11 3 2
9 1 15 4 15 13 10 0 9 2
19 15 13 0 1 11 2 3 13 1 1 11 7 11 2 13 3 2 8 2
7 3 4 15 13 10 9 2
4 11 2 11 2
2 11 2
2 11 2
3 11 11 2
4 11 11 11 2
6 15 4 3 13 9 2
54 1 1 15 2 6 2 15 13 10 0 9 2 13 10 0 9 1 11 11 2 13 10 0 9 2 15 13 14 13 10 0 9 3 2 10 12 2 9 0 11 11 13 13 15 10 9 2 2 15 13 2 10 0 2
11 4 15 13 9 1 7 1 10 0 9 2
5 4 15 13 0 2
6 1 10 0 9 9 2
5 3 13 15 9 2
7 13 14 13 3 1 9 2
14 10 9 15 13 1 1 11 11 7 11 11 1 9 2
1 11
5 8 1 12 12 9
2 11 2
6 0 11 11 2 9 2
5 13 10 13 0 2
5 4 15 13 15 2
1 11
20 11 11 13 15 16 15 13 10 9 9 2 0 7 0 2 1 10 11 9 2
25 15 4 13 14 13 0 9 1 10 11 11 9 2 3 11 2 7 13 15 9 4 13 3 0 2
7 4 15 13 15 10 9 2
17 15 4 13 1 11 11 1 11 7 15 4 13 1 10 9 9 2
6 13 15 1 15 9 2
2 9 2
1 11
70 2 16 2 2 2 8 2 0 9 0 1 9 9 1 15 0 9 13 10 9 7 10 0 9 1 2 10 9 14 4 13 1 9 9 2 2 13 7 14 13 1 10 0 9 9 2 9 7 10 9 9 2 4 4 3 13 7 13 7 10 2 9 2 4 4 13 1 0 9 2
1 3
2 11 11
3 12 12 9
19 11 2 3 13 10 9 9 15 13 1 11 11 2 11 11 7 11 11 2
9 15 13 15 13 7 9 7 9 2
10 15 13 1 10 9 9 7 9 0 2
21 16 10 9 13 14 4 13 1 11 2 15 4 13 15 1 11 2 11 7 11 2
1 9
2 11 11
3 12 12 9
20 11 11 13 15 16 15 13 10 9 9 2 0 7 0 2 1 10 11 9 2
25 15 4 13 14 13 0 9 1 10 11 11 9 2 3 11 2 7 13 15 9 4 13 3 0 2
7 4 15 13 15 10 9 2
17 15 4 13 1 11 11 1 11 7 15 4 13 1 10 9 9 2
6 13 15 1 15 9 2
2 9 2
1 11
24 6 13 10 13 9 14 13 16 15 4 13 10 1 10 9 10 15 13 0 16 13 1 11 2
14 15 4 13 1 11 11 1 11 2 11 12 2 12 2
3 13 15 2
1 11
4 11 2 8 2
3 12 12 9
19 9 2 13 4 10 13 9 10 13 0 9 1 10 9 1 12 7 12 2
15 10 9 4 3 4 13 1 10 9 9 3 3 16 0 2
19 13 15 1 15 9 7 15 13 15 4 13 10 0 9 14 13 10 9 2
6 2 11 11 0 9 9
3 2 5 2
14 13 16 10 9 13 0 2 13 1 11 14 9 9 2
11 2 11 2 11 2 11 2 2 2 8 2
3 12 12 9
7 0 9 9 1 11 9 12
6 9 9 12 9 9 2
14 13 4 11 14 9 9 12 2 9 12 2 9 9 2
17 15 13 15 13 0 1 10 9 7 9 15 4 13 1 10 9 2
25 1 10 9 2 10 9 2 2 13 10 0 9 9 9 1 9 9 1 10 9 12 1 12 2 2
19 2 13 9 9 9 9 1 12 0 1 0 9 1 9 1 9 9 2 2
12 2 13 1 13 9 9 9 1 9 9 2 2
40 2 13 10 12 9 5 0 9 1 0 9 16 13 9 9 1 0 9 2 13 10 9 16 10 9 14 13 14 13 0 9 9 7 0 11 2 13 9 2 2
40 2 13 9 14 13 9 7 13 13 9 1 9 9 9 2 7 13 10 9 9 13 14 13 10 9 1 10 9 1 10 9 12 9 2 12 5 12 2 2 2
26 2 13 10 0 9 1 9 9 2 1 10 12 5 9 14 13 7 9 7 10 9 1 13 9 9 2
27 10 13 9 4 13 0 3 1 0 9 1 10 9 1 9 7 13 9 1 1 0 9 7 0 9 2 2
21 2 13 10 9 9 1 10 9 7 9 9 2 16 3 0 1 10 0 9 2 2
28 2 13 10 12 2 9 0 9 1 9 9 9 13 1 12 2 16 9 9 13 10 0 9 1 0 9 2 2
10 2 13 10 9 9 9 1 10 9 2
51 11 3 13 16 10 9 9 9 9 2 9 2 4 13 0 1 9 14 9 2 7 4 13 10 3 0 9 9 13 14 13 13 9 1 9 9 7 14 13 10 12 2 9 1 12 2 9 0 9 9 2
39 15 3 4 13 1 10 9 16 10 10 2 9 9 4 13 1 11 14 9 1 11 11 1 11 12 7 12 2 14 13 10 9 7 14 13 1 15 9 2
12 15 13 3 16 13 15 9 7 13 15 9 2
31 10 13 9 13 10 9 12 9 9 2 10 9 2 10 9 1 11 14 13 9 9 12 2 2 7 10 9 1 13 9 2
19 3 2 6 13 16 10 9 9 7 10 9 13 1 2 11 12 2 9 2
22 15 4 13 0 14 13 10 0 9 1 10 0 9 1 11 2 1 9 1 0 9 2
12 15 13 3 16 13 15 1 11 12 5 12 2
17 1 10 9 2 15 13 15 0 9 1 10 0 7 0 9 9 2
12 11 11 11 11 2 12 2 12 2 12 2 12
26 2 8 8 8 8 8 8 9 2 2 8 8 8 9 2 2 8 8 8 8 8 8 8 8 9 2
4 9 11 11 2
36 15 13 14 13 16 10 9 1 11 11 4 13 14 13 10 9 1 10 9 1 9 9 9 9 1 10 9 14 9 13 1 11 9 7 9 2
3 13 15 2
2 3 2
6 11 11 9 2 11 11
14 13 4 10 9 1 10 9 9 1 10 9 14 9 2
3 0 9 2
13 15 9 13 3 14 4 13 1 12 5 12 9 2
15 11 11 2 15 0 9 2 4 13 10 9 1 15 9 2
23 11 11 4 13 1 10 0 9 1 15 9 7 15 4 13 15 3 1 9 9 3 9 2
25 9 4 4 13 1 15 1 9 2 9 2 12 2 2 9 2 12 2 2 7 9 2 12 2 2
17 15 4 13 10 9 9 1 9 14 0 9 2 12 9 11 2 2
7 10 13 1 9 13 12 2
4 9 13 12 2
13 10 9 14 9 13 9 1 12 9 2 11 2 2
2 11 11
5 13 1 2 11 11
3 12 12 9
14 13 4 10 9 1 10 9 9 1 10 9 14 9 2
3 0 9 2
13 15 9 13 3 14 4 13 1 12 5 12 9 2
15 11 11 2 15 0 9 2 4 13 10 9 1 15 9 2
23 11 11 4 13 1 10 0 9 1 15 9 7 15 4 13 15 3 1 9 9 3 9 2
25 9 4 4 13 1 15 1 9 2 9 2 12 2 2 9 2 12 2 2 7 9 2 12 2 2
17 15 4 13 10 9 9 1 9 14 0 9 2 12 9 11 2 2
7 10 13 1 9 13 12 2
4 9 13 12 2
13 10 9 14 9 13 9 1 12 9 2 11 2 2
3 0 9 2
7 13 14 13 10 0 9 2
7 15 13 10 3 0 9 2
6 15 4 13 10 9 2
2 0 2
1 11
2 11 11
3 12 12 9
2 11 2
60 3 16 13 10 0 9 9 2 12 7 12 5 2 15 13 15 4 13 16 10 2 0 2 9 4 13 0 7 4 1 9 13 0 2 7 16 10 0 9 1 9 4 13 0 7 0 1 3 13 1 9 7 9 2 7 3 13 1 9 2
20 1 0 2 15 4 14 13 3 0 1 10 9 7 15 13 15 13 1 15 2
11 3 2 15 13 15 4 13 10 9 3 2
18 15 13 1 10 9 16 13 10 9 14 13 15 1 10 0 0 9 2
38 7 16 10 2 3 0 2 9 13 3 0 1 15 9 1 10 9 1 11 7 11 2 15 13 14 13 3 10 9 1 9 1 10 9 2 9 3 2
15 9 2 10 9 14 13 9 1 2 9 9 2 4 13 2
13 10 9 13 9 0 16 13 10 2 9 9 2 2
22 10 9 9 13 0 0 9 1 11 7 15 7 15 9 13 7 13 10 0 9 3 2
14 15 9 9 13 10 9 13 10 9 1 2 9 2 2
29 1 15 9 2 11 11 13 11 7 11 14 13 15 1 10 9 1 10 9 15 13 14 13 15 9 3 1 9 2
8 7 11 11 14 9 13 0 2
25 1 10 11 9 2 10 0 11 2 11 2 7 10 0 11 2 11 2 13 9 16 13 1 9 2
9 11 13 10 2 9 2 9 9 2
25 10 9 3 13 1 11 14 13 10 2 0 2 9 2 1 9 2 9 2 9 9 2 10 9 2
21 1 10 0 9 2 10 11 9 13 11 2 15 9 2 7 15 9 1 10 9 2
25 11 13 3 3 16 10 9 1 11 14 9 9 13 15 0 14 13 1 10 0 9 1 10 9 2
26 15 3 13 16 3 9 4 3 13 1 15 0 9 2 9 2 13 1 10 13 9 13 1 10 9 2
16 9 2 15 13 0 16 11 14 13 3 15 9 16 4 13 2
14 1 10 0 9 2 10 9 1 10 2 9 2 13 2
23 1 10 9 2 10 0 9 1 11 13 10 0 9 13 14 13 3 10 9 16 4 13 2
35 1 10 0 9 2 9 13 16 11 2 1 9 2 2 13 1 10 9 2 2 7 10 9 13 2 7 11 13 1 10 9 1 11 9 2
6 15 13 0 2 11 2
20 9 4 14 13 3 16 13 10 9 9 3 1 10 9 2 13 14 13 15 2
7 9 3 3 1 10 9 2
38 11 3 13 10 0 9 2 4 14 13 10 9 1 9 9 1 15 9 2 3 13 16 10 9 9 13 14 13 3 2 13 7 13 1 9 7 9 2
5 4 13 10 9 2
2 8 8
3 12 12 9
9 15 13 10 9 1 15 9 9 2
20 10 9 7 9 9 4 13 1 10 11 2 0 9 13 9 9 9 0 9 2
19 1 1 9 9 2 3 13 9 1 10 11 9 4 13 14 13 15 9 2
20 3 2 15 13 12 9 1 11 2 11 9 7 12 9 1 11 2 11 9 2
8 6 13 15 13 1 15 9 2
7 9 9 4 13 16 13 2
5 9 2 11 1 11
10 9 2 11 2 11 9 11 2 11 9
6 9 12 9 9 12 9
7 3 2 1 9 11 1 11
8 9 2 12 5 12 12 5 12
6 9 2 11 11 2 13
4 11 11 2 13
4 11 11 2 13
4 11 11 2 13
26 1 10 9 16 15 13 9 9 7 4 14 13 2 10 9 1 10 9 7 9 9 4 4 3 13 2
21 1 3 2 13 15 1 15 9 7 6 13 15 1 9 12 16 15 13 10 9 2
4 11 11 9 9
5 0 1 15 3 2
6 15 4 14 13 9 2
1 0
1 11
8 2 11 11 11 2 2 8 2
3 12 12 9
10 6 4 14 13 15 11 9 1 9 2
4 13 1 9 2
1 11
5 9 1 10 9 2
6 4 15 13 10 9 2
2 11 11
3 12 12 9
1 3
31 11 11 2 11 11 7 11 11 1 11 4 13 1 9 1 10 11 0 1 0 9 0 11 2 11 9 7 9 9 9 2
27 10 9 9 4 3 13 14 13 11 13 0 9 9 9 7 9 0 9 9 14 13 10 9 9 9 9 2
25 3 16 15 13 1 11 14 0 9 9 15 4 13 0 9 1 9 9 9 3 1 0 9 9 2
35 15 4 3 13 1 10 9 2 0 12 2 1 10 11 9 10 13 11 2 9 2 2 11 7 11 1 11 11 11 9 12 7 9 12 2
29 10 0 9 9 13 9 1 12 5 12 12 9 1 0 9 7 15 13 0 9 14 13 12 9 13 1 9 12 2
22 9 4 13 14 13 10 11 9 9 1 12 5 12 9 9 7 12 5 12 5 9 2
22 9 13 14 13 10 0 9 1 11 14 11 11 9 12 9 7 3 13 10 9 3 2
12 11 4 13 1 3 11 9 12 13 1 3 2
24 11 14 9 4 13 14 13 16 15 13 10 9 16 13 10 9 1 7 10 13 7 13 9 2
14 10 9 4 4 13 1 10 11 14 9 7 10 11 2
37 15 13 3 3 0 14 13 11 14 13 1 10 0 7 0 9 2 7 11 13 14 13 15 0 7 2 7 0 9 1 11 3 10 9 13 0 2
23 10 9 13 14 13 11 9 1 15 12 9 11 2 11 9 1 9 1 10 0 9 9 2
23 4 9 1 15 9 6 13 15 10 0 8 13 0 9 1 10 9 1 9 1 11 12 2
2 6 13
2 8 8
3 12 12 9
12 6 13 2 7 15 4 13 1 9 3 3 2
11 15 3 3 13 9 3 9 4 13 1 2
1 11
2 11 11
3 12 12 9
36 13 1 1 15 9 9 2 1 10 9 1 9 2 15 4 14 13 15 13 0 14 13 10 10 9 1 15 9 14 9 14 13 1 10 9 2
25 15 13 0 9 9 7 13 10 9 4 13 15 14 13 9 16 0 9 4 14 13 0 0 9 2
41 10 0 9 15 13 10 9 13 1 10 9 3 10 9 13 10 9 9 1 10 0 2 0 9 2 13 5 12 12 2 7 3 13 16 15 13 14 10 0 9 2
9 1 15 9 2 15 4 3 13 2
16 15 4 13 10 9 1 9 7 15 0 9 4 13 1 9 2
10 3 15 4 14 13 14 13 10 9 2
18 3 16 15 13 2 15 9 4 13 1 10 9 2 3 10 0 9 2
21 10 9 16 13 9 13 3 0 1 10 9 1 10 9 13 14 13 15 9 1 2
9 13 1 10 12 9 9 1 15 2
17 13 15 0 14 13 10 0 9 7 15 9 1 10 0 0 9 2
23 16 13 3 1 10 0 9 3 15 4 13 10 9 16 10 9 9 13 3 12 2 9 2
2 6 13
1 8
3 12 12 9
4 0 11 11 2
9 13 15 3 3 1 15 0 9 2
5 13 4 15 9 2
9 15 13 10 0 9 1 10 9 2
20 10 9 13 1 10 9 9 9 9 2 0 2 9 7 9 2 11 11 11 2
26 15 4 13 1 11 12 2 7 10 0 9 9 13 16 16 15 13 3 1 10 9 2 15 13 0 2
9 13 3 16 13 15 9 2 9 2
2 9 2
1 11
2 2 9
2 6 2
10 10 9 14 9 13 1 10 0 9 2
11 15 13 14 0 3 15 4 4 13 15 2
5 3 4 9 13 2
6 10 9 1 10 9 2
2 8 8
3 12 12 9
3 15 13 2
41 3 13 10 9 2 16 15 4 13 1 10 9 9 2 12 9 2 14 13 1 9 2 10 9 13 15 7 13 16 15 4 13 0 15 9 13 1 10 0 9 2
12 10 9 4 13 3 1 9 7 4 14 13 2
24 15 4 14 13 6 2 3 11 2 10 0 9 2 12 9 0 2 7 15 13 1 10 9 2
14 15 13 3 2 12 7 15 13 10 9 1 15 9 2
12 1 9 1 9 2 15 13 9 1 12 9 2
7 10 15 3 13 15 13 2
13 15 13 16 11 4 3 13 14 13 1 15 0 2
17 15 13 15 16 15 13 10 9 10 4 13 14 13 1 15 9 2
10 15 13 15 9 7 13 9 1 15 2
5 3 0 2 6 2
22 10 9 10 13 1 11 13 7 15 3 13 3 1 15 2 7 15 4 14 13 15 2
21 3 2 15 13 10 0 9 16 15 4 13 14 13 15 1 9 2 12 9 2 2
9 15 13 3 12 9 0 1 9 2
9 15 13 1 10 9 1 10 9 2
15 1 9 15 13 3 1 9 9 7 1 9 15 9 13 2
11 15 13 10 9 9 3 14 13 15 1 2
11 15 13 15 9 1 10 9 1 10 9 2
16 7 15 13 0 3 11 13 14 13 15 13 15 13 3 0 2
12 6 13 10 9 1 10 11 9 9 3 3 2
2 9 2
1 11
2 11 11
3 12 12 9
10 3 2 11 4 13 1 10 9 9 2
9 15 13 1 15 0 1 15 9 2
10 13 15 9 0 1 11 10 4 13 2
5 6 13 15 13 2
2 9 2
9 11 2 6 13 9 1 15 1 11
2 11 11
3 12 12 9
2 10 2
18 10 9 7 9 9 13 15 13 0 9 9 10 13 14 4 13 3 2
38 16 15 13 0 0 9 13 11 10 9 2 0 11 2 7 3 2 11 2 15 13 15 0 14 13 10 1 10 0 9 1 10 1 2 9 9 9 2
20 15 4 13 10 9 1 11 2 11 12 7 4 13 3 12 9 14 4 13 2
18 15 4 13 16 15 13 10 9 1 10 0 9 2 9 7 3 2 2
18 15 4 13 0 9 9 1 10 9 7 10 0 9 9 1 10 9 2
29 15 13 16 9 14 13 7 1 10 9 2 12 9 5 12 9 2 7 9 2 12 9 5 12 9 2 0 9 2
16 6 13 15 9 13 10 9 3 7 13 15 9 1 10 9 2
29 1 9 2 15 4 13 10 9 10 13 0 9 14 13 16 13 12 7 0 1 10 9 4 15 4 13 10 9 2
7 9 1 9 1 15 9 2
3 13 15 2
1 11
14 3 13 15 12 5 2 10 12 12 9 2 13 1 2
8 4 15 13 15 1 0 9 2
5 0 9 2 9 2
2 11 11
3 12 12 9
4 0 9 9 2
25 10 9 13 16 11 3 13 10 0 9 1 9 9 10 4 4 13 1 0 9 7 0 9 9 2
1 11
2 8 8
2 12 12
3 3 13 9
15 0 1 11 11 11 11 2 5 12 2 5 12 5 9 2
15 0 1 11 3 5 12 2 11 12 5 9 3 5 12 2
13 11 0 9 3 13 11 14 9 9 9 13 5 12
7 14 0 1 10 0 9 2
1 11
9 11 2 6 13 9 1 15 1 11
8 11 2 10 13 13 15 9 2
18 8 2 1 9 12 2 15 4 13 10 9 1 9 1 10 0 9 2
31 8 2 1 9 12 2 1 10 0 9 1 10 9 13 2 9 2 1 10 9 2 9 2 7 1 10 9 2 9 2 2
14 8 2 1 9 12 2 13 12 9 9 1 12 9 2
14 3 2 13 10 9 1 10 9 1 9 2 12 2 2
22 8 2 1 9 12 15 4 3 13 16 10 9 9 9 15 13 13 3 10 0 9 2
25 8 2 1 9 12 2 9 2 9 2 4 4 13 14 13 1 10 9 1 10 9 1 10 9 2
17 8 2 13 10 9 2 9 2 1 10 9 1 0 0 9 9 2
16 8 2 13 10 9 1 9 16 15 4 3 13 1 9 12 2
11 8 2 3 4 10 13 9 9 9 13 2
15 8 2 1 10 9 2 10 9 9 4 3 13 1 9 2
29 3 2 1 10 0 9 1 10 9 13 10 9 2 9 2 1 10 9 2 9 2 7 1 10 9 2 9 2 2
16 8 2 1 9 9 2 13 10 9 1 9 1 10 0 9 2
9 15 4 3 13 9 2 9 9 2
23 8 2 1 9 1 9 2 9 2 9 2 13 1 10 9 9 10 15 13 14 0 13 2
17 1 9 2 9 2 2 13 10 2 9 2 2 1 10 9 9 2
15 8 2 9 4 4 13 16 15 4 3 13 1 9 12 2
16 8 2 1 9 2 9 1 9 2 13 10 9 2 9 2 2
6 15 4 13 9 9 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
2 8 8
3 12 12 9
2 11 2
28 15 4 13 14 13 10 9 10 11 4 13 1 15 0 9 9 9 10 11 4 13 1 9 1 10 0 9 2
18 13 6 13 10 9 0 9 2 1 10 9 9 9 2 1 15 9 2
8 6 13 10 13 16 15 13 2
68 8 2 10 0 9 4 14 13 10 9 13 16 15 13 9 9 2 10 1 15 0 9 13 16 15 4 13 1 9 14 9 9 7 16 15 4 13 10 9 0 0 1 9 7 10 0 1 10 9 2 7 13 0 1 15 9 2 7 13 10 9 3 1 10 9 14 9 2
42 8 2 15 4 14 13 10 2 9 2 9 1 10 9 2 3 16 10 0 9 1 10 9 2 15 4 14 2 7 4 10 9 2 13 10 9 1 9 1 10 9 2
16 16 15 13 3 16 15 13 10 9 9 2 15 4 13 3 2
45 8 2 10 9 1 9 9 13 10 9 3 1 10 0 9 2 10 9 3 13 16 10 0 9 9 13 3 0 7 3 0 2 7 15 4 13 0 9 13 15 1 10 9 2 2
52 13 1 9 10 9 1 9 2 15 13 14 13 0 9 2 13 15 9 14 13 15 9 1 1 10 9 1 9 2 9 7 9 1 10 2 9 9 9 2 1 10 9 14 13 10 9 2 13 10 9 2 2
39 3 15 4 14 13 9 1 10 9 9 1 10 9 1 10 9 1 9 16 10 0 9 13 2 3 2 3 1 10 9 16 2 13 9 2 1 9 0 2
27 13 15 13 15 9 1 10 9 7 16 15 13 0 16 15 13 15 1 0 9 16 10 9 9 4 13 2
17 16 15 13 0 2 15 4 13 10 9 1 15 0 0 9 9 2
9 9 3 1 15 9 1 10 9 2
1 11
48 9 6 13 0 14 13 11 11 7 11 11 1 15 9 2 15 4 4 13 10 9 1 15 2 9 2 2 15 4 13 1 11 1 11 1 10 9 2 7 4 13 1 1 9 1 3 12 2
8 15 4 13 1 3 1 11 2
2 11 2
19 15 4 13 1 15 10 9 1 9 2 15 13 9 9 7 10 9 9 2
18 15 4 13 1 10 9 7 4 13 15 1 15 3 1 9 7 9 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
3 11 11 11
3 12 12 9
2 11 2
22 15 9 1 9 9 4 13 3 0 16 15 13 10 1 10 9 10 13 10 9 0 2
6 13 15 0 1 15 2
9 16 3 2 13 15 0 14 13 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
1 8
3 12 12 9
2 11 2
15 15 13 16 15 4 3 13 10 9 10 13 10 0 9 2
13 3 4 15 13 1 1 10 13 9 1 10 9 2
2 11 2
23 1 9 1 15 0 9 1 10 8 9 9 9 2 15 13 15 4 13 10 0 9 9 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
4 11 7 11 2
7 4 15 13 9 1 12 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
2 11 2
26 16 15 13 1 15 9 2 11 11 1 11 11 2 9 9 2 4 13 14 13 15 9 1 15 9 2
23 15 13 0 9 1 10 9 2 8 2 9 9 2 7 4 13 14 13 1 15 1 15 2
10 15 9 13 12 7 9 9 13 8 2
14 16 15 13 1 10 9 2 15 4 13 10 9 9 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
3 11 11 11
3 12 12 9
9 3 13 9 10 13 1 12 3 2
6 11 11 11 12 12 9
8 15 13 14 13 10 0 9 2
2 9 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
3 11 11 11
3 12 12 9
22 4 15 13 12 7 3 7 4 15 13 14 13 10 1 11 16 15 4 14 4 13 2
13 3 13 15 13 7 15 4 13 15 10 0 9 2
6 11 11 11 12 12 9
2 11 2
25 4 9 9 1 10 0 9 9 13 14 4 13 7 13 10 9 10 15 13 1 15 10 0 9 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
1 8
3 12 12 9
2 11 2
24 15 13 11 11 2 15 9 9 2 7 11 11 4 3 13 10 0 0 9 1 10 9 9 2
53 15 13 1 11 11 10 9 2 15 13 3 0 1 10 9 1 10 9 1 10 9 2 7 15 13 10 0 9 2 9 9 1 9 12 0 1 10 9 1 9 1 9 1 9 10 11 4 13 1 11 3 3 2
38 3 3 16 10 9 13 2 10 0 13 9 10 15 13 0 1 2 3 16 13 10 9 2 13 16 15 4 13 13 10 9 13 10 9 1 0 9 2
13 13 16 15 4 3 13 10 9 13 3 0 9 2
2 11 11
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
3 11 11 11
3 12 12 9
10 15 4 13 9 9 12 1 15 9 2
6 15 13 11 9 12 2
3 4 13 2
2 11 2
9 9 3 3 1 15 9 1 15 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
3 11 11 11
3 12 12 9
10 15 4 13 9 11 12 1 15 9 2
6 15 13 11 9 12 2
3 4 13 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
3 11 11 11
3 12 12 9
10 15 4 13 9 9 12 1 15 9 2
6 15 13 11 9 12 2
3 4 13 2
2 11 2
9 15 4 13 10 9 1 15 9 2
6 13 15 0 14 13 2
13 15 13 1 1 10 9 9 7 4 13 3 9 2
4 6 13 15 2
2 9 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
1 8
3 12 12 9
2 11 2
15 15 9 9 4 14 13 3 10 9 9 13 14 4 13 2
20 15 3 13 1 10 0 9 9 1 10 9 9 10 13 10 9 1 9 3 2
10 13 15 10 0 9 10 15 4 13 2
2 11 2
9 15 9 1 10 9 9 13 0 2
12 1 9 1 10 9 2 15 4 13 10 9 2
9 15 9 4 14 13 10 0 9 2
4 13 15 10 2
1 11
2 6 2
14 11 11 11 11 12 12 2 9 2 12 2 9 2 8
2 10 2
9 6 13 10 13 9 9 1 11 2
17 15 13 15 10 14 13 10 9 16 15 15 13 13 10 0 9 2
12 15 13 10 3 0 2 3 0 9 1 11 2
8 11 4 13 7 13 10 9 2
29 15 4 13 16 11 4 13 10 2 9 9 2 10 13 3 15 4 13 11 1 10 9 1 1 10 0 11 9 2
20 16 9 13 10 9 7 9 1 10 9 1 10 9 2 6 13 15 10 9 2
52 3 2 15 4 13 10 9 4 14 13 0 1 10 9 9 9 9 2 7 14 13 15 2 15 4 13 9 1 9 12 10 13 15 3 16 10 11 3 13 3 14 13 16 10 9 13 0 1 10 9 9 2
15 11 11 1 10 9 9 4 13 1 15 14 13 10 9 2
9 15 13 14 13 10 9 10 9 2
11 16 15 13 10 9 2 6 13 15 13 2
15 1 9 2 15 4 13 10 0 9 1 15 1 15 9 2
2 9 2
2 11 12
10 2 9 2 8 8 8 8 8 9 2
2 11 2
36 15 4 13 16 13 10 9 9 1 15 9 2 3 2 15 13 15 4 13 14 13 3 12 9 1 9 1 11 14 13 1 11 14 9 2 2
36 16 15 13 1 15 2 16 1 10 9 15 4 14 13 11 9 2 15 4 13 14 13 1 9 9 10 4 13 14 13 10 9 1 15 9 2
9 15 1 2 9 9 13 11 12 2
41 16 15 13 16 11 12 4 13 0 1 16 13 10 9 2 9 1 10 0 9 1 1 10 9 10 13 4 13 1 15 1 1 0 11 9 2 6 13 15 13 2
29 11 4 3 13 15 16 15 4 13 13 9 2 9 1 15 9 16 15 13 13 10 1 2 9 9 1 11 12 2
4 9 2 11 2
1 11
23 4 10 9 2 15 7 11 9 2 9 2 4 13 7 3 13 10 13 3 2 9 9 2
1 9
3 11 11 12
2 10 2
9 6 13 10 13 9 9 1 11 2
17 15 13 15 10 14 13 10 9 16 15 15 13 13 10 0 9 2
12 15 13 10 3 0 2 3 0 9 1 11 2
8 11 4 13 7 13 10 9 2
29 15 4 13 16 11 4 13 10 2 9 9 2 10 13 3 15 4 13 11 1 10 9 1 1 10 0 11 9 2
20 16 9 13 10 9 7 9 1 10 9 1 10 9 2 6 13 15 10 9 2
52 3 2 15 4 13 10 9 4 14 13 0 1 10 9 9 9 9 2 7 14 13 15 2 15 4 13 9 1 9 12 10 13 15 3 16 10 11 3 13 3 14 13 16 10 9 13 0 1 10 9 9 2
15 11 11 1 10 9 9 4 13 1 15 14 13 10 9 2
9 15 13 14 13 10 9 10 9 2
11 16 15 13 10 9 2 6 13 15 13 2
15 1 9 2 15 4 13 10 0 9 1 15 1 15 9 2
2 9 2
2 11 12
10 2 9 2 8 8 8 8 8 9 2
8 13 15 3 1 10 9 3 2
33 15 4 13 11 9 10 9 16 13 11 1 11 2 11 12 1 11 2 11 7 13 1 11 2 11 12 1 11 1 11 2 11 2
8 9 9 13 5 12 1 9 2
7 11 7 11 13 1 9 2
7 4 15 7 11 13 15 2
19 11 7 11 4 14 13 0 14 13 3 1 12 1 1 11 14 0 9 2
8 6 13 15 2 13 15 13 2
2 9 2
2 11 12
16 11 2 0 1 10 0 9 2 7 15 13 15 4 13 3 2
42 15 13 1 10 9 0 9 7 15 4 13 2 15 4 14 13 16 15 13 3 7 14 2 7 15 4 13 16 15 4 4 3 13 3 1 9 10 13 0 2 9 2
2 11 2
42 10 9 9 13 10 0 11 9 9 7 9 0 1 9 2 15 13 10 9 9 13 10 9 7 11 11 13 10 0 9 7 9 16 10 9 9 9 14 13 1 9 2
20 3 0 9 4 15 13 14 13 10 11 9 16 13 10 0 11 9 9 9 2
32 15 4 13 10 9 9 1 16 13 10 9 1 10 9 9 2 15 4 3 13 1 10 0 9 10 4 13 10 9 1 9 2
9 4 15 13 15 13 14 13 0 2
4 9 2 11 11
4 6 2 9 2
4 15 13 0 2
12 15 3 4 14 13 16 15 13 15 7 11 2
4 9 2 11 2
2 11 2
29 10 0 11 9 4 13 11 10 13 9 9 1 10 9 1 10 9 9 1 9 7 10 0 9 10 13 10 9 2
8 10 0 9 9 9 13 12 2
21 15 13 1 10 9 16 11 11 4 13 15 1 10 9 2 11 4 3 13 0 2
2 11 11
16 11 2 0 1 10 0 9 2 7 15 13 15 4 13 3 2
42 15 13 1 10 9 0 9 7 15 4 13 2 15 4 14 13 16 15 13 3 7 14 2 7 15 4 13 16 15 4 4 3 13 3 1 9 10 13 0 2 9 2
2 11 2
42 10 9 9 13 10 0 11 9 9 7 9 0 1 9 2 15 13 10 9 9 13 10 9 7 11 11 13 10 0 9 7 9 16 10 9 9 9 14 13 1 9 2
20 3 0 9 4 15 13 14 13 10 11 9 16 13 10 0 11 9 9 9 2
32 15 4 13 10 9 9 1 16 13 10 9 1 10 9 9 2 15 4 3 13 1 10 0 9 10 4 13 10 9 1 9 2
9 4 15 13 15 13 14 13 0 2
4 9 2 11 11
4 3 15 13 2
2 11 2
5 13 10 13 9 2
9 13 15 13 16 15 13 10 9 2
2 11 2
16 10 9 13 3 0 1 10 9 15 13 3 10 0 9 3 2
7 13 15 0 1 10 9 2
3 10 9 2
8 10 9 2 15 4 3 13 2
2 9 2
2 11 2
21 13 4 10 11 0 12 9 1 9 1 10 9 12 14 4 13 1 10 9 9 2
2 9 2
10 0 9 13 1 12 13 5 12 12 2
15 10 9 1 9 13 13 1 10 0 9 13 5 12 12 2
9 10 9 13 3 1 1 10 13 2
23 5 12 12 2 13 9 9 2 11 2 11 2 11 2 11 2 7 11 11 2 2 5 13
11 5 12 12 2 11 9 9 2 5 14 13
19 5 12 12 2 0 9 1 11 9 1 1 9 9 13 1 12 2 5 13
8 9 1 10 9 4 13 3 2
22 3 2 9 1 10 9 13 13 9 1 11 1 9 1 11 14 9 9 4 13 3 2
9 6 13 15 1 9 16 15 13 9
2 9 2
1 11
2 11 2
7 0 16 3 13 15 9 2
5 11 13 3 0 2
10 6 13 7 13 15 13 15 15 13 2
10 13 15 13 16 15 13 3 0 11 2
2 9 2
2 11 2
2 11 2
19 3 13 10 9 9 7 10 0 9 1 10 9 15 13 1 15 0 11 2
19 16 15 4 13 15 4 13 9 1 10 3 0 9 1 9 7 0 9 2
15 15 4 3 13 9 15 13 3 0 1 15 0 0 9 2
22 16 15 13 9 15 4 13 10 9 13 15 14 13 15 7 2 7 13 15 15 9 2
4 13 15 11 2
1 11
35 11 11 11 9 9 1 0 9 11 11 11 11 12 11 11 2 9 2 12 11 2 11 12 9 2 12 9 2 12 9 2 12 9 2 12
2 11 2
4 13 15 13 2
2 11 2
1 11
16 10 1 2 9 9 1 11 12 2 4 13 3 0 14 13 2
28 1 10 9 9 2 9 4 13 3 0 14 13 9 0 16 15 4 13 2 11 2 11 2 11 2 0 2 2
11 15 13 10 9 1 9 13 1 10 9 2
22 11 4 13 0 14 13 9 2 7 10 1 10 9 4 13 1 1 10 12 9 9 2
18 2 1 9 11 13 7 13 1 1 2 9 4 13 12 9 3 3 2
19 15 4 13 1 11 1 10 9 1 10 9 7 9 4 13 12 9 3 2
33 11 4 14 13 1 1 9 16 15 13 1 10 9 7 10 0 9 7 9 13 14 13 10 9 1 10 9 10 4 14 4 13 2
7 14 10 0 9 1 9 2
34 10 9 9 13 1 10 11 9 7 15 13 0 1 15 9 9 2 11 7 11 13 10 0 12 9 14 13 1 12 5 1 9 2 2
11 4 13 9 9 7 9 9 1 11 3 2
33 15 4 13 14 13 10 9 1 10 0 1 2 9 9 0 2 7 16 9 16 15 13 2 10 0 9 4 13 11 12 2 12 2
12 16 15 13 9 7 9 2 6 13 15 13 2
1 9
3 11 11 12
2 11 2
36 15 4 13 16 13 10 9 9 1 15 9 2 3 2 15 13 15 4 13 14 13 3 12 9 1 9 1 11 14 13 1 11 14 9 2 2
36 16 15 13 1 15 2 16 1 10 9 15 4 14 13 11 9 2 15 4 13 14 13 1 9 9 10 4 13 14 13 10 9 1 15 9 2
9 15 1 2 9 9 13 11 12 2
41 16 15 13 16 11 12 4 13 0 1 16 13 10 9 2 9 1 10 0 9 1 1 10 9 10 13 4 13 1 15 1 1 0 11 9 2 6 13 15 13 2
29 11 4 3 13 15 16 15 4 13 13 9 2 9 1 15 9 16 15 13 13 10 1 2 9 9 1 11 12 2
2 9 2
2 11 2
29 13 1 10 11 9 1 9 11 13 15 4 13 9 1 10 0 9 2 2 0 9 2 9 2 3 1 9 12 2
35 15 9 13 16 1 3 7 3 11 2 10 9 13 10 9 7 9 14 13 10 9 1 9 2 10 4 13 0 1 9 2 9 14 9 2
26 9 4 13 15 11 13 1 9 7 9 2 13 1 9 1 0 2 7 11 4 9 2 13 10 9 2
2 0 2
12 13 15 4 13 15 2 7 13 14 13 0 2
10 15 13 3 10 9 1 9 4 13 2
17 15 13 2 15 13 1 10 9 7 4 14 13 3 15 4 13 2
10 15 4 13 16 15 4 13 14 13 2
2 9 2
2 0 2
1 11
16 9 1 10 9 2 10 0 9 1 15 9 4 13 1 9 2
15 16 15 4 14 13 2 11 4 13 15 13 9 1 9 2
14 15 4 13 2 9 2 16 3 15 4 3 13 3 2
7 15 4 13 15 10 9 2
2 0 2
1 11
6 13 10 2 9 9 2
16 9 2 10 9 13 1 9 9 7 10 9 1 10 11 11 2
4 11 12 2 12
3 1 11 11
4 10 11 11 11
1 11
35 10 9 11 9 4 13 9 14 13 13 12 9 1 9 9 7 9 15 13 11 14 9 9 14 13 16 15 13 1 9 14 13 9 9 2
49 10 0 9 2 13 1 9 11 11 11 2 11 2 11 11 2 4 13 1 10 9 1 9 0 9 13 1 0 0 9 9 7 9 16 15 4 13 10 9 1 10 11 2 2 10 9 9 2 2
46 9 7 9 9 13 16 10 9 2 13 1 10 9 15 13 10 9 14 9 9 2 13 10 11 9 9 2 13 10 9 1 10 9 2 13 9 7 13 13 9 1 9 1 9 9 2
41 10 0 9 1 10 9 9 13 16 11 11 2 10 9 1 10 11 11 11 2 13 3 3 15 13 9 14 13 0 9 9 13 14 13 10 9 9 9 4 13 2
27 11 13 15 0 9 7 11 11 11 3 15 13 10 12 2 9 9 14 13 10 9 2 9 7 9 13 2
21 2 15 4 14 13 3 10 9 4 4 13 9 1 10 0 9 2 2 13 11 2
32 10 9 4 13 15 13 2 13 11 2 14 13 13 9 1 10 9 1 10 9 2 7 14 13 1 9 2 0 9 7 9 2
17 11 9 11 11 13 10 11 13 2 0 2 1 10 9 1 11 2
26 2 10 11 13 15 13 10 13 9 2 3 15 13 10 13 9 13 1 10 0 9 2 2 11 13 2
13 11 13 9 2 13 10 9 1 10 0 9 9 2
14 11 9 11 11 13 11 14 9 4 13 10 0 9 2
20 10 9 4 13 1 11 0 9 16 12 9 1 9 2 14 13 10 9 3 2
18 1 10 9 2 9 4 13 14 13 9 1 11 1 1 10 9 9 2
10 2 15 13 10 9 2 2 11 13 2
8 2 15 13 14 13 9 2 2
31 15 13 0 1 10 9 9 13 1 11 12 3 11 9 9 13 1 0 9 1 10 9 1 9 9 9 4 13 1 9 2
28 10 9 4 13 9 3 0 1 5 12 1 9 2 3 12 9 1 10 5 12 1 9 9 1 12 9 3 2
37 2 15 2 9 9 2 13 7 13 10 5 12 9 9 2 7 10 0 9 1 11 13 3 0 2 2 13 11 2 15 9 4 4 13 1 11 2
7 2 10 9 13 3 2 2
29 9 13 16 1 11 12 2 9 9 7 9 9 13 9 1 10 11 11 11 11 2 13 16 10 0 9 4 13 2
22 10 9 2 12 1 10 2 4 13 1 12 9 1 10 0 7 13 9 1 9 9 2
43 2 16 3 13 3 2 10 2 11 2 9 9 4 13 9 1 10 9 2 13 9 7 13 0 9 1 9 9 2 2 13 12 9 13 1 11 11 9 9 11 11 12 2
34 16 15 13 9 0 16 10 9 13 3 14 13 1 9 9 2 11 13 10 9 7 0 9 1 10 0 9 13 0 9 1 9 9 2
28 15 13 10 0 9 1 10 9 4 13 14 13 16 9 13 14 2 13 2 9 2 10 4 13 0 9 9 2
29 1 10 11 12 9 2 9 9 13 0 9 16 16 9 9 4 14 13 15 4 13 1 10 9 1 10 9 9 2
6 10 9 13 15 9 2
13 10 0 9 2 10 0 9 13 10 0 9 9 2
16 15 4 13 1 9 13 10 5 12 9 9 13 12 9 3 2
23 9 9 3 13 15 9 16 13 10 9 2 13 15 4 14 13 10 9 3 1 10 9 2
30 15 13 14 13 9 1 11 2 7 1 11 12 10 11 13 15 0 9 12 9 7 13 1 9 2 10 4 3 13 2
22 15 13 10 0 9 4 13 1 10 11 7 11 14 13 10 0 9 1 10 9 9 2
35 11 2 15 1 15 9 1 9 7 0 13 9 1 10 11 2 13 10 12 2 9 9 9 2 13 0 9 14 13 10 5 12 9 9 2
12 0 9 16 13 10 9 13 1 10 0 9 2
27 7 10 11 9 2 10 4 13 10 9 9 2 7 10 9 13 1 11 14 9 16 10 9 4 4 13 2
36 1 9 2 10 9 15 13 13 10 9 9 2 11 11 2 13 1 10 9 1 9 1 10 11 7 11 9 9 3 9 16 10 9 4 13 2
8 15 4 14 13 9 1 15 2
14 2 1 9 2 15 4 4 13 15 2 2 11 13 2
17 16 10 9 9 0 2 10 9 13 9 1 0 9 13 0 9 2
39 2 10 11 9 13 1 10 9 1 10 9 14 0 9 9 1 9 9 2 3 13 10 9 1 9 10 4 13 1 1 10 3 0 9 2 2 11 13 2
14 2 15 13 1 9 16 15 13 14 13 9 3 0 2
25 10 9 13 10 9 14 9 1 9 7 13 10 11 14 13 10 9 1 10 9 2 13 9 2 2
25 9 1 9 13 1 10 9 1 5 12 10 9 1 5 12 10 9 1 12 9 2 11 9 13 2
12 11 13 10 13 9 1 9 13 5 12 12 2
18 11 13 10 9 2 13 12 9 1 10 9 2 13 1 1 13 11 2
12 9 2 15 13 2 4 14 13 1 10 9 2
21 3 15 13 10 13 9 1 0 9 2 10 4 13 14 13 9 9 14 13 9 2
21 11 13 10 9 9 13 10 11 14 13 9 4 9 1 9 4 13 1 0 9 2
16 2 15 13 10 9 15 13 13 10 0 9 2 2 11 13 2
18 2 1 15 9 2 15 4 14 13 15 13 7 13 0 10 0 9 2
17 15 13 15 13 15 0 16 15 13 10 9 1 9 7 9 2 2
37 11 11 2 11 2 15 13 10 11 9 9 1 10 9 7 0 9 1 10 9 10 13 9 9 2 13 11 4 14 13 15 16 13 10 9 9 2
19 11 2 11 3 13 15 13 0 16 9 1 10 9 2 9 9 4 13 2
21 2 11 13 15 1 15 2 2 13 11 2 11 2 0 9 1 10 11 11 11 2
20 2 15 13 15 15 13 13 14 4 13 1 10 9 14 13 10 9 13 2 2
16 10 11 9 13 10 9 9 10 0 9 13 11 13 15 9 2
28 10 9 9 13 14 13 11 13 2 7 15 13 9 0 9 4 13 1 0 9 2 10 11 14 9 11 13 2
22 11 11 11 2 10 0 11 11 11 11 9 2 13 13 10 11 9 7 3 13 11 2
22 2 15 13 10 9 9 2 7 15 13 14 3 14 13 11 13 0 2 2 11 13 2
16 2 15 2 11 9 2 13 15 10 0 9 9 4 13 2 2
14 15 11 14 9 13 14 13 13 3 10 10 9 13 2
19 15 13 9 7 9 1 10 9 1 11 14 11 12 9 4 13 0 9 2
24 2 15 4 14 13 3 15 13 15 15 13 2 7 15 13 0 14 13 1 2 2 11 13 2
25 2 11 13 15 13 10 9 1 10 9 1 11 2 7 15 13 10 9 13 10 9 1 9 2 2
25 15 4 13 11 11 14 9 7 13 15 1 10 9 1 10 9 14 13 13 10 9 1 10 9 2
10 15 4 13 15 1 16 15 4 13 2
4 11 7 11 2
34 15 4 13 10 9 1 11 7 11 11 1 11 14 13 15 9 1 10 9 14 13 15 0 9 1 11 2 1 9 3 1 9 2 2
9 4 15 13 15 9 7 3 3 2
33 15 9 13 16 10 9 4 13 0 1 15 2 3 2 2 7 15 9 12 9 13 14 13 14 13 10 11 9 13 1 10 9 2
11 10 9 16 3 11 7 11 4 13 3 2
2 9 2
3 13 0 2
35 15 13 10 2 0 9 2 1 10 9 2 0 9 7 9 1 10 9 2 7 1 1 10 9 2 10 9 1 10 13 9 1 12 9 2
5 13 15 10 9 2
10 15 4 13 1 11 14 13 10 9 2
25 16 15 13 2 11 2 11 7 15 3 13 1 12 9 2 7 15 13 0 14 13 1 10 9 2
2 0 2
1 11
5 4 15 13 9 2
11 7 16 6 2 15 13 10 9 7 9 2
1 11
8 2 11 11 11 2 2 8 2
3 12 12 9
10 15 13 10 12 9 9 2 3 3 2
8 4 15 13 10 9 16 13 2
22 15 13 9 0 1 10 0 9 2 7 9 3 0 16 13 12 10 13 3 1 9 2
10 3 1 10 9 1 10 9 1 15 2
12 3 13 10 2 0 2 9 1 10 9 9 2
67 16 15 4 13 9 2 15 13 15 4 13 11 1 9 16 15 9 13 14 1 9 1 10 9 2 16 15 13 1 10 9 2 7 16 15 9 13 3 10 0 9 10 4 13 1 10 9 2 16 11 3 4 14 13 15 0 9 1 10 9 2 4 3 13 15 2 2
36 3 2 10 0 9 13 1 9 13 16 15 9 2 10 0 9 7 3 10 9 15 13 14 13 2 13 7 13 14 10 0 9 1 10 9 2
4 15 13 15 2
1 9
2 8 8
3 12 12 9
30 1 11 11 9 2 4 15 6 13 15 10 9 2 9 1 9 15 13 1 11 11 11 1 10 9 1 11 7 11 2
41 1 9 2 4 15 13 1 10 9 3 14 13 16 15 13 10 0 9 1 15 9 10 13 9 1 11 2 16 15 4 13 15 13 10 1 15 13 9 1 11 2
5 9 1 15 9 2
14 2 11 11 2 4 15 13 10 9 1 9 7 9 2
19 2 11 11 2 4 15 13 10 9 1 9 9 7 9 2 0 9 9 2
13 9 2 11 11 2 11 11 2 11 11 2 11 11
19 0 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11
14 0 9 2 11 11 2 11 11 2 11 11 2 11 11
4 9 2 11 11
12 9 2 9 2 11 11 2 11 11 2 11 11
4 9 2 11 11
1 11
2 13 0
3 11 11 11
3 12 12 9
2 11 2
5 3 4 15 13 2
34 16 15 4 13 10 0 9 1 11 11 9 2 15 4 13 14 13 16 15 13 1 11 11 16 13 15 13 1 11 14 9 1 9 2
7 9 1 15 9 10 9 2
1 11
25 1 10 12 9 15 4 13 3 2 15 13 0 1 10 11 2 11 0 9 9 1 10 9 9 2
3 9 0 2
7 16 3 2 6 13 11 2
2 8 8
3 12 12 9
28 11 2 15 13 10 9 1 10 0 9 9 11 13 13 1 11 7 15 4 13 11 11 15 13 0 9 3 2
17 15 4 13 10 9 15 13 7 13 15 13 14 13 10 9 3 2
24 11 4 15 13 10 0 9 9 13 1 10 9 1 11 7 13 15 0 1 10 11 4 13 2
17 15 13 11 11 0 9 7 15 4 14 13 13 10 0 9 9 2
9 15 13 3 2 10 0 9 3 2
1 11
2 11 2
8 4 15 13 15 9 1 11 2
34 15 13 10 9 1 10 15 4 13 15 9 13 2 2 8 2 4 15 13 10 0 9 1 10 9 1 0 9 9 13 1 11 11 2
18 2 8 2 13 15 0 16 11 13 12 9 1 0 9 9 1 11 2
16 2 8 2 13 15 0 1 10 9 9 1 11 15 13 15 2
12 6 13 15 10 9 16 15 4 13 14 13 2
1 11
15 14 3 15 13 3 2 7 15 13 14 3 10 0 9 2
4 11 7 11 2
14 13 15 0 14 13 10 2 0 9 2 9 9 9 2
45 16 15 13 10 9 9 2 15 4 13 3 0 16 12 1 15 4 13 15 10 9 14 13 10 9 2 15 13 15 4 13 1 11 14 9 3 1 15 1 9 1 3 0 9 2
1 11
1 5
5 10 9 13 0 2
17 15 4 3 13 0 7 3 13 1 9 9 9 7 0 0 9 2
34 16 15 4 13 15 1 9 6 13 15 13 1 9 7 3 13 15 1 15 9 2 15 4 14 13 10 9 7 13 15 9 1 9 2
1 5
9 13 15 1 11 11 1 15 9 2
2 9 2
2 8 8
3 12 12 9
2 11 2
10 1 15 9 9 2 3 13 10 9 2
23 16 15 13 2 6 13 15 13 3 15 13 0 2 7 15 4 13 9 14 13 15 1 2
6 13 15 1 15 9 2
2 11 12
1 8
5 11 11 2 8 2
3 12 12 9
3 6 11 2
13 4 15 13 16 10 11 4 13 0 11 11 3 2
16 3 2 13 15 1 11 14 9 2 16 15 4 13 15 3 2
9 13 15 8 11 9 4 13 3 2
1 11
2 2 9
16 16 15 4 13 1 10 9 1 15 9 2 15 4 4 13 2
9 6 13 15 14 13 10 9 9 2
3 8 8 8
3 12 12 9
23 3 16 11 13 1 15 9 2 4 15 13 14 13 15 13 10 9 9 1 11 1 15 2
10 15 4 13 15 10 9 1 15 9 2
5 13 15 14 13 2
2 11 11
3 12 12 9
24 1 1 9 2 15 4 14 13 9 1 0 16 13 1 11 11 14 9 13 11 12 2 12 2
11 15 4 13 10 9 1 5 12 1 12 2
16 11 2 6 13 15 13 15 15 13 14 13 3 14 13 9 2
5 8 1 12 12 9
12 10 13 9 4 4 13 1 15 1 11 11 2
9 2 13 13 9 2 8 8 9 2
4 2 8 8 9
3 11 11 11
3 12 12 9
10 15 4 13 15 10 9 1 15 9 2
5 13 15 14 13 2
2 11 11
3 12 12 9
24 1 1 9 2 15 4 14 13 9 1 0 16 13 1 11 11 14 9 13 11 12 2 12 2
11 15 4 13 10 9 1 5 12 1 12 2
16 11 2 6 13 15 13 15 15 13 14 13 3 14 13 9 2
8 4 11 13 16 13 10 9 2
1 8
3 12 12 9
21 3 13 10 13 9 1 10 9 2 9 2 7 9 9 1 11 14 9 14 13 2
17 16 15 4 13 2 15 13 15 13 10 9 1 10 9 14 9 2
19 15 4 4 13 10 9 9 3 16 15 4 13 14 13 1 1 15 9 2
38 15 13 3 1 11 11 15 9 13 9 11 4 13 13 3 10 9 14 9 1 9 1 10 9 2 9 1 10 9 9 7 10 9 10 9 4 13 2
11 16 15 13 3 2 15 4 13 15 3 2
12 13 14 13 10 9 1 10 9 14 9 9 2
2 9 2
2 6 2
8 13 1 11 7 10 9 9 2
14 10 9 14 13 4 3 13 1 11 12 1 12 9 2
18 10 9 14 9 9 13 3 0 11 12 7 11 9 13 0 11 12 2
10 15 13 15 9 13 10 9 11 13 2
6 15 13 10 1 3 2
2 2 11
3 2 9 2
20 10 9 13 1 10 9 9 4 13 3 1 9 1 10 9 7 9 13 3 2
44 16 10 9 1 10 9 13 14 10 13 9 2 7 10 9 7 9 0 14 13 15 1 10 13 9 2 15 4 3 13 16 10 9 2 9 7 9 1 10 9 4 3 13 2
25 16 15 4 13 10 9 1 9 2 6 3 13 15 1 9 2 12 2 2 7 13 10 0 9 2
3 13 15 2
7 2 11 11 2 2 8 2
3 12 12 9
4 0 11 11 2
1 2
29 16 15 13 10 15 10 9 9 1 10 9 1 15 9 2 15 13 15 4 13 15 10 0 9 1 9 3 3 2
1 2
15 15 13 3 3 0 16 13 11 13 15 9 9 9 9 2
41 15 4 13 0 9 1 9 0 1 11 2 11 11 2 11 11 7 11 11 2 7 15 4 13 0 14 13 10 9 15 4 13 1 10 0 9 1 15 0 9 2
26 10 0 9 1 15 9 2 3 2 13 0 1 10 9 15 4 13 14 13 10 0 9 1 10 9 2
27 15 13 10 9 1 10 9 9 10 4 4 13 10 11 11 11 14 9 9 9 7 9 1 9 9 9 2
23 1 10 9 15 4 13 3 0 13 9 14 13 10 1 15 9 7 13 15 0 9 9 2
29 3 15 9 9 2 1 1 3 12 1 15 9 9 2 4 13 14 13 1 10 9 1 11 9 1 10 10 9 2
28 3 10 9 4 13 1 12 1 12 9 1 9 2 9 2 7 9 16 16 15 13 0 0 9 1 15 9 2
27 1 10 9 15 4 13 15 1 10 0 9 1 15 13 9 9 7 10 9 1 9 1 9 1 10 9 2
26 10 0 9 1 10 9 4 13 16 3 15 4 13 10 9 14 13 10 9 1 9 13 1 9 9 2
14 15 13 3 0 16 13 9 10 13 0 1 10 9 2
22 15 4 13 14 13 1 11 12 7 2 11 12 2 16 9 1 15 9 13 3 0 2
25 6 13 15 13 15 13 0 2 7 13 0 14 13 15 10 9 16 15 13 10 9 2 12 2 2
1 2
2 9 2
2 5 11
12 11 11 9 9 11 11 11 2 12 2 12 12
8 2 11 11 11 2 2 8 2
3 12 12 9
4 9 2 11 2
9 4 15 13 10 9 9 1 11 2
2 9 2
2 8 8
3 12 12 9
19 15 4 13 10 9 1 10 9 13 1 10 9 3 3 16 15 13 15 2
1 11
8 2 11 2 11 2 2 8 2
3 12 12 9
3 6 9 2
7 6 2 3 15 13 0 2
6 7 15 13 3 0 2
48 10 9 1 11 11 14 0 0 7 9 9 9 4 4 13 14 13 1 10 0 9 7 9 1 11 9 9 1 10 9 14 13 10 9 9 10 4 13 11 11 7 10 9 1 11 10 9 2
18 10 9 9 4 4 13 14 13 10 9 9 9 9 14 4 13 9 2
6 3 2 12 9 5 9
25 3 2 12 11 11 11 2 1 11 7 11 2 9 12 11 11 1 11 2 11 2 11 7 11 12
15 15 2 9 1 10 13 9 4 4 13 0 1 10 9 2
18 11 14 0 9 7 10 9 9 4 13 0 14 13 9 1 10 9 2
17 15 13 0 16 15 4 13 10 9 1 10 11 9 9 3 9 2
1 2
19 2 9 13 10 0 9 2 1 1 10 9 16 15 13 1 15 0 9 2
21 11 11 0 9 11 11 14 11 11 12 11 11 9 12 11 11 2 11 12 12 8
11 10 9 1 9 7 9 2 15 13 15 2
25 9 13 2 1 7 1 15 2 10 0 9 2 7 15 3 3 13 1 9 7 9 3 3 13 2
11 3 4 15 13 10 10 9 2 13 15 2
24 13 1 15 7 13 10 10 9 13 9 9 9 3 3 15 4 14 4 13 2 7 15 13 2
12 15 13 10 9 15 13 11 11 1 10 9 2
28 15 13 10 9 15 4 13 9 2 1 1 10 9 10 0 9 4 13 1 10 8 0 9 2 15 13 3 2
12 7 15 4 13 16 13 15 15 13 10 9 2
15 14 3 2 9 13 15 9 13 7 4 13 15 15 13 2
11 15 13 3 9 13 7 9 13 1 15 2
6 15 4 3 3 13 2
43 15 13 10 0 9 3 3 15 13 1 15 9 7 4 14 13 14 13 16 16 15 13 14 13 9 2 15 13 3 9 14 13 1 7 13 10 0 9 9 1 10 9 2
6 3 0 9 13 15 2
24 7 15 13 10 0 9 1 10 3 0 2 0 2 9 9 13 9 0 9 10 4 13 15 2
57 3 15 13 15 10 1 9 2 15 13 9 14 14 13 9 7 3 3 3 3 15 13 9 1 13 1 9 15 4 3 13 2 13 2 13 9 2 13 10 9 7 10 9 9 3 16 15 13 3 0 14 13 15 15 4 13 2
16 9 1 15 4 3 13 15 9 2 7 4 15 13 15 9 2
9 13 1 15 9 2 13 15 15 2
4 3 15 13 2
3 13 15 2
16 13 13 14 13 15 9 1 1 9 14 2 13 10 9 2 2
32 15 13 10 9 14 13 10 9 2 15 4 14 13 10 9 16 15 13 3 2 15 13 10 9 10 15 13 7 15 13 9 2
3 0 9 2
21 3 16 15 13 0 2 4 14 13 15 10 9 14 13 1 10 10 9 1 15 2
29 10 9 15 4 13 1 10 10 0 9 0 9 3 2 9 2 13 1 16 13 9 7 13 1 9 1 10 9 2
11 15 13 10 0 9 15 13 2 9 2 2
6 15 4 4 13 1 2
3 2 8 2
3 2 8 2
24 15 13 16 11 13 0 14 13 3 1 15 0 9 1 10 11 9 10 13 3 12 9 3 2
28 3 2 11 9 7 9 13 3 0 1 2 9 2 9 16 10 0 9 1 10 0 9 1 10 11 9 13 2
62 10 3 0 9 13 14 16 11 13 3 0 14 13 1 0 9 9 7 9 9 2 7 16 10 9 15 4 13 1 10 0 9 3 0 1 11 7 11 2 9 10 13 1 1 10 9 9 10 13 9 7 13 9 1 9 2 9 7 9 2 9 2
4 15 13 3 2
27 13 10 2 11 2 9 4 13 3 0 2 15 13 1 1 15 3 1 10 9 3 15 13 1 11 2 2
21 15 4 14 13 10 9 16 13 10 9 13 9 10 13 15 9 13 1 10 9 2
37 3 12 9 15 4 13 9 9 2 2 3 15 4 13 1 10 0 9 2 16 15 4 13 16 11 13 0 9 3 16 13 14 13 10 0 9 2
36 15 4 13 14 13 11 9 1 10 9 16 15 4 13 10 2 9 16 13 9 2 9 10 3 13 1 10 9 16 13 9 1 10 11 9 2
29 3 15 4 13 9 14 13 3 16 15 13 10 0 9 2 16 15 13 0 16 13 9 4 13 1 0 9 2 2
10 7 9 4 13 10 0 9 9 1 2
24 3 2 10 9 4 13 3 16 13 10 0 9 13 1 10 0 7 3 0 2 0 0 9 2
31 10 0 9 3 2 9 9 1 10 11 11 11 13 10 9 2 0 9 1 9 1 12 0 9 16 10 0 9 14 13 2
26 15 13 10 0 9 14 13 9 1 10 0 2 0 9 16 1 9 2 9 10 11 9 4 4 13 2
21 10 0 13 10 0 9 9 2 13 2 1 11 14 14 13 3 0 9 1 9 2
11 11 13 10 9 9 14 13 1 10 9 2
33 7 13 15 13 1 15 9 2 7 10 9 1 10 9 9 3 3 2 16 15 4 13 15 9 7 13 10 9 1 9 9 3 2
2 11 2
1 2
11 13 1 11 11 1 11 11 1 12 12 9
4 13 10 0 9
38 1 11 11 14 0 9 2 11 2 9 13 10 9 13 1 10 0 9 9 14 13 9 13 12 0 9 1 10 0 9 0 16 2 9 13 9 2 2
9 15 13 10 9 16 13 1 9 2
73 12 1 15 3 13 9 13 10 9 16 15 13 3 0 9 1 10 9 14 13 15 0 9 7 1 10 0 9 15 13 3 12 2 16 15 13 10 9 1 15 7 15 2 15 13 3 3 1 10 9 13 9 2 15 0 9 2 10 9 7 10 9 2 10 9 7 10 9 2 10 1 15 2
27 15 4 13 10 9 3 16 13 10 9 3 9 3 13 10 0 9 16 13 15 0 9 2 9 7 9 2
18 13 1 10 9 2 16 15 4 2 1 12 0 9 7 12 0 9 2
9 15 9 13 1 15 9 7 9 2
8 10 0 9 7 15 10 13 2
11 10 9 1 10 0 9 13 15 10 3 2
26 13 1 1 9 1 9 13 10 0 9 2 1 15 13 10 10 9 15 4 13 14 13 1 1 9 2
39 15 13 3 3 0 1 15 0 2 15 13 3 3 0 1 10 0 1 15 2 13 9 7 13 1 10 9 13 15 10 9 16 15 13 0 13 10 9 2
16 3 10 0 13 10 9 1 9 7 9 15 13 15 10 3 2
35 3 15 0 3 3 14 13 9 13 10 9 1 9 7 9 1 15 1 15 15 13 2 3 3 4 15 13 15 2 7 15 4 13 15 2
13 15 13 10 9 1 10 0 9 15 10 13 1 2
14 15 15 13 4 3 13 3 14 7 13 7 13 15 2
31 15 4 3 13 1 10 9 1 15 9 1 10 9 2 15 9 1 10 0 1 10 0 2 7 15 9 1 9 1 9 2
16 11 13 16 15 15 13 10 0 1 10 9 15 13 1 15 2
11 15 4 15 13 1 10 0 1 10 9 2
14 16 15 13 3 1 10 9 3 2 13 15 13 3 2
27 13 16 15 15 13 1 15 13 15 7 9 0 2 13 16 15 15 13 1 15 7 9 0 13 15 9 2
28 3 3 10 9 15 13 1 9 16 13 0 2 15 4 3 13 0 9 16 15 3 13 14 13 10 0 9 2
17 3 9 4 13 15 9 3 16 15 0 0 9 4 14 13 3 2
12 1 10 0 9 0 9 4 13 14 4 13 2
22 4 15 13 14 13 1 9 1 10 9 7 13 7 13 1 10 9 1 9 7 9 2
23 4 15 13 14 13 1 9 7 9 7 13 3 13 7 13 16 13 1 1 9 7 9 2
12 15 13 10 9 1 9 7 10 9 1 9 2
2 11 12
7 11 11 2 11 11 2 11
8 11 11 9 2 9 0 0 9
4 12 0 9 2
4 12 0 9 2
6 15 4 15 13 1 2
4 0 0 9 2
6 0 9 1 15 9 2
3 0 9 2
8 9 1 10 9 1 0 9 2
44 16 15 4 13 1 10 9 2 9 9 14 13 13 1 15 9 7 15 4 13 1 10 9 13 16 13 1 9 1 10 0 9 9 2 11 13 10 9 10 4 13 15 13 2
20 11 13 10 0 9 7 4 3 13 14 13 10 0 9 1 10 9 9 9 2
11 10 9 4 13 10 3 0 9 1 9 2
11 13 13 9 1 10 0 9 2 13 9 2
2 0 9
11 11 13 10 3 0 9 1 9 13 9 2
14 10 9 4 13 10 0 7 0 9 9 1 0 9 2
13 10 0 9 9 9 13 0 0 9 9 1 9 2
29 1 10 9 9 2 15 9 4 3 13 13 10 9 1 10 9 9 16 10 9 1 9 2 9 7 9 4 13 2
14 3 3 4 10 10 0 9 13 0 16 13 0 9 2
5 13 10 9 9 2
10 10 9 13 2 1 1 9 7 9 2
14 0 9 9 1 10 0 9 2 10 9 7 9 9 2
9 0 9 9 2 13 10 9 9 2
9 0 1 15 1 9 13 9 7 9
11 0 2 3 0 2 9 1 10 9 13 0
2 0 9
12 11 4 13 10 0 9 9 10 13 3 0 2
20 15 13 15 9 16 10 9 9 4 13 10 1 10 0 9 1 9 9 9 2
21 10 9 4 14 4 13 1 10 9 2 10 9 2 10 9 2 7 10 13 9 2
6 15 13 10 0 9 2
6 15 13 0 9 9 2
7 15 13 14 3 9 9 2
23 16 15 13 14 13 5 12 12 7 3 3 13 5 12 12 2 15 13 14 0 9 9 2
23 12 9 3 15 9 4 3 13 10 0 7 0 2 13 10 9 1 0 2 9 0 9 2
21 10 11 9 9 13 10 9 10 13 10 9 4 4 13 1 15 15 13 1 15 2
6 13 15 0 1 11 2
10 13 9 14 13 10 0 9 1 11 2
20 10 9 4 13 10 9 1 0 9 9 2 7 15 9 7 9 2 11 11 2
5 10 9 4 13 2
74 15 4 13 2 2 3 14 13 10 9 1 0 9 2 2 3 11 13 10 0 9 14 13 15 9 2 2 10 0 0 9 1 10 9 2 2 3 10 2 9 2 9 2 13 0 9 9 3 2 2 10 9 9 1 9 14 13 15 13 3 2 7 2 10 9 14 13 1 10 2 9 2 9 2
7 3 13 10 9 14 13 2
3 12 7 12
7 10 9 14 13 13 2 12
8 9 2 11 2 11 12 2 12
7 9 2 12 9 11 11 11
4 9 2 9 9
11 12 9 2 12 9 2 12 9 2 12 9
6 15 4 13 15 3 2
4 11 11 12 12
8 9 2 2 11 2 2 8 2
1 6
3 6 10 2
16 15 3 13 10 9 9 2 10 13 0 1 7 1 9 9 2
15 15 13 15 14 13 10 9 2 16 15 13 0 0 9 2
10 15 13 10 9 1 7 9 7 9 2
1 11
1 2
14 9 13 10 9 10 4 13 1 12 1 11 11 11 2
15 15 13 10 0 9 7 13 10 9 16 13 9 7 9 2
7 9 13 3 0 1 9 2
23 15 4 13 1 7 13 10 9 1 9 2 13 10 9 0 7 13 10 0 9 1 9 2
16 9 13 1 10 11 9 2 9 2 13 9 7 9 1 9 2
17 10 9 1 10 9 13 13 1 10 0 9 1 9 2 9 2 2
27 3 9 13 10 9 1 10 9 2 9 9 2 1 15 9 14 13 10 9 1 10 9 2 0 9 2 2
9 10 9 4 3 13 1 1 9 2
1 2
2 10 9
11 13 10 10 9 7 9 1 9 1 9 2
3 13 9 2
7 13 1 0 9 1 9 2
6 10 9 4 13 0 2
15 9 1 10 9 2 9 2 9 7 0 9 4 4 13 2
14 9 1 10 9 2 9 2 9 7 9 4 4 13 2
7 10 9 13 0 7 0 2
7 9 1 9 4 4 13 2
6 0 9 4 13 0 2
10 9 1 10 9 7 9 4 4 13 2
6 13 9 1 10 9 2
10 13 9 7 9 1 10 9 7 9 2
3 13 9 2
3 13 9 2
3 13 9 2
3 13 9 2
6 9 9 4 4 13 2
5 9 4 4 13 2
11 13 1 9 2 9 7 13 15 14 9 2
20 0 9 2 9 2 9 2 9 1 9 2 0 9 2 0 9 4 4 13 2
21 13 9 7 9 9 9 2 0 9 2 9 2 9 2 9 2 9 7 9 9 2
13 13 10 9 14 13 1 12 5 12 9 1 9 2
1 2
2 10 9
10 10 12 9 1 10 9 4 13 3 2
18 3 10 9 13 1 10 9 9 2 10 9 3 7 13 1 10 9 2
35 3 1 10 9 1 2 6 2 6 2 2 2 6 2 6 2 2 10 9 13 15 9 2 13 10 0 9 1 10 9 1 10 0 9 2
16 1 10 0 12 9 2 10 9 3 13 15 9 1 10 9 2
12 9 4 4 13 1 3 0 9 16 15 13 2
1 2
2 10 9
25 3 10 9 13 10 9 1 10 9 1 2 6 2 6 2 2 2 10 0 9 4 3 4 13 2
5 3 13 10 9 2
28 10 12 9 3 13 7 13 3 13 2 2 3 15 4 13 14 13 10 9 1 9 9 2 0 9 2 2 2
17 13 1 10 9 13 2 2 15 13 10 0 9 14 13 15 2 2
16 13 1 10 9 13 2 2 15 13 3 14 13 15 9 2 2
12 13 3 13 2 2 15 3 13 1 15 2 2
17 13 3 13 2 2 15 13 0 14 13 10 9 10 4 13 2 2
16 10 0 12 9 13 2 2 6 11 15 13 15 0 9 2 2
5 11 13 11 9 9
2 11 2
32 10 11 9 4 13 10 11 11 1 9 1 11 16 13 12 9 16 13 1 10 0 9 1 10 9 9 12 9 3 1 11 11
40 11 11 11 2 12 2 1 11 2 11 2 13 10 9 9 14 13 10 0 9 1 11 11 2 3 3 1 10 11 11 2 14 13 12 9 15 4 4 13 2
41 2 10 1 10 9 7 10 1 10 9 15 13 13 1 1 10 9 13 10 9 16 15 13 9 1 10 11 2 11 2 9 3 15 4 13 2 2 11 11 13 2
39 11 11 2 10 9 2 13 15 13 3 3 12 0 9 1 10 0 9 1 11 11 1 11 12 3 15 13 15 15 13 13 10 9 13 1 15 9 9 2
14 2 15 0 9 13 14 13 15 3 2 2 15 13 2
29 2 10 0 9 3 15 9 13 10 9 1 10 9 14 9 1 10 9 9 7 3 15 13 13 1 10 9 2 2
11 10 0 9 13 3 0 1 0 0 9 2
20 10 0 3 13 0 9 10 9 7 10 0 9 13 9 10 9 2 9 13 2
35 10 12 13 14 13 10 9 7 13 15 9 1 10 9 0 9 3 7 10 9 13 1 10 9 7 13 13 12 2 9 2 0 11 11 2
10 2 15 9 13 2 2 11 11 13 2
17 2 15 13 15 9 7 15 9 7 13 15 9 7 13 3 2 2
21 10 9 13 10 12 2 9 2 12 11 11 2 13 15 1 10 9 2 15 13 2
37 11 11 13 10 0 9 1 10 9 2 13 15 7 13 11 14 13 7 15 3 13 1 12 2 9 2 0 11 11 2 15 13 1 10 0 9 2
17 3 11 11 13 9 1 10 9 7 3 15 9 13 0 14 13 2
14 2 10 9 13 9 7 15 13 9 2 2 15 13 2
18 2 1 10 9 2 11 13 7 10 9 13 15 7 13 1 15 9 2
27 15 13 1 10 9 14 9 7 15 13 15 1 10 0 9 1 10 9 1 10 9 10 9 1 9 2 2
5 10 9 13 3 2
27 16 15 13 10 9 7 9 1 10 12 2 9 9 2 11 11 13 15 4 14 13 15 13 10 0 3 2
13 7 11 11 7 11 11 2 3 2 4 13 3 2
18 11 11 7 15 9 13 12 9 3 7 13 12 9 1 10 11 11 2
16 11 11 13 10 12 9 1 9 14 13 9 1 10 0 9 2
31 7 11 11 7 11 11 4 13 1 10 9 7 13 2 16 11 11 13 10 9 1 10 9 1 15 9 2 11 11 13 2
15 11 11 13 12 1 12 9 14 13 10 11 11 1 11 2
28 10 9 9 4 13 1 9 15 2 13 15 9 1 10 0 9 16 13 7 13 14 13 10 9 1 9 2 2
41 10 0 0 9 1 10 9 13 11 11 11 2 12 2 1 11 2 15 4 13 11 12 2 12 2 16 13 14 13 10 11 9 9 9 1 10 9 13 10 9 2
16 11 11 13 0 9 1 10 9 16 15 4 13 1 10 9 2
25 11 9 11 11 13 10 9 9 1 12 16 4 13 1 9 9 1 10 9 9 10 13 12 9 2
12 10 9 13 1 10 5 12 2 11 2 9 2
5 0 9 1 0 9
2 11 11
10 15 13 10 0 9 1 9 11 11 2
36 15 13 12 9 0 16 13 10 9 1 10 9 2 7 15 13 14 13 15 9 11 11 16 10 0 9 4 14 13 10 0 9 1 12 9 2
1 11
9 15 13 14 10 9 16 3 13 2
7 15 13 0 1 11 11 2
1 11
20 10 9 4 13 16 13 9 2 1 9 2 7 9 14 13 10 0 0 9 2
1 11
13 10 9 4 13 1 10 9 14 9 11 11 11 2
7 15 13 1 11 11 11 2
1 11
22 10 9 13 1 10 9 13 1 10 9 1 9 10 9 2 9 4 13 0 14 13 2
21 15 4 3 13 2 11 2 2 10 9 1 10 9 13 1 12 13 1 12 9 2
29 16 9 2 11 9 9 11 11 7 11 11 13 15 9 1 10 9 9 2 15 13 10 9 13 1 1 2 11 2
1 11
20 9 11 11 13 10 9 16 13 9 1 10 9 1 10 9 3 1 10 9 2
48 3 11 11 13 3 1 10 9 9 1 10 9 9 2 15 13 10 9 1 9 13 1 2 9 2 7 3 13 1 11 16 15 13 10 9 2 9 2 2 10 9 9 13 14 13 9 9 2
11 15 4 3 13 1 1 11 1 0 9 2
2 11 11
26 11 11 7 11 11 13 10 9 14 13 16 10 9 15 13 4 4 13 11 2 11 7 11 2 11 2
1 11
36 11 11 7 11 11 13 14 13 15 0 9 2 11 11 2 7 15 4 3 13 1 10 9 9 3 15 13 14 13 1 10 9 1 0 9 2
4 11 2 11 2
19 11 11 13 10 9 1 15 9 1 2 10 9 9 2 7 2 9 2 2
14 11 13 14 13 10 9 1 11 11 1 11 11 11 2
1 11
15 13 1 11 11 14 13 10 9 10 13 0 1 9 9 2
15 3 13 11 2 11 2 10 2 5 2 4 13 3 3 2
1 11
17 9 11 11 13 3 1 10 9 3 15 9 13 13 9 1 9 2
11 10 0 9 9 1 10 9 4 13 11 2
1 11
20 11 11 7 11 11 4 13 1 10 9 9 1 10 11 2 11 11 11 2 2
28 10 9 9 1 10 9 4 13 11 2 10 11 13 15 1 10 9 14 13 9 1 10 9 7 9 0 2 2
15 10 9 4 13 14 13 13 10 3 13 9 9 1 11 2
22 10 9 3 4 13 7 11 7 11 13 14 13 15 15 13 7 13 15 1 10 9 2
11 15 13 10 9 11 7 13 10 11 9 2
10 3 15 13 10 0 9 1 10 9 2
1 11
28 15 13 1 10 11 9 2 9 2 13 9 2 7 2 9 2 10 9 13 1 11 14 13 1 10 0 9 2
1 11
16 13 1 12 11 11 9 2 11 13 10 9 1 11 11 11 2
34 9 11 13 10 9 2 11 11 13 15 7 11 11 14 13 9 13 1 15 2 7 11 11 14 13 10 11 2 0 9 1 10 9 2
1 11
18 10 9 4 13 1 11 11 7 13 1 15 9 2 11 14 11 2 2
16 15 13 10 9 15 13 0 1 9 7 9 7 13 3 0 2
16 11 9 11 11 7 11 11 13 10 9 16 15 13 15 9 2
5 15 13 1 11 2
9 9 2 8 9 2 5 12 9 2
3 6 10 2
21 15 13 3 0 9 1 10 9 13 16 13 11 11 2 3 3 13 10 0 9 2
5 15 13 3 14 2
26 10 0 9 13 11 13 3 0 1 10 0 9 7 15 4 13 13 16 15 4 14 13 14 13 3 2
15 15 4 13 0 9 9 3 13 1 9 7 1 10 9 2
20 3 15 13 16 10 9 1 10 9 4 3 3 13 10 9 1 9 4 13 2
29 15 13 2 10 9 1 10 9 4 13 1 11 7 3 4 13 0 7 15 4 3 13 15 0 9 14 13 5 2
27 15 13 9 0 1 10 0 9 1 10 9 15 7 15 13 16 10 9 4 13 10 9 1 0 9 9 2
2 9 2
1 11
2 6 2
4 0 9 9 2
9 15 4 3 13 3 1 11 11 2
6 9 13 10 9 9 2
2 11 12
26 11 12 13 10 13 9 9 2 16 11 11 4 13 1 9 1 11 2 3 11 12 4 13 11 12 2
23 3 2 15 13 14 13 10 9 7 10 9 4 13 15 3 15 13 1 1 12 9 9 2
14 6 6 2 15 4 13 15 3 15 13 1 1 11 2
8 9 13 11 12 1 10 9 2
25 7 15 13 16 15 4 13 3 3 16 15 13 14 13 1 10 10 9 3 15 3 13 3 3 2
32 3 3 1 8 9 13 1 7 15 13 10 9 1 0 9 10 13 15 15 13 3 10 0 9 10 15 4 13 15 1 1 2
13 7 10 0 9 16 13 10 9 2 9 9 6 5
12 15 13 3 3 0 2 15 3 13 11 11 2
7 15 4 14 13 1 15 2
15 13 1 10 11 11 9 9 1 1 0 9 1 10 9 2
9 15 13 10 0 9 9 9 9 2
28 10 9 13 1 10 9 10 1 10 0 9 15 4 3 13 1 10 9 7 15 4 4 13 1 10 9 9 2
6 15 13 0 10 9 2
17 15 13 10 9 7 4 3 13 13 10 0 9 14 13 0 9 2
14 15 4 13 1 10 10 9 9 9 7 10 9 9 2
8 10 9 13 3 12 5 0 2
15 15 4 14 13 15 3 13 0 14 13 10 11 12 9 2
9 0 9 1 10 1 10 11 9 2
17 15 13 11 11 7 15 13 1 10 11 11 11 11 1 11 11 2
28 15 13 10 9 1 0 0 9 10 4 13 1 12 1 11 7 15 4 3 13 11 1 10 9 1 9 13 2
8 10 9 13 10 3 0 9 2
28 15 4 13 14 13 0 0 9 15 13 3 3 0 14 13 3 1 10 9 7 13 15 0 9 14 13 1 2
31 15 13 10 0 9 0 16 15 13 16 9 13 10 0 9 7 10 0 9 7 3 13 0 14 13 1 10 1 10 9 2
32 15 13 3 10 9 15 4 13 1 9 1 15 0 0 9 13 11 1 11 2 10 13 10 9 1 10 9 1 10 0 9 2
15 15 13 1 10 9 1 10 9 7 15 9 13 15 9 2
14 15 4 13 14 3 13 10 1 15 14 13 15 9 2
20 15 13 9 1 9 2 7 1 15 9 15 13 9 1 9 1 9 1 9 2
23 15 4 4 13 14 13 2 7 3 15 4 13 3 1 10 13 15 9 9 7 13 15 2
12 15 4 4 13 1 0 9 1 10 0 9 2
23 15 4 13 14 13 15 13 15 1 10 9 7 15 4 13 10 9 1 15 2 3 3 2
18 16 15 13 15 1 15 9 2 15 4 13 15 3 1 15 11 9 2
15 15 13 15 9 1 10 1 15 1 0 9 2 7 9 2
11 13 7 13 6 2 15 4 4 3 13 2
18 15 4 3 13 1 10 0 9 2 3 15 4 13 3 1 10 9 2
11 15 4 13 3 15 13 3 7 13 3 2
13 15 13 10 0 9 2 7 3 2 9 1 9 2
1 11
16 0 9 2 9 2 9 2 9 2 9 2 9 2 8 8 2
4 15 13 3 2
14 13 15 7 14 2 1 9 7 9 2 15 13 3 2
4 15 13 15 2
26 15 13 10 0 7 0 2 10 9 2 13 2 10 13 9 2 9 7 9 9 2 10 0 7 0 2
11 15 13 10 9 1 9 2 0 7 0 2
13 15 13 7 4 13 9 1 15 0 2 9 3 2
16 15 13 9 2 0 2 0 2 1 0 9 7 13 0 9 2
14 15 13 10 9 16 15 4 13 10 0 9 1 15 2
5 7 15 13 15 2
11 15 15 13 10 0 9 1 0 1 9 2
19 15 15 13 16 9 4 13 1 9 7 9 9 16 15 13 10 9 9 2
44 9 2 0 9 2 0 9 2 9 2 9 2 9 2 10 9 4 13 1 10 9 2 0 9 2 0 9 2 13 10 9 2 0 9 2 9 9 2 9 9 2 9 9 2
9 7 15 13 15 14 13 1 15 2
25 9 13 0 16 10 10 9 13 15 2 1 1 10 9 2 2 10 9 2 10 9 2 10 9 2
9 6 13 15 15 13 10 0 9 2
5 4 15 13 0 2
3 3 0 2
19 3 1 10 0 9 1 10 13 9 1 9 2 15 4 13 15 7 15 2
11 4 15 13 1 10 0 9 7 13 9 2
24 1 10 9 2 4 15 13 10 11 1 11 7 11 11 2 7 4 15 3 13 10 0 9 2
8 15 13 3 9 15 13 3 2
33 6 13 16 15 13 3 14 13 10 9 15 13 15 9 14 13 10 9 2 10 9 2 10 9 2 10 9 2 7 10 0 9 2
22 0 1 15 3 13 9 1 15 3 3 0 1 10 0 9 2 9 7 9 2 9 2
11 0 1 15 13 16 13 9 7 13 9 2
43 0 1 15 4 13 1 10 9 14 13 10 0 9 1 9 2 10 0 9 3 3 3 0 1 15 15 13 1 2 7 0 1 15 4 14 13 16 15 13 10 0 9 2
24 4 15 13 16 3 12 12 11 13 7 13 2 1 9 2 1 9 7 3 13 1 10 9 2
25 10 1 10 12 12 13 9 2 9 2 9 2 7 3 3 7 3 4 10 9 13 1 10 9 2
10 4 14 15 13 15 13 9 15 13 2
4 13 15 0 2
17 4 15 13 16 10 9 15 4 13 13 1 10 0 7 0 9 2
18 4 15 13 10 9 14 13 0 9 16 3 13 16 3 15 13 3 2
23 15 13 16 10 1 15 13 2 7 16 10 1 15 13 2 7 15 13 15 13 15 9 2
11 15 13 15 9 3 16 15 13 15 9 2
23 15 13 3 3 2 3 3 10 0 9 2 10 0 9 1 15 9 2 13 3 14 13 2
3 1 9 2
14 11 11 2 1 11 2 9 9 12 11 2 11 12 11
17 9 2 15 4 13 14 13 10 0 9 9 9 14 13 10 9 2
4 9 13 0 2
4 9 4 13 2
29 10 13 9 1 10 9 2 13 10 9 1 11 11 1 2 10 11 11 2 9 12 9 12 2 9 12 5 12 2
2 2 2
40 9 2 3 4 15 13 10 0 9 14 13 10 2 0 2 9 9 13 1 15 9 10 4 13 9 1 10 9 1 9 2 2 3 2 9 2 9 2 8 2
15 15 13 10 9 1 9 0 1 10 9 1 10 9 9 2
22 16 9 1 1 15 4 14 13 15 15 13 2 13 15 0 9 9 2 7 10 9 2
19 9 1 9 9 2 7 9 1 9 9 9 4 13 3 1 9 7 9 2
2 2 2
14 9 2 15 13 2 9 1 10 11 9 2 9 2 2
26 15 13 1 10 13 9 1 10 11 9 1 10 11 11 11 2 7 3 0 9 9 2 1 0 9 2
11 10 2 9 2 4 13 14 13 10 1 15
8 9 2 2 11 2 2 8 2
3 9 2 9
6 9 2 0 9 13 2
7 3 0 0 9 2 1 11
11 1 2 11 11 11 12 2 12 9 2 12
5 0 9 2 9 2
34 15 13 11 11 11 2 9 1 10 0 11 1 10 11 11 1 11 11 11 11 11 2 7 3 13 1 11 1 10 11 11 1 11 2
17 10 9 4 13 15 16 15 4 14 13 7 1 9 7 1 9 2
40 15 13 14 13 1 15 1 15 9 1 10 0 7 0 9 14 13 10 3 0 9 9 2 10 13 10 9 1 10 0 9 1 9 1 10 9 13 0 9 2
26 15 4 13 15 1 0 9 3 14 13 15 9 16 13 9 9 10 4 3 13 1 10 9 1 11 2
49 15 9 7 15 13 15 9 16 13 10 9 13 1 15 9 2 15 4 3 4 3 13 1 10 9 1 9 1 10 11 11 1 11 2 7 3 13 15 9 1 9 1 10 11 11 11 11 11 2
52 1 10 9 1 10 12 2 9 2 15 9 2 3 9 2 9 1 10 11 11 1 11 2 13 14 13 1 10 0 9 1 10 11 1 10 11 1 11 14 13 13 9 9 9 1 10 13 11 11 1 11 2
40 10 0 9 4 3 13 1 10 9 2 9 1 15 0 9 2 15 13 14 13 0 9 9 9 1 10 13 9 1 11 2 10 3 2 13 11 2 0 9 2
25 15 9 13 10 9 9 1 11 1 12 1 10 9 1 12 2 12 12 11 9 2 5 12 2 2
44 1 1 10 9 2 12 2 12 12 9 2 5 12 2 4 13 1 11 11 2 11 1 11 11 7 0 11 11 9 2 7 12 12 9 2 5 12 2 1 0 7 0 9 2
21 7 15 9 14 0 0 9 9 13 1 9 1 10 11 1 11 7 15 9 9 2
40 15 9 4 13 1 15 0 9 16 13 10 9 1 10 11 1 10 11 1 11 7 13 10 9 9 1 15 9 2 1 9 1 10 9 16 13 15 1 9 2
54 3 2 15 9 1 12 13 14 0 14 13 10 9 1 10 0 9 2 10 1 15 0 9 4 13 10 9 1 12 12 1 12 12 9 2 5 12 5 5 12 2 2 7 1 10 0 9 7 1 0 2 9 9 2
22 1 10 9 1 15 12 9 2 15 4 14 13 0 14 13 10 9 9 13 1 11 2
15 15 13 3 15 9 7 15 9 4 3 13 15 0 9 2
62 15 0 9 1 10 9 9 13 10 13 9 1 10 11 11 1 11 2 11 11 2 15 13 10 0 9 1 10 11 9 7 0 9 1 10 11 9 9 2 7 11 11 2 15 0 9 1 10 9 4 13 1 10 9 1 10 11 9 9 1 15 2
35 15 4 13 15 14 13 10 9 13 12 1 12 2 12 9 2 12 5 12 5 2 1 15 0 9 1 15 9 14 13 1 10 0 9 2
17 10 11 11 11 1 10 11 11 1 11 4 13 1 15 13 9 2
19 15 13 16 15 13 10 9 1 10 9 2 9 2 1 10 9 1 11 2
15 15 13 16 10 9 1 10 9 4 13 9 0 7 0 2
17 7 15 4 13 15 16 10 4 13 0 1 10 9 1 10 9 2
13 10 0 9 13 4 14 4 13 2 15 13 15 2
13 6 4 4 13 16 10 9 9 13 12 5 0 2
22 16 15 4 14 13 14 13 1 10 9 2 6 13 15 0 9 14 3 13 10 9 2
8 15 13 16 15 13 15 9 2
10 15 9 7 15 9 4 13 3 0 2
11 6 13 1 0 9 1 10 9 9 3 2
5 3 1 0 9 2
15 11 11 11 9 2 12 9 2 12 9 2 12 9 2 8
6 11 13 14 13 9 9
3 13 10 9
26 9 9 1 10 0 11 4 13 14 13 9 1 11 11 2 10 3 0 9 14 13 10 9 1 9 2
20 9 1 9 4 13 0 1 11 2 7 10 11 9 1 11 11 4 3 13 2
12 10 9 9 13 9 13 0 14 13 10 0 2
12 2 15 4 3 13 15 3 2 2 15 13 2
20 1 13 9 2 9 13 14 13 10 11 11 9 3 1 1 12 9 13 9 2
12 10 11 9 13 1 9 2 7 9 4 13 2
5 9 1 0 11 11
17 2 15 13 10 3 2 3 0 9 2 2 11 11 11 11 13 2
9 2 10 9 13 16 13 10 9 2
15 12 9 1 11 11 13 13 1 10 9 13 2 9 2 2
10 2 15 4 13 2 13 2 13 9 2
15 15 13 0 9 2 2 11 11 13 10 11 11 9 9 2
34 15 13 14 13 15 9 1 10 9 1 15 9 9 16 9 9 13 1 10 9 1 10 10 12 9 2 0 1 10 13 1 9 9 2
1 9
36 9 13 9 1 1 10 9 2 0 9 4 4 13 2 7 9 9 4 13 9 14 13 12 9 2 12 9 2 9 7 9 9 1 10 9 2
33 16 10 9 13 2 15 4 13 2 15 9 1 11 2 4 13 15 9 2 9 2 12 9 9 7 0 9 7 15 4 13 3 9
5 11 11 11 2 11
3 15 11 9
2 13 11
29 11 11 9 11 11 13 1 1 12 5 1 10 9 4 13 2 1 10 9 1 9 12 9 2 12 9 2 0 2
8 15 13 9 9 4 3 13 2
28 2 10 9 1 10 9 10 13 0 3 4 13 12 7 12 9 2 10 12 9 2 1 9 2 2 15 13 2
38 10 11 11 11 1 11 13 15 4 13 10 9 14 13 10 9 9 2 7 10 9 14 9 9 9 4 13 9 3 14 13 14 13 3 1 15 9 2
18 10 11 14 11 11 1 11 11 13 15 13 9 16 0 9 13 1 2
19 3 0 9 4 4 13 14 13 10 9 1 0 9 14 13 9 1 9 2
18 16 10 9 4 13 0 9 2 9 4 3 13 14 13 9 7 9 2
4 2 9 0 2
10 10 9 13 14 13 3 0 1 11 2
20 2 15 4 13 14 4 13 1 9 0 1 10 9 2 2 10 9 9 13 2
9 2 10 9 13 16 13 10 9 2
13 9 13 1 9 4 4 13 1 10 9 7 3 2
18 9 1 9 13 0 2 7 9 13 15 4 13 9 16 9 4 13 2
30 2 15 4 3 13 16 15 13 15 11 13 1 12 9 3 2 2 13 11 11 11 11 16 13 10 9 1 10 9 2
16 9 4 4 13 10 10 9 2 13 12 9 15 13 15 9 2
21 11 11 1 11 13 10 9 1 11 11 16 15 13 1 11 7 11 16 13 3 2
11 11 9 3 13 12 9 13 1 10 9 2
29 1 11 2 12 9 4 13 0 1 12 9 1 9 10 4 13 1 10 12 9 2 12 9 2 2 9 9 2 2
19 10 9 14 9 9 4 13 2 1 10 9 2 2 0 9 11 11 13 2
1 9
21 11 14 11 11 13 9 14 13 11 1 9 7 13 15 10 9 4 3 4 13 2
4 13 11 14 9
28 10 11 11 11 4 13 9 1 9 1 15 0 2 3 0 9 9 7 0 9 9 4 4 13 1 13 9 2
28 11 11 11 11 2 15 4 13 15 9 12 9 0 2 4 13 1 11 14 13 1 10 11 11 7 0 9 2
23 9 9 1 0 1 5 12 12 13 15 4 13 10 11 9 9 14 3 0 0 9 3 2
31 10 9 1 0 9 1 10 0 9 13 10 0 5 12 10 9 1 1 10 9 1 9 7 9 9 1 10 11 1 11 2
16 10 11 9 9 4 13 16 9 4 4 13 1 9 9 9 2
4 13 1 10 9
15 9 9 9 2 9 2 9 7 9 2 9 13 1 9 9
7 9 2 11 13 10 9 2
6 2 13 2 12 9 2
1 9
7 9 2 11 13 10 9 2
5 9 2 9 2 9
6 13 1 2 11 2 11
5 9 9 2 5 12
7 13 2 12 11 12 12 9
7 13 2 12 11 12 12 9
4 9 9 2 12
11 3 0 9 4 10 11 13 11 1 9 2
1 9
9 9 2 1 2 11 13 10 9 2
12 13 1 2 11 2 11 1 12 11 12 12 9
5 6 11 2 11 2
24 1 11 12 2 12 2 10 11 11 11 11 13 5 12 12 1 9 1 11 1 0 9 12 2
16 15 13 10 5 12 12 9 16 15 11 13 1 0 9 12 2
5 11 11 11 1 11
2 9 9
4 11 12 2 12
41 2 11 11 7 11 11 2 11 2 2 4 13 1 5 12 12 2 10 9 1 5 12 12 1 10 9 13 9 2 7 10 9 1 5 12 12 1 10 9 9 2
21 10 0 5 12 12 1 9 9 4 13 1 11 1 10 9 14 9 1 10 9 2
24 2 10 9 1 9 9 1 10 9 9 4 13 1 5 12 12 2 10 13 9 1 10 9 2
12 2 10 11 11 11 4 13 1 5 12 12 2
25 10 9 13 11 9 1 5 12 12 1 1 10 13 13 9 1 10 11 1 3 3 9 1 9 2
7 2 10 11 2 11 9 2
15 2 10 11 11 11 2 11 2 4 13 1 5 12 12 2
12 2 10 0 9 9 4 13 1 5 12 12 2
10 2 5 12 12 4 13 1 11 11 2
24 11 11 11 2 11 2 2 4 13 1 5 12 12 2 10 0 1 9 7 10 9 9 2 2
1 8
4 11 13 11 13
29 2 10 11 11 11 13 10 3 0 9 11 14 13 11 14 0 9 12 9 1 5 12 12 16 15 11 11 13 2
37 10 9 13 14 13 11 5 12 12 1 12 2 3 5 12 12 0 16 15 10 11 13 7 3 5 12 12 0 16 15 11 9 13 1 11 2 2
9 15 13 15 4 13 10 9 0 2
15 16 15 13 10 9 2 6 13 9 0 16 13 10 9 2
1 11
4 11 9 9 2
2 11 9
7 9 13 1 14 13 10 9
9 9 2 1 2 11 13 10 9 2
11 1 2 11 2 11 1 12 11 12 12 9
4 0 9 11 2
7 13 15 13 10 0 9 2
14 15 4 13 9 1 11 9 3 2 1 15 0 9 2
19 3 2 1 15 0 9 2 9 3 11 13 0 2 1 10 0 9 9 2
28 15 13 16 15 13 9 3 0 16 3 11 13 15 9 15 4 13 3 12 4 13 10 9 1 11 2 11 2
60 13 15 13 15 10 9 2 16 15 4 13 11 3 2 13 10 0 9 2 13 1 10 9 2 13 10 9 1 0 9 2 13 10 9 2 13 10 9 2 13 10 0 9 2 8 3 15 4 3 3 13 10 9 10 11 4 13 1 15 2
17 3 11 13 10 0 9 9 1 9 2 10 9 13 15 13 0 2
4 0 2 11 2
20 9 2 1 2 11 13 10 9 2 1 2 11 2 11 1 12 11 12 12 9
37 15 13 16 11 13 10 0 9 1 9 9 14 9 2 7 15 13 3 0 0 9 1 9 9 9 2 16 15 13 15 0 3 14 13 1 15 2
29 15 3 13 10 11 11 1 10 11 13 10 9 2 7 15 13 15 4 3 13 15 9 13 1 10 11 1 11 2
37 3 3 2 1 10 0 9 2 9 9 14 9 4 13 1 10 9 1 0 9 9 2 7 9 1 10 0 2 7 15 13 0 1 10 0 9 2
29 1 9 1 11 14 9 2 4 15 3 13 16 13 9 1 9 9 1 10 9 13 10 0 9 14 13 10 9 2
3 7 9 2
8 15 13 15 3 0 14 13 2
26 15 13 15 4 4 4 13 1 10 3 3 9 0 9 2 3 3 1 0 2 0 2 9 2 11 2
5 3 15 12 9 2
4 9 16 13 2
8 6 13 10 9 14 13 15 2
28 15 13 16 15 4 13 0 2 7 15 13 0 1 15 9 7 13 0 14 13 9 14 13 15 0 0 9 2
15 15 13 3 9 2 7 4 13 3 12 9 1 15 9 2
15 15 13 14 10 9 2 16 3 0 1 10 9 3 13 2
28 1 0 9 2 11 11 2 10 0 9 1 15 9 2 4 13 10 9 1 10 9 9 15 9 4 13 1 2
36 10 9 13 0 1 10 0 9 10 13 10 5 12 0 9 2 10 15 4 13 14 13 1 9 14 13 15 1 10 9 9 10 15 4 13 2
14 3 13 10 9 1 9 13 10 0 0 1 10 9 2
22 15 15 4 13 14 13 13 13 9 1 10 9 2 1 9 14 13 15 1 0 9 2
24 15 13 3 1 0 9 2 7 13 15 9 16 16 10 9 9 4 4 13 1 10 0 9 2
16 15 4 13 1 10 13 9 2 15 4 3 13 10 0 9 2
18 6 13 10 9 14 13 1 10 9 3 7 13 15 9 1 11 11 2
11 13 15 1 9 1 15 9 1 10 9 2
18 3 2 6 13 15 3 1 9 15 13 2 7 10 1 15 9 9 2
12 15 13 10 9 1 10 9 14 13 15 1 2
4 10 9 9 13
15 15 4 13 10 9 1 10 1 15 1 10 11 11 9 2
4 10 9 13 2
21 10 9 9 1 11 1 10 11 13 2 7 15 13 10 10 9 13 1 10 9 2
22 15 4 13 15 1 3 3 2 14 13 16 15 13 3 0 2 7 1 10 0 9 2
38 11 13 15 0 9 2 7 15 4 13 14 13 9 1 15 10 9 15 4 2 3 10 9 9 13 0 14 13 15 13 14 13 15 9 2 13 9 2
14 0 9 2 7 4 11 13 15 10 7 13 15 0 2
28 3 13 10 9 15 4 13 2 1 1 10 9 1 10 9 9 9 15 4 13 1 11 2 3 1 15 9 2
2 11 2
24 15 4 13 15 10 9 10 15 4 13 3 13 10 9 14 13 10 9 1 10 9 9 9 2
32 16 15 4 13 10 9 3 2 7 13 9 15 13 14 13 15 1 15 9 2 8 2 15 4 13 10 9 16 13 15 1 2
2 9 2
1 11
2 11 2
12 15 4 13 10 9 13 10 9 15 4 13 2
9 15 13 10 9 1 10 9 9 2
10 10 9 16 13 15 4 4 3 13 2
8 15 13 3 1 10 0 9 2
25 11 13 14 13 1 11 11 3 10 9 1 10 9 2 7 15 9 1 10 0 9 9 4 13 2
22 15 4 14 13 10 9 14 13 1 10 9 2 7 1 10 9 2 15 9 13 0 2
8 15 13 15 13 10 0 9 2
26 3 13 15 9 14 13 15 3 1 15 9 2 7 3 3 2 16 16 10 9 14 13 15 13 3 2
18 15 4 13 1 0 9 1 9 14 13 10 5 12 1 10 9 9 2
12 13 15 3 3 16 13 3 14 13 15 9 2
1 11
7 9 9 7 9 1 11 11
12 3 2 11 12 2 12 2 12 9 1 12 9
5 3 2 11 11 11
6 9 2 9 1 10 9
17 11 11 13 15 0 9 15 13 0 9 2 7 15 13 15 9 2
26 15 9 1 10 9 13 9 15 13 4 13 1 2 7 15 13 14 13 15 14 13 14 13 10 9 2
16 11 13 12 0 0 9 2 7 9 15 13 15 7 13 15 2
10 6 13 15 14 13 15 13 10 9 2
11 1 15 9 2 15 13 15 4 13 15 2
19 15 4 13 12 9 2 7 11 11 4 13 2 9 1 9 7 0 9 2
11 15 13 10 9 15 4 14 13 14 13 2
35 9 2 9 2 7 9 4 13 1 11 11 2 15 4 4 13 1 10 11 1 10 11 11 1 10 11 11 11 1 11 11 1 11 12 2
27 10 9 1 10 9 4 13 5 12 2 10 11 11 13 14 13 1 9 14 13 15 1 10 11 11 9 2
14 6 13 15 16 13 1 10 11 1 10 11 9 1 2
19 13 10 9 1 11 11 2 7 13 15 13 11 1 15 9 13 9 3 2
10 9 4 3 4 13 1 11 11 11 2
13 13 9 0 1 11 11 9 2 1 11 1 11 11
3 1 11 11
5 2 13 2 12 2
33 11 14 0 9 1 9 4 13 9 1 0 7 0 9 1 10 9 16 15 13 0 9 1 9 1 3 3 3 1 11 7 11 2
32 10 9 1 0 0 9 1 10 0 0 9 0 9 7 10 9 9 1 11 13 10 0 3 0 9 1 11 14 13 0 9 2
12 13 9 9 1 11 4 13 10 0 9 1 9
39 10 9 2 3 2 13 1 10 9 13 0 9 1 11 11 11 14 13 0 9 9 3 2 3 9 10 4 14 4 13 1 11 1 9 1 9 1 11 2
22 10 9 9 4 13 1 1 10 2 0 9 2 1 10 0 9 2 10 13 1 11 2
47 7 3 1 10 9 10 11 14 11 2 10 9 9 2 4 13 16 9 1 10 11 11 11 1 10 12 9 13 2 3 10 9 1 10 9 1 11 7 11 1 10 9 1 0 9 2 2
37 10 11 9 9 13 9 1 10 0 9 2 9 7 9 9 1 10 9 10 9 13 4 13 1 1 12 9 10 9 16 3 13 9 1 10 9 2
13 10 9 2 3 2 4 13 0 9 1 10 9 2
26 7 10 11 11 7 11 13 3 3 0 1 10 3 3 0 9 1 11 14 9 1 2 9 9 2 2
20 1 11 2 11 13 14 13 10 9 14 13 9 1 11 1 10 9 1 11 2
25 15 4 13 5 12 12 1 10 0 9 14 9 9 2 10 13 15 1 12 9 9 1 15 9 2
32 3 2 10 9 2 15 13 16 15 13 9 14 13 11 14 0 9 2 9 1 10 11 11 11 11 1 10 11 11 11 11 2
38 10 9 3 2 11 14 3 0 9 9 9 4 13 10 5 12 12 9 1 9 7 0 9 9 1 11 2 10 3 13 12 9 9 1 11 14 9 2
18 11 13 15 0 9 1 9 7 0 9 7 3 13 10 0 9 9 2
28 7 16 15 9 4 13 1 10 9 1 12 9 9 1 9 1 10 0 12 9 2 3 13 15 9 1 9 2
19 10 9 15 13 11 1 10 9 14 3 0 9 1 9 2 1 10 11 2
40 15 13 9 2 13 1 10 0 9 1 9 9 3 3 1 10 9 14 13 9 1 13 9 1 9 9 2 4 13 1 10 9 1 10 9 1 9 10 9 2
12 9 4 3 13 1 9 9 1 10 0 9 2
42 16 11 11 13 9 2 13 9 9 14 2 13 3 2 14 13 9 2 15 4 13 13 1 9 1 10 11 11 11 2 3 3 1 10 9 10 11 13 1 15 9 2
16 11 13 2 1 10 9 2 16 10 9 4 13 10 0 9 2
13 10 12 13 3 0 14 13 1 11 14 9 9 2
28 11 13 0 16 11 4 13 15 1 15 9 14 13 10 9 1 10 9 10 11 13 14 13 1 10 11 11 2
19 11 13 10 9 1 10 9 2 13 9 14 4 13 1 7 11 7 11 2
21 11 13 10 0 9 1 15 0 9 2 10 4 13 15 0 9 16 9 13 1 2
22 3 2 9 4 13 16 11 14 9 4 13 16 15 13 0 7 3 1 15 0 9 2
28 11 11 2 10 0 9 1 10 11 11 11 1 11 2 13 10 9 1 10 11 11 11 13 3 0 10 9 2
24 2 9 13 16 15 4 13 10 9 1 9 7 9 1 10 9 1 10 9 2 2 15 13 2
20 2 15 4 13 10 0 0 9 7 15 4 14 13 10 9 9 13 0 2 2
49 11 11 2 10 11 11 2 13 9 1 0 9 2 13 15 9 9 13 1 16 11 4 13 10 10 13 9 1 15 9 1 11 16 10 9 1 10 9 15 13 1 1 13 12 9 10 9 9 2
48 2 16 11 14 9 13 2 10 2 1 15 9 2 13 3 0 2 3 9 9 4 13 2 7 1 15 2 10 9 1 10 9 10 13 15 2 2 11 11 2 11 14 0 11 9 2 13 2
33 2 11 4 13 1 1 10 0 9 11 9 2 3 15 4 13 14 13 3 13 0 9 1 10 9 16 15 15 13 1 15 2 2
22 11 14 0 9 14 13 9 7 9 13 10 0 9 1 15 0 9 1 10 0 9 2
11 2 11 13 10 0 9 2 2 15 13 2
40 2 15 13 10 0 9 1 0 9 3 11 4 13 14 13 15 9 9 1 10 11 11 11 1 10 9 13 1 10 11 11 7 13 1 11 7 11 11 2 2
3 9 2 8
6 9 1 10 0 13 9
1 2
34 16 15 13 16 15 3 13 10 9 1 0 9 14 13 10 9 13 10 9 1 9 2 13 10 13 16 13 1 10 3 0 9 3 2
14 9 4 13 1 0 9 2 7 9 13 0 1 15 2
10 9 13 14 13 16 15 4 13 9 2
28 15 13 3 0 14 13 1 10 0 0 9 9 1 10 9 1 9 13 1 10 9 9 10 13 1 10 9 2
14 13 10 0 9 1 10 9 7 13 1 15 9 13 2
29 13 15 9 12 1 9 1 10 0 1 15 9 2 13 15 9 0 2 9 13 7 9 1 10 9 1 15 9 2
12 15 9 4 13 0 7 0 2 1 10 9 2
18 13 10 9 7 3 13 1 15 9 2 13 10 9 13 1 15 9 2
5 8 2 0 9 9
7 13 14 13 3 7 3 2
38 1 10 9 2 13 10 9 1 15 9 13 0 7 0 2 7 3 15 0 9 7 0 9 4 13 16 15 4 13 1 10 9 1 10 0 0 9 2
13 13 10 9 13 3 16 15 13 13 3 7 3 2
18 13 15 13 1 10 0 2 0 9 13 1 10 9 1 10 9 2 2
28 13 10 0 2 0 9 1 10 9 2 15 9 7 9 2 2 10 9 1 1 15 2 7 10 9 1 15 2
9 13 15 13 1 10 9 7 9 2
24 16 15 13 1 10 9 2 10 9 1 10 0 9 13 15 9 7 13 15 13 0 7 0 2
4 15 13 15 2
8 10 0 9 13 0 7 0 2
11 3 15 13 3 1 10 9 2 1 9 2
7 9 1 15 13 3 0 2
12 7 2 15 13 9 7 10 9 1 10 9 2
15 15 13 14 13 15 9 1 10 0 0 9 10 13 15 2
18 13 14 13 1 10 0 9 16 15 9 14 13 1 10 10 0 9 2
24 7 16 13 3 13 13 10 9 9 9 9 2 13 3 1 9 9 2 13 3 1 9 2 2
8 13 15 1 12 1 12 9 2
9 3 13 3 1 11 3 2 3 2
10 13 15 13 1 10 9 3 7 3 2
7 15 9 13 0 7 0 2
14 13 15 9 13 3 1 10 9 13 10 0 9 3 2
14 10 9 14 9 7 9 13 3 1 15 2 13 15 2
10 15 13 1 10 9 1 9 7 9 2
17 1 10 9 2 13 15 9 7 13 16 15 13 0 2 1 9 2
19 13 14 13 10 9 1 10 9 3 1 15 9 2 13 15 3 7 3 2
24 15 13 14 13 9 3 1 15 1 15 0 9 9 3 15 13 15 9 13 1 10 0 9 2
21 15 4 13 10 9 1 10 9 2 10 0 9 7 9 1 9 7 10 0 9 2
23 13 10 9 1 15 9 13 1 10 0 9 2 13 10 9 7 13 3 3 1 10 9 2
15 10 0 2 0 9 13 1 15 9 7 13 15 3 3 2
10 13 15 9 7 9 13 3 1 9 2
20 3 13 15 13 16 3 15 13 2 13 15 9 7 9 10 0 2 13 15 2
4 13 15 9 2
4 8 2 9 9
6 10 9 15 4 13 2
23 13 15 4 13 1 9 1 10 9 2 7 16 15 13 10 3 0 9 15 4 13 1 2
17 13 16 15 4 13 3 1 0 9 2 3 1 9 1 10 9 2
12 3 13 16 0 9 4 13 15 1 10 9 2
12 13 15 4 3 13 1 10 0 9 7 9 2
14 3 13 14 13 1 15 9 10 9 2 9 9 9 2
10 15 9 13 2 0 9 13 3 2 2
34 13 10 9 2 4 14 3 13 1 15 0 9 7 13 14 13 1 11 2 9 9 9 2 1 10 0 9 2 0 9 7 9 2 2
19 13 3 2 3 2 3 1 9 2 1 10 9 2 16 15 4 13 15 2
5 15 4 13 9 2
14 15 13 0 14 13 10 9 2 3 3 10 0 9 2
16 13 3 1 10 9 13 15 13 9 2 15 13 10 0 9 2
19 3 2 13 14 13 7 13 1 0 9 13 10 0 9 2 10 0 9 2
32 13 15 4 13 1 0 9 7 9 2 7 13 16 15 0 9 1 9 13 1 0 9 1 10 0 9 7 9 3 1 15 2
23 15 4 13 3 7 13 16 15 9 9 2 10 9 1 10 0 9 2 4 13 1 9 2
13 13 1 3 3 16 15 13 2 3 13 15 9 2
7 6 15 13 3 0 5 2
20 10 0 9 13 14 13 10 0 9 1 15 9 7 10 0 9 7 0 9 2
18 4 14 13 16 15 13 9 13 1 10 9 7 9 2 15 13 0 2
16 15 13 10 9 7 9 14 13 0 14 13 1 10 12 9 2
8 10 0 9 13 14 13 13 2
10 16 15 4 14 13 2 3 9 13 2
25 6 3 10 9 4 13 2 7 13 15 13 15 15 13 0 9 7 3 13 0 9 1 9 9 2
1 2
7 11 11 11 11 1 11 11
22 16 15 15 13 1 10 9 9 2 12 4 3 13 16 10 11 13 0 1 0 9 2
7 7 15 13 14 10 9 2
45 0 9 10 9 13 10 11 11 11 11 1 11 11 4 13 14 13 3 10 9 16 3 3 10 9 1 9 13 14 0 16 13 10 9 7 9 1 0 9 1 0 2 9 9 2
37 12 1 2 11 14 2 0 9 13 14 13 9 1 10 13 2 9 1 0 9 2 2 10 4 13 7 4 3 13 13 1 9 1 10 11 9 2
47 15 13 10 9 1 9 9 7 13 2 2 15 4 13 16 10 11 4 14 13 1 0 2 9 9 15 13 14 13 7 13 3 7 3 1 10 9 2 9 2 7 9 1 0 9 2 2
49 10 9 14 13 10 11 9 14 13 0 9 4 13 0 9 7 3 4 4 13 1 10 12 0 9 2 3 15 13 10 0 9 1 0 9 1 10 2 0 2 9 2 9 2 9 1 10 9 2
17 1 15 11 9 10 11 11 13 3 14 13 15 9 1 10 9 2
13 15 9 11 7 15 9 11 3 4 13 10 9 2
20 3 2 10 11 13 3 14 13 10 9 1 9 1 10 11 9 1 10 9 2
41 2 16 10 9 4 13 16 13 1 2 0 9 2 2 9 15 4 14 13 15 2 0 9 2 4 13 1 2 9 1 10 11 11 11 11 1 11 11 2 2 2
21 6 13 16 10 9 13 3 0 9 2 15 13 9 1 0 9 7 9 13 9 2
26 16 15 13 10 9 6 13 0 14 13 15 2 1 11 10 9 2 3 15 4 13 1 10 9 2 2
23 13 2 1 9 4 13 0 1 10 9 1 11 12 7 11 12 2 7 15 4 13 15 2
30 15 4 13 9 7 9 9 2 7 0 9 2 1 9 1 11 1 9 1 15 2 9 9 2 1 11 1 11 12 2
9 13 15 1 15 9 1 10 9 2
9 1 10 11 1 10 11 11 11 2
4 11 11 12 8
1 2
15 11 11 11 11 1 11 11 9 1 0 9 11 12 2 12
30 10 3 0 0 9 2 1 10 9 1 9 2 9 7 9 2 13 10 9 1 9 7 10 0 9 1 0 0 9 2
11 15 13 3 3 0 3 15 13 10 9 2
19 15 4 13 1 15 9 14 13 0 2 14 13 0 2 1 10 9 9 2
37 10 9 14 13 7 13 10 9 13 3 0 16 15 11 11 11 13 15 1 13 1 15 9 14 2 13 10 9 1 9 1 15 7 15 9 2 2
37 10 11 11 11 3 13 10 2 0 9 2 1 0 9 1 2 9 2 9 2 10 9 1 10 9 1 15 0 9 2 7 10 9 1 9 2 2
29 1 9 2 9 4 13 16 16 13 10 9 1 13 9 14 13 7 13 9 2 15 4 13 10 9 1 10 9 2
28 5 1 10 0 9 1 9 1 11 2 10 9 16 13 9 14 13 13 0 1 10 9 1 10 0 0 9 2
15 10 0 9 13 0 9 2 3 13 1 2 13 3 0 2
23 9 1 10 9 1 9 1 15 15 4 3 13 15 9 13 0 7 0 9 7 0 9 2
10 15 13 13 14 13 7 13 10 9 2
24 1 0 9 2 9 7 0 9 2 15 4 13 1 9 14 13 1 9 1 15 0 0 9 2
20 15 13 10 9 1 0 9 7 0 9 14 13 0 9 1 0 2 9 9 2
18 1 0 9 15 13 10 9 1 9 1 10 0 9 14 13 7 13 2
49 15 13 16 10 9 2 3 10 9 2 4 13 14 13 9 1 9 7 13 12 13 9 2 16 1 10 0 7 13 9 2 16 13 10 9 9 10 13 15 13 3 3 0 2 3 3 3 0 2
26 15 13 10 9 16 9 7 9 13 1 0 1 15 0 9 1 1 10 0 2 0 7 0 9 13 2
16 3 2 15 13 1 15 0 9 9 14 13 1 10 0 9 2
35 15 4 13 16 10 9 4 14 13 1 0 2 9 9 15 13 14 13 7 13 3 7 3 1 10 9 2 9 2 7 9 1 0 9 2
9 15 13 9 1 9 1 10 9 2
22 15 13 16 10 9 4 14 13 0 9 14 13 1 2 7 13 2 0 2 9 9 2
29 3 2 10 9 1 9 0 9 13 10 0 9 1 10 9 7 9 15 13 1 2 7 13 2 0 2 9 9 2
31 10 9 4 14 13 10 9 1 12 0 9 1 10 16 13 9 15 0 9 14 13 7 14 13 10 9 13 1 0 9 2
29 1 9 9 2 15 13 15 1 0 9 2 9 2 9 2 7 0 9 1 10 9 1 10 9 7 9 14 13 2
1 2
7 11 11 11 11 2 11 12
7 9 2 11 11 2 8 2
13 10 12 9 3 10 11 4 13 10 9 1 11 11
19 15 4 13 1 15 9 1 9 7 9 2 13 3 3 0 9 1 10 11
4 15 0 11 2
48 16 0 1 15 4 4 13 2 11 11 4 13 10 0 2 9 0 9 13 11 11 14 13 10 0 9 1 10 11 11 11 11 2 14 13 10 9 13 1 10 9 1 10 9 1 10 9 2
33 1 15 9 2 10 9 4 14 13 9 16 7 16 10 11 11 11 13 15 9 2 16 13 1 15 9 2 9 12 2 9 12 2
18 10 9 1 10 9 2 1 9 3 1 10 0 9 2 4 13 1 8
21 9 11 11 13 3 3 0 1 10 1 10 0 9 13 14 13 9 1 10 9 2
7 15 13 10 3 0 9 2
18 15 13 3 3 1 15 9 2 1 11 9 7 1 9 9 1 11 2
24 15 13 10 0 7 0 9 2 13 0 9 1 10 0 9 9 2 10 0 9 1 11 11 2
20 15 13 0 9 1 9 1 0 11 11 9 2 7 15 4 13 9 1 9 2
30 15 13 10 0 2 0 9 2 2 13 0 2 0 2 0 2 0 1 10 9 2 0 1 15 9 2 0 1 9 2
5 15 9 13 15 2
6 15 0 9 13 15 2
5 15 9 13 15 2
5 11 11 13 15 2
23 6 2 15 13 0 16 10 9 4 14 13 10 9 15 13 15 4 13 1 10 11 11 2
28 7 0 9 4 13 10 9 15 13 15 4 13 2 7 10 9 15 13 15 13 14 13 10 9 15 13 15 2
47 3 3 10 11 4 13 0 14 13 3 2 16 16 14 13 15 7 14 2 7 1 10 9 2 9 1 11 12 2 12 2 15 13 16 15 13 0 1 10 12 2 12 9 13 1 9 2
38 10 11 13 3 0 14 13 3 3 7 13 10 9 2 16 15 3 3 13 14 13 11 11 1 10 11 11 2 14 4 13 10 9 11 13 0 1 2
21 3 15 13 10 9 1 13 2 1 9 1 10 11 14 13 15 0 9 1 9 2
21 15 13 10 0 9 10 13 1 10 9 2 2 13 1 9 2 13 1 9 2 2
19 3 15 4 13 10 0 9 3 3 2 3 13 15 1 0 9 14 13 2
102 15 13 15 13 0 14 13 1 9 11 11 2 1 15 9 2 16 15 13 12 0 9 2 10 3 0 0 9 1 15 9 2 10 13 15 3 0 1 10 9 1 11 11 9 2 15 4 14 3 13 1 10 9 1 2 9 7 9 2 13 1 10 9 2 7 15 13 0 14 13 13 15 1 1 9 14 13 10 2 11 11 11 2 2 10 13 1 3 2 13 0 9 1 10 9 1 11 7 10 11 11 2
9 7 1 1 10 0 9 2 2 2
22 2 15 4 13 1 15 9 1 9 7 9 2 13 3 3 0 9 1 10 11 2 2
23 1 15 0 9 2 15 13 12 9 1 10 11 11 2 10 0 2 0 2 7 0 9 2
30 7 10 0 9 1 10 9 7 9 15 13 13 16 16 12 9 1 10 9 13 0 2 10 0 12 4 13 15 3 2
99 7 11 11 13 1 10 3 2 13 0 9 2 13 10 2 11 11 11 2 2 10 13 16 10 11 4 13 0 9 1 10 0 9 2 7 16 10 0 9 4 13 1 9 1 3 9 10 10 9 3 13 2 13 10 9 1 10 0 9 10 4 13 14 13 0 1 0 9 2 7 10 9 2 10 13 2 10 4 13 2 7 10 4 13 1 0 9 13 1 10 9 1 11 2 3 1 10 11 2
16 10 9 13 14 9 1 10 0 9 2 15 13 10 0 9 2
57 2 11 1 11 2 4 14 13 16 15 13 10 9 1 10 9 2 3 16 15 13 10 9 2 3 16 15 13 10 9 1 10 0 9 2 13 16 2 13 3 2 10 10 9 13 1 11 7 10 10 9 13 1 10 11 11 2
27 1 10 11 11 11 2 10 9 1 11 7 9 1 10 11 11 13 10 0 9 16 10 11 13 1 15 2
21 7 3 11 7 10 11 11 13 0 9 1 10 11 2 1 10 0 9 1 15 2
30 7 10 11 13 10 9 2 0 1 9 1 10 9 2 13 1 1 10 0 9 2 10 4 13 3 1 15 0 9 2
39 7 3 10 11 11 1 11 2 10 9 1 10 0 7 10 9 1 10 0 2 13 3 10 0 9 2 3 0 1 11 11 7 0 11 1 11 11 12 2
14 7 10 13 3 10 11 4 13 10 9 1 11 11 2
11 1 9 7 0 9 2 6 13 10 9 2
3 9 1 8
5 9 7 9 1 8
4 9 1 15 2
6 4 11 13 15 10 2
6 7 4 11 13 11 2
8 11 11 11 2 9 8 7 8
8 9 1 10 9 4 13 3 2
19 16 15 13 14 13 2 6 13 15 1 9 15 13 15 13 14 13 15 2
3 8 7 8
1 5
20 13 11 11 2 11 11 11 2 12 11 11 11 9 12 11 2 11 12 12 8
1 13
16 11 7 9 9 2 13 14 13 9 9 9 10 9 1 0 9
29 10 9 4 13 1 11 7 9 1 9 1 11 7 0 9 13 9 4 13 3 16 4 13 1 10 9 9 3 2
33 9 13 10 0 9 2 11 7 9 14 13 2 9 9 2 9 2 13 14 13 2 13 2 13 7 13 10 9 9 1 10 9 2
15 15 4 3 13 1 0 2 0 2 0 2 7 0 9 2
33 9 3 0 7 14 13 13 9 2 11 7 9 14 13 2 9 9 2 9 3 3 10 9 13 10 0 2 13 7 0 9 9 2
15 15 4 3 13 1 0 2 0 2 0 2 7 0 9 2
20 0 2 11 7 9 14 13 2 9 9 2 9 14 13 10 9 1 0 9 2
23 15 13 3 10 9 9 9 1 11 7 9 7 3 4 14 13 9 13 10 9 9 9 2
56 10 9 1 11 7 11 3 14 13 1 12 10 10 0 9 9 9 13 1 10 9 2 1 10 9 1 10 9 9 2 3 13 15 7 13 3 1 10 9 9 9 2 13 10 0 9 1 9 9 1 9 9 1 0 9 2
7 11 13 15 0 0 9 9
12 0 9 13 9 1 10 9 1 10 9 14 9
3 1 11 11
4 9 12 11 11
1 11
19 11 13 11 11 2 15 0 0 9 2 3 9 1 0 11 14 11 11 2
29 10 9 1 0 9 13 1 11 14 3 0 9 9 3 9 2 13 1 9 1 10 9 9 10 4 13 12 9 2
28 10 9 1 10 11 11 9 4 13 1 11 11 2 12 2 7 11 11 2 12 2 1 11 14 0 9 9 2
23 10 0 9 1 10 11 11 11 11 1 0 11 13 10 0 9 1 11 11 1 11 12 2
32 15 12 2 9 9 13 15 0 9 1 10 0 9 1 0 9 2 11 7 10 11 11 2 10 4 13 7 13 9 1 9 2
20 0 9 13 11 13 14 13 10 0 9 9 1 15 0 1 10 0 0 9 2
22 7 15 13 0 16 16 11 13 14 13 10 11 11 1 10 9 1 15 0 9 9 2
20 11 11 4 13 11 14 13 1 10 9 1 12 1 10 0 9 1 0 9 2
43 11 14 2 13 14 10 13 2 1 2 9 9 2 2 13 11 11 2 11 2 10 9 1 0 9 15 13 9 9 1 10 0 9 1 10 11 11 11 1 11 2 11 2
8 2 15 13 14 1 10 9 2
16 15 13 10 9 10 4 13 10 9 2 2 11 2 11 13 2
21 2 15 4 14 13 14 13 15 2 16 15 4 14 13 15 14 13 10 9 9 2
14 9 4 13 10 0 9 1 10 9 1 15 9 2 2
54 11 14 9 14 13 10 11 2 13 9 14 13 10 12 2 9 0 9 9 4 4 13 1 0 1 10 9 1 10 9 1 9 2 13 10 0 9 14 0 9 9 7 9 15 4 13 9 10 4 13 10 9 9 2
10 10 9 13 3 1 11 14 12 9 2
42 11 13 1 12 9 13 14 13 10 9 1 11 2 13 9 9 1 11 14 9 14 13 10 9 1 9 1 10 0 9 1 10 9 1 11 7 0 2 0 9 9 2
16 2 15 13 11 14 9 9 2 2 11 9 11 11 13 11 2
12 2 15 13 15 10 0 9 1 15 9 2 2
19 15 13 2 3 2 16 11 4 14 13 10 9 14 0 9 1 0 9 2
36 1 0 2 15 13 10 9 1 0 9 1 0 9 14 13 10 11 9 9 7 14 13 10 9 1 11 14 13 10 9 9 9 2 11 13 2
28 10 9 1 11 7 11 4 13 10 9 1 10 13 9 1 10 12 2 9 0 9 9 2 11 2 11 13 2
31 10 0 9 2 15 13 2 4 13 10 9 1 10 0 9 10 4 13 10 9 9 1 9 3 10 12 9 13 1 11 2
20 10 0 9 14 0 9 4 13 9 1 0 9 7 9 1 9 7 9 9 2
17 10 0 9 4 13 10 9 7 9 1 10 0 2 9 9 9 2
26 3 3 12 9 13 11 14 9 4 13 10 9 9 14 13 10 9 1 9 1 11 14 13 0 9 2
33 2 10 11 4 13 0 14 13 3 2 2 13 11 11 11 2 9 1 10 11 2 11 2 13 8 2 10 0 0 9 9 9 2
26 2 15 13 3 10 9 15 4 13 15 1 2 13 15 13 16 15 13 14 9 9 2 2 11 13 2
32 1 10 11 7 0 0 9 1 10 11 11 2 11 13 10 0 9 16 13 10 9 1 10 11 11 9 1 10 12 11 9 2
14 16 15 13 1 2 10 11 3 13 15 1 10 9 2
17 2 2 11 2 4 13 10 0 9 14 13 15 2 2 11 13 2
12 2 15 4 13 1 9 1 9 1 10 11 2
18 7 15 4 14 13 14 13 1 10 9 14 13 15 3 10 9 2 2
40 11 14 9 13 13 1 11 14 9 1 10 0 0 2 9 9 2 10 11 11 11 2 7 10 9 1 10 0 9 9 9 1 11 11 1 10 11 11 11 2
42 10 12 9 2 15 13 2 4 3 13 11 14 9 9 14 13 1 10 9 3 9 4 13 7 13 1 11 14 9 10 9 0 16 13 10 9 1 9 7 13 3 2
1 8
8 9 2 2 11 2 2 8 2
21 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9
22 15 13 10 9 1 10 0 9 9 9 2 7 13 0 9 1 0 9 7 10 9 2
65 3 2 15 13 10 9 10 13 10 0 9 9 9 13 1 1 0 9 15 13 15 1 9 7 13 10 9 1 10 9 1 1 12 9 1 9 2 16 16 15 4 3 13 10 9 1 1 15 9 7 13 15 1 0 9 15 13 15 14 13 10 9 1 9 2
48 10 9 3 13 2 10 13 16 10 9 13 3 0 2 15 13 3 0 1 15 2 9 2 16 15 4 13 2 3 16 13 10 9 13 1 10 9 2 1 10 9 1 9 2 9 2 9 2
27 3 15 13 10 9 9 2 7 15 13 10 9 1 10 9 10 3 13 10 9 10 9 1 10 9 13 2
37 15 13 9 14 2 9 2 1 10 9 2 7 15 4 3 13 15 1 10 9 2 13 7 13 10 0 9 7 9 10 10 9 4 16 15 13 2
36 3 3 2 16 15 4 13 1 15 9 13 10 9 2 10 0 2 0 2 0 9 2 4 13 2 3 1 10 0 9 10 0 2 0 9 2
30 10 0 9 15 13 10 9 13 14 13 9 13 15 16 15 13 1 10 9 15 4 13 13 10 9 1 10 9 9 2
7 15 13 0 16 13 9 2
14 16 15 13 9 3 3 2 3 4 14 15 13 9 2
27 15 4 14 13 14 13 1 11 1 9 9 7 13 14 13 3 15 4 14 13 9 1 15 1 15 9 2
6 10 9 4 4 13 2
8 3 13 10 9 1 10 9 2
3 6 3 2
42 15 13 10 9 9 9 1 10 0 9 3 2 7 9 2 3 15 9 13 15 1 15 2 15 13 15 2 7 13 1 10 9 1 10 9 10 9 1 10 9 13 2
51 6 2 3 3 2 3 15 13 10 9 2 13 2 2 15 13 10 0 9 10 0 0 9 1 11 4 13 2 15 13 1 1 15 0 2 0 0 9 2 7 13 16 15 13 14 13 9 1 10 9 2
16 3 2 16 9 4 13 15 10 9 2 15 4 3 13 15 2
22 15 13 1 9 2 15 7 15 1 15 15 13 1 11 4 13 10 0 9 1 15 2
3 15 4 2
18 15 4 13 10 9 1 15 15 4 14 13 7 4 13 14 13 15 2
13 15 4 3 13 10 9 3 10 9 4 4 13 2
33 15 4 13 2 16 16 15 4 13 3 2 13 7 13 15 2 10 0 0 9 4 4 13 1 9 1 9 1 10 0 9 9 2
8 7 15 4 15 13 1 15 2
7 1 2 11 11 2 8 2
10 9 2 11 2 12 11 12 12 2 12
6 1 2 11 2 8 2
10 9 2 9 9 2 11 11 5 10 9
55 15 13 15 0 9 13 1 10 9 2 3 15 13 3 0 16 2 13 2 10 9 15 13 2 7 15 13 15 13 0 16 15 4 3 13 1 0 9 9 1 10 9 1 0 9 1 9 2 7 10 9 1 0 9 2
47 15 13 14 0 16 10 1 15 13 0 1 9 9 2 7 14 13 15 15 4 14 13 2 15 4 13 11 11 2 9 1 11 11 7 11 11 1 0 0 9 9 2 13 9 7 9 2
27 2 15 3 3 13 15 14 13 1 9 9 9 16 11 11 13 1 10 9 1 9 13 1 0 9 2 2
17 10 9 13 1 10 9 13 2 11 7 2 10 11 11 11 2 2
31 16 9 13 10 0 9 2 13 15 2 16 15 13 10 3 0 9 10 10 9 2 9 4 13 7 14 13 15 0 9 2
10 7 15 13 15 15 13 1 9 9 2
20 2 1 10 9 2 13 10 9 1 10 9 9 2 10 3 0 7 0 9 2
25 9 9 4 13 7 13 1 0 9 1 13 9 2 3 10 9 4 13 1 1 12 11 1 9 2
11 15 4 13 1 10 9 16 15 3 13 2
6 15 13 10 0 9 2
18 10 9 13 10 9 14 13 10 9 10 13 0 1 10 9 1 9 2
33 9 2 10 4 13 1 15 9 3 10 9 1 3 3 16 15 4 8 13 2 13 10 9 1 9 13 10 9 3 1 10 9 2
12 2 10 9 13 15 2 9 2 1 9 2 2
26 3 11 14 9 2 2 9 13 3 9 1 10 9 2 10 9 13 9 2 2 4 13 1 10 9 2
22 14 13 12 1 10 3 0 9 15 13 2 9 1 9 4 13 1 15 0 9 2 2
21 10 9 2 7 3 10 9 2 13 15 3 14 13 14 13 10 9 1 10 9 2
28 16 9 13 0 16 13 1 10 9 2 7 16 13 15 9 2 16 15 13 0 7 0 2 15 4 13 15 2
27 7 15 3 13 10 9 13 10 9 14 13 2 3 16 15 13 10 9 9 3 0 15 2 12 12 2 2
7 10 9 1 10 9 13 8
17 16 15 13 10 0 9 2 9 2 15 13 15 9 9 13 0 2
16 3 2 16 9 13 14 13 11 14 0 9 2 13 15 13 2
7 15 13 3 1 10 9 2
32 15 13 3 10 9 3 15 13 15 10 0 0 1 10 9 3 2 7 15 13 12 1 10 0 9 1 15 16 13 3 0 2
6 15 13 10 13 0 2
4 6 1 3 2
2 11 11
4 9 9 2 12
15 2 9 1 11 2 4 15 13 15 9 4 13 15 9 2
5 11 13 14 0 2
2 9 2
3 2 11 2
1 2
4 5 13 0 5
4 13 9 2 2
6 10 13 14 10 9 2
27 15 13 15 1 10 9 9 7 13 14 13 15 2 15 4 14 13 1 10 0 0 9 10 9 3 13 2
8 10 15 13 13 2 15 13 2
4 13 0 9 2
4 6 13 15 2
12 1 12 9 2 15 13 13 9 1 10 9 2
4 15 13 0 2
15 15 13 15 4 13 3 2 7 10 9 3 13 13 3 2
11 1 15 0 9 2 15 13 3 5 12 2
18 1 10 9 1 10 0 9 15 4 13 10 9 1 0 1 5 12 2
16 1 10 0 9 15 13 0 1 5 12 7 15 4 3 13 2
22 15 13 3 15 0 9 7 15 4 13 10 9 1 5 12 7 15 4 3 13 3 2
24 15 13 3 1 5 12 7 12 9 2 7 15 4 13 0 1 15 1 10 9 16 3 13 2
15 13 15 13 15 3 15 13 7 3 3 2 3 15 13 2
25 3 13 0 15 13 15 3 3 2 16 15 4 13 10 9 1 1 15 2 16 15 4 13 15 2
27 15 13 15 16 16 15 13 10 9 3 1 15 4 13 13 0 9 16 15 13 0 16 13 9 3 0 2
8 9 2 13 10 0 9 3 2
8 2 13 15 1 7 13 15 2
11 13 10 0 9 7 13 10 9 13 3 2
4 15 13 0 2
4 15 13 0 2
13 7 2 15 9 13 3 5 12 2 7 9 2 2
2 0 2
27 15 13 14 10 9 2 9 2 15 13 0 2 15 13 0 2 7 15 13 3 10 9 2 15 3 13 2
15 16 10 10 13 9 4 13 1 2 15 4 13 0 9 2
3 6 13 2
20 6 13 10 9 3 2 7 5 12 7 0 4 13 15 1 12 1 12 9 2
14 10 9 13 0 1 1 10 9 7 9 1 10 9 2
11 6 13 15 9 16 3 13 1 10 9 2
12 15 4 3 13 10 9 1 10 9 9 9 2
10 15 13 1 10 9 16 13 9 9 2
13 0 0 9 13 0 14 13 0 9 1 0 9 2
30 3 2 10 9 13 1 10 9 9 13 0 1 9 10 4 13 16 9 1 15 7 15 13 14 4 13 1 10 9 2
9 3 13 10 12 0 9 1 9 2
3 9 12 2
25 13 12 0 9 1 9 7 13 10 13 1 10 9 1 9 2 6 13 15 1 15 9 9 2 2
35 3 13 12 11 5 12 9 7 13 12 1 1 10 1 10 12 9 1 9 16 10 9 4 14 4 13 1 10 9 2 14 13 9 2 2
15 3 2 13 12 9 1 10 1 10 12 9 7 13 15 2
30 15 3 4 13 12 13 9 2 10 1 10 9 1 9 13 10 3 9 2 15 9 7 9 2 7 10 5 12 9 2
9 15 15 4 13 13 13 10 9 2
6 10 13 3 0 2 2
13 15 4 13 10 0 9 7 15 4 13 1 15 2
20 1 0 1 15 15 13 10 0 0 7 0 0 1 10 0 9 1 15 10 2
22 3 15 13 15 1 1 10 11 11 11 2 12 2 7 15 13 16 15 13 3 0 2
9 13 10 12 9 1 10 13 9 2
13 8 2 11 11 12 2 12 11 11 11 11 12 11
13 8 2 11 11 9 9 12 11 11 2 11 12 11
18 8 2 11 11 7 11 11 12 11 11 2 9 12 11 2 11 12 11
11 8 2 11 11 11 11 12 12 11 11 11
14 8 2 11 11 12 11 11 11 9 12 11 2 11 12
45 9 12 2 3 13 10 9 12 9 1 10 9 10 15 13 3 2 13 10 0 9 3 2 12 13 12 2 12 13 12 2 7 8 2 7 13 15 9 1 9 12 1 10 9 2
3 9 12 2
18 13 9 15 13 14 7 13 14 13 10 9 3 0 1 0 16 0 2
13 3 13 15 13 9 1 3 3 12 9 9 2 5
10 2 15 13 15 13 0 1 12 9 2
20 10 15 13 13 12 2 7 13 2 10 0 15 13 2 10 0 9 15 13 2
5 15 13 3 0 2
20 16 15 13 10 9 2 13 1 9 12 9 12 7 12 1 10 0 9 9 2
23 13 10 9 1 10 9 1 15 7 3 15 13 9 2 15 4 13 15 3 2 7 3 2
24 6 13 16 10 9 13 0 1 1 10 9 7 9 1 10 9 7 16 15 3 13 1 9 2
6 13 1 15 10 9 2
24 16 15 13 1 9 2 10 9 4 13 7 10 9 10 3 0 9 4 13 4 13 15 9 2
30 9 2 15 4 13 14 13 10 9 7 9 13 1 15 2 7 1 10 9 7 0 9 7 13 10 9 9 13 15 2
10 15 13 16 15 4 3 13 10 9 2
27 2 3 2 15 4 13 10 0 9 14 13 10 5 12 9 1 0 9 14 13 10 9 1 9 9 2 2
30 3 2 16 10 9 4 13 7 10 9 3 13 2 10 9 4 4 13 1 15 9 1 10 9 9 1 12 9 10 2
28 15 9 4 13 1 10 9 3 16 16 3 15 9 13 10 9 12 9 15 4 4 13 9 1 9 1 9 2
20 10 10 9 1 3 5 12 2 5 12 1 10 1 10 0 12 9 13 3 2
17 13 15 3 2 13 15 0 9 1 10 9 7 15 13 1 9 2
11 2 9 16 3 14 13 1 9 9 2 2
18 9 12 2 15 4 14 13 14 13 10 0 9 14 13 15 0 9 2
31 3 13 15 9 1 10 9 1 10 9 7 13 15 9 1 10 9 1 10 9 2 7 13 2 9 2 1 10 9 9 2
12 15 4 13 10 0 9 1 10 9 14 9 2
3 9 12 2
19 13 10 0 2 9 2 9 7 13 15 9 1 10 9 1 10 0 9 2
11 1 10 2 9 2 9 13 2 9 2 2
22 15 4 13 10 9 1 10 9 1 10 9 16 16 15 4 13 15 9 1 10 9 2
3 9 12 2
10 13 15 0 9 9 1 10 9 9 2
22 16 15 13 14 13 15 9 1 0 9 2 15 4 3 13 10 9 14 13 3 1 2
3 9 12 2
26 13 9 9 7 13 10 9 1 10 0 9 16 13 10 9 1 10 9 7 13 9 1 10 9 9 2
32 13 1 10 9 2 15 4 13 10 9 10 9 13 16 15 13 1 10 9 1 9 1 10 0 9 2 13 10 13 9 9 2
4 15 13 0 2
2 9 2
4 10 13 15 2
11 10 15 13 14 13 2 7 15 3 13 2
2 0 9
11 11 11 2 15 13 11 1 11 11 11 2
3 1 11 11
3 11 11 11
10 11 2 11 2 11 12 2 11 2 2
36 3 16 15 13 1 11 11 11 14 9 7 13 1 10 9 1 12 2 9 1 10 11 11 11 2 10 11 11 11 4 13 10 3 0 9 2
39 1 0 1 1 10 9 2 10 0 9 4 3 13 1 10 0 12 9 1 10 9 2 1 1 10 0 9 9 1 11 11 11 11 1 11 14 11 11 2
12 10 0 9 4 13 1 11 11 11 1 12 2
32 0 9 7 9 9 2 1 15 9 10 9 9 4 13 2 3 13 15 9 1 10 9 7 13 15 1 1 10 9 3 13 2
18 15 9 4 13 2 15 9 4 13 7 3 10 0 9 4 4 13 2
18 1 10 0 9 2 9 2 9 1 1 11 7 11 13 3 1 9 2
18 1 9 7 11 2 0 9 13 14 13 0 0 9 2 3 1 11 2
28 1 10 9 2 10 9 13 10 9 1 10 11 9 3 13 10 0 9 2 3 13 15 3 15 9 13 0 2
13 16 3 2 10 0 9 4 14 4 13 1 3 2
31 9 3 13 15 10 0 9 13 10 13 9 1 11 7 13 15 1 10 9 3 1 10 9 2 13 14 13 10 13 9 2
7 16 0 2 10 9 13 2
13 1 9 2 10 9 14 9 13 14 13 15 9 2
23 3 2 10 9 1 9 13 16 13 10 9 3 1 15 0 9 9 1 10 0 11 11 2
37 10 9 13 1 10 9 2 13 16 12 9 4 13 1 11 1 12 1 10 11 11 7 11 11 2 16 1 10 0 7 3 2 13 9 1 9 2
28 10 9 9 4 13 2 7 3 15 13 10 13 12 9 13 10 0 11 2 3 3 12 9 3 15 13 9 2
34 12 0 9 1 9 13 10 9 13 1 10 9 9 2 10 9 10 13 10 9 2 9 7 9 1 10 0 9 1 9 1 15 9 2
16 10 0 9 13 1 11 11 11 4 13 0 9 1 10 9 2
57 11 9 9 11 11 7 11 11 4 13 16 9 3 13 9 2 9 9 2 16 15 4 13 10 9 10 0 9 1 2 10 9 1 9 2 2 9 10 13 1 10 0 9 13 1 10 9 14 9 1 11 11 7 10 11 11 2
40 15 13 16 9 1 11 13 14 13 0 1 0 9 7 9 13 1 10 9 1 9 2 10 9 10 13 10 9 16 13 0 9 7 13 10 9 1 9 9 2
43 1 9 2 3 2 11 7 11 4 13 2 9 1 10 9 3 4 13 10 9 16 13 3 0 9 1 9 9 2 3 15 13 3 1 10 0 2 7 13 1 10 9 2
33 2 10 15 13 14 13 13 13 1 10 9 2 2 11 11 2 9 9 9 1 10 11 11 7 11 11 2 13 11 14 11 11 2
8 2 15 13 2 2 6 2 2
19 10 9 10 13 14 13 0 1 10 9 9 13 3 10 9 1 9 2 2
12 10 0 9 4 13 10 0 0 9 1 11 2
15 0 0 9 7 9 4 13 0 9 1 9 2 1 9 2
24 3 15 4 13 3 12 9 9 1 10 9 14 0 9 16 10 9 13 2 3 15 13 12 2
17 2 15 4 13 0 1 10 9 1 9 2 2 11 13 11 11 2
18 2 15 13 10 9 1 9 1 9 7 15 13 2 2 15 13 2 2
9 7 15 4 4 13 1 0 9 2
34 1 9 9 2 9 9 2 9 7 9 13 9 1 0 9 2 9 2 10 0 9 1 0 9 2 9 2 13 9 10 13 4 13 2
11 15 13 0 1 9 1 10 9 1 9 2
11 10 9 13 9 7 9 9 1 9 9 2
8 9 13 0 1 9 9 2 2
15 11 13 10 0 9 9 2 12 1 10 0 1 10 9 2
24 11 13 16 10 9 1 9 4 14 13 3 3 16 10 9 13 3 2 15 9 13 3 0 2
16 2 15 13 3 0 16 13 0 9 2 2 3 2 15 13 2
7 2 9 13 3 3 0 2
9 15 4 3 13 3 1 12 9 2
12 1 12 0 9 15 4 13 10 0 9 2 2
41 9 9 1 10 0 11 4 13 3 0 10 11 7 11 11 4 13 14 13 10 9 14 9 1 9 1 9 7 2 3 2 14 13 15 1 10 0 9 9 3 2
20 11 13 10 9 4 13 0 9 9 1 10 0 11 2 16 13 1 0 9 2
24 10 9 13 10 9 13 16 9 4 13 1 0 9 2 13 11 2 11 7 11 2 1 9 2
18 1 11 12 2 11 11 11 11 11 11 11 11 13 14 13 1 15 2
12 15 13 10 11 9 14 13 10 9 14 9 2
10 11 13 15 9 4 3 13 10 9 2
18 3 1 10 9 14 0 9 2 15 0 9 1 0 9 3 13 0 2
6 9 4 13 0 9 2
25 10 11 9 4 13 0 2 13 1 10 9 2 1 10 11 9 0 9 2 0 12 9 1 9 2
20 3 2 15 9 13 14 4 13 2 16 11 13 10 2 3 0 0 9 2 2
19 15 13 3 3 12 9 1 10 0 2 7 15 13 10 13 12 9 9 2
15 9 1 9 2 9 9 13 0 9 7 0 9 1 9 2
19 15 3 3 13 9 2 10 9 4 14 2 1 10 9 1 10 11 11 2
17 7 9 13 0 2 3 0 2 14 13 9 9 2 1 10 9 2
18 15 13 14 4 13 16 15 4 13 10 0 9 1 10 13 0 9 2
14 13 10 9 1 9 13 1 11 0 1 10 0 9 2
9 15 13 14 13 3 10 2 9 2
18 0 2 15 13 3 12 9 7 9 9 13 1 9 1 10 11 11 2
37 15 3 13 0 9 4 13 10 1 10 9 1 10 9 13 15 4 13 2 1 9 2 10 9 1 11 11 13 9 1 10 0 9 14 3 3 2
23 11 13 10 9 4 14 13 14 13 1 10 9 2 3 2 7 15 10 3 3 4 13 2
37 15 13 1 12 9 1 9 9 1 0 11 9 2 9 4 14 13 10 0 9 10 4 14 13 1 12 1 10 9 10 9 13 2 7 15 9 2
1 2
22 11 11 13 10 0 9 13 10 9 1 9 1 10 9 2 1 9 0 9 11 11 2
3 9 2 8
7 9 2 9 13 2 9 13
3 1 11 11
3 11 11 11
10 11 2 11 2 11 12 2 11 2 2
41 9 4 13 3 15 13 1 3 0 9 11 2 7 11 2 10 9 4 13 7 15 10 9 13 2 7 3 11 14 9 2 9 7 9 4 14 13 1 10 9 2
15 15 3 4 13 15 9 1 9 1 9 16 15 4 13 2
43 15 13 1 12 1 10 0 9 1 10 13 9 13 10 9 1 10 0 0 9 1 13 9 2 7 9 15 13 10 9 4 13 0 1 10 9 10 9 4 13 0 9 2
38 11 11 11 2 10 9 9 7 9 1 10 9 9 11 11 2 13 10 12 9 1 10 11 1 10 11 11 1 11 1 15 12 2 9 0 0 9 2
15 9 13 10 9 14 9 7 9 9 2 10 9 1 9 2
31 11 14 9 1 12 9 13 16 3 0 1 12 2 9 4 13 1 0 9 0 9 3 1 1 10 0 9 1 15 9 2
14 9 13 3 1 15 9 1 10 9 7 9 13 3 2
14 10 0 9 4 13 1 3 12 9 16 15 13 14 2
12 10 9 9 4 13 1 0 11 3 1 11 2
14 9 1 10 12 9 11 13 13 10 9 0 1 9 2
8 1 11 2 10 9 13 3 2
31 10 9 1 12 9 9 1 10 11 11 13 3 12 2 9 4 13 15 9 12 1 12 9 3 16 15 4 12 9 3 2
66 2 12 1 10 0 2 3 3 2 13 7 0 9 1 9 1 10 0 9 4 13 10 0 9 1 9 16 13 10 0 9 1 9 7 0 9 2 2 13 10 9 13 2 13 11 1 11 11 11 1 10 11 11 2 2 13 1 10 11 11 1 11 11 0 9 2
19 11 9 13 1 3 12 9 10 4 13 10 9 16 16 9 4 13 9 2
44 2 9 1 10 9 13 0 9 1 10 0 9 1 10 0 9 7 9 9 2 2 13 11 11 2 10 11 1 11 2 11 9 7 12 1 10 9 14 13 9 1 10 9 2
14 10 9 4 13 1 10 9 2 11 13 11 14 11 2
20 2 1 10 11 11 2 10 0 9 1 9 14 9 4 13 2 2 15 13 2
20 11 4 13 0 1 15 9 13 10 9 9 2 10 13 1 11 7 0 11 2
12 10 13 9 3 4 13 1 10 1 15 9 2
16 2 0 9 13 1 9 16 13 10 0 9 2 2 15 13 2
24 2 15 4 13 0 9 1 9 9 1 11 7 0 11 1 9 3 10 9 13 3 0 2 2
43 13 1 11 14 0 9 2 12 9 9 2 1 9 2 4 13 3 10 9 9 13 3 3 2 13 1 10 13 9 9 2 3 4 13 1 10 0 9 1 15 0 9 2
16 1 10 11 11 2 15 13 2 2 9 13 3 12 9 0 2
8 9 9 4 13 12 9 3 2
12 0 9 4 13 1 1 11 7 10 11 11 2
20 9 7 9 9 4 13 0 2 0 0 9 13 3 1 11 7 10 11 2 2
27 16 10 11 9 13 2 2 0 9 3 13 14 13 16 10 9 1 9 9 13 3 0 1 11 9 2 2
21 0 9 13 9 7 2 1 10 9 2 9 1 9 7 9 1 9 9 1 9 2
15 10 9 3 13 9 1 9 9 0 1 9 9 7 9 2
66 10 0 9 2 1 9 2 4 13 16 13 10 9 9 1 9 9 2 13 7 13 0 9 1 10 9 16 15 13 2 1 2 13 10 9 9 1 9 2 13 0 9 16 4 13 2 16 0 9 4 13 0 9 9 3 13 1 10 9 14 13 7 13 9 2 2
18 10 11 9 13 1 10 9 1 11 1 10 2 11 11 11 11 2 2
31 10 11 2 1 9 1 10 11 11 2 11 2 11 2 11 2 11 2 11 2 10 11 11 7 11 2 4 13 1 12 2
21 2 10 9 1 0 9 4 13 9 3 1 10 11 2 2 13 11 9 11 11 2
17 2 10 11 4 13 10 1 10 3 0 7 0 9 9 1 11 2
23 10 9 1 9 9 1 10 9 7 10 9 4 13 14 13 3 1 10 9 14 13 2 2
33 10 11 13 0 9 9 4 13 12 9 1 12 9 11 1 10 0 12 9 7 4 13 3 3 3 3 3 1 10 0 12 9 2
32 0 9 9 9 4 13 1 12 9 1 10 9 1 10 0 9 2 10 9 13 2 16 10 9 13 0 9 1 9 9 9 2
33 2 4 10 11 11 13 9 2 0 1 9 2 15 13 0 16 0 9 7 10 9 9 4 4 13 1 9 2 2 10 9 13 2
15 1 1 3 0 9 9 2 3 9 13 1 10 0 9 2
42 10 0 9 2 2 10 11 1 11 11 2 10 11 1 10 11 2 2 13 1 10 11 2 13 11 11 11 7 13 3 3 1 10 0 12 2 13 3 1 10 9 2
28 1 10 12 9 2 10 11 9 13 2 9 9 3 13 16 10 9 9 1 10 11 4 3 13 10 0 9 2
31 15 13 3 1 10 0 11 3 10 9 9 4 13 14 13 3 1 10 9 16 10 9 9 1 0 9 4 3 13 2 2
21 1 10 0 9 2 10 9 13 10 9 4 14 13 3 0 1 10 11 11 9 2
22 2 10 9 1 0 9 1 9 9 7 9 13 0 14 13 2 2 10 11 9 13 2
24 2 10 9 1 10 9 13 13 3 0 16 14 14 13 0 1 10 9 1 10 11 11 2 2
35 10 0 0 9 10 3 4 13 1 9 13 9 2 9 2 9 2 9 2 0 9 7 0 9 1 9 7 9 2 0 1 10 11 9 2
19 0 9 10 3 4 13 13 9 2 9 2 11 9 7 10 9 1 9 2
32 13 1 10 9 9 2 7 1 10 9 1 9 13 1 10 11 9 2 4 12 1 10 0 9 13 9 1 10 0 9 9 2
22 10 11 9 13 0 9 9 2 7 15 13 0 0 9 2 0 1 9 7 0 9 2
19 1 10 0 0 9 2 3 2 10 9 4 13 9 4 13 10 0 9 2
19 10 9 13 16 15 13 15 13 1 10 0 9 2 9 9 7 0 9 2
10 10 11 9 13 14 13 10 0 9 2
24 15 13 10 9 2 0 2 1 0 9 2 7 16 13 3 13 10 9 9 10 9 3 0 2
33 10 9 2 1 2 9 16 13 0 9 13 10 9 10 3 4 13 14 4 13 1 9 2 16 9 7 9 4 13 3 3 3 2
37 2 3 9 4 13 10 9 1 11 1 11 9 2 15 13 9 14 13 1 10 0 9 1 9 2 2 13 11 11 1 2 10 11 11 11 2 2
45 2 13 3 1 10 9 2 13 15 9 1 10 9 2 13 1 10 9 1 9 7 9 2 7 3 15 4 13 15 2 10 9 1 10 9 9 2 3 3 3 1 10 11 2 2
4 7 3 14 2
1 2
15 11 13 10 0 9 1 11 13 10 9 1 0 9 9 2
2 9 8
10 9 1 11 13 1 10 9 3 3 2
22 13 0 14 13 7 13 7 13 15 9 2 16 10 9 13 10 0 9 13 10 9 2
1 5
7 3 4 11 13 10 11 2
18 15 4 13 10 13 9 1 11 11 7 15 4 4 13 1 10 9 2
30 9 9 4 13 14 13 9 1 9 1 13 9 16 9 4 13 14 13 9 1 11 11 13 10 9 1 9 7 9 2
42 1 10 9 9 2 9 13 16 11 4 13 10 0 9 1 10 9 10 11 4 13 1 9 7 3 2 3 13 10 9 1 9 7 0 9 15 13 10 9 4 13 2
20 3 2 11 11 11 11 4 13 15 4 13 10 9 16 3 10 9 4 13 2
7 3 4 11 13 10 11 2
6 4 15 13 15 9 2
12 4 10 9 13 10 9 0 9 13 10 11 2
8 13 15 15 9 13 10 9 2
1 5
6 10 1 10 0 9 2
47 2 1 10 11 2 15 4 13 14 13 10 9 14 13 10 10 2 11 7 11 9 2 16 15 4 13 1 10 9 1 2 9 2 10 4 13 10 9 1 15 9 14 13 15 0 9 2
33 15 15 13 1 11 11 13 10 0 9 1 10 9 1 10 9 9 2 10 9 1 9 10 0 1 10 9 13 13 10 0 9 2
6 15 4 13 10 9 2
12 15 9 13 15 13 9 2 7 15 13 14 2
11 15 13 10 9 9 10 13 11 11 2 2
6 2 11 2 11 2 11
26 2 15 4 3 13 1 10 9 1 10 11 2 9 2 2 6 9 2 7 15 4 13 15 13 2 2
24 10 0 9 13 16 11 13 10 9 0 1 10 9 1 0 9 1 10 0 9 1 15 9 2
16 3 3 15 4 14 13 10 9 1 0 0 9 2 9 2 2
4 2 11 2 11
104 2 15 4 14 13 15 4 13 10 11 9 10 13 15 4 13 2 3 3 10 9 13 2 9 2 1 10 9 15 4 13 10 9 3 1 10 0 9 1 10 9 7 13 14 13 2 3 10 0 9 2 10 13 15 13 15 13 1 10 9 1 0 9 2 4 13 15 9 2 3 14 13 9 1 1 15 9 7 13 1 15 9 2 0 9 1 10 9 13 15 2 2 9 2 13 14 10 9 9 7 9 9 2 2
4 2 11 2 11
10 2 10 9 4 3 3 13 10 11 2
11 9 13 14 15 15 13 1 10 0 9 2
17 3 2 9 13 3 0 2 7 15 4 13 14 13 12 2 3 2
3 2 11 2
23 2 10 11 4 13 15 9 1 10 9 1 10 9 7 15 4 13 9 1 12 0 9 2
13 13 15 1 15 9 2 7 11 13 3 0 2 2
7 2 11 11 2 11 2 11
12 2 11 4 13 3 14 13 1 15 9 3 2
3 2 11 2
11 15 13 3 0 10 9 10 9 4 13 2
15 3 2 9 1 10 11 1 0 9 4 13 10 0 9 2
24 15 4 14 13 16 9 15 13 16 11 13 10 9 1 9 4 13 15 9 1 10 0 9 2
18 15 13 10 9 15 13 3 1 11 16 13 10 0 9 1 10 9 2
17 6 2 15 7 15 9 13 0 14 13 10 0 9 1 10 9 2
14 15 9 13 10 9 1 10 11 3 10 9 1 0 2
17 2 13 15 7 14 2 15 13 10 9 1 12 9 14 13 2 2
27 10 9 10 4 13 1 11 14 13 13 10 0 9 1 10 9 10 11 4 13 1 10 9 1 0 9 2
10 3 1 10 9 0 7 10 0 9 2
18 15 13 2 15 4 13 1 10 11 2 11 11 9 0 1 15 9 2
13 3 14 1 11 2 15 13 1 11 7 11 11 2
53 15 13 10 9 1 0 9 1 10 1 10 9 2 7 15 4 13 1 10 9 2 13 15 9 3 15 13 1 11 2 7 3 15 13 3 7 13 1 10 0 9 13 0 2 0 1 12 5 2 1 0 11 2
37 10 9 13 2 3 15 13 13 1 9 1 11 11 2 3 15 3 13 15 0 2 9 1 11 7 11 2 15 13 0 1 10 9 1 0 9 2
38 15 4 14 13 14 13 10 9 2 7 3 15 4 13 1 15 9 1 11 2 11 11 2 7 9 0 13 3 3 1 15 2 15 13 3 3 0 2
14 3 2 6 2 11 13 9 10 13 3 0 1 9 2
30 3 2 13 10 9 1 11 7 11 1 10 0 9 2 15 4 13 15 3 13 1 10 9 1 10 9 1 12 9 2
16 3 2 15 13 3 14 4 13 2 13 15 1 9 7 9 2
12 10 13 14 13 2 7 3 0 13 0 14 2
17 6 2 15 13 10 0 9 1 11 2 15 4 13 9 1 15 2
21 3 2 11 11 3 13 0 0 9 2 9 15 13 9 3 16 15 13 10 9 2
15 15 4 14 13 16 15 4 13 0 9 14 9 1 11 2
21 15 13 15 4 14 13 3 2 7 15 3 13 3 0 9 9 13 1 10 9 2
12 15 4 13 16 15 4 13 10 9 1 11 2
25 15 13 16 0 1 10 13 9 2 15 0 7 15 3 2 4 13 1 10 9 15 4 13 1 2
33 10 12 12 9 15 4 4 13 1 9 7 9 9 1 11 4 13 14 13 11 2 11 2 11 11 7 11 2 7 10 13 9 2
29 6 2 10 4 13 2 7 15 13 10 9 16 16 0 13 14 13 9 7 0 9 2 15 4 13 0 16 13 2
13 15 13 0 16 15 11 4 13 1 1 12 9 2
16 4 0 9 13 15 9 1 11 16 10 9 4 13 9 3 2
22 7 4 10 3 9 2 0 9 13 3 0 1 15 15 4 3 13 9 1 15 9 2
22 4 10 9 9 1 11 13 13 16 10 9 1 10 9 13 1 1 10 9 1 9 2
22 4 9 10 13 0 1 12 4 13 10 9 9 1 1 15 9 16 13 10 9 9 2
16 15 4 10 0 9 13 14 13 9 1 10 9 7 9 9 2
11 15 13 10 1 10 9 15 4 4 13 2
1 11
4 9 13 3 2
11 15 9 13 0 7 13 9 0 1 9 2
1 11
26 6 2 15 13 0 1 10 9 7 3 4 14 13 11 2 3 15 9 9 13 0 7 15 13 15 2
28 15 3 13 1 10 9 7 16 15 9 7 9 13 16 3 0 13 9 16 9 13 9 3 15 13 10 9 2
17 15 15 13 13 16 15 13 10 0 9 15 9 13 1 11 11 2
18 15 9 4 14 13 9 9 2 3 15 13 10 9 13 7 13 3 2
30 10 9 3 2 11 2 13 14 13 10 9 9 1 3 1 11 2 16 15 4 13 3 16 9 4 13 1 3 3 2
16 10 9 4 14 4 13 16 10 9 13 0 1 15 0 9 2
21 10 9 13 16 9 13 1 10 9 4 13 10 9 9 7 13 16 9 13 0 2
14 15 13 11 12 2 7 3 12 9 9 4 4 13 2
22 15 15 13 13 9 1 9 9 13 10 4 4 4 13 14 13 9 15 13 10 9 2
38 15 15 13 13 10 11 1 11 11 2 13 16 15 4 14 13 10 9 7 9 0 14 4 13 16 15 4 13 1 9 0 14 13 15 15 14 13 2
18 3 0 9 13 10 9 9 1 9 7 0 9 9 15 4 15 13 2
7 3 2 11 13 10 9 2
18 3 12 9 1 15 9 2 15 13 13 10 9 9 3 12 0 9 2
24 3 15 3 13 1 13 7 15 13 10 15 4 13 14 13 15 9 3 1 10 3 13 9 2
15 3 15 4 14 13 16 15 4 13 1 10 0 9 3 2
30 15 13 16 15 13 10 9 10 13 10 0 9 3 2 15 4 14 13 7 13 15 1 10 9 15 9 4 13 0 2
20 3 2 10 9 10 4 4 13 13 0 7 10 0 4 13 1 9 3 3 2
39 10 9 1 15 10 13 16 11 4 13 1 0 9 14 13 0 9 2 3 15 15 4 13 13 13 9 16 13 10 11 0 1 11 7 0 9 8 3 2
29 15 13 10 9 2 16 15 4 13 14 13 9 1 9 13 2 9 2 3 14 13 10 9 13 10 1 15 0 2
28 0 1 9 2 0 1 9 9 2 7 0 1 0 9 10 4 13 15 0 1 10 0 9 9 2 15 2 2
15 15 13 0 15 13 15 13 14 13 3 15 13 15 1 2
20 1 10 9 15 13 3 13 9 10 4 4 13 0 1 10 9 1 10 0 2
5 1 15 15 13 2
5 11 1 12 2 9
22 16 15 13 10 9 1 12 2 10 0 12 14 13 4 13 2 13 1 10 9 2 2
23 12 4 13 10 9 1 9 7 9 2 7 3 10 0 4 13 0 14 13 16 13 0 2
17 10 11 9 4 13 14 13 15 9 7 13 15 9 1 0 9 2
12 15 4 13 14 13 15 3 7 13 15 9 2
31 15 4 13 1 10 0 14 13 1 0 0 9 14 13 0 9 1 15 2 16 15 9 4 13 1 10 10 2 9 9 2
19 15 4 13 3 0 7 0 1 0 2 7 9 4 13 3 1 15 9 2
20 16 15 13 14 13 10 0 0 9 7 9 9 2 15 9 4 4 13 3 2
15 12 4 13 15 13 3 3 2 7 13 14 13 3 3 2
5 11 1 12 2 9
12 2 9 2 13 10 0 9 1 15 2 11 2
25 1 0 9 7 9 2 15 4 13 3 3 12 0 9 10 4 13 1 15 9 1 10 0 9 2
33 15 13 10 9 15 4 13 14 13 9 1 15 9 7 13 15 16 15 4 13 10 9 15 13 14 13 1 10 9 1 15 9 2
14 16 10 9 13 2 10 3 0 15 9 7 9 13 2
20 1 10 9 2 15 9 13 2 7 15 0 9 4 13 0 9 1 15 9 2
34 1 10 9 1 10 9 2 15 4 13 10 0 0 9 1 9 7 9 9 2 13 0 9 7 13 3 15 0 9 10 9 7 12 2
5 11 1 12 2 9
38 15 9 16 13 1 10 9 1 0 9 4 13 1 10 9 2 11 2 7 3 15 4 13 14 13 13 10 9 10 2 9 2 4 13 1 15 9 2
11 16 12 13 2 10 9 3 4 13 0 2
18 15 3 13 15 1 15 14 13 10 9 1 9 1 15 10 15 13 2
10 10 9 7 9 3 13 9 7 9 2
24 15 9 1 9 1 10 9 13 1 0 9 9 2 13 15 9 1 10 0 0 9 10 9 2
32 1 10 9 1 12 15 4 13 10 0 0 9 1 9 1 15 9 7 15 9 9 2 7 10 0 0 9 14 13 15 1 2
5 11 1 12 2 9
19 13 10 9 1 15 0 7 0 9 4 13 12 1 10 9 14 0 9 2
28 1 10 0 9 2 15 0 9 10 9 4 13 1 9 7 9 2 13 9 1 0 9 1 9 1 0 9 2
8 13 10 0 9 3 15 4 2
7 10 0 9 4 13 0 2
33 15 4 4 13 0 9 1 15 9 9 2 7 15 4 13 10 9 0 1 15 2 7 1 10 9 15 4 13 15 13 0 15 2
19 15 9 9 13 0 2 7 10 9 1 9 7 9 9 13 1 10 9 2
27 1 10 9 1 12 2 15 4 13 3 0 2 3 0 2 7 3 3 0 16 13 10 9 13 1 15 2
5 11 1 12 2 9
31 13 10 0 9 2 1 1 10 0 0 7 0 9 2 4 13 0 10 9 16 15 4 1 10 0 9 1 15 2 11 2
22 10 3 0 9 4 13 13 10 9 13 10 0 1 15 2 7 3 14 13 15 9 2
15 15 4 13 0 14 13 9 1 9 3 1 1 0 9 2
22 9 1 12 4 13 15 10 9 14 13 2 7 15 4 13 10 9 1 10 15 9 2
6 9 13 3 7 3 2
11 9 4 3 13 0 1 10 3 0 9 2
31 7 2 15 13 10 9 1 10 9 15 4 13 3 2 7 1 10 9 1 12 2 15 4 13 3 1 0 9 7 9 2
5 11 1 12 2 9
13 15 9 9 4 14 13 3 3 10 9 2 11 2
15 1 9 1 12 2 15 4 4 13 15 9 1 10 9 2
12 1 10 0 9 2 15 9 4 13 3 0 2
17 3 4 14 13 15 1 13 2 15 3 13 14 13 0 10 9 2
28 15 9 9 4 13 1 0 1 10 9 2 7 10 9 13 7 13 1 12 13 3 0 14 13 10 0 9 2
12 7 2 15 4 13 14 13 10 0 0 9 2
31 1 9 1 10 9 1 9 1 15 9 2 1 10 9 14 9 2 15 4 13 16 12 4 13 15 9 1 9 7 9 2
5 11 1 12 2 9
15 13 15 9 2 9 11 2 7 13 1 10 3 0 9 2
21 1 0 11 1 15 9 2 15 13 3 15 9 2 3 3 15 0 9 13 0 2
6 9 7 9 13 3 2
23 16 15 13 14 3 0 2 7 13 14 13 2 15 3 4 13 1 10 9 1 10 9 2
26 15 13 10 9 15 4 13 14 4 13 10 9 1 9 7 13 1 15 9 2 16 9 13 10 9 2
30 10 12 9 1 9 10 4 14 3 13 3 0 16 15 4 13 4 13 15 9 2 3 9 4 13 0 7 9 0 2
20 1 9 14 9 2 15 4 13 15 3 13 10 0 9 2 10 1 10 0 2
5 11 1 12 2 9
26 11 2 15 4 3 13 9 2 3 0 9 2 1 15 9 10 9 2 3 1 10 9 1 0 9 2
26 16 15 13 3 0 1 10 9 1 15 9 2 15 4 13 15 13 1 1 0 0 9 1 15 9 2
15 15 9 4 13 1 10 3 0 9 15 4 3 13 1 2
10 15 4 3 13 15 9 1 10 9 2
30 16 15 13 10 9 1 10 0 9 13 1 10 9 2 7 15 4 13 0 1 0 9 2 9 1 9 4 13 3 2
6 13 0 1 0 9 2
12 15 4 14 13 0 2 7 15 4 13 0 2
16 4 14 13 1 10 9 2 3 2 13 1 10 9 1 12 2
5 11 1 12 2 9
8 13 15 0 14 13 0 9 2
8 16 14 2 15 4 13 3 2
24 15 13 9 2 11 2 4 13 1 10 0 9 1 11 2 13 2 0 9 2 2 1 12 2
15 15 13 3 0 9 13 1 10 9 16 15 13 3 0 2
15 15 4 13 10 0 9 13 10 9 14 13 15 0 9 2
24 15 4 13 0 9 16 13 15 9 1 10 9 16 13 0 9 10 13 15 14 13 3 3 2
29 1 10 0 9 1 10 9 2 15 4 3 13 0 9 1 10 0 0 9 10 4 13 15 1 10 0 12 9 2
23 7 2 10 9 15 13 3 4 13 10 3 0 9 2 6 2 1 10 9 1 15 9 2
14 3 2 12 13 0 14 13 10 9 15 4 14 13 2
5 11 1 12 2 9
16 15 4 13 9 1 0 9 13 15 9 1 12 2 9 11 2
34 10 3 13 9 15 4 13 1 15 9 9 13 1 10 9 2 7 1 10 9 1 10 9 15 4 13 3 0 1 15 9 1 0 2
20 3 2 15 4 13 10 0 9 2 16 10 0 9 4 13 15 13 10 9 2
19 15 9 9 4 13 3 2 7 15 13 0 14 13 9 7 9 10 9 2
40 1 9 2 10 9 1 15 9 7 9 9 4 13 0 2 7 13 13 15 4 13 1 15 0 2 7 0 2 1 3 2 16 0 4 13 7 13 1 12 2
5 11 1 12 2 9
14 12 13 15 13 15 0 7 0 9 3 3 2 11 2
34 10 9 1 10 9 13 14 13 7 13 15 2 16 15 13 15 0 9 1 10 0 9 0 1 15 9 2 3 13 9 1 10 9 2
27 12 13 0 14 13 3 3 12 0 9 1 10 9 9 2 7 15 9 4 4 13 1 0 9 7 9 2
22 14 3 10 2 7 9 2 9 2 7 0 9 13 0 9 1 10 9 1 15 9 2
27 1 9 14 9 2 15 0 9 2 9 4 4 13 15 1 0 0 9 2 7 10 0 0 9 1 3 2
7 11 1 12 2 9 2 9
11 15 13 10 0 9 1 15 2 9 11 2
18 3 3 2 1 12 15 4 13 15 13 3 7 3 3 1 10 9 2
15 15 4 13 10 0 9 1 9 7 13 9 1 0 9 2
29 13 9 1 9 7 0 9 10 9 2 16 11 13 10 0 1 15 9 2 15 9 9 2 7 10 9 1 0 2
31 1 10 9 1 10 9 2 15 4 13 1 10 0 9 2 13 1 10 0 9 9 2 7 3 13 10 9 1 15 9 2
33 15 13 0 16 15 13 9 7 9 1 9 1 15 14 13 2 16 10 9 1 9 1 15 0 7 0 9 4 13 0 7 0 2
15 13 0 7 0 2 7 9 13 3 0 14 13 1 12 2
11 2 13 10 0 2 2 7 13 10 9 2
10 2 9 13 1 9 2 3 1 10 9
4 11 2 2 2
5 13 9 9 2 2
7 13 15 9 2 8 2 8
4 13 15 2 12
6 13 1 15 2 8 2
6 2 13 3 3 3 2
1 8
3 12 12 9
1 2
28 10 0 11 11 4 13 1 10 0 0 0 9 11 11 15 13 5 11 11 13 10 11 5 2 12 5 12 2
2 2 2
1 2
19 1 11 11 11 2 10 9 2 13 1 15 11 9 11 7 11 14 9 2
1 2
10 11 0 9 2 11 12 2 12 9 11
11 11 13 1 11 2 11 12 2 12 9 11
11 11 14 11 11 13 2 11 12 2 12 11
9 11 13 11 2 11 12 2 12 11
8 11 13 2 11 12 2 12 11
10 11 11 14 9 2 11 12 2 12 11
10 11 11 11 13 2 11 12 2 12 11
14 2 9 1 11 2 11 11 13 2 11 12 2 12 11
12 2 11 2 4 11 13 3 2 11 2 6 2
9 2 11 9 12 2 9 12 2 2
10 11 13 1 9 2 11 12 2 12 11
8 11 13 2 11 12 2 12 11
9 11 13 2 11 12 2 12 11 11
11 11 11 14 9 2 11 12 2 12 11 11
16 9 1 5 10 11 7 10 11 5 2 11 12 2 12 11 11
8 11 11 2 11 12 2 12 11
13 0 11 11 13 2 11 12 2 12 11 5 11 2
1 2
13 2 1 10 9 1 11 2 11 10 11 4 13 2
21 1 10 0 9 15 13 11 2 13 10 0 9 1 9 2 7 13 10 0 9 2
26 7 13 10 9 3 0 1 15 9 11 2 7 1 10 0 9 15 13 11 2 2 2 11 11 2 11
1 2
14 11 11 12 5 12 2 11 11 14 0 11 1 11 2
24 2 16 2 11 14 11 4 13 2 15 13 10 9 11 11 11 11 2 0 1 9 7 9 2
59 10 0 9 2 11 11 2 13 11 1 12 7 13 0 1 11 7 11 11 2 1 15 1 10 9 15 13 14 4 13 1 9 1 9 2 10 4 14 13 3 3 2 7 10 11 13 3 0 9 7 9 16 15 13 0 1 9 9 2
18 1 12 11 13 7 13 10 9 1 10 13 9 1 2 11 11 2 2
48 1 10 9 11 4 13 11 11 2 10 9 1 11 2 7 13 1 15 2 2 15 13 3 0 2 3 0 2 3 0 2 3 0 2 16 15 13 2 3 0 2 16 15 4 13 15 2 2
7 2 9 12 2 9 12 2
31 14 13 10 9 3 0 7 0 2 11 11 13 2 10 3 0 7 0 9 2 2 7 3 3 13 15 1 15 9 9 2
13 10 9 1 11 14 9 3 13 11 1 11 2 2
1 2
16 11 11 11 2 9 12 2 9 12 2 11 2 12 11 12 2
7 1 2 11 11 2 8 2
10 9 2 11 2 12 11 12 12 5 12
13 9 2 1 2 9 2 9 1 9 2 11 2 11
14 2 15 13 10 11 1 11 14 13 1 1 10 9 2
65 0 2 7 12 1 11 10 15 13 1 13 10 9 1 10 11 9 2 11 11 2 15 4 13 9 1 11 14 9 2 9 2 10 11 1 11 2 4 3 13 10 0 11 1 10 3 0 9 2 7 11 11 2 15 13 10 9 1 11 11 1 10 0 9 2
33 14 13 0 2 7 11 7 11 13 9 2 7 15 4 13 1 1 11 16 13 2 16 15 3 13 2 3 3 3 2 11 2 2
1 2
24 2 11 11 11 2 12 5 12 2 13 10 0 0 9 13 1 11 16 13 14 13 11 11 2
23 10 12 9 0 11 11 4 13 0 7 4 3 13 7 13 1 11 12 2 12 1 11 2
45 3 3 2 11 12 2 11 11 4 13 10 0 9 9 1 11 11 7 10 0 9 4 13 14 13 10 9 9 1 11 11 2 13 16 15 4 2 3 2 13 1 10 9 2 2
23 10 0 9 2 12 2 10 0 9 13 11 11 3 13 10 9 1 10 9 9 1 11 2
32 11 14 12 9 2 8 8 8 8 8 8 8 8 8 8 8 2 13 10 9 1 9 9 2 13 10 9 10 13 15 9 2
1 2
5 9 9 12 5 12
2 2 2
10 12 11 2 11 13 1 11 2 11 2
6 0 9 7 13 9 2
13 12 11 2 11 9 1 11 2 13 7 13 9 2
16 12 11 2 11 2 3 11 11 2 10 11 2 13 1 11 2
21 12 11 2 11 11 11 2 11 1 11 2 13 16 13 9 1 15 9 1 11 2
8 12 11 11 1 11 13 9 2
5 12 9 4 13 2
11 12 11 11 13 11 7 13 10 10 9 2
9 12 0 9 9 13 12 0 9 2
14 12 11 11 13 10 12 2 9 9 14 13 10 9 2
9 12 11 11 13 15 9 1 9 2
5 13 10 9 9 2
5 2 11 2 12 2
14 12 11 11 2 10 0 9 2 13 9 1 15 9 2
10 12 11 9 11 2 11 13 1 11 2
6 9 1 0 9 9 2
10 12 11 11 13 0 0 9 1 11 2
14 12 11 7 11 13 11 7 11 1 9 1 11 11 2
8 12 11 13 11 11 1 11 2
14 12 1 10 11 1 11 2 10 9 1 9 4 13 2
12 12 11 13 9 2 7 13 15 9 13 9 2
12 12 11 11 11 1 11 13 10 0 9 9 2
5 12 11 9 13 2
12 12 11 10 11 13 16 13 10 9 1 9 2
14 12 11 14 9 13 1 11 1 11 7 13 1 11 2
1 2
102 2 2 15 4 13 15 2 9 2 2 13 10 9 2 2 16 15 4 13 14 13 15 0 9 2 7 16 1 3 2 13 9 9 1 9 2 9 2 7 9 4 13 1 10 9 1 15 15 4 14 13 2 7 4 14 13 2 7 13 0 1 13 2 3 9 1 10 9 4 13 14 4 13 2 1 10 9 16 2 15 3 13 10 9 2 15 4 13 9 3 0 16 14 13 10 1 15 1 0 9 2 2
85 2 2 6 3 2 2 13 11 11 2 2 10 0 9 13 1 10 9 7 9 1 10 9 2 3 10 13 9 2 9 9 2 7 2 1 0 2 10 10 9 10 4 4 13 1 10 9 2 7 3 15 13 3 2 15 13 14 13 3 9 13 2 9 13 15 10 1 10 9 10 13 12 1 10 0 2 7 10 13 0 1 10 9 2 2
90 2 10 0 9 2 2 13 11 2 2 16 14 3 0 3 16 15 4 13 15 10 7 10 10 9 2 3 3 1 10 0 9 1 10 9 1 9 2 3 2 3 3 16 10 9 13 2 10 9 13 15 0 0 9 2 7 3 10 9 4 13 15 4 3 13 2 13 1 7 13 3 2 7 13 1 1 10 9 2 10 13 3 16 13 9 1 10 9 2 2
19 2 15 4 13 3 0 7 3 0 10 9 2 11 2 2 13 11 11 2
47 2 6 2 2 13 11 2 2 15 4 13 16 10 1 15 9 14 9 13 1 15 2 9 10 2 1 15 2 13 0 7 0 2 4 13 14 13 0 9 16 15 13 15 7 13 15 2
1 2
24 1 10 11 13 9 2 0 2 0 2 0 2 8 2 2 2 11 14 13 10 3 3 0 2
6 11 10 11 1 10 11
51 2 16 4 13 3 3 2 11 11 11 2 10 0 9 1 10 0 9 2 13 3 7 13 1 10 13 9 1 10 9 1 12 9 1 10 11 1 11 11 2 13 1 11 11 2 10 0 9 1 11 2
36 10 3 0 9 1 10 0 9 13 14 13 3 2 1 10 9 1 12 9 2 1 10 9 1 10 9 1 9 1 10 9 1 15 0 9 2
70 13 1 1 10 9 2 11 4 13 1 10 9 3 0 16 15 4 13 7 10 9 7 10 9 2 7 3 10 9 1 10 9 2 7 15 13 14 10 9 2 16 16 10 0 9 1 10 0 9 2 13 1 10 9 1 10 9 2 4 13 15 0 3 3 1 0 2 2 2 2
4 15 13 3 2
28 15 4 13 3 3 10 0 7 0 9 2 10 13 14 13 10 9 1 0 9 1 10 0 9 1 10 9 2
41 2 2 2 7 0 1 15 0 9 2 4 13 1 10 0 9 1 11 11 11 2 0 7 0 2 1 0 9 7 13 1 0 9 16 16 1 10 0 9 2 2
1 2
2 11 11
37 2 15 4 13 0 1 10 9 2 7 11 13 10 9 7 3 13 3 1 1 15 9 11 2 7 11 16 15 4 13 1 10 9 1 15 9 2
16 1 9 2 3 2 15 13 3 2 7 10 9 4 13 15 2
31 1 10 0 9 2 10 4 4 13 2 15 13 15 9 0 9 2 7 10 9 13 3 1 10 9 7 3 13 15 9 2
42 15 13 14 13 16 10 9 13 0 7 10 9 1 10 0 7 0 9 1 10 9 10 13 10 9 13 14 13 9 16 10 13 0 7 16 10 9 4 3 4 13 2
8 2 7 9 13 0 1 15 2
14 1 10 9 15 4 13 10 9 1 11 2 10 9 2
17 15 13 3 1 15 7 13 1 15 3 16 15 4 13 10 9 2
19 15 7 15 9 13 15 1 15 9 7 13 9 1 15 1 10 13 9 2
24 3 7 3 15 4 4 13 15 9 1 15 4 15 4 13 3 14 13 10 9 1 10 9 2
15 3 2 1 0 9 2 15 13 16 15 9 13 3 0 2
10 7 15 13 14 13 0 3 1 11 2
18 15 4 13 15 2 7 11 13 15 9 3 16 15 13 15 10 9 2
19 15 13 16 15 4 4 13 15 3 4 15 13 15 15 4 13 1 11 2
29 11 13 10 9 10 15 4 13 2 13 15 1 15 9 2 9 2 7 13 15 1 10 9 1 10 9 2 11 2
29 3 15 13 15 15 4 14 13 2 16 16 15 13 11 14 9 15 13 15 1 2 7 11 4 13 14 13 15 2
23 15 13 15 4 4 13 1 10 9 9 1 10 10 9 13 7 13 15 1 16 15 13 2
52 1 3 15 13 1 10 9 14 13 15 13 10 9 7 14 13 15 1 10 13 9 2 7 15 13 16 16 15 4 13 1 1 10 9 15 0 9 4 3 3 4 3 13 7 15 4 13 0 1 0 9 2
23 1 10 9 1 11 2 10 9 4 13 2 16 10 10 9 4 13 9 1 10 9 2 2
1 2
2 11 11
16 10 9 9 13 1 10 9 2 12 2 9 1 10 11 2 2
66 15 13 1 11 2 15 13 10 9 9 1 10 11 2 13 1 11 1 1 10 0 9 1 11 11 2 3 1 11 2 2 2 14 3 11 4 13 15 9 2 2 3 3 10 9 2 7 3 10 9 1 10 9 7 3 10 9 13 1 10 11 13 1 11 2 2
48 10 9 9 13 1 10 9 10 13 10 9 14 4 13 1 10 9 7 1 10 9 9 7 1 10 9 9 0 1 9 9 2 9 7 9 2 1 15 1 11 11 2 9 1 10 11 2 2
68 15 13 1 10 9 15 9 11 11 13 10 11 16 16 9 4 4 13 7 1 10 9 13 0 14 13 0 9 1 10 0 9 1 15 9 7 0 9 1 10 0 9 7 1 13 11 13 10 9 1 12 9 1 9 2 11 11 2 2 3 3 12 2 9 1 10 11 2
17 15 13 13 14 13 16 10 9 4 13 2 10 11 14 11 2 2
51 1 10 9 1 10 9 1 11 1 10 9 2 10 9 1 11 2 10 3 3 2 13 11 11 2 13 15 9 1 10 0 9 2 10 2 11 11 2 10 13 2 10 11 1 11 2 2 2 0 3 2
51 10 11 11 11 2 12 1 10 11 14 0 9 14 13 9 2 0 7 0 9 7 14 13 10 9 1 9 2 4 13 11 11 2 10 0 9 9 1 10 11 2 1 10 9 1 10 9 3 1 11 2
15 10 9 3 11 13 1 9 9 1 1 11 11 14 9 2
8 11 11 13 9 13 10 9 2
41 10 0 9 10 13 11 11 13 2 14 3 11 4 13 15 9 2 13 1 11 11 11 2 1 11 2 9 9 1 10 11 2 13 2 2 11 13 1 10 9 2
6 15 4 13 7 13 2
10 15 13 3 0 1 11 7 11 2 2
15 15 13 10 9 3 11 14 11 13 1 10 9 1 9 2
25 12 9 1 10 9 2 3 12 9 3 2 11 11 2 9 1 10 11 9 2 13 1 10 9 2
21 1 3 3 2 10 11 13 14 13 0 1 0 9 7 14 13 15 1 10 9 2
66 11 11 14 9 13 2 3 3 1 15 13 10 9 1 0 9 2 3 3 16 14 13 10 9 2 3 10 2 11 14 11 2 4 4 13 2 0 9 1 11 11 2 7 1 10 0 9 11 11 13 10 9 13 1 0 9 3 15 13 14 13 15 0 9 9 2
39 13 10 9 1 10 11 14 9 1 9 10 4 13 2 1 9 2 0 9 0 16 2 15 13 10 11 2 7 0 0 0 9 1 2 11 11 12 2 2
68 1 10 0 9 2 10 11 13 1 15 0 0 9 1 2 11 1 10 11 2 15 13 3 10 9 1 10 11 11 1 11 13 10 9 1 10 9 1 10 9 2 10 9 11 11 2 15 13 14 13 10 9 1 10 11 2 2 13 1 9 13 1 11 11 2 10 9 2
51 11 11 11 13 10 11 14 9 13 9 0 1 2 11 13 10 9 1 10 15 13 15 9 2 15 4 14 13 1 11 2 8 2 8 2 2 2 11 2 7 2 7 10 9 3 2 2 2 13 2 2
159 11 11 11 13 14 13 1 11 11 2 7 3 15 13 10 9 7 13 14 13 10 0 9 1 11 3 1 11 11 1 10 11 11 9 13 2 9 2 2 13 3 3 15 4 13 1 10 0 9 15 13 7 13 15 13 14 13 16 15 11 13 3 15 13 1 10 9 1 2 10 11 1 11 7 11 2 2 2 10 9 9 4 13 2 15 4 13 14 13 15 2 2 2 10 9 1 11 1 11 11 13 3 1 10 9 1 9 7 9 10 13 11 13 10 9 1 10 2 11 11 2 9 2 9 13 1 10 2 11 13 2 9 2 3 15 13 16 3 3 9 4 13 1 15 13 2 15 13 3 3 2 1 15 2 13 1 11 2 2
12 10 9 1 11 13 3 16 15 4 13 0 2
28 15 13 0 14 13 16 15 4 13 12 9 2 13 12 2 3 3 1 12 2 10 0 9 1 0 9 9 2
52 16 11 11 2 13 3 1 10 9 13 1 15 9 1 11 1 11 2 2 15 13 14 13 1 10 9 1 9 2 2 15 4 13 9 9 1 11 1 1 10 9 2 10 13 9 7 13 3 1 0 9 2
72 1 11 11 15 9 14 9 13 10 9 13 1 10 9 16 16 15 13 10 9 2 7 15 4 4 3 3 13 1 15 9 9 1 10 9 16 15 4 13 2 11 2 2 3 1 11 3 10 9 9 4 13 11 2 3 3 16 15 13 9 1 10 9 2 2 11 13 9 1 10 9 2
70 10 9 9 16 3 3 15 13 11 2 9 15 9 15 4 14 13 2 2 4 13 3 15 4 13 16 11 13 10 9 1 11 11 2 11 14 0 9 2 1 15 11 13 1 10 9 1 11 11 7 1 15 15 13 9 7 9 2 16 15 4 3 13 1 15 2 0 11 2 2
27 1 10 0 9 11 4 13 3 1 11 11 2 15 13 11 14 9 1 0 9 2 1 1 15 13 9 2
33 11 4 13 3 1 11 2 7 1 9 1 10 9 15 13 10 0 9 14 9 13 14 13 1 11 2 1 10 8 0 0 9 2
55 11 13 16 15 13 11 13 10 9 2 7 15 4 14 13 16 15 13 16 15 13 0 1 10 9 1 1 15 0 9 7 0 9 7 3 16 1 15 9 15 0 9 13 14 10 0 2 3 16 15 4 3 13 0 2
95 10 0 9 13 10 9 1 9 1 11 7 15 9 7 11 7 15 9 7 15 13 15 13 14 13 1 0 11 1 10 9 1 10 9 1 9 1 15 9 7 13 11 11 13 15 0 1 15 9 1 9 7 13 9 2 15 13 10 9 10 15 13 1 10 2 13 15 13 2 9 7 13 14 13 9 1 0 9 1 10 0 9 2 13 10 9 15 4 14 4 13 1 10 9 2
36 15 13 0 14 13 10 9 1 11 3 15 13 2 2 15 4 13 10 9 2 10 9 15 4 14 13 2 2 1 9 1 11 1 10 9 2
29 2 15 3 13 10 9 10 15 0 9 11 11 4 13 15 3 15 13 15 0 1 15 0 9 7 0 9 2 2
70 11 13 10 10 0 9 9 1 10 9 2 1 1 15 0 9 2 9 7 9 7 1 1 15 13 9 2 16 15 13 15 10 0 9 1 3 12 9 2 16 16 15 4 13 1 2 13 3 0 16 10 0 9 4 13 15 13 10 9 1 0 9 3 2 16 11 7 11 13 2
16 15 13 9 10 15 9 9 1 0 0 9 4 14 13 3 2
15 15 13 3 0 16 9 7 9 4 14 13 9 7 9 2
35 16 13 10 9 2 11 11 13 0 9 1 9 11 11 14 13 15 0 16 13 14 13 10 9 1 10 11 2 9 1 10 15 3 13 2
71 1 1 10 9 10 15 0 9 1 11 11 4 13 15 2 15 13 9 0 1 2 2 15 4 13 10 9 7 10 9 2 12 9 15 4 14 13 13 3 15 13 0 3 2 7 13 9 1 10 2 11 11 2 9 13 16 2 3 15 13 0 9 14 13 3 0 1 10 9 2 2
17 10 11 4 3 3 13 1 9 0 1 15 1 15 9 7 9 2
15 12 1 10 9 1 15 9 13 10 9 1 0 11 11 2
24 10 9 13 1 10 9 3 11 11 13 11 11 1 10 11 9 1 10 9 16 13 15 13 2
63 3 11 13 11 16 15 4 13 9 16 3 9 4 13 1 11 1 15 9 1 10 11 7 11 13 16 15 13 9 12 1 10 0 9 9 2 11 13 1 10 0 9 2 2 6 2 2 1 11 2 2 2 16 16 11 13 10 0 9 7 9 0 2
35 1 10 11 14 9 2 13 3 2 15 13 0 11 14 2 13 3 16 3 15 3 13 2 2 16 16 11 13 14 10 9 1 0 9 2
37 3 3 2 11 13 11 1 10 11 9 16 10 0 9 13 10 9 1 9 7 0 9 2 7 1 10 9 15 4 4 3 13 9 1 10 11 2
25 10 0 9 13 1 10 9 1 11 14 9 13 16 15 13 10 0 9 15 4 3 13 10 9 2
33 10 3 13 9 13 1 10 9 1 9 1 10 9 1 11 14 9 2 11 11 2 13 1 15 1 10 0 9 14 13 3 1 2
41 10 9 1 2 11 11 2 2 10 0 9 9 9 1 11 11 13 2 2 15 4 14 13 10 9 1 10 9 3 7 15 4 14 13 14 13 9 1 15 2 2
37 15 13 0 14 13 16 10 9 4 13 0 1 10 0 9 9 1 1 10 9 7 9 1 11 11 2 15 13 16 10 9 9 4 4 13 15 2
14 15 9 13 1 10 9 3 3 15 15 13 10 0 2
10 11 11 13 16 11 11 13 10 9 2
16 11 11 13 16 15 13 0 16 13 16 9 13 1 11 11 2
66 11 11 13 1 10 9 16 2 11 13 10 3 0 9 7 15 4 14 4 13 3 3 2 2 10 1 15 13 10 9 2 7 10 11 13 3 10 9 1 3 0 9 2 16 9 3 3 2 15 4 3 13 10 9 1 0 9 9 7 15 13 3 0 1 11 2
33 10 11 1 10 9 1 10 2 11 2 13 3 3 3 1 11 7 10 0 0 9 1 10 9 1 10 11 13 1 1 11 11 2
15 1 11 11 10 11 4 4 13 3 10 0 9 1 11 2
52 11 11 13 3 16 15 13 16 13 9 2 7 15 13 9 1 9 2 13 16 1 10 9 15 4 13 1 10 9 1 11 10 13 1 15 7 10 13 15 9 14 9 1 1 15 11 7 9 1 0 9 2
20 15 13 15 4 13 9 1 10 9 2 16 16 10 0 11 4 14 4 13 2
14 13 10 0 11 13 14 13 1 0 1 9 1 9 2
17 11 13 9 3 3 2 16 3 0 0 9 1 9 1 10 9 2
76 16 10 11 13 15 0 9 1 10 0 2 11 14 11 2 1 15 12 0 9 2 11 2 11 11 2 2 15 13 10 0 9 1 0 0 0 9 1 10 8 0 9 7 13 15 9 1 9 2 15 13 15 9 1 9 2 9 1 9 2 9 1 9 9 2 9 2 0 9 2 9 2 8 2 8 2
43 10 9 16 0 9 9 0 1 10 11 7 10 11 11 13 10 10 0 9 10 14 3 10 0 0 9 4 13 2 13 16 10 9 1 11 13 1 9 2 13 10 9 2
89 10 3 0 9 2 13 9 2 0 0 9 2 0 7 0 9 1 0 9 2 8 0 9 9 2 9 9 2 0 0 9 2 0 9 1 9 2 8 9 1 9 2 13 9 2 9 2 9 2 9 2 0 7 0 9 7 10 0 9 1 0 9 2 13 1 1 10 0 9 10 11 13 1 15 0 9 10 11 7 10 11 11 2 1 10 11 14 11 2
36 16 15 13 3 15 13 9 7 9 1 15 9 2 15 13 16 15 13 10 9 2 9 7 10 9 0 1 10 13 1 11 11 7 11 11 2
23 15 13 15 14 13 10 9 1 1 15 9 13 1 9 0 1 10 11 14 0 12 9 2
5 15 4 4 13 2
4 10 0 9 2
5 2 10 12 9 2
15 1 10 9 1 9 2 15 4 13 15 9 1 15 9 2
6 9 2 11 2 8 2
9 9 2 9 2 9 2 9 2 9
7 9 1 11 2 10 13 9
4 1 11 11 11
10 8 8 8 8 8 8 8 9 2 9
4 11 12 11 12
23 10 9 4 4 13 1 1 10 9 9 1 9 16 10 11 9 4 13 10 9 1 11 2
47 2 10 11 9 4 13 15 11 9 1 10 0 0 9 1 13 0 9 1 11 1 10 11 11 2 13 1 0 9 9 2 13 0 0 9 1 10 0 9 2 2 13 11 1 11 9 2
52 2 10 11 0 11 11 10 9 2 2 13 11 2 2 13 2 11 9 9 2 15 13 16 10 11 9 4 4 13 16 10 11 11 4 3 13 10 9 16 13 10 9 2 13 9 1 9 2 13 0 9 2
25 10 2 10 9 13 0 2 9 4 13 11 11 11 11 14 3 13 9 1 10 0 12 9 2 2
14 10 9 1 10 9 1 10 10 9 13 3 1 9 2
5 8 2 9 1 11
33 10 0 9 1 11 4 13 1 10 9 1 3 0 0 9 2 3 10 11 11 7 10 11 11 1 11 11 1 11 2 11 2 2
19 7 11 7 11 13 0 9 1 10 0 0 9 1 11 10 13 3 9 2
14 1 9 2 11 3 13 10 0 9 1 10 0 9 2
20 4 10 11 11 13 0 9 1 11 2 10 9 1 11 4 13 0 7 0 2
31 1 10 0 12 9 1 11 2 12 11 9 4 4 13 1 11 2 13 1 10 12 9 1 10 11 11 9 9 1 11 2
37 0 1 10 9 13 1 0 9 4 13 1 0 0 9 10 13 15 0 9 2 13 10 0 9 13 10 9 2 7 13 0 0 9 1 10 9 2
35 16 10 11 13 11 2 15 13 0 16 0 9 2 3 13 1 9 1 0 9 2 4 3 13 9 9 1 11 1 0 9 0 1 11 2
45 10 9 4 13 10 0 9 1 11 7 0 9 2 11 9 4 4 13 14 13 15 3 1 15 9 2 7 11 9 4 13 15 13 14 13 10 0 9 15 3 13 13 1 9 2
13 11 2 3 10 13 9 2 4 13 3 1 9 2
5 8 2 11 14 9
31 1 11 2 11 4 14 13 10 0 12 9 13 15 0 9 13 1 1 0 9 2 13 9 2 7 12 0 2 13 9 2
42 16 11 14 0 9 13 14 15 15 13 1 10 9 1 10 11 2 11 9 2 15 9 4 13 7 10 9 1 10 0 9 4 13 2 10 9 13 0 0 9 3 2
31 13 1 10 9 13 1 10 11 1 11 7 11 11 1 11 1 12 2 11 2 13 10 12 9 1 9 7 3 12 9 2
14 15 13 12 11 11 11 13 1 9 7 0 0 9 2
43 11 14 9 3 13 9 1 12 0 9 9 2 12 0 0 9 9 2 12 9 9 2 12 9 9 2 12 9 9 2 12 9 2 12 9 9 2 7 12 0 9 2 2
26 2 11 13 3 10 0 0 0 9 10 13 10 0 0 0 9 1 11 9 2 2 13 10 11 9 2
17 2 11 13 0 9 1 0 9 2 7 13 10 0 9 1 9 2
24 15 13 0 9 16 15 4 13 7 10 0 2 9 9 9 7 10 9 1 9 1 0 9 2
23 15 4 3 3 13 15 9 1 0 9 2 7 10 9 1 15 0 9 9 13 0 2 2
29 10 11 9 13 1 11 12 13 2 2 1 1 15 9 1 10 11 11 2 11 4 3 13 10 9 1 10 9 2
29 10 3 13 2 9 2 9 1 10 0 9 13 11 3 1 10 9 1 10 9 13 14 13 9 1 1 10 9 2
49 3 10 0 9 10 11 13 1 9 13 0 3 14 13 9 2 7 0 9 1 0 9 9 1 9 9 9 1 10 9 1 10 9 13 15 0 0 0 9 1 10 0 9 4 13 3 0 2 2
22 2 3 0 2 2 13 10 11 9 2 2 13 10 9 13 16 13 7 13 15 9 2
51 10 11 9 13 0 9 3 11 4 13 9 13 10 3 0 9 2 0 9 9 2 2 11 4 13 0 0 9 7 9 9 9 1 11 2 9 9 1 11 11 2 9 1 11 2 7 0 9 2 2 2
24 15 13 11 14 9 9 10 13 10 0 9 1 0 9 1 10 9 2 3 1 10 11 11 2
25 11 14 9 13 10 11 11 13 10 13 9 1 9 10 13 3 1 10 0 9 13 1 10 9 2
23 10 9 15 3 13 12 9 2 10 11 1 11 2 10 4 3 13 1 10 0 0 9 2
12 1 9 2 11 13 10 0 9 1 10 9 2
16 9 9 13 1 10 9 4 13 0 9 1 10 9 13 3 2
24 1 10 10 9 1 11 14 9 2 10 3 0 13 10 0 2 13 11 2 11 2 11 11 2
14 10 9 13 2 3 2 10 0 0 9 1 10 9 2
10 10 11 4 13 11 12 1 0 9 2
21 15 0 0 2 9 9 13 9 12 2 10 12 9 0 1 10 0 2 13 11 2
12 10 11 13 12 0 9 14 13 15 0 9 2
25 10 9 14 9 13 16 12 7 12 9 4 13 10 9 2 7 12 9 4 13 10 12 9 9 2
10 10 11 13 3 0 1 10 11 9 2
20 13 16 15 13 12 11 10 13 10 11 11 1 9 1 12 2 13 12 9 2
10 10 11 4 14 13 15 14 13 15 2
20 10 11 9 9 11 11 4 3 13 1 10 11 11 2 1 10 12 9 3 2
27 13 1 10 11 13 10 11 11 11 11 2 10 13 10 11 11 2 10 11 11 2 7 10 11 11 11 2
10 10 11 11 4 3 13 1 10 9 2
37 10 11 9 2 1 15 0 9 7 9 14 13 9 9 2 4 13 0 9 10 9 16 11 13 14 13 1 10 9 1 10 0 9 1 15 9 2
20 1 10 0 9 13 10 9 16 11 13 15 0 9 1 10 0 9 1 11 2
23 3 2 10 11 4 13 10 0 9 1 9 13 0 9 2 9 2 13 9 7 9 9 2
20 10 0 0 9 4 13 12 9 7 9 1 9 1 0 1 10 9 1 9 2
21 10 9 1 11 4 13 10 9 9 2 10 9 10 4 13 0 1 10 12 9 2
44 16 11 13 14 13 10 7 10 1 15 12 0 9 9 2 1 1 10 7 10 1 15 3 12 2 0 9 2 1 10 11 9 2 10 9 1 10 11 11 4 13 3 0 2
5 8 2 10 0 9
25 1 11 1 12 2 11 7 11 13 1 10 0 9 9 14 13 2 9 7 9 2 1 10 9 2
42 15 13 10 0 9 1 10 0 9 1 11 2 7 10 9 1 11 14 9 1 11 1 10 9 1 0 11 11 11 11 2 10 4 3 13 1 10 9 13 1 11 2
23 10 9 1 11 4 13 10 0 9 9 2 7 4 3 13 11 1 0 9 1 0 9 2
12 1 11 2 11 14 9 13 9 14 13 1 2
19 3 10 0 9 13 11 13 1 10 0 0 9 1 10 11 11 1 11 2
22 11 4 13 9 1 9 16 13 0 0 9 14 13 1 10 9 1 11 14 0 9 2
21 1 1 12 2 11 13 10 12 9 1 9 2 12 9 2 7 10 0 9 9 2
25 10 0 11 11 4 13 1 12 1 12 9 2 9 9 7 12 9 9 2 13 3 1 12 9 2
23 11 3 13 12 1 10 0 9 1 0 9 1 10 9 2 13 3 1 11 2 13 9 2
20 11 2 11 11 7 11 4 13 0 9 1 9 2 1 2 10 2 9 9 2
23 13 15 13 10 3 2 13 9 16 11 13 3 10 3 0 0 9 9 1 10 11 11 2
7 8 2 11 7 10 11 9
41 16 10 0 9 1 13 0 9 2 9 1 10 9 2 7 0 9 13 0 16 10 11 13 11 2 10 13 1 9 1 10 9 1 11 1 10 11 2 11 9 2
22 11 14 9 4 13 2 13 3 1 15 0 9 1 9 7 0 9 14 13 15 9 2
25 1 10 0 0 9 2 11 4 13 9 1 11 1 5 12 12 9 9 1 0 9 7 0 9 2
41 11 4 13 12 12 9 1 13 0 9 1 11 1 10 0 12 9 2 4 13 10 0 11 9 9 1 11 2 7 4 13 12 9 1 9 1 9 1 10 9 2
29 11 4 13 10 9 1 10 9 1 11 1 10 11 11 2 3 15 4 13 1 10 13 9 13 1 11 1 11 2
19 10 11 9 1 11 4 4 13 1 11 1 10 0 9 1 15 0 9 2
24 3 2 10 9 1 10 11 11 4 13 10 9 13 11 14 13 0 9 1 10 11 1 11 2
29 4 11 13 14 13 1 10 11 14 13 15 9 7 0 9 9 1 11 2 10 11 4 4 13 1 10 0 9 2
24 10 9 13 14 3 1 10 0 9 2 16 11 4 13 10 9 1 10 11 1 9 1 11 2
19 3 3 2 11 13 10 0 9 1 10 0 9 1 10 9 1 15 9 2
44 11 11 11 2 13 1 10 11 11 2 13 1 11 1 12 16 2 1 10 9 1 0 9 1 0 9 9 1 10 11 11 2 10 0 9 13 9 9 1 3 5 12 12 2
11 11 14 9 1 9 13 3 5 12 12 2
8 11 11 13 3 5 12 12 2
12 10 9 13 10 9 0 9 1 10 11 11 2
24 16 13 10 9 1 15 9 2 10 9 4 13 10 9 1 0 9 7 13 11 9 9 13 2
32 11 4 3 13 14 13 11 7 11 14 13 0 9 2 7 1 10 9 1 11 2 1 11 2 1 9 2 11 13 10 9 2
18 11 7 11 2 7 10 9 1 0 2 13 0 9 9 16 15 13 2
17 15 4 13 10 9 13 10 0 9 10 9 16 10 9 13 2 2
21 2 10 0 9 1 11 2 2 13 11 2 2 4 13 3 11 4 13 15 9 2
38 3 11 14 9 13 14 4 13 2 0 9 1 11 2 11 2 3 12 9 1 10 9 1 10 9 4 13 1 11 2 4 13 15 13 1 11 11 2
12 9 9 4 13 10 0 9 1 0 0 9 2
28 16 15 13 1 13 9 9 7 10 9 1 10 9 9 2 0 9 4 13 10 0 9 1 10 11 11 2 2
12 1 0 2 11 13 10 0 9 1 10 9 2
12 4 15 13 14 13 2 15 4 3 13 15 2
38 11 14 0 9 1 15 3 13 1 10 0 9 2 11 13 10 0 9 1 10 11 11 11 11 2 7 4 13 10 9 1 11 13 1 10 11 11 2
4 8 2 0 9
23 0 9 4 1 9 13 15 1 10 9 16 15 9 4 13 7 13 10 9 1 10 9 2
12 10 0 9 1 10 0 11 11 13 10 9 2
16 10 0 12 9 1 10 11 9 2 3 2 4 13 10 9 2
22 3 2 10 9 4 13 0 9 1 10 9 1 10 0 9 2 13 10 9 1 9 2
18 9 1 13 9 1 11 7 11 2 9 13 1 10 10 2 9 9 2
13 9 1 0 9 7 9 2 9 4 13 14 13 2
14 1 10 9 2 10 0 9 4 13 1 10 9 9 2
34 12 0 9 2 12 10 11 11 9 7 10 0 10 3 0 9 9 2 13 13 10 9 1 9 7 13 10 9 9 1 10 11 9 2
48 13 1 11 11 1 11 7 11 11 11 11 11 1 11 11 2 10 0 9 1 10 11 9 4 13 1 5 12 12 7 5 12 12 2 13 1 9 1 9 10 9 13 3 1 10 11 9 2
32 16 10 9 1 11 13 15 9 1 11 2 7 13 14 13 11 2 15 9 4 3 13 1 10 9 16 13 3 0 9 3 2
29 13 1 15 10 0 9 13 1 11 2 7 10 0 9 0 1 10 0 9 1 10 9 1 11 9 1 10 9 2
40 16 11 7 11 2 1 15 0 9 2 9 9 7 13 0 9 9 2 13 14 13 1 10 3 0 11 9 1 11 2 15 9 3 4 13 9 1 10 9 2
20 11 14 9 1 10 9 4 13 9 1 9 7 9 9 1 9 10 0 9 2
43 1 10 0 2 9 9 2 10 3 2 13 0 9 1 9 13 10 9 1 0 9 14 13 10 13 7 13 9 4 13 1 9 2 13 10 0 9 1 0 7 0 9 2
8 9 2 13 10 1 15 0 2
27 10 9 4 4 13 3 3 16 0 2 10 9 1 9 4 13 10 9 3 0 1 9 7 0 0 9 2
32 15 13 0 14 13 10 9 1 10 9 10 4 13 10 11 11 1 10 0 7 0 9 1 11 2 11 2 11 7 11 3 2
27 11 4 13 1 0 9 16 13 1 10 9 1 0 9 2 7 3 10 9 4 4 13 1 10 0 9 2
34 3 2 0 11 11 11 3 13 16 11 4 14 13 15 0 9 1 10 9 1 0 9 9 2 7 13 14 13 13 11 1 10 9 2
16 3 2 10 9 1 11 14 0 9 4 13 11 1 10 9 2
11 11 3 13 13 16 13 9 1 10 9 2
32 10 9 0 1 10 9 1 10 9 2 3 2 13 14 3 13 10 9 4 4 13 1 10 3 2 13 2 9 1 9 2 2
23 3 2 10 10 9 1 10 9 13 10 9 1 10 9 2 9 1 10 9 2 13 9 2
11 10 9 1 9 4 13 10 10 0 9 2
8 13 3 3 1 12 11 11 2
25 11 11 11 7 15 9 4 3 13 3 0 9 1 9 1 9 14 13 0 9 1 10 9 9 2
19 13 10 0 9 9 13 3 1 10 9 3 0 0 9 13 1 10 9 2
6 3 3 2 13 11 2
27 11 11 2 11 14 3 0 9 2 3 13 11 1 10 9 1 10 12 9 14 2 13 1 10 9 2 2
24 10 9 1 11 13 0 0 9 1 10 11 3 3 1 10 9 2 7 1 10 12 0 9 2
24 10 9 1 0 9 4 4 13 1 10 9 1 11 2 7 1 10 9 1 9 1 10 9 2
13 10 9 13 1 12 3 2 0 9 2 11 11 2
27 10 11 9 13 14 13 10 10 3 2 13 11 9 1 11 2 7 10 12 9 13 0 1 10 9 3 2
7 13 10 1 15 10 9 2
15 9 13 6 2 7 9 3 13 10 9 1 0 0 9 2
29 10 9 16 10 11 9 4 13 0 14 13 11 7 13 10 0 9 1 10 9 1 0 9 13 1 12 0 9 2
8 15 13 15 3 3 1 11 2
18 1 11 11 2 13 1 2 15 15 4 13 2 2 13 1 11 11 2
21 12 2 0 9 1 9 13 1 10 0 7 0 9 9 10 9 1 12 7 12 2
16 12 2 9 1 0 9 3 13 1 10 11 9 16 13 9 2
19 12 2 9 1 9 10 4 13 0 1 12 16 10 0 2 9 9 13 2
28 12 2 9 1 9 11 13 0 9 2 0 9 2 0 9 2 9 7 9 1 15 12 9 1 10 9 9 2
21 15 9 13 10 0 9 14 13 1 10 0 9 1 10 9 9 16 13 10 9 2
27 12 2 9 1 9 13 1 0 9 1 10 11 14 12 2 9 2 9 9 1 10 9 2 13 1 12 2
36 12 2 9 1 9 16 13 9 3 11 13 3 14 13 10 11 11 2 10 0 9 14 13 9 9 1 3 12 9 9 1 12 9 1 12 2
13 10 11 11 13 14 13 15 9 1 12 9 9 2
15 12 10 9 1 10 11 11 3 1 9 1 9 9 9 2
16 12 2 9 1 0 0 9 9 9 10 11 11 13 0 1 2
24 12 2 9 1 9 16 13 9 3 11 13 1 15 9 9 14 13 9 9 9 1 9 9 2
34 12 2 9 9 9 9 4 13 1 10 0 12 9 1 11 14 0 0 2 9 9 2 10 9 1 12 9 9 1 15 12 9 2 2
25 12 2 9 1 9 10 11 9 13 1 12 16 0 9 4 4 3 13 16 0 9 4 4 13 2
32 5 12 12 2 9 10 11 2 11 12 9 7 10 11 11 11 13 1 9 1 10 9 9 2 9 2 9 2 7 9 9 2
20 12 2 9 1 9 9 13 7 13 0 9 1 11 14 0 12 9 1 9 2
39 12 2 9 1 11 9 9 15 13 9 1 10 9 9 2 13 12 9 9 2 10 12 3 0 11 11 9 2 7 0 1 12 0 0 2 9 9 2 2
49 12 5 0 9 1 9 9 7 9 9 0 1 10 9 10 4 4 13 1 10 11 9 1 11 1 12 9 2 10 9 10 13 15 3 3 0 16 9 9 14 13 10 9 1 10 0 0 9 2
17 12 2 9 9 1 11 11 11 9 9 1 9 1 11 14 9 2
15 12 2 9 9 1 0 9 1 0 9 16 11 13 9 2
15 12 2 9 9 1 0 9 1 0 9 16 11 13 9 2
20 5 12 12 2 9 10 11 3 13 10 0 9 3 13 0 9 1 13 9 2
22 5 12 12 2 9 10 11 13 10 0 9 3 13 9 1 13 9 1 10 11 9 2
21 12 2 9 1 9 1 11 14 12 2 9 11 11 11 1 9 1 0 9 9 2
15 12 2 9 1 9 13 14 13 11 14 11 11 11 9 2
20 12 2 9 1 9 1 12 11 3 11 14 11 11 11 13 11 14 9 9 2
12 12 2 9 1 10 9 14 9 10 13 0 2
12 12 2 9 1 10 9 14 9 13 1 11 2
12 12 2 9 1 10 9 14 9 10 13 0 2
12 12 2 9 1 10 9 14 9 13 1 11 2
16 12 2 9 1 9 10 11 11 13 1 12 2 10 0 9 2
17 12 2 13 9 1 0 9 10 4 13 1 11 14 11 11 9 2
17 12 2 9 1 11 11 11 9 1 10 9 2 9 9 1 12 2
23 12 2 9 1 0 9 10 11 9 2 10 9 14 0 9 2 13 1 10 9 10 9 2
28 5 12 12 2 9 1 10 11 9 9 1 0 9 9 2 9 1 12 2 10 9 2 9 13 2 9 13 2
21 5 12 2 9 1 0 9 1 10 11 9 9 1 0 9 9 2 9 1 12 2
27 12 2 13 9 1 9 9 13 0 9 1 0 2 9 9 10 13 0 1 10 0 9 1 10 11 9 2
18 12 2 9 1 10 9 10 11 3 13 14 13 10 9 14 13 3 2
29 12 2 9 1 13 9 1 11 11 15 3 13 1 0 2 9 9 9 2 3 9 1 15 4 14 13 9 9 2
15 12 2 9 1 9 1 11 11 15 3 13 1 9 9 2
20 12 2 9 1 9 1 11 11 15 3 13 1 9 2 9 2 7 9 9 2
36 12 2 9 9 1 11 11 13 12 9 0 1 10 9 1 11 2 11 2 3 10 11 11 11 9 13 12 1 10 0 11 9 1 11 9 2
26 12 2 9 1 11 9 0 9 1 0 9 13 1 12 11 12 7 12 11 12 10 13 11 2 11 2
24 12 2 9 1 11 9 0 9 1 0 9 7 9 1 10 0 9 10 13 11 7 11 11 2
22 12 2 9 1 11 9 0 9 1 0 9 7 9 1 10 0 9 10 13 9 9 2
24 12 2 9 1 11 9 0 9 1 0 9 7 9 1 10 0 9 10 13 9 1 0 9 2
19 12 2 9 1 9 11 13 11 11 11 1 15 12 9 1 10 9 9 2
20 12 2 9 1 9 3 11 13 9 7 9 1 15 12 9 1 10 9 9 2
27 12 2 9 1 9 11 13 11 2 11 2 7 9 2 1 1 9 2 1 15 12 9 1 10 9 9 2
37 5 12 12 2 13 9 1 10 9 10 11 11 11 1 11 11 2 11 2 13 1 11 11 2 11 11 14 9 1 10 11 11 7 11 9 9 2
18 12 2 9 1 9 11 13 11 11 1 15 12 9 1 10 9 9 2
20 12 2 9 9 1 12 7 12 1 0 0 9 1 0 9 1 10 11 11 2
14 12 2 9 1 10 12 11 9 15 13 1 11 11 2
22 12 2 9 1 12 11 9 15 9 9 13 1 0 11 2 0 2 11 11 2 9 2
24 12 2 9 1 11 2 13 9 1 10 11 11 9 2 13 1 11 11 3 3 1 12 11 2
33 12 2 9 1 11 7 11 11 2 11 2 9 13 14 13 1 12 13 0 9 1 10 11 11 1 9 3 11 2 11 13 0 2
22 5 12 12 2 9 10 11 11 13 0 14 13 10 12 9 14 13 10 12 11 9 2
15 5 12 2 11 13 1 11 11 14 13 0 11 0 9 2
15 5 12 12 2 9 11 13 1 10 11 14 13 9 9 2
18 5 12 12 2 9 13 1 10 9 10 13 1 10 11 9 9 9 2
16 5 12 12 2 9 10 12 0 9 4 13 14 13 13 9 2
20 12 2 9 1 11 9 13 1 10 11 9 1 9 7 9 12 16 13 0 2
5 11 11 2 0 9
29 12 2 9 3 11 13 3 1 15 9 9 1 10 11 11 11 2 3 12 9 16 15 12 2 9 9 13 3 2
22 5 12 2 9 10 9 1 9 13 1 12 1 9 15 4 13 11 14 11 9 9 2
17 12 5 12 2 9 1 9 15 13 1 11 14 9 1 10 9 2
19 12 2 9 1 9 1 10 9 15 13 3 1 9 1 11 14 9 9 2
69 12 2 9 1 9 3 11 11 2 11 2 11 11 11 2 10 11 11 2 11 11 2 10 9 9 11 2 11 11 2 10 0 9 1 10 11 11 11 2 11 11 2 7 10 11 11 11 1 11 2 11 11 2 10 0 9 1 10 9 1 11 2 13 1 9 2 13 2 2
25 12 2 9 1 0 0 7 11 9 9 15 13 10 9 15 13 0 9 9 13 1 9 1 11 2
22 12 2 9 1 9 1 10 11 11 7 11 1 11 15 13 10 9 13 1 10 9 2
31 12 2 9 1 9 10 10 11 13 13 10 9 15 4 13 10 11 2 10 9 2 1 10 9 1 10 9 1 10 9 2
20 12 2 9 9 1 9 1 12 7 12 1 11 11 9 2 9 14 9 2 2
2 0 9
18 12 2 9 1 9 10 11 11 4 13 7 13 1 16 13 1 9 2
25 12 2 0 9 1 9 2 1 1 10 9 1 12 13 1 10 11 11 2 1 10 11 0 9 2
17 12 2 9 1 10 0 9 14 0 9 10 10 11 13 1 9 2
15 2 15 13 1 12 2 10 9 1 10 9 1 11 2 2
10 5 12 12 2 13 0 9 1 12 2
3 9 1 11
31 12 2 10 9 1 10 11 11 2 11 11 14 0 9 1 10 11 11 2 13 11 11 10 9 1 0 9 1 10 9 2
31 12 2 9 1 9 16 11 13 16 11 11 11 13 10 9 1 10 12 11 9 3 15 13 1 9 14 2 13 2 11 2
29 12 2 0 9 1 0 9 1 11 13 1 0 11 9 9 1 12 7 11 12 2 13 1 10 11 11 11 11 2
34 12 12 2 13 9 1 9 3 15 13 1 10 9 1 12 11 12 2 1 9 1 10 9 1 11 2 10 0 0 9 1 9 9 2
22 5 12 12 2 13 0 9 1 11 0 9 1 11 13 1 10 11 11 1 11 12 2
23 5 12 12 2 0 0 9 1 10 11 0 9 1 11 13 1 11 1 11 11 1 12 2
21 5 12 12 2 9 1 10 9 13 1 10 0 9 14 13 10 9 9 1 11 2
31 5 12 2 9 10 0 9 13 2 13 11 14 13 9 2 14 13 10 0 9 2 16 9 13 10 0 9 16 13 15 2
26 12 2 9 3 11 13 15 9 1 9 1 11 9 9 9 13 2 15 4 14 13 9 1 11 2 2
16 5 12 12 2 0 9 1 9 13 1 11 1 11 7 11 2
14 5 12 12 2 13 9 1 11 9 9 13 1 11 2
12 5 12 12 2 9 1 11 11 9 1 11 2
20 5 12 12 2 9 10 9 7 15 9 4 13 14 13 1 10 12 0 9 2
30 12 2 9 1 9 1 10 10 11 11 13 0 9 16 15 13 14 13 9 13 11 9 1 9 1 10 11 11 11 2
17 12 2 9 1 11 14 0 9 1 9 1 0 9 1 0 12 2
17 12 2 9 1 11 14 0 9 1 9 1 0 9 1 0 12 2
14 12 2 9 1 10 0 9 15 13 0 1 10 9 2
16 12 2 9 1 10 0 9 15 13 0 10 9 1 10 9 2
17 12 2 9 1 0 9 9 1 11 1 10 11 9 1 11 12 2
22 12 2 9 9 1 11 9 1 11 1 11 12 2 10 9 9 9 2 3 2 13 2
20 12 2 9 1 9 1 0 9 13 3 10 10 11 9 4 13 14 4 13 2
21 12 2 9 1 0 9 1 10 13 0 10 11 4 13 1 10 9 1 10 9 2
5 10 9 14 0 9
30 12 2 9 1 9 1 11 12 9 1 9 1 10 9 3 1 11 9 2 13 14 13 10 9 1 10 11 2 12 2
15 5 12 12 2 13 9 16 13 10 12 9 1 11 9 2
18 12 2 9 1 9 9 10 9 9 13 4 14 13 3 1 9 12 2
19 12 2 9 1 9 10 13 0 9 1 10 0 9 9 13 14 13 0 2
31 12 2 9 1 11 1 11 14 13 1 9 0 16 13 11 2 12 9 7 13 1 9 9 7 9 1 10 9 1 12 2
4 13 10 9 0
18 5 12 2 0 9 13 1 9 3 1 10 0 9 1 9 9 9 2
14 5 12 2 9 13 1 9 1 9 9 1 11 11 2
21 5 12 2 9 13 1 9 1 9 9 1 11 2 11 2 11 11 14 9 9 2
12 5 12 2 9 13 1 9 1 11 11 9 2
12 5 12 2 9 13 1 9 1 11 11 11 2
23 5 12 2 9 13 1 9 1 11 11 2 11 2 9 1 11 11 2 11 14 9 9 2
35 12 2 9 1 12 9 13 1 10 11 11 1 11 1 0 12 10 13 3 14 13 10 9 1 0 9 9 9 1 15 0 2 9 9 2
25 12 2 9 1 0 11 9 1 10 9 1 12 10 10 11 11 11 13 4 14 3 13 9 3 2
16 12 2 9 1 9 13 0 9 10 13 1 11 11 10 9 2
19 12 2 13 9 1 11 9 9 10 4 13 2 13 9 13 1 9 9 2
15 12 2 9 1 0 9 10 13 1 10 11 11 1 9 2
11 12 2 9 1 10 9 13 1 0 9 2
16 5 12 12 2 13 9 14 13 3 11 9 1 10 0 9 2
12 5 12 2 9 11 13 1 9 9 1 12 2
16 5 12 12 2 9 10 11 9 4 13 1 9 9 1 12 2
12 12 2 9 1 0 0 9 1 10 11 11 2
22 12 2 9 1 11 0 9 3 10 9 9 4 13 10 9 1 0 1 12 12 9 2
31 12 2 9 1 0 9 7 9 1 2 9 9 2 13 1 10 11 1 11 11 10 4 4 13 7 13 1 12 11 12 2
7 13 10 9 3 1 10 0
18 5 12 12 2 0 9 1 10 9 1 11 14 0 12 2 9 9 2
19 12 2 9 1 11 0 1 11 14 0 12 9 1 0 9 7 9 9 2
25 5 12 2 0 9 9 1 11 14 9 13 1 12 1 10 9 1 9 1 0 9 7 9 9 2
37 12 2 9 1 0 9 1 10 11 0 9 11 7 11 10 11 4 13 1 0 9 2 13 10 11 11 11 11 11 11 7 11 9 11 11 2 2
18 12 2 9 1 11 14 0 12 9 15 3 13 1 15 9 14 9 2
7 10 9 1 10 9 1 9
20 5 12 12 2 9 1 0 0 9 10 11 2 11 12 9 13 2 10 9 2
29 5 12 12 2 9 1 0 9 13 1 10 11 9 2 10 0 9 2 9 9 13 1 10 11 2 11 12 9 2
23 2 9 13 14 13 3 3 5 12 16 13 3 9 1 1 1 5 12 1 9 7 9 2
25 9 4 13 9 2 10 4 13 1 10 9 2 13 10 9 14 13 9 16 15 13 3 0 2 2
5 11 11 2 9 9
18 12 12 2 9 1 9 10 4 13 1 11 14 0 12 9 1 9 2
15 12 2 10 0 9 1 0 9 1 10 9 1 10 9 2
20 5 12 12 2 10 11 9 9 1 12 2 10 0 1 9 1 10 0 9 2
21 5 12 12 2 13 0 9 13 1 10 9 1 10 9 3 11 13 9 1 12 2
10 5 12 12 2 11 0 9 1 9 2
5 11 11 2 9 9
22 12 2 9 1 0 9 1 11 12 15 13 15 4 13 10 9 1 11 14 9 9 2
23 12 2 9 1 9 9 10 4 13 1 10 0 12 9 9 1 0 9 3 3 13 1 2
22 12 2 9 1 11 1 11 12 15 13 16 15 9 4 3 13 3 16 11 13 9 2
31 12 2 9 1 0 9 15 4 13 0 1 5 12 1 15 12 0 9 1 10 9 1 12 9 1 0 9 7 9 9 2
12 5 12 2 9 11 15 13 1 9 1 12 2
2 9 9
11 12 12 2 9 1 11 0 1 11 12 2
19 12 12 2 9 1 11 15 13 15 9 1 0 12 9 1 10 11 9 2
15 12 12 2 9 1 9 13 1 11 14 12 9 1 9 2
4 9 1 10 0
20 12 12 2 9 1 11 13 1 10 9 9 2 12 1 12 1 10 9 2 2
15 12 12 2 9 1 9 1 10 9 7 3 13 1 0 2
22 12 12 2 9 1 11 10 10 9 13 1 2 9 0 2 2 1 0 9 2 0 2
23 5 12 12 2 9 13 1 10 0 9 10 13 9 1 0 9 16 15 4 13 15 9 2
20 12 2 9 1 9 1 10 11 11 13 1 10 0 12 9 9 1 10 9 2
18 12 2 9 1 9 1 11 13 1 10 0 9 8 9 1 10 9 2
6 11 11 7 15 0 9
17 5 12 12 2 9 1 11 9 2 13 10 0 9 1 11 9 2
21 5 12 12 2 9 11 9 11 11 13 1 9 9 9 1 10 12 2 9 9 2
19 5 12 12 2 9 11 13 16 13 15 11 9 3 16 10 9 13 0 2
21 5 12 2 9 10 11 9 13 11 1 12 9 1 15 0 9 1 10 12 9 2
31 12 2 9 1 9 1 9 1 11 14 9 7 11 2 15 10 11 13 2 11 11 2 2 3 3 4 13 1 10 9 2
4 11 11 2 9
17 12 2 0 9 1 9 11 13 13 0 9 9 16 9 1 11 2
13 12 2 9 1 0 0 9 3 11 13 1 9 2
15 12 2 9 1 0 0 9 1 12 9 1 10 11 9 2
24 12 2 9 1 10 5 12 12 11 13 14 13 9 1 11 10 4 13 1 9 2 3 9 2
3 10 0 9
22 12 2 9 1 13 11 2 11 9 10 10 11 11 13 4 13 1 11 11 2 11 2
11 12 2 9 1 9 1 10 9 1 11 2
28 12 2 9 1 9 9 4 13 2 13 2 7 13 14 13 0 9 2 9 2 7 9 1 15 9 1 11 2
12 12 2 9 1 13 9 9 1 11 11 9 2
18 12 2 9 1 9 1 9 4 13 1 9 1 11 14 0 0 9 2
5 10 9 2 0 9
25 12 12 2 9 1 11 1 9 9 1 10 9 1 12 2 0 1 12 9 9 1 10 9 2 2
19 12 12 2 9 1 11 15 13 15 9 9 1 11 14 0 9 1 9 2
5 9 9 1 10 11
24 12 2 9 1 0 2 9 9 13 1 10 11 11 14 13 10 9 1 10 11 3 1 12 2
21 12 2 9 1 0 2 9 9 13 1 10 11 11 14 13 11 9 3 1 12 2
46 12 2 9 1 10 11 11 1 9 13 14 13 10 0 9 1 9 9 13 1 10 12 11 11 11 9 2 11 2 11 2 7 11 11 4 13 3 0 2 11 4 13 3 0 2 2
17 5 12 12 2 9 10 11 11 13 1 0 9 7 9 1 12 2
17 5 12 12 2 9 10 11 11 13 1 0 9 7 9 1 12 2
17 12 2 9 1 11 15 13 10 0 9 1 10 11 11 1 12 2
4 0 2 9 9
22 12 2 9 1 11 15 13 1 10 9 11 4 13 15 9 1 11 1 12 11 12 2
22 12 2 9 1 11 15 13 1 10 9 11 4 13 15 9 1 11 1 12 11 12 2
23 12 2 9 1 11 15 13 1 10 9 11 4 13 15 9 1 11 1 12 11 2 12 2
22 12 2 9 1 11 15 13 1 10 9 11 4 13 15 9 1 11 1 12 11 12 2
21 12 2 9 1 11 15 13 1 10 9 11 4 13 15 9 1 11 1 11 12 2
10 3 0 10 0 16 15 4 13 14 13
24 12 2 9 1 9 9 11 13 1 11 12 2 10 3 2 0 9 1 10 9 1 11 9 2
7 2 9 9 11 11 2 2
13 12 2 9 1 9 9 10 0 11 13 10 9 2
34 12 2 9 1 9 9 11 13 1 11 12 2 10 9 15 13 10 12 11 0 0 9 13 2 11 11 11 0 14 13 11 9 2 2
45 12 2 9 1 9 11 4 13 10 7 9 1 15 9 3 1 10 11 11 1 15 9 1 11 2 11 2 15 9 14 9 1 11 2 11 2 7 11 11 1 1 12 11 12 2
8 10 9 3 15 13 1 10 9
26 12 2 9 1 9 9 1 15 0 12 9 1 9 1 10 11 13 1 9 16 13 2 9 2 9 2
4 9 1 15 9
13 12 2 9 1 9 10 13 10 11 9 9 9 2
32 12 2 9 1 9 13 1 10 12 9 9 10 4 13 1 11 11 7 11 2 10 0 9 2 9 9 2 10 0 0 9 2
21 12 2 9 1 9 10 4 4 13 1 9 9 9 10 4 14 13 10 9 9 2
23 12 2 1 12 11 12 2 10 11 13 10 9 16 4 13 11 11 4 3 13 1 12 2
21 5 12 12 2 9 13 1 10 11 2 11 12 9 2 10 0 1 0 0 9 2
22 5 12 12 2 9 13 1 10 11 2 11 12 9 9 2 1 10 9 1 11 12 2
19 5 12 12 2 9 10 10 11 2 11 12 9 13 14 13 1 11 12 2
26 12 9 1 11 2 11 9 2 9 15 4 13 9 9 2 16 13 5 12 10 2 1 1 11 12 2
27 12 2 9 1 11 2 11 9 2 9 15 4 13 9 9 2 16 13 5 12 10 2 1 1 11 12 2
20 5 12 12 2 10 9 9 7 9 4 13 1 11 2 11 1 1 11 12 2
17 12 2 9 1 11 15 4 14 13 10 11 11 1 10 11 11 2
27 12 2 9 1 11 15 13 10 11 11 14 9 1 11 12 16 11 11 13 3 0 1 10 12 11 9 2
23 12 2 9 1 11 15 13 1 11 12 16 11 14 2 9 1 0 9 2 4 4 13 2
20 12 2 9 1 11 15 13 1 11 12 16 11 4 13 15 9 1 11 9 2
21 12 2 9 1 0 0 9 15 4 14 13 11 2 11 2 7 11 1 10 9 2
18 12 2 9 1 0 0 9 15 4 14 13 10 11 11 1 10 9 2
18 12 2 9 1 0 0 9 15 4 14 13 10 9 1 10 11 11 2
18 12 2 9 1 0 0 9 15 4 14 13 10 9 1 10 11 11 2
18 12 2 9 1 0 0 9 15 4 14 13 10 11 11 1 10 9 2
19 12 2 9 1 11 15 13 16 2 9 7 9 13 3 0 14 13 2 2
5 10 9 1 15 9
32 12 12 2 13 9 1 11 15 13 15 1 11 15 13 11 11 1 15 0 9 7 15 13 10 11 1 10 0 9 1 11 2
13 12 12 2 9 1 11 15 13 1 11 1 12 2
15 12 12 2 9 1 9 1 0 15 13 1 11 1 12 2
14 12 2 9 1 9 15 13 15 1 13 2 3 11 2
20 12 2 9 1 9 10 4 14 13 10 9 2 9 2 1 0 9 9 9 2
7 15 9 3 4 14 13 2
14 6 15 9 13 3 0 2 15 3 4 14 13 9 2
22 15 13 12 9 7 3 13 15 9 2 15 13 10 0 9 1 10 9 1 12 9 2
26 3 15 13 10 0 7 15 3 13 15 9 3 3 15 10 13 15 7 15 13 15 13 10 0 9 2
30 15 13 3 1 2 6 15 4 13 3 0 14 3 13 15 2 15 13 15 13 15 2 2 7 15 4 14 3 13 2
17 15 13 3 13 1 10 9 1 3 0 9 4 13 15 13 0 2
12 6 2 10 9 4 3 13 1 15 2 9 2
33 4 14 13 15 6 2 15 13 0 7 13 14 13 15 9 1 10 1 15 14 13 1 15 2 6 13 7 9 16 15 13 9 2
11 15 13 0 1 15 2 15 13 10 0 9
6 0 9 11 13 9 2
21 4 9 13 15 10 9 10 9 10 4 13 12 2 9 7 9 13 2 1 7 2
5 0 9 2 9 7
2 0 9
15 10 9 13 9 1 11 1 16 15 15 13 1 9 9 2
18 11 11 2 15 13 3 1 10 9 0 9 2 13 9 1 0 9 2
14 15 0 9 13 14 13 1 11 7 13 10 9 9 2
7 11 11 1 11 1 11 2
6 11 11 1 11 2 11
29 11 11 2 15 13 15 13 10 9 2 7 16 15 13 15 3 15 4 13 3 1 10 0 9 2 2 1 11 2
20 13 1 10 11 9 2 13 1 9 9 7 13 1 10 9 15 13 14 13 2
27 15 4 13 15 10 0 9 1 10 10 9 10 13 10 9 15 13 2 7 10 10 9 15 13 14 13 2
12 1 1 11 2 15 0 13 10 11 0 1 2
2 0 9
79 15 4 14 13 10 9 15 13 0 2 16 15 13 15 15 9 13 1 11 15 4 13 2 13 9 0 13 15 13 0 3 1 1 10 9 15 13 15 2 10 9 15 13 7 13 9 2 7 10 9 15 13 2 3 16 15 4 14 13 0 2 0 9 3 1 10 0 9 1 11 2 11 2 11 11 2 7 11 2
34 1 9 11 13 0 14 13 9 1 10 9 15 13 15 14 11 7 13 10 11 14 13 1 10 9 16 15 13 10 9 1 10 9 2
37 15 13 14 4 13 1 10 9 7 16 15 13 14 3 15 4 4 13 13 10 9 14 13 15 9 2 16 15 4 13 1 10 0 9 9 1 9
8 13 10 9 9 1 10 9 2
10 4 15 13 13 1 11 1 10 9 2
34 15 4 4 13 10 9 14 13 1 11 2 11 2 0 9 1 9 1 15 9 2 16 15 13 1 11 2 15 13 10 9 7 9 2
9 7 4 15 13 15 1 10 9 2
21 10 11 13 3 0 1 11 2 7 3 10 9 15 13 9 1 11 3 13 3 2
19 11 13 10 0 9 9 2 15 13 9 3 2 15 4 4 13 1 9 2
12 1 9 2 15 3 4 14 3 13 14 13 2
6 11 13 15 1 12 2
19 16 15 13 2 0 9 2 13 1 9 1 11 2 7 3 1 10 9 2
44 11 13 10 10 0 9 2 9 2 9 9 2 9 9 2 0 9 2 15 13 3 1 12 9 3 1 9 2 7 11 13 15 3 3 2 15 4 14 13 2 7 4 15 2
6 15 13 3 15 9 2
11 15 11 11 13 1 0 9 9 15 13 2
5 4 15 4 13 2
16 15 3 13 10 11 2 7 10 9 13 3 3 10 12 9 2
13 7 15 4 14 3 13 10 0 9 1 9 9 2
14 14 1 10 9 2 16 15 13 15 9 16 13 0 9
19 15 13 0 14 7 13 1 10 9 9 2 7 13 12 10 4 14 13 2
5 11 11 4 13 2
7 4 15 13 13 9 9 2
8 13 10 0 9 1 11 11 2
14 3 15 4 13 10 0 9 1 11 11 7 11 11 2
8 10 9 13 1 9 7 9 2
11 7 15 4 3 13 10 9 9 9 9 2
9 15 4 13 11 11 7 11 11 2
13 15 13 3 0 7 13 1 10 9 10 10 9 2
21 1 10 11 11 9 15 13 10 9 13 3 0 7 15 13 10 9 13 10 9 2
6 13 15 13 1 15 2
12 13 10 9 7 9 1 11 10 0 0 9 2
6 7 3 0 13 15 2
4 15 13 12 2
27 15 4 3 13 1 10 11 9 7 9 3 3 2 15 4 13 10 9 1 10 0 9 1 15 9 9 2
21 3 15 13 11 1 11 2 0 9 2 15 13 10 0 9 15 13 10 11 9 2
8 4 9 13 15 9 1 15 2
59 15 4 13 0 7 0 2 3 3 0 2 3 0 1 9 1 9 9 9 9 2 9 9 7 9 2 1 3 1 10 9 9 15 13 0 9 2 3 10 9 1 10 9 13 10 9 14 13 3 7 9 14 13 10 9 1 10 9 2
17 10 9 13 15 9 7 0 9 7 10 9 15 13 1 13 9 2
26 15 4 3 13 3 0 3 10 0 9 13 3 2 7 15 13 9 1 0 9 7 0 9 1 9 2
18 15 13 10 0 9 9 10 13 3 0 1 15 0 9 1 10 9 2
13 15 9 13 3 0 1 15 0 9 1 10 9 2
13 15 13 14 13 12 9 7 13 10 0 7 13 2
22 3 4 15 13 1 15 14 13 1 15 12 9 2 13 9 2 7 13 3 7 3 2
41 13 1 10 9 1 9 7 16 15 13 10 9 9 2 15 13 1 10 9 3 15 13 15 13 9 2 13 15 1 10 9 7 13 1 15 9 14 13 15 13 2
27 16 15 13 1 10 9 3 1 10 9 15 4 13 15 1 7 10 9 13 0 14 13 15 1 10 9 2
52 13 15 1 10 9 1 9 2 13 15 9 1 10 9 1 10 9 7 13 15 9 3 2 13 13 15 16 15 13 1 10 9 13 10 0 9 0 9 2 16 15 4 13 0 9 14 13 0 7 0 2 9
8 15 0 11 11 0 9 2 2
44 6 9 2 3 13 15 9 1 15 0 11 11 0 9 2 6 2 15 3 13 14 13 12 1 11 2 7 3 2 13 1 13 11 11 1 15 9 2 4 9 3 13 15 2
7 3 13 15 9 1 15 2
12 13 15 10 0 9 1 0 2 0 9 9 2
6 15 1 15 9 9 2
9 13 15 0 1 11 9 7 14 2
14 15 13 12 8 9 9 2 9 12 5 0 0 9 2
11 15 9 7 9 4 4 3 13 2 9 2
19 11 11 2 12 12 9 0 9 13 9 7 4 13 10 9 1 0 9 2
9 15 13 3 0 0 1 10 9 2
5 15 13 3 0 2
10 10 0 9 1 10 0 9 7 9 2
17 15 9 13 16 15 4 14 13 9 9 3 2 15 13 1 11 2
11 13 15 11 1 9 16 13 3 3 6 2
6 0 9 1 15 9 2
44 3 13 14 13 2 15 13 10 11 9 2 15 4 13 3 16 15 13 15 9 9 6 3 12 5 12 9 2 15 4 13 10 0 9 2 13 15 9 0 1 15 9 9 2
2 9 2
3 7 15 2
14 6 13 15 2 7 15 4 15 13 14 13 10 9 2
5 7 15 13 0 2
11 13 15 0 15 13 14 9 1 10 9 2
11 13 10 9 1 0 9 7 13 9 1 9
29 13 10 9 1 10 3 0 9 9 0 1 10 9 13 0 9 7 0 9 15 13 2 8 13 1 10 9 1 9
19 15 4 13 1 10 9 16 15 13 9 16 15 4 13 10 0 9 1 9
7 9 13 14 13 10 9 13
35 15 4 13 10 9 9 9 1 10 9 10 4 13 0 1 15 2 0 9 13 10 0 0 7 13 9 2 10 3 13 1 1 0 9 2
1 11
6 11 11 0 9 9 2
48 16 15 13 1 10 0 9 9 14 9 7 15 4 13 4 15 13 14 13 9 1 10 0 9 1 15 9 1 15 9 7 4 15 13 1 0 9 16 15 4 14 13 9 1 15 0 9 2
21 15 4 13 10 9 1 10 11 9 9 7 4 14 13 10 9 2 4 9 13 2
10 13 1 10 9 4 13 2 15 0 9
14 15 4 13 0 7 15 4 14 13 2 4 13 9 0
11 15 13 1 10 9 1 15 0 9 9 2
17 15 9 4 13 16 7 3 15 4 13 14 13 1 10 0 9 2
22 16 15 9 4 14 13 15 16 13 10 9 1 11 11 3 15 4 13 1 10 9 2
33 15 3 13 16 15 13 10 9 1 9 7 16 15 4 3 13 1 11 11 7 13 10 9 1 15 9 14 13 15 0 9 9 2
15 1 11 2 15 13 10 0 9 14 13 1 1 10 9 2
6 9 11 2 11 2 11
12 13 10 0 9 1 11 2 3 15 13 3 2
8 13 12 9 3 13 3 3 2
9 13 12 0 9 3 13 10 9 2
12 15 4 13 1 10 9 13 2 11 11 2 2
5 0 9 7 0 2
4 0 9 3 2
2 11 14
18 14 3 10 9 7 15 15 13 3 15 13 3 7 10 9 15 13 2
10 10 9 4 13 3 0 1 10 9 2
17 15 4 13 9 3 1 10 0 9 7 13 3 3 0 10 9 2
9 7 10 0 9 13 14 13 9 2
17 13 1 8 9 1 9 15 4 13 1 10 9 7 13 1 9 2
23 15 3 4 13 14 13 2 0 9 2 9 7 13 9 13 9 3 1 10 0 0 9 2
22 14 16 15 13 9 0 1 15 16 15 3 13 0 9 10 13 7 13 1 10 9 2
8 13 15 10 9 1 9 9 2
57 15 13 10 0 9 9 13 3 1 15 9 14 9 2 7 16 15 13 0 14 13 15 3 3 2 3 9 13 1 10 9 1 9 2 2 7 16 15 4 13 0 2 15 13 15 4 13 1 9 9 2 16 15 9 13 15 2
22 15 13 16 10 9 4 3 13 2 7 15 4 13 16 15 13 10 9 1 9 9 2
17 15 3 13 14 13 10 0 9 13 10 0 0 9 10 9 5 2
8 16 13 10 0 9 2 6 2
16 10 0 9 13 9 7 15 3 13 14 10 9 14 13 15 2
19 13 10 9 1 10 9 9 7 13 15 13 9 14 13 10 9 1 9 2
29 6 2 15 4 13 10 9 1 10 9 9 13 1 9 7 9 16 15 13 10 0 3 0 9 9 1 0 9 2
12 10 0 9 4 13 11 7 11 1 15 9 2
6 11 9 2 9 9 2
2 6 2
25 3 15 13 10 3 0 9 1 9 15 13 14 13 11 9 1 7 12 1 15 13 15 0 9 2
7 15 13 9 7 0 9 2
17 15 13 3 0 3 15 13 15 4 13 14 13 15 10 9 9 2
15 15 4 14 13 0 9 3 15 13 11 9 2 9 9 2
8 15 4 13 10 9 13 3 2
10 10 9 13 2 15 13 10 0 9 2
11 8 2 15 13 15 1 16 13 10 9 9
12 7 1 12 9 3 15 13 15 13 3 0 2
9 2 6 3 14 1 10 0 9 2
8 13 15 10 9 14 13 15 2
14 8 2 10 9 1 9 4 15 13 14 13 10 9 2
20 8 2 13 15 10 0 9 14 13 15 10 9 16 15 13 15 1 10 9 2
28 9 9 9 13 1 9 2 10 9 13 10 0 9 9 2 3 15 4 13 10 9 9 3 2 13 1 0 9
12 13 0 9 1 15 1 10 9 1 1 9 2
3 0 9 2
15 15 13 10 12 5 12 9 0 9 7 15 13 1 11 2
22 15 4 13 1 15 9 14 1 11 11 7 15 4 13 13 1 10 9 1 11 11 2
12 15 9 13 10 0 9 7 15 13 15 3 2
8 15 13 3 0 1 10 9 2
5 4 15 13 15 2
13 16 3 3 3 4 15 13 1 10 9 9 3 2
1 9
7 15 13 15 9 11 13 2
4 15 13 15 2
22 7 15 13 10 0 2 0 9 2 3 12 15 13 2 9 4 13 12 0 9 2 2
21 15 4 13 1 10 9 2 9 1 0 9 7 15 13 14 13 10 9 9 3 2
20 16 15 9 4 14 13 14 13 10 9 9 2 15 4 13 10 9 13 15 2
2 6 2
28 13 15 9 3 3 4 13 15 1 7 15 4 13 0 2 0 2 0 2 7 4 14 13 14 13 1 15 2
11 10 9 4 15 13 16 13 1 15 9 2
11 10 9 4 15 13 14 13 1 15 9 2
5 4 11 13 0 2
6 16 14 2 15 13 2
16 15 0 9 4 3 13 10 11 9 2 15 4 14 13 9 2
24 16 15 4 13 10 9 2 11 4 13 0 16 10 9 10 15 13 15 9 1 13 3 13 2
15 15 4 13 9 1 10 3 0 9 2 7 15 13 11 2
14 3 13 10 9 0 1 10 9 16 0 9 14 13 2
8 15 13 1 10 9 1 11 2
19 3 10 9 9 2 15 13 9 2 10 13 3 0 1 9 4 13 3 2
10 11 7 10 9 1 0 9 13 0 2
30 15 13 11 11 2 15 13 0 2 3 4 14 13 9 9 7 9 9 3 13 15 2 15 13 15 2 13 2 9 2
20 8 16 9 15 13 13 10 0 7 13 9 15 4 13 7 3 13 10 9 2
19 9 2 13 15 0 14 13 14 13 10 9 16 15 13 3 3 0 2 2
10 15 4 14 13 14 13 10 9 6 5
13 15 4 14 13 14 13 15 2 15 13 3 3 2
11 15 4 14 13 15 14 13 9 7 9 6
2 6 11
6 6 6 6 6 6 6
6 15 13 3 14 15 2
1 6
7 15 13 14 10 1 15 6
5 15 13 15 11 2
5 15 4 14 13 2
5 3 4 15 13 2
7 15 13 14 15 13 15 2
23 15 4 3 13 3 15 13 1 9 7 3 15 13 14 3 0 15 3 13 1 0 9 5
4 15 13 15 6
2 15 2
9 6 7 15 4 14 13 15 9 5
30 9 2 15 13 3 15 13 15 13 14 11 7 4 14 13 15 13 15 2 15 13 15 10 13 15 15 4 13 1 2
7 9 2 3 15 13 0 2
7 9 2 3 4 15 13 2
10 6 15 3 13 14 3 3 0 1 15
8 7 15 9 13 0 1 15 2
25 4 15 13 10 9 1 11 7 3 13 15 1 11 11 7 13 10 0 13 2 13 9 1 15 2
39 15 13 14 13 10 9 1 15 9 1 11 2 4 15 13 0 14 3 13 10 9 15 13 1 15 9 7 13 15 3 1 10 9 7 15 13 1 0 2
2 9 9
15 6 3 10 9 13 9 0 10 13 15 4 13 15 3 2
16 7 10 9 13 1 10 11 7 10 11 13 11 12 1 9 2
15 15 4 14 13 10 9 16 0 9 4 13 14 13 0 2
32 7 9 1 9 16 15 4 13 15 9 10 9 13 0 15 13 10 0 9 7 3 9 1 11 2 11 2 11 2 11 8 2
5 3 10 9 9 2
6 6 3 3 15 4 2
15 15 13 0 9 10 13 9 13 1 10 11 10 13 15 3
25 16 1 9 15 13 9 9 3 6 9 9 13 10 0 8 3 15 13 5 13 15 13 15 9 2
11 3 4 15 13 9 1 15 0 9 9 2
21 15 13 0 16 15 0 9 4 13 15 2 7 15 4 14 13 15 14 13 15 2
17 15 4 13 3 12 1 15 7 15 3 13 1 10 12 9 9 2
34 15 4 13 10 10 9 1 10 9 9 9 7 13 10 1 10 0 9 2 3 10 9 2 1 10 0 9 14 13 10 9 4 13 2
12 13 10 9 12 5 12 9 10 9 1 9 2
15 13 9 1 9 9 1 9 2 9 2 8 1 10 9 2
24 15 13 0 16 10 9 14 4 13 1 9 7 16 10 1 15 13 15 9 4 13 3 0 2
17 13 1 10 9 13 1 2 9 9 2 7 2 0 9 9 2 2
8 10 9 1 0 9 15 13 2
38 10 9 4 14 13 15 9 1 10 0 9 9 9 1 9 4 14 13 15 9 16 15 13 7 15 4 13 10 9 9 1 10 0 9 7 13 15 9
9 15 13 10 9 1 11 14 11 2
3 6 13 2
4 16 15 4 2
3 12 9 2
14 6 2 15 13 16 11 14 13 9 13 1 3 3 2
12 7 15 13 14 13 10 9 13 10 9 9 2
8 7 10 9 13 0 9 9 2
8 16 0 9 13 15 12 9 2
13 3 0 1 10 9 7 9 15 13 3 13 12 2
27 3 4 9 6 13 10 1 10 9 10 13 10 9 9 2 7 10 9 1 9 9 15 13 1 10 9 2
2 6 2
23 10 9 15 3 13 15 2 7 13 15 1 10 3 1 15 9 4 4 13 1 12 9 2
3 6 13 2
4 13 15 2 5
12 13 3 7 10 9 13 10 9 15 4 13 5
1 8
3 12 9 2
5 2 12 9 11 11
3 2 0 9
3 12 9 2
3 2 11 11
5 2 12 9 11 11
4 2 0 9 9
3 2 11 9
6 2 11 2 1 2 11
3 2 9 9
5 2 11 11 2 9
5 2 9 7 9 9
4 0 9 9 2
27 9 1 10 0 9 7 4 10 9 2 9 2 10 15 13 15 2 1 15 9 7 9 9 3 13 0 2
17 7 4 15 3 13 14 13 16 15 13 16 9 4 13 14 13 15
4 11 13 0 2
31 15 4 13 9 1 1 12 9 7 15 13 15 10 10 9 2 15 4 14 13 0 1 9 0 7 15 13 14 9 0 2
27 15 13 15 14 13 0 2 4 15 13 14 13 10 9 2 16 15 13 10 9 2 15 13 15 4 14 2
23 15 13 3 14 13 0 7 0 7 15 4 13 15 10 9 16 15 4 13 15 3 3 5
6 15 13 14 3 0 2
6 9 13 3 3 0 2
29 15 4 13 15 13 14 13 1 9 2 16 3 15 4 13 1 15 9 9 14 13 15 13 0 1 9 7 9 2
14 15 4 14 13 16 15 13 0 0 14 13 1 15 2
8 15 3 13 3 1 10 9 2
8 15 4 10 9 9 13 1 2
20 13 1 10 9 1 9 10 13 3 0 9 16 13 2 13 7 13 9 9 2
27 15 13 10 9 9 1 10 0 9 9 7 10 9 13 15 14 13 15 0 9 1 15 9 1 15 9 2
32 15 13 14 3 0 1 10 9 9 16 15 3 13 12 9 2 16 10 0 9 13 12 7 12 9 1 10 14 13 10 9 2
23 10 0 10 9 2 10 0 10 9 7 10 0 10 9 10 0 10 9 1 10 9 3 2
20 0 1 0 9 15 4 14 13 0 0 9 7 10 9 14 13 12 9 3 2
7 1 9 10 13 0 9 2
11 15 3 13 15 10 0 9 7 9 9 2
14 15 13 0 1 9 10 13 10 0 0 1 10 9 2
13 15 13 15 13 0 2 7 15 13 1 10 9 2
26 10 9 13 14 13 0 9 3 3 2 16 15 4 14 13 14 13 3 3 1 10 9 1 15 2 5
10 3 3 14 13 1 1 10 11 11 2
16 15 13 14 13 1 1 10 11 9 2 3 12 5 12 5 5
29 15 13 3 12 7 15 13 3 12 9 10 9 1 9 2 3 10 9 0 2 15 13 14 13 12 9 10 9 5
22 15 9 13 1 11 7 15 13 3 2 12 7 0 16 15 13 15 9 14 3 2 6
5 0 0 9 5 12
3 11 5 12
3 7 6 2
27 4 9 13 3 3 15 4 13 15 14 13 1 1 10 11 9 7 10 0 9 14 13 2 13 9 2 5
2 6 2
14 13 0 15 13 10 9 2 0 1 15 3 13 9 5
18 15 13 10 11 9 9 2 1 10 0 0 9 2 3 10 9 9 2
17 15 13 3 5 12 0 2 10 13 15 13 10 0 9 7 3 2
8 3 13 10 9 9 9 2 8
6 4 14 13 1 15 2
22 16 15 4 14 3 13 0 9 2 15 4 3 13 1 3 14 13 10 9 9 3 2
6 6 9 15 13 15 13
14 4 10 9 9 9 13 1 16 15 14 13 1 9 2
19 15 13 1 10 9 9 2 15 13 14 13 15 10 9 15 4 13 9 2
89 13 10 9 1 9 14 13 16 9 13 3 9 2 9 1 11 7 6 9 1 11 4 13 3 3 16 15 4 14 13 1 9 2 1 9 2 16 15 4 13 1 9 2 2 10 9 15 4 9 2 2 14 13 9 2 10 13 3 0 2 15 13 10 0 9 0 1 9 14 13 0 0 9 7 15 13 14 13 10 9 3 15 4 4 13 9 2 9 2
6 9 1 11 13 12 9
15 2 15 3 13 2 13 0 1 0 3 13 1 7 0 7
15 2 15 13 1 2 13 10 9 10 4 13 1 10 0 9
47 1 9 2 10 0 9 9 10 13 14 4 13 1 9 9 9 4 13 0 2 15 13 0 13 10 9 1 1 10 9 2 16 10 0 9 9 13 1 9 9 4 13 0 7 0 0 8
11 0 9 13 3 0 9 1 9 1 9 2
77 15 4 13 10 0 9 9 7 15 4 3 13 1 15 11 7 15 13 16 15 13 14 13 1 10 9 1 9 16 15 4 13 15 9 7 15 13 15 6 16 15 13 15 13 0 1 9 7 15 9 13 3 0 9 1 15 7 15 13 15 13 9 10 4 14 13 9 3 3 15 4 13 10 9 1 15 2
46 15 13 3 0 2 15 4 14 3 13 14 13 10 2 10 15 13 14 13 2 13 14 13 10 9 1 10 9 2 7 3 13 10 9 1 15 9 2 10 9 10 4 13 10 9 2
3 15 4 13
6 11 11 11 11 11 11
9 15 9 2 5 12 1 12 11 2
5 13 3 13 3 2
15 15 13 10 0 9 15 13 15 9 7 4 14 13 15 2
17 15 13 3 3 0 9 2 16 15 13 7 13 7 13 2 3 2
5 9 13 3 0 2
17 10 0 9 1 10 9 13 0 1 10 0 9 1 10 0 9 2
5 9 1 9 9 2
18 3 4 15 13 15 9 9 1 10 9 15 13 10 9 3 1 9 2
14 15 9 9 13 11 2 7 15 13 14 13 1 11 2
10 4 15 9 13 11 3 13 1 11 2
15 16 6 2 15 4 14 13 14 13 15 16 15 13 3 2
15 16 6 2 15 4 13 14 13 1 12 1 10 9 9 2
16 1 11 3 13 10 9 14 9 9 3 15 13 11 3 3 2
11 15 4 14 13 1 10 9 15 13 3 2
21 15 4 13 15 7 15 13 3 1 10 9 9 1 11 3 13 10 0 0 9 2
25 3 16 15 4 14 13 10 9 14 9 15 4 13 0 1 10 0 9 9 1 10 0 9 9 2
12 15 13 3 15 4 13 7 13 0 9 9 2
34 6 16 15 13 9 9 13 1 0 1 12 7 12 9 1 10 0 9 9 2 3 10 9 4 13 15 9 7 13 10 9 1 9 2
6 3 3 13 1 9 9
5 13 10 0 9 2
10 15 4 13 1 1 10 10 9 9 2
3 11 9 2
135 15 9 13 11 11 11 7 15 13 12 9 0 7 15 13 1 0 1 11 9 1 10 9 7 15 13 9 7 15 13 0 16 13 7 15 13 9 1 15 0 9 10 13 11 14 11 7 15 13 10 11 7 15 4 13 14 13 10 0 9 10 9 4 13 14 13 7 15 13 0 14 13 3 15 13 15 7 15 13 1 9 1 10 9 7 15 13 10 9 14 9 10 9 1 12 7 15 13 15 9 13 15 16 15 13 3 3 7 15 4 14 13 16 3 0 15 9 13 7 15 4 4 13 1 10 9 3 16 15 4 13 7 15 13 9
9 6 2 13 1 15 9 7 9 2
6 15 13 10 0 9 2
23 10 9 4 13 14 13 15 16 15 4 14 3 13 2 3 16 15 13 10 0 9 9 2
9 9 9 7 9 13 14 13 0 2
17 10 9 4 13 14 13 15 3 16 15 13 0 1 9 7 9 2
12 6 2 15 4 13 10 9 1 10 0 9 2
1 6
11 0 9 9 2 4 15 13 1 0 9 2
23 15 13 14 13 10 9 9 14 13 1 11 2 15 13 12 10 13 0 1 11 1 12 2
88 9 13 2 1 10 9 2 10 9 9 13 3 16 15 4 2 3 15 13 9 10 9 2 9 4 13 1 15 3 12 9 16 9 13 3 15 4 14 13 2 2 3 15 3 3 13 14 13 1 10 9 2 16 15 3 4 13 15 3 1 11 1 12 2 2 15 13 10 9 10 13 15 1 11 12 2 4 15 13 10 0 9 10 4 13 1 15 2
7 7 4 15 13 14 13 2
45 2 1 10 9 15 2 15 4 14 13 9 16 10 9 15 4 13 14 13 2 7 9 13 2 10 9 3 1 11 13 14 3 0 7 4 3 13 10 9 2 2 10 9 6 2
23 9 7 9 9 4 13 1 9 7 11 11 2 7 10 9 13 9 4 4 13 1 15 2
18 3 0 9 13 14 13 1 10 11 9 7 13 2 13 15 2 2 8
12 3 4 15 13 10 0 9 13 1 10 9 2
28 15 4 13 10 0 9 9 7 15 13 9 1 11 16 15 13 7 16 15 9 13 3 15 9 4 13 1 2
24 4 15 13 13 10 9 9 7 10 0 13 3 9 16 15 4 14 13 15 4 13 15 10 9
38 15 4 3 13 10 0 9 7 15 4 13 10 0 9 1 15 9 9 15 13 10 9 9 1 15 3 15 13 1 11 11 7 3 15 4 14 3 2
40 6 15 4 13 12 0 9 1 9 7 12 13 0 9 15 13 1 10 9 7 13 3 1 10 9 7 13 0 14 13 10 9 3 6 10 0 9 4 13 0
1 6
15 15 13 10 9 15 13 10 13 3 3 0 14 13 1 2
1 8
18 15 13 10 9 2 15 13 0 14 13 2 3 0 7 0 1 10 9
15 9 13 0 3 2 7 13 10 9 9 1 10 0 9 2
21 9 9 13 14 0 1 9 3 2 16 10 9 13 0 1 10 10 9 1 15 2
7 9 7 13 9 1 15 9
1 11
10 9 14 9 2 1 10 0 7 0 2
6 15 13 12 9 0 2
9 15 4 14 13 3 1 15 9 2
13 15 13 10 0 9 7 13 14 13 10 0 9 2
6 15 13 3 0 3 2
11 15 4 14 13 10 0 9 16 13 15 2
10 4 15 13 0 16 15 14 13 9 2
5 13 1 0 9 2
5 15 13 1 11 2
6 15 13 14 13 13 2
24 15 9 4 14 13 15 2 15 3 13 15 16 15 4 13 15 1 1 9 3 15 13 12 2
12 15 4 14 3 13 14 13 1 15 3 3 2
12 7 3 3 15 13 10 3 0 9 14 13 2
5 6 9 1 9 2
9 15 13 10 0 9 16 13 15 2
7 9 1 9 4 13 0 2
15 9 13 0 1 9 7 15 4 3 13 9 1 9 9 2
16 15 13 14 13 3 3 5 15 4 14 13 10 13 9 3 2
12 13 10 9 9 7 9 9 7 0 0 9 2
4 9 13 0 2
8 0 2 0 2 7 3 0 2
4 13 10 9 2
12 15 4 3 13 1 0 9 3 15 13 0 2
12 4 13 10 9 9 16 13 1 1 15 0 2
7 0 9 14 9 2 11 2
11 15 3 13 11 7 11 13 10 0 9 2
16 10 0 11 9 11 11 13 0 9 7 13 15 15 0 9 2
12 6 2 15 4 14 13 10 13 9 1 15 2
15 7 15 0 9 2 11 13 10 0 0 9 9 2 9 2
19 3 2 11 13 10 9 1 0 9 1 0 9 1 11 2 3 1 11 2
7 11 4 13 1 10 0 2
24 1 11 2 3 10 9 4 13 2 15 4 4 13 2 0 9 2 13 1 15 1 15 9 2
22 15 13 0 1 10 9 1 9 2 1 9 2 10 9 13 9 7 14 1 13 9 2
2 8 2
37 0 9 1 10 9 13 2 2 11 11 11 2 5 0 9 1 10 9 2 9 3 13 2 11 2 2 2 1 9 2 2 11 11 11 11 2 2
30 7 16 10 9 4 13 1 0 3 15 4 13 1 0 9 7 3 13 2 9 9 2 1 9 14 13 1 15 9 2
9 15 13 3 0 16 11 13 0 2
7 15 13 10 0 13 0 2
11 15 13 14 0 3 15 0 9 13 1 2
13 15 13 10 9 2 9 1 15 9 7 9 9 2
42 15 13 12 9 13 1 10 0 9 7 10 9 10 4 13 1 12 1 10 9 7 10 9 2 15 4 3 13 10 9 3 3 3 15 4 13 10 0 9 1 12 2
17 3 4 15 3 13 15 3 16 15 4 14 13 10 0 9 13 2
17 4 15 13 0 16 15 13 10 9 7 13 10 0 9 3 3 2
38 13 10 9 1 7 13 16 10 9 13 3 3 2 4 13 9 1 10 9 2 16 10 9 13 3 3 16 10 9 3 3 10 9 13 14 10 9 2
38 16 10 0 13 3 16 10 9 3 2 3 13 0 16 9 1 10 9 4 13 2 15 4 13 10 9 9 2 9 9 2 9 9 2 9 2 8 2
30 16 9 4 13 2 7 15 3 13 10 9 2 13 13 10 9 2 16 15 13 3 3 2 13 13 1 1 10 9 2
33 15 13 7 10 9 1 10 9 1 10 9 9 2 7 10 0 9 9 10 13 10 10 9 2 1 10 9 10 10 9 9 13 2
15 0 9 14 13 12 9 9 1 11 12 16 3 7 3 2
42 15 4 13 15 11 12 14 13 12 9 9 7 15 13 16 15 4 14 13 10 9 3 2 15 13 14 13 10 9 1 10 9 2 1 10 9 2 14 13 10 9 2
17 15 4 0 11 9 13 3 15 13 14 13 9 3 15 4 13 2
10 4 15 3 13 10 9 9 1 15 2
6 15 13 10 0 9 2
10 6 10 9 9 4 13 10 0 9 2
16 15 13 9 0 7 13 0 15 13 10 9 3 13 10 9 2
14 15 4 13 3 7 13 0 15 9 4 14 13 8 2
21 15 13 3 0 14 13 10 9 10 13 3 0 7 0 1 15 3 15 13 3 2
15 10 9 9 13 3 7 4 14 13 0 9 1 15 9 2
17 10 9 9 9 13 10 0 9 16 13 15 13 9 1 10 9 2
9 0 0 9 13 15 2 1 11 2
1 8
21 15 13 10 0 3 14 9 1 0 12 9 9 1 10 12 9 1 15 11 9 2
1 8
14 1 0 9 1 0 2 9 9 2 13 13 15 9 2
1 8
8 4 10 9 1 11 4 13 2
25 15 13 10 9 1 0 9 13 10 9 1 0 9 7 15 9 4 13 15 13 10 9 1 11 2
21 15 9 13 15 13 9 7 3 4 14 4 13 15 4 13 15 13 15 15 13 0
11 6 2 15 13 3 10 9 1 10 0 9
16 10 9 1 11 4 1 12 9 1 10 9 13 9 1 10 9
47 10 9 9 1 10 9 9 1 11 2 11 11 9 4 13 16 15 13 10 9 9 1 10 13 9 9 1 0 9 1 10 9 7 10 0 9 13 16 15 13 2 9 2 1 10 9 2
40 15 4 14 13 15 13 1 1 0 9 13 10 3 0 9 2 9 13 1 9 7 9 7 10 3 0 9 10 13 1 1 9 9 1 9 1 9 1 9 2
6 6 2 15 13 9 2
16 15 9 13 15 13 1 1 15 9 7 13 14 13 15 9 2
42 13 15 13 15 2 13 3 15 13 1 9 7 4 13 10 0 9 1 15 9 2 13 3 3 13 15 9 15 2 15 13 10 0 9 16 15 13 14 13 15 9 2
5 0 9 1 11 2
23 15 4 13 15 9 3 1 15 0 9 9 9 7 15 10 13 16 15 13 10 0 9 2
16 15 4 13 1 10 9 1 11 11 11 3 15 13 9 0 2
12 15 4 13 10 9 13 3 1 9 1 9 2
28 15 4 3 13 1 10 9 9 1 10 0 9 1 10 9 1 10 9 7 15 4 13 15 1 1 12 9 2
20 15 4 3 13 1 10 1 10 9 3 10 9 7 7 9 4 13 3 0 2
17 15 4 13 1 1 11 7 11 2 11 14 2 7 11 11 14 2
7 9 1 9 1 10 9 2
29 9 2 15 13 0 1 10 11 11 2 11 11 2 10 11 2 10 11 11 2 11 14 2 11 11 14 2 8 2
23 15 4 13 10 9 7 13 10 12 10 15 4 13 14 13 3 15 9 7 15 0 9 2
10 6 3 9 1 10 12 15 13 3 2
3 0 9 2
11 15 13 3 0 1 11 14 7 11 11 2
19 15 4 3 13 1 10 9 15 4 13 7 4 15 13 1 9 15 13 2
7 15 13 15 13 15 9 2
8 6 2 13 10 0 0 9 2
12 9 2 4 10 9 13 0 13 1 10 9 2
7 1 15 9 1 10 9 2
11 7 4 10 9 1 10 9 13 10 9 2
2 9 11
33 16 9 13 0 2 7 15 4 13 15 1 3 14 4 13 3 1 0 9 2 3 15 4 13 3 15 4 13 14 13 15 3 2
8 15 13 10 9 14 13 3 2
36 9 13 0 9 1 15 9 14 13 15 9 2 7 15 13 14 4 13 3 2 7 15 9 4 13 1 9 1 10 9 1 9 1 15 9 2
39 3 15 13 10 9 9 7 13 1 9 2 15 9 4 13 9 2 10 9 4 13 0 1 15 2 7 4 14 13 0 14 13 10 9 3 16 15 4 2
21 15 4 3 13 14 13 0 16 9 13 1 10 9 7 9 2 9 15 4 13 2
14 15 3 4 14 13 15 13 3 0 1 15 3 3 2
37 3 2 15 13 14 10 0 9 2 7 15 4 13 15 0 7 13 15 1 16 15 13 10 9 14 13 15 10 0 9 15 4 13 1 1 15 2
12 15 4 13 10 9 16 10 9 4 3 13 2
8 15 4 3 13 15 3 3 2
12 15 13 10 3 0 9 14 13 1 11 11 2
16 15 4 13 15 9 1 11 7 11 11 13 12 1 10 9 2
13 10 9 7 9 4 13 3 0 14 13 1 11 2
5 13 1 11 9 2
19 15 13 3 0 9 1 3 2 7 15 13 0 16 15 4 13 15 2 5
23 16 15 4 13 1 11 2 3 15 4 3 13 10 0 9 13 2 2 10 11 11 2 2
24 15 13 10 3 0 9 1 3 2 7 3 0 9 2 9 13 14 13 9 7 9 1 3 2
6 15 13 3 0 9 2
24 3 2 4 14 13 14 13 1 11 14 0 9 9 2 2 11 11 2 11 2 7 11 11 2
5 9 13 15 2 5
4 11 11 2 8
8 2 15 13 3 7 3 2 2
4 11 11 2 8
18 2 15 13 3 3 7 10 9 13 3 10 9 1 10 0 11 2 2
4 11 11 2 8
7 2 10 0 9 9 2 2
4 11 9 2 8
5 13 15 13 2 5
5 13 9 1 11 2
7 10 9 13 11 2 11 9
11 15 13 3 0 3 2 15 4 13 15 9
6 15 13 3 1 9 3
13 15 13 10 0 0 0 9 2 9 15 13 2 2
6 15 4 15 13 15 2
24 15 13 10 0 0 9 1 15 9 2 15 9 13 0 2 3 15 4 3 13 9 1 15 2
27 15 13 0 0 2 10 9 7 9 7 9 2 15 4 14 13 10 9 1 9 15 13 2 3 10 9 2
6 15 4 15 13 15 2
6 13 0 9 9 0 2
38 2 16 3 15 9 13 3 0 2 15 13 10 9 4 13 0 16 15 4 14 13 10 0 9 2 13 15 10 0 9 15 4 13 1 10 9 9 2
8 2 11 2 11 2 2 9 2
21 9 13 10 9 1 9 2 15 13 9 9 2 15 4 14 13 9 2 7 9 2
13 13 0 16 15 13 10 0 9 1 9 1 15 2
7 16 15 4 13 10 9 2
13 15 13 10 0 6 9 9 1 11 14 2 9 2
11 15 13 11 14 11 7 11 15 13 2 2
9 6 15 13 15 1 15 9 3 2
5 6 10 0 9 2
6 7 13 0 9 9 2
3 15 4 13
27 16 15 13 10 9 9 3 13 10 9 2 9 9 7 3 13 9 9 4 13 2 7 4 14 13 9 2
12 3 4 15 13 1 11 11 11 1 11 11 2
4 15 13 12 9
8 13 10 11 7 10 11 11 9
14 4 9 13 15 16 10 11 13 3 1 11 1 11 2
9 16 14 10 9 4 15 13 1 2
1 6
6 1 10 11 2 11 2
15 1 10 9 2 13 10 9 10 13 2 11 1 9 2 2
6 13 10 9 1 11 2
13 15 4 13 15 1 10 11 9 9 13 1 9 2
15 13 1 15 1 10 2 11 2 11 11 2 11 2 9 2
15 13 3 1 10 11 12 9 13 1 2 11 11 11 2 2
10 13 3 1 10 2 11 11 2 9 2
6 1 10 11 11 9 2
15 16 15 13 2 10 9 13 15 1 1 10 11 1 11 2
15 15 4 3 13 14 13 10 9 7 10 11 3 1 11 2
16 1 10 9 2 13 1 9 12 13 1 2 11 11 11 2 2
7 13 10 9 1 10 9 2
12 13 1 10 9 1 10 2 11 11 2 9 2
11 1 10 11 2 13 1 10 11 1 11 2
15 13 10 12 9 1 2 11 2 1 10 2 11 2 9 2
22 13 3 1 10 12 9 1 2 11 11 2 7 13 15 1 10 2 11 11 2 9 2
10 15 13 0 0 7 0 9 14 9 2
13 15 13 3 0 9 1 0 0 0 7 0 9 2
13 15 13 11 7 15 4 14 13 15 2 13 0 2
10 3 13 12 1 15 9 1 0 7 0
1 8
9 10 9 10 15 13 6 13 5 9
8 15 4 3 13 15 1 11 2
22 15 4 13 15 10 9 0 9 2 3 3 1 9 16 3 15 0 7 0 9 13 2
9 13 15 9 16 15 13 3 1 9
11 13 10 0 9 7 13 10 9 1 9 2
17 13 10 9 9 1 2 9 2 15 4 13 15 9 0 7 0 2
12 13 9 5 9 7 13 10 9 14 9 9 2
14 15 4 13 10 9 7 9 1 0 9 1 10 9 2
17 1 0 9 1 10 9 1 0 9 13 1 10 11 9 9 2 8
16 1 0 9 16 13 9 1 11 13 1 10 11 9 9 2 8
4 13 15 13 2
7 11 13 0 7 3 0 2
17 7 0 13 3 11 11 7 16 15 13 1 10 11 15 13 11 5
21 13 15 15 13 1 2 0 7 0 2 2 0 9 4 13 10 0 0 7 0 2
9 13 9 1 11 10 13 0 9 2
6 0 0 9 1 11 2
32 15 13 14 13 1 11 14 13 15 9 9 1 11 11 7 13 1 10 0 9 3 3 0 1 15 9 1 10 9 14 9 2
16 3 10 9 4 13 10 9 13 10 0 9 14 13 10 9 2
20 0 9 13 1 1 10 0 9 7 4 14 13 10 9 15 4 13 1 2 2
13 4 15 3 13 14 13 15 9 1 10 9 9 2
6 15 13 15 4 14 2
21 15 13 14 13 1 12 1 10 0 9 10 13 10 9 1 11 11 7 11 11 2
18 4 15 13 10 0 9 1 15 0 9 9 7 3 10 0 9 3 2
8 3 10 2 0 2 13 0 2
21 3 15 13 0 9 15 4 3 13 9 2 0 9 7 9 10 13 0 9 3 2
15 16 15 13 1 15 4 13 1 0 9 16 15 13 3 2
18 11 11 13 10 0 9 7 10 9 4 13 15 9 1 9 1 9 2
18 3 13 10 0 9 4 13 0 1 10 9 10 13 0 7 3 0 2
1 8
13 10 0 2 0 9 2 0 9 13 1 11 11 2
5 15 13 0 9 2
9 13 10 9 1 10 9 1 9 2
14 15 9 9 4 14 13 9 3 10 9 1 10 9 2
20 3 15 13 10 9 1 9 1 9 15 13 1 10 9 7 13 10 9 13 2
6 15 4 13 15 1 2
2 3 2
20 16 15 13 10 9 1 2 9 2 15 13 1 13 9 9 15 4 13 15 2
15 15 4 13 10 9 1 9 15 13 14 13 10 13 9 2
12 3 15 13 10 9 15 13 0 14 13 3 2
15 15 4 13 9 1 12 9 7 15 3 13 15 0 9 2
12 15 4 13 3 3 7 13 10 0 9 3 2
12 15 13 0 0 9 7 15 13 3 3 0 2
24 13 9 13 3 0 1 1 10 0 9 7 15 4 13 1 10 0 9 9 3 1 9 9 2
11 15 13 10 9 1 0 9 0 9 9 2
6 13 10 9 1 9 2
6 15 9 4 13 3 2
7 15 4 3 13 0 9 2
11 15 4 13 0 13 15 1 10 9 14 13
11 16 15 3 13 15 2 6 1 10 9 2
40 15 0 9 7 0 9 13 15 2 15 3 13 10 9 7 13 1 10 0 9 1 15 1 9 9 2 13 2 1 10 0 9 2 10 9 9 1 10 0 2
14 3 16 15 13 15 1 10 9 15 4 14 13 15 2
9 15 13 15 0 9 1 9 9 2
10 15 0 9 13 13 8 3 7 13 2
22 15 13 3 15 3 13 1 3 0 10 9 15 9 3 13 2 7 3 0 15 13 2
20 16 15 13 10 11 2 9 9 1 10 9 9 2 15 3 4 14 13 15 2
8 15 4 13 3 0 7 0 2
26 15 4 14 13 3 0 15 9 13 2 7 3 3 15 4 13 2 7 3 3 15 13 10 13 9 2
16 15 13 13 3 3 13 15 13 2 7 3 0 15 9 13 2
12 15 13 10 9 3 15 13 0 9 9 3 2
29 9 13 9 14 13 15 9 1 9 7 13 3 10 9 2 3 13 10 10 9 1 10 9 16 15 9 13 0 2
8 15 13 14 13 10 9 13 2
12 7 15 4 14 13 12 13 2 1 9 9 2
16 15 13 3 10 0 9 3 15 13 9 9 2 0 7 14 2
18 0 2 3 15 4 13 1 10 0 9 1 15 15 4 3 13 9 2
19 13 10 9 7 0 9 10 16 15 13 0 15 4 13 3 0 7 0 2
13 15 4 13 0 0 9 1 7 9 7 0 9 2
14 3 9 4 13 1 10 9 7 15 3 13 7 13 2
2 0 2
6 12 9 9 9 9 2
23 15 13 10 12 9 9 9 1 12 9 1 0 9 9 2 7 12 9 1 0 0 9 2
14 15 13 0 1 10 9 13 16 13 10 9 10 9 2
10 15 4 3 13 10 9 9 1 12 2
9 15 13 10 12 9 9 1 15 2
10 15 3 13 10 9 2 13 10 3 2
31 15 13 10 0 9 2 3 15 13 14 13 10 9 9 2 7 15 13 10 9 16 3 10 9 9 7 9 9 4 13 2
13 3 4 15 13 14 13 10 9 1 10 12 9 2
11 4 15 13 10 9 9 7 10 0 9 2
1 9
39 16 10 9 13 10 13 1 9 9 2 10 15 13 0 15 13 14 2 3 15 13 14 13 12 1 10 13 1 9 9 9 16 16 15 4 13 10 9 2
13 10 9 4 13 3 1 15 9 1 10 9 9 2
27 1 10 0 9 1 10 9 2 15 4 13 10 0 9 9 1 10 9 10 13 10 9 3 1 15 9 2
28 16 15 4 13 14 13 1 10 9 16 13 10 9 1 10 9 2 13 10 9 9 4 14 13 10 0 9 2
26 10 11 11 11 13 10 0 9 9 9 2 15 13 10 1 2 9 9 10 4 3 13 1 15 9 2
6 11 11 7 11 11 2
12 16 15 15 13 15 13 3 3 10 0 9 2
25 10 1 10 0 9 15 13 13 10 9 9 2 0 9 9 2 7 0 9 10 10 11 11 13 2
14 4 10 9 13 10 0 9 1 9 13 1 10 11 2
9 15 4 14 13 10 11 7 11 2
15 15 3 13 10 9 10 13 10 0 9 0 16 3 13 2
28 6 2 15 13 1 10 11 11 7 15 13 14 15 15 13 5 4 15 13 9 14 13 1 10 9 12 9 2
6 7 3 13 10 11 2
21 6 15 3 13 10 11 11 2 7 15 13 14 13 16 15 13 3 0 1 15 2
8 15 13 1 10 0 9 15 2
30 3 15 13 1 15 13 3 1 10 11 11 2 15 13 3 0 3 2 16 15 13 15 11 11 1 10 0 9 9 2
13 3 15 13 15 4 13 1 10 3 0 11 11 2
10 15 13 3 0 15 4 13 0 15 2
3 13 9 2
14 13 1 11 11 14 9 15 4 13 14 13 3 0 2
19 3 11 11 15 13 0 9 2 3 0 9 7 10 0 9 7 10 9 2
1 8
21 9 11 11 2 11 7 11 11 11 2 11 7 11 11 11 2 11 11 2 11 11
1 8
4 11 1 11 2
21 6 3 2 15 4 13 14 13 10 9 1 11 14 13 15 9 9 1 15 9 2
25 15 13 3 3 10 2 15 13 0 11 2 0 9 1 9 2 0 0 2 2 9 1 9 2 2
42 15 13 14 13 15 3 3 15 4 13 14 13 0 9 2 0 9 2 9 2 3 10 9 2 9 9 4 13 0 2 2 0 9 2 7 3 3 10 0 9 2 5
17 15 4 13 1 9 1 9 15 13 10 11 9 7 10 9 9 2
23 15 3 13 1 10 9 1 11 10 9 1 9 3 3 15 13 14 10 9 1 10 9 2
8 10 0 9 13 3 0 2 5
7 13 15 1 15 9 9 2
12 6 6 2 15 13 10 9 1 10 0 9 2
22 13 1 10 0 9 7 9 9 2 7 13 10 9 14 9 1 10 2 11 11 2 2
12 15 13 3 1 10 0 9 2 9 7 9 2
10 15 13 9 3 1 10 9 7 9 2
7 13 15 9 10 0 9 2
32 16 15 4 13 1 10 0 9 2 10 0 9 2 15 13 14 13 1 2 2 2 7 0 9 2 13 1 11 7 11 14 2
8 6 6 6 2 15 13 0 2
18 16 15 13 2 13 0 15 13 10 9 9 2 15 4 14 13 15 5
8 3 14 13 10 0 0 9 2
23 15 4 13 10 12 9 1 15 9 9 7 15 3 13 14 13 3 14 3 13 15 1 2
6 15 13 3 10 9 2
15 10 7 10 9 16 15 15 13 14 13 7 13 4 13 2
2 9 2
38 3 15 13 10 9 13 0 15 13 10 9 2 1 0 9 2 3 15 13 10 9 2 1 3 9 3 2 13 1 10 10 9 10 4 13 1 9 2
16 13 3 0 9 16 0 9 4 13 1 15 9 14 0 9 2
12 15 13 10 9 7 13 9 9 1 10 9 2
28 13 1 15 9 2 9 9 13 10 0 1 9 2 7 13 1 10 9 7 13 15 1 9 1 12 5 12 2
11 13 3 12 9 7 12 7 13 15 9 2
15 16 9 4 13 0 15 4 13 15 9 1 15 0 9 2
28 9 13 0 16 9 13 10 9 13 1 1 9 3 7 10 9 9 13 14 0 16 15 13 9 1 10 9 2
17 13 10 9 13 15 10 9 3 15 4 13 15 1 2 15 4 13
10 13 9 1 10 9 15 13 1 15 2
7 13 0 10 9 13 0 2
17 4 14 13 15 0 9 3 1 10 9 7 9 13 1 15 9 2
6 9 0 4 13 0 2
15 13 0 16 15 13 0 9 16 15 13 3 1 12 10 2
11 13 15 0 14 13 9 1 1 15 9 2
6 15 4 13 14 13 3
10 15 13 15 4 3 13 1 10 9 2
8 15 13 14 4 13 0 3 2
5 15 13 0 2 5
14 3 1 0 9 7 9 2 9 9 9 2 9 2 5
1 8
18 13 16 15 13 9 7 9 1 9 9 16 15 13 15 1 15 9 2
28 16 15 13 3 0 2 9 9 4 14 13 3 3 0 7 0 16 10 9 3 4 14 13 1 1 10 9 2
9 3 2 15 4 13 14 13 3 2
1 8
11 13 9 9 3 3 16 13 10 9 9 2
9 9 9 13 10 3 0 1 9 2
20 10 9 4 13 1 10 9 9 7 13 10 9 1 10 9 14 13 15 1 2
16 13 15 9 1 10 13 9 7 13 15 1 15 0 9 9 2
15 15 13 12 9 9 1 0 7 0 7 0 1 0 9 2
1 8
11 13 10 9 16 13 9 9 1 0 9 2
14 0 0 9 13 10 9 13 1 10 9 1 10 9 2
16 10 9 4 13 1 8 9 2 0 1 9 9 7 9 9 2
1 8
13 13 14 13 10 9 9 1 10 9 1 10 9 2
12 15 13 12 9 10 13 10 9 1 10 9 2
5 13 10 9 3 2
23 13 10 9 7 13 15 9 9 13 1 10 9 1 10 9 9 10 13 1 10 9 9 2
9 12 9 0 9 9 0 1 9 2
27 15 13 10 12 9 0 9 9 7 15 13 16 15 2 15 9 4 14 13 1 15 1 10 9 1 9 2
28 15 13 14 13 16 15 3 13 10 9 1 10 9 0 1 10 2 9 9 2 16 15 7 10 9 4 13 2
39 15 13 3 0 14 13 1 10 9 7 13 10 9 7 15 3 4 13 3 3 1 10 9 1 15 7 13 15 10 9 3 3 2 3 10 9 13 3 2
13 15 13 15 13 0 1 10 9 3 15 13 15 2
28 15 13 3 10 9 1 15 0 2 10 9 13 0 7 15 4 14 13 1 10 9 14 13 1 15 1 9 2
5 15 13 10 9 2
20 13 15 10 0 9 1 10 9 2 16 15 2 15 4 13 0 3 0 9 2
20 15 13 14 13 16 10 9 4 14 13 1 15 7 9 2 15 2 15 13 2
14 9 13 9 13 9 7 15 4 13 10 9 13 0 2
20 3 10 9 13 15 9 3 10 9 13 0 1 15 13 15 4 14 13 9 2
18 15 13 0 2 3 13 0 16 10 9 10 9 13 1 4 13 0 2
20 16 10 9 13 0 3 2 10 15 13 0 15 13 3 2 15 4 13 0 2
14 3 13 14 13 0 10 9 4 3 13 1 10 9 2
9 13 10 9 1 15 2 3 2 5
10 4 15 13 1 11 1 10 11 11 2
37 6 3 15 13 14 10 0 9 2 7 15 9 13 4 15 13 1 10 11 11 9 3 15 13 1 11 2 4 15 13 9 1 10 11 11 9 2
8 7 4 15 4 13 1 15 2
12 15 13 0 16 15 4 14 13 10 9 3 2
7 15 13 9 13 15 15 13
4 1 0 6 2
6 3 14 1 10 9 2
23 16 15 2 11 2 9 13 10 9 1 10 0 0 9 2 15 9 7 9 4 13 3 2
9 15 4 2 3 2 13 10 9 2
22 10 0 9 14 13 1 0 13 14 13 12 2 7 15 9 9 9 9 2 7 13 2
29 10 9 7 9 13 0 2 3 10 0 9 15 4 14 13 4 13 16 15 13 2 6 2 10 0 9 9 9 2
19 6 15 4 2 7 15 4 13 15 9 1 9 16 15 13 10 0 9 2
14 6 15 4 13 1 11 1 10 11 1 10 11 9 2
5 10 9 4 13 2
6 15 13 9 1 9 2
14 15 4 13 14 13 10 0 9 1 15 9 1 11 2
15 13 15 10 0 9 14 13 7 4 15 9 3 13 9 2
10 9 3 0 16 15 13 10 9 9 2
26 3 15 13 0 14 13 16 15 4 13 10 0 9 7 10 1 10 9 9 13 13 10 1 15 9 2
17 13 15 13 10 9 15 4 13 10 2 9 2 9 1 15 9 2
8 15 13 9 1 15 0 9 2
19 6 2 15 13 15 0 9 2 11 2 3 9 7 16 15 4 13 14 13
9 15 14 13 14 13 15 0 9 2
37 16 15 13 1 10 0 9 15 4 13 1 10 9 1 10 9 7 15 4 13 13 3 16 15 4 13 7 15 13 14 13 7 15 13 0 3 2
38 3 3 15 13 14 13 1 9 1 15 3 15 13 10 9 1 9 7 15 13 15 1 15 9 2 15 13 3 3 7 15 3 13 3 1 15 9 2
34 3 2 3 4 15 13 1 8 9 1 15 15 4 3 14 13 10 9 10 15 13 1 7 15 13 1 13 3 7 13 14 13 3 2
8 6 13 15 13 0 1 15 2
2 9 2
3 13 1 2
13 3 2 15 9 4 14 13 1 2 15 13 9 2
15 3 2 15 13 0 9 16 15 13 10 9 1 10 9 2
14 3 2 3 13 15 9 1 15 9 7 13 15 3 2
17 15 4 3 13 7 13 15 7 3 15 4 13 15 10 0 9 2
4 13 15 13 2
4 13 15 9 2
6 15 3 13 15 9 2
8 15 13 3 3 0 7 0 2
20 16 15 4 3 13 1 2 13 0 1 10 0 9 7 9 15 4 13 0 2
23 16 15 13 3 0 1 15 9 2 3 15 4 13 13 15 7 13 14 13 10 0 3 2
8 7 3 13 15 9 1 3 2
9 13 11 10 0 9 14 13 1 2
16 15 9 7 15 4 13 14 13 1 11 1 10 9 1 9 2
20 3 15 3 13 14 13 16 15 13 10 0 9 14 13 1 7 1 10 9 2
22 3 16 2 15 13 1 10 0 0 9 11 4 13 3 0 1 11 2 13 15 0 2
20 15 4 13 0 16 9 13 2 3 9 15 4 13 1 11 7 13 3 2 5
4 15 13 3 2
23 2 15 4 4 13 1 11 15 0 9 7 15 4 13 16 15 4 13 1 10 0 9 2
25 15 13 12 4 13 14 13 10 0 9 1 11 16 15 13 10 9 1 9 14 4 13 1 12 2
6 9 14 13 1 11 2
16 15 13 1 9 7 9 3 15 4 13 1 9 7 1 9 2
20 2 9 2 9 9 2 9 2 9 13 10 1 10 9 15 4 13 1 9 2
16 7 3 15 4 13 10 9 1 11 7 11 1 12 9 3 2
30 3 2 6 15 13 14 3 0 1 11 2 7 15 13 0 7 3 0 2 7 15 4 3 13 1 11 1 12 9 2
9 6 13 15 13 16 15 13 9 0
6 13 11 3 1 11 2
9 9 1 11 2 7 3 4 13 2
23 4 14 13 10 9 1 11 7 11 13 3 0 3 15 4 14 13 14 13 1 1 15 2
23 16 15 13 10 0 9 15 13 2 7 0 9 9 16 13 2 15 4 13 3 1 15 2
7 13 15 10 0 9 9 2
14 15 4 14 13 4 15 13 11 7 11 2 11 11 2
8 7 3 11 2 11 7 11 2
20 15 13 10 0 0 3 15 13 9 7 11 2 11 3 10 0 9 13 1 2
9 2 0 1 11 2 11 7 11 2
27 11 11 4 4 13 3 3 1 10 11 3 10 9 13 3 1 9 16 10 11 11 4 13 3 0 9 2
18 11 4 14 13 15 0 9 3 16 15 4 13 14 13 1 10 9 2
12 3 3 3 15 13 15 4 13 10 0 9 2
53 15 13 11 2 11 13 10 3 0 9 15 13 15 6 12 9 2 15 13 3 0 1 0 9 7 3 0 15 13 3 0 1 10 9 9 7 10 9 2 16 15 4 14 13 14 13 10 9 10 13 15 9 2
6 11 11 13 3 0 2
15 9 2 15 13 10 0 1 10 2 3 13 10 0 9 2
31 15 4 14 13 1 10 11 9 7 15 4 13 16 11 4 13 15 4 14 13 10 9 12 16 13 3 3 1 15 9 2
28 16 15 13 11 15 13 3 3 15 9 16 13 10 0 11 3 15 4 14 13 16 13 10 9 1 10 9 2
48 15 4 13 15 4 3 13 10 0 11 3 7 15 4 14 13 15 11 4 13 1 11 7 3 2 16 15 13 10 11 2 10 15 3 13 13 10 0 3 2 15 4 13 0 1 10 9 2
9 15 13 10 0 9 1 10 9 2
10 15 9 13 10 9 9 7 13 0 2
28 1 9 10 9 1 10 9 15 13 14 13 0 1 12 9 7 10 2 7 3 15 13 3 16 9 4 13 2
21 15 13 10 9 9 14 13 3 3 9 4 13 2 3 0 9 13 3 0 9 2
7 15 9 13 12 9 0 2
12 1 15 9 3 3 4 9 4 9 3 13 2
33 13 15 1 15 0 9 7 13 15 0 16 15 4 13 3 1 10 12 9 16 4 13 1 10 1 10 9 15 4 4 13 1 2
15 1 15 9 1 15 9 12 5 12 9 13 1 10 9 2
12 1 12 9 2 15 9 4 13 10 0 9 2
14 0 9 10 4 3 13 1 3 13 12 5 12 9 2
18 0 13 3 13 14 13 0 9 9 2 3 15 9 4 13 3 3 2
11 0 9 3 3 13 1 12 5 12 9 2
11 9 1 9 13 0 1 12 9 13 0 2
26 15 4 13 9 1 12 9 7 10 0 9 15 4 3 13 13 10 12 9 0 0 7 15 13 0 2
25 1 9 2 0 9 13 10 9 9 1 12 5 12 9 13 16 3 0 9 13 1 10 0 9 2
29 13 1 10 9 9 2 10 9 9 1 10 0 9 13 10 9 1 11 2 11 15 3 13 1 10 9 1 12 2
12 15 13 10 9 10 13 1 15 9 0 12 2
7 9 1 12 13 10 9 2
9 13 7 13 15 9 14 9 2 2
25 15 13 16 15 4 13 15 9 14 9 2 7 3 15 4 14 13 1 15 3 15 13 15 9 2
5 15 4 15 13 2
8 4 9 13 16 13 15 9 2
15 9 13 0 14 13 9 1 2 7 15 4 13 3 3 2
14 10 0 9 9 4 4 13 16 15 13 0 1 15 2
19 13 1 15 9 7 13 10 2 9 9 2 1 15 9 13 10 0 9 2
11 9 13 7 13 1 15 9 2 3 9 2
25 13 15 9 0 7 13 1 15 9 2 7 13 10 9 2 8 7 3 15 4 13 3 1 15 2
25 13 15 13 1 15 0 9 2 4 14 13 1 15 2 7 3 3 13 1 0 9 1 15 9 2
18 15 4 13 15 9 2 7 15 3 4 14 13 10 9 14 13 12 2
6 9 13 10 9 2 5
21 15 4 3 13 10 0 2 0 2 0 9 2 7 15 4 3 13 10 0 9 2
7 7 3 3 15 4 13 2
5 10 9 13 0 2
44 1 15 9 2 15 3 13 15 7 13 15 2 7 3 15 13 10 9 14 13 15 3 2 15 13 1 15 2 15 13 15 4 13 14 13 15 3 7 15 4 14 13 15 2
30 10 9 4 13 16 3 15 13 10 9 9 15 13 16 15 4 13 15 1 10 9 2 7 9 4 14 3 13 9 2
21 3 2 15 4 14 13 10 9 4 14 13 15 2 7 3 4 14 13 10 9 2
8 3 14 13 10 9 9 9 2
10 6 15 13 10 0 9 1 9 9 2
20 15 9 13 9 7 9 3 2 7 15 13 9 7 9 16 3 14 13 15 2
22 15 4 13 3 12 9 1 9 3 13 0 10 9 13 14 3 0 16 15 4 13 2
11 7 15 13 14 13 3 14 13 10 9 2
18 6 13 15 3 0 16 15 4 7 15 9 13 14 3 14 3 3 2
4 9 4 13 2
19 9 2 16 15 13 10 9 10 15 13 15 4 13 15 0 3 3 7 3
7 11 9 2 9 2 9 9
21 13 1 9 9 2 13 9 2 13 0 9 2 0 9 2 7 0 0 9 9 2
20 13 1 3 0 9 15 13 2 3 13 0 9 9 1 9 7 9 1 9 2
18 13 9 1 9 2 13 9 7 13 9 2 13 1 9 9 7 9 2
23 15 13 0 0 9 2 10 15 4 13 14 13 1 16 15 13 1 9 7 9 7 9 2
52 13 9 9 7 9 9 1 0 9 1 9 9 9 7 9 9 9 2 15 13 9 9 9 2 9 2 3 0 9 14 13 9 3 2 0 9 2 9 2 9 2 9 2 9 2 9 9 2 9 2 9 9
38 9 4 13 1 9 9 7 9 9 2 7 9 2 9 2 7 9 2 7 13 12 1 12 7 9 2 15 4 13 11 11 7 9 9 1 0 9 2
1 8
1 8
1 8
1 8
1 8
1 8
1 2
13 3 4 15 13 15 9 14 13 13 3 15 13 2
11 15 13 10 9 15 3 13 12 9 9 2
15 15 13 10 0 9 2 3 3 15 13 15 13 3 3 2
22 3 10 9 15 4 3 13 15 1 1 12 9 1 10 9 2 13 14 13 15 9 2
14 7 3 15 13 15 15 13 15 13 15 4 13 2 5
21 15 13 3 16 15 13 14 13 15 9 3 2 7 13 15 10 9 16 15 13 2
7 15 13 0 1 15 3 2
4 10 0 9 2
7 4 15 13 15 4 13 2
7 15 4 13 1 1 9 2
13 6 2 15 13 16 10 9 15 9 9 13 0 2
8 10 9 2 15 4 14 13 2
24 15 4 13 9 2 10 9 9 2 9 1 9 2 9 2 9 2 10 0 9 9 2 8 2
13 15 4 3 3 13 1 1 15 7 13 10 9 2
17 3 15 13 15 1 1 15 9 2 15 13 3 3 7 0 9 2
14 15 4 4 13 7 15 4 14 13 15 4 4 13 2
19 3 13 15 9 10 15 4 13 1 10 13 15 10 9 14 13 15 9 1
31 6 4 14 13 10 9 14 9 0 15 4 13 15 8 9 2 15 13 3 10 9 7 15 13 3 0 2 13 15 9 2
51 9 1 15 2 9 9 13 3 2 3 3 15 13 15 1 10 9 13 15 1 1 15 9 2 14 13 15 16 15 4 14 13 15 2 15 4 13 15 2 15 4 3 3 13 2 16 9 13 15 0 9
6 10 9 9 13 0 2
16 6 2 15 13 14 13 10 0 9 9 7 13 10 9 9 2
21 2 3 1 10 9 9 10 15 4 13 14 13 2 10 1 10 12 9 13 0 2
1 8
1 8
9 15 4 14 13 1 9 7 9 2
1 8
7 10 9 13 0 1 9 2
12 15 3 13 14 13 3 3 1 3 1 9 2
5 15 13 14 13 2
29 15 4 13 14 13 10 9 9 16 15 13 2 7 13 9 9 1 10 9 2 16 10 0 9 4 13 7 13 2
10 10 9 4 13 3 12 5 12 9 2
11 10 13 0 9 3 13 1 10 0 12 2
23 16 15 13 10 9 15 13 0 14 13 10 9 9 3 7 13 15 1 9 7 10 0 2
38 15 13 12 1 10 9 0 9 1 10 9 7 15 13 14 3 0 14 13 0 2 3 3 13 2 10 9 9 13 0 7 15 4 14 13 3 3 2
7 3 13 10 0 9 3 2
1 8
1 8
1 8
1 8
1 8
45 15 13 3 10 9 3 0 1 15 9 7 16 15 11 13 10 9 15 4 13 0 14 13 12 0 9 2 0 13 1 10 0 9 12 1 0 9 1 10 0 13 0 9 3 2
7 10 0 9 13 3 0 2
13 15 13 10 0 9 2 13 1 10 0 11 9 2
28 15 13 3 0 7 10 11 9 13 13 0 0 1 12 9 2 7 15 4 13 10 9 1 12 1 15 3 5
14 13 1 9 9 7 9 9 9 0 1 10 9 9 2
34 15 4 13 10 9 1 10 9 9 15 13 1 15 12 9 9 1 15 9 7 15 13 15 4 4 13 1 10 9 7 1 10 9 2
23 15 13 14 0 16 13 10 9 15 9 13 1 16 15 4 13 15 1 1 10 9 3 2
52 1 15 9 2 16 15 4 13 1 10 9 2 15 9 13 13 15 9 16 15 13 7 13 3 1 9 1 10 9 1 10 9 16 15 13 10 1 10 9 9 14 13 1 10 9 2 7 15 13 0 9 9
46 16 15 13 1 10 9 15 4 14 13 14 13 16 13 15 1 2 7 10 9 4 3 13 15 16 15 13 1 10 9 1 10 9 7 15 3 13 16 15 4 14 13 9 3 3 2
7 15 13 15 9 7 9 2
10 15 13 9 1 10 1 15 13 9 2
24 15 4 13 16 15 13 3 0 2 15 13 14 1 10 9 9 10 15 4 13 1 10 9 2
16 15 3 13 15 0 0 9 1 10 9 7 15 13 3 0 2
21 15 13 3 12 9 2 9 2 7 9 7 4 3 13 10 9 1 10 9 9 2
13 1 10 9 13 10 9 2 13 15 1 10 9 2
3 0 9 2
17 9 16 15 13 0 16 10 9 13 15 13 9 1 15 1 9 2
18 15 3 13 10 12 9 9 7 9 9 1 15 7 15 13 14 13 15
19 13 10 9 1 10 9 15 4 13 15 7 10 10 0 9 15 4 13 9
10 15 13 0 9 14 13 9 1 2 2
17 15 9 13 11 5 7 15 13 14 13 9 2 9 1 15 9 2
35 15 4 13 14 13 10 9 9 10 9 7 15 9 4 13 13 15 0 9 3 9 13 15 7 10 0 9 15 13 13 11 14 7 11 2
21 6 7 3 15 13 1 11 11 13 1 9 1 6 10 11 9 7 11 8 6 5
12 15 4 3 13 2 10 11 11 2 1 11 2
12 15 4 3 13 1 10 0 9 1 0 9 2
8 4 14 13 1 10 9 3 2
5 3 13 7 13 2
7 15 13 0 0 9 3 2
16 10 11 11 7 11 4 3 13 3 12 9 1 10 11 11 2
15 15 13 3 9 1 9 1 10 9 7 1 15 0 9 2
20 16 15 4 3 13 1 9 2 3 13 1 15 9 1 15 9 2 9 9 2
20 9 1 9 1 10 9 2 1 10 9 6 13 1 10 0 9 1 10 9 2
13 9 1 10 11 2 13 10 11 9 1 10 11 2
11 13 12 9 3 7 13 10 9 1 11 2
10 13 12 9 1 11 7 13 10 9 2
10 15 13 1 10 9 1 11 7 11 2
5 10 11 11 7 11
3 12 11 11
4 11 2 11 12
2 12 9
2 13 15
4 9 1 9 2
3 11 1 11
5 12 9 5 12 9
3 11 7 11
5 12 9 5 12 9
2 0 9
3 11 1 11
5 12 9 5 12 9
3 5 12 9
3 5 12 9
5 5 12 11 7 11
22 16 15 13 16 13 0 1 10 0 9 15 4 13 14 13 15 3 1 10 11 9 2
8 9 1 10 9 1 10 11 2
32 1 10 9 1 10 11 1 12 2 13 15 10 9 13 16 16 9 4 13 0 9 14 13 9 1 10 9 16 15 4 13 2
12 16 6 2 13 11 0 1 10 9 2 9 2
12 6 2 15 13 3 3 0 16 13 10 9 2
27 11 2 11 1 11 1 11 2 2 10 13 10 0 0 9 2 13 3 1 9 1 10 9 1 10 11 2
19 9 2 15 13 10 0 9 9 13 3 10 9 2 3 1 9 1 9 2
29 16 15 3 13 1 10 9 9 2 15 4 4 13 14 13 10 11 9 9 2 9 9 2 1 12 9 1 9 2
11 0 9 13 10 9 16 3 13 10 9 2
33 11 13 3 3 10 9 1 9 1 9 2 13 0 9 9 2 9 2 7 9 2 9 2 9 9 2 9 9 2 7 3 3 2
33 15 13 3 0 9 1 1 9 1 1 11 2 7 15 13 16 10 0 13 1 1 10 11 9 2 10 9 1 11 13 3 15 2
1 8
1 2
50 9 2 3 15 13 14 13 3 2 0 2 16 14 10 2 9 9 3 13 9 9 3 2 7 15 13 3 0 14 13 15 14 3 13 10 9 1 10 9 1 9 1 15 9 3 15 13 1 9 2
23 15 3 3 13 10 9 13 0 7 4 13 16 13 2 7 13 10 9 0 16 13 15 2
5 15 4 14 13 3
4 4 14 13 2
12 3 13 10 0 9 15 13 16 10 9 13 2
4 12 9 3 2
12 15 13 10 0 9 15 4 13 16 1 11 2
22 15 4 13 1 11 1 3 10 9 3 15 4 13 15 13 10 0 9 15 4 13 2
16 15 13 10 12 9 0 0 13 1 15 3 15 4 13 9 2
12 1 10 0 9 9 10 15 3 4 13 1 2
8 3 13 10 9 9 1 11 2
17 13 15 10 0 9 10 13 0 9 2 7 3 10 9 3 3 2
15 15 4 14 13 14 13 0 15 4 13 10 9 1 9 2
1 9
15 10 0 9 15 4 13 1 11 13 14 13 1 10 9 2
22 3 2 15 4 13 15 15 4 13 1 0 9 1 11 2 1 9 2 9 2 8 2
10 7 15 4 13 9 7 9 1 11 2
8 6 3 15 4 13 13 11 2
6 13 1 10 9 9 2
9 13 1 10 9 2 9 9 9 2
4 13 11 11 2
17 11 13 3 0 1 10 9 1 11 2 16 3 3 15 13 9 2
12 10 0 9 9 13 3 13 13 1 10 9 2
11 15 13 10 9 1 11 2 10 13 0 2
21 15 4 13 10 9 1 0 9 7 13 10 3 0 2 0 9 2 9 9 3 2
9 13 10 0 9 3 16 15 4 2
6 15 13 10 0 9 2
12 15 13 14 13 16 15 13 0 9 1 11 2
18 15 13 0 1 10 9 14 1 14 13 10 9 2 10 9 2 8 2
17 15 4 13 14 13 15 0 9 16 13 10 9 2 9 2 3 2
23 15 0 9 4 3 13 14 13 10 9 1 10 11 11 11 9 7 13 10 9 1 11 2
8 11 13 14 10 3 0 9 2
9 0 9 12 1 11 9 12 9 2
25 15 4 13 10 9 9 10 13 10 9 12 11 9 2 7 1 10 9 15 13 12 2 9 9 2
14 15 9 13 15 3 13 0 2 9 7 0 1 11 2
4 15 9 13 2
15 8 2 15 10 13 9 1 10 0 9 7 11 9 12 2
14 8 2 4 11 9 9 13 10 12 2 9 9 9 2
41 14 13 9 11 11 13 16 10 9 1 10 0 9 2 9 4 13 1 9 1 10 0 9 13 10 0 2 0 2 9 1 9 13 1 9 1 10 9 2 12 2
23 15 3 13 16 10 9 3 13 10 2 15 13 9 2 9 10 13 13 10 9 16 13 2
20 3 10 9 4 13 10 9 4 13 15 13 9 2 13 2 10 15 13 14 2
12 1 10 9 15 13 10 9 16 10 9 13 2
37 16 10 9 13 13 10 9 3 2 3 1 10 0 9 2 10 11 11 9 2 12 13 1 14 13 10 0 9 1 10 9 15 4 4 13 1 2
39 10 9 2 9 13 10 9 1 9 15 13 13 3 15 13 9 2 9 2 7 11 13 9 1 3 10 9 2 9 2 3 1 9 1 9 1 10 9 2
17 9 14 9 4 14 13 10 9 1 9 2 7 13 3 3 0 2
8 8 2 0 9 12 13 0 2
11 11 9 12 13 14 13 1 7 3 13 2
12 8 2 10 9 9 13 7 0 7 8 0 2
6 10 9 13 12 9 2
6 15 13 3 0 11 5
5 0 9 12 13 0
9 13 16 13 1 11 11 1 11 2
11 13 15 0 14 13 1 11 1 10 9 2
8 13 10 9 3 3 7 13 2
5 13 15 3 9 2
9 13 16 13 1 11 7 11 11 2
12 13 15 0 14 13 1 11 2 1 10 9 2
4 11 13 0 2
26 15 4 13 15 13 1 9 1 10 11 9 2 4 14 13 2 15 13 3 0 2 3 9 4 13 5
30 1 1 11 2 6 10 9 4 3 13 2 7 15 13 3 0 2 15 4 13 15 2 7 15 4 14 13 10 9 2
17 16 9 1 9 4 3 13 3 2 3 15 4 13 0 14 13 2
27 3 10 11 13 13 1 1 10 9 16 10 9 1 15 13 3 9 7 9 7 4 14 4 13 1 3 2
30 15 13 0 16 15 4 13 10 9 10 4 13 1 10 11 9 2 7 16 14 3 15 4 13 10 1 0 3 9 2
28 1 10 9 15 4 13 13 1 11 2 3 1 10 9 7 3 15 4 13 3 9 3 9 4 13 1 9 2
6 13 9 1 11 11 2
28 2 9 15 4 13 15 4 13 1 1 11 2 7 16 15 13 9 2 4 15 13 11 11 11 11 7 11 2
17 3 3 13 15 0 9 15 13 3 3 2 15 13 3 0 2 8
24 9 1 9 13 0 9 2 16 15 13 3 0 2 15 4 3 13 3 1 10 9 1 9 2
22 1 9 1 10 9 2 13 1 10 9 9 7 4 14 13 3 16 0 9 4 13 2
5 6 15 13 0 2
6 6 2 6 7 9 2
4 9 0 1 11
2 9 2
7 10 9 9 4 15 13 2
33 15 13 3 12 9 12 5 12 9 12 2 12 9 0 7 15 4 13 10 9 9 15 4 13 10 15 4 14 13 1 1 3 2
1 9
1 11
26 15 4 13 15 3 13 1 15 9 9 2 10 9 15 13 0 16 13 2 7 13 16 13 2 8 2
12 7 15 4 13 1 10 9 9 1 12 9 2
24 15 13 2 0 2 13 15 13 0 1 10 9 2 7 15 13 1 10 0 9 1 10 9 2
43 15 13 15 9 3 15 13 12 7 15 13 3 12 9 12 5 12 9 12 2 3 15 13 13 3 15 13 12 9 12 9 7 15 9 13 1 12 7 12 9 2 11 2
24 3 4 14 13 0 14 13 9 10 0 0 1 2 0 2 3 16 9 15 13 10 9 9 2
14 10 0 9 4 14 3 13 10 9 15 4 14 13 2
5 13 15 1 9 2
25 3 13 1 9 16 15 13 14 13 0 14 13 3 1 10 9 2 16 15 3 13 14 2 8 2
31 15 3 13 14 13 0 15 4 13 7 13 3 7 10 9 15 13 0 0 16 16 10 9 15 13 2 15 4 13 15 2
52 15 13 12 9 12 5 12 9 7 13 12 6 4 13 1 11 7 15 9 13 12 9 7 15 13 0 9 1 15 15 4 13 3 3 1 10 9 9 2 3 1 10 9 16 6 15 4 14 0 2 14 3
17 16 15 4 14 13 14 13 1 1 15 3 13 10 12 9 12 2
24 9 0 15 4 13 1 2 9 0 4 13 3 0 7 0 14 13 7 13 2 3 3 13 2
4 13 15 13 5
7 3 1 10 9 13 11 2
2 11 11
35 3 13 14 13 12 1 10 3 0 9 1 10 9 2 10 11 11 1 10 9 1 11 7 11 2 13 10 3 4 13 9 1 10 9 2
37 10 9 1 10 9 4 13 3 1 2 11 11 11 2 2 10 11 14 11 2 2 3 10 0 9 1 9 13 10 0 9 1 9 1 10 9 2
29 16 10 9 13 3 1 10 9 2 13 10 9 1 10 9 2 15 13 10 0 9 14 13 10 9 11 11 9 2
34 3 2 13 10 1 15 9 1 10 9 1 10 9 2 16 1 0 15 13 3 12 9 10 13 3 1 3 12 9 1 10 11 11 2
28 10 11 11 13 3 0 7 2 0 1 15 9 9 7 9 2 15 4 13 1 10 9 1 7 9 7 9 2
31 10 0 9 1 10 9 13 11 11 1 11 2 3 12 9 1 10 9 2 7 11 11 11 1 11 2 10 13 3 0 2
24 10 9 13 9 10 4 13 3 1 10 0 9 0 1 11 11 2 11 11 11 7 11 11 2
33 10 9 13 3 10 0 9 2 7 13 3 1 11 11 10 9 13 10 0 12 9 2 16 10 9 13 3 0 1 0 13 9 2
16 10 9 9 3 1 11 11 13 10 0 9 13 3 12 9 2
37 11 1 10 0 9 13 10 0 9 2 3 10 4 13 3 14 13 1 9 1 10 9 7 0 9 2 7 3 13 10 9 1 9 1 10 9 2
32 1 15 1 10 0 9 1 10 9 7 10 0 9 2 15 13 10 9 9 3 0 1 10 9 1 9 1 9 1 10 9 2
7 11 7 11 16 13 3 2
30 15 4 13 14 13 7 13 3 7 13 3 15 4 13 15 4 14 13 3 4 15 13 4 13 10 0 9 14 13 2
5 3 4 15 13 2
16 15 4 3 13 3 8 1 15 9 1 11 11 11 6 13 2
3 3 11 2
10 15 13 10 9 7 4 13 0 9 2
14 10 0 13 14 13 1 1 10 11 7 13 15 3 2
13 11 13 10 0 9 14 13 7 0 14 13 1 2
11 15 4 13 0 14 13 10 0 9 3 2
1 8
15 16 15 13 1 10 11 15 4 13 3 0 9 1 11 2
14 11 13 11 1 15 9 1 13 11 7 0 0 9 2
31 15 4 13 14 13 10 9 16 15 13 9 1 15 9 2 3 15 4 2 13 1 2 15 9 2 2 7 14 13 9 2
15 15 4 13 14 13 0 11 14 13 10 0 9 1 11 2
8 3 2 1 11 9 13 0 2
13 9 13 10 11 2 3 10 11 4 14 13 11 2
10 11 11 13 0 2 3 1 10 11 2
10 15 13 0 7 10 9 13 3 0 2
36 15 13 14 13 1 11 1 12 9 7 15 13 1 3 12 1 15 0 9 14 13 1 10 9 2 15 4 13 1 12 9 1 12 9 2 2
13 9 1 10 9 13 0 7 10 9 13 3 0 2
24 3 2 16 15 4 13 10 9 7 15 13 10 0 2 9 9 2 3 13 1 11 2 11 2
7 15 13 3 1 12 9 2
16 16 15 11 13 0 2 0 2 3 13 1 11 1 10 9 2
10 15 3 3 13 13 1 10 0 9 2
21 15 13 15 1 9 12 1 11 2 11 7 15 13 10 3 0 9 1 15 9 2
13 4 10 11 13 14 4 13 3 14 13 1 11 2
9 15 13 10 0 9 1 10 11 2
9 15 13 10 9 13 1 0 9 9
1 8
22 2 0 3 1 9 9 2 10 11 11 11 2 11 2 13 10 9 14 3 13 9 2
45 3 13 1 10 11 11 11 2 11 14 11 11 2 11 14 11 11 2 11 14 11 11 7 0 0 9 1 2 15 13 14 13 9 1 15 9 7 15 4 14 13 15 13 2 2
8 13 15 13 15 3 3 3 2
18 15 13 10 0 9 3 3 2 3 2 15 13 10 9 9 9 2 2
1 8
11 2 15 13 10 0 9 1 11 11 11 2
9 6 13 2 15 13 10 0 9 2
13 15 13 10 0 9 2 1 10 9 1 10 9 2
9 15 13 10 9 1 10 9 2 2
26 10 0 9 1 11 4 13 15 13 10 0 9 1 10 11 1 11 7 9 13 1 15 13 10 9 8
39 3 13 16 15 4 14 3 13 10 9 0 9 16 15 9 14 4 13 2 15 0 9 2 9 2 9 9 2 8 7 16 15 4 14 13 16 13 9 2
27 10 9 4 14 13 14 13 15 2 10 0 9 1 10 9 13 14 13 15 9 3 14 13 15 9 7 9
8 13 10 11 11 14 13 15 8
2 6 2
9 11 3 13 1 10 9 1 9 2
4 12 5 9 2
11 13 1 10 9 7 13 1 15 11 9 2
50 15 13 10 0 9 1 10 11 7 2 11 11 11 2 2 15 13 12 5 10 9 2 16 10 0 9 13 2 13 1 10 7 10 9 1 10 9 2 15 13 14 15 7 15 15 4 13 14 13 2
19 10 0 9 1 10 11 9 13 15 2 15 13 10 0 1 11 2 3 2
1 8
9 3 4 15 13 15 9 9 13 2
32 15 13 10 0 9 7 9 15 13 3 10 9 7 3 13 9 3 3 16 15 13 4 9 13 15 13 1 3 14 13 15 13
15 15 13 10 9 2 15 4 13 14 2 13 2 15 13 2
11 15 13 16 13 14 13 12 9 4 13 2
5 15 4 14 13 2
7 3 15 13 10 0 9 2
16 13 16 15 12 3 3 13 10 0 2 3 15 13 9 3 2
19 3 15 13 14 13 0 2 3 3 2 0 0 2 7 0 0 14 13 2
22 15 4 13 3 12 2 12 1 15 0 9 9 2 3 12 5 12 9 1 10 9 2
4 3 10 9 2
15 0 9 2 10 0 9 2 0 9 9 7 3 0 9 2
16 10 9 13 15 15 13 14 13 2 7 15 13 0 1 15 2
13 13 15 0 2 7 15 4 13 3 15 13 0 2
13 15 4 14 13 15 13 2 15 4 3 13 15 2
1 11
10 9 9 13 14 10 0 9 14 13 2
14 0 1 10 9 12 13 3 0 1 13 1 10 0 2
23 9 13 10 12 10 13 14 3 0 7 13 15 0 1 10 9 9 1 12 5 12 9 2
33 10 9 4 13 10 9 9 0 0 1 12 9 2 7 10 9 1 15 2 7 3 3 12 9 0 0 1 12 0 14 13 1 2
9 10 9 9 4 13 12 5 12 2
27 3 13 10 12 1 10 9 9 3 0 9 2 9 7 2 7 9 16 15 4 13 1 12 5 12 9 2
6 3 13 10 0 9 2
26 15 4 14 13 3 3 7 15 4 13 3 10 0 12 4 13 1 12 1 9 9 16 15 4 13 2
14 3 10 9 14 0 9 13 2 15 13 0 14 13 2
13 10 12 13 15 9 1 10 9 15 13 1 15 2
8 13 10 9 9 1 1 12 9
9 6 13 1 15 9 14 9 9 2
12 15 13 10 12 12 2 12 9 0 0 9 2
29 3 15 4 13 10 9 13 10 0 9 16 15 3 13 12 9 9 7 15 13 15 4 13 15 3 13 12 9 2
8 3 15 4 4 13 10 9 2
12 15 4 13 13 10 10 9 9 7 3 10 2
13 15 4 3 13 1 10 9 7 3 15 13 3 2
23 15 4 14 13 10 9 14 13 15 1 10 9 3 3 7 15 4 13 14 13 10 9 2
14 15 13 14 13 10 9 12 5 12 9 10 9 3 2
14 15 4 13 10 9 7 4 15 13 10 9 9 3 2
28 15 13 15 7 13 14 13 15 7 15 4 14 13 3 15 4 13 0 14 13 15 1 1 9 5 6 13 2
20 3 1 10 2 15 13 3 0 14 13 15 4 13 10 9 1 15 9 2 5
9 0 9 13 10 9 1 0 9 2
25 9 7 0 9 9 13 12 0 9 2 7 15 3 13 0 9 2 16 0 9 1 9 4 13 2
25 16 15 13 9 1 10 9 2 7 10 9 13 14 13 1 9 2 3 15 13 3 10 0 9 2
15 7 15 9 4 13 10 9 1 9 2 7 15 13 0 2
32 13 10 9 15 9 4 3 13 12 9 2 15 4 13 10 0 9 9 4 13 9 9 2 10 0 4 13 1 0 0 9 2
26 9 1 15 4 13 0 14 13 2 7 16 15 13 0 1 15 9 15 4 3 13 14 13 10 9 2
8 9 2 0 9 2 7 9 2
19 9 4 13 3 10 9 10 10 9 3 13 1 4 13 1 10 9 9 2
23 15 13 15 13 3 0 2 7 13 15 1 10 9 13 10 0 9 15 4 13 1 15 2
14 1 10 9 13 0 15 13 9 1 9 0 1 15 2
10 15 13 14 13 1 11 13 9 9 2
11 15 13 3 12 9 16 12 9 13 9 2
7 4 15 13 1 12 9 2
33 13 1 10 11 7 11 11 9 9 1 8 2 15 13 2 9 2 15 4 13 10 0 9 16 15 9 14 13 0 1 13 2 2
17 3 2 10 0 9 9 3 13 16 2 10 0 9 9 13 12 2
6 10 9 9 4 13 2
12 15 4 13 1 0 9 1 10 0 9 2 2
12 10 11 11 9 13 15 0 9 1 0 9 2
21 7 1 10 9 15 13 15 9 7 10 9 15 13 2 10 0 9 4 13 3 2
9 3 2 10 9 13 1 15 9 2
16 7 15 13 0 16 15 13 1 10 9 14 13 10 0 9 2
10 3 13 13 3 3 1 10 0 9 2
16 0 9 2 15 13 10 9 9 13 1 11 11 11 1 8 2
6 3 13 15 15 13 3
21 2 8 2 4 15 13 1 10 11 11 9 3 16 15 13 0 1 12 9 2 2
58 2 16 10 11 11 11 11 13 16 10 9 9 4 14 3 13 15 9 14 13 3 13 1 11 2 10 11 11 11 11 4 13 15 7 15 0 9 2 13 1 1 13 9 2 7 13 15 9 3 16 15 13 0 1 12 9 2 2
11 13 10 0 9 1 10 9 9 1 9 2
5 6 15 4 13 2
14 10 9 9 13 1 10 9 14 13 1 10 0 9 2
25 15 9 4 3 13 1 10 9 1 9 2 3 10 1 15 3 2 13 1 9 2 1 10 9 2
8 13 3 2 13 1 15 9 2
4 9 1 11 2
19 12 13 10 0 9 2 9 1 15 4 13 1 10 2 0 9 9 2 2
14 3 13 10 2 9 2 16 15 4 13 14 4 13 2
2 11 11
2 11 2
11 15 13 0 7 4 14 13 15 14 13 2
3 6 13 2
26 6 2 3 15 9 4 4 13 15 14 13 15 9 9 1 10 0 9 7 15 3 13 3 1 15 2
44 2 15 3 13 15 13 15 14 13 12 1 10 9 9 9 3 2 3 15 3 13 15 2 7 15 13 10 9 9 1 11 11 13 15 10 9 9 1 15 9 9 1 11 2
5 15 13 3 0 2
9 15 13 15 13 1 11 7 3 2
25 3 15 13 13 7 3 15 13 10 9 2 15 13 1 8 9 11 7 13 3 8 9 9 2 5
20 3 15 13 15 3 3 3 13 13 7 3 3 3 13 3 13 1 10 9 2
14 2 15 13 1 11 3 2 15 13 0 7 0 3 2
19 4 14 13 15 0 15 13 14 13 2 7 1 12 9 5 15 13 3 2
20 15 4 13 10 12 9 9 3 1 10 0 9 1 11 7 13 3 12 9 2
16 2 6 2 14 13 14 13 0 7 13 1 7 15 13 3 2
11 4 9 6 13 15 13 0 1 10 9 2
6 3 3 15 4 13 2
12 13 10 12 9 15 0 16 3 13 3 3 2
35 7 15 4 13 0 12 9 16 15 4 0 13 1 10 9 1 0 9 2 15 4 13 14 13 3 13 0 15 13 10 9 14 13 2 5
15 6 2 15 13 2 15 4 14 13 14 13 0 1 15 2
11 3 3 15 13 14 13 1 11 1 11 2
16 7 2 13 3 12 9 13 15 13 15 15 13 1 15 9 2
9 2 9 0 4 13 2 2 9 2
24 13 15 16 15 4 2 7 3 16 15 9 13 15 15 4 13 3 1 10 0 9 1 9 2
16 16 15 4 14 13 15 2 15 4 3 13 12 9 2 13 2
8 13 15 13 10 9 1 9 2
7 2 1 10 0 9 2 2
6 15 13 0 0 11 2
10 13 10 9 1 15 2 15 4 13 2
48 8 2 10 11 11 13 10 0 9 1 10 11 2 10 9 1 0 0 9 7 9 1 11 10 13 10 9 1 10 9 1 10 0 9 1 3 12 2 13 10 9 1 0 7 0 0 11 2
28 10 9 11 13 1 9 10 0 9 10 13 1 9 1 10 0 9 2 1 10 9 1 9 0 1 11 11 2
57 16 10 9 1 10 9 10 4 13 3 1 10 0 9 1 0 9 7 9 4 4 13 1 10 0 9 1 10 0 9 2 0 9 1 0 9 7 9 13 3 0 2 10 11 4 14 13 1 0 9 1 10 9 1 10 9 2
40 10 9 11 2 11 1 11 2 13 2 9 2 2 7 10 9 13 3 13 1 10 13 9 1 10 9 1 0 9 1 10 9 10 11 9 13 10 11 11 2
29 10 9 2 16 0 2 4 13 1 10 0 2 7 1 10 0 9 1 10 9 9 4 3 13 1 10 11 11 2
29 8 2 10 9 0 11 2 1 9 9 2 13 10 9 9 13 14 13 10 9 1 10 0 9 1 10 0 11 2
51 10 0 11 9 4 3 13 14 13 1 10 9 2 1 11 14 9 1 10 11 11 1 11 7 10 9 1 11 11 11 1 11 2 7 14 4 13 1 12 1 10 9 1 11 1 10 9 1 11 11 2
36 10 9 4 3 13 1 11 2 8 2 1 10 0 0 9 2 7 13 15 9 1 10 2 0 9 2 1 9 7 9 13 1 11 11 11 2
39 2 8 2 1 10 0 12 9 2 9 1 10 9 4 4 3 13 1 0 9 9 16 13 0 9 2 13 0 9 2 7 13 3 1 10 0 0 9 2
3 2 8 2
4 13 15 13 2
20 15 13 0 7 15 4 13 1 10 11 1 10 0 9 2 15 4 15 13 2
36 15 3 13 14 13 1 10 10 0 15 4 13 1 10 11 3 16 16 15 13 15 13 3 13 1 10 9 7 16 13 1 9 9 7 9 2
12 4 15 13 15 9 14 9 3 1 10 9 2
14 15 4 13 16 11 3 13 10 12 9 9 14 9 2
12 4 15 13 14 13 1 10 0 9 3 3 2
3 9 9 2
3 9 9 2
13 7 4 15 3 13 15 9 7 13 1 10 9 2
30 15 4 13 1 10 9 10 13 16 10 0 9 13 10 9 1 9 7 0 13 15 13 10 9 9 3 13 10 9 2
38 15 3 13 10 9 15 14 13 7 13 1 7 13 3 14 13 0 9 1 10 1 10 9 13 1 10 9 2 10 15 3 4 14 13 10 9 1 2
20 15 13 3 0 16 15 13 10 9 15 14 13 1 7 13 9 14 13 3 2
23 10 0 9 4 13 15 3 1 10 9 2 15 13 10 9 1 10 9 2 1 12 9 2
13 15 13 10 0 9 7 9 9 7 9 1 15 2
13 15 4 14 13 14 13 10 9 14 13 0 9 2
1 8
27 3 13 10 9 1 10 11 1 11 9 9 2 10 4 13 15 10 10 9 10 15 13 2 13 9 9 2
4 15 13 0 2
16 15 3 13 0 1 12 9 1 10 9 3 15 13 10 11 2
18 15 4 13 0 1 3 10 9 2 16 15 4 13 3 1 12 9 2
13 15 4 3 13 1 10 0 9 16 15 13 3 2
11 15 13 14 0 3 3 15 13 10 9 2
12 15 4 13 10 0 9 2 3 10 9 3 2
24 15 13 11 2 11 2 7 11 11 14 3 3 2 7 15 4 13 3 3 7 1 0 9 2
18 3 13 9 0 16 15 4 13 14 4 13 2 7 15 4 13 0 2
6 10 0 3 13 15 2
15 15 4 15 13 16 15 13 10 9 9 7 10 9 9 2
25 15 13 10 9 9 7 10 9 9 15 13 12 9 15 4 10 9 9 7 10 9 9 4 13 2
21 16 15 13 10 9 1 15 9 15 4 13 14 13 15 14 13 15 1 15 9 2
14 10 9 13 1 9 4 13 10 13 2 9 2 9 2
22 15 13 10 9 1 9 1 9 1 10 9 7 9 2 3 10 9 4 13 1 9 2
28 15 4 14 13 10 9 9 7 9 15 4 13 1 3 15 4 14 13 10 9 15 9 4 13 0 14 13 2
13 3 2 15 4 13 10 9 15 4 2 4 13 2
3 9 9 2
5 9 13 0 9 2
5 9 13 0 9 2
18 10 9 1 10 9 4 13 0 9 2 16 0 9 13 10 0 9 2
13 9 11 2 9 13 0 9 9 2 10 13 0 2
11 9 13 0 9 10 4 13 0 7 0 2
12 10 9 0 7 0 0 9 13 10 0 9 2
10 9 4 13 0 7 0 1 10 9 2
28 9 2 9 2 16 15 9 13 10 9 2 9 10 9 4 13 10 9 3 3 2 16 10 9 13 3 0 2
19 0 9 2 9 2 9 4 13 0 9 2 9 16 15 13 3 3 0 2
18 9 2 9 4 3 13 10 0 9 1 16 15 13 10 3 0 9 2
28 9 9 2 9 13 9 9 10 13 3 3 12 9 9 2 9 7 9 2 9 13 3 3 2 7 13 0 2
20 3 13 1 10 11 15 4 13 10 9 2 9 2 9 2 7 0 13 9 2
8 12 9 2 9 13 12 9 2
5 9 13 12 9 2
25 13 3 2 12 9 13 3 0 2 9 4 13 14 13 10 0 9 1 10 2 7 3 12 9 2
11 9 9 13 0 9 2 7 3 0 13 2
19 9 13 0 9 16 15 13 0 2 4 13 3 2 7 13 0 1 9 2
3 0 9 2
3 11 2 11
13 15 13 10 9 1 15 9 9 1 15 11 9 2
8 15 4 15 13 1 10 9 2
21 8 8 8 15 13 10 9 1 15 9 9 1 15 11 9 2 13 9 3 2 2
8 15 4 15 13 1 10 9 2
17 10 9 13 14 10 0 2 7 10 9 13 1 0 1 15 9 2
24 13 10 9 3 15 4 14 13 10 9 4 14 13 15 0 9 2 15 13 1 15 0 9 2
20 15 13 14 13 1 0 9 2 9 2 9 2 7 13 16 13 10 9 3 2
21 2 9 2 7 15 4 13 3 0 1 9 2 16 15 4 13 0 1 15 9 2
12 6 2 15 4 13 15 3 0 9 9 3 2
20 3 15 13 0 16 9 13 15 13 15 9 1 10 9 7 15 13 14 15 9
12 3 0 2 7 3 0 0 9 1 15 9 2
3 1 9 2
21 1 10 9 1 10 9 2 10 9 15 4 13 1 13 1 9 0 1 10 9 2
22 15 13 3 10 0 9 9 1 10 9 9 7 15 13 1 10 9 9 1 10 9 2
36 1 10 9 9 2 1 10 9 2 15 13 10 9 1 10 9 13 3 2 10 9 1 9 1 10 0 0 9 7 15 13 1 10 9 9 2
23 1 10 9 1 10 9 2 10 13 9 1 10 9 13 3 0 3 3 1 10 9 9 2
30 3 2 10 12 13 14 15 9 2 15 4 13 13 10 0 9 16 15 4 14 13 13 15 1 1 10 9 13 0 2
8 15 4 13 10 9 2 3 2
42 15 9 13 14 13 0 9 16 15 4 13 1 1 10 9 7 16 0 2 13 1 10 9 2 13 1 10 9 2 13 15 15 13 14 13 14 13 0 1 0 9 2
15 13 10 3 0 9 13 3 0 16 13 1 0 9 9 2
23 15 4 13 10 0 0 9 13 15 16 15 13 9 1 10 9 15 4 14 13 3 3 2
8 15 13 10 0 9 1 11 2
18 3 3 16 15 13 0 15 3 0 9 4 13 10 2 9 9 2 2
26 1 10 15 9 15 4 3 13 9 1 15 7 4 3 13 1 10 0 9 3 15 13 15 1 9 2
21 16 10 9 13 2 15 9 4 2 13 2 1 15 9 1 3 12 5 12 9 2
34 1 10 9 9 4 13 1 10 9 2 13 15 9 1 10 0 7 15 9 7 13 10 9 1 9 1 9 1 10 9 7 10 9 2
20 10 9 3 13 10 9 9 3 9 7 9 13 1 1 10 9 1 10 9 2
16 9 13 0 7 3 7 3 1 10 9 1 11 7 11 3 2
7 7 3 3 1 10 9 2
39 10 0 0 9 15 4 13 13 16 1 10 9 1 11 12 9 1 10 9 4 3 13 1 10 9 10 9 1 10 9 2 10 9 13 1 10 0 9 2
15 10 0 9 2 7 10 13 9 1 15 2 13 10 11 2
44 10 11 13 10 9 13 1 10 9 1 10 0 9 10 13 7 13 10 9 1 9 2 13 1 3 2 2 1 10 9 14 13 1 10 0 9 1 9 10 11 4 13 1 2
33 11 13 10 9 14 13 0 2 0 7 1 10 9 1 10 9 9 2 13 10 13 12 12 9 3 13 11 11 1 10 0 9 2
19 15 8 15 13 12 7 13 16 10 9 13 0 14 13 1 10 0 9 2
30 10 11 11 7 10 9 1 11 11 4 4 13 1 10 14 14 13 10 0 9 7 3 13 10 9 14 4 13 12 2
29 10 9 1 10 9 1 11 4 3 3 13 1 11 1 10 11 7 1 9 1 15 13 10 0 13 9 1 11 2
6 9 9 7 10 9 2
26 10 0 9 15 13 1 15 9 13 2 15 13 9 9 1 11 2 9 9 7 9 2 9 1 11 2
6 11 9 1 11 9 2
12 4 9 13 9 1 10 9 9 16 9 13 2
12 4 9 13 9 1 10 9 9 16 9 13 2
30 15 13 0 1 15 2 16 3 15 13 10 0 1 9 9 1 15 9 7 15 4 14 13 16 13 10 9 1 9 2
43 15 13 16 10 9 2 3 13 10 9 2 8 2 4 13 14 13 10 9 9 9 13 1 9 2 0 1 0 9 2 9 9 2 7 0 13 9 10 13 4 14 13 2
31 3 3 16 15 13 2 10 9 4 13 3 0 2 7 15 9 13 2 4 9 3 13 10 9 13 1 10 9 1 9 2
13 3 2 4 9 13 9 1 9 1 15 2 9 2
34 16 3 2 3 4 15 13 16 16 15 13 10 0 9 7 15 9 2 9 2 9 13 1 10 0 9 1 15 15 4 3 13 0 2
23 15 4 14 13 2 15 4 14 3 13 0 9 2 7 15 4 14 13 15 1 15 9 2
30 3 2 15 4 14 13 16 0 9 4 13 9 1 10 0 9 2 15 13 0 15 4 13 3 2 7 13 15 0 2
5 3 15 1 9 2
6 4 9 13 13 9 2
19 6 2 9 13 10 9 1 13 9 10 4 13 3 14 13 10 13 9 2
32 10 9 4 13 1 10 9 1 3 12 9 2 10 13 3 0 15 13 14 13 16 15 14 13 15 1 10 13 2 0 9 2
32 1 10 9 2 13 9 13 10 9 16 13 10 0 0 0 9 16 15 9 9 13 14 13 1 10 9 1 12 1 12 9 2
16 3 15 13 10 9 13 3 7 8 3 15 13 0 1 15 2
20 3 9 13 16 16 15 9 13 14 13 9 2 15 13 3 1 1 10 9 2
18 13 13 10 9 14 0 9 2 7 15 4 13 15 1 10 9 9 2
4 6 15 13 2
22 15 13 3 0 16 15 4 13 9 1 10 9 9 16 15 9 13 9 1 10 9 9
11 3 0 4 15 4 13 1 1 9 9 2
26 15 13 12 9 13 1 9 1 10 12 9 9 2 7 10 9 13 3 12 9 3 16 3 15 13 2
29 10 9 3 15 4 13 13 14 0 14 13 14 13 15 3 3 2 7 15 4 14 13 10 9 16 13 15 15 2
18 3 15 13 14 13 9 2 7 0 9 2 14 13 15 1 10 9 2
18 16 15 13 3 0 15 13 0 14 13 2 15 13 10 0 9 9 2
11 15 13 10 9 10 13 5 12 1 9 2
4 13 1 0 2
61 0 14 13 2 7 15 13 15 4 13 14 13 1 9 9 1 10 0 9 10 15 4 13 7 13 10 9 1 15 2 7 10 1 9 1 10 9 14 9 7 9 2 16 15 13 0 14 13 9 1 10 7 0 2 15 4 13 10 9 3 2
9 13 16 15 13 15 15 13 1 2
13 12 9 13 14 0 2 7 15 4 13 0 9 2
24 10 9 13 0 14 13 15 9 2 7 15 3 13 0 9 10 13 14 10 0 1 10 9 2
32 13 2 13 9 1 10 9 2 0 9 2 0 9 3 1 0 9 4 3 13 13 0 2 1 3 3 0 2 1 15 9 2
20 15 13 15 9 13 1 11 1 11 7 15 13 1 10 0 2 0 9 9 2
11 15 13 0 3 15 13 3 7 13 9 2
41 1 3 2 15 3 13 10 0 9 9 9 1 9 15 13 1 15 9 14 13 10 9 1 15 2 13 10 0 9 1 9 2 7 15 9 3 13 3 0 9 2
18 10 9 15 4 13 13 1 15 1 3 13 0 7 0 3 15 13 2
11 15 4 13 11 11 11 7 13 10 9 2
26 3 16 15 4 14 13 14 13 15 2 15 4 13 15 10 9 1 15 15 4 13 7 15 13 0 2
4 13 9 3 2
18 13 0 10 9 9 15 13 4 13 2 13 7 13 9 1 0 9 2
6 4 15 13 15 3 2
10 15 13 14 13 10 9 1 10 9 2
9 15 13 3 1 10 9 16 0 2
22 3 3 16 15 13 3 1 10 0 9 3 0 4 15 13 15 4 13 3 10 9 2
17 3 13 15 10 9 14 3 3 13 10 9 15 13 14 13 1 2
7 6 15 4 13 10 9 2
17 7 16 14 3 13 6 7 15 13 15 13 6 12 1 3 3 2
13 8 2 3 13 10 9 10 13 9 9 13 9 2
1 8
30 9 13 2 3 2 4 3 13 1 12 9 1 10 9 2 7 15 4 3 13 10 0 2 0 9 2 9 1 9 2
21 2 12 9 1 10 9 4 13 0 3 2 3 9 9 13 15 0 14 13 3 2
19 15 4 13 0 14 13 3 1 10 9 16 15 13 0 9 1 11 2 2
24 8 2 0 16 13 15 0 9 7 9 2 15 4 14 13 10 9 15 4 13 15 0 9 2
3 0 9 2
17 0 9 9 1 0 1 10 0 9 9 2 3 12 9 1 9 2
21 13 1 15 0 15 4 13 14 13 0 16 9 4 13 1 10 9 1 0 9 2
8 10 9 14 13 9 1 9 2
46 13 3 12 9 1 9 16 10 9 9 13 9 3 1 10 9 8 3 1 11 2 11 2 2 11 1 11 2 11 2 2 11 1 11 2 11 2 2 11 1 11 1 11 9 8 2
17 6 15 13 0 1 10 9 9 2 3 13 1 10 3 0 9 2
22 3 2 15 4 13 16 16 15 13 12 9 1 10 9 2 3 16 15 13 3 15 2
16 3 10 9 15 13 2 13 15 13 2 5 12 12 3 3 2
62 7 6 15 4 14 13 10 0 16 15 13 0 0 9 1 10 9 1 9 3 3 1 9 2 6 13 10 11 11 9 2 3 13 1 11 7 13 15 1 3 7 13 1 11 3 13 1 11 14 13 10 11 16 13 1 11 14 13 10 0 9 2
14 13 10 11 11 11 11 3 0 3 1 10 0 9 2
2 6 2
42 15 4 13 10 0 0 9 1 10 11 11 11 1 10 0 9 2 10 11 3 13 10 0 9 1 11 3 1 11 2 15 13 9 1 0 15 4 4 13 1 11 2
14 10 0 11 11 7 10 0 9 1 10 11 13 0 2
8 10 11 13 3 0 2 0 2
15 16 10 11 11 7 11 13 3 2 15 13 1 10 9 2
51 3 2 10 11 11 4 13 3 0 3 1 10 0 9 2 9 4 4 13 14 13 10 0 9 7 15 13 16 0 9 3 3 13 0 7 0 1 10 9 13 11 3 15 13 15 10 9 13 9 1 2
35 10 0 9 4 14 3 13 1 9 3 2 7 3 2 15 4 3 13 10 9 9 1 10 9 1 3 1 10 3 0 2 0 9 9 2
20 11 11 13 3 0 7 0 1 10 13 0 11 11 9 13 1 1 0 9 2
17 15 13 14 3 3 16 0 9 9 1 9 13 14 13 10 9 2
15 15 3 13 0 11 9 2 0 9 2 0 9 1 3 2
5 15 13 10 9 2
12 0 9 4 14 13 1 10 9 1 10 9 2
14 15 4 14 13 0 9 1 0 9 1 10 0 9 2
11 15 13 0 9 13 1 10 0 9 3 2
17 15 13 0 0 9 1 10 9 1 9 3 0 9 4 14 13 2
22 3 11 13 10 0 9 2 0 9 7 13 9 1 1 9 7 9 9 1 10 9 2
24 11 11 4 13 1 10 0 7 0 9 1 3 0 9 1 1 10 0 9 15 13 0 9 2
17 15 4 3 13 10 0 2 0 0 9 16 11 4 13 1 11 2
26 15 13 10 0 0 9 1 10 9 16 15 13 3 7 15 4 14 13 10 9 16 11 11 4 13 2
16 11 11 13 3 0 7 0 7 0 1 10 9 1 9 3 2
15 10 9 1 11 11 13 3 0 1 11 11 1 10 9 2
24 9 2 15 9 4 14 13 0 3 15 4 13 10 3 0 9 1 9 0 15 13 10 9 2
7 4 9 7 9 13 3 2
22 15 4 13 16 13 10 9 1 10 9 2 7 15 9 13 16 15 13 14 13 3 2
18 15 3 13 12 9 10 4 13 1 10 9 1 15 9 2 9 9 2
51 15 13 3 10 0 9 9 10 15 4 13 1 10 0 9 9 4 13 3 3 7 15 4 13 16 13 10 9 1 10 9 1 10 9 2 7 13 10 9 1 10 9 7 10 9 1 10 9 1 9 2
21 3 2 1 10 9 9 4 15 13 0 16 10 9 14 13 3 1 1 10 9 2
29 15 13 10 9 9 1 9 7 9 1 10 9 2 7 15 13 9 10 10 9 4 14 13 0 14 13 3 3 2
21 3 2 4 9 7 9 13 3 3 3 16 15 13 0 9 1 15 9 7 9 2
45 2 10 9 9 4 13 10 9 3 0 0 1 10 9 2 10 9 4 14 13 0 14 13 1 10 9 9 2 3 2 13 15 0 16 10 9 3 13 10 0 9 1 9 9 2
14 15 0 9 13 15 10 0 9 2 7 15 13 0 2
9 15 3 13 14 13 0 2 9 2
44 6 2 7 13 0 16 15 9 13 3 9 2 15 13 3 9 2 2 9 4 13 9 7 9 15 13 13 2 3 13 0 1 15 2 9 13 0 1 3 10 9 1 9 2
25 1 15 9 9 2 7 9 2 13 3 0 1 9 2 9 9 2 9 2 9 2 9 2 8 2
10 13 0 3 14 13 15 9 0 9 2
45 15 13 15 13 1 0 9 7 15 13 0 1 9 2 3 10 9 2 4 14 13 10 1 15 1 12 9 16 9 9 13 0 1 15 1 9 2 0 9 4 13 9 1 15 2
12 3 2 4 14 13 10 1 15 1 12 9 2
3 0 9 2
26 6 15 13 7 9 4 3 13 10 9 7 10 9 4 13 1 3 7 10 9 4 13 10 0 9 2
17 3 13 3 0 7 10 9 4 13 0 1 9 7 0 1 9 2
16 9 4 13 3 3 4 14 13 0 16 9 4 13 1 9 2
13 9 13 0 7 4 13 9 3 13 1 1 15 2
6 13 9 4 14 13 2
15 15 9 7 15 4 13 14 13 9 14 13 10 0 9 2
72 15 4 13 10 9 1 0 2 15 13 10 9 9 9 1 10 9 1 10 9 13 10 9 1 9 9 1 10 9 1 15 1 10 9 1 10 9 2 13 10 9 1 9 9 2 13 10 9 1 9 13 15 1 7 13 9 1 10 9 1 10 9 2 9 13 3 0 7 4 14 13 2
5 15 4 15 13 3
28 15 4 13 14 13 1 9 3 0 1 9 2 9 2 9 7 9 2 15 10 13 10 3 3 0 9 9 2
8 15 4 3 13 10 0 9 2
17 0 9 13 3 0 7 3 15 13 13 9 7 13 9 7 9 2
20 3 16 15 4 13 15 2 15 13 15 13 10 9 16 13 15 7 13 15 2
15 15 13 3 3 0 1 10 9 2 7 1 9 7 9 2
15 3 10 9 9 4 13 15 2 16 15 4 14 13 9 2
17 9 13 0 16 15 15 4 13 2 7 15 13 1 10 9 9 2
28 15 4 13 14 13 1 9 3 0 1 9 2 9 2 9 7 9 2 15 10 13 10 3 3 0 9 9 2
22 9 13 10 3 0 9 9 1 9 7 15 4 13 15 9 3 4 14 13 0 0 2
35 15 13 15 3 4 13 9 16 15 4 13 1 9 10 4 14 13 3 0 1 0 9 2 3 1 9 15 13 9 2 3 9 9 2 2
35 15 4 13 10 0 9 1 9 9 2 7 3 13 14 13 15 0 9 2 7 15 13 15 9 13 3 3 0 7 4 14 13 0 0 2
41 15 4 13 0 9 1 9 1 10 9 1 10 0 9 9 2 3 0 1 10 9 9 2 7 15 4 4 13 1 10 9 9 15 4 13 1 10 9 9 2 2
7 15 13 9 7 13 15 8
18 9 13 1 3 1 12 11 10 13 10 0 0 9 2 3 3 0 2
1 8
29 15 4 13 0 14 13 10 9 1 15 9 13 2 7 15 4 13 10 10 9 1 9 7 10 9 1 13 9 2
14 15 13 9 1 10 9 7 10 9 15 13 8 7 8
13 4 10 11 9 7 15 9 7 9 13 0 9 2
14 10 9 1 15 13 11 1 11 16 1 9 0 9 2
15 15 4 14 13 10 9 7 9 9 10 13 0 13 9 2
13 15 13 0 1 15 9 16 15 3 13 0 9 2
37 3 16 15 13 10 9 1 10 9 14 15 4 14 13 3 15 13 1 10 9 2 1 9 10 9 4 4 4 13 13 10 9 13 16 13 9 2
37 15 13 3 14 3 10 9 16 13 9 2 9 7 3 4 13 14 13 0 13 9 2 7 10 9 7 15 9 4 14 4 4 13 1 13 9 2
19 9 1 11 4 13 14 13 9 9 7 4 13 9 1 9 1 10 9 2
16 15 10 13 13 10 9 3 13 10 9 7 9 16 1 9 2
8 3 9 13 14 13 13 9 2
23 15 13 14 0 16 10 9 13 14 13 16 13 9 16 10 9 4 13 0 9 1 15 2
31 15 13 15 13 3 0 16 3 10 9 4 13 3 3 12 0 9 7 9 7 3 12 9 10 0 9 9 4 13 0 2
12 3 15 13 1 11 2 10 10 9 13 0 2
29 15 4 14 13 0 9 2 3 13 15 2 15 13 1 9 10 13 14 10 9 9 2 15 13 9 1 0 9 2
25 15 4 14 13 1 15 9 7 13 15 13 7 13 10 9 1 9 10 9 15 13 14 13 15 2
51 3 15 13 1 10 9 2 15 13 1 15 9 1 9 7 15 9 2 16 15 4 14 13 15 2 15 13 3 14 13 3 1 10 9 2 7 15 13 15 9 9 13 3 0 14 13 1 2 6 2 2
42 9 7 9 3 13 10 0 9 1 0 9 9 3 2 15 3 13 0 1 9 9 2 0 1 13 9 2 0 1 0 9 2 8 2 3 1 9 9 7 9 9 2
2 6 2
13 14 13 9 9 2 0 9 13 0 7 0 9 2
13 11 13 12 2 7 10 11 4 13 10 0 9 2
11 15 4 13 11 9 1 10 9 1 9 2
11 15 4 14 13 10 9 13 14 13 3 2
17 16 9 13 15 13 10 9 9 3 15 4 13 13 0 0 9 2
13 3 14 13 15 9 14 13 15 13 10 9 9 2
9 15 4 14 13 9 1 9 9 2
17 3 15 13 15 9 15 13 15 4 3 13 10 9 1 15 9 2
12 15 13 10 9 1 9 7 4 3 13 12 2
19 15 13 10 15 9 7 13 3 13 14 13 12 2 15 13 12 1 10 9
7 13 10 9 1 15 9 2
20 3 16 15 13 3 0 9 7 9 15 4 13 16 13 10 9 15 4 13 2
20 13 15 15 13 1 12 9 10 9 2 16 3 10 0 2 14 13 15 0 2
26 13 0 1 10 9 14 13 16 3 16 15 4 14 13 1 15 15 16 15 13 0 14 13 1 15 2
37 16 15 4 13 15 1 10 9 13 14 13 15 1 10 9 9 7 13 12 1 10 9 14 13 10 9 13 15 9 3 0 7 0 15 4 13 2
13 3 3 13 14 13 15 9 14 13 15 10 9 2
29 15 9 13 0 1 9 3 15 3 13 2 15 13 15 1 12 1 15 9 9 9 7 15 13 1 9 1 15 2
18 13 0 2 7 4 14 13 15 1 15 16 15 4 13 15 3 3 2
3 0 9 2
13 15 0 13 15 9 14 13 15 13 10 9 9 2
5 8 2 13 0 2
24 13 10 15 9 16 4 13 2 13 9 1 10 13 9 2 13 15 9 0 2 7 3 3 2
26 13 2 1 15 9 14 9 2 16 15 2 7 15 2 4 13 10 9 3 13 9 1 15 0 9 2
18 8 2 13 1 2 7 13 2 16 16 15 13 0 1 15 0 9 2
6 8 2 13 1 15 2
21 13 14 13 0 9 2 13 1 15 9 1 10 9 1 0 9 2 9 1 15 2
7 8 2 13 10 9 9 2
57 16 15 4 13 10 9 1 10 9 2 7 10 10 9 13 14 13 0 1 16 15 4 13 7 10 2 15 4 13 0 14 13 15 9 16 2 13 15 10 0 9 2 3 15 4 14 13 0 14 13 15 16 13 10 0 9 2
16 1 10 9 9 2 13 15 16 13 1 10 9 9 1 15 2
14 16 15 13 3 2 13 16 15 4 13 10 9 9 2
16 16 15 4 13 15 2 13 14 13 15 14 13 2 13 15 2
13 15 9 14 9 13 3 0 2 15 4 15 13 2
20 3 9 15 13 10 9 9 1 15 0 9 9 11 2 13 1 11 11 2 2
18 0 9 15 13 10 9 9 15 13 10 9 7 15 9 13 15 3 2
14 7 9 2 15 13 10 9 7 13 16 15 13 0 2
17 15 3 4 13 15 9 16 15 13 3 10 0 0 2 13 9 2
16 3 15 0 9 13 1 15 2 3 4 15 13 10 9 1 2
31 16 15 13 15 1 10 9 7 3 0 15 4 13 3 2 4 15 13 15 1 10 9 16 10 9 4 13 1 15 9 2
13 15 3 4 13 9 7 9 2 7 3 0 9 2
4 6 3 2 5
6 0 9 4 13 9 5
72 15 4 3 13 15 1 10 9 7 13 15 9 13 10 0 9 1 3 2 9 9 13 1 10 9 1 10 9 2 3 3 14 13 15 10 0 9 2 7 16 15 4 13 15 13 15 15 4 3 13 15 1 10 9 7 9 2 6 15 4 14 13 2 15 13 1 15 3 13 15 2 6
16 6 3 16 15 9 4 13 0 2 15 4 2 13 15 2 2
25 3 13 10 9 1 10 13 9 9 1 10 9 7 13 16 15 13 1 7 13 7 3 13 15 2
34 16 15 4 14 13 0 7 15 3 13 0 3 15 4 13 10 9 1 10 9 7 13 15 1 10 0 9 2 1 10 9 7 9 2
40 15 4 14 13 10 9 3 2 15 13 15 13 3 0 7 16 3 13 3 15 4 13 1 3 13 10 9 7 14 13 15 3 14 13 0 9 1 15 9 2
13 15 4 13 10 9 9 3 2 0 7 3 0 2
39 15 4 3 3 13 16 10 9 13 1 1 3 12 9 7 3 13 15 2 1 10 9 2 15 4 3 13 10 9 1 10 9 9 7 13 3 3 0 2
24 7 3 3 13 13 10 9 1 9 9 16 15 9 4 13 10 0 9 7 9 1 15 9 2
3 0 9 2
33 3 15 9 3 2 10 9 2 13 15 9 1 13 2 13 4 13 14 13 3 0 1 15 7 0 1 15 9 1 10 0 9 2
12 15 9 2 13 15 16 15 15 13 0 2 5
6 13 14 13 1 11 2
23 15 13 10 12 9 0 0 9 7 15 4 13 1 9 1 9 0 1 10 9 11 9 2
15 11 13 1 11 11 3 15 4 3 13 10 0 9 9 2
3 10 9 2
10 13 0 7 13 1 11 13 3 0 2
13 15 4 13 10 11 11 1 11 11 2 3 9 2
10 15 13 0 1 9 0 2 9 2 2
12 7 2 15 4 13 8 3 15 9 13 15 2
29 1 0 9 2 13 3 3 0 15 13 14 13 10 9 1 10 9 2 15 4 3 13 14 13 1 10 9 9 2
6 7 2 4 15 13 2
15 13 10 0 13 15 10 9 3 15 13 16 13 1 11 2
11 13 15 9 3 2 16 15 4 14 3 2
19 2 13 10 11 13 14 0 2 15 4 14 13 1 3 3 12 9 2 2
1 8
24 10 0 9 9 2 16 15 13 10 0 9 7 10 2 13 2 9 13 1 12 5 12 9 2
27 13 14 13 2 7 13 15 12 9 9 4 13 1 0 9 7 10 9 9 14 13 1 11 2 14 0 2
7 13 15 13 0 1 15 2
12 3 2 13 14 13 1 11 2 13 14 0 2
20 15 4 13 2 14 13 10 9 2 7 13 14 4 13 2 1 10 0 9 2
46 15 9 2 10 0 10 0 2 7 15 0 9 9 2 13 1 10 0 11 7 11 11 9 2 7 10 0 0 9 2 10 9 7 0 0 9 1 10 11 2 4 3 13 1 9 2
31 15 13 10 9 2 7 15 4 4 13 1 9 1 9 1 9 2 1 3 1 10 9 2 1 10 9 1 10 9 9 2
25 16 15 4 14 13 10 9 9 3 5 15 13 3 12 1 12 9 3 16 4 13 1 11 11 2
9 3 4 14 13 15 9 2 3 2
15 10 15 13 2 4 14 13 14 13 3 8 1 0 9 2
35 15 4 14 13 0 14 13 9 7 13 10 9 2 1 11 2 8 16 13 14 13 15 11 11 7 0 11 11 11 9 1 10 0 9 2
21 13 10 11 7 1 10 2 9 2 15 4 4 13 3 3 16 15 13 3 3 2
13 13 15 3 2 7 3 2 7 15 4 13 0 2
2 11 11
2 11 2
6 3 14 13 15 9 2
9 15 13 10 12 9 9 9 9 2
8 3 15 4 13 9 13 15 2
24 15 4 3 3 13 13 1 9 2 10 9 15 13 10 9 1 2 15 4 13 14 13 15 2
11 7 15 4 14 13 15 3 15 4 13 2
15 15 13 9 1 9 1 15 2 7 3 15 4 14 13 2
14 13 15 10 9 4 13 15 13 3 14 13 1 9 2
23 7 10 9 15 13 8 9 15 4 13 1 9 7 13 1 15 2 4 14 13 1 15 2
9 15 13 3 0 1 9 15 13 2
5 3 14 13 15 2
48 0 9 13 10 9 15 13 1 10 9 7 9 0 1 15 2 15 4 13 14 13 3 2 16 15 4 14 2 15 4 13 10 10 9 16 15 13 15 13 3 2 15 4 15 13 1 15 2
5 9 13 10 9 2
5 13 15 3 3 2
11 6 2 15 13 10 9 9 1 12 9 2
12 15 13 14 13 15 4 13 10 9 9 9 2
32 10 9 1 9 13 1 10 9 14 9 7 9 7 13 10 9 1 10 9 3 1 10 9 1 10 9 1 9 1 9 9 2
13 10 9 2 15 4 14 13 10 9 14 13 15 2
30 3 15 13 15 9 14 13 1 15 3 2 13 15 3 2 6 6 2 3 13 15 1 10 0 9 7 13 15 9 2
15 13 15 3 7 3 7 15 4 13 14 13 1 10 9 2
6 9 13 10 9 3 2
16 15 13 10 0 9 7 4 13 1 9 7 9 1 15 9 2
17 7 3 2 3 13 1 9 7 0 9 2 3 13 7 3 13 2
6 3 13 1 1 9 2
16 15 13 15 9 14 13 15 1 15 9 9 2 14 13 15 2
6 0 9 1 15 9 2
4 10 10 0 2
14 13 15 1 9 9 9 7 13 10 0 9 9 2 5
21 3 4 14 15 13 10 9 10 15 13 7 3 13 15 15 3 15 13 9 3 2
21 7 2 16 15 13 1 0 9 1 9 2 13 10 9 9 9 7 9 3 3 2
28 13 14 13 15 14 13 2 10 13 14 13 1 15 16 15 13 14 13 1 10 9 2 7 15 4 13 15 2
33 7 15 4 3 13 10 13 9 1 10 9 7 15 4 13 1 10 9 7 3 2 16 15 13 3 3 2 4 13 1 10 9 2
22 10 9 1 9 4 15 13 14 13 1 11 11 2 11 2 11 1 5 12 1 9 2
3 6 9 2
35 15 4 13 14 13 11 1 10 9 1 10 9 1 11 0 9 7 15 4 13 10 9 1 9 15 4 13 1 5 12 1 9 1 9 2
28 15 4 13 12 1 15 3 15 4 3 4 13 1 12 9 9 1 5 12 2 3 1 10 9 1 10 9 2
40 15 4 13 1 10 13 2 3 9 16 15 13 14 13 10 9 16 13 10 9 10 13 0 2 3 13 1 9 1 10 9 2 7 13 1 10 9 15 13 2
8 9 1 9 16 13 15 9 2
23 6 2 3 13 14 13 2 4 15 13 0 14 13 2 1 1 10 9 3 1 8 13 2
8 1 11 15 4 13 11 11 2
9 13 1 11 3 7 13 3 3 2
7 9 13 1 12 1 9 2
6 10 9 13 3 0 2
16 4 13 2 1 11 15 13 0 14 13 0 9 2 9 9 2
11 15 4 13 10 9 1 10 11 11 9 2
21 15 13 1 10 9 13 1 10 9 2 0 9 9 3 7 10 9 13 3 0 2
19 7 1 0 2 11 13 10 0 9 14 13 10 0 0 9 1 10 9 2
7 1 11 15 4 14 13 2
19 15 4 13 1 10 3 0 9 3 2 7 15 4 13 10 9 7 11 2
18 3 2 16 13 13 9 3 15 4 13 7 16 15 13 10 9 9 2
20 1 11 15 4 13 1 10 9 0 9 13 2 15 13 15 1 10 11 11 2
9 15 13 0 7 0 1 10 11 2
8 15 13 3 0 14 13 9 2
9 2 4 14 13 1 11 3 3 2
6 12 9 13 0 2 2
6 15 13 0 9 3 2
16 15 4 13 12 1 10 0 9 3 7 15 13 0 7 0 2
7 0 9 2 13 15 9 2
33 15 4 13 10 0 9 9 1 5 12 1 9 1 10 9 15 13 2 10 9 3 4 13 15 14 13 0 9 1 11 7 11 2
1 8
15 14 13 1 11 2 11 11 11 13 0 14 13 1 11 2
6 15 13 1 11 11 2
29 10 0 9 1 3 1 11 11 11 11 2 11 11 2 7 11 11 11 7 11 11 7 11 11 13 3 1 15 2
15 14 13 1 11 2 11 11 7 11 11 13 0 1 15 2
5 15 4 3 13 2
11 14 13 1 11 2 11 11 13 15 9 2
10 10 12 1 1 15 13 10 0 9 2
16 10 9 2 10 9 2 10 9 2 10 9 7 10 9 9 2
9 7 3 13 10 12 10 0 9 2
5 13 10 9 9 2
13 15 13 10 9 2 7 9 7 9 13 14 13 2
22 10 9 9 13 0 16 15 13 10 9 0 1 10 9 2 9 2 9 2 7 9 2
23 3 16 15 13 15 2 15 13 0 14 13 2 16 0 9 3 13 14 13 1 15 9 2
7 3 15 9 13 9 9 2
9 2 7 15 4 14 13 3 3 2
13 13 16 15 15 13 1 10 9 2 14 13 0 2
26 3 13 1 10 9 15 13 2 3 0 9 15 4 13 10 9 2 3 0 9 15 4 13 2 8 2
12 15 4 13 9 1 10 1 10 9 1 9 2
9 15 9 4 13 14 13 10 9 2
12 15 13 3 0 2 3 0 2 7 3 0 2
28 15 13 14 2 13 1 10 9 2 3 1 15 9 7 13 14 13 1 15 9 7 13 1 1 15 9 9 2
19 10 0 9 13 15 4 4 13 1 9 7 9 7 13 10 3 0 9 2
13 15 13 9 2 9 2 7 15 13 0 9 9 2
35 15 0 9 4 13 14 13 10 9 9 2 3 3 3 0 1 9 1 9 2 3 3 15 13 14 2 7 3 3 1 0 9 7 9 2
11 3 2 9 7 9 7 3 0 9 9 2
15 15 2 3 2 13 0 9 9 7 4 13 10 10 9 2
15 15 4 13 15 9 2 7 15 13 0 7 13 15 9 2
12 15 4 3 13 10 9 10 4 14 13 15 2
7 3 13 2 13 10 9 2
5 13 10 9 9 2
4 15 13 12 2
9 15 13 0 7 13 14 4 13 2
13 15 13 14 13 12 16 15 4 14 13 3 3 2
7 13 0 15 13 12 9 2
12 12 9 4 13 7 15 3 4 14 13 9 2
21 9 9 2 3 13 9 2 13 0 9 7 13 0 1 10 9 7 13 1 9 2
21 15 4 13 3 15 13 15 1 10 9 16 15 14 13 15 10 9 1 9 9 2
15 15 13 9 7 9 9 7 9 2 9 2 9 2 9 2
25 4 14 13 15 9 2 9 2 9 2 9 2 9 9 2 15 13 3 3 0 16 15 14 13 2
13 3 15 4 14 13 9 2 15 13 0 1 15 2
30 16 15 13 10 9 0 15 4 14 13 7 15 4 13 13 1 9 1 15 2 3 13 15 1 15 9 7 13 15 2
9 13 12 9 0 9 7 13 15 2
3 13 9 2
15 15 13 14 13 7 13 9 2 7 13 14 13 13 9 2
23 15 13 15 0 9 7 15 13 12 12 9 0 9 3 3 7 13 1 15 9 14 9 2
23 15 4 14 13 14 13 14 13 15 1 16 15 13 12 9 0 7 15 4 13 15 9 2
26 15 13 9 3 2 3 3 15 9 2 2 2 7 4 3 13 14 13 3 9 2 13 15 0 9 2
10 15 9 7 9 13 3 0 1 9 2
17 15 13 15 13 0 7 16 9 4 13 2 7 15 13 3 0 2
23 15 9 3 13 0 3 16 15 4 13 1 15 9 9 3 3 3 10 9 1 3 3 2
17 10 9 7 0 9 14 13 15 10 3 0 9 4 4 3 13 2
11 15 13 3 3 10 9 15 13 2 6 2
11 13 15 1 12 9 1 0 14 13 9 2
10 16 15 13 13 9 2 13 10 9 2
13 13 0 15 13 9 1 9 9 10 4 13 3 2
18 13 1 10 9 1 9 2 15 4 3 13 3 0 1 12 1 9 2
18 15 4 13 10 9 1 9 7 3 13 3 10 9 15 4 13 0 2
15 1 10 9 15 13 15 3 14 13 3 14 13 1 9 2
13 3 16 15 13 9 2 13 1 1 15 9 9 2
9 15 4 13 9 7 9 7 9 2
9 15 4 13 1 15 9 7 9 2
19 1 10 9 15 4 2 4 13 13 15 3 14 13 15 9 7 9 3 2
20 7 1 10 9 2 3 13 9 7 0 9 9 15 4 4 13 1 10 9 2
6 3 13 9 1 15 2
18 13 9 1 9 7 13 0 15 13 9 3 14 13 10 9 15 13 2
15 13 13 10 9 10 0 9 10 9 1 0 9 1 9 2
19 13 14 13 1 3 1 10 0 9 1 9 7 13 15 16 15 15 13 2
16 16 15 3 4 14 13 10 9 2 13 10 0 9 13 0 2
25 15 4 13 9 9 1 0 9 1 0 9 2 0 2 13 1 9 2 13 10 0 9 2 8 2
8 15 13 10 9 13 3 0 2
29 3 15 4 14 13 7 13 2 15 4 14 13 3 3 0 9 2 15 4 14 13 3 3 0 9 9 2 8 5
11 13 9 13 14 15 9 7 13 15 1 2
10 7 13 0 9 16 15 13 0 9 5
8 13 10 9 3 1 10 9 2
17 3 13 9 9 1 10 0 9 2 13 9 2 13 10 9 8 2
14 15 13 10 9 14 13 1 10 9 9 9 1 11 2
15 15 13 10 0 9 14 13 1 10 9 9 9 1 11 2
4 13 9 7 9
10 15 13 16 16 15 3 13 10 9 2
32 10 9 13 10 9 3 1 10 9 2 1 10 0 9 2 15 13 14 13 15 9 14 9 1 10 9 9 2 9 14 9 2
11 15 0 12 9 4 13 1 0 11 9 2
9 10 9 9 4 13 3 1 9 2
10 15 0 9 2 4 13 1 0 11 2
35 15 4 14 13 16 15 4 14 13 15 1 10 0 9 1 9 15 4 13 1 1 10 9 7 4 13 14 13 1 9 9 1 12 9 2
22 12 9 3 3 15 13 3 16 13 1 15 9 9 2 15 13 1 15 4 3 13 2
53 15 13 14 13 10 11 1 10 11 11 1 11 11 2 13 9 1 10 0 9 9 13 3 1 15 2 16 15 4 14 13 10 0 9 1 15 3 2 13 15 1 2 13 15 3 2 3 13 1 15 9 9 2
24 16 15 4 3 13 1 10 9 9 1 10 0 9 2 15 13 0 14 13 15 1 10 9 2
21 1 5 12 15 4 3 13 15 13 7 4 13 1 12 9 9 7 15 9 3 2
19 15 13 1 11 3 3 2 10 9 4 13 3 0 1 0 9 2 9 2
25 15 3 13 0 9 2 7 13 10 0 9 1 10 9 4 10 9 13 1 2 15 13 10 9 2
21 9 2 3 13 8 1 10 9 9 7 13 10 10 9 15 13 14 13 15 9 2
24 15 4 3 13 14 13 15 14 13 0 9 2 7 3 13 1 10 9 7 13 15 10 9 2
10 15 4 3 13 15 10 3 2 3 2
9 13 3 16 15 4 13 1 11 2
1 8
9 16 15 4 13 3 2 13 3 2
1 8
2 0 9
20 15 9 4 14 13 1 15 9 9 16 15 13 12 7 13 15 1 9 9 2
16 15 13 10 9 14 13 13 10 9 4 13 1 10 0 9 2
35 15 13 15 3 16 15 4 13 10 9 15 4 13 14 13 9 16 13 1 15 9 9 3 15 4 3 3 13 1 11 7 1 0 9 2
19 3 10 9 4 13 1 11 10 9 4 13 16 10 9 4 13 10 9 2
15 3 3 16 15 4 13 15 4 13 1 15 1 10 9 2
25 10 0 9 13 10 9 10 13 10 9 1 10 11 3 13 16 3 15 4 13 15 4 13 15 2
6 11 11 7 11 9 2
11 3 16 15 4 13 1 1 2 10 2 2
11 15 13 14 13 10 15 13 3 7 3 2
5 13 10 9 13 2
3 2 0 9
4 2 0 0 9
3 2 0 9
8 2 7 3 0 11 15 13 3
8 6 13 10 11 7 11 9 2
14 11 7 11 11 13 12 0 9 9 10 13 0 9 2
12 10 9 9 13 14 13 1 12 7 10 0 2
8 13 15 10 0 9 1 15 2
10 13 10 9 4 13 15 9 10 3 2
22 1 15 9 15 13 1 12 0 9 2 10 11 11 7 10 11 11 11 1 10 11 2
27 9 10 9 13 1 0 9 1 11 2 11 11 2 11 2 11 11 2 10 11 7 11 11 2 11 11 2
18 10 11 3 13 15 0 9 11 11 11 2 11 11 2 7 11 11 2
22 10 11 1 10 11 13 1 15 0 9 11 11 7 11 2 10 0 9 1 11 2 2
30 15 13 0 1 10 9 10 10 1 10 9 13 7 4 14 13 16 15 4 13 10 0 9 16 13 1 10 9 9 2
10 9 10 9 15 13 10 9 1 9 2
16 3 15 13 10 0 9 7 10 9 1 9 3 7 3 3 2
15 15 13 16 10 0 9 1 10 11 1 10 11 13 0 2
11 1 10 11 15 13 10 9 7 9 9 2
24 16 15 13 13 10 9 2 11 11 13 0 1 10 0 9 7 11 13 3 0 1 10 9 2
19 9 9 15 13 10 9 1 10 9 9 1 10 11 7 11 1 10 11 2
17 15 13 16 10 9 13 10 0 0 9 1 10 11 1 10 11 2
15 9 1 9 10 11 7 11 1 10 11 10 13 0 9 2
17 15 4 13 12 9 10 13 3 1 12 1 15 9 1 10 11 2
33 15 13 10 3 0 9 1 10 11 2 7 13 16 10 9 13 10 0 9 7 16 15 4 14 13 10 0 9 16 13 10 9 2
20 9 10 11 1 10 11 7 11 10 13 9 9 9 2 10 0 9 9 13 2
9 15 10 13 9 1 9 7 9 2
13 15 13 10 11 14 9 3 16 12 13 10 9 2
15 16 15 13 9 2 15 4 13 9 10 15 4 3 13 2
12 9 15 13 10 9 1 10 11 7 13 15 2
13 15 4 14 13 10 9 1 10 11 1 10 11 2
12 3 15 4 14 13 3 3 13 10 9 9 2
14 11 11 13 0 2 7 10 0 9 13 11 11 11 2
5 13 1 15 9 8
3 11 11 2
10 11 4 4 13 10 11 1 9 9 2
9 10 9 13 10 0 14 13 1 2
10 15 3 13 14 13 3 15 13 9 2
8 3 1 10 11 4 15 13 2
4 3 1 11 2
6 4 15 3 13 3 2
10 3 3 4 15 13 1 1 10 9 2
9 2 15 13 12 9 1 9 2 2
9 7 3 3 0 9 4 15 13 2
7 3 15 4 13 13 3 6
2 9 5
15 15 13 3 15 13 7 6 2 9 2 6 1 10 9 2
4 13 11 11 2
29 14 10 0 9 14 13 1 1 10 0 9 16 15 4 3 13 3 7 15 4 14 13 3 15 4 4 13 1 2
5 1 10 11 11 2
4 9 1 9 2
22 15 13 12 1 15 2 12 13 1 11 1 11 7 11 1 11 11 7 3 1 3 2
22 15 13 12 0 13 1 1 10 0 9 1 11 3 1 10 9 7 11 1 10 11 2
7 15 4 15 13 14 13 2
14 0 9 1 11 11 2 11 2 11 1 10 11 11 2
17 9 7 11 1 11 7 10 8 11 9 1 11 2 11 2 11 2
8 10 0 9 1 11 2 11 2
12 0 9 1 11 2 11 2 11 11 7 11 2
18 11 11 0 9 1 11 2 11 2 11 11 2 11 11 7 11 11 2
2 11 2
10 3 3 0 1 10 9 1 10 11 2
7 4 15 13 10 0 9 2
9 15 4 13 10 9 1 11 3 2
9 1 11 1 11 1 11 7 11 2
13 11 1 10 9 9 2 11 7 10 3 0 11 2
34 10 9 9 1 11 7 10 11 1 11 1 10 9 9 1 10 11 7 10 9 1 11 16 13 3 1 11 7 11 7 11 7 11 2
30 15 4 13 1 10 1 10 9 7 4 3 13 10 9 1 15 9 13 1 9 2 0 9 13 2 15 9 7 9 2
11 9 1 9 4 13 0 1 3 0 9 2
22 4 15 13 14 13 10 10 9 7 3 10 0 9 7 1 15 9 1 10 0 9 2
15 4 15 9 13 15 16 3 3 15 4 13 1 10 9 2
27 15 13 10 9 1 9 1 9 2 9 2 13 10 9 2 9 2 0 9 2 15 13 15 7 9 13 2
40 16 15 13 10 9 7 10 9 1 10 9 3 15 4 13 0 14 13 1 3 15 4 13 2 1 3 3 15 4 13 7 15 15 4 13 3 15 13 3 2
7 12 9 1 9 7 9 2
3 0 9 2
17 15 13 13 10 0 0 11 7 13 9 1 10 11 15 9 13 2
11 15 4 14 13 10 9 16 15 15 13 2
4 13 1 11 2
6 11 2 10 0 9 2
5 7 3 1 11 2
4 11 9 9 2
6 0 1 10 9 9 2
12 3 4 15 13 15 9 13 1 10 0 9 2
16 15 7 15 9 4 13 1 10 0 9 3 1 10 0 9 2
25 15 4 3 13 10 9 1 10 9 1 10 9 13 1 9 7 10 0 9 13 1 10 0 9 2
16 15 4 13 10 9 1 12 9 7 4 14 13 14 13 15 2
11 3 4 15 13 15 13 1 10 0 9 2
14 15 4 14 3 13 9 2 15 9 4 13 15 9 2
40 9 13 3 0 1 9 2 7 15 13 3 0 3 15 13 1 10 0 9 2 10 0 9 4 13 0 1 9 2 7 0 9 2 6 3 3 15 13 3 2
26 15 4 13 14 13 15 3 10 0 9 14 13 2 16 15 4 13 15 15 9 2 7 13 0 3 2
15 3 2 15 4 13 10 9 14 13 1 3 15 13 0 2
30 15 4 13 14 13 15 9 7 9 2 7 10 9 7 9 13 15 2 7 13 1 9 2 7 13 15 1 10 9 2
34 10 9 15 13 1 13 0 2 13 15 3 0 16 15 4 13 4 13 10 9 16 9 13 0 2 2 7 9 4 13 3 3 3 2
13 13 10 9 2 7 13 15 1 3 1 10 9 2
17 15 4 13 3 0 1 10 12 9 2 1 1 10 0 0 9 2
22 15 4 13 10 9 2 13 9 1 15 9 2 7 13 14 13 15 13 1 15 9 2
40 15 4 13 15 16 10 0 9 13 1 3 2 7 16 10 0 9 4 13 3 2 15 13 0 16 15 13 1 9 0 14 9 3 15 13 1 10 0 9 2
22 1 10 9 14 9 2 15 4 4 13 15 15 2 7 4 4 13 0 0 1 0 2
11 13 15 1 1 10 10 9 2 14 13 2
6 3 13 15 3 3 2
18 15 4 4 13 1 2 3 13 3 1 15 9 4 13 15 3 0 2
31 13 10 9 15 13 3 10 9 2 7 1 10 0 9 2 3 13 15 1 15 9 1 9 2 16 15 13 0 14 13 2
20 3 15 4 13 10 0 9 15 2 7 15 13 10 12 0 9 14 13 1 2
20 13 14 13 1 15 16 15 13 1 10 9 2 7 13 15 3 0 15 13 2
33 13 14 13 15 10 9 15 13 14 13 16 10 9 13 15 2 13 15 2 7 15 4 13 0 1 10 0 9 1 10 0 9 2
10 15 4 3 13 13 1 9 1 9 2
12 0 9 1 15 0 9 7 1 15 0 9 2
19 13 15 13 3 15 13 15 9 13 14 13 10 0 9 16 15 13 0 2
10 1 9 3 15 2 15 4 13 2 5
8 15 3 13 15 1 15 0 2
15 15 3 13 10 12 9 0 9 0 9 1 0 0 9 2
13 0 9 2 15 13 10 12 9 0 0 0 9 2
33 2 15 13 12 9 2 15 4 14 13 1 10 9 2 7 15 0 9 13 16 15 4 14 13 3 1 9 2 7 3 1 15 2
19 15 4 13 3 7 15 4 13 1 10 9 7 13 1 15 7 13 3 2
14 15 0 0 9 13 16 15 4 14 13 1 15 9 2
20 15 4 13 10 9 7 13 14 13 15 1 3 10 9 2 15 4 14 13 2
10 15 4 14 3 13 3 1 10 9 2
11 16 15 13 1 15 2 15 4 13 3 2
12 3 4 15 13 15 14 13 0 1 15 9 2
12 7 14 3 13 3 2 7 14 13 1 9 2
8 15 4 14 13 9 1 9 2
5 15 13 3 0 2
15 15 13 10 12 9 0 0 9 10 15 13 1 10 9 2
5 15 13 15 15 2
58 15 13 9 13 2 9 13 2 7 4 13 2 13 3 2 13 2 13 2 13 2 7 4 3 13 1 10 0 9 16 15 13 10 9 1 10 9 7 3 3 3 1 15 9 2 7 15 4 14 13 15 16 15 13 15 10 9 2
10 6 2 9 1 9 7 9 1 9 2
14 15 3 4 14 13 3 14 13 15 1 10 13 9 2
9 15 13 15 1 16 15 13 9 2
40 2 7 3 2 15 15 13 13 10 0 9 15 13 1 15 9 2 9 1 9 2 9 1 9 2 9 1 9 2 9 1 9 2 7 9 1 9 2 6 2
8 13 15 10 9 15 4 13 2
7 3 13 10 9 1 9 2
10 15 13 14 13 1 9 1 10 9 2
16 15 13 9 14 13 15 0 9 0 1 10 9 7 13 3 2
7 15 4 13 1 10 9 2
16 13 10 9 1 10 9 7 3 13 1 10 9 10 0 9 2
12 3 13 10 9 1 7 13 9 0 1 15 2
5 3 13 15 3 2
26 3 10 9 13 0 1 15 2 3 13 10 9 7 13 1 10 9 2 13 10 9 0 10 10 9 2
5 13 9 0 3 2
13 13 15 9 13 3 3 15 13 14 1 10 9 2
6 4 14 13 10 9 2
11 13 15 13 3 7 3 1 10 0 9 2
23 1 10 9 15 4 13 0 1 15 7 15 4 3 13 10 9 7 14 1 3 3 3 2
13 13 10 9 7 13 15 1 7 13 3 15 13 2
10 16 15 13 15 2 15 4 3 13 2
16 16 13 3 2 13 10 9 1 7 3 13 15 1 10 9 2
8 15 4 13 14 3 13 15 2
8 9 3 4 13 1 10 9 2
4 13 9 9 2
22 13 9 1 15 2 15 3 13 15 7 15 13 3 15 4 13 16 15 13 15 3 2
15 3 4 15 13 10 0 9 1 10 11 11 1 0 9 2
26 4 3 13 1 11 11 11 1 12 9 7 15 4 13 1 10 12 9 7 12 9 9 1 11 11 2
18 15 4 4 13 3 3 7 13 9 13 3 0 7 10 9 13 0 2
9 4 15 3 13 7 13 3 3 2
12 7 13 15 0 16 15 13 16 15 13 3 2
20 16 15 13 2 4 10 9 15 13 3 1 0 9 13 10 0 9 9 9 2
12 3 2 10 9 9 4 13 3 0 3 3 2
3 13 15 2
13 16 15 13 0 7 0 2 13 11 11 2 11 2
18 15 4 13 3 1 12 11 11 11 1 10 9 1 10 9 9 9 2
10 15 4 13 10 9 7 15 13 0 2
18 15 13 10 9 1 10 9 9 10 13 0 7 10 9 9 13 0 2
15 15 4 14 13 10 0 9 7 13 13 3 0 15 13 2
16 3 2 11 11 4 13 3 1 10 0 9 7 13 3 0 2
11 7 6 2 15 4 14 13 1 15 2 5
7 15 13 3 10 0 9 2
10 7 4 14 13 14 13 1 10 9 2
10 10 9 13 14 1 10 0 9 9 2
7 3 0 9 7 9 9 2
7 6 2 16 15 13 0 2
7 11 11 13 14 10 9 2
13 15 13 10 9 9 7 15 13 15 0 9 8 2
3 9 9 12
3 13 9 2
19 15 13 14 0 14 13 1 10 11 2 15 13 10 9 3 10 9 9 2
25 16 15 13 0 15 4 13 10 9 7 9 9 1 15 11 2 16 3 15 13 2 7 11 11 2
18 1 10 1 10 9 2 15 4 13 3 7 13 10 9 1 10 9 2
17 0 1 10 9 10 15 4 13 1 13 9 1 10 11 11 9 2
32 15 13 10 9 1 10 9 2 3 13 10 9 13 2 13 1 10 0 9 2 13 9 7 13 0 9 10 4 13 1 9 2
24 10 9 13 3 0 2 3 16 15 13 10 0 9 2 7 9 2 14 13 14 13 10 9 2
22 9 2 16 15 13 15 1 11 11 11 11 2 13 10 9 1 15 9 11 14 9 2
16 15 4 13 11 11 7 15 13 1 10 9 1 11 11 11 2
34 15 13 10 0 0 14 13 1 1 9 2 15 4 13 10 9 2 7 15 4 13 9 14 9 2 13 15 3 1 10 9 7 0 2
16 15 13 10 9 1 11 11 7 15 4 13 1 9 1 3 2
18 15 4 13 1 10 0 9 1 10 9 1 15 2 7 10 9 9 2
11 13 10 0 9 8 2 3 15 13 1 2
24 15 13 1 11 1 10 9 1 15 11 1 11 11 9 2 7 15 4 13 10 12 9 3 2
46 15 13 10 0 9 7 13 10 9 3 15 13 9 9 2 13 10 0 9 10 4 13 1 10 9 9 2 13 1 13 9 9 7 13 10 0 9 16 15 13 14 13 10 0 9 2
20 11 13 0 16 13 15 3 1 10 3 0 9 7 13 15 9 10 0 9 2
5 9 7 9 2 2
27 15 13 10 9 9 9 1 12 1 15 9 14 9 9 7 15 13 15 13 3 3 0 15 0 9 13 2
14 15 13 15 1 15 9 7 15 13 14 13 13 9 2
10 7 15 13 3 3 0 9 7 9 2
29 10 0 9 7 9 2 15 13 0 14 13 10 9 3 3 16 15 13 1 5 12 2 14 13 3 1 9 9 2
15 15 3 13 10 0 9 13 15 9 7 15 0 9 13 2
14 16 15 4 14 13 16 13 3 5 12 1 10 0 9
11 15 3 13 9 9 10 13 1 15 9 2
61 15 4 13 9 1 9 1 10 9 2 10 12 9 9 15 13 1 11 2 15 13 15 4 13 2 9 1 9 9 9 2 13 1 10 9 2 15 13 16 13 0 9 1 15 9 7 9 9 7 14 3 1 10 9 15 13 15 9 7 9 2
11 3 13 15 15 13 3 7 15 3 13 2
37 3 15 3 13 3 15 13 12 9 7 13 15 3 3 14 13 15 9 1 15 9 7 13 15 3 1 12 9 1 10 9 1 10 0 9 9 2
9 3 10 0 9 1 10 0 9 2
29 3 12 9 1 10 9 1 10 9 16 10 15 9 13 1 3 3 16 15 4 2 16 15 4 14 13 10 9 2
23 3 10 9 13 9 2 12 9 3 3 3 16 15 4 7 10 0 3 2 3 13 9 2
34 15 4 3 13 13 2 3 12 9 2 3 12 1 10 9 2 3 3 12 3 12 13 0 10 9 4 13 1 10 9 1 15 9 2
26 16 10 9 4 13 1 15 9 2 15 13 15 9 3 2 13 10 9 3 1 10 9 1 15 9 2
11 13 10 9 13 9 2 7 10 0 9 2
28 10 10 4 13 15 13 10 9 3 2 13 0 9 7 13 15 9 3 2 14 13 15 9 1 10 0 9 2
20 3 15 4 14 13 15 9 13 1 9 2 15 4 13 1 10 9 10 9 2
13 3 15 3 13 13 15 15 4 13 15 10 9 2
14 3 15 3 13 15 3 7 3 10 9 7 16 13 2
14 3 3 3 13 15 9 0 2 7 15 9 4 13 2
7 15 4 15 13 9 1 2
35 15 4 14 13 1 9 15 4 13 3 1 9 7 13 15 9 2 13 3 2 1 10 9 2 15 13 3 10 9 14 13 1 15 9 2
11 15 13 3 1 15 9 9 2 3 3 2
9 6 15 3 4 14 13 1 10 9
22 3 10 9 9 4 13 2 3 15 9 3 13 1 15 7 15 4 13 16 13 12 2
68 1 15 9 9 2 3 13 13 10 15 9 1 15 9 7 13 1 1 3 15 9 2 13 15 9 1 13 15 1 9 10 3 15 13 3 10 3 15 13 5 13 15 9 9 2 3 13 13 1 10 9 1 15 9 2 1 10 9 1 15 9 2 7 13 14 13 10 9
21 15 4 14 13 14 13 0 1 5 12 7 3 15 13 10 0 9 16 13 9 2
7 15 3 4 14 13 15 2
8 15 14 13 15 9 1 9 2
11 15 9 4 13 0 1 3 12 9 3 2
14 15 4 4 13 9 3 7 15 13 14 13 0 9 2
18 15 13 15 4 13 16 15 13 14 13 9 7 4 14 13 10 9 2
18 15 13 15 1 10 11 11 7 15 13 9 9 7 9 13 3 0 2
6 10 9 7 9 0 2
26 10 9 13 15 13 9 7 13 15 9 1 15 9 2 10 9 1 9 9 1 1 10 13 3 9 2
5 3 15 9 13 2
13 13 15 0 16 9 14 13 1 9 16 13 9 2
6 7 4 10 9 13 2
19 15 4 13 14 13 15 9 7 15 4 14 13 15 2 15 4 15 13 2
22 15 4 14 13 15 14 13 0 7 3 4 15 13 14 13 15 10 0 9 1 9 2
7 2 10 9 4 13 0 2
3 13 15 5
20 15 4 14 13 9 2 9 15 13 15 7 15 3 4 4 13 10 0 9 2
26 15 13 1 9 16 13 15 7 16 15 15 4 13 3 15 4 14 4 13 9 1 10 0 0 9 2
12 15 4 13 15 10 9 7 13 15 15 13 2
6 13 15 1 10 9 2
26 6 3 15 13 1 10 9 7 15 13 15 13 15 0 9 7 13 9 7 3 10 0 1 10 9 2
23 16 15 13 10 9 0 9 15 13 3 14 13 1 13 9 1 3 3 10 9 1 9 2
35 15 13 3 1 9 14 13 1 15 7 15 4 13 12 3 15 4 3 13 3 7 13 15 9 5 9 9 1 10 9 15 4 3 13 2
7 14 13 15 9 1 9 2
20 8 2 15 13 14 0 16 9 14 4 13 2 3 3 14 13 9 1 15 2
24 3 2 16 15 4 4 13 0 9 2 3 10 9 4 13 1 1 9 1 10 9 7 9 2
17 15 4 3 13 11 2 10 9 0 9 2 7 10 9 1 9 2
11 4 15 9 13 9 2 9 2 9 2 2
18 8 2 15 9 4 14 13 15 16 15 4 14 13 15 4 13 0 2
18 8 2 16 15 13 10 9 1 9 2 3 13 15 3 1 15 9 2
12 15 4 13 1 1 9 7 10 9 1 9 2
17 15 4 13 0 0 2 3 16 15 13 14 13 7 13 9 2 2
18 1 3 15 13 1 1 9 9 2 10 4 13 1 9 7 9 9 2
15 7 13 0 2 13 2 7 13 9 3 4 14 13 0 2
6 8 2 13 15 9 2
24 15 4 4 13 10 0 9 1 15 2 13 10 9 1 9 7 3 0 14 13 1 10 9 2
35 15 13 16 15 9 4 13 16 4 13 2 7 13 1 9 9 14 13 15 9 2 13 10 9 9 2 7 14 13 16 15 13 14 13 2
16 15 4 3 13 15 9 1 3 14 13 9 15 13 9 1 2
14 15 4 13 15 9 2 7 13 3 0 1 15 9 2
15 10 9 3 4 13 0 14 13 15 3 16 15 9 4 2
9 15 13 14 13 15 9 10 9 2
8 13 0 9 7 13 9 9 2
3 0 9 2
3 10 9 2
20 15 9 13 15 3 10 9 4 13 10 9 2 15 4 13 10 9 1 9 2
8 4 15 13 10 9 2 9 2
13 15 4 14 13 16 13 9 13 0 1 10 9 2
15 15 4 13 15 9 3 7 13 15 15 13 0 7 14 2
4 0 9 9 2
22 15 4 3 13 14 13 15 10 0 7 15 15 4 13 10 0 1 13 9 1 15 2
11 15 13 1 15 9 7 3 13 1 11 2
24 13 1 10 8 2 0 9 15 9 1 9 13 2 13 10 9 2 13 15 1 2 8 2 2
17 3 2 15 4 13 1 10 9 16 10 0 9 9 13 3 0 2
17 1 15 2 9 4 3 13 13 1 9 7 9 2 3 13 1 2
31 1 9 2 1 15 9 12 2 1 2 12 9 13 9 10 13 3 3 7 3 2 3 2 3 2 1 15 8 2 11 2
11 15 13 3 3 0 16 13 1 10 9 2
19 15 3 2 13 3 1 10 0 2 16 15 4 13 10 0 9 1 9 2
4 13 15 0 2
14 15 4 13 10 0 9 15 13 15 2 7 15 13 2
11 15 13 0 3 15 13 10 0 1 9 2
10 15 13 3 0 3 15 13 3 0 2
19 3 2 3 15 13 1 9 7 3 15 13 9 3 15 13 14 13 15 2
22 15 3 13 14 13 15 3 15 13 15 1 1 10 9 2 1 10 9 15 13 13 2
15 15 9 13 15 13 10 9 1 15 7 3 13 15 3 2
11 7 10 9 15 13 13 14 13 10 0 2
10 4 15 3 13 9 1 10 0 9 2
20 15 15 4 13 1 10 9 13 3 0 7 3 3 15 4 14 13 10 9 2
36 15 13 14 0 1 10 9 2 3 10 2 9 2 7 2 9 2 4 14 13 1 15 3 15 13 16 13 1 10 9 1 9 1 0 9 2
14 16 15 15 13 10 9 13 1 10 9 13 3 0 2
25 15 4 14 13 15 3 16 15 4 3 13 15 7 13 0 0 14 13 15 14 13 13 15 1 2
24 15 4 3 13 0 1 0 16 15 4 14 13 14 13 15 7 15 13 15 1 10 0 9 2
34 15 13 15 13 15 7 15 13 15 1 10 9 7 3 1 10 9 2 7 15 4 14 13 15 13 15 7 13 14 13 1 1 15 2
20 1 9 15 4 14 13 14 4 13 1 10 9 13 1 15 2 10 13 0 2
29 13 10 9 16 15 15 13 2 15 13 10 9 16 15 13 9 1 9 2 7 15 4 14 13 14 13 9 3 2
31 2 8 2 2 13 2 8 2 2 7 2 15 4 13 15 2 7 15 4 13 15 0 1 15 9 9 3 1 9 2 2
7 11 13 15 10 0 9 2
8 15 4 13 1 10 0 9 2
42 15 15 13 14 13 13 16 15 13 0 1 11 14 13 13 9 9 1 9 2 15 13 9 0 16 9 7 9 13 3 9 2 10 13 3 15 10 9 13 1 15 2
45 15 3 13 15 9 0 1 10 9 7 15 13 14 15 9 1 10 9 7 15 4 13 14 13 15 1 10 9 9 2 7 13 14 13 15 13 16 15 4 14 13 14 13 3 2
33 16 15 13 0 3 15 13 0 15 4 13 15 13 16 1 0 9 15 4 13 0 16 9 4 14 13 16 15 4 13 15 9 2
26 15 4 13 10 2 13 10 9 13 1 9 1 15 2 7 13 0 16 15 3 13 10 9 1 9 2
24 0 1 10 9 16 9 4 14 13 10 9 1 9 2 7 15 13 10 9 15 0 9 13 2
8 4 4 13 9 16 15 13 2
12 3 14 3 13 15 9 7 13 15 15 9 2
14 0 7 0 2 13 10 0 11 11 13 13 10 9 2
8 15 13 10 9 1 10 9 2
23 15 4 3 13 14 13 1 15 9 16 15 4 13 1 11 7 13 9 1 10 9 9 2
10 13 15 10 9 1 15 9 14 9 2
4 5 11 11 2
9 15 13 12 9 1 10 0 9 2
22 9 15 13 1 9 13 14 13 1 9 1 3 3 16 0 16 15 13 3 9 0 2
15 9 13 14 13 10 9 7 13 3 2 1 11 2 8 2
18 15 13 3 10 9 1 15 2 9 1 9 2 0 9 2 8 2 2
26 15 9 4 14 13 9 7 13 15 16 15 4 13 14 13 5 12 1 9 1 10 9 15 13 12 2
4 3 2 9 2
3 5 11 2
6 15 3 13 15 9 2
5 15 13 3 0 2
20 15 4 3 13 13 10 9 2 7 15 13 14 10 9 15 4 13 1 1 2
10 15 3 13 15 4 13 1 10 9 2
33 15 4 14 13 15 4 4 13 12 2 7 15 13 10 11 11 9 1 0 9 2 3 15 9 13 3 0 16 15 13 15 13 2
8 3 15 13 3 3 0 3 2
14 15 13 2 15 13 14 0 3 14 13 1 10 9 2
8 7 6 2 15 4 13 0 2
2 6 2
3 5 11 2
12 2 13 2 3 15 4 14 13 10 0 9 2
9 4 15 13 15 13 0 1 9 2
5 3 4 15 13 2
2 13 2
17 15 9 13 3 0 2 7 15 13 14 0 1 0 0 9 9 2
5 10 0 8 0 2
15 1 15 9 2 3 3 0 9 13 1 9 13 0 9 2
23 6 9 1 9 7 9 9 13 0 2 7 3 0 9 13 3 3 1 9 1 10 9 2
24 15 4 13 14 13 10 9 2 3 15 13 16 15 4 3 13 9 3 3 3 15 13 0 2
24 15 4 13 14 13 3 0 7 1 11 2 7 3 3 15 4 13 3 0 15 4 13 0 2
23 15 4 3 13 10 9 14 9 3 15 4 13 3 7 13 0 9 7 13 10 0 9 2
19 15 3 13 16 15 4 14 4 13 3 3 0 1 11 16 15 4 3 2
23 7 15 13 14 3 16 3 0 15 13 2 9 1 9 13 3 0 1 0 9 1 11 2
19 13 13 1 11 1 10 9 14 9 2 3 13 15 1 9 1 11 11 2
14 15 3 13 14 13 1 1 10 10 0 9 1 11 2
17 15 13 3 14 10 0 9 14 13 13 7 13 10 0 9 9 2
14 1 10 9 3 13 10 9 2 7 15 4 3 13 2
14 7 15 4 3 13 9 16 15 15 4 3 13 1 2
21 7 15 4 13 16 13 0 14 13 9 15 4 13 10 9 14 13 13 15 1 2
29 1 10 9 16 15 13 3 15 4 3 13 3 1 11 11 1 10 0 9 1 9 16 15 4 13 15 13 1 2
14 7 10 10 9 15 13 3 15 4 4 13 1 9 2
13 15 4 14 13 3 13 10 9 14 13 1 11 2
23 15 13 15 13 3 0 16 15 13 10 9 10 13 3 12 1 15 9 9 1 15 9 2
11 7 15 13 3 7 15 4 3 13 3 2
24 15 13 3 3 0 0 9 3 3 15 13 16 15 4 13 3 10 9 4 13 1 15 9 2
4 15 12 9 2
4 13 10 9 2
5 15 4 13 3 2
18 16 9 9 13 0 1 10 9 2 4 14 13 15 13 0 1 11 2
27 9 4 4 13 10 9 1 3 10 9 9 1 9 1 10 0 12 5 9 2 3 15 13 14 9 0 2
8 15 13 16 15 15 13 1 2
7 12 9 9 4 14 13 2
10 15 13 13 15 13 2 15 13 9 2
10 3 4 15 0 9 9 13 14 13 2
8 15 13 10 0 0 9 9 2
15 15 4 13 9 15 4 14 13 15 14 13 7 15 13 2
18 15 13 10 0 9 2 1 9 7 9 1 9 9 7 10 9 9 2
20 3 3 16 15 13 2 9 13 3 0 16 15 4 13 3 15 9 13 0 2
12 13 1 10 9 2 15 13 0 7 13 0 2
11 15 4 4 13 1 10 9 16 15 4 2
17 2 15 13 16 9 10 13 9 13 1 10 9 4 14 13 2 2
55 15 4 4 13 9 2 15 13 3 0 15 4 4 13 15 1 1 15 9 2 7 3 15 4 4 13 15 9 7 15 4 14 3 13 15 10 9 1 15 2 15 3 13 15 9 1 10 9 7 15 13 15 1 2 2
7 15 13 15 10 0 9 2
27 15 13 0 2 16 0 9 9 13 2 7 15 13 10 3 0 0 3 2 15 3 13 14 13 7 9 2
7 15 3 13 15 1 9 2
11 15 4 14 13 3 15 4 14 13 3 2
20 15 4 13 13 15 12 7 12 0 9 7 12 7 12 0 2 13 2 9 2
16 15 4 3 13 13 15 10 9 10 13 3 3 16 15 13 2
29 15 4 13 13 15 1 10 0 9 7 13 15 1 10 0 9 1 10 9 7 3 7 15 4 14 13 10 9 2
14 15 13 1 9 1 15 7 4 14 13 14 13 15 2
11 15 4 14 13 14 13 16 15 13 9 2
27 15 4 13 2 13 2 7 9 7 0 9 2 7 13 15 1 14 13 15 9 2 7 15 4 14 13 2
19 15 4 13 13 7 0 7 13 9 1 9 9 2 7 1 0 9 9 2
22 15 4 13 10 0 9 9 9 7 4 13 13 10 9 1 9 1 10 9 14 9 2
8 15 4 14 3 13 14 13 2
15 15 13 3 0 7 0 7 15 4 14 13 15 14 13 2
9 15 4 14 13 1 10 0 9 2
12 15 4 3 13 14 13 15 12 1 10 9 2
14 15 13 3 10 0 9 2 1 10 9 1 10 9 2
6 4 9 3 0 13 2
12 3 15 13 15 3 0 9 4 15 13 15 2
13 16 15 13 15 3 0 15 4 3 14 13 0 2
19 16 15 4 14 13 0 1 15 3 3 15 4 13 15 13 3 14 0 2
16 15 9 13 12 7 3 15 13 0 15 13 10 9 3 3 2
20 15 4 13 15 3 15 13 0 15 13 15 15 13 7 3 4 14 13 15 2
9 13 9 4 13 10 9 16 13 2
31 1 10 9 2 15 4 3 13 3 3 7 13 10 9 2 0 9 13 9 2 10 4 13 1 10 0 9 7 13 9 2
15 9 9 3 13 13 2 3 1 10 0 9 1 10 9 2
8 15 13 10 0 9 14 13 2
27 16 10 9 13 14 0 7 13 2 7 15 9 4 3 13 2 10 9 1 9 3 13 10 9 1 9 2
16 9 13 0 2 7 10 9 1 9 10 4 13 14 4 13 2
14 10 9 10 4 13 10 9 9 14 13 13 13 9 2
20 15 4 13 3 15 9 9 13 0 14 13 2 16 15 9 4 13 0 13 2
9 15 9 4 13 0 13 2 3 2
13 1 10 0 9 10 9 4 13 14 13 15 9 2
25 1 9 2 10 9 4 3 13 1 15 9 1 7 10 9 7 9 2 13 3 1 9 7 9 2
23 15 13 0 7 3 3 16 15 4 14 13 10 0 9 1 15 9 13 9 14 13 1 2
16 15 13 2 10 9 1 10 0 9 4 3 13 1 15 9 2
11 15 13 0 7 0 7 15 9 13 0 2
4 13 15 13 2
11 15 13 3 15 13 0 14 13 10 9 2
13 15 13 3 15 9 7 13 10 9 3 10 9 2
8 4 15 12 9 13 7 13 2
6 3 0 13 3 0 2
2 13 2
22 15 13 10 12 7 10 9 9 0 0 13 9 7 10 0 12 9 0 13 0 9 2
21 10 0 9 15 13 15 3 15 13 10 13 1 10 9 9 7 13 15 1 15 2
65 10 0 9 15 13 15 1 1 10 9 16 15 4 13 10 0 1 2 7 10 9 13 3 1 10 0 12 9 16 13 10 0 7 3 15 3 3 13 7 15 4 4 13 2 13 10 0 1 7 1 10 9 2 13 3 1 10 9 7 13 1 10 0 2 2
36 3 3 15 13 16 15 0 9 4 13 1 15 9 7 3 15 9 7 15 4 13 3 3 7 13 3 3 15 13 1 7 3 15 13 0 2
5 4 15 9 13 2
6 7 4 15 3 13 2
35 15 4 4 2 13 2 1 15 9 7 9 3 16 15 13 16 15 13 7 9 3 15 4 13 16 15 13 10 0 3 3 10 12 9 2
4 10 9 13 2
13 15 4 14 13 10 0 9 1 10 9 3 3 2
21 15 13 14 13 15 1 3 3 10 9 2 7 3 10 9 1 0 9 4 13 2
26 13 10 0 9 15 0 0 9 4 13 15 14 13 0 7 4 13 15 10 9 14 13 1 3 0 2
22 3 3 2 15 9 4 13 1 10 9 2 7 15 13 16 10 1 10 9 13 15 2
16 13 15 1 1 10 9 2 7 13 10 9 0 1 10 9 2
8 3 13 15 1 1 12 9 2
14 13 15 12 10 0 9 2 3 12 2 7 3 3 2
25 15 4 13 12 9 2 10 0 9 4 13 15 9 1 10 9 1 15 9 2 13 15 15 9 2
18 15 4 13 14 13 1 7 13 0 2 15 4 13 15 4 14 3 2
23 15 13 15 4 13 9 0 14 9 2 7 4 14 13 15 2 7 13 8 9 14 13 2
10 15 4 13 0 14 13 16 13 0 2
17 3 3 2 15 9 4 13 0 14 13 16 15 9 4 14 13 2
23 3 10 9 13 2 15 4 13 16 10 9 9 13 15 2 7 15 4 13 0 1 15 2
7 10 9 9 4 4 13 2
38 15 9 4 13 15 14 13 15 1 15 9 2 13 15 9 13 9 7 13 10 9 13 10 9 9 13 3 13 2 14 13 10 9 1 1 15 9 2
5 15 13 14 0 2
27 13 15 9 14 13 1 15 9 2 7 16 15 13 10 0 9 1 2 13 10 9 1 9 1 10 9 2
29 15 4 13 9 0 1 15 9 2 7 15 13 14 4 13 16 15 3 13 15 2 7 13 15 9 1 15 9 2
16 15 4 13 14 13 15 2 7 15 4 13 3 0 1 15 2
10 3 15 13 13 2 15 4 14 13 2
9 16 15 13 2 15 4 14 13 2
22 16 15 13 2 7 12 13 2 15 4 13 15 2 7 15 4 13 10 9 1 15 2
10 9 13 0 2 16 15 13 14 13 2
13 16 15 13 2 13 15 2 7 13 15 9 3 2
18 13 10 9 1 15 9 4 13 15 13 3 0 2 7 15 4 13 2
3 0 9 2
13 10 9 13 3 10 2 13 10 9 3 2 9 2
8 15 13 15 4 13 3 3 2
11 3 15 13 13 15 13 15 4 3 13 2
40 16 15 4 13 3 3 7 6 0 13 2 14 13 3 3 16 15 4 2 2 7 0 13 2 14 13 3 3 16 15 4 1 15 9 2 3 15 4 13 2
27 15 13 12 9 2 7 3 3 15 13 1 10 0 16 9 13 3 0 2 7 3 15 4 13 7 13 2
23 10 9 13 3 10 9 13 2 15 13 15 13 0 7 15 13 10 0 9 14 13 3 2
6 15 13 15 4 13 2
20 3 15 4 3 13 1 10 0 7 15 9 4 13 15 13 16 15 4 13 2
10 15 4 13 3 15 13 0 3 2 5
12 15 13 10 9 1 11 11 1 10 11 11 2
28 3 11 13 9 1 12 15 4 13 1 10 0 15 4 13 10 9 2 12 9 3 12 9 14 13 11 11 2
27 15 13 14 13 15 7 13 10 9 14 13 10 9 1 12 1 12 9 2 1 10 0 9 1 12 2 2
12 15 4 14 13 15 10 9 1 9 15 13 2
38 15 13 11 1 0 9 2 3 15 13 10 13 7 13 9 3 1 10 13 7 13 9 10 13 2 1 10 0 9 2 10 0 9 16 13 10 9 2
6 9 13 2 15 13 2
42 10 11 4 14 13 10 0 9 1 10 0 11 2 10 9 9 2 2 15 4 4 13 1 10 0 9 11 2 10 13 0 9 2 7 10 11 11 11 2 11 2 2
46 3 10 11 13 3 1 15 13 7 13 9 10 11 3 13 15 4 14 13 1 1 10 11 9 2 7 10 0 9 4 13 14 13 10 9 7 13 0 1 10 9 1 11 7 11 2
18 10 10 0 9 1 10 9 1 11 13 0 2 10 11 4 4 13 2
18 3 2 11 4 14 13 10 9 13 10 9 7 13 1 10 11 9 2
25 15 4 13 16 15 4 13 1 10 0 9 7 4 3 13 10 9 2 7 15 13 15 0 9 2
4 10 11 13 2
7 15 4 14 13 10 11 2
36 3 2 15 15 13 14 13 1 10 11 11 13 14 13 1 10 11 7 13 10 11 1 10 0 9 3 15 4 13 13 0 13 7 13 9 2
40 10 11 13 15 4 13 10 11 2 13 10 9 1 10 0 0 9 2 7 10 9 4 3 13 1 10 0 9 7 13 10 11 13 1 10 9 1 0 9 2
5 10 13 10 9 2
3 15 13 2
20 10 11 13 10 9 14 13 10 0 9 7 4 3 13 9 1 10 0 9 2
10 10 11 13 3 1 9 9 7 13 2
17 1 12 9 10 11 9 4 4 13 1 1 10 0 9 1 11 2
6 10 9 4 14 13 2
6 7 10 0 0 9 2
9 3 13 10 0 9 2 15 13 2
6 1 10 0 0 9 2
12 11 13 10 0 0 7 0 9 1 10 11 2
15 15 4 13 3 1 11 7 11 16 10 11 1 0 9 2
43 10 9 13 15 9 14 13 10 9 2 7 1 10 9 7 9 10 11 9 2 7 10 11 2 13 11 10 9 15 4 13 15 14 13 1 10 9 2 9 15 13 15 2
27 10 15 13 14 13 1 10 0 9 13 13 10 9 14 13 1 11 7 11 7 13 1 10 0 11 9 2
24 7 11 13 3 0 15 4 14 13 15 13 10 9 3 15 4 13 1 15 1 10 0 9 2
36 3 15 13 10 0 1 2 13 10 9 1 11 11 2 13 1 10 0 9 2 7 13 10 9 1 15 9 1 9 13 14 13 1 11 11 2
13 15 13 1 16 3 13 15 9 3 15 13 15 2
33 10 0 9 4 14 13 10 1 15 2 7 13 11 11 14 13 10 9 11 4 13 2 14 14 13 16 10 0 9 4 13 2 2
15 1 10 9 11 13 15 9 1 2 2 9 1 9 2 2
6 7 15 13 10 9 2
12 14 13 10 9 2 7 15 13 10 0 9 2
10 14 13 10 9 0 1 10 0 9 2
8 1 15 2 15 3 3 13 2
33 1 11 2 10 9 13 0 7 0 1 10 9 1 11 16 16 10 9 1 0 9 4 13 1 10 9 16 13 10 11 7 11 2
39 11 13 15 0 16 10 9 13 10 0 9 16 13 3 16 10 11 13 15 4 13 10 11 7 16 10 11 13 3 0 14 13 0 9 14 13 15 9 2
18 15 13 10 3 0 9 1 10 9 10 4 13 1 11 11 11 11 2
14 13 9 14 13 10 9 16 15 4 13 14 13 15 2
5 0 9 9 2 2
8 15 3 13 10 9 12 9 2
36 15 13 10 9 9 9 10 13 15 13 10 0 9 10 13 12 5 0 0 2 9 7 13 0 9 9 0 1 10 0 0 2 9 1 15 2
23 15 9 13 4 15 13 15 13 15 3 3 10 9 2 7 10 2 9 9 2 15 13 2
12 15 3 4 13 3 3 4 10 9 13 3 2
22 10 9 1 11 11 13 12 9 2 7 1 9 1 10 9 15 13 12 1 12 9 2
15 15 4 13 0 1 15 0 9 2 7 4 14 13 3 2
12 15 13 0 9 9 9 7 13 2 13 9 2
7 10 9 4 4 3 13 2
6 13 15 1 15 9 2
41 13 15 13 14 13 15 1 3 3 16 15 4 2 0 2 0 1 10 9 9 2 9 1 10 0 9 13 12 9 1 2 9 2 2 9 2 9 2 7 9 2
23 10 9 9 13 9 9 4 13 9 2 13 9 9 2 15 13 10 0 9 14 13 1 2
14 9 1 10 0 9 4 3 4 13 1 10 0 9 2
40 9 4 3 13 10 0 9 1 10 9 9 2 16 15 13 10 9 2 9 9 9 2 10 13 10 0 9 9 9 10 4 13 7 9 7 9 1 12 9 2
40 15 3 13 16 15 4 14 13 0 2 0 9 9 16 15 4 13 14 13 0 9 9 7 2 7 9 1 9 3 14 13 15 13 9 13 9 9 1 9 2
43 10 0 9 9 9 13 0 2 1 11 14 11 9 2 8 13 14 13 9 9 13 1 10 9 14 9 1 10 9 10 9 4 3 3 13 9 3 16 0 9 3 13 2
36 3 2 14 13 15 9 2 6 2 16 15 3 13 10 9 10 13 15 13 11 3 15 4 14 13 2 10 9 14 9 2 10 15 13 13 2
11 15 13 14 3 13 10 9 1 11 9 2
42 10 9 1 11 13 3 0 2 1 9 15 13 3 10 0 9 14 3 13 15 0 9 9 9 13 15 2 15 4 14 13 10 0 9 9 13 13 0 9 9 9 2
31 11 7 13 9 2 4 13 3 12 11 1 10 9 2 12 11 1 10 9 2 4 13 0 1 12 5 12 9 10 9 2
19 13 13 9 13 14 10 0 9 9 9 2 15 13 14 13 0 9 9 2
25 0 9 13 0 9 2 15 13 14 13 10 9 13 14 13 10 13 9 2 3 3 15 13 9 2
12 11 9 13 3 0 1 0 9 1 0 0 2
34 9 2 9 9 2 0 9 2 7 0 9 9 2 1 13 2 9 2 9 2 7 9 2 13 0 9 1 9 9 14 13 15 13 2
18 11 9 7 0 9 4 3 4 13 1 0 9 2 1 9 14 9 2
22 15 4 3 13 16 15 13 1 10 0 13 9 14 13 0 15 13 9 13 1 3 2
1 8
1 8
26 6 15 13 1 10 9 1 15 9 7 9 7 10 15 13 15 1 2 3 3 3 16 15 13 0 2
74 16 15 13 0 9 15 4 13 1 2 1 9 10 12 5 12 5 12 9 1 9 1 12 9 2 3 15 4 13 15 0 10 0 12 5 12 9 2 16 15 13 10 0 9 7 15 4 14 13 10 9 3 12 5 12 3 3 1 10 9 1 3 3 12 5 12 9 1 10 9 3 10 9 2
40 10 9 15 3 13 14 13 10 9 1 10 9 16 15 4 13 10 9 9 9 1 11 9 1 15 9 1 10 9 3 7 1 0 9 15 4 13 10 0 2
24 1 16 15 10 9 13 15 13 11 13 2 10 13 0 1 9 1 9 16 15 13 1 9 2
17 10 9 1 11 13 10 9 1 10 9 1 15 11 13 2 6 2
18 6 2 15 13 15 10 2 9 9 2 0 2 15 13 15 11 13 2
27 7 15 4 13 3 12 5 12 9 2 3 16 10 9 4 13 3 1 12 5 12 9 1 15 0 9 2
13 1 1 10 9 2 3 13 0 14 13 10 9 2
35 3 2 11 3 4 14 13 9 10 4 14 13 2 3 15 13 9 14 9 16 7 3 15 4 13 10 13 2 13 9 7 10 13 9 2
17 15 13 3 15 9 15 4 13 15 2 7 4 14 13 1 15 2
11 3 13 0 9 9 2 1 9 7 9 2
4 0 1 9 2
8 13 10 9 7 10 9 0 2
67 15 4 13 10 11 9 1 15 9 7 15 4 13 14 13 1 10 9 7 15 13 10 0 9 10 15 13 2 7 15 4 13 2 10 4 14 13 3 2 7 10 13 0 9 14 13 1 9 7 15 13 14 13 10 4 13 0 15 3 4 14 13 7 15 9 13 2
4 6 13 15 2
10 6 7 6 13 3 12 13 0 9 2
3 6 3 2
5 6 13 10 9 2
5 3 13 15 9 2
11 15 13 10 0 9 10 15 13 1 11 2
12 15 13 1 13 10 9 1 9 9 1 11 2
9 1 3 15 13 3 0 7 10 2
10 15 4 13 7 13 15 8 0 9 2
11 1 10 9 1 9 15 13 0 1 15 2
13 15 13 3 0 7 15 4 14 13 7 13 15 2
14 15 4 13 14 13 15 7 15 3 4 14 4 13 2
10 15 4 14 13 14 4 13 7 13 2
12 15 13 10 9 10 15 4 13 7 13 9 2
10 15 3 13 15 7 15 4 13 3 2
11 10 9 1 9 16 15 13 9 2 9 2
10 15 13 0 15 13 0 9 7 9 2
4 15 13 15 2
8 3 1 10 15 13 3 0 2
7 15 13 15 1 12 9 2
10 15 4 13 9 7 15 13 14 0 2
6 10 0 9 13 15 2
7 15 9 3 13 1 15 2
9 15 13 10 0 9 1 15 9 2
9 15 13 15 13 15 1 15 9 2
9 15 13 3 3 10 0 9 9 2
10 3 13 10 9 13 1 10 0 9 2
58 2 10 0 10 0 14 13 2 13 1 0 0 9 2 9 2 7 0 9 9 2 10 9 1 10 9 2 0 9 9 13 10 9 13 14 0 2 13 1 10 0 9 1 10 9 2 10 0 9 13 10 9 9 1 15 9 2 2
24 13 1 10 9 1 9 1 15 9 10 13 1 10 9 7 13 3 1 10 9 1 10 9 2
11 10 9 13 1 9 10 0 9 10 0 2
13 2 13 1 10 13 9 6 2 13 1 0 9 2
19 16 15 13 10 9 10 9 2 10 9 9 1 10 9 2 4 13 0 2
8 10 9 13 7 0 7 0 2
9 15 4 13 16 15 13 12 9 2
13 7 13 7 12 9 7 12 9 2 7 12 9 2
6 4 14 13 12 9 2
28 15 3 4 14 13 3 2 15 13 3 10 9 13 6 6 7 1 0 3 2 12 9 13 14 13 10 9 2
12 15 13 12 0 9 7 10 0 7 0 9 2
5 15 13 10 0 2
18 16 15 13 14 13 10 9 15 13 10 9 10 15 13 14 13 15 2
21 3 16 15 13 16 13 12 2 3 13 0 1 12 1 10 0 9 15 13 9 2
17 15 9 13 15 3 14 13 15 7 15 13 3 0 1 10 9 2
23 15 13 15 12 9 14 13 10 0 9 14 13 0 14 13 1 7 13 1 1 15 9 2
7 15 13 10 9 15 13 2
11 3 15 4 13 1 15 3 1 15 9 2
7 3 15 4 13 1 15 2
18 8 2 3 15 13 10 9 2 13 15 7 15 7 15 1 10 9 2
15 13 15 1 3 1 9 7 9 7 0 1 3 12 9 2
10 8 2 3 13 15 9 1 10 9 2
12 15 13 10 9 7 13 15 3 1 10 9 2
19 3 15 13 1 10 9 2 13 12 9 1 10 9 2 13 10 9 9 2
26 2 10 9 15 4 13 15 9 1 9 2 7 9 13 9 6 2 3 15 13 1 10 9 7 13 2
22 10 9 15 4 13 16 15 9 13 0 7 15 4 14 13 14 13 15 7 13 15 2
7 13 15 1 3 12 9 2
19 2 15 4 13 9 16 15 13 14 2 7 13 10 9 1 3 12 9 2
19 8 2 1 3 9 12 2 15 4 13 1 13 10 9 9 1 15 9 2
26 2 4 14 13 1 10 9 9 1 10 9 2 15 4 13 15 1 10 9 15 13 1 15 9 2 2
20 3 13 15 9 7 13 15 1 15 9 2 1 9 1 15 9 7 13 3 2
11 13 15 9 1 15 9 3 7 13 3 2
43 2 10 0 9 1 9 15 4 13 3 1 10 9 7 3 3 16 15 4 14 13 3 7 13 15 4 13 0 1 15 2 15 4 13 10 9 16 14 13 1 15 9 2
22 3 15 13 16 15 4 14 13 15 2 15 4 13 1 1 15 9 3 15 13 3 2
20 8 2 16 15 4 14 13 3 1 3 15 3 13 14 13 13 7 13 13 2
10 4 14 13 2 13 2 7 13 15 2
4 15 13 9 2
5 4 14 13 1 2
50 1 10 9 1 9 15 13 3 15 13 9 15 13 14 13 1 15 9 2 3 15 13 3 15 13 14 13 3 1 15 9 2 3 15 13 3 7 3 15 13 1 1 15 9 7 1 1 10 9 2
14 7 3 15 13 13 3 15 13 14 13 1 10 9 2
3 0 9 2
12 15 13 1 15 7 15 13 15 13 1 15 2
4 15 13 0 2
15 7 15 13 15 9 3 15 4 13 10 9 1 10 9 2
4 10 9 13 0
2 9 2
14 15 13 3 0 7 15 13 0 14 13 9 1 15 2
5 15 13 3 0 2
8 15 13 10 9 13 11 2 5
10 3 13 10 0 9 14 13 1 11 2
11 15 9 7 15 4 13 14 13 1 11 2
18 15 13 1 10 9 2 7 3 15 4 13 14 13 1 3 7 9 2
30 15 4 14 13 3 0 9 2 7 16 15 4 3 13 1 1 9 15 4 13 3 1 10 9 1 11 1 0 11 2
50 15 4 14 13 15 14 13 3 0 2 14 0 3 3 15 9 13 2 7 15 10 9 13 3 1 3 1 15 9 9 2 2 7 15 4 14 13 16 15 13 14 13 3 1 10 9 1 9 3 2
30 15 13 3 1 15 0 9 7 3 13 14 13 10 0 9 16 15 13 3 0 7 16 15 9 13 14 13 3 0 2
20 4 9 13 15 10 9 16 3 10 0 9 16 15 14 13 1 11 4 13 2
16 9 4 14 13 1 11 1 9 1 10 9 2 15 13 0 2
19 12 9 15 4 13 0 1 1 0 9 13 3 0 15 4 13 0 1 2
20 15 4 13 9 7 9 1 11 2 7 9 9 1 11 7 3 1 10 9 2
7 7 3 3 13 10 9 2
22 11 13 10 9 1 9 2 16 0 9 13 10 9 3 0 1 12 9 1 10 9 2
7 11 11 13 10 3 13 2
12 10 9 13 10 0 2 13 10 3 0 9 2
36 10 0 9 13 1 10 2 12 9 1 10 9 2 9 2 10 8 3 13 16 15 4 14 13 10 9 3 15 13 1 10 9 1 10 9 2
10 10 0 9 2 3 2 4 4 13 2
39 1 9 2 1 11 1 11 2 10 9 13 3 0 7 2 3 3 2 3 0 2 1 10 9 1 9 15 4 14 13 14 13 1 9 1 1 12 9 2
33 15 13 3 0 9 9 2 10 13 15 13 3 0 9 3 3 3 1 10 3 0 9 1 10 9 2 7 9 13 1 15 0 2
26 14 3 2 0 1 10 0 9 13 1 10 9 16 16 14 13 9 1 10 9 7 10 3 0 9 2
43 9 2 11 1 11 2 7 11 2 11 1 11 2 13 0 9 2 16 10 9 14 3 2 13 9 1 10 9 9 4 3 13 10 9 1 8 2 7 0 2 9 9 2
39 3 2 15 13 10 0 9 1 10 9 7 9 2 7 10 9 4 13 3 0 1 11 7 11 1 1 11 2 3 2 15 13 3 9 1 10 9 9 2
12 11 9 13 10 3 2 0 11 11 14 11 2
33 16 9 4 14 3 13 1 9 2 9 2 11 1 11 2 4 13 0 2 1 0 9 1 10 9 2 10 9 7 9 1 0 2
74 9 13 1 15 0 2 7 0 1 10 9 14 9 9 7 9 13 1 1 11 7 4 14 13 1 11 2 10 3 13 9 1 10 3 0 9 16 3 11 4 13 1 0 1 10 0 2 15 13 0 2 0 7 0 1 12 9 2 7 15 13 3 10 9 14 13 1 3 10 9 13 13 3 2
32 10 9 14 13 13 14 13 10 0 9 1 15 2 9 16 15 4 13 1 16 15 13 0 7 13 1 9 3 15 13 1 2
10 0 9 7 9 13 0 7 10 9 2
21 16 10 0 11 11 11 13 2 15 13 10 0 9 1 0 9 3 10 0 9 2
43 0 15 4 14 13 3 0 2 15 13 3 10 9 1 9 9 2 16 16 10 9 13 3 0 3 10 0 0 9 4 13 1 10 0 0 0 9 7 9 7 3 3 2
13 16 15 13 10 11 1 11 2 11 2 3 3 2
22 10 9 3 13 3 3 0 1 0 1 10 11 2 4 15 13 1 10 11 2 2 2
19 15 9 13 10 0 1 10 10 9 1 10 0 9 7 15 4 13 9 2
16 15 4 13 3 0 1 11 3 13 1 9 13 15 0 9 2
4 11 1 9 2
24 13 10 9 7 13 10 9 9 3 1 11 13 10 9 7 15 4 13 10 9 1 10 9 2
45 14 13 10 0 9 15 4 13 14 13 0 3 14 13 10 9 16 0 9 13 0 7 3 13 3 3 1 10 0 9 2 9 2 0 0 9 4 14 13 10 9 7 9 9 2
30 15 4 13 1 10 9 7 13 10 9 9 1 6 10 11 1 11 7 11 11 7 15 4 13 1 10 10 0 9 2
25 1 9 0 9 4 13 1 10 0 9 3 15 4 13 14 13 1 1 10 0 9 1 10 9 2
41 0 9 10 0 9 1 9 4 13 1 0 11 5 0 11 7 15 4 13 1 9 1 9 1 9 1 10 9 1 10 9 3 13 0 1 0 9 2 9 8 2
25 15 3 13 10 0 0 9 10 9 2 3 12 11 1 10 0 9 2 3 1 12 11 0 9 2
9 15 13 15 9 1 3 12 9 2
20 11 13 1 8 11 3 3 3 16 10 9 13 16 14 3 13 1 10 9 2
15 10 9 13 14 13 7 15 13 3 0 2 0 7 0 2
26 15 13 9 1 11 3 15 4 14 13 13 3 1 10 9 14 13 0 2 9 9 13 15 0 9 2
11 15 4 13 15 13 3 0 14 13 11 2
23 15 4 13 14 13 10 0 12 9 13 1 1 9 2 9 2 9 2 9 7 9 9 2
13 13 3 1 0 13 3 0 13 1 11 15 13 2
6 9 9 9 9 9 2
7 15 13 12 9 9 9 2
13 12 1 15 13 3 0 7 13 3 12 9 0 2
15 12 1 15 13 3 0 7 13 3 12 5 12 9 0 2
14 10 0 9 13 0 3 7 15 13 3 12 9 0 2
11 15 13 15 9 2 7 0 9 0 3 2
17 4 15 13 15 10 0 9 16 13 15 7 13 9 1 10 9 2
4 9 1 9 2
2 6 2
14 16 15 13 0 14 13 9 0 2 15 13 3 0 2
17 15 13 1 15 9 9 2 9 3 7 9 0 3 1 10 9 2
20 9 2 7 9 2 13 3 0 1 9 2 9 0 16 13 9 7 13 9 2
15 15 13 16 15 13 16 15 0 7 0 0 9 13 9 2
22 16 15 4 13 0 16 13 1 11 11 13 10 9 1 10 9 1 10 0 9 3 2
8 16 15 13 9 1 15 9 2
6 15 9 4 3 13 2
25 16 9 13 0 2 12 2 12 9 2 7 10 9 13 3 3 13 16 15 13 2 15 4 13 2
16 2 15 4 3 13 10 9 1 9 13 9 1 10 13 9 2
12 16 15 13 14 13 9 13 10 0 9 9 2
6 13 1 10 0 9 2
22 15 13 0 9 16 15 4 13 15 9 2 3 3 7 10 9 13 0 3 1 15 2
24 13 10 3 13 9 9 2 10 9 2 0 9 9 7 3 10 9 1 0 9 14 13 15 2
56 15 13 10 9 9 15 4 13 9 2 9 13 7 9 13 15 1 12 9 2 13 9 1 10 9 7 13 15 1 10 9 1 0 2 0 9 7 13 1 10 9 1 10 13 9 7 13 15 16 10 9 4 13 3 3 2
51 16 15 13 10 9 14 13 10 9 2 8 2 7 9 2 8 2 2 7 13 15 3 1 0 9 2 2 13 16 15 4 13 0 12 5 9 9 2 3 15 13 15 3 15 4 13 10 9 0 9 2
23 3 13 1 9 2 7 16 10 9 13 3 3 2 15 4 13 12 5 12 9 10 9 2
29 1 0 9 7 3 13 2 13 2 13 2 13 9 3 1 10 9 2 15 4 13 12 5 12 9 1 10 9 2
12 13 7 13 3 0 9 2 15 4 13 0 2
32 13 10 9 10 9 1 10 9 2 9 4 3 13 7 13 7 3 13 1 9 2 4 13 15 14 13 7 13 15 0 9 2
14 15 3 13 10 9 1 10 9 7 9 1 15 9 2
8 10 9 9 13 1 15 3 2
10 15 3 4 13 14 13 10 9 9 2
14 10 9 7 9 2 9 2 13 14 0 1 10 9 2
29 3 3 15 13 0 14 13 10 3 13 9 1 0 9 9 1 10 9 14 13 0 9 10 13 3 1 10 9 2
24 3 13 10 9 1 9 13 10 9 1 9 3 1 10 9 9 7 13 0 14 2 13 2 2
30 13 10 9 1 10 9 0 9 1 15 4 13 10 9 14 9 1 9 7 15 13 3 0 14 13 9 7 9 0 2
12 16 10 9 4 14 13 9 2 13 10 13 2
23 8 2 4 10 9 9 2 0 1 10 0 9 7 10 9 7 0 9 2 13 10 9 2
11 8 2 4 15 13 1 1 0 9 9 2
11 8 2 13 15 3 0 9 1 10 9 2
10 9 9 13 0 2 13 1 0 11 2
10 15 13 16 15 13 1 0 9 9 2
28 3 16 15 4 13 15 9 9 14 13 10 9 7 9 2 0 13 9 2 9 2 15 4 13 15 10 9 2
30 13 15 10 0 3 2 10 9 1 12 1 3 12 9 2 9 1 9 2 7 12 1 12 9 4 13 0 1 9 2
26 9 9 2 10 0 9 14 9 9 4 4 13 16 15 4 13 12 1 15 0 9 9 14 0 9 2
29 15 13 10 9 1 9 3 7 15 4 13 1 10 9 1 15 4 13 15 9 9 2 9 2 9 7 9 2 2
10 10 9 1 9 13 14 1 0 9 2
40 3 16 15 13 10 0 9 1 9 9 2 0 9 2 15 4 13 1 10 9 2 9 2 1 10 9 7 13 9 14 13 3 7 13 10 9 7 9 2 2
27 3 3 15 13 0 1 3 13 9 1 0 9 9 1 10 9 14 13 0 9 10 13 3 1 10 9 2
24 3 13 10 9 1 9 13 10 9 1 9 3 1 10 9 9 7 13 0 14 2 13 2 2
16 16 15 13 9 1 10 9 1 10 9 9 2 15 13 0 2
19 7 13 10 9 1 2 3 13 1 0 9 9 7 3 1 10 9 9 2
11 1 9 10 9 4 13 1 10 9 9 2
54 16 10 9 1 9 13 13 1 2 9 9 2 1 13 9 2 10 1 10 3 0 9 9 13 13 16 1 12 5 12 9 1 9 2 15 4 13 10 12 5 9 9 2 16 10 9 13 2 15 4 13 9 9 2
21 10 9 13 16 3 0 9 4 13 7 10 9 4 13 3 7 13 10 10 9 2
28 10 9 13 1 10 3 0 11 9 14 13 1 10 9 2 16 15 4 13 0 9 1 1 10 9 7 9 2
9 9 4 13 10 9 1 11 0 2
20 16 10 9 13 0 2 15 4 13 7 3 13 0 16 10 0 9 13 1 2
6 13 15 3 3 3 2
10 13 15 13 0 9 1 10 9 3 2
7 11 9 9 1 0 9 2
11 15 4 4 13 15 12 7 12 9 9 2
8 15 13 10 0 9 1 9 2
6 4 15 13 10 9 2
11 10 9 7 9 14 13 15 10 0 9 2
2 9 2
5 15 13 9 9 2
10 0 9 13 0 14 13 10 0 9 2
11 15 13 1 9 13 2 0 7 0 9 2
16 15 4 13 0 9 2 15 4 13 0 9 13 1 15 9 2
6 15 13 10 0 9 2
21 3 16 15 4 13 14 13 9 9 1 9 7 9 2 10 0 9 15 4 13 2
10 11 9 2 13 10 0 9 1 15 2
21 15 13 0 9 14 13 11 9 13 10 0 9 16 15 14 13 10 0 9 9 2
20 1 12 3 2 1 15 9 11 9 4 13 0 7 13 14 13 0 7 0 2
18 15 13 10 0 9 2 10 3 0 9 1 9 14 13 15 9 9 2
12 10 9 4 13 3 2 1 0 0 9 9 2
16 4 15 13 16 10 9 1 10 0 9 4 13 3 0 9 2
22 6 2 10 0 9 7 9 13 9 1 10 11 9 13 3 0 1 9 1 10 9 2
26 15 13 10 9 2 15 4 13 10 9 1 9 1 9 14 13 1 15 0 9 2 1 2 9 9 2
13 9 0 9 7 9 9 4 13 1 10 0 9 2
11 15 13 12 9 2 11 11 7 11 11 2
12 10 4 13 13 1 9 10 9 1 10 9 2
22 11 9 13 12 2 9 9 9 2 7 10 9 13 0 14 13 15 10 9 15 13 2
12 15 4 13 3 0 9 2 13 3 7 3 2
7 15 4 13 3 7 3 2
10 10 9 13 9 1 9 2 3 13 2
15 9 9 2 9 7 0 0 9 13 3 1 0 9 3 2
14 15 13 0 0 9 1 0 9 1 10 9 3 3 2
12 15 13 0 9 3 7 3 13 1 10 9 2
11 15 4 13 0 9 13 10 11 11 9 2
9 10 9 9 13 10 9 1 9 2
13 9 9 2 9 9 2 0 9 7 0 0 9 2
9 15 13 3 10 9 1 10 9 2
16 10 0 9 1 9 7 9 4 13 10 0 9 1 10 9 2
6 15 13 0 9 3 2
28 15 13 9 1 9 7 9 2 9 9 2 9 9 1 10 0 2 3 13 0 9 3 7 0 0 0 9 2
16 3 15 4 13 15 9 1 10 9 7 13 10 9 1 9 2
12 14 13 7 14 13 11 9 13 10 0 9 2
13 15 13 0 0 9 13 10 9 9 1 0 9 2
18 15 4 13 10 0 9 7 9 9 16 13 10 9 0 1 10 9 2
16 0 9 13 0 2 3 2 10 11 9 13 3 3 3 13 2
15 15 4 13 10 0 9 2 7 3 9 9 7 0 9 2
13 15 4 3 13 14 13 11 9 7 10 11 9 2
33 15 3 13 15 9 2 9 1 10 9 2 9 1 9 2 13 3 3 13 7 13 9 2 3 2 15 13 10 10 9 3 0 2
19 1 0 9 2 15 4 3 13 10 9 7 9 9 16 15 4 13 3 2
13 13 1 10 9 14 9 3 3 16 15 13 3 2
9 4 14 13 0 16 13 15 3 2
18 15 13 10 9 3 10 3 15 13 3 2 10 3 15 4 13 9 2
37 15 13 13 10 0 9 9 2 16 15 13 0 9 14 13 9 7 9 7 16 15 9 13 2 3 1 9 2 15 4 13 10 0 9 1 9 2
13 13 10 9 1 9 7 0 0 9 1 15 9 2
26 10 1 10 9 13 14 13 0 7 13 2 9 2 1 15 9 13 15 7 15 9 13 15 9 3 2
23 15 4 3 13 9 1 10 9 1 15 9 2 9 2 16 3 15 13 1 10 13 9 2
28 9 9 4 14 13 1 9 7 15 13 15 10 2 9 2 9 2 9 1 9 1 15 9 10 4 13 3 2
23 10 9 15 4 13 10 2 9 2 13 10 11 10 13 10 1 10 9 1 10 0 9 2
31 15 3 13 15 1 9 7 13 10 9 15 13 15 2 13 2 14 13 7 10 13 15 13 16 13 1 9 16 3 13 2
6 10 9 4 13 0 2
19 0 9 9 4 3 13 0 1 9 16 9 4 13 0 1 10 0 9 2
28 15 9 7 15 2 1 15 9 1 10 9 2 3 13 10 12 9 9 7 10 9 9 13 9 0 14 13 2
5 15 13 10 9 2
13 15 13 10 3 9 7 15 13 15 15 4 13 2
26 15 13 3 0 9 14 13 16 15 4 3 13 15 9 1 9 7 10 0 9 1 10 9 4 13 2
30 10 9 4 4 13 1 7 13 1 1 10 0 9 1 0 9 3 15 4 13 10 9 1 0 9 1 10 0 9 2
13 10 9 1 9 4 4 13 16 13 10 9 9 2
47 15 13 10 9 9 2 10 13 9 2 1 0 9 3 1 9 2 3 13 10 9 9 1 15 15 13 9 13 2 3 10 9 9 2 3 15 13 10 9 1 9 3 16 9 3 13 2
17 15 4 3 13 3 0 1 15 9 16 15 13 1 10 11 9 2
16 16 15 13 1 15 9 9 2 10 9 13 9 7 10 9 2
16 10 0 9 13 16 15 4 13 10 0 9 1 10 0 9 2
28 15 9 3 13 10 9 16 15 13 9 9 7 3 0 9 16 15 9 14 9 13 1 9 7 3 0 9 2
22 16 15 13 15 9 2 15 3 3 13 3 1 15 9 9 7 13 3 0 15 13 2
15 3 15 13 10 0 9 9 13 9 1 9 15 13 15 2
14 16 15 4 13 10 9 2 15 3 13 10 0 9 2
11 7 9 13 3 0 7 15 13 3 0 2
12 15 13 15 13 12 9 1 15 9 0 9 2
8 15 13 1 15 9 2 9 2
8 15 13 3 15 4 13 3 2
2 9 2
17 15 13 15 1 9 7 9 3 2 3 15 4 3 13 7 13 2
10 6 2 15 4 13 14 13 15 0 2
20 15 4 13 10 9 1 10 0 9 2 7 15 4 3 13 0 9 7 9 2
26 15 13 15 9 2 13 15 9 14 9 2 3 15 13 3 10 9 16 15 13 14 13 15 10 9 2
20 6 2 3 12 9 3 15 13 3 7 13 15 9 14 9 7 13 3 0 2
27 15 3 13 15 3 15 13 2 7 15 13 15 3 3 12 0 2 0 2 9 13 9 16 15 13 3 2
15 15 4 3 3 13 1 15 9 14 0 9 7 15 13 2
29 2 6 2 16 15 3 3 13 14 13 15 15 4 13 3 7 13 15 1 7 3 15 4 13 10 9 3 2 2
20 15 4 3 13 3 3 15 4 3 13 1 10 9 16 15 13 10 0 0 2
2 6 2
62 6 2 3 15 13 1 13 12 9 1 1 15 9 14 9 2 15 4 3 13 16 10 9 13 15 2 7 13 15 14 13 15 1 10 0 9 2 3 15 13 10 9 2 3 15 13 10 0 9 6 2 7 15 4 13 3 3 7 13 15 3 2
14 15 13 15 14 13 14 13 6 12 9 16 15 13 2
37 3 2 15 13 10 9 14 13 16 15 13 0 7 15 13 14 13 15 13 3 1 10 9 3 15 13 3 0 1 9 15 13 14 13 1 3 5
25 6 2 3 15 13 12 9 3 3 15 13 7 13 10 9 2 7 15 3 4 14 13 1 3 2
14 15 4 14 13 16 15 4 13 15 3 9 7 14 2
34 15 13 10 9 1 9 13 14 13 16 15 13 15 2 7 15 13 0 16 15 13 10 9 7 3 15 13 10 15 13 1 10 9 2
28 1 10 0 9 3 2 16 15 13 10 9 15 4 3 4 13 1 1 3 16 15 4 14 13 10 9 13 2
22 15 4 14 13 15 9 3 16 15 13 10 0 9 15 4 13 15 3 1 15 9 2
8 15 13 10 9 7 9 9 2
12 6 2 15 4 13 10 9 1 15 3 3 2
9 13 15 1 9 16 15 13 2 5
33 6 2 6 3 3 16 15 13 10 0 9 16 13 10 9 3 2 15 13 14 10 9 2 15 13 3 3 13 9 1 10 9 2
20 15 4 13 10 9 3 0 16 10 9 13 3 16 15 4 13 12 0 9 2
29 10 9 15 13 15 4 14 13 10 9 3 13 16 15 2 4 14 13 14 13 15 2 1 15 9 14 0 9 2
21 15 13 3 10 0 9 15 4 13 15 9 14 9 16 15 3 13 3 1 15 2
28 10 0 9 15 13 3 1 15 1 10 0 9 13 16 15 0 9 15 13 1 15 4 13 1 1 15 0 2
24 3 2 15 13 15 9 1 10 9 1 12 9 2 3 15 13 15 15 13 10 0 9 2 2
16 10 2 15 4 13 13 10 0 9 10 13 13 1 10 9 2
10 3 2 3 15 13 3 1 10 9 2
21 6 2 13 1 2 15 13 14 16 15 13 10 9 10 13 3 7 13 15 6 2
10 15 4 13 10 9 1 3 12 9 2
16 15 13 12 2 3 6 15 13 3 9 3 15 13 10 0 2
9 15 13 10 0 9 0 1 15 2
8 7 6 2 15 4 13 15 2
22 14 13 11 11 2 6 15 4 13 1 15 5 15 13 15 13 10 15 4 13 1 2
31 1 10 0 9 2 15 4 3 3 3 13 15 7 13 6 15 13 0 3 3 2 15 4 13 15 3 15 4 13 3 2
13 7 3 3 16 13 9 13 2 15 13 10 9 2
9 15 4 3 13 15 3 3 3 2
20 15 13 3 3 2 6 2 15 9 13 14 4 13 2 3 13 10 9 2 2
10 7 15 3 13 3 1 10 0 9 2
9 15 4 13 15 1 15 13 0 2
7 13 16 15 3 13 15 2
13 7 15 13 14 13 15 4 15 13 10 0 9 2
11 4 15 13 13 1 2 9 2 1 15 2
7 7 13 15 14 15 9 2
5 7 13 15 0 2
8 16 15 13 15 15 4 13 2
23 15 4 13 16 15 4 14 13 15 1 1 11 13 15 3 15 4 4 13 0 14 13 2
27 15 13 15 13 10 9 1 1 10 9 1 10 9 14 13 3 7 13 15 6 15 4 13 15 11 11 2
20 9 2 15 3 4 14 13 15 9 13 1 9 16 4 13 16 12 9 13 2
32 15 4 13 9 13 9 1 15 0 7 13 3 3 16 12 9 13 3 16 15 4 13 3 12 7 12 15 4 4 13 3 2
29 15 3 4 13 15 13 10 9 3 1 1 10 9 14 9 9 7 15 13 10 13 9 15 4 13 14 13 15 3
43 3 15 13 0 1 15 0 9 15 9 13 10 9 13 11 2 2 1 15 15 4 14 13 15 13 10 9 13 15 9 1 15 9 2 0 1 10 9 1 9 1 9 2
37 15 13 1 15 9 0 7 13 12 9 2 7 15 10 13 3 1 10 0 2 7 10 12 1 15 13 10 9 7 13 1 0 1 10 9 2 5
10 3 3 13 15 15 4 4 13 1 2
6 7 15 13 9 3 2
9 15 13 10 9 16 13 15 9 2
35 6 12 9 15 13 1 15 15 13 15 4 14 13 9 16 15 4 13 3 13 1 15 9 14 0 0 9 2 7 15 13 6 6 6 2
24 15 13 0 15 9 4 13 15 16 15 4 14 13 15 0 9 15 13 15 9 4 3 13 2
45 6 12 9 3 3 15 13 3 3 15 4 3 13 1 15 9 14 0 11 7 15 13 3 7 6 15 13 9 1 15 9 1 10 0 9 15 13 1 13 7 15 13 6 15 2
21 15 13 1 6 15 4 13 15 9 9 2 15 13 1 6 4 15 13 15 9 2
16 15 13 10 0 9 14 13 2 7 15 13 15 13 15 9 2
38 7 16 15 13 9 3 13 1 15 2 10 0 9 15 13 15 15 4 13 15 15 13 14 4 13 1 10 9 15 15 13 1 16 15 13 15 1 2
15 15 13 0 2 7 3 13 15 13 14 10 9 1 15 2
75 6 15 4 13 0 1 15 2 15 9 3 13 15 9 1 15 2 3 10 0 9 16 15 13 10 9 7 12 9 2 6 2 15 13 16 15 4 13 3 0 3 15 4 13 10 9 3 7 16 3 10 9 13 15 10 9 7 4 14 13 10 9 16 15 4 14 13 14 3 13 16 15 14 13 2
23 1 10 9 1 9 1 10 9 2 7 9 2 9 9 2 15 4 13 10 3 0 9 2
15 13 9 3 16 15 4 13 7 13 15 13 3 3 3 2
48 0 7 14 2 15 4 13 10 0 9 16 15 4 13 10 0 9 1 9 15 13 14 4 13 15 0 1 2 16 15 4 13 7 13 14 13 15 3 7 14 2 15 4 14 13 9 3 2
27 15 13 2 3 3 2 15 9 2 7 16 15 13 15 14 13 10 9 3 1 9 4 15 13 0 9 2
7 9 2 9 13 1 15 2
5 4 13 9 0 2
16 15 13 10 9 14 13 1 10 3 0 12 9 9 1 0 2
12 15 13 14 0 2 7 15 4 4 13 9 2
8 3 13 15 10 9 4 13 2
24 15 13 10 12 9 9 10 13 10 1 15 9 9 1 10 0 9 1 12 5 12 9 3 2
30 15 13 15 1 1 0 0 9 2 16 15 13 15 10 9 13 7 10 0 9 9 13 0 7 15 13 10 9 9 2
18 3 15 13 15 1 10 9 10 9 1 11 14 4 13 1 10 9 2
31 15 13 15 3 10 9 1 10 9 7 15 4 13 10 9 7 13 15 16 4 13 9 2 15 13 15 14 13 10 2 2
24 15 4 3 13 10 9 9 1 10 0 9 1 15 9 7 13 14 4 13 9 1 10 9 2
13 13 15 1 10 9 9 7 15 13 10 9 9 2
25 15 4 13 10 15 9 7 4 14 13 10 2 7 4 14 13 9 1 9 1 9 14 13 15 2
14 15 13 0 13 1 15 9 9 7 4 13 9 9 2
23 10 0 0 9 10 15 13 13 16 15 3 13 15 9 7 3 13 0 1 15 0 9 2
24 10 9 15 4 13 1 10 9 9 3 1 10 13 9 9 13 1 1 15 0 9 1 9 2
12 15 4 14 13 14 13 15 13 0 1 15 2
25 6 2 15 4 14 13 10 9 9 7 4 13 10 0 9 9 7 15 9 13 10 0 0 9 2
15 15 13 14 14 13 10 9 9 16 15 13 10 0 9 2
17 15 4 3 13 10 9 0 1 10 9 9 2 7 10 9 9 2
27 15 13 10 1 15 9 7 15 3 13 15 10 9 14 13 15 13 1 1 10 9 1 9 1 15 9 2
13 3 15 4 13 10 9 7 13 15 15 4 13 2
28 15 4 4 13 1 15 9 3 7 16 15 4 13 15 2 13 10 0 9 9 13 1 9 7 10 9 9 2
17 4 4 13 10 9 1 10 9 9 10 9 4 3 13 3 3 2
7 15 0 9 4 13 9 2
22 15 4 4 13 15 0 9 2 9 3 14 13 10 9 3 3 16 15 4 13 15 2
4 3 10 9 2
6 13 15 4 13 15 2
2 11 2
9 9 13 1 1 9 7 14 0 2
11 9 13 0 14 13 15 8 3 1 15 2
11 15 4 4 13 15 9 7 9 1 15 2
26 0 13 1 0 2 15 13 1 1 10 5 5 7 13 14 13 15 1 3 7 13 10 0 9 9 2
13 15 4 3 0 3 7 14 13 0 9 1 9 2
31 15 13 10 9 10 15 3 4 14 13 0 14 13 7 3 16 15 13 12 12 1 9 15 13 3 1 1 15 9 9 2
20 15 13 15 10 9 4 13 1 9 12 7 12 2 15 13 14 15 14 13 2
22 15 13 10 9 10 4 14 13 14 13 9 0 1 15 16 9 15 4 14 13 3 2
25 15 4 13 9 7 15 3 13 10 9 9 1 15 9 1 10 9 16 15 4 14 13 0 9 2
22 15 4 14 13 15 4 13 0 14 13 15 9 3 3 3 16 15 4 13 10 9 2
15 15 4 14 13 14 13 13 1 10 9 15 4 14 13 2
11 15 13 0 14 13 10 9 9 7 13 2
9 10 9 13 10 9 15 13 0 2
21 15 4 3 4 13 15 0 9 3 15 13 10 9 7 9 14 13 15 1 9 2
32 11 13 3 15 13 14 13 0 9 7 10 9 7 9 3 13 15 13 3 10 9 9 1 9 1 10 9 1 10 0 9 2
35 15 4 3 13 9 9 7 10 9 9 2 1 10 0 9 9 7 10 9 1 9 1 10 0 9 2 10 4 7 4 14 4 13 2 2
7 10 9 13 14 1 9 2
5 15 4 14 13 2
4 15 4 13 9
7 10 9 13 14 1 9 2
5 15 4 14 13 2
24 15 4 13 9 2 7 3 1 15 13 16 13 1 10 9 14 7 4 13 3 1 12 9 2
8 15 4 14 13 15 3 3 2
18 15 13 16 15 13 10 9 16 13 15 7 3 13 14 13 15 1 2
18 1 10 0 9 15 4 13 9 15 4 13 9 13 3 3 1 9 2
9 15 13 15 4 13 14 13 0 2
9 15 13 0 14 13 15 10 9 2
22 11 2 15 4 3 13 10 0 9 7 4 13 1 9 9 1 10 9 9 3 3 2
9 13 1 9 2 9 9 7 0 2
10 15 4 13 10 9 9 13 16 13 2
27 10 9 2 9 4 13 3 14 13 10 9 1 9 10 4 3 13 1 0 9 7 4 4 13 1 9 2
14 16 15 13 10 9 3 9 4 14 13 14 13 15 2
10 15 13 3 12 1 10 0 9 1 9
39 15 13 15 13 3 0 16 15 4 13 1 10 9 9 0 7 4 13 10 9 1 0 9 2 7 10 9 1 9 2 16 15 13 14 13 10 9 1 2
35 15 4 13 10 11 9 13 14 13 1 15 9 9 16 15 4 14 13 3 13 10 9 1 1 10 9 7 13 15 0 0 9 13 9 2
21 0 9 9 15 13 1 9 7 16 13 9 1 9 15 13 14 13 10 9 1 2
8 13 15 9 15 13 1 1 2
24 16 3 13 1 15 7 15 4 13 15 10 10 0 9 15 4 16 15 13 1 15 13 3 2
26 15 13 0 14 13 14 13 10 9 1 7 3 13 14 13 15 1 2 7 10 9 13 0 10 9 2
18 16 15 13 10 9 13 0 15 3 15 13 15 9 4 13 9 1 2
17 1 1 9 16 11 13 13 1 11 15 4 13 14 13 1 15 2
8 3 3 10 0 9 4 3 2
25 15 0 13 9 9 13 3 3 15 13 10 9 1 10 11 7 3 10 0 9 9 9 1 11 2
12 15 13 10 9 1 11 7 13 15 13 3 2
13 10 9 13 1 9 7 15 4 14 13 0 9 2
19 15 4 13 10 0 1 3 2 7 9 16 15 9 9 13 13 1 11 2
41 15 13 10 9 16 15 13 0 7 9 4 13 10 0 9 16 13 1 9 3 16 15 13 9 13 9 2 7 15 4 14 13 10 9 9 1 3 3 12 9 2
26 15 4 13 10 1 15 9 9 4 13 3 3 15 4 13 0 9 16 11 13 7 3 13 1 9 2
13 12 9 3 13 15 9 9 16 4 13 1 9 2
19 15 4 3 13 0 0 9 10 13 3 1 9 9 1 12 2 12 9 2
20 10 0 9 15 13 13 16 10 9 9 13 14 13 3 1 10 0 9 3 2
33 15 4 3 13 9 7 10 9 10 0 0 9 1 10 3 0 9 13 10 9 1 0 9 14 13 10 0 9 1 10 0 9 2
5 15 4 14 13 2
15 11 13 10 9 1 9 9 1 16 3 0 15 13 3 2
23 15 4 13 14 13 16 15 4 13 1 9 1 15 9 9 7 13 10 9 1 10 9 2
17 15 13 15 13 0 9 13 16 11 11 13 3 4 13 13 9 2
29 15 13 15 13 10 0 9 13 10 0 9 1 0 9 9 3 2 7 15 4 13 10 9 16 10 9 4 13 2
16 10 9 16 15 13 10 9 9 1 9 4 15 13 11 11 2
15 11 11 4 13 9 0 9 7 4 14 3 13 10 9 2
9 13 15 13 15 15 13 14 13 2
25 15 13 14 13 0 4 13 2 7 3 15 4 14 13 15 4 13 1 10 9 3 3 10 9 2
11 3 15 13 15 4 3 13 16 13 3 2
17 15 4 13 15 9 3 16 15 13 16 15 13 10 9 7 14 2
42 16 15 13 10 0 9 2 10 15 13 0 15 13 2 1 15 2 15 4 13 0 16 16 10 9 13 0 1 10 9 2 14 3 0 15 15 13 14 13 1 15 2
37 3 16 15 4 13 1 15 13 0 1 10 0 9 2 15 13 3 10 9 1 9 7 3 9 3 15 4 13 14 13 13 3 3 1 10 9 2
16 3 10 1 10 2 13 10 9 1 9 16 13 1 10 9 2
20 10 0 13 1 1 9 3 4 3 13 15 9 16 10 9 13 1 15 9 2
13 4 15 4 13 10 9 1 10 9 13 10 9 2
5 7 10 0 9 2
6 13 15 3 1 15 2
7 7 4 15 13 1 9 2
12 15 3 13 16 15 4 4 13 10 0 9 2
21 15 13 16 15 4 14 13 14 13 15 13 16 15 4 14 13 15 1 10 9 2
14 15 13 15 10 9 4 13 2 7 15 4 13 0 2
4 3 0 9 9
17 4 14 13 1 10 9 2 3 16 15 13 14 13 15 9 13 2
29 15 13 10 3 0 9 1 15 9 7 13 3 0 3 15 13 3 14 13 15 3 15 4 14 13 1 15 9 2
7 0 2 0 2 0 9 2
2 0 9
19 11 11 13 15 9 1 10 9 9 7 13 3 3 0 1 10 0 9 2
24 15 4 14 13 9 9 7 0 9 2 15 13 15 9 9 10 13 0 7 10 9 13 0 2
5 15 9 13 0 2
7 15 13 15 15 4 13 2
3 15 9 12
12 15 3 13 15 9 1 12 7 13 3 0 2
13 11 7 9 13 10 10 15 13 7 12 9 0 2
6 10 9 13 8 0 2
18 16 15 13 10 9 10 13 0 7 0 14 13 1 15 13 10 9 2
5 9 3 11 14 2
1 11
3 0 9 9
15 15 3 13 10 9 13 1 11 7 15 4 14 13 0 2
9 15 13 3 0 16 15 3 13 2
16 10 9 13 0 2 10 9 13 0 7 10 9 13 0 9 2
16 15 4 3 13 10 9 1 9 13 14 13 10 0 9 13 2
3 0 7 0
10 15 13 14 13 9 1 10 9 15 2
12 7 15 13 10 9 0 7 10 9 3 0 2
17 3 13 10 9 1 10 9 7 13 15 3 0 3 9 13 0 2
6 13 10 9 7 9 2
12 1 1 10 9 15 13 15 1 10 12 9 2
3 0 9 9
20 15 4 13 11 11 11 0 9 3 7 15 4 13 0 9 1 15 12 9 2
10 11 13 0 7 13 0 9 1 9 2
19 10 0 9 13 14 1 3 3 15 13 15 9 7 3 3 15 13 15 2
5 15 3 13 15 2
31 15 13 11 11 11 7 11 7 11 7 11 11 11 7 11 11 1 11 2 11 13 15 11 11 11 11 1 3 0 9 2
18 15 13 15 9 7 15 4 13 1 9 9 7 11 9 9 1 0 2
6 9 1 11 11 11 2
5 10 9 13 0 2
12 15 13 15 9 9 1 3 0 1 10 9 2
25 10 9 13 1 9 7 4 14 13 10 9 2 15 13 3 14 13 7 13 10 9 3 7 3 2
13 15 4 14 13 3 0 1 10 9 15 9 13 2
4 0 9 9 2
2 9 5
34 15 4 13 11 11 10 9 5 16 10 9 13 0 1 9 0 2 15 13 15 9 3 10 0 9 2 7 10 9 15 13 13 0 2
21 15 13 10 9 14 13 9 1 15 1 15 9 2 15 4 13 15 13 1 15 2
1 11
5 10 9 13 0 2
8 9 3 13 3 0 7 0 2
23 15 13 0 14 13 15 4 13 0 9 2 0 9 2 7 1 10 0 9 10 1 12 2
15 15 4 13 9 15 13 3 7 15 10 13 10 0 9 2
10 15 4 4 13 3 1 9 14 13 2
3 0 9 11
19 11 0 9 11 11 13 3 0 16 3 13 15 9 7 13 10 0 9 2
33 1 10 0 0 9 9 2 15 4 13 10 0 0 2 9 2 2 13 10 9 0 2 1 15 9 14 13 10 3 0 9 0 2
3 9 13 0
24 15 4 13 3 12 1 12 9 7 10 9 9 15 13 13 13 1 7 13 16 15 13 15 2
12 15 13 15 9 0 10 9 3 0 7 0 2
6 9 7 9 13 0 2
14 15 4 13 0 16 15 4 13 3 9 13 13 0 2
1 11
4 0 7 0 9
16 15 13 1 11 14 1 11 7 13 15 0 9 14 9 13 2
22 15 13 0 1 9 1 10 9 1 10 0 9 15 13 2 7 15 9 13 0 9 2
7 3 1 9 7 0 9 2
11 13 3 14 13 10 0 9 13 10 9 2
4 15 13 11 11
9 15 13 11 7 15 9 13 15 2
11 15 3 13 14 13 1 9 1 10 9 2
20 15 4 13 15 0 9 1 9 7 13 3 16 13 15 9 7 9 10 9 2
14 15 9 13 0 10 9 3 15 13 1 7 13 1 2
5 11 11 0 7 0
40 15 13 11 11 11 7 1 12 9 11 4 13 1 15 9 7 9 13 10 15 15 13 10 11 9 9 9 9 2 7 13 10 9 1 3 12 9 1 9 2
7 0 2 0 7 0 9 2
3 3 0 2
3 3 13 2
4 15 0 9 2
21 15 13 1 11 11 14 13 1 9 2 7 15 9 4 13 15 9 9 1 3 2
7 15 13 0 7 13 3 2
19 3 16 15 13 3 2 15 13 15 0 9 14 13 9 1 9 7 9 2
9 9 3 2 0 9 1 10 9 2
4 15 13 11 14
6 0 9 7 0 9 2
23 15 13 3 3 10 9 14 13 9 1 15 7 15 9 7 10 9 1 11 14 13 0 2
6 15 13 0 7 0 2
17 15 4 3 13 10 9 1 15 9 16 15 3 13 1 10 9 2
4 15 13 0 2
58 13 10 9 9 1 10 9 2 13 10 9 9 1 10 9 9 1 11 2 7 15 9 3 13 15 1 10 0 9 2 3 15 13 12 12 9 9 1 10 11 11 11 14 13 10 9 16 13 9 2 7 13 15 3 0 7 0 2
3 0 9 2
7 11 11 13 10 0 9 2
7 15 4 13 15 1 9 2
19 15 4 13 0 9 9 1 10 9 15 4 3 13 7 3 13 14 13 2
26 15 13 1 10 9 9 1 12 5 12 1 12 7 15 13 0 14 13 1 10 11 3 10 9 3 2
2 0 9
6 11 11 13 10 0 2
5 0 2 0 9 2
3 0 9 2
3 0 9 2
13 3 3 4 0 4 13 1 10 9 1 10 9 2
18 15 4 13 15 3 2 13 2 1 2 13 16 15 3 13 9 3 2
11 15 4 13 10 0 14 13 0 1 15 2
7 0 9 14 13 15 0 9
11 15 4 3 13 10 0 9 13 1 11 2
11 15 13 9 9 12 15 4 13 1 15 2
23 15 13 7 13 11 11 7 13 16 15 4 3 13 0 9 1 15 7 13 1 15 9 2
8 13 15 3 1 0 9 9 2
5 11 11 11 9 9
35 11 1 11 11 11 11 2 13 10 3 0 9 3 3 2 10 9 2 13 10 9 1 15 7 15 13 15 3 3 2 0 9 0 9 2
3 3 13 2
3 9 11 2
12 11 2 0 11 11 11 9 2 1 0 9 2
58 1 10 0 0 9 13 3 0 14 13 9 3 0 9 0 9 9 10 9 9 15 13 10 10 10 9 1 9 3 0 15 3 13 10 15 9 4 14 4 13 1 0 9 10 15 13 10 9 1 9 14 13 1 9 1 10 9 9
2 0 9
15 13 10 9 1 10 9 7 15 13 14 13 15 13 0 2
36 15 13 14 13 12 1 10 0 9 10 15 4 13 1 1 10 0 9 2 10 9 13 0 7 15 13 10 3 0 9 7 10 0 9 9 2
11 0 9 0 9 7 15 0 4 15 13 2
3 0 0 0
14 10 9 13 1 3 10 0 11 9 15 4 13 1 2
22 10 9 13 3 0 2 10 9 13 3 3 0 2 7 10 10 9 13 13 10 9 2
10 3 0 7 15 4 14 13 1 15 2
14 13 15 10 0 11 14 13 1 1 11 2 11 11 2
5 0 0 9 9 2
29 11 11 11 13 9 2 13 15 0 9 16 13 0 7 0 9 9 2 9 2 9 2 9 9 9 2 7 0 2
11 15 13 0 9 1 9 7 13 1 9 2
16 15 13 13 1 10 0 7 0 9 9 7 4 13 1 9 2
2 0 9
7 15 13 9 9 13 3 2
7 11 11 7 9 13 0 2
18 15 13 0 1 15 9 7 13 1 15 9 14 13 9 1 10 9 2
14 11 11 13 10 9 1 9 7 13 15 9 1 15 2
9 9 13 9 9 7 13 3 0 2
5 9 13 3 0 2
6 10 0 1 10 9 2
21 15 4 13 1 10 10 0 9 9 1 10 9 7 11 11 13 1 3 10 0 2
13 15 13 3 0 1 10 9 10 15 13 1 15 2
11 10 9 13 0 7 10 9 13 3 0 2
13 15 4 13 10 9 1 9 13 14 13 10 9 2
9 11 2 12 9 1 11 11 11 2
11 10 9 4 13 10 0 9 1 15 9 2
13 15 4 13 10 12 1 15 9 13 11 11 11 2
21 10 9 4 3 13 7 15 4 13 3 0 1 10 9 2 10 9 7 10 9 2
7 0 9 2 11 11 11 2
4 0 9 7 9
6 10 9 13 3 0 2
17 15 13 10 0 9 1 9 1 3 1 10 9 1 10 0 9 2
27 10 9 13 15 13 3 0 7 13 3 0 2 16 15 13 3 0 7 4 14 13 9 3 3 1 9 2
9 13 1 15 9 9 10 11 9 2
2 9 5
7 0 9 9 7 0 9 2
16 10 9 1 11 11 13 15 9 13 1 3 1 15 13 9 2
19 15 13 0 1 2 0 2 9 1 2 13 2 9 7 13 3 0 9 2
18 10 10 0 9 3 3 16 9 9 7 11 11 7 11 3 1 9 2
6 13 14 13 1 1 9
16 15 13 3 15 13 1 15 2 3 3 1 15 13 9 9 2
16 15 9 13 0 2 0 7 13 16 15 4 13 1 10 9 2
6 15 4 14 13 9 2
7 15 13 10 9 9 9 2
13 10 9 13 10 9 1 11 2 0 1 10 9 2
13 3 3 4 15 13 1 5 12 7 13 10 9 2
10 0 9 1 0 9 3 3 1 11 2
14 15 4 13 1 10 0 9 7 10 0 9 9 9 2
28 15 4 13 12 9 3 1 11 7 4 13 0 1 0 9 5 9 7 4 14 13 10 9 1 9 7 9 2
7 13 1 10 12 2 9 9
6 15 4 14 13 15 2
27 10 9 13 0 2 1 10 0 9 7 0 9 2 7 10 9 13 0 2 7 3 15 9 9 9 2 2
24 6 2 10 9 13 10 0 0 2 7 13 3 2 4 15 3 13 3 14 13 1 11 3 2
17 15 4 3 13 0 9 1 11 2 15 4 13 7 13 10 9 2
37 15 3 13 11 2 15 13 10 0 9 2 15 2 13 2 10 9 15 13 15 9 2 3 0 7 13 13 15 9 14 13 0 15 9 13 0 2
8 15 3 13 13 15 9 9 2
6 0 0 9 1 10 9
12 10 9 3 13 0 7 0 1 1 10 9 2
12 10 9 4 13 3 1 10 12 9 1 9 2
16 10 9 9 13 0 9 16 0 9 4 13 1 3 5 12 2
21 15 13 0 10 9 1 9 1 10 9 2 10 9 13 0 7 10 9 13 0 2
3 0 9 2
22 15 13 10 0 9 2 15 4 4 13 11 1 3 12 9 7 4 14 13 3 3 2
24 15 13 10 9 1 9 7 10 9 1 10 9 13 1 11 10 13 10 9 3 1 10 9 2
15 10 9 13 3 13 7 13 0 16 13 10 9 1 9 2
58 15 13 10 9 1 9 1 15 9 9 7 16 15 4 14 13 15 1 10 9 2 16 15 9 9 13 1 10 0 9 2 2 15 13 15 1 9 1 0 9 1 10 9 9 9 7 3 15 4 3 13 11 1 15 0 9 9 2
2 3 13
7 15 3 13 3 7 3 2
24 1 9 2 15 3 13 14 13 15 9 2 7 15 13 1 1 15 9 14 13 9 1 15 2
21 3 2 3 15 13 9 2 15 9 2 2 15 13 15 9 1 1 10 13 9 2
9 15 4 13 12 5 0 7 0 2
3 3 13 2
3 9 9 9
16 3 2 4 15 13 13 14 13 1 10 0 0 9 1 9 2
25 15 4 4 13 14 16 16 10 9 10 9 15 13 15 4 14 13 0 9 1 9 1 10 9 2
13 11 11 13 3 7 13 15 9 9 1 10 0 2
4 7 15 13 2
4 13 15 11 11
6 0 2 0 9 1 9
9 15 13 12 11 9 10 15 13 2
12 15 13 10 9 1 9 13 10 0 9 9 2
24 15 3 13 16 9 9 13 0 1 9 9 7 14 3 11 9 2 9 7 3 0 2 9 2
13 7 10 9 13 10 0 9 9 15 4 13 3 2
8 13 10 9 2 15 13 10 0
3 3 0 2
11 0 2 13 9 2 0 9 2 0 9 2
11 9 13 3 0 2 13 15 1 10 9 2
8 4 14 13 1 10 0 9 2
13 4 4 13 3 10 7 10 9 15 13 3 3 2
14 3 2 11 13 10 0 9 15 4 13 10 0 9 2
3 9 13 3
5 15 13 11 11 2
54 11 11 10 9 7 9 13 0 9 1 15 9 2 16 15 13 1 0 9 2 3 0 2 0 9 15 13 0 9 1 11 11 16 15 13 3 0 9 4 13 0 0 9 3 15 13 11 3 7 15 4 3 13 15
7 0 9 2 4 14 13 2
10 4 14 15 13 10 0 9 1 9 2
16 15 13 3 0 2 7 15 13 10 0 9 3 7 3 3 2
8 10 9 13 0 7 3 0 2
10 10 9 1 9 7 9 4 13 15 2
6 13 10 9 2 9 2
13 11 7 11 12 13 15 3 2 3 4 14 15 2
3 9 13 9
16 15 3 13 1 10 9 3 1 9 14 13 1 10 11 9 2
11 15 13 10 9 2 10 9 7 10 9 2
16 9 13 1 10 9 13 9 10 3 13 10 9 1 9 2 2
12 10 11 2 11 2 7 11 14 13 15 9 2
10 7 9 1 15 4 3 13 3 3 2
6 10 9 3 13 0 2
16 16 10 0 9 13 2 10 9 9 4 13 1 10 0 9 2
13 15 13 12 5 0 1 11 11 14 0 9 9 2
19 10 0 9 13 15 13 10 9 13 0 2 7 9 3 13 0 0 0 2
10 13 3 3 3 16 15 9 13 3 2
1 8
2 0 2
9 6 15 9 12 9 4 3 13 2
9 15 13 0 14 13 15 5 12 2
6 7 15 13 5 12 2
10 15 13 15 16 13 14 13 1 11 2
17 11 13 14 13 1 15 9 7 15 4 14 13 14 13 1 15 2
6 12 9 8 13 15 2
3 0 9 2
7 15 4 13 15 1 9 2
4 0 0 9 2
20 15 4 14 13 3 1 11 9 2 3 16 15 13 10 10 0 9 1 9 2
25 0 9 9 7 0 9 7 13 15 13 10 9 0 1 15 9 9 2 16 9 13 10 0 9 2
18 2 0 9 2 9 9 2 9 2 0 9 2 7 9 7 0 9 2
7 15 9 7 9 13 0 2
6 7 9 13 3 0 2
6 9 1 9 3 0 2
5 3 13 10 9 2
6 3 3 13 0 9 2
7 3 0 1 10 9 9 2
6 9 9 13 3 0 2
6 3 16 15 13 1 2
14 14 13 10 9 15 4 13 14 13 1 9 1 9 2
5 7 3 13 3 2
3 14 0 2
57 11 1 11 1 11 13 15 9 16 15 13 15 9 13 7 13 1 10 9 15 13 3 0 7 10 9 13 0 7 15 4 4 13 3 3 1 12 9 3 0 7 15 13 1 15 9 13 15 9 13 1 15 9 15 13 0 2
7 7 15 9 13 3 0 2
4 0 9 1 9
17 15 13 10 9 3 11 11 4 13 0 9 1 10 0 0 9 2
6 9 3 13 3 0 2
7 9 13 0 7 13 3 2
19 10 9 9 13 1 0 2 15 13 15 9 3 15 13 1 10 9 2 2
13 16 15 13 0 9 3 11 13 10 9 14 13 2
41 15 4 14 13 1 13 15 9 3 2 7 15 4 13 10 9 15 13 1 15 13 3 0 2 15 13 0 14 13 10 9 1 10 9 10 13 10 9 1 15 2
26 3 15 4 13 15 9 1 9 7 0 0 9 9 1 0 2 3 16 15 4 14 13 15 9 3 2
5 10 0 9 1 9
16 16 15 13 9 1 11 2 13 0 15 13 1 11 14 3 2
22 15 9 13 0 2 3 15 15 13 1 10 13 9 4 3 13 0 3 1 10 9 2
11 15 13 15 1 13 9 9 7 9 9 2
14 13 15 2 15 13 3 3 7 15 4 3 13 3 2
3 0 9 9
12 15 9 4 13 9 10 9 1 10 0 9 2
21 15 13 10 9 9 3 15 13 14 0 15 15 4 13 1 3 15 13 1 9 2
18 10 9 13 3 0 7 13 15 3 15 15 13 1 15 0 9 9 2
7 10 9 1 11 13 0 2
7 15 4 13 15 1 9 2
10 0 9 7 9 1 10 3 0 9 2
9 10 9 13 0 9 7 3 0 2
12 15 4 13 15 9 3 7 13 10 0 9 2
20 15 4 3 13 3 10 9 1 9 14 13 10 9 3 7 9 13 3 0 2
17 9 16 13 3 0 9 1 15 0 9 1 9 10 3 13 0 2
8 13 11 1 11 1 12 9 2
13 3 1 9 7 3 1 9 3 0 9 10 9 2
12 10 9 4 14 3 13 10 9 1 9 9 2
27 9 2 15 13 0 9 1 10 9 2 1 12 7 12 9 2 7 3 13 3 14 13 15 9 1 9 2
9 15 13 14 10 9 14 4 13 2
35 15 13 10 0 9 7 13 0 14 13 15 0 9 3 15 13 10 9 9 9 7 15 4 13 15 3 13 1 15 9 7 13 15 13 2
28 1 3 15 4 13 14 13 15 13 15 0 9 9 3 3 16 15 13 0 7 4 3 3 13 10 10 9 2
3 0 9 2
22 15 3 13 15 9 13 1 11 11 7 4 13 16 15 13 3 0 1 10 0 9 2
32 1 10 9 1 9 13 1 15 14 13 9 1 10 0 9 2 1 10 9 1 10 9 9 1 10 0 9 1 10 9 15 2
7 15 13 9 0 14 13 2
8 3 0 16 15 13 1 15 2
3 10 9 9
24 9 13 14 4 13 10 0 9 13 7 13 1 10 0 2 16 15 7 0 9 4 3 13 2
21 10 9 1 10 9 13 3 1 10 9 7 3 13 14 13 10 9 9 14 9 2
20 15 13 14 16 15 13 1 7 13 1 10 9 1 9 13 4 15 13 15 2
6 4 14 13 15 9 3
10 15 13 10 9 1 11 1 10 9 2
6 6 2 15 13 15 2
17 3 2 1 10 9 2 15 13 15 15 4 14 13 15 9 13 2
24 3 2 15 13 15 0 9 2 0 1 9 9 9 2 16 16 15 9 4 13 15 3 3 2
7 15 13 1 13 3 0 2
5 4 15 13 15 2
6 15 4 14 13 15 2
15 0 7 0 9 2 13 2 2 2 0 9 2 0 9 2
18 15 13 1 10 9 7 15 13 10 9 1 9 1 15 9 9 9 2
10 10 9 15 13 10 0 9 13 0 2
17 16 15 13 10 0 10 11 13 14 13 2 15 13 1 1 3 2
13 15 13 1 10 11 1 12 13 1 10 0 9 2
19 11 11 13 15 16 15 9 13 1 9 7 16 15 4 13 15 1 11 2
21 15 4 13 10 9 1 11 11 1 12 9 7 4 13 9 1 9 1 9 8 2
9 15 13 9 1 0 9 1 11 2
8 4 14 13 1 11 11 11 2
2 0 9
14 1 10 9 1 15 15 4 13 10 9 1 0 9 2
39 15 15 13 13 10 5 12 5 9 9 14 13 10 9 1 10 0 12 5 12 9 5 9 10 15 4 3 13 14 13 9 8 2 13 2 10 9 2 2
15 3 1 15 10 9 13 1 10 0 9 7 10 9 13 0
6 13 15 13 1 10 9
8 13 3 1 11 3 11 11 2
9 15 3 13 10 9 1 10 9 2
8 15 13 0 14 13 10 9 2
22 16 15 4 13 1 9 7 13 10 9 9 0 15 13 15 13 2 1 12 9 3 2
14 7 3 1 10 15 9 13 1 10 9 3 10 9 2
4 13 3 3 2
6 13 1 9 2 3 2
3 3 13 2
24 11 13 10 9 9 1 15 9 9 7 15 13 10 3 0 9 7 0 2 0 7 0 9 2
5 10 9 1 9 2
3 3 0 2
3 0 9 2
16 15 3 13 11 7 15 9 9 9 1 0 9 9 7 9 2
5 15 13 15 9 2
3 11 2 11
2 3 0
14 15 13 1 11 2 11 1 10 9 9 1 11 11 2
19 15 13 3 7 10 9 13 3 0 1 15 9 7 10 9 15 13 1 2
12 10 9 13 3 0 2 13 10 9 7 9 2
23 15 13 10 0 9 2 7 15 13 15 4 13 14 13 15 9 2 1 2 9 1 11 2
5 0 9 7 9 2
17 11 11 13 10 9 9 7 15 7 10 9 1 10 9 13 0 2
15 15 13 14 13 15 3 13 3 16 15 13 10 9 9 2
18 16 15 13 3 1 9 3 11 4 13 3 14 13 15 1 3 13 2
9 15 13 16 15 13 10 9 2 2
7 9 4 14 13 3 0 2
4 0 9 1 11
29 10 0 13 2 0 13 9 7 15 0 9 13 10 9 0 2 3 13 2 3 13 9 1 10 3 0 1 9 2
19 13 15 9 2 9 2 10 15 4 13 1 16 13 1 15 0 9 9 2
17 15 13 10 0 9 1 10 9 15 4 13 1 10 1 0 11 2
12 11 11 13 10 0 9 14 13 15 9 13 2
15 15 13 3 0 2 9 13 0 2 7 15 4 3 13 2
23 15 13 10 0 9 1 10 9 2 9 9 10 13 3 5 12 7 15 3 13 12 9 2
4 15 13 15 2
5 9 13 3 0 2
5 13 10 9 1 2
8 15 13 15 4 14 4 13 2
6 0 9 1 10 0 9
5 11 13 3 0 2
17 15 13 15 0 9 1 10 0 9 7 13 15 9 9 3 0 2
33 15 13 3 0 14 13 1 7 13 15 9 9 3 0 7 15 13 10 0 9 2 3 3 1 15 2 7 1 15 9 7 9 2
4 15 13 0 2
7 15 4 13 15 1 9 2
4 3 3 0 2
2 0 2
18 11 12 2 12 0 9 13 1 11 11 11 7 15 13 10 0 9 2
23 1 10 0 9 9 1 10 9 9 9 7 10 9 7 13 1 9 2 10 13 9 13 2
11 3 0 15 13 1 1 10 9 9 9 2
8 3 0 9 15 4 13 15 2
4 9 13 0 2
1 11
3 13 1 11
25 0 9 2 1 10 9 16 13 15 9 10 9 4 13 7 13 3 3 12 9 16 15 4 13 2
25 3 1 15 1 9 1 15 13 9 15 4 14 13 1 9 1 10 9 14 3 13 10 0 9 2
18 15 9 1 10 13 15 4 13 1 10 9 2 6 13 15 13 14 2
7 9 4 13 10 0 9 2
23 11 14 0 12 13 10 0 0 3 3 2 7 10 0 9 9 4 13 9 1 10 9 2
9 10 9 3 3 13 14 4 13 2
11 13 3 7 13 11 10 0 9 3 3 2
23 15 13 10 0 9 16 0 9 14 13 0 1 7 10 10 9 1 12 4 13 3 0 2
3 0 9 2
10 11 11 7 15 9 1 9 13 0 2
27 15 4 4 13 1 9 9 1 3 12 9 7 4 13 1 0 9 2 9 2 9 7 9 1 10 9 2
14 15 13 10 11 9 3 12 9 14 13 15 13 0 2
14 7 3 12 9 1 15 0 9 15 13 0 1 3 2
3 9 9 2
9 15 4 4 13 10 9 7 13 2
10 15 9 7 15 13 3 1 10 9 2
15 15 13 1 10 0 9 9 2 15 13 3 0 7 0 2
11 15 9 13 3 0 7 10 9 13 0 2
18 15 9 4 13 10 0 9 2 3 15 13 10 0 9 1 0 9 2
12 15 13 10 0 2 0 9 1 10 1 15 2
3 0 0 0
26 13 1 3 7 13 15 9 13 13 3 1 10 0 9 3 13 15 3 14 4 13 1 15 10 9 2
22 15 4 14 3 13 15 13 10 9 16 13 15 7 13 15 3 15 4 4 13 15 2
6 15 4 14 13 3 2
7 15 13 14 13 10 9 2
10 13 9 9 7 15 13 3 0 3 2
13 15 13 0 14 13 10 10 10 9 1 9 9 2
29 16 15 13 10 9 1 9 2 11 2 7 13 10 1 10 9 2 8 2 15 4 13 15 13 15 10 9 3 2
28 3 16 13 10 9 1 9 2 15 4 13 16 15 13 10 9 3 0 16 15 13 0 2 9 5 12 2 2
13 10 15 4 13 13 16 15 13 0 15 13 3 2
12 10 9 13 0 1 9 7 10 9 13 0 2
11 10 9 13 1 9 2 3 13 10 9 2
6 10 9 9 13 0 2
21 16 13 1 10 9 7 13 9 9 2 15 13 10 9 15 4 14 13 3 3 2
11 15 4 13 3 7 13 9 1 10 9 2
3 13 15 2
34 15 3 13 10 9 16 15 13 0 14 13 10 0 9 1 9 15 13 2 10 9 2 7 13 15 10 0 9 7 3 10 0 9 2
22 9 0 15 13 10 13 15 4 13 15 7 13 14 13 15 0 7 13 15 0 9 2
7 15 13 10 9 9 3 2
11 15 13 11 11 7 15 13 0 15 13 2
5 10 9 13 0 2
8 15 13 0 2 0 7 0 2
25 10 9 13 0 7 10 9 1 10 9 13 14 3 0 2 6 2 10 9 13 14 3 0 2 2
19 10 9 4 4 13 9 3 2 7 15 3 1 15 2 13 3 9 2 2
20 15 4 13 3 3 1 10 0 9 7 4 14 13 3 7 4 14 13 15 2
11 0 9 1 9 2 0 9 2 0 9 5
9 6 15 13 15 11 1 12 9 2
11 15 4 14 13 7 13 10 9 9 9 2
23 15 4 14 13 9 0 0 14 13 15 3 15 13 15 3 7 15 13 15 1 5 12 2
12 9 9 13 3 3 7 9 1 10 0 9 2
10 0 2 0 9 9 5 13 1 9 2
6 11 14 1 11 2 6
25 15 13 10 0 11 14 9 2 13 1 10 0 9 1 10 0 9 2 7 10 9 13 3 3 2
11 9 1 0 9 7 15 13 13 0 9 2
10 13 1 9 9 2 10 9 4 13 2
13 15 13 0 0 9 1 15 9 9 3 3 3 2
10 3 3 11 14 2 15 4 4 13 2
12 15 13 3 0 1 10 9 1 11 11 11 2
17 15 9 9 13 3 0 16 15 13 10 9 14 13 7 13 15 2
11 15 13 0 9 16 15 13 14 13 15 2
10 15 13 1 9 7 13 15 9 3 2
10 15 13 3 0 3 0 13 15 9 2
14 16 15 13 10 9 1 15 9 2 15 4 13 15 2
7 0 9 3 1 9 9 2
13 15 13 1 1 9 1 10 9 7 13 15 9 2
3 6 6 2
14 15 13 3 12 9 1 9 7 10 9 13 3 0 2
18 15 13 10 9 1 9 1 15 7 13 15 1 10 0 9 1 9 2
18 15 13 15 4 3 13 0 1 10 9 15 4 4 13 10 0 9 2
4 9 11 11 2
1 0
11 15 13 10 0 9 14 13 15 9 13 2
23 15 4 13 3 9 7 9 3 3 15 13 14 13 15 9 13 7 3 15 13 10 9 2
21 3 15 13 15 9 13 3 2 15 13 0 9 9 16 15 4 14 13 15 9 2
19 10 9 13 0 7 1 9 15 13 14 13 0 2 7 10 9 13 0 2
2 3 13
20 15 4 13 1 11 1 15 9 9 7 0 9 1 9 7 4 3 4 13 2
17 3 3 10 9 15 13 1 3 15 13 2 15 3 13 13 0 2
29 15 4 3 3 13 15 1 10 0 9 2 9 7 9 13 9 2 15 13 0 14 13 1 1 15 9 7 3 2
5 15 3 13 15 2
5 0 9 1 11 11
10 10 10 0 9 2 15 13 10 9 2
12 14 10 0 0 9 10 10 10 0 9 13 2
12 15 9 13 3 0 2 0 9 2 0 9 2
37 15 3 13 10 0 9 15 3 13 2 14 3 3 1 10 9 15 13 1 10 9 9 2 15 13 1 8 3 3 16 15 13 0 1 10 9 2
2 10 0
18 11 11 7 15 9 4 13 10 0 9 1 10 9 1 10 15 9 2
22 11 11 13 3 0 7 0 1 10 9 2 7 3 0 7 1 10 9 1 10 9 2
12 15 13 10 0 9 14 13 1 15 14 9 2
22 3 16 15 13 3 3 1 15 9 15 3 13 10 9 16 15 9 4 13 10 0 2
25 15 9 7 15 13 13 10 3 0 0 9 1 15 9 1 0 9 1 1 0 9 7 9 13 2
18 15 3 13 11 1 11 7 15 13 10 9 7 0 1 15 7 0 2
22 15 13 0 2 0 2 0 2 0 7 3 10 0 0 9 15 3 13 1 15 9 2
10 15 4 13 15 9 3 5 3 0 2
2 0 9
12 15 4 13 9 9 13 9 9 1 15 9 2
12 15 13 15 2 3 14 3 13 1 10 9 2
12 11 11 7 10 9 13 9 1 9 1 9 2
8 15 13 1 14 13 15 9 2
29 3 15 4 13 0 9 2 7 15 4 13 15 16 1 15 9 9 15 4 4 13 10 0 1 11 11 11 11 2
15 15 4 13 3 12 9 7 10 12 9 15 4 13 0 2
15 15 4 13 1 15 9 7 2 10 9 13 3 14 0 2
24 15 13 11 1 0 0 9 7 1 10 9 10 11 13 3 3 13 1 9 7 3 0 2 5
8 15 13 15 13 15 9 0 2
16 15 4 13 14 13 15 12 0 9 1 0 0 9 7 13 2
16 15 13 15 1 10 9 7 15 13 15 3 15 13 15 9 2
7 15 13 3 0 7 0 2
29 6 4 14 13 10 9 9 16 15 4 14 13 14 2 13 2 13 9 7 10 0 9 1 10 9 1 15 9 2
27 15 4 13 15 10 0 9 1 10 9 7 1 10 9 1 15 9 15 4 13 10 9 2 15 13 15 2
12 15 4 13 11 13 10 0 9 13 15 9 2
32 15 4 13 15 14 13 3 10 9 3 16 15 13 15 9 16 3 15 4 13 15 1 3 10 9 7 10 9 10 12 9 2
7 0 1 0 1 10 9 2
27 13 13 12 2 9 9 2 15 13 3 3 3 7 4 14 13 10 3 0 9 16 10 2 9 2 13 2
11 10 9 13 10 0 9 7 9 14 9 2
20 3 0 9 9 9 9 1 9 10 15 3 4 14 13 1 10 9 1 9 2
18 15 13 3 3 0 7 15 4 14 13 10 0 9 13 10 0 9 2
12 15 13 10 10 9 16 15 13 15 0 9 2
18 3 3 15 4 3 13 10 9 1 3 3 15 13 3 14 13 15 2
6 0 9 2 9 2 11
6 0 9 1 0 9 2
16 15 13 15 0 11 9 9 7 10 15 13 14 13 13 6 2
15 9 1 9 2 0 0 9 9 2 9 2 9 9 8 2
11 15 13 15 13 10 0 9 1 9 11 2
9 9 2 0 2 0 7 0 9 2
14 15 4 13 15 1 10 9 9 7 9 9 7 9 11
6 0 9 0 9 0 9
8 15 13 14 13 9 0 3 2
4 10 9 13 2
19 13 15 9 11 1 15 7 15 13 10 13 9 9 7 13 15 13 0 2
11 15 3 13 10 9 9 9 2 0 3 2
11 15 13 10 9 9 9 7 15 13 0 2
20 15 3 13 10 11 9 10 13 0 2 3 10 9 13 12 1 1 12 9 2
5 4 14 13 3 2
15 15 13 14 13 15 9 13 11 2 1 11 12 13 0 2
34 15 13 14 0 1 10 9 15 13 2 3 0 2 0 9 2 7 1 10 9 1 12 2 15 13 10 9 1 10 9 1 10 9 2
26 15 3 13 10 9 2 7 15 13 15 9 3 0 2 12 1 15 0 9 13 16 15 4 13 0 2
3 10 9 2
30 15 13 3 10 9 1 0 9 1 9 14 3 10 9 1 0 9 7 15 13 14 13 10 0 9 3 1 11 11 2
15 0 2 0 2 0 3 13 10 0 1 10 9 7 9 2
14 3 0 2 3 0 2 7 3 10 9 1 11 11 2
8 3 4 10 9 13 1 9 2
12 10 9 13 10 9 9 7 15 13 14 15 2
3 0 0 9
17 15 9 7 15 13 1 10 11 0 9 2 7 15 9 13 0 2
13 9 15 13 4 13 1 9 2 7 4 13 3 2
16 10 9 2 13 9 2 7 9 9 13 10 0 15 3 13 2
17 3 10 9 13 2 7 15 13 9 3 10 0 9 15 3 13 2
13 15 4 13 15 1 1 2 15 13 0 10 9 2
5 0 0 9 3 2
11 15 13 10 0 0 9 15 4 3 13 2
21 10 10 9 13 0 2 7 1 10 0 9 1 9 7 10 9 2 15 13 0 2
11 10 9 13 3 13 3 3 9 7 0 2
18 10 9 15 13 2 11 2 10 9 2 4 3 13 15 9 7 15 2
15 3 2 15 13 3 9 0 2 7 15 13 15 1 9 2
2 9 9
5 11 11 13 0 2
14 15 13 11 7 11 13 3 14 13 15 9 9 13 2
6 10 9 13 3 0 2
18 11 13 3 1 12 9 16 15 13 1 10 12 1 12 0 11 9 2
22 16 15 13 9 14 13 15 1 1 15 9 9 2 15 3 4 13 11 11 7 11 2
5 3 10 0 9 2
7 15 9 7 15 13 15 2
2 15 13
4 13 3 3 2
11 13 14 13 10 11 11 7 10 11 11 2
19 16 13 3 7 3 1 10 9 2 15 4 13 1 9 2 7 15 13 2
10 9 9 13 2 9 9 13 3 0 2
34 15 13 12 9 1 11 11 2 7 15 13 12 9 3 1 11 11 1 11 2 13 1 10 9 2 11 2 7 4 3 13 9 1 2
3 0 7 0
28 11 1 11 11 4 3 13 10 0 9 9 2 1 15 9 7 9 1 10 9 1 15 9 9 7 9 9 2
20 15 9 7 9 13 13 10 9 1 10 9 9 2 13 9 1 10 9 9 2
15 16 15 4 13 11 15 4 14 13 14 13 1 9 0 2
12 15 3 4 13 15 9 1 9 1 15 9 2
33 15 13 1 3 12 7 15 13 1 12 7 13 14 13 10 9 7 15 13 3 1 10 9 3 15 4 13 13 3 16 15 13 2
24 13 10 9 9 10 13 0 2 9 1 9 10 13 0 7 0 7 9 9 10 13 3 0 2
11 3 13 14 13 3 7 13 10 9 3 2
11 11 13 3 0 7 13 3 10 9 13 2
3 0 9 3
17 1 10 0 0 11 15 4 13 15 16 15 13 14 0 0 9 2
10 3 2 15 3 13 10 9 10 9 2
10 3 10 9 2 9 9 2 7 9 2
4 9 13 0 2
7 15 0 9 13 10 9 2
13 15 13 14 13 0 2 3 4 15 9 13 15 2
7 9 4 14 13 0 5 2
6 2 9 2 3 13 2
5 15 13 10 9 2
4 13 15 13 15
20 15 13 3 0 0 0 9 14 13 1 11 2 4 14 2 13 15 9 3 2
6 15 13 10 9 9 2
15 10 9 13 0 7 10 9 4 14 13 0 2 3 3 2
9 1 9 15 9 13 1 15 9 2
13 3 15 13 10 0 9 7 15 9 3 13 0 2
13 9 13 0 7 0 2 15 13 1 10 0 9 2
7 15 4 14 13 10 9 2
2 9 9
12 15 9 4 13 10 0 9 3 10 9 13 2
15 11 11 13 10 9 15 13 7 13 10 9 3 7 3 2
17 15 3 13 15 0 9 14 13 16 15 13 9 0 10 13 9 2
14 15 13 10 0 9 14 13 16 9 13 1 15 9 2
19 3 10 0 9 13 3 2 15 4 14 13 14 13 11 1 11 11 11 2
3 0 0 9
14 10 0 9 13 0 7 13 15 16 13 9 9 9 2
32 1 15 9 5 12 9 2 0 9 3 1 9 2 1 10 9 1 11 13 9 3 2 7 9 15 13 5 12 7 0 9 2
11 15 13 15 1 15 2 3 0 11 14 2
20 3 9 13 10 9 2 0 7 0 16 11 11 0 9 2 13 15 9 9 9
5 0 9 1 0 9
27 11 11 13 3 0 1 15 9 2 7 11 11 13 10 9 14 13 15 13 10 0 9 15 4 13 1 2
23 15 3 13 10 12 2 1 2 12 9 3 1 10 9 15 4 13 1 0 9 7 9 2
26 16 15 13 15 4 14 13 10 9 1 10 9 9 3 2 16 15 13 15 4 3 13 10 9 3 2
45 13 15 9 1 10 0 9 7 4 3 13 1 15 9 2 13 10 9 9 3 16 9 4 13 14 13 9 2 7 10 0 9 1 15 9 2 1 11 2 11 2 13 16 13 2
18 10 9 15 13 3 16 13 7 13 1 10 9 7 1 10 0 9 2
10 4 3 13 1 9 13 0 9 9 2
4 11 2 11 2
5 15 13 15 9 2
18 11 11 13 10 0 9 1 10 9 1 15 9 9 15 13 1 3 2
22 16 15 13 0 16 13 1 1 10 0 0 9 3 15 4 13 10 0 9 14 13 2
36 15 13 10 3 0 9 15 4 3 13 1 2 16 15 13 14 13 1 15 9 4 14 13 0 3 15 13 3 0 13 1 11 11 4 13 2
2 0 2
5 10 9 13 0 2
22 15 13 0 14 13 2 7 10 0 9 13 0 2 3 0 16 13 1 1 10 9 2
5 10 9 13 0 2
16 15 13 1 10 13 9 1 15 9 2 7 4 14 13 15 2
25 3 2 10 9 4 14 13 1 9 9 2 7 9 2 1 11 14 9 2 10 9 13 0 9 2
10 10 9 9 2 13 10 9 1 15 2
27 15 13 9 1 10 9 7 11 11 13 3 7 9 13 0 3 15 13 10 13 1 9 1 2 5 12 2
11 13 11 2 12 9 7 9 9 7 9 2
31 15 13 3 0 1 10 9 9 7 3 3 0 1 10 9 9 2 14 13 9 9 9 7 9 1 10 9 1 10 9 2
14 15 13 3 0 7 4 3 13 3 7 13 1 3 2
12 13 1 10 11 11 0 9 7 0 11 9 2
12 3 15 13 9 2 9 7 9 15 13 15 2
20 0 9 2 9 9 1 11 11 7 15 13 10 9 7 9 14 13 15 1 2
17 3 15 13 1 11 15 4 13 10 0 9 10 13 7 13 3 2
18 16 15 9 13 10 9 7 15 3 13 15 13 7 13 9 13 0 2
3 11 11 8
6 0 9 1 10 0 9
27 15 3 13 3 7 4 13 0 1 10 0 9 2 15 13 10 0 12 7 15 4 4 3 13 1 15 2
35 10 9 13 3 3 0 2 10 0 9 12 15 13 13 1 10 11 9 7 15 3 13 14 4 13 10 0 3 2 7 15 13 3 0 2
15 15 9 9 9 13 12 1 10 0 9 15 4 3 13 2
3 0 9 2
8 3 0 9 1 10 9 9 2
11 15 13 3 0 1 10 9 7 1 9 2
21 15 13 3 1 15 16 15 13 0 9 2 16 15 13 15 9 3 3 3 13 2
16 3 10 9 4 13 3 16 13 3 0 1 9 13 9 13 2
10 15 4 3 13 9 1 11 11 3 2
15 13 11 15 13 9 1 11 9 14 13 1 1 10 9 2
5 15 13 10 0 9
12 15 4 13 3 3 7 10 9 13 3 0 2
17 15 13 10 0 9 1 9 14 13 1 7 15 9 13 3 0 2
40 15 13 13 3 16 15 4 3 13 3 3 2 15 4 4 13 9 14 13 10 9 1 0 9 7 15 4 3 13 1 10 0 7 1 15 10 0 13 3 2
11 15 13 15 14 13 7 13 15 0 9 2
52 11 11 7 11 13 3 0 9 2 7 10 9 15 13 1 15 9 2 10 0 0 9 13 3 2 7 9 7 9 13 3 1 10 9 2 16 7 3 15 13 15 1 3 1 9 13 3 10 9 1 9 2
16 10 0 9 2 16 15 13 0 1 3 10 0 9 1 9 2
16 13 15 10 9 16 13 10 9 2 14 13 16 15 13 15 2
11 15 4 14 13 14 13 0 16 13 9 2
27 13 3 9 2 15 4 13 14 13 1 12 0 11 9 2 3 15 13 14 9 2 13 10 9 1 9 2
4 10 9 13 2
10 13 15 13 3 0 1 12 9 9 2
7 15 13 10 0 9 3 2
25 4 14 13 9 2 3 13 12 9 3 3 1 11 11 2 15 3 4 13 14 13 15 9 3 2
6 13 3 10 9 9 2
18 15 13 14 10 0 9 9 9 2 0 1 10 9 11 13 1 11 2
16 3 2 16 15 13 10 9 7 9 2 6 2 15 13 0 2
12 16 15 13 10 9 0 9 2 15 13 0 2
17 16 15 13 10 9 2 6 2 10 13 14 10 0 1 11 11 2
18 3 0 7 16 15 4 13 10 11 11 9 9 2 10 13 3 15 2
1 11
9 0 9 14 13 1 10 11 9 2
32 10 9 13 0 2 0 9 1 9 3 3 2 7 1 0 10 9 13 0 2 10 9 3 13 10 0 9 1 10 9 3 2
15 13 1 1 3 0 9 7 3 4 14 13 1 10 9 2
15 7 10 9 13 0 9 10 15 4 13 1 10 0 9 2
16 16 15 13 10 9 9 9 2 15 13 10 0 9 14 13 2
3 0 9 7
17 15 13 1 10 11 11 1 0 12 7 15 4 13 10 13 9 2
12 15 13 14 13 1 11 7 15 13 10 9 2
19 10 9 2 11 2 13 3 3 0 3 15 13 10 9 0 1 0 9 2
16 15 13 3 0 7 15 4 3 13 3 1 10 9 7 9 2
19 7 15 13 10 0 9 7 0 9 1 10 9 10 13 10 0 13 9 2
9 0 9 2 9 2 13 10 0 9
22 15 4 13 10 9 1 0 9 2 13 9 1 9 2 13 9 9 2 7 9 9 2
11 15 13 10 0 9 3 7 0 9 9 2
22 12 9 13 10 9 0 2 7 15 13 10 9 3 3 16 15 9 14 9 13 0 2
19 7 15 13 3 0 14 13 15 1 10 9 2 9 2 7 15 13 0 2
5 3 2 0 9 2
7 10 0 9 13 10 9 2
5 10 0 9 3 2
22 10 9 0 2 3 15 4 14 13 3 3 2 7 15 13 3 10 9 3 15 13 2
8 10 9 13 0 15 15 13 2
18 15 4 13 15 13 3 1 1 9 16 15 4 14 13 10 9 9 2
29 15 4 13 10 9 13 14 13 15 9 1 1 10 9 2 16 15 4 13 10 9 3 14 13 10 9 3 3 2
7 3 0 9 2 3 0 9
31 15 15 13 3 1 10 9 2 3 1 10 9 2 13 16 13 3 13 15 13 16 15 13 1 10 0 9 3 1 11 2
39 10 9 13 3 0 2 15 13 0 9 1 10 0 9 2 7 10 9 14 13 3 1 10 9 2 3 1 10 9 16 15 13 3 10 9 2 13 0 2
11 12 1 15 0 12 9 14 13 1 11 2
1 0
23 10 9 13 0 1 10 11 11 11 2 3 15 13 15 4 13 5 13 1 10 0 9 2
17 10 9 13 0 3 3 2 7 3 0 13 10 9 9 7 9 2
15 4 14 3 13 15 13 16 3 0 15 13 14 13 3 2
31 15 4 13 3 12 9 16 15 3 13 2 7 10 9 4 13 0 10 9 2 10 9 3 13 3 1 3 0 7 0 2
12 9 12 9 12 9 12 9 12 2 11 12 2
12 13 10 0 0 9 1 10 9 1 12 9 2
4 9 13 0 2
4 9 13 0 2
4 9 13 0 2
37 15 4 13 10 9 1 10 9 3 15 13 10 9 10 13 3 0 7 10 9 13 0 7 16 15 13 1 9 3 2 15 4 3 13 10 9 2
8 10 0 9 1 10 0 9 2
9 9 1 2 0 9 2 13 3 2
3 0 9 2
3 3 0 2
29 15 13 15 2 13 15 9 1 10 9 15 13 1 15 9 2 7 13 15 1 10 9 10 15 13 1 0 9 2
11 13 7 4 13 1 9 1 10 0 9 2
11 15 13 3 0 1 10 9 1 11 11 2
21 15 13 0 2 13 0 9 1 10 9 2 7 13 10 0 9 16 13 10 9 2
11 15 3 13 15 1 10 1 15 9 2 2
14 0 9 2 13 13 1 15 9 16 13 1 10 9 2
16 15 13 10 12 9 0 0 9 0 9 1 10 11 11 11 2
21 10 9 13 3 0 16 13 10 0 9 1 15 7 10 9 15 9 13 13 0 2
20 16 15 13 1 10 9 1 10 0 9 9 4 14 13 14 13 1 10 9 2
16 15 9 13 10 0 9 7 4 13 10 0 9 1 15 9 2
5 9 0 2 9 0
23 10 9 2 13 1 10 9 1 15 9 14 9 7 9 13 1 13 14 13 15 9 9 2
12 13 1 9 2 9 2 9 9 3 13 15 2
11 3 13 3 1 15 16 15 13 15 9 2
14 13 14 13 10 10 9 9 14 9 15 14 13 9 2
12 3 12 9 2 3 0 13 1 9 15 13 2
12 9 13 0 2 7 9 13 10 9 1 15 2
12 11 11 15 13 10 0 9 15 4 3 13 2
10 15 13 0 2 0 2 0 7 0 2
38 15 13 15 13 15 1 15 9 3 3 1 15 9 2 3 15 9 4 4 13 10 9 0 16 15 13 3 2 3 15 13 0 15 13 15 9 3 2
6 3 16 15 13 0 2
9 13 15 16 13 14 13 15 9 2
13 15 13 0 1 15 9 7 15 13 1 15 9 2
2 9 9
11 15 13 15 9 3 1 10 0 9 9 2
26 15 13 15 13 15 1 10 0 9 2 7 13 14 13 16 15 9 4 14 13 16 15 13 10 9 2
21 12 9 3 2 15 13 15 9 1 10 9 7 15 13 10 9 9 1 13 9 2
23 16 15 13 10 9 1 9 2 4 13 1 2 7 9 9 2 15 13 10 9 1 15 2
7 16 14 2 13 3 3 2
2 0 9
19 3 16 15 4 3 13 11 11 7 15 13 1 0 9 16 15 13 0 2
34 15 13 7 13 1 10 9 1 9 9 7 10 9 7 9 15 13 10 9 13 14 13 15 2 7 3 3 13 15 10 0 9 9 2
17 15 13 15 14 13 1 10 9 7 3 15 4 13 15 10 9 2
8 10 9 1 0 9 13 15 2
11 15 4 14 13 14 13 15 9 1 15 2
4 0 9 9 2
7 3 3 15 13 1 11 2
2 11 2
4 6 2 11 2
4 3 1 11 2
3 3 11 2
18 7 10 0 9 1 10 12 2 9 9 13 10 0 7 3 0 9 2
24 10 0 7 0 2 13 9 13 1 0 9 1 10 0 9 1 10 9 3 1 10 0 9 2
12 0 9 13 1 9 2 3 3 13 9 9 2
14 10 0 9 14 13 1 9 1 10 9 1 9 9 2
5 0 9 7 0 9
26 9 9 13 1 9 14 9 2 9 4 3 3 13 2 15 13 14 13 12 9 1 10 9 9 2 2
36 7 15 13 3 0 14 13 16 10 11 11 14 9 13 0 2 1 10 0 9 13 1 0 9 9 2 10 9 13 12 5 12 5 0 2 2
15 10 9 13 3 0 2 0 2 0 7 0 16 13 0 2
4 4 3 13 2
2 3 0
23 10 9 1 9 2 13 1 10 9 1 15 9 2 13 15 10 0 0 9 15 4 13 2
42 13 15 1 9 1 10 9 15 13 3 2 0 1 15 3 0 16 15 13 2 1 10 9 1 0 9 1 9 2 16 15 13 2 2 2 2 3 3 16 15 4 2
23 16 15 4 13 15 2 13 0 7 13 0 14 13 2 16 15 4 13 3 3 15 4 2
7 0 9 2 0 9 9 2
17 13 1 10 11 11 10 0 9 1 9 7 9 2 9 13 0 2
20 13 14 13 1 9 16 10 9 2 9 13 2 15 13 0 15 13 15 9 2
13 3 2 16 15 4 13 2 10 9 4 13 0 2
11 9 13 0 2 9 0 2 7 9 0 2
12 15 13 10 0 9 9 10 10 9 3 13 2
11 13 1 10 11 11 2 15 4 13 0 2
13 15 4 13 10 0 9 16 15 4 13 1 11 2
31 7 15 9 7 15 3 13 3 13 15 4 13 0 9 2 13 9 1 9 2 2 7 15 13 1 14 13 10 0 9 2
20 7 2 15 4 13 2 15 13 12 1 15 0 9 14 13 1 10 1 11 2
2 0 2
25 4 14 13 10 0 9 9 13 15 2 15 13 10 0 7 0 9 2 12 9 3 2 3 3 2
6 0 9 2 0 9 9
14 15 3 13 10 9 9 9 1 15 9 1 11 14 2
29 15 13 12 9 1 10 9 2 7 9 13 3 1 10 9 0 1 3 3 10 9 2 7 10 0 9 3 3 2
24 10 9 13 0 14 13 1 1 10 9 9 2 7 10 9 1 10 9 7 9 9 13 0 2
18 15 3 13 11 14 1 9 13 10 0 9 1 9 2 9 7 9 2
3 0 9 2
12 15 13 1 10 9 16 10 9 13 15 9 2
18 15 4 13 1 10 0 11 11 11 9 2 1 11 1 1 11 11 2
9 10 9 4 13 1 9 7 9 2
10 10 0 9 13 13 0 7 3 0 2
9 10 9 13 15 11 13 3 1 2
14 3 2 15 13 10 9 0 9 7 10 4 13 0 2
17 15 9 7 9 13 0 7 15 4 3 4 13 1 15 9 3 2
5 0 9 2 0 9
16 15 4 13 14 13 10 9 10 13 11 11 11 13 0 9 2
19 15 13 15 14 13 16 10 9 3 13 9 13 9 1 3 2 0 11 2
12 10 9 7 9 15 13 10 9 13 0 9 2
33 15 4 13 0 9 1 15 7 15 4 3 13 3 0 1 15 16 15 13 1 0 9 1 9 1 10 0 9 1 15 9 9 2
5 15 13 15 3 2
13 4 14 3 13 3 2 14 3 16 15 9 13 2
14 15 9 13 14 13 1 3 2 9 13 0 7 0 2
11 15 13 3 0 1 15 9 7 15 9 2
21 15 4 14 13 10 9 9 7 3 16 15 9 13 2 15 4 14 13 15 3 2
6 4 14 3 13 3 2
14 15 13 11 11 11 1 10 0 9 1 10 0 9 2
8 7 15 13 14 13 10 9 2
7 4 14 13 3 2 13 15
1 0
21 15 4 4 13 15 9 3 1 12 9 3 7 13 3 14 13 12 9 13 1 2
26 15 13 3 1 12 9 0 9 1 10 9 2 12 9 0 9 1 10 9 2 7 12 1 10 9 2
9 15 9 13 0 7 15 13 0 2
11 10 9 4 4 13 1 11 2 16 15 2
16 15 13 10 0 9 7 15 13 16 10 9 0 13 1 15 2
13 13 8 15 10 9 7 4 14 13 1 10 9 2
6 10 0 11 11 9 2
24 15 3 13 10 11 1 10 0 3 13 9 2 3 2 15 13 14 13 10 9 1 15 9 2
11 15 13 10 9 1 15 0 9 2 11 2
17 15 13 10 9 9 1 10 9 7 13 10 9 4 3 13 3 2
15 15 13 15 14 13 15 7 15 3 13 16 15 13 0 2
8 0 0 9 13 3 0 9 2
14 4 14 13 2 7 15 4 13 3 14 13 15 9 2
1 0
20 10 0 2 15 13 1 11 3 7 13 3 0 1 0 9 9 7 0 9 2
17 15 13 10 9 1 12 7 9 1 15 13 3 0 1 15 9 2
17 11 13 3 1 9 7 13 3 0 9 1 10 9 1 15 9 2
17 15 13 15 0 9 0 7 10 9 9 15 13 14 13 3 13 2
21 16 15 4 13 13 9 1 9 1 15 9 16 15 9 4 3 0 16 15 13 2
2 3 13
22 15 13 3 14 13 15 0 9 1 12 9 1 9 7 13 9 1 9 7 10 9 2
13 10 9 13 0 1 0 7 10 9 13 3 0 2
20 15 9 1 9 7 9 3 13 1 10 0 9 13 15 10 9 15 13 3 2
35 15 4 3 13 3 3 3 1 10 9 7 15 13 0 10 0 9 2 16 10 9 13 13 15 9 2 3 1 10 0 0 9 9 3 2
3 0 2 2
18 15 13 14 13 10 1 10 0 9 15 4 3 13 10 9 16 13 2
13 10 9 13 0 2 0 1 12 9 1 10 0 2
11 15 3 13 10 9 1 12 1 10 9 2
12 15 13 0 9 7 9 7 15 3 13 9 2
11 15 13 11 11 9 7 15 13 14 15 2
9 15 13 9 1 11 11 9 9 2
12 15 13 9 7 15 13 10 0 7 0 9 2
9 15 4 14 13 10 9 1 9 2
19 0 9 3 15 9 13 0 3 0 3 15 13 11 11 11 11 9 9 2
15 15 13 1 15 9 1 10 9 7 13 13 1 10 9 2
17 15 13 3 0 7 13 0 14 13 15 3 15 13 0 1 15 2
22 16 15 13 15 15 13 10 1 15 9 1 10 9 7 3 13 15 10 0 9 3 2
20 15 13 16 16 15 9 9 13 14 4 13 2 15 4 4 13 11 11 11 11
8 15 4 13 0 1 10 9 2
15 11 11 4 13 1 9 16 15 13 0 9 9 1 11 2
18 10 9 9 2 11 11 2 13 10 0 9 9 1 15 3 13 11 2
19 9 13 10 0 9 7 3 10 9 13 16 15 4 13 1 9 1 9 2
15 10 9 13 0 2 13 3 3 7 10 9 14 13 1 2
20 15 13 15 9 7 15 4 14 13 14 13 15 14 13 0 9 4 13 0 2
9 0 9 15 3 13 13 10 9 2
28 0 9 2 3 3 4 15 13 10 0 9 15 13 8 1 12 9 7 10 9 9 3 13 15 3 1 9 2
5 3 0 7 0 2
19 15 3 13 10 9 16 15 4 14 13 14 13 1 9 7 13 0 9 2
23 15 4 3 13 12 9 1 10 9 2 10 0 9 13 1 11 7 10 9 13 1 11 2
11 10 13 0 9 9 15 13 15 9 3 2
18 10 9 4 13 10 0 9 16 13 9 1 10 0 9 1 15 9 2
38 15 3 3 13 14 13 3 1 10 3 9 9 2 7 3 13 10 0 9 0 9 3 13 15 2 2 10 9 9 13 14 3 9 2 2 1 9 2
39 9 15 13 1 11 11 7 15 13 12 9 1 9 1 15 1 9 2 7 15 13 3 1 1 3 3 3 2 3 13 9 14 13 10 9 1 15 9 2
4 3 0 7 0
22 1 0 2 9 9 9 2 15 9 7 15 13 11 11 1 11 11 11 2 3 0 2
16 15 13 1 15 1 1 10 9 2 13 15 13 15 0 9 2
26 11 14 9 1 10 9 7 9 1 15 9 9 2 13 15 13 0 1 15 9 14 13 3 15 13 2
16 15 4 3 13 11 1 9 13 1 10 9 1 10 11 11 2
9 15 13 15 9 2 9 7 9 2
2 0 9
33 3 2 10 0 9 3 4 3 13 1 11 14 2 7 15 4 13 16 11 3 13 5 12 1 10 9 10 13 3 3 9 9 2
19 15 4 4 13 1 11 1 12 9 3 3 16 15 4 13 9 1 9 2
16 15 13 0 9 7 15 3 13 15 9 14 13 15 13 0 2
26 10 1 10 0 9 10 13 3 13 10 9 8 0 2 7 16 15 13 1 11 2 15 4 13 0 2
2 6 2
16 13 10 0 2 3 13 2 9 9 2 10 0 9 1 15 2
8 13 10 9 2 15 13 0 2
12 13 10 9 1 7 13 15 0 1 0 9 2
2 6 2
24 15 13 10 9 7 10 9 13 2 7 13 16 15 13 0 2 7 13 15 13 14 15 9 2
8 15 3 13 14 13 10 9 2
10 15 13 15 9 2 7 13 14 3 2
10 0 9 13 0 9 13 1 10 9 2
7 15 4 3 13 3 3 3
12 1 0 0 9 2 15 13 10 9 14 13 2
24 15 13 14 13 1 9 1 11 11 7 11 11 1 11 2 11 2 9 0 7 3 3 0 2
16 3 2 15 4 14 13 0 9 0 16 15 13 1 10 9 2
11 10 0 9 15 4 13 1 10 0 9 2
20 15 4 14 13 1 11 11 11 3 2 7 9 13 3 0 7 10 9 0 2
16 3 15 13 14 13 1 10 9 14 13 10 9 2 0 9 2
3 0 9 2
11 15 9 13 0 1 11 11 7 11 11 2
7 11 11 13 9 1 0 2
15 15 13 15 13 16 15 13 10 3 0 9 1 10 9 2
7 11 13 15 13 3 0 2
11 13 15 1 0 9 7 13 0 9 13 2
13 13 1 10 9 15 4 13 14 13 0 7 0 2
7 9 13 9 1 10 9 2
23 15 4 13 9 14 13 13 11 11 7 11 11 14 13 10 10 0 9 15 13 14 13 2
30 11 13 10 0 7 0 9 2 15 13 10 0 9 7 9 1 15 9 14 9 7 10 9 15 13 15 9 14 13 2
23 3 2 15 13 9 3 3 2 15 9 13 0 2 7 15 4 14 13 15 9 1 9 2
6 11 13 0 14 13 2
34 1 3 12 5 12 13 9 2 15 13 3 3 0 16 13 1 0 9 1 11 9 3 14 9 7 4 3 13 15 0 9 1 9 2
2 2 11
6 15 13 15 0 9 2
16 15 4 13 14 13 15 1 10 9 9 15 13 1 15 9 2
22 9 4 13 1 10 0 9 7 9 4 13 7 13 1 10 9 3 10 9 13 0 2
14 15 3 13 10 9 3 11 13 1 10 9 10 9 2
18 7 3 10 9 13 0 10 9 4 13 1 7 13 1 10 0 9 2
10 15 4 14 13 14 13 11 11 3 2
11 15 4 3 13 15 1 10 1 15 9 2
1 6
83 15 3 13 10 9 10 9 15 13 10 0 9 13 1 7 15 13 3 0 7 15 13 6 3 0 7 3 15 13 10 0 9 10 13 3 0 7 15 13 6 3 0 15 4 13 10 9 2 7 3 15 13 10 9 15 3 13 3 0 7 15 3 13 15 0 9 15 13 3 0 1 10 0 9 9 15 13 15 4 13 14 13 2
12 3 15 13 3 1 15 9 7 13 9 7 9
3 3 0 2
14 15 3 13 3 1 11 9 7 3 13 10 9 3 2
32 15 9 1 9 13 15 1 10 0 0 9 9 1 9 2 15 13 3 0 15 3 13 14 13 7 13 15 1 1 8 15 2
6 15 9 9 13 0 2
11 15 9 13 0 1 9 15 4 3 13 2
4 3 1 11 2
22 15 4 3 13 10 9 1 9 13 1 10 0 9 2 0 9 2 7 0 9 9 2
6 13 15 11 11 11 2
22 15 13 12 1 10 0 9 15 4 13 2 15 13 15 9 0 7 13 1 10 11 2
28 3 16 15 3 13 15 10 9 15 13 7 4 14 13 2 15 13 1 10 13 10 9 1 1 10 9 9 2
17 10 0 9 13 10 9 13 16 15 4 13 10 12 9 9 9 2
8 0 9 13 1 10 0 9 2
7 10 0 9 13 10 9 2
19 3 1 15 2 13 10 9 2 1 10 9 11 9 2 15 13 10 9 2
4 0 9 1 11
27 15 13 3 1 12 9 3 10 9 13 10 0 0 5 10 9 13 3 0 7 0 2 7 1 0 9 2
19 15 3 13 10 9 1 11 2 3 10 9 11 13 3 3 0 7 0 2
6 10 9 9 13 0 2
28 10 0 9 10 15 13 1 12 9 16 13 3 13 16 10 9 13 3 0 2 3 15 4 13 15 9 9 2
8 15 4 13 10 9 1 9 2
6 15 3 13 13 3 2
5 10 0 9 3 2
7 15 4 3 13 0 9 2
13 15 9 13 1 7 9 13 15 9 1 11 11 2
15 15 13 15 1 7 13 15 3 3 7 13 1 10 9 2
7 9 13 0 7 3 0 2
19 10 9 9 3 13 15 10 9 3 7 13 15 1 3 15 9 13 0 2
16 10 9 13 15 1 1 9 7 13 1 10 9 1 15 9 2
8 15 13 10 9 10 9 5 2
11 15 4 3 4 13 15 9 3 1 9 2
4 9 1 11 2
3 4 13 2
2 10 5
6 10 9 13 10 0 2
13 15 13 9 3 7 3 15 4 14 13 13 15 2
7 0 11 2 7 0 9 2
8 9 1 3 13 14 13 15 2
14 15 9 9 13 1 1 10 9 7 9 13 3 0 2
10 15 13 3 3 3 12 9 10 9 2
18 15 13 0 9 9 0 9 1 10 0 9 7 3 13 10 9 9 2
3 9 5 2
8 11 7 11 15 13 15 11 2
5 2 10 9 2 5
4 0 2 0 9
12 10 12 2 9 9 1 12 13 1 1 9 2
20 15 13 10 9 1 9 10 9 1 9 3 7 9 13 7 0 7 3 0 2
17 10 9 13 14 13 3 0 2 9 9 2 0 9 2 0 9 2
8 10 9 4 14 13 1 9 2
36 15 13 10 0 9 3 0 9 4 13 1 10 0 9 2 1 1 0 0 9 2 2 7 16 15 13 0 1 15 2 10 9 13 3 0 2
4 13 10 9 2
7 10 0 0 9 1 10 9
6 10 0 9 1 11 2
6 4 15 13 10 9 2
12 3 16 15 13 1 10 9 16 15 13 11 2
14 10 9 13 10 0 7 3 15 13 15 1 10 9 2
14 10 9 9 9 2 9 9 2 13 14 14 4 13 2
17 9 9 13 0 7 3 15 13 10 9 9 10 13 3 1 9 2
25 13 0 9 1 10 9 2 10 0 9 15 13 3 15 4 13 16 13 10 0 3 1 10 9 2
13 11 11 13 12 1 10 0 9 9 15 4 13 2
21 10 0 9 15 13 15 15 13 1 9 7 13 9 1 15 1 10 9 15 13 2
20 10 9 9 10 13 1 11 11 13 3 0 7 0 7 13 10 9 15 13 2
19 15 4 13 9 1 15 10 0 9 7 15 13 3 3 0 1 10 9 2
26 16 15 4 13 1 9 9 10 4 13 15 10 0 13 9 9 2 3 11 11 13 10 9 1 15 2
6 10 3 0 0 9 2
15 1 10 3 0 0 9 2 15 3 13 11 11 11 11 2
17 15 13 0 2 0 2 7 13 0 9 7 9 16 13 15 9 2
39 3 3 13 15 9 7 15 3 0 2 7 15 3 13 10 9 9 9 13 3 1 10 9 9 10 15 3 13 2 16 7 16 11 11 11 13 15 9 2
21 13 1 10 9 9 2 10 9 9 13 16 10 9 1 15 9 13 2 0 2 2
7 10 0 9 1 11 11 2
6 15 13 11 14 11 2
17 1 10 9 10 0 9 14 13 10 0 0 9 7 10 9 9 2
16 11 14 4 13 10 11 11 9 1 12 9 7 1 0 9 2
19 9 13 7 13 13 0 10 9 13 0 7 10 9 9 2 13 1 9 2
18 15 3 13 13 1 10 9 1 15 0 0 9 9 2 3 10 0 2
18 16 15 4 13 1 11 11 2 9 13 15 13 1 15 9 9 3 2
3 11 11 11
36 0 9 1 11 11 13 12 10 0 9 9 2 15 4 13 1 15 1 15 9 2 15 13 3 0 15 13 15 1 15 9 9 2 7 9 2
19 15 13 3 0 2 0 2 13 10 9 1 9 2 7 3 1 15 9 2
41 11 12 1 9 13 0 2 15 13 10 0 9 2 7 13 1 9 2 15 4 3 13 13 15 7 13 15 1 0 9 15 4 1 1 10 0 9 15 13 15 2
4 0 9 9 2
9 0 9 2 0 9 2 0 9 2
16 15 13 10 9 1 0 9 3 13 15 0 13 9 9 12 2
14 16 13 1 12 0 9 15 3 13 11 1 11 11 2
32 3 3 13 15 10 0 9 7 15 9 7 9 13 1 15 9 10 9 15 13 2 13 15 13 10 0 9 15 4 3 13 2
13 7 15 13 1 15 0 9 7 11 13 10 9 2
12 13 16 15 13 10 9 1 9 1 10 9 2
4 0 10 9 2
5 15 0 9 1 11
23 15 4 4 13 1 10 11 2 11 1 1 12 9 1 9 9 7 3 13 10 11 3 2
6 15 13 15 12 9 2
11 15 4 14 13 15 13 10 12 9 9 2
21 15 4 13 3 13 10 0 9 1 11 2 10 9 13 9 10 15 4 13 1 2
25 15 13 10 9 1 11 7 9 2 10 13 15 13 1 10 12 9 9 1 10 9 1 10 9 2
12 15 13 10 9 1 9 7 15 13 3 0 2
5 3 1 11 2 11
18 16 3 1 11 6 13 10 9 14 13 11 11 11 11 7 15 9 2
16 15 13 7 3 4 13 10 0 9 1 11 10 15 4 13 2
12 15 4 3 13 10 9 16 13 10 11 9 2
21 15 4 3 13 10 9 16 13 10 0 0 9 2 10 15 4 13 1 9 1 2
27 15 4 8 2 3 13 3 0 1 15 9 7 9 10 15 0 9 13 15 3 15 13 3 1 12 9 2
3 9 3 2
52 15 4 3 13 10 9 14 13 10 9 7 13 10 9 3 2 7 1 10 9 15 4 13 1 1 10 9 1 9 1 10 9 2 15 9 15 13 14 13 11 11 2 15 4 3 14 13 10 9 1 9 2
22 16 10 9 4 13 1 10 0 9 10 9 4 13 3 15 13 10 9 14 4 13 2
27 9 4 4 13 1 1 15 3 1 3 0 15 9 4 4 13 7 15 4 4 13 1 1 15 0 9 2
5 0 9 9 1 11
8 15 13 10 11 1 10 9 2
16 10 9 9 13 3 0 1 10 9 1 10 9 15 13 1 2
15 15 13 3 0 7 0 16 13 10 9 16 13 10 9 2
9 10 9 13 10 3 0 7 0 2
19 15 13 14 13 15 9 9 3 3 16 0 16 15 4 14 13 15 9 2
14 3 2 15 13 3 0 1 10 9 9 7 15 9 2
15 16 15 4 13 14 13 10 9 2 3 13 15 10 9 2
6 15 13 10 0 9 2
13 15 4 13 10 9 1 11 9 7 15 13 0 2
23 15 4 3 13 10 12 9 9 10 15 13 1 13 1 10 9 7 0 9 1 10 9 2
22 6 2 15 13 14 13 2 7 9 13 10 9 9 10 13 10 3 9 13 9 3 2
7 10 9 4 13 10 0 2
17 3 3 16 4 13 1 10 9 9 2 15 4 14 13 15 9 2
9 1 10 9 15 13 1 9 9 2
17 15 13 10 0 9 7 3 0 16 15 13 9 1 10 11 9 2
2 0 9
26 15 13 0 9 1 10 11 9 2 16 9 7 9 13 15 16 15 4 3 13 10 9 1 10 11 2
21 11 11 13 3 3 0 1 10 11 2 7 3 13 0 14 3 13 9 1 15 2
20 15 13 3 0 1 10 9 15 13 2 13 15 9 1 0 9 14 13 1 2
17 13 1 10 9 15 13 10 9 1 0 2 11 11 13 10 0 2
13 15 3 13 10 9 10 9 0 9 1 0 9 2
7 15 4 13 15 1 9 2
1 0
12 10 9 13 10 0 12 15 4 3 13 1 2
12 15 13 15 1 12 9 2 7 15 13 0 2
25 15 13 9 3 1 10 9 2 9 3 13 1 10 9 2 7 10 0 9 1 10 9 13 0 2
37 10 9 7 10 9 13 0 2 15 4 14 13 1 10 9 2 7 15 13 1 0 9 2 15 13 9 2 16 10 9 13 1 10 9 14 2 2
20 10 9 13 0 3 3 2 13 9 10 9 2 7 4 14 13 15 9 3 2
7 0 9 9 7 0 9 2
30 15 13 10 0 9 14 13 15 9 9 2 15 13 14 13 10 0 9 1 9 10 13 1 9 9 14 13 10 9 2
6 15 13 12 9 3 2
22 15 4 14 13 0 14 13 10 9 9 9 1 11 3 10 4 13 0 14 13 15 2
12 2 15 4 13 1 3 3 12 9 3 2 2
29 16 15 13 9 14 13 1 11 16 15 13 1 10 9 9 2 15 4 3 16 15 4 13 10 9 13 3 3 2
13 3 0 1 0 11 11 11 2 3 16 13 0 9
30 16 13 3 1 9 7 13 14 13 9 1 10 11 2 15 4 13 1 10 11 11 11 11 1 10 9 1 0 9 2
35 10 0 9 13 15 14 13 1 9 1 9 1 15 0 9 9 16 16 15 4 13 9 1 12 1 12 7 10 9 9 13 3 15 9 2
24 15 13 3 0 16 3 0 0 9 4 13 3 3 1 12 9 7 15 13 14 13 10 9 2
2 9 5
29 10 9 4 3 13 9 9 0 2 7 16 15 4 13 1 10 0 9 7 13 14 10 9 2 4 14 13 15 2
23 10 0 9 15 13 15 15 4 13 14 13 11 3 15 13 15 15 4 13 1 10 9 2
16 15 13 15 15 13 7 13 10 9 16 15 13 14 10 9 2
25 15 13 14 13 15 15 13 3 15 13 13 15 16 15 13 15 9 13 1 7 15 13 10 9 2
16 3 15 13 14 3 0 1 10 9 1 9 13 1 10 9 2
8 0 7 0 9 15 4 13 3
10 15 9 7 15 13 3 1 9 9 2
16 10 9 1 15 4 3 13 2 3 15 13 15 4 13 15 2
10 0 9 2 10 9 13 0 7 0 2
10 15 10 13 13 14 13 9 15 13 2
35 10 0 9 15 13 0 13 10 9 9 2 15 3 13 1 2 15 13 13 2 15 13 10 13 9 14 13 0 2 15 0 9 13 0 2
19 4 14 13 10 9 1 9 2 1 9 2 13 15 9 7 13 3 3 2
3 8 13 2
22 15 13 14 10 9 1 8 2 7 12 1 15 9 13 11 13 10 9 13 0 9 2
17 15 13 1 15 7 1 0 12 9 15 4 13 15 9 1 11 2
44 16 15 4 13 1 0 9 9 14 13 16 10 9 4 13 0 9 7 14 2 7 15 4 13 16 15 13 0 0 9 1 11 3 11 3 13 10 9 9 1 15 0 9 2
10 10 9 1 9 15 13 13 3 0 2
10 15 4 13 14 13 15 0 9 1 8
5 11 11 1 10 11
4 9 11 11 2
12 15 4 4 13 10 0 11 11 1 10 11 2
14 10 1 15 4 13 0 1 15 0 9 1 10 9 2
10 0 9 2 0 11 9 1 10 9 2
8 0 11 9 9 1 10 9 2
12 0 9 2 9 9 3 2 11 11 2 9 2
7 9 9 9 9 2 9 2
8 3 13 1 11 7 10 9 2
7 9 9 9 9 2 11 2
8 3 13 1 11 7 10 9 2
7 9 9 9 9 2 11 2
8 3 13 1 11 7 10 9 2
3 0 7 0
22 16 15 13 0 0 9 13 3 1 9 1 0 9 2 15 13 14 10 9 1 15 2
19 16 15 13 3 13 0 9 10 13 10 0 0 9 2 15 4 13 11 2
21 9 2 3 10 0 9 7 9 15 4 3 13 2 7 15 4 13 10 9 2 2
20 10 9 13 0 2 10 9 13 9 2 0 2 10 9 4 14 4 13 0 2
23 15 4 13 1 9 1 0 2 9 9 7 15 4 3 3 13 15 9 4 3 3 13 2
6 0 9 2 0 9 2
30 15 4 13 1 10 9 3 2 3 1 10 9 7 3 1 10 9 9 2 7 15 3 13 1 1 15 9 2 11 2
19 15 13 10 9 1 9 0 1 9 9 2 9 9 2 9 9 2 8 2
15 10 9 13 2 15 3 13 0 9 9 1 3 0 9 2
14 15 13 3 0 9 7 9 1 9 16 15 4 13 2
20 10 9 13 10 0 9 7 15 4 13 15 9 1 15 7 10 1 15 9 2
7 0 9 2 10 10 9 2
3 11 13 0
13 11 13 10 3 0 7 0 9 10 15 4 13 2
13 15 13 0 14 13 10 15 13 1 15 1 9 2
18 15 13 0 7 13 3 9 4 14 13 13 1 9 1 15 9 9 2
15 7 10 9 7 9 9 10 15 13 1 15 13 3 0 2
9 15 13 10 9 3 1 15 3 2
8 15 4 3 13 11 1 9 2
6 15 4 13 15 9 2
25 15 4 14 3 13 9 15 13 9 1 1 15 7 15 4 14 3 13 16 15 13 10 9 3 2
3 14 3 0
18 15 9 3 13 10 9 3 1 10 9 15 4 3 13 15 10 9 2
13 15 13 10 0 9 7 15 13 10 9 1 9 2
8 7 3 10 9 10 9 13 2
22 15 13 15 3 7 15 4 14 13 10 9 7 13 15 13 15 9 1 1 15 9 2
23 3 15 4 13 14 13 15 1 0 9 7 13 14 13 15 3 16 3 13 15 10 9 2
5 10 13 3 0 2
16 15 13 1 10 0 9 3 7 15 3 13 15 12 9 3 2
5 11 13 14 3 0
4 3 0 1 9
30 15 4 4 13 15 9 1 10 0 9 3 7 4 13 10 9 7 3 1 1 10 9 10 15 4 13 15 4 13 2
21 10 9 3 13 14 13 3 1 0 7 0 2 7 15 13 0 1 15 9 9 2
22 3 13 10 9 16 15 4 13 15 10 9 1 10 9 2 3 16 15 13 10 9 2
5 15 13 3 0 2
21 15 13 14 13 3 3 16 15 4 1 15 3 16 15 3 13 1 10 9 9 2
9 15 4 14 13 12 9 1 15 2
3 0 9 2
19 13 10 9 14 13 15 13 1 10 9 14 13 9 9 7 13 10 9 2
23 15 13 1 9 15 13 15 13 9 1 9 7 4 14 13 15 0 9 7 13 10 9 2
30 3 15 13 10 9 14 13 2 15 13 15 13 10 9 4 14 13 1 9 7 16 10 0 9 13 3 0 9 3 2
11 3 16 13 15 13 14 13 15 9 3 2
9 3 15 13 10 9 1 10 9 2
8 14 3 13 3 7 13 1 2
9 15 4 3 13 9 1 10 9 2
2 3 2
6 9 9 13 0 7 0
42 15 4 13 14 13 10 9 1 15 9 14 13 10 9 7 10 9 9 0 9 13 11 13 15 10 9 2 7 16 15 13 0 15 9 15 4 4 13 13 15 9 2
30 15 13 9 7 13 1 9 2 6 2 4 15 13 1 9 14 0 9 10 9 4 4 13 1 10 9 14 13 9 2
29 1 10 0 9 9 15 4 13 1 9 13 14 13 10 9 1 10 9 7 3 13 16 15 13 3 1 10 9 2
6 13 3 1 10 9 2
7 10 9 13 10 9 2 9
20 15 13 10 9 3 14 13 10 2 13 9 2 9 13 3 1 11 1 12 2
22 15 13 15 13 2 9 7 9 2 7 13 15 5 12 14 13 10 9 2 13 9 2
22 15 13 3 3 0 7 15 13 15 13 1 1 10 9 16 13 9 1 1 10 9 2
25 10 9 13 1 13 10 9 9 9 9 2 12 9 2 7 10 9 9 9 2 12 9 9 2 2
9 15 13 10 9 15 1 5 12 2
10 15 13 10 9 1 10 9 1 9 2
22 15 9 7 15 13 10 9 1 10 9 16 15 4 14 13 14 13 1 9 1 11 2
11 15 10 0 9 2 10 9 13 10 9 2
7 9 8 15 13 3 0 2
31 9 8 10 9 13 0 7 0 2 1 10 0 9 1 10 0 9 9 2 7 2 3 3 2 9 8 10 9 13 0 2
14 15 13 0 0 9 2 0 9 3 13 7 13 3 2
21 10 9 13 0 7 15 13 3 1 0 1 10 9 1 12 9 1 10 9 9 2
9 13 10 9 2 15 4 13 15 2
9 13 15 16 13 15 13 3 0 2
15 15 13 3 7 13 11 11 3 10 9 3 16 13 9 2
17 15 13 14 13 15 16 15 4 14 13 12 7 4 14 13 12 2
23 15 13 10 0 9 10 15 4 3 13 7 15 13 10 15 9 16 15 4 13 15 3 2
9 15 13 10 9 1 15 1 15 2
17 11 11 2 16 15 13 15 2 13 15 16 13 15 13 3 0 2
19 15 13 0 7 13 16 15 13 0 9 0 1 15 3 16 15 4 3 2
7 15 4 14 13 15 3 2
16 11 1 11 2 9 0 9 1 9 1 9 9 7 9 8 2
29 15 4 13 10 9 7 9 1 11 1 11 1 3 1 12 9 3 7 15 3 13 15 9 9 10 12 9 3 2
30 11 13 10 13 9 1 10 9 7 15 4 4 13 16 15 4 13 14 13 10 15 9 9 1 10 3 9 0 9 2
36 15 4 13 3 0 1 10 9 7 13 2 1 9 15 4 13 1 15 1 10 9 2 9 3 0 9 9 9 13 1 11 7 15 9 11 2
3 15 9 9
25 6 15 9 13 11 7 15 4 13 10 9 1 15 0 9 9 1 11 2 11 7 1 11 11 2
17 15 13 10 13 0 9 9 7 15 13 1 9 1 0 9 9 2
10 15 13 0 2 0 7 13 9 9 2
10 15 9 13 0 2 0 2 7 0 2
13 6 13 15 9 14 13 0 1 15 9 1 8 2
10 15 13 10 13 9 1 0 9 9 2
6 13 15 0 9 3 2
18 15 4 13 9 1 9 15 4 13 1 15 3 1 10 0 9 9 2
3 0 1 9
18 16 15 13 9 7 13 3 10 0 9 9 15 15 4 13 10 9 2
14 15 13 3 5 12 7 1 9 3 12 0 9 9 2
16 15 13 9 7 9 9 1 10 9 7 15 13 15 13 9 2
29 15 13 15 12 9 0 7 15 13 7 13 3 2 3 3 15 4 13 2 13 7 2 13 2 10 9 7 9 2
11 10 9 13 3 3 0 7 0 1 15 2
17 1 10 9 10 13 0 14 13 13 9 2 9 7 3 10 9 2
8 0 2 0 7 9 1 9 2
2 6 2
23 15 4 14 13 0 0 9 1 11 7 10 0 9 15 4 13 1 15 7 15 9 11 2
14 11 13 3 0 14 13 15 16 15 13 14 13 15 2
13 15 4 3 13 3 1 11 3 1 0 9 9 2
25 15 4 13 9 1 15 0 9 1 3 12 9 3 7 15 4 14 13 11 13 1 9 1 15 2
13 15 13 0 2 0 2 7 3 0 1 15 9 2
26 15 4 13 15 10 9 2 15 13 0 10 9 14 13 16 15 9 13 1 0 9 1 11 11 11 2
6 0 9 15 4 3 13
19 15 13 15 13 9 0 14 13 1 10 9 2 7 3 2 15 13 14 2
8 8 2 9 7 9 13 0 2
20 8 2 10 9 3 13 3 1 9 7 13 3 0 1 10 9 16 13 0 2
21 2 1 7 15 7 9 2 8 2 15 4 3 13 3 0 9 13 1 10 9 2
8 8 2 10 9 13 3 0 2
18 10 9 13 14 0 2 3 15 13 0 14 13 15 15 4 13 1 2
15 15 4 13 14 13 15 9 7 9 7 13 10 0 9 2
5 11 13 10 0 2
13 11 13 10 3 13 7 3 0 9 9 1 11 2
11 15 4 4 13 3 1 1 12 9 3 2
18 10 9 13 3 0 7 0 7 10 9 2 11 2 13 10 0 9 2
19 10 9 9 13 0 13 16 10 9 13 0 14 13 7 3 13 1 11 2
33 1 9 2 10 9 13 1 3 0 9 1 10 9 1 11 11 2 10 4 13 3 3 16 0 1 9 13 1 0 9 1 11 2
11 11 13 3 0 7 0 3 1 15 9 2
5 13 3 1 11 2
1 0
24 11 3 13 10 9 1 15 9 3 1 1 15 9 1 11 11 2 7 15 4 14 13 15 2
26 10 9 3 13 12 9 7 2 10 9 13 14 1 1 9 1 10 9 9 7 10 9 10 9 13 2
31 10 9 15 13 13 0 7 15 13 14 3 0 16 15 4 4 13 2 13 16 15 4 13 1 15 9 3 1 15 9 2
7 10 0 9 13 3 0 2
19 5 12 1 10 9 10 13 3 12 0 9 9 7 13 0 1 9 9 2
7 15 4 14 13 3 3 2
6 11 13 1 10 9 2
16 1 10 9 15 13 10 9 2 15 13 15 13 10 9 0 2
12 10 9 13 0 2 7 10 9 13 3 0 2
23 15 3 13 10 12 2 9 9 9 2 10 13 15 9 1 9 7 9 14 13 15 9 2
44 3 2 16 15 13 1 9 2 11 13 10 9 1 7 9 2 9 2 7 9 14 13 3 10 9 2 7 1 12 9 2 13 15 0 9 1 0 2 10 9 9 2 2 2
17 16 15 13 14 0 2 11 4 13 15 10 9 15 4 3 13 2
7 10 9 13 14 0 7 0
11 15 4 13 1 11 11 9 1 12 9 2
8 15 13 10 9 7 10 9 2
14 15 13 10 0 9 7 15 13 0 13 3 1 9 2
6 10 9 9 13 0 2
9 7 10 9 13 3 0 2 3 2
19 6 2 15 3 13 10 0 9 2 7 15 4 13 14 13 3 15 13 2
11 10 0 9 10 15 4 13 13 10 9 2
6 15 13 10 0 9 2
19 15 13 15 13 0 2 7 15 4 14 13 15 1 1 9 2 0 9 2
11 0 1 15 2 15 4 13 13 3 2 5
9 10 9 13 10 9 14 4 13 2
17 10 9 9 4 13 10 10 9 1 9 7 13 1 0 1 0 2
16 10 0 13 2 1 9 9 1 10 9 3 13 1 10 9 2
10 15 4 13 10 9 1 10 10 9 2
18 15 3 13 16 10 9 13 10 9 16 15 4 13 1 1 15 9 2
18 16 15 4 13 7 13 1 10 9 3 15 13 10 0 9 1 15 2
23 3 15 13 14 0 15 14 13 1 10 9 1 9 7 15 0 9 14 13 1 10 9 2
10 15 13 10 0 9 7 3 0 15 2
6 11 2 0 0 11 11
11 15 4 13 10 11 11 12 9 1 12 2
26 1 11 11 2 1 10 9 1 10 11 9 2 2 15 4 13 3 2 10 9 1 0 9 7 9 2
16 15 13 9 3 2 1 9 10 0 9 4 13 1 10 9 2
11 15 13 0 9 1 10 9 1 10 9 2
14 7 3 3 2 15 9 4 14 13 1 10 0 9 2
10 15 4 4 13 0 16 15 4 13 2
12 11 7 11 2 10 9 13 10 9 1 9 2
10 0 2 0 2 0 2 0 7 0 2
6 15 13 14 13 3 2
3 9 9 2
42 3 0 9 2 15 4 13 3 1 9 13 15 4 13 3 1 10 9 9 7 6 2 15 13 10 0 9 1 11 11 9 13 1 10 9 13 9 7 13 10 9 2
37 10 9 9 9 3 13 2 3 2 7 10 9 15 13 14 13 10 0 1 10 9 2 3 1 10 0 1 10 9 13 15 15 4 13 0 9 2
14 15 13 16 10 9 13 1 9 15 13 15 15 13 2
2 6 2
21 9 9 2 11 2 3 3 1 10 9 9 15 4 4 4 13 9 0 14 9 2
14 10 9 7 15 3 13 15 12 7 12 9 9 3 2
66 16 15 13 14 3 0 0 1 15 9 2 9 9 2 0 9 7 10 0 0 9 14 13 1 2 2 15 13 3 3 15 13 1 12 9 1 10 9 9 7 13 1 13 10 0 9 3 2 3 15 4 13 10 0 0 9 16 15 4 4 16 9 4 13 3 2
21 15 13 14 10 0 9 2 7 15 13 0 16 15 13 7 10 9 13 3 0 2
18 1 5 12 15 13 10 0 9 1 10 9 1 9 3 1 10 9 2
6 13 15 9 1 9 2
23 15 13 12 9 13 1 9 1 9 13 14 13 15 11 14 13 7 13 10 9 15 4 2
13 15 13 3 14 13 1 3 15 13 11 7 11 2
16 15 13 1 10 9 16 13 15 11 10 15 13 1 7 0 2
29 10 9 1 10 11 11 13 1 7 1 10 9 1 9 7 13 15 3 10 9 15 4 13 3 7 3 13 13 2
9 15 4 14 13 0 1 10 9 2
8 15 4 13 15 9 1 9 2
16 13 15 10 9 2 13 10 9 3 7 13 13 15 9 3 2
4 10 0 9 2
14 15 13 14 13 10 9 2 7 15 3 13 3 0 2
10 0 9 13 1 10 9 13 0 9 2
50 1 10 9 9 1 10 9 2 15 13 13 1 10 9 2 13 11 9 2 1 11 2 7 10 3 0 9 9 1 10 9 1 10 11 11 2 7 3 9 16 15 13 15 1 10 9 1 10 9 2
41 15 13 10 0 9 1 9 15 4 3 13 10 9 2 10 3 4 13 0 2 3 3 13 16 15 15 13 2 7 15 13 0 15 4 13 15 0 14 13 0 2
1 6
38 6 2 13 0 14 13 10 9 2 16 10 0 9 13 0 2 1 10 0 9 2 15 13 16 10 9 13 3 7 13 3 15 9 13 1 15 9 2
7 10 9 13 1 10 0 2
20 15 9 13 3 0 15 13 15 10 12 5 9 2 7 15 13 0 10 9 2
9 10 9 13 9 13 10 9 0 2
44 15 3 13 15 13 10 9 3 1 15 9 2 13 15 0 2 16 15 4 13 1 10 0 9 1 10 0 9 7 9 1 10 9 11 11 4 13 15 9 12 5 12 9 2
7 11 13 3 10 0 9 2
31 15 4 13 1 10 11 11 11 9 1 0 9 2 7 15 3 13 10 9 13 3 16 10 9 13 15 14 13 11 3 2
9 15 13 3 0 1 15 9 3 2
9 10 1 10 9 13 0 7 0 2
10 15 13 9 2 9 2 7 10 9 2
6 15 13 10 0 9 2
22 3 13 3 0 7 0 2 7 15 4 13 15 13 15 15 4 13 3 1 10 9 2
13 15 9 13 0 2 7 15 13 9 10 10 9 2
10 15 3 13 10 9 7 11 1 9 2
6 15 4 14 4 13 2
4 0 7 3 0
21 3 15 3 13 16 10 9 13 3 0 3 16 10 9 13 15 13 0 7 0 2
30 15 4 13 16 15 13 10 0 9 7 10 15 13 13 16 15 13 10 9 9 1 10 0 0 9 1 0 0 9 2
26 10 9 9 13 3 12 9 1 10 0 9 1 15 10 13 3 1 15 16 15 13 12 9 13 3 2
38 16 15 13 1 9 7 13 10 9 1 9 15 13 13 3 7 16 15 4 13 1 10 0 3 0 9 4 14 13 10 9 13 15 7 13 3 3 2
15 0 2 7 3 10 0 0 0 9 0 13 1 1 11 2
23 15 4 13 7 13 1 11 2 10 13 10 0 0 0 2 0 2 0 2 8 2 9 2
28 3 0 1 9 2 16 11 9 4 13 1 7 13 0 9 2 7 0 9 9 13 9 1 15 0 9 9 2
32 6 2 15 4 3 13 1 10 9 2 7 13 10 9 1 0 0 9 2 11 11 13 10 9 13 1 14 13 10 0 9 2
20 10 15 13 14 13 14 13 15 0 0 9 2 13 13 10 0 9 1 9 2
3 10 9 2
9 10 0 11 9 15 4 3 13 2
19 15 13 16 15 13 1 9 3 15 13 1 10 0 9 1 10 0 9 2
12 10 9 13 1 0 9 7 10 9 13 0 2
7 10 9 13 0 7 0 2
16 15 3 13 10 8 0 9 7 10 9 14 9 1 10 9 2
13 15 13 12 1 10 0 9 15 4 3 13 1 2
12 15 4 13 15 10 11 11 1 10 0 9 2
29 15 13 9 1 15 9 7 9 1 10 9 14 9 15 13 11 2 13 15 10 9 1 11 2 7 13 10 11 2
6 9 11 11 11 11 2
4 9 2 0 2
50 15 4 4 13 9 1 3 15 0 9 7 15 4 3 13 1 10 9 9 1 11 11 7 1 10 9 7 3 10 0 9 1 11 2 7 3 15 13 10 9 9 2 15 13 10 0 9 9 3 2
25 10 1 10 9 9 13 10 0 1 15 2 3 15 13 12 1 10 0 13 10 9 7 10 9 2
11 10 9 3 13 0 13 1 10 0 9 2
17 10 0 8 9 1 10 9 9 13 10 9 16 13 9 1 11 2
13 13 14 13 9 16 15 4 14 13 9 7 9 2
4 13 15 13 2
32 13 10 0 9 1 10 9 3 2 11 11 2 15 13 0 2 0 7 4 14 13 10 0 9 1 10 9 10 4 13 3 2
34 15 13 14 0 16 13 1 10 9 1 9 1 15 2 15 13 14 13 15 10 9 1 15 13 9 3 16 13 15 4 13 10 9 2
38 15 3 4 14 13 9 7 13 16 15 13 11 10 0 2 0 9 14 13 2 10 12 4 14 4 13 15 9 2 7 15 9 14 2 7 15 9 2
18 15 13 3 0 14 13 10 9 13 3 0 2 3 3 15 13 0 2
2 3 13
8 15 13 1 10 0 9 9 2
21 16 15 13 10 0 9 15 3 13 9 1 10 0 9 3 15 13 15 13 0 2
33 15 13 15 1 10 9 12 9 3 12 1 15 9 13 1 10 9 1 10 9 9 7 13 0 9 10 15 13 14 0 14 13 2
15 3 4 15 13 16 15 4 3 4 13 15 9 3 3 2
21 15 13 15 1 10 3 0 9 13 1 10 9 9 14 9 2 13 1 9 9 2
17 15 13 15 14 13 3 0 2 0 2 0 2 7 0 3 3 2
6 15 4 13 15 3 2
10 15 4 14 13 10 0 9 1 15 2
42 3 2 13 15 13 16 16 15 13 1 11 2 15 13 14 1 11 2 15 4 14 13 1 9 7 15 3 13 11 1 9 2 3 0 2 3 0 2 3 0 2 2
8 15 13 2 15 13 10 9 2
27 10 9 13 3 3 3 0 16 15 4 13 1 11 2 15 13 15 13 0 2 7 10 9 13 3 0 2
29 10 9 13 10 9 14 4 13 7 10 9 13 15 10 10 9 11 13 0 3 13 1 10 0 9 1 10 9 2
8 3 15 13 15 13 15 9 3
31 3 15 13 1 11 11 1 12 2 15 4 13 7 13 1 1 10 9 9 2 11 11 2 1 10 3 0 7 0 9 2
16 15 13 1 15 15 15 13 7 16 15 3 13 1 11 11 2
9 11 11 13 10 9 1 10 9 2
17 15 13 15 2 10 9 2 15 4 13 10 9 7 13 3 2 2
16 11 11 13 15 10 0 9 1 10 9 7 10 9 1 9 2
12 11 11 4 13 10 0 9 9 1 10 9 2
19 15 13 10 11 11 10 11 9 7 10 1 0 11 9 14 13 13 11 2
4 0 9 9 2
4 0 2 0 9
13 15 13 15 12 11 11 3 14 13 10 13 9 2
18 10 9 13 5 12 14 13 15 7 10 5 12 14 13 10 0 9 2
28 11 11 13 16 0 1 10 9 10 9 13 13 14 4 13 13 0 7 15 13 14 4 13 13 3 5 12 2
17 15 13 3 0 1 10 9 7 9 1 11 7 9 1 11 11 2
15 15 13 10 9 1 1 10 9 7 15 13 0 10 9 2
9 15 4 3 13 10 0 15 13 2
21 7 15 13 0 16 15 4 14 13 10 9 9 14 13 10 9 2 9 13 9 2
2 11 11
8 11 13 10 9 1 10 9 2
8 2 11 11 2 13 10 9 2
18 1 10 9 15 13 1 15 1 15 0 9 2 15 4 14 4 13 2
12 0 9 13 9 1 10 13 1 9 11 11 2
6 15 4 3 13 15 2
19 10 0 9 15 13 16 13 0 1 9 2 15 4 14 13 14 13 15 2
7 11 11 13 0 7 0 2
23 15 3 4 14 3 13 12 5 1 10 9 10 10 1 10 0 0 9 13 1 10 9 2
14 15 4 4 3 13 9 16 15 13 15 9 9 0 2
9 3 13 9 11 2 7 3 0 2
2 0 9
12 15 4 14 13 10 0 9 1 2 11 11 2
28 1 10 9 2 15 13 14 13 15 0 9 2 10 15 4 3 13 0 16 15 4 13 1 10 9 9 9 2
28 15 13 15 13 0 16 10 15 13 15 0 9 1 0 9 2 3 2 15 4 14 3 13 15 1 15 9 2
11 15 13 0 1 15 13 15 0 9 3 2
17 15 13 15 4 4 13 0 14 13 15 9 16 13 15 0 9 2
19 13 16 15 13 14 13 15 15 9 7 3 15 13 9 9 13 14 0 2
6 15 13 3 0 3 2
4 15 4 13 15
10 15 4 13 15 9 13 1 12 9 2
9 15 13 16 15 4 14 13 15 2
17 1 10 9 2 9 13 14 3 0 2 7 15 3 13 3 0 2
20 3 1 15 9 2 15 9 13 14 13 2 7 3 15 4 14 13 3 3 2
23 15 4 13 9 15 4 13 1 9 9 2 14 13 1 0 9 9 3 1 11 11 11 2
16 15 3 13 15 15 4 13 1 7 4 13 10 0 9 3 2
27 15 4 13 0 9 10 10 9 4 14 13 2 16 16 15 4 13 0 9 9 16 15 13 15 14 13 2
9 3 0 9 1 10 10 0 9 2
13 15 4 13 1 11 1 11 1 0 1 12 9 2
19 15 4 14 13 15 3 3 15 4 13 1 15 9 2 9 7 9 2 2
28 15 3 13 11 14 9 9 16 15 4 3 13 1 10 9 7 13 2 15 13 15 9 2 15 13 15 2 2
10 0 2 0 2 0 9 1 0 9 2
26 15 4 13 14 13 0 3 15 13 1 10 9 7 15 4 3 13 10 0 1 0 9 7 9 9 2
10 15 9 4 3 13 10 0 2 3 2
8 15 4 14 13 10 9 3 2
3 9 11 2
4 15 9 1 11
29 15 9 13 13 1 11 11 2 15 13 3 0 2 15 13 3 0 2 7 10 9 13 0 2 3 0 7 0 2
34 3 15 13 0 14 13 9 1 10 9 1 9 1 10 9 2 7 15 13 1 10 12 2 9 9 2 7 10 9 15 13 3 0 2
27 16 15 4 14 13 1 10 9 2 3 15 4 13 1 10 9 9 14 9 2 7 13 1 1 11 11 2
5 10 9 13 0 2
17 13 0 14 13 10 0 9 1 15 9 3 16 15 13 15 9 2
12 2 15 13 1 10 9 2 1 10 9 9 2
3 0 9 2
24 15 4 13 1 2 3 13 1 16 15 13 16 15 4 13 1 15 9 12 5 12 9 3 2
51 15 13 16 15 13 3 1 15 9 7 15 4 13 14 13 3 3 3 16 15 4 16 15 13 15 9 1 9 1 12 9 2 7 10 9 4 13 1 15 13 15 4 13 14 13 10 9 3 1 12 2
7 0 2 0 2 3 9 2
23 13 16 10 15 13 1 13 10 9 7 13 9 1 9 2 10 9 1 10 9 3 3 2
12 13 10 0 9 1 9 16 15 13 3 0 2
9 15 4 3 13 1 10 9 3 2
2 0 9
19 15 13 11 11 1 15 0 9 14 9 9 16 15 4 4 13 1 15 2
27 15 13 3 0 16 15 13 1 14 13 11 2 15 13 10 0 9 15 13 9 1 9 7 9 1 15 2
30 10 9 13 10 10 15 13 15 4 13 2 15 4 13 0 9 1 3 3 7 10 9 15 13 1 11 13 15 10 2
31 15 13 3 0 2 10 9 4 13 3 7 3 2 15 13 3 0 14 13 10 9 1 9 3 0 7 0 13 1 9 2
15 13 15 11 15 13 14 13 15 1 10 9 1 0 9 2
4 0 0 9 2
56 15 13 12 2 7 15 9 13 0 2 7 3 2 0 2 16 12 1 10 9 13 2 2 15 3 13 16 15 15 13 7 13 15 9 1 9 16 3 14 13 15 9 16 15 4 13 15 14 13 10 9 15 13 15 14 2
14 15 3 13 15 9 7 13 10 9 14 13 15 3 2
12 15 13 9 7 3 4 14 13 15 14 13 2
15 15 13 10 0 9 1 10 3 0 2 0 2 0 9 2
15 15 4 3 13 15 7 4 4 13 3 1 15 0 9 2
2 6 2
13 7 9 13 5 12 3 2 4 14 13 1 15 2
3 9 14 9
9 6 2 10 9 13 14 3 0 2
17 15 9 9 2 12 0 9 7 12 0 9 13 3 14 4 13 2
31 10 9 13 16 15 4 13 7 10 9 9 4 13 1 10 9 7 15 13 10 9 1 9 3 14 13 14 13 15 1 2
4 7 9 13 2
10 15 13 12 9 1 10 9 13 9 2
11 16 15 4 14 13 2 4 14 13 3 2
21 15 9 13 1 0 9 9 7 15 13 14 13 0 10 0 9 16 15 13 3 2
25 15 4 14 13 12 9 16 13 10 0 9 9 7 15 13 3 1 10 9 10 9 7 10 9 2
5 0 9 2 0 9
22 15 13 14 13 3 3 10 9 16 15 13 1 10 9 7 13 15 9 7 9 9 2
7 11 9 9 13 0 3 2
26 3 1 10 2 10 9 13 0 1 15 9 7 3 1 0 9 2 3 13 15 1 12 9 7 0 2
21 1 10 9 2 10 9 2 5 12 5 5 12 2 13 14 13 10 0 1 9 2
13 10 9 13 14 13 9 7 13 15 9 3 3 2
18 9 1 10 0 9 4 14 13 15 9 7 9 2 7 15 3 13 2
21 15 13 14 10 11 7 11 2 15 13 10 9 9 9 7 10 0 12 1 15 2
4 13 10 9 2
13 4 3 3 3 13 10 9 7 13 10 9 9 2
9 15 13 10 0 9 2 1 9 2
6 0 2 0 7 0 2
12 13 3 1 0 9 1 10 9 1 0 9 2
16 10 9 1 10 9 13 0 2 15 13 15 1 10 9 9 2
12 15 13 10 9 10 4 13 3 1 10 9 2
7 11 13 0 1 10 9 2
19 15 13 0 1 11 2 3 3 15 9 13 1 10 9 2 13 15 3 2
27 0 1 10 9 2 15 13 10 9 2 4 14 13 14 13 15 15 13 3 10 2 0 2 9 2 2 2
12 13 3 3 3 3 7 15 4 13 1 9 2
11 0 7 3 16 15 13 1 10 0 9 2
29 15 7 15 9 13 1 11 1 10 11 11 2 15 9 9 2 1 10 11 11 7 1 9 12 1 10 9 9 2
15 15 13 10 11 11 9 3 15 13 0 16 10 11 13 2
26 10 11 11 13 0 3 0 2 15 13 12 9 1 10 9 2 15 13 0 10 0 7 10 0 9 2
36 15 13 10 12 9 9 13 10 0 9 3 16 10 9 13 16 15 13 0 7 16 15 3 13 7 13 3 1 12 1 12 14 13 11 11 2
16 7 16 15 3 3 13 3 15 4 14 13 3 0 1 10 9
10 15 13 10 11 7 15 9 13 0 2
24 15 13 9 9 9 1 11 7 13 11 2 11 13 10 9 7 13 3 2 3 0 7 0 2
23 15 3 3 13 16 11 13 10 9 1 14 13 13 2 7 15 4 13 10 9 1 11 2
16 15 13 0 7 11 13 1 9 1 12 9 14 13 10 9 2
19 15 13 13 1 11 2 7 13 0 16 3 10 9 4 13 1 10 9 2
11 10 9 13 3 7 10 9 13 3 0 2
15 15 4 3 13 11 2 7 4 13 10 9 1 15 9 2
11 9 11 7 11 1 15 9 7 0 9 2
4 11 11 2 11
8 15 4 14 13 15 9 3 2
14 15 13 10 9 1 10 9 13 10 9 1 11 12 2
28 15 3 13 16 10 9 13 1 10 9 4 14 13 14 13 15 9 15 4 13 14 13 15 13 1 10 9 2
4 6 2 3 2
36 1 10 10 9 9 3 3 2 10 0 9 2 9 13 3 2 7 15 4 13 14 13 10 12 2 12 9 9 13 3 16 15 13 9 0 2
5 3 0 1 15 2
38 16 15 13 15 7 14 2 16 15 9 13 1 10 9 2 0 1 9 2 8 10 0 9 15 4 13 13 13 10 9 4 13 16 15 4 14 13 2
2 0 9
27 15 4 3 13 1 11 1 15 9 9 7 13 10 0 9 2 7 15 13 1 10 11 11 1 15 9 2
23 0 9 13 15 13 0 7 15 4 13 15 2 7 15 13 10 9 3 0 1 9 0 2
4 11 13 0 2
26 15 13 3 1 9 2 0 2 1 10 9 2 7 13 15 1 10 9 15 13 1 15 0 9 9 2
19 15 3 13 1 10 9 2 13 3 9 9 7 13 15 9 1 10 9 2
9 15 4 14 3 13 10 9 3 2
25 0 9 7 2 0 9 1 10 9 7 15 13 15 1 0 9 16 15 4 14 13 15 15 13 2
17 15 4 13 10 0 9 2 3 15 13 10 0 9 1 10 9 2
8 10 9 13 0 7 3 0 2
11 10 9 13 9 1 9 3 1 0 9 2
19 10 9 13 0 2 15 9 13 13 15 9 3 16 15 13 15 0 9 2
15 14 13 15 13 10 9 7 9 9 2 15 13 3 0 2
6 15 4 4 13 3 2
14 15 13 15 9 3 2 9 2 9 9 2 7 9 2
12 9 13 0 2 3 0 1 10 9 7 9 2
15 15 4 3 13 0 9 3 0 2 15 13 3 3 0 2
14 3 15 13 9 1 7 15 4 14 13 1 9 3 2
4 15 13 11 11
3 4 13 3
34 9 2 2 11 2 10 9 2 13 3 0 7 3 13 1 15 9 2 3 0 9 2 0 9 2 3 15 0 9 9 2 15 13 2
18 4 14 13 3 3 15 4 13 0 9 9 7 10 1 10 0 9 2
31 9 2 2 9 13 14 3 0 2 3 0 9 1 10 13 9 2 13 9 2 9 2 13 3 12 9 1 9 1 9 2
11 10 10 9 7 9 13 0 1 10 9 2
9 0 9 2 4 13 10 9 3 2
12 15 4 13 10 9 3 0 9 13 15 3 2
18 15 9 9 13 0 2 3 15 4 13 15 9 2 7 10 0 9 2
5 3 0 2 3 0
11 10 9 1 11 11 13 3 0 7 0 2
41 15 4 13 1 10 9 7 4 14 3 13 15 15 13 7 15 13 3 0 7 13 10 9 14 3 13 1 15 15 9 13 7 13 15 0 9 14 13 10 9 2
18 15 13 3 0 16 13 15 13 10 0 9 3 1 3 13 10 9 2
16 15 9 1 15 13 0 2 0 9 2 3 0 7 3 0 2
23 16 13 10 9 15 13 15 13 10 9 14 13 1 10 9 7 13 15 3 0 16 0 2
9 1 9 1 9 15 13 0 9 2
13 15 4 3 13 13 10 9 1 1 15 0 9 2
7 10 9 9 13 10 9 2
8 15 13 3 10 9 9 3 2
20 16 15 4 14 13 4 13 2 13 7 13 1 3 15 13 10 9 1 15 2
11 15 4 13 10 9 14 13 7 13 15 2
14 15 13 1 9 1 9 14 13 15 9 9 1 9 2
44 1 10 9 15 13 9 1 12 1 1 12 0 9 9 1 10 0 9 7 13 10 9 1 10 9 1 10 9 1 9 15 13 4 14 13 9 1 0 13 9 1 10 9 2
20 15 3 13 10 9 1 12 0 9 7 15 13 15 13 10 9 1 15 9 2
11 11 13 10 9 16 15 13 10 0 5 2
3 0 9 2
23 15 4 13 3 10 0 9 1 9 9 7 3 13 15 9 2 9 7 9 9 13 9 2
30 15 13 15 3 7 15 13 3 0 1 9 7 3 13 9 1 15 9 10 4 13 10 9 7 13 15 0 9 9 2
15 15 3 13 1 0 9 7 9 1 10 9 1 10 9 2
36 15 13 15 0 13 16 15 13 9 16 16 15 4 14 13 14 13 3 7 13 9 1 1 9 14 13 3 7 3 7 13 14 13 10 9 2
9 0 9 2 0 9 7 3 0 2
21 15 3 4 14 13 16 15 13 14 13 15 10 9 1 9 10 15 4 14 13 2
5 13 15 9 1 11
24 15 13 1 11 11 1 11 12 1 10 12 2 9 9 7 4 3 13 15 1 10 12 9 2
18 10 9 1 11 7 11 1 10 9 9 2 3 11 2 13 3 0 2
12 15 4 13 3 0 3 15 4 13 1 9 2
21 16 10 9 13 13 11 11 7 0 1 10 11 11 11 2 10 9 13 3 0 2
14 15 4 3 13 10 9 1 0 9 7 9 1 9 2
18 10 9 13 1 9 9 1 11 11 14 2 11 11 2 7 0 9 2
11 10 3 2 13 2 0 9 13 10 9 2
14 0 9 14 13 16 15 13 1 7 3 3 11 11 2
9 15 13 0 9 1 10 9 9 2
48 11 11 13 1 7 15 13 12 9 2 10 15 13 13 12 5 9 9 2 15 13 10 0 2 15 13 9 12 3 15 4 4 13 9 3 2 13 1 10 10 9 10 13 15 13 0 2 2
31 14 3 4 15 13 13 1 16 15 3 13 16 15 15 13 2 10 15 13 0 1 13 15 13 10 9 3 3 7 3 2
14 3 0 0 9 7 1 10 9 1 0 9 0 9 2
18 15 13 0 15 13 15 9 7 4 14 4 13 16 13 9 1 15 2
16 13 9 15 13 10 3 13 15 7 13 14 13 10 9 3 2
8 4 14 13 15 9 7 9 2
30 15 13 15 12 9 0 9 3 1 10 9 7 14 13 0 2 3 1 10 9 9 2 15 13 15 13 9 7 0 2
31 3 13 1 9 10 9 16 15 12 9 0 13 14 13 0 1 10 9 3 2 15 13 15 3 1 12 9 9 1 9 2
16 16 15 4 13 1 10 11 11 15 4 14 3 13 1 15 2
32 16 15 13 3 0 1 9 14 13 10 9 7 13 0 14 13 1 10 0 9 1 5 12 1 12 12 9 3 13 1 15 2
23 2 1 10 9 15 4 14 13 15 13 15 12 9 2 15 4 14 13 12 1 15 2 2
15 11 11 7 11 11 2 15 4 14 13 11 11 11 3 2
19 15 13 10 0 9 16 13 10 9 16 15 13 7 4 13 1 11 11 2
16 15 3 13 15 1 9 7 15 0 9 4 13 3 9 0 2
21 15 0 9 4 4 13 7 15 3 3 13 10 9 9 3 15 0 9 13 0 2
41 1 9 1 10 9 9 2 11 11 4 13 15 3 1 15 9 7 9 1 10 3 2 9 1 15 9 2 15 0 9 13 1 10 0 9 1 9 1 10 9 2
20 15 13 3 0 14 13 10 0 9 14 13 16 10 9 9 4 13 1 3 2
2 11 11
5 0 9 2 6 2
15 16 15 9 4 13 1 2 15 13 15 10 9 1 9 2
20 10 9 13 15 16 15 13 10 0 9 15 4 3 13 2 7 15 13 0 2
3 10 9 2
50 15 13 14 13 13 15 1 3 1 10 9 2 7 11 2 15 13 10 9 3 5 10 9 3 2 15 13 10 3 0 9 2 15 13 10 0 9 13 10 9 9 10 12 9 9 7 15 13 3 2
23 3 0 2 4 14 13 15 0 2 7 15 9 13 0 7 0 3 15 13 3 1 9 2
23 7 10 9 2 13 0 14 13 1 10 9 7 13 9 1 9 3 2 15 4 13 15 2
5 11 11 13 15 9
9 6 2 11 11 13 14 3 0 2
13 15 13 15 0 9 1 15 7 15 13 3 0 2
44 15 13 1 10 9 1 10 9 7 16 15 13 7 15 13 15 1 1 10 9 9 15 13 16 0 9 1 10 9 3 13 9 13 1 11 11 1 0 9 7 13 3 0 2
26 16 15 13 15 3 1 9 2 10 0 9 7 15 4 3 13 10 9 13 9 1 15 9 3 3 2
28 6 2 15 3 13 15 1 10 9 2 5 12 2 7 13 10 9 14 13 15 10 5 12 2 9 2 9 2
9 15 3 13 15 1 10 9 9 2
5 13 1 10 9 2
5 12 1 10 0 9
16 10 9 7 15 9 9 11 11 13 10 0 9 14 13 1 2
29 10 9 13 0 14 13 16 15 4 13 2 15 13 10 9 0 1 10 9 1 9 2 7 3 13 1 15 9 2
43 15 13 14 13 3 1 3 12 9 3 7 10 9 2 15 13 14 13 10 9 2 13 15 9 13 1 10 9 2 7 15 4 14 13 14 13 15 1 10 9 1 9 2
14 15 13 10 12 9 16 13 15 9 7 15 13 0 2
33 1 15 9 10 9 4 4 13 1 1 10 9 9 2 7 9 15 13 0 1 15 9 7 9 4 3 13 1 10 0 0 9 2
6 13 3 1 9 1 9
2 6 2
7 15 13 14 13 10 9 2
14 7 3 16 15 13 9 1 10 9 2 9 4 13 2
23 15 4 13 3 1 11 1 15 9 7 0 9 15 13 1 15 2 15 13 15 9 9 2
8 0 15 13 10 9 1 15 2
19 1 9 15 4 14 13 0 16 7 13 10 9 7 13 1 10 0 9 2
19 2 10 0 9 9 13 0 14 13 2 15 4 14 3 13 1 11 2 2
17 13 1 10 9 1 9 7 13 10 9 2 15 4 13 0 9 2
29 3 2 16 11 13 12 9 1 0 9 1 1 9 1 10 0 0 9 9 2 15 4 13 0 14 13 1 11 2
14 9 7 15 13 14 13 10 9 7 13 9 7 0 2
14 15 13 11 1 3 12 7 13 10 9 15 3 13 2
14 15 4 13 16 15 4 14 9 16 15 4 13 3 2
16 15 13 10 0 9 14 13 15 13 15 9 4 4 13 3 2
33 15 13 15 10 9 9 7 13 9 3 14 13 1 14 13 15 9 0 13 15 7 15 4 13 14 13 3 7 13 1 10 9 2
13 15 13 12 9 3 7 13 15 9 1 10 9 2
3 15 13 2
5 0 9 3 3 2
19 1 12 9 15 13 15 10 9 4 4 13 2 10 0 9 15 13 14 2
11 0 9 1 9 13 9 7 13 9 9 2
11 9 13 10 9 7 10 9 13 10 9 2
8 13 1 10 9 3 8 0 2
10 15 4 14 13 10 9 15 4 13 2
27 15 13 14 13 3 15 0 9 7 15 13 14 13 16 15 14 13 15 16 15 13 14 3 15 4 13 2
18 13 3 16 13 15 4 13 15 13 10 9 1 9 6 15 13 14 2
5 9 13 8 0 2
18 13 3 15 13 10 9 4 14 13 1 10 9 13 3 1 10 9 2
7 8 0 16 9 14 13 2
37 13 1 10 9 9 15 4 14 13 14 13 10 9 9 3 3 15 13 10 0 0 9 16 13 9 15 4 14 13 0 14 13 3 1 10 9 2
2 13 2
4 15 4 13 9
13 10 9 13 9 16 15 4 13 9 1 0 9 2
35 15 13 9 1 9 16 15 13 10 0 9 2 3 1 9 15 13 10 3 0 9 3 3 2 15 13 3 10 0 9 9 1 10 9 2
37 15 13 9 10 13 14 3 9 2 13 9 10 13 10 9 13 1 10 0 9 3 15 13 14 2 10 0 9 1 9 9 2 7 3 7 3 2
8 1 0 1 0 9 14 13 2
18 3 4 14 4 13 3 2 13 15 9 0 16 15 13 14 13 3 2
28 1 10 0 9 2 10 11 11 9 4 13 1 15 9 9 2 15 9 9 2 7 15 9 1 10 0 9 2
2 3 3
26 4 14 13 3 16 15 13 14 13 2 13 2 13 7 4 13 14 13 3 1 10 9 1 12 9 2
31 15 4 14 3 13 9 14 13 10 0 9 16 4 13 14 13 7 16 15 13 1 0 9 15 9 4 13 1 10 9 2
20 15 13 10 0 9 15 4 3 13 7 4 13 14 13 16 0 9 4 13 2
16 15 4 13 14 13 15 9 14 13 16 15 13 14 13 15 2
15 6 2 7 15 9 9 13 0 3 10 0 9 7 9 2
25 7 10 9 13 9 9 2 13 9 13 14 13 10 0 9 9 14 13 15 9 2 9 7 9 2
10 13 0 9 1 10 11 11 11 3 2
9 15 13 15 13 15 15 13 1 2
22 15 13 14 13 3 1 10 0 9 1 15 9 2 3 15 13 1 10 0 9 9 2
22 15 13 3 2 7 15 4 13 1 10 0 2 9 2 1 10 9 1 12 0 9 2
21 16 15 13 15 10 9 2 15 13 15 0 9 13 1 7 4 14 13 15 9 2
22 3 15 4 13 1 10 9 1 10 0 9 1 10 9 2 3 1 1 10 9 9 2
16 15 4 13 10 0 9 10 13 3 16 15 13 1 15 9 2
32 3 15 3 13 9 1 10 9 15 4 13 11 2 15 13 15 9 2 7 15 3 4 14 13 10 0 9 15 4 2 13 2
5 15 13 3 0 2
13 15 13 10 9 16 10 9 1 15 9 13 3 2
24 15 13 10 0 0 9 1 10 9 14 13 9 2 15 13 14 10 0 15 13 7 3 0 2
29 10 0 9 13 15 13 15 0 9 13 1 3 10 0 9 10 0 9 4 13 3 14 13 10 9 9 7 9 2
20 15 13 10 9 0 1 3 10 10 9 13 10 13 15 7 15 9 3 0 2
21 15 4 13 9 1 9 1 15 9 3 9 13 3 2 15 4 4 13 10 9 2
8 3 0 9 7 0 9 3 2
9 0 9 15 4 13 1 9 3 2
15 15 3 13 10 9 13 9 9 14 13 10 9 10 9 2
5 0 9 9 13 0
20 10 11 11 11 4 13 1 15 11 11 9 1 10 0 9 1 11 11 11 2
21 10 0 11 13 12 9 13 7 3 13 10 0 0 9 9 9 1 11 1 11 2
29 10 9 13 10 9 7 9 9 2 1 9 2 0 2 9 2 9 2 9 2 9 9 2 9 2 9 7 9 2
39 15 4 13 8 11 11 11 1 1 10 9 7 3 13 10 0 7 0 9 15 4 13 9 7 0 3 3 1 10 9 13 0 9 9 13 10 11 9 2
29 15 13 14 3 0 14 13 10 9 3 3 2 15 4 13 15 12 1 1 12 7 12 9 1 10 9 11 7 11
14 15 13 10 12 2 9 0 0 0 11 1 10 9 2
17 10 9 15 13 3 3 2 15 13 16 10 0 9 13 10 9 2
11 2 15 4 13 10 9 16 13 1 9 2
10 3 0 15 13 10 0 9 9 2 2
18 15 13 16 15 4 4 13 9 1 10 9 1 0 9 1 9 9 2
12 2 7 15 13 10 0 9 1 10 9 2 2
10 3 15 13 10 9 3 10 0 9 2
22 15 13 15 16 15 13 14 1 9 7 13 14 13 15 5 12 3 14 13 10 9 2
14 15 13 3 0 15 13 15 14 13 14 13 10 9 2
4 15 13 3 2
10 3 15 9 13 16 3 13 10 9 2
7 13 3 3 3 16 0 2
2 0 9
20 16 15 4 13 10 11 11 11 15 13 10 0 7 0 9 1 9 1 9 2
31 9 13 0 1 10 9 1 10 9 15 2 13 15 1 15 9 7 13 10 0 9 2 7 3 7 3 16 15 13 3 2
27 9 9 9 4 3 13 14 13 15 7 3 15 7 15 13 15 10 9 16 15 13 7 13 0 1 15 2
21 10 9 15 13 0 2 0 7 3 0 7 15 3 13 16 15 13 1 0 9 2
28 15 0 9 2 11 11 11 13 3 10 0 9 7 3 0 7 1 10 9 15 13 7 10 9 15 4 13 2
13 9 13 3 0 16 15 4 14 13 14 13 3 2
1 11
5 0 9 1 0 9
23 15 13 15 9 9 1 10 11 14 11 2 7 15 13 12 1 10 0 9 10 15 13 2
35 15 13 10 0 9 2 15 13 10 0 9 1 9 2 7 15 9 7 15 13 12 9 1 9 7 10 9 13 3 3 0 16 15 13 2
8 15 4 3 13 9 7 9 2
26 15 13 10 0 9 2 3 12 9 7 3 2 7 3 9 4 13 3 7 15 10 13 10 0 9 2
32 3 16 15 4 3 13 14 13 10 0 9 1 9 2 3 9 13 1 10 0 9 2 15 4 13 3 1 10 9 1 15 2
19 15 3 13 11 14 16 13 10 0 9 3 0 1 15 0 9 7 9 2
1 0
11 15 13 1 11 16 13 10 1 10 9 2
20 15 13 1 9 1 10 9 7 3 13 16 15 13 3 14 13 15 9 13 2
13 15 13 15 13 9 14 13 1 7 13 10 9 2
11 11 13 15 9 7 15 13 15 15 13 2
12 15 13 0 9 7 15 13 1 15 9 9 2
15 15 13 10 0 9 15 4 13 10 9 16 15 9 0 2
27 3 15 13 13 15 1 7 15 13 14 13 16 15 13 15 14 13 15 15 4 13 1 1 15 0 9 2
30 7 15 13 10 0 9 13 15 13 15 15 4 13 1 10 9 7 13 15 9 1 10 9 15 4 13 15 1 9 2
6 15 13 14 3 0 2
5 15 4 3 13 3
26 16 3 13 1 11 11 2 15 4 13 1 10 0 2 0 2 7 0 9 1 11 11 14 11 9 2
25 15 13 0 1 10 9 9 1 1 10 0 9 7 9 1 10 9 2 7 9 1 10 11 11 2
17 10 9 13 3 0 7 13 9 2 3 16 13 10 0 11 9 2
16 10 0 9 13 0 0 9 7 10 11 0 9 13 3 0 2
53 1 15 9 2 15 9 13 15 10 9 1 10 9 9 3 15 4 13 15 4 13 10 5 12 5 9 14 13 7 13 1 10 9 2 1 10 9 15 4 3 13 10 9 3 7 4 13 14 13 15 9 9 2
11 15 13 10 0 1 0 9 1 11 14 2
12 13 1 10 9 2 15 4 13 3 0 1 2
6 12 9 13 3 0 2
16 0 9 13 13 9 3 1 10 13 7 15 13 15 4 13 2
43 15 4 3 13 1 10 9 1 10 9 3 10 9 13 0 2 10 9 13 0 1 0 9 14 9 1 15 2 10 9 9 13 13 7 0 7 10 9 13 0 1 9 2
37 15 13 9 14 13 16 15 13 10 9 10 9 13 1 7 4 13 2 15 13 10 11 11 2 3 10 11 2 7 10 0 3 13 1 1 15 2
14 14 13 15 14 13 3 1 10 9 3 13 14 0 2
23 15 13 14 12 9 1 9 0 7 9 15 4 13 1 10 0 9 1 9 4 4 13 2
5 9 7 0 9 9
15 16 13 11 16 13 11 9 4 13 1 10 11 13 9 2
10 15 4 13 10 0 9 16 13 9 2
14 13 10 9 9 2 13 12 0 9 13 10 0 9 2
11 13 9 9 1 9 13 3 10 0 9 2
7 3 11 4 13 10 9 2
12 11 13 15 14 13 10 9 1 10 0 9 2
25 9 1 9 9 7 0 9 1 9 1 0 9 1 9 1 9 2 9 7 9 13 3 0 3 2
12 3 3 4 15 13 14 13 0 9 1 9 2
21 9 13 12 9 7 0 9 9 13 12 9 14 9 3 0 15 9 9 4 13 2
5 1 9 2 0 2
13 1 9 2 15 13 10 9 14 13 15 9 13 2
7 4 14 13 14 13 3 2
14 15 13 1 3 10 0 9 10 15 4 3 13 1 2
25 15 13 1 11 11 1 10 0 9 7 15 9 13 1 10 11 11 16 10 15 9 14 13 1 2
15 15 4 14 4 13 3 13 2 3 0 7 3 3 13 2
18 10 9 13 0 1 10 9 2 1 0 9 1 11 7 15 0 9 2
18 9 13 3 0 7 3 13 1 1 15 9 14 13 0 9 13 3 2
42 15 4 14 13 14 13 3 1 11 11 7 1 10 0 9 2 3 15 12 9 0 2 15 13 9 1 11 11 7 10 10 9 2 7 4 13 1 15 16 15 13 2
15 15 4 3 13 10 11 11 1 15 0 9 1 11 11 2
16 0 9 2 15 13 1 11 11 7 13 12 1 15 13 9 2
15 11 13 3 2 13 5 12 9 3 14 13 1 10 9 2
32 15 13 10 9 1 15 9 2 10 9 13 3 0 3 15 13 3 13 2 13 10 9 7 13 10 0 9 1 10 0 9 2
34 10 0 9 13 5 12 2 0 1 9 16 15 11 13 2 14 13 7 13 15 1 10 9 1 10 9 9 2 10 11 13 14 2 2
18 15 9 13 3 1 10 10 9 1 11 1 10 0 9 7 0 9 2
11 13 1 15 16 11 13 3 0 16 0 2
27 3 0 1 11 11 3 3 2 15 13 16 15 13 15 9 1 9 7 9 1 9 2 3 15 13 14 2
9 11 11 1 11 11 1 11 2 11
22 3 13 15 13 1 16 13 2 16 15 4 13 3 0 9 1 11 11 1 11 11 2
18 15 13 3 0 16 10 9 4 13 1 11 2 16 15 13 1 11 2
19 15 13 3 12 9 3 7 13 10 0 9 10 15 4 13 1 15 9 2
14 15 13 12 1 15 7 15 4 13 3 1 10 9 2
12 15 13 15 9 1 10 9 7 15 13 0 2
6 15 4 13 15 1 2
11 15 3 13 15 9 16 13 15 9 3 2
12 16 10 9 13 12 9 2 15 13 10 9 2
18 10 0 9 13 10 0 9 2 10 13 9 9 1 10 9 1 9 2
15 9 1 15 4 4 13 15 9 3 2 10 13 10 9 2
5 0 9 2 0 9
11 11 13 0 7 0 1 9 1 2 9 2
18 15 13 0 14 13 1 15 1 15 0 9 7 13 10 9 1 9 2
21 10 9 4 13 1 10 9 9 7 15 13 3 0 7 0 13 2 10 15 13 2
21 10 9 9 13 16 3 15 13 10 9 1 9 1 10 9 1 0 9 2 9 2
13 15 13 1 11 1 12 9 7 13 9 7 9 2
20 10 9 13 0 7 15 13 0 1 15 7 4 14 13 10 9 1 15 9 2
33 15 13 15 4 13 10 9 1 9 7 4 14 13 10 9 2 7 1 12 9 15 13 16 15 13 14 3 0 10 9 2 9 2
14 2 15 13 3 10 0 0 1 10 10 13 9 2 2
6 0 2 0 7 0 9
18 10 9 13 3 0 2 7 13 15 0 9 1 9 7 9 9 9 2
16 0 9 13 0 7 0 2 3 0 9 14 13 7 13 2 2
17 10 0 9 10 4 13 10 9 1 12 9 2 0 0 0 9 2
38 0 7 0 9 2 10 9 0 3 9 4 13 3 3 1 10 9 3 2 7 15 4 14 13 3 3 16 15 4 3 3 13 3 1 10 9 3 2
6 10 9 13 3 0 2
21 15 13 3 1 11 11 11 7 10 12 9 9 1 11 11 10 13 0 1 9 2
19 15 13 0 1 9 9 1 11 11 2 11 11 2 7 10 0 9 9 2
15 15 3 13 15 9 7 4 3 13 1 10 11 11 3 2
5 11 11 13 15 2
22 13 0 7 0 2 3 13 15 9 13 10 9 2 15 4 13 10 0 9 1 0 2
8 15 3 13 15 15 4 13 2
45 10 9 13 1 15 9 7 13 1 15 9 14 9 2 15 13 10 9 7 13 3 0 0 7 0 2 15 4 13 1 10 9 16 10 9 4 14 13 2 15 13 15 3 2 2
22 15 13 10 0 9 2 13 15 13 10 9 13 15 10 9 2 15 13 10 9 9 2
22 3 15 9 14 9 7 9 4 3 13 3 3 2 3 15 13 16 13 10 0 9 2
28 3 6 2 15 4 14 13 16 13 10 9 1 11 11 1 0 0 9 9 2 13 15 11 11 1 15 9 2
8 15 13 3 9 1 11 11 2
31 15 4 13 2 15 13 0 1 10 9 1 10 9 9 7 9 2 7 15 13 16 15 4 13 10 9 3 1 10 9 2
14 15 13 10 9 1 9 2 11 2 11 11 7 9 2
19 10 13 0 2 7 15 13 10 9 13 9 10 13 0 1 10 0 9 2
52 1 15 9 7 9 2 15 13 1 10 9 1 15 11 11 11 2 15 4 13 15 13 0 2 1 10 0 9 7 15 13 10 11 9 3 13 1 15 2 15 13 15 13 0 2 15 13 3 0 7 0 2
14 16 15 13 1 11 15 13 14 13 13 10 9 1 2
12 10 0 9 15 13 1 10 9 13 10 9 2
9 15 13 1 10 9 1 11 2 2
3 9 9 9
15 15 9 4 13 15 12 11 11 3 1 10 0 9 9 2
30 10 9 9 1 10 9 9 2 10 9 13 3 2 10 0 9 9 9 4 13 1 3 2 7 10 9 4 13 3 2
24 13 1 10 9 13 10 9 2 7 3 9 4 13 3 2 15 4 3 13 1 1 10 9 2
15 15 4 13 2 3 4 14 13 2 0 9 1 10 9 2
9 10 1 15 13 1 15 9 9 2
25 16 15 13 15 9 15 13 10 9 7 9 9 1 15 9 14 9 7 13 15 3 14 13 15 2
19 15 4 14 13 10 9 1 9 2 3 3 9 3 0 1 10 9 9 2
16 7 15 4 13 15 1 3 3 9 2 7 13 16 13 15 2
5 9 2 0 9 2
10 13 15 11 3 3 1 0 9 9 2
10 10 0 9 15 13 14 13 0 9 2
17 3 2 15 4 3 13 10 9 16 15 1 15 14 13 15 9 2
10 15 13 16 15 4 13 1 10 9 2
11 15 13 15 14 13 15 3 1 12 9 2
8 15 13 15 3 1 12 9 2
14 15 2 13 2 10 9 7 13 15 10 9 13 0 2
18 15 13 1 15 4 14 3 13 10 9 2 13 15 13 1 15 3 2
15 15 3 4 14 13 10 9 1 15 14 13 15 9 9 2
31 15 3 13 3 14 13 9 0 1 10 9 9 2 10 0 9 2 2 7 3 15 13 10 9 3 15 13 10 0 9 2
10 15 4 3 13 10 9 1 11 11 2
2 0 9
19 15 13 14 13 16 11 13 10 0 9 1 15 9 1 15 9 1 9 2
14 10 15 9 13 3 12 9 3 7 11 13 3 0 2
26 15 13 10 3 0 9 1 15 9 7 15 7 11 13 10 9 14 13 10 7 10 12 12 1 15 2
27 15 13 3 0 1 15 9 1 10 9 7 7 15 3 13 9 14 13 0 16 15 15 4 3 13 1 2
22 15 13 0 15 13 14 10 9 16 10 9 9 13 10 0 9 1 10 10 0 9 2
21 15 9 13 3 3 1 15 9 2 7 15 9 13 3 1 10 0 9 1 9 2
11 10 15 9 13 3 0 16 4 4 13 2
11 13 15 11 1 10 15 9 3 7 3 2
3 10 11 9
2 0 9
19 16 15 13 10 9 13 1 0 9 2 11 2 2 15 4 13 15 3 2
9 15 13 15 9 1 3 12 9 2
7 15 13 12 9 1 15 2
10 10 9 13 15 13 3 12 9 9 2
26 3 2 15 13 7 13 7 1 10 8 9 2 13 12 9 1 9 3 3 13 3 16 13 15 9 2
19 10 13 1 9 4 13 1 10 9 2 10 9 2 13 15 9 3 2 2
15 15 13 14 13 10 9 2 15 13 15 9 1 0 11 2
8 15 4 14 13 10 15 9 2
15 15 4 3 13 15 16 15 4 13 10 9 15 13 3 2
29 15 9 13 16 15 4 3 13 3 16 15 13 14 13 3 3 10 9 7 13 10 9 0 9 4 13 1 15 2
5 9 3 13 1 2
20 11 9 2 15 4 13 1 1 11 14 12 9 9 2 9 9 1 11 2 2
11 15 3 13 12 9 3 16 10 9 13 2
7 10 9 4 14 13 1 2
9 15 13 1 12 9 7 3 13 2
22 15 13 12 1 15 9 2 7 10 0 9 13 3 1 10 9 9 13 1 10 9 2
16 6 2 3 3 15 4 13 16 15 13 3 0 1 10 9 2
9 15 13 15 0 9 1 15 9 2
32 1 9 14 0 9 2 15 13 10 9 16 10 9 3 14 3 4 13 15 10 9 9 7 9 16 15 4 13 14 13 0 2
18 1 10 9 9 2 15 13 0 15 13 3 0 16 10 9 13 9 2
13 7 3 9 4 13 15 1 10 0 9 1 11 2
2 0 2
2 3 2
5 15 13 14 13 2
7 10 9 13 0 3 3 2
12 3 3 0 7 13 3 16 13 0 9 0 2
17 15 13 3 0 2 7 3 0 1 15 9 1 9 1 15 9 2
47 15 13 3 13 14 13 9 1 12 1 10 0 9 2 16 6 2 15 13 14 10 0 2 7 10 0 9 1 10 9 1 12 9 1 10 13 0 3 15 13 10 0 9 13 14 13 2
34 15 4 14 13 14 13 15 9 1 9 13 1 9 2 7 15 4 14 13 14 13 1 9 15 4 14 13 3 14 13 15 1 9 2
20 13 10 9 2 1 0 9 7 10 3 0 9 1 0 2 0 2 7 0 2
18 3 2 10 0 9 1 10 9 2 10 9 1 10 1 1 9 9 2
5 0 9 1 9 2
2 6 2
6 10 9 13 10 0 2
13 15 13 0 2 0 9 2 7 13 3 7 3 2
18 15 3 13 14 13 1 10 9 2 7 15 13 10 9 10 0 9 2
29 15 13 15 9 10 15 4 4 3 4 13 1 2 7 13 0 9 14 13 1 15 3 15 13 15 1 10 9 2
19 13 10 9 13 10 0 16 15 13 10 9 1 10 9 13 10 0 9 2
23 15 4 13 0 7 4 14 13 15 13 15 2 16 15 9 1 9 3 13 15 15 13 2
24 15 13 10 9 9 10 13 1 1 10 9 2 7 15 9 13 1 10 9 9 1 10 9 2
19 3 15 4 14 13 15 14 3 13 10 1 10 9 10 15 13 10 9 2
7 15 3 3 13 15 9 2
8 3 13 13 1 10 9 3 2
13 15 13 12 9 0 7 13 0 9 15 0 9 2
12 1 10 9 1 12 15 13 13 1 10 9 2
10 15 9 7 9 1 0 9 13 15 2
13 15 13 10 10 9 15 4 13 14 13 10 9 2
13 1 10 0 9 1 15 9 2 15 3 13 3 2
11 15 13 3 13 16 13 3 7 3 13 2
17 11 11 7 15 0 9 13 10 3 0 9 15 4 3 13 1 2
22 15 13 15 13 0 16 15 15 4 13 2 7 13 15 1 10 9 1 15 0 9 2
7 15 3 13 9 7 9 2
19 10 9 14 13 7 13 3 4 3 4 13 1 10 3 0 9 1 9 2
15 13 15 11 11 2 11 11 2 11 11 7 10 0 9 2
10 11 11 11 0 9 2 11 11 11 11
4 0 9 7 9
16 3 3 13 10 9 3 0 16 15 15 13 2 15 13 0 2
47 1 10 9 2 15 13 10 9 7 15 13 0 9 7 0 9 16 15 13 0 9 2 7 15 13 10 9 2 2 2 10 9 4 13 1 9 7 10 9 13 10 9 1 10 0 9 2
22 9 15 13 1 10 9 2 1 9 2 3 10 9 13 0 2 1 3 12 0 9 2
22 15 13 3 12 9 16 15 9 14 13 3 7 1 10 9 15 12 9 0 13 15 2
12 4 15 3 13 3 3 1 10 9 7 9 2
30 15 13 10 9 1 9 7 10 0 9 13 14 13 9 1 0 9 1 9 2 16 15 13 10 0 14 13 15 9 2
13 15 4 14 13 13 10 9 3 7 3 13 3 2
6 11 11 13 3 0 2
5 9 7 9 9 2
10 15 13 10 9 16 10 9 13 0 2
63 7 15 13 15 9 13 1 15 13 5 0 9 7 9 9 7 10 9 15 13 15 1 13 3 1 10 10 9 7 10 9 3 2 7 12 9 3 15 13 14 13 15 1 15 0 9 16 10 9 1 10 9 1 11 13 10 0 9 7 15 13 9 2
42 15 9 3 13 15 13 14 15 9 15 13 10 9 10 13 10 9 2 3 15 4 14 13 13 10 9 16 15 13 10 0 12 9 7 3 1 9 7 10 9 9 2
22 15 4 13 15 4 13 10 0 9 7 15 4 14 13 16 15 4 4 13 0 9 2
5 10 13 3 0 2
23 3 14 13 10 9 16 15 13 15 15 9 3 3 3 12 9 16 15 13 3 1 9 2
3 9 9 2
10 15 13 10 0 9 1 10 0 9 2
17 15 9 9 2 11 11 2 11 11 13 10 9 7 9 13 0 2
9 3 15 13 10 9 1 5 12 2
13 10 9 14 9 13 16 9 4 4 2 13 2 2
9 11 11 13 10 9 1 10 9 2
15 10 9 13 15 9 14 13 15 15 13 1 11 2 11 2
18 15 3 13 15 1 1 10 9 9 7 3 4 14 3 13 10 9 2
35 15 3 13 14 3 13 10 9 3 16 10 9 4 3 4 13 2 7 3 10 9 9 4 13 14 13 10 9 1 5 12 4 13 3 2
6 15 13 10 0 9 2
7 3 0 4 15 3 13 2
21 3 3 4 15 4 13 1 9 15 4 14 13 2 10 9 9 13 0 14 13 2
11 15 13 10 9 13 10 0 9 9 9 2
24 15 4 4 13 14 13 11 11 3 7 4 14 13 9 0 14 13 15 9 2 9 2 8 2
17 15 4 13 1 10 9 1 0 9 16 15 9 4 3 4 13 2
10 15 13 10 0 9 7 0 9 9 2
15 1 12 9 2 15 13 15 13 7 13 1 10 0 9 2
7 15 13 15 1 10 9 2
6 15 3 13 15 9 2
15 15 13 10 9 10 4 4 4 13 16 13 16 15 13 2
16 15 13 7 13 1 15 14 13 15 16 16 15 4 13 0 2
8 15 3 13 15 10 0 9 2
12 15 13 12 9 2 15 3 13 12 7 0 2
19 16 15 13 9 14 13 12 2 15 13 10 0 9 2 7 13 15 3 2
18 15 13 10 9 1 9 7 9 10 13 0 9 13 1 10 0 9 2
9 15 13 10 9 1 9 1 15 2
1 9
10 15 13 10 9 16 13 1 10 9 2
13 15 13 12 9 9 1 10 9 1 10 13 9 2
21 15 3 13 9 13 10 9 13 0 7 2 15 13 9 3 0 1 10 9 2 2
14 6 15 13 10 13 9 13 1 10 9 1 9 6 2
12 3 15 9 13 15 16 15 4 13 15 3 2
23 10 0 9 15 13 15 1 12 9 9 7 15 10 13 15 10 0 9 2 9 13 9 2
15 15 13 7 13 10 0 9 1 9 7 9 13 15 3 2
38 1 10 0 9 2 15 9 4 3 13 14 13 12 9 1 9 10 13 10 9 14 13 7 13 15 9 3 15 13 15 13 3 10 9 1 9 9 2
14 16 15 13 12 9 15 4 13 15 1 7 12 9 2
6 0 9 15 9 13 2
11 13 15 9 9 0 1 15 12 9 9 2
5 0 9 9 1 11
20 11 2 10 0 11 2 11 9 9 7 9 9 2 3 13 10 0 9 3 2
28 15 13 3 1 10 9 7 9 1 11 11 7 10 4 13 15 16 15 4 13 1 1 11 11 7 11 14 2
13 15 13 3 1 15 9 9 9 9 9 1 11 2
13 15 13 10 0 0 9 13 1 9 1 9 9 2
33 9 2 9 9 2 9 2 7 10 9 14 13 3 7 13 1 9 14 13 15 0 9 7 16 10 0 15 9 9 9 4 13 2
36 15 13 10 9 15 13 1 9 10 2 15 4 4 13 2 2 9 14 13 15 13 16 11 4 13 10 0 9 16 13 13 10 9 1 11 2
15 15 13 1 13 10 9 9 7 4 3 13 3 1 0 2
12 9 2 9 2 9 2 9 2 9 2 13 2
5 13 1 1 15 9
6 13 1 1 15 9 2
8 10 9 13 0 1 15 9 2
31 15 13 15 16 13 10 9 7 9 9 9 1 0 9 7 15 3 13 15 4 13 14 13 15 1 1 10 13 0 9 2
21 1 10 0 9 9 10 15 4 13 2 15 13 3 9 1 9 1 15 0 9 2
30 10 0 9 13 16 15 4 14 3 13 3 1 10 9 15 13 1 2 15 3 13 2 9 2 1 9 1 10 9 2
60 15 4 13 1 9 15 4 13 1 15 15 13 9 0 14 13 1 10 9 3 3 7 1 9 13 0 14 13 9 1 15 3 16 15 3 13 16 15 13 11 11 4 13 15 9 1 1 10 9 7 13 0 14 13 15 9 16 13 15 2
12 4 13 2 15 4 13 15 1 9 15 4 2
3 13 15 2
8 15 13 10 0 9 1 11 2
6 15 13 3 10 0 2
32 1 10 11 11 2 11 2 12 11 2 11 14 2 11 2 7 11 1 9 3 2 11 13 10 1 10 0 9 9 1 9 2
18 11 13 10 9 12 9 9 1 11 2 7 13 1 9 7 0 9 2
19 10 11 2 10 11 9 9 2 3 13 10 11 0 12 10 9 2 3 2
44 11 3 13 0 2 9 9 1 9 7 9 2 7 10 0 7 13 2 1 9 1 10 9 13 3 0 1 9 2 9 2 7 3 9 13 14 13 1 10 0 2 0 9 2
25 11 13 3 9 1 9 11 2 11 11 2 11 2 11 11 2 11 11 2 7 10 11 11 11 2
15 15 13 10 0 9 1 11 7 3 13 0 9 10 9 2
10 10 11 1 11 4 3 13 2 3 2
5 11 13 10 9 2
4 4 14 13 2
32 15 9 7 15 4 13 1 1 10 9 1 10 9 1 15 9 1 0 9 15 4 13 3 12 9 7 4 13 1 10 9 2
23 3 15 13 1 10 9 2 16 15 4 13 14 4 16 15 13 10 9 2 2 9 13 2
28 3 2 10 0 9 2 3 15 2 1 0 0 0 9 2 13 14 13 1 10 9 2 15 13 14 13 3 2
54 3 3 10 2 7 15 13 15 2 1 15 9 2 16 15 13 15 9 14 13 1 10 0 9 1 10 9 1 10 9 7 13 10 9 9 16 10 9 13 2 3 16 15 9 13 9 10 0 9 14 13 10 9 2
18 11 13 14 0 2 15 13 14 10 0 9 2 7 10 9 13 0 2
13 14 13 9 1 9 2 15 13 14 13 15 9 2
4 4 14 13 2
11 11 13 10 0 0 9 2 9 5 1 12
9 15 13 15 9 1 11 11 11 2
41 15 13 3 0 9 1 10 9 2 0 9 9 2 1 0 9 7 9 1 0 9 2 0 9 2 7 10 3 2 13 9 9 2 15 13 1 10 9 9 2 2
16 3 2 3 3 2 15 13 10 0 9 2 1 3 0 9 2
5 10 1 10 9 2
32 1 15 15 13 2 10 0 9 1 10 15 9 13 3 1 12 2 9 9 2 0 1 15 13 1 10 0 12 1 11 11 2
31 16 15 13 2 9 13 1 11 2 11 11 2 11 2 11 2 11 7 11 2 11 2 11 2 7 11 11 2 1 9 2
14 0 9 13 1 11 2 13 15 9 2 13 9 9 2
24 10 9 13 2 11 13 15 10 9 14 13 15 1 10 0 9 2 7 15 13 14 13 3 2
9 3 10 0 0 9 1 10 9 2
48 15 4 13 1 10 0 0 9 12 9 13 2 7 15 13 14 13 15 13 12 1 10 0 9 9 15 4 3 13 1 10 9 2 7 15 4 3 13 15 1 10 0 9 15 4 13 1 2
31 10 0 9 1 15 9 7 15 13 3 10 0 9 10 9 1 10 9 2 7 10 9 7 9 4 3 13 12 2 9 2
29 10 9 13 3 0 2 10 9 2 9 13 10 0 9 2 10 9 13 3 0 2 7 10 9 7 9 13 0 2
21 15 13 10 9 3 2 9 9 2 1 10 0 9 2 7 10 9 1 10 9 2
25 10 9 13 3 3 13 2 7 10 9 13 3 0 2 15 13 3 3 16 13 9 10 9 2 5
20 15 3 4 14 13 3 1 10 9 2 15 13 3 10 0 9 0 13 1 2
6 15 9 0 9 1 11
17 15 4 4 13 0 1 10 0 9 2 9 3 1 1 0 9 2
42 15 13 0 9 2 9 2 6 6 15 13 10 9 7 4 14 13 13 3 2 15 13 3 3 3 3 10 9 7 3 15 13 1 10 9 1 10 0 9 7 9 2
7 10 9 13 0 7 0 2
13 15 4 14 13 10 0 11 7 0 14 13 3 2
27 15 13 9 3 3 2 15 4 14 13 15 9 10 13 10 9 15 13 15 2 7 10 9 13 3 0 2
27 15 13 10 0 9 9 1 15 9 1 9 2 9 2 9 2 7 9 7 9 7 0 9 7 13 9 2
6 7 15 9 13 0 2
19 15 4 14 13 3 0 10 9 7 9 9 7 10 9 13 14 13 1 2
12 13 3 7 13 10 9 15 4 14 13 15 2
10 10 9 1 9 1 11 11 1 11 2
3 3 0 2
20 15 4 4 13 1 11 11 1 10 9 1 9 7 4 3 13 15 1 9 2
71 15 4 13 10 1 10 9 3 7 4 13 14 13 16 6 2 1 10 0 9 14 9 15 13 3 10 9 2 13 16 15 0 9 4 4 13 1 2 7 10 1 10 9 7 9 10 4 13 4 13 0 2 3 16 15 4 13 1 10 0 0 9 3 16 15 4 14 13 9 2 2
22 15 4 13 0 1 10 9 1 10 9 7 4 14 3 4 13 9 1 9 7 9 2
39 15 4 14 13 1 15 7 10 9 7 9 15 13 13 3 1 10 0 9 1 15 2 10 9 2 7 15 13 10 9 14 13 9 10 15 13 1 15 2
25 15 3 4 13 0 9 7 16 15 4 3 13 1 10 9 9 2 11 11 13 10 9 1 15 2
5 14 15 15 13 2
24 15 13 10 0 9 16 13 7 13 0 9 2 7 1 15 9 15 4 14 13 1 10 9 2
37 2 15 13 3 12 9 14 4 13 1 15 9 2 16 3 15 13 10 12 9 14 13 15 9 7 10 0 12 9 16 15 9 13 1 15 9 2
66 3 0 1 10 9 10 13 12 9 7 13 3 0 1 10 9 2 6 15 13 10 9 7 9 14 13 15 0 2 16 15 13 1 10 9 15 13 15 9 14 13 1 7 15 13 15 13 1 15 9 7 13 3 14 13 15 7 15 13 0 14 13 9 14 9 2
18 9 13 0 7 10 9 9 13 0 7 10 0 1 10 9 13 0 2
18 1 9 1 15 3 15 13 14 13 15 9 9 3 14 13 15 1 2
17 4 14 13 3 16 15 13 10 9 1 9 10 9 0 7 0 2
9 0 9 2 3 0 2 0 9 2
10 11 11 4 13 10 9 1 15 9 2
22 9 4 13 10 9 9 1 9 7 9 10 15 13 7 13 10 9 16 13 15 13 2
8 10 9 13 3 0 7 0 2
32 15 3 13 16 15 13 9 1 15 9 2 2 1 9 1 15 2 2 15 13 10 9 1 10 9 7 13 0 9 14 13 2
35 15 4 14 3 13 15 9 3 7 13 3 2 7 3 13 9 1 10 0 9 1 10 9 7 3 13 14 13 10 9 16 13 1 9 2
12 10 9 1 9 2 9 7 9 13 0 3 2
18 10 9 15 13 15 13 14 13 10 0 9 7 12 10 13 9 0 2
17 9 4 13 3 0 2 9 13 0 7 10 9 9 13 3 0 2
23 9 13 0 2 2 9 14 9 13 3 12 2 7 11 15 13 9 9 9 2 15 13 2
8 0 9 2 9 2 7 9 9
66 15 13 15 9 7 15 13 10 0 9 9 14 13 10 9 9 3 1 12 13 1 10 9 9 2 7 10 9 13 15 13 10 9 1 11 14 7 3 0 9 13 15 1 1 10 0 0 9 9 2 11 13 1 1 10 9 7 13 0 14 13 10 0 0 9 2
42 3 3 4 15 13 0 2 7 10 9 13 0 2 10 9 13 14 3 0 14 8 13 10 9 2 7 10 9 15 13 3 3 0 2 7 0 2 7 3 0 3 2
40 16 15 4 13 14 13 10 0 1 1 15 9 14 13 3 2 15 4 3 13 15 13 16 16 15 4 13 0 1 15 3 1 15 15 4 3 13 10 9 2
9 2 3 15 13 10 3 0 9 2
16 7 15 13 10 0 9 3 3 2 15 13 0 3 3 2 2
7 15 13 0 12 9 9 2
9 9 9 0 7 9 9 1 9 9
6 15 13 10 9 9 2
20 1 9 2 15 9 9 13 2 1 1 9 2 10 13 15 14 13 13 1 2
22 15 13 10 0 9 1 9 9 2 3 12 5 2 7 9 1 9 1 10 0 9 2
17 15 3 13 12 9 1 15 0 9 7 12 9 1 15 0 9 2
4 15 13 0 2
20 15 13 3 3 1 9 7 15 9 9 13 3 12 5 0 1 3 12 9 2
23 16 13 1 9 9 15 13 10 0 9 1 9 7 3 13 16 15 9 14 9 13 15 2
12 15 13 3 3 2 13 3 1 9 1 9 2
14 15 15 13 3 1 11 11 13 16 15 13 3 0 2
8 15 13 1 15 1 10 9 2
11 15 4 13 15 3 13 7 13 14 13 2
10 15 13 3 0 14 4 13 11 11 2
13 3 15 13 3 0 13 15 9 9 1 10 9 2
4 10 9 1 11
23 1 10 0 9 2 12 0 9 1 9 0 1 10 11 9 9 13 10 0 2 9 9 2
7 11 4 13 10 9 3 2
20 10 9 13 1 10 0 9 9 2 10 13 10 9 3 1 10 11 11 9 2
16 10 9 1 11 13 14 13 9 0 16 13 15 13 3 3 2
9 10 9 4 3 13 10 13 9 2
26 15 13 9 1 9 2 7 15 4 3 13 10 9 1 9 9 15 4 14 13 13 7 13 15 9 2
10 3 1 10 2 15 13 10 9 2 2
7 3 9 7 10 0 9 2
16 13 14 13 0 9 2 7 10 9 15 13 1 10 0 9 2
14 7 16 15 13 13 1 10 9 2 15 4 13 11 2
32 10 9 3 13 10 0 9 1 11 2 15 4 13 10 9 1 10 9 2 7 0 9 4 13 9 16 15 13 10 9 9 2
8 10 0 9 1 10 0 9 2
5 13 15 2 11 2
4 9 9 1 9
8 15 0 9 13 3 0 9 2
13 15 4 4 13 10 9 7 14 13 10 10 9 2
21 15 4 13 9 9 7 13 3 10 0 9 1 9 7 13 0 0 9 3 3 2
22 15 13 10 9 14 9 9 7 16 13 10 9 9 15 4 13 7 13 1 0 9 2
11 10 9 2 11 2 4 13 3 12 9 2
4 10 10 9 2
19 15 13 10 3 0 2 0 7 3 2 13 9 1 10 0 9 1 9 2
25 15 3 13 13 15 7 0 14 13 15 13 1 11 7 13 10 9 1 10 0 10 9 9 9 2
19 10 9 13 10 0 9 7 13 0 14 13 10 0 9 7 10 0 9 2
37 1 10 9 2 11 2 10 9 9 2 13 9 1 9 2 9 2 0 2 9 2 13 9 2 0 9 2 9 2 10 9 1 0 9 1 9 2
7 0 9 1 10 0 9 2
3 13 3 2
3 11 11 12
6 10 12 11 13 0 2
13 15 13 10 0 9 1 10 3 0 12 11 11 2
32 15 4 3 13 10 9 3 16 10 9 1 11 11 13 15 7 15 13 15 15 13 15 3 7 16 9 13 3 0 1 15 2
18 15 13 15 15 15 13 1 7 15 3 13 15 15 13 10 9 9 2
40 15 13 10 9 1 7 13 3 7 13 1 10 9 15 13 11 7 15 13 15 3 3 3 13 15 9 2 15 13 10 9 0 16 9 4 13 3 0 9 2
39 15 13 16 13 7 15 13 15 13 1 7 15 9 13 1 11 7 15 13 9 1 9 1 10 9 10 15 13 13 2 2 13 15 13 14 13 15 2 2
24 15 13 15 4 13 1 1 15 9 9 7 15 3 13 1 15 7 3 15 4 4 13 0 2
19 11 7 11 13 3 0 16 15 15 13 7 13 3 3 14 13 10 9 2
5 3 13 13 15 2
6 9 7 9 2 0 9
49 13 10 11 9 12 9 3 2 16 15 13 1 12 0 9 1 0 9 2 4 13 15 4 13 10 2 0 9 9 9 2 14 13 9 7 13 10 0 2 13 2 9 2 0 1 9 9 2 2
12 4 13 5 12 3 0 1 9 9 2 8 2
11 10 9 2 13 16 15 4 13 10 9 2
4 4 13 0 2
34 13 10 9 13 1 2 13 9 2 3 3 3 3 10 9 4 14 13 10 13 9 7 15 13 5 12 7 3 5 12 1 10 9 2
17 15 4 13 10 9 1 3 5 12 10 4 13 15 10 13 9 2
8 3 1 5 12 1 5 12 2
4 13 15 0 2
31 15 13 16 15 4 14 13 15 10 9 16 15 13 3 10 9 7 3 16 15 13 10 0 9 15 13 12 9 10 9 2
22 7 10 9 4 14 13 9 16 15 15 4 13 2 7 0 2 15 4 13 7 13 2
10 15 13 10 0 9 13 1 10 9 2
35 3 16 9 13 1 10 9 2 3 1 9 9 2 10 11 11 13 14 0 7 15 13 3 0 1 10 1 10 9 9 15 4 13 1 2
13 6 2 15 13 0 2 7 0 13 14 3 0 2
49 15 13 15 1 10 13 7 13 9 2 13 3 1 10 9 14 9 1 0 9 3 7 13 3 3 13 2 0 9 1 0 9 9 2 15 4 3 13 15 3 2 1 12 0 0 9 9 2 2
19 10 9 13 3 0 7 15 4 13 15 9 1 10 11 11 1 10 9 2
24 4 14 13 3 16 15 13 15 9 1 15 0 9 7 13 15 3 3 7 1 15 0 9 2
45 16 15 9 1 10 9 2 3 4 15 13 15 9 13 2 2 13 14 13 2 2 1 10 9 9 1 11 2 2 15 4 3 13 10 9 3 13 2 2 1 10 11 11 2 2
3 13 15 2
23 15 3 13 10 9 9 1 10 9 7 15 13 0 16 3 3 11 7 15 9 4 13 2
14 15 13 1 10 9 14 13 16 15 9 9 4 13 2
39 15 13 14 13 15 1 10 9 1 12 9 7 15 4 13 14 13 1 9 9 3 3 16 15 13 16 3 3 3 0 9 15 13 15 4 14 13 15 2
18 6 15 13 3 0 1 15 7 13 15 1 9 3 13 9 1 9 2
23 1 10 9 15 13 0 14 13 3 0 9 15 13 2 3 10 9 1 13 14 13 9 2
23 15 4 3 13 15 13 15 10 9 14 13 1 15 16 3 10 9 1 10 9 13 0 2
14 15 4 3 13 1 10 9 3 3 16 15 13 9 2
18 15 13 3 12 9 3 7 7 15 4 3 13 10 9 14 13 15 2
23 1 9 15 13 3 16 13 15 9 1 10 9 3 1 16 3 15 9 7 15 4 13 2
7 6 2 3 13 10 9 2
8 15 13 10 9 1 10 11 2
10 10 9 13 0 2 10 9 13 0 2
24 15 13 15 13 3 1 10 9 16 3 15 13 3 9 13 3 7 13 2 3 1 10 9 2
15 1 15 9 10 9 4 13 0 2 1 10 0 9 2 2
50 3 2 10 9 2 9 3 13 14 4 13 2 16 15 3 13 10 14 13 1 2 7 13 12 9 2 3 13 1 9 3 0 9 4 14 3 13 7 14 13 3 3 3 14 13 16 9 4 13 2
23 1 10 9 10 9 13 1 1 9 2 1 10 9 10 9 3 4 14 13 2 13 3 2
26 15 4 3 13 9 14 13 9 2 9 0 2 16 15 13 14 9 9 3 3 3 15 13 15 3 2
14 15 3 13 14 13 15 15 4 13 1 3 15 13 2
24 0 0 9 2 0 9 2 3 9 2 2 7 4 14 13 16 15 13 10 0 9 1 9 2
4 13 10 11 9
25 15 3 13 10 11 9 1 10 15 9 2 15 4 4 13 3 1 9 7 4 3 13 3 3 2
18 10 9 13 3 0 7 3 13 1 10 9 9 3 1 13 15 9 2
29 15 13 3 10 3 0 9 7 15 13 9 0 7 10 9 1 9 4 3 13 0 15 13 3 1 10 0 9 2
20 15 13 1 10 1 10 0 9 7 13 16 9 13 16 10 9 13 1 15 2
8 1 10 9 1 10 9 9 2
27 11 13 10 3 0 9 9 1 9 7 15 13 15 16 15 13 15 15 13 0 3 8 3 15 13 0 2
25 3 15 4 13 3 10 9 13 7 13 15 13 3 1 10 0 9 7 14 13 15 1 10 9 2
22 15 4 13 13 1 11 1 11 16 15 13 12 1 10 3 0 9 9 1 10 9 2
22 3 13 15 9 13 1 15 13 14 13 10 0 7 10 11 13 3 9 15 4 13 2
53 15 13 14 13 10 9 0 9 16 15 13 16 15 13 10 0 9 1 10 9 3 1 10 0 9 2 0 9 9 2 1 9 9 1 9 9 2 9 9 2 7 9 1 15 13 3 0 7 0 10 9 9 2
32 3 15 13 10 11 11 9 2 0 9 7 9 9 2 7 0 9 9 9 2 5 12 2 5 12 2 7 5 12 3 2 2
41 10 0 9 9 9 13 3 10 0 9 2 0 7 0 2 10 0 9 15 13 10 15 4 13 13 3 0 15 7 10 0 9 2 7 15 3 13 0 9 2 2
14 10 0 9 13 14 3 3 0 2 3 13 15 9 2
17 10 0 9 13 16 10 9 13 14 0 7 13 3 0 2 0 2
25 10 9 13 0 2 10 9 13 0 7 0 1 10 1 2 1 2 9 0 2 9 9 13 9 2
11 7 15 4 13 3 16 10 9 4 13 2
7 15 13 3 14 0 15 2
6 4 14 13 9 7 9
13 15 4 13 1 12 9 1 10 9 1 11 12 2
19 1 12 9 1 9 9 12 2 10 9 9 7 9 9 13 1 15 9 2
7 15 13 14 9 9 9 2
14 3 15 13 1 2 15 13 10 0 0 2 0 9 2
10 15 13 10 0 9 7 13 10 9 2
21 16 13 1 9 1 9 7 9 7 13 9 2 15 13 14 3 13 1 7 13 2
27 10 9 9 3 13 1 15 2 13 16 10 0 9 4 13 1 2 16 16 15 4 13 15 1 2 2 2
27 15 3 13 16 3 10 12 9 9 9 4 13 2 3 3 12 9 4 13 2 10 0 9 1 15 2 2
28 10 0 9 13 10 9 3 2 7 3 13 14 13 15 10 9 1 10 9 16 15 13 15 1 15 12 9 2
18 10 9 13 0 0 2 7 15 13 10 0 9 1 10 9 7 9 2
13 4 14 13 3 16 15 13 14 13 1 10 9 2
10 0 9 2 9 1 9 2 4 14 13
33 15 13 13 11 11 3 1 12 7 4 13 10 0 9 1 10 9 1 9 2 9 2 9 9 2 7 3 10 0 9 1 9 2
26 10 0 9 13 1 10 9 9 2 3 10 9 13 3 0 7 13 10 9 15 3 13 1 10 9 2
49 15 13 15 3 12 9 14 13 10 0 9 2 7 0 9 1 15 9 1 1 15 9 1 9 7 9 2 14 16 15 13 10 9 1 10 9 2 7 15 13 14 3 3 13 14 13 0 2 2
49 3 2 15 4 13 14 13 15 9 9 13 1 15 2 7 15 3 13 2 7 1 10 0 9 14 13 11 11 1 10 9 14 13 15 1 15 9 2 15 3 13 1 7 13 1 10 0 9 2
20 6 4 14 13 3 16 15 13 0 2 0 2 0 0 9 15 4 13 1 2
17 13 15 10 9 2 9 7 9 7 13 10 3 0 9 2 9 2
21 10 9 9 4 3 13 1 11 2 7 13 3 1 11 2 11 2 13 11 11 2
39 3 10 9 13 2 12 9 3 16 13 2 15 13 16 15 13 14 13 10 10 9 15 13 13 1 11 7 0 5 12 16 15 14 13 3 1 15 9 2
13 15 13 14 1 9 3 2 7 15 3 13 15 2
9 7 10 5 12 16 13 10 9 2
12 3 13 5 12 3 1 9 16 10 9 13 2
12 13 15 2 13 14 1 10 0 9 3 3 2
30 15 4 13 1 1 12 9 9 7 15 13 1 12 0 9 12 9 14 13 10 9 2 1 12 9 5 12 9 2 2
22 10 0 9 15 4 13 12 9 3 1 12 7 12 2 15 4 13 2 9 4 13 2
18 3 15 3 4 13 15 7 13 13 3 3 0 16 15 13 15 3 2
14 12 0 9 2 15 4 14 13 10 9 9 7 9 2
15 15 13 14 13 9 3 16 15 13 13 9 1 15 9 2
3 0 9 3
15 15 13 3 1 12 9 2 10 0 9 7 3 13 0 2
16 3 2 10 0 9 15 13 1 11 2 10 0 10 9 13 2
28 15 4 3 13 15 9 13 1 2 15 13 3 9 13 9 1 10 9 2 3 16 15 4 13 14 4 13 2
36 10 9 4 13 14 13 1 12 7 15 4 13 9 3 3 1 12 13 2 13 9 7 13 15 2 13 2 15 1 10 0 9 1 10 9 2
55 3 2 3 15 13 1 2 15 13 10 9 9 1 9 2 15 13 3 7 13 14 13 15 1 12 9 9 2 7 15 3 13 15 9 3 2 7 0 9 2 10 4 3 13 2 15 13 9 9 7 9 1 15 2 2
39 11 13 10 0 9 15 4 3 13 1 7 15 13 1 1 10 1 10 0 2 0 9 10 13 3 2 3 10 0 9 10 3 13 10 9 16 13 9 2
10 4 14 13 3 2 15 4 13 15 2
5 10 0 9 3 2
20 15 4 13 1 11 11 1 11 7 11 2 7 15 13 1 1 10 0 9 2
37 15 4 13 1 15 1 10 9 2 15 4 14 13 10 0 9 1 11 2 7 13 16 11 13 0 14 13 1 1 15 9 1 9 1 10 9 2
10 15 13 15 4 13 10 9 10 9 2
26 3 2 16 13 10 13 5 12 2 8 0 2 9 16 13 10 9 7 9 2 15 13 0 15 13 2
12 15 13 10 9 1 9 3 2 11 13 0 2
18 15 13 9 9 2 7 9 1 9 3 2 10 10 13 3 1 9 2
22 1 10 9 15 13 1 10 9 15 13 15 15 4 13 1 2 15 13 3 10 9 2
8 3 9 7 10 9 1 9 2
4 15 13 10 2
13 10 9 13 3 3 0 1 9 14 13 1 15 2
23 6 9 2 13 9 7 4 14 4 13 1 1 10 9 16 11 7 11 13 1 10 9 2
15 15 13 3 10 9 16 15 14 13 15 9 1 15 0 9
2 0 2
2 0 2
28 3 15 13 3 2 10 9 1 9 13 2 2 6 6 2 15 4 13 2 15 13 1 10 9 1 9 2 2
16 1 10 0 0 9 2 15 13 2 2 15 4 15 13 2 2
11 3 1 1 15 9 15 13 16 15 13 2
9 15 13 16 10 9 13 9 9 2
15 15 3 13 2 6 2 15 13 10 5 12 9 3 2 2
10 3 3 15 13 15 1 10 9 9 2
22 3 15 13 15 3 13 2 1 10 9 3 9 4 13 1 15 4 13 15 3 2 2
23 15 13 9 9 1 15 16 10 9 3 13 16 15 13 10 0 9 1 10 9 2 9 2
8 15 3 13 1 10 9 9 2
12 15 13 2 15 13 9 1 2 9 2 2 2
8 13 10 9 13 9 1 9 2
8 15 3 13 15 1 15 9 2
11 15 13 15 4 13 10 0 7 0 9 2
17 15 13 10 9 16 14 13 7 4 13 15 3 3 16 15 4 2
5 4 14 13 3 2
13 15 13 14 13 1 10 9 13 10 9 9 3 2
20 15 9 7 15 13 14 13 3 1 10 9 9 2 13 1 1 15 9 9 2
20 15 13 1 12 9 1 10 9 7 13 14 13 3 1 15 9 1 10 9 2
23 3 15 9 7 15 13 14 13 15 12 9 0 9 1 10 9 7 15 4 14 13 15 2
16 15 9 13 10 9 14 13 15 9 3 3 16 15 13 15 2
22 15 13 16 15 13 14 4 13 1 10 9 3 16 15 4 14 13 1 10 12 9 2
19 15 13 15 3 10 0 9 16 13 15 11 1 7 15 3 4 14 13 2
13 9 13 0 2 15 13 2 7 15 13 10 9 2
15 15 13 12 9 14 13 1 10 9 2 3 10 9 3 2
9 15 13 12 9 2 3 10 9 2
23 1 12 1 10 9 15 13 10 9 1 10 9 14 10 13 15 9 2 10 9 13 9 2
8 15 3 13 11 11 7 9 2
30 15 13 0 15 13 10 0 9 14 13 16 13 10 0 9 2 7 16 9 0 13 1 15 9 2 15 4 14 13 2
1 0
17 6 15 13 10 11 11 15 4 4 13 1 9 1 11 2 11 2
13 15 13 10 11 13 3 0 1 0 11 9 9 2
25 15 13 14 13 10 0 9 10 0 9 13 1 10 0 9 2 7 15 13 14 13 10 0 9 2
14 15 13 15 4 13 14 13 16 15 13 3 1 11 2
14 6 3 15 13 1 10 9 1 11 7 4 13 3 2
12 15 13 10 9 7 15 13 1 10 0 9 2
28 15 13 15 4 13 10 0 9 2 0 9 2 13 1 10 9 2 16 10 9 13 1 10 9 1 10 9 2
9 15 13 13 0 9 9 7 9 2
6 3 15 13 10 9 2
9 15 13 16 15 3 13 3 3 2
19 15 4 14 13 3 15 13 15 2 7 0 9 2 15 13 10 0 9 2
19 15 13 10 9 16 13 10 9 16 13 11 9 16 10 11 3 13 15 2
14 15 4 13 2 15 4 14 13 3 15 9 9 13 2
23 15 4 13 14 13 10 9 14 13 10 9 9 1 10 9 2 11 11 13 0 1 15 2
9 0 9 2 0 9 9 2 0 9
20 15 13 1 12 1 9 15 13 10 9 9 1 10 11 11 14 1 11 11 2
11 10 9 13 0 2 7 3 13 15 9 2
42 3 15 13 9 14 13 10 9 3 3 2 15 4 14 13 15 13 10 1 10 9 1 10 9 2 10 15 4 13 1 10 0 9 15 4 13 10 9 9 1 2 2
12 15 3 13 16 15 4 13 9 3 1 9 2
25 10 9 13 14 13 13 1 10 9 2 15 4 13 1 10 9 13 1 15 9 15 4 13 3 2
9 15 9 13 0 7 9 3 0 2
6 0 16 13 15 13 2
18 10 9 13 3 0 2 0 7 13 15 13 16 15 4 13 15 9 2
39 15 13 10 0 9 0 2 15 3 13 15 9 9 14 13 10 9 9 2 7 15 13 15 1 7 13 15 1 10 9 9 16 13 15 1 10 9 9 2
10 15 4 14 4 13 11 11 14 3 2
19 15 13 0 9 1 9 3 3 0 1 9 10 13 9 7 9 3 3 2
4 13 1 11 11
16 11 11 13 3 0 9 2 16 10 9 13 3 1 10 9 2
6 15 13 3 0 9 2
14 1 10 0 9 10 9 9 13 14 0 7 0 9 2
12 3 2 15 4 14 13 9 3 1 10 9 2
13 3 2 15 4 3 13 12 9 13 15 15 9 2
21 15 13 14 10 0 9 7 15 13 14 13 15 9 3 16 15 13 14 13 15 2
20 15 13 14 13 10 9 15 13 15 9 7 15 3 13 3 14 13 15 13 2
8 15 13 14 13 1 15 9 2
22 3 15 3 13 3 10 9 13 14 3 0 2 15 13 3 10 9 1 9 13 3 2
9 15 13 3 1 11 9 2 12 2
23 15 13 3 3 1 11 9 12 2 3 15 9 14 11 9 13 3 16 10 9 1 15 2
34 10 9 13 3 7 13 15 13 0 7 13 10 0 9 1 9 2 15 13 15 4 14 3 13 9 16 10 9 4 3 13 7 13 2
17 1 15 9 4 4 3 13 1 10 9 1 10 9 1 10 9 2
7 7 9 13 15 0 9 2
4 9 9 3 2
11 15 9 9 13 3 0 1 10 9 9 2
16 15 13 1 10 9 9 2 7 15 3 13 9 7 9 3 2
14 15 13 16 15 13 0 3 2 7 15 13 3 14 2
25 3 2 15 4 13 15 3 1 9 2 7 3 13 14 13 1 15 9 2 7 13 15 13 2 2
19 15 13 1 1 10 9 9 2 16 15 4 13 0 9 16 15 4 13 2
22 15 3 13 12 9 1 10 9 9 2 16 15 13 14 13 0 0 9 1 10 9 2
15 15 9 13 10 9 0 1 15 2 7 15 13 3 0 2
19 15 13 10 0 9 3 15 13 10 9 1 9 1 9 1 5 12 0 2
11 3 2 10 9 9 2 15 4 13 15 2
14 15 13 15 3 12 9 7 15 13 13 9 1 9 2
17 2 9 2 13 1 9 1 11 11 2 15 4 13 9 13 3 2
21 15 13 3 1 12 7 12 7 15 4 14 13 3 0 9 15 4 13 15 13 2
19 3 15 4 14 13 3 2 7 10 9 1 10 9 9 3 13 10 9 2
19 15 12 9 2 9 4 13 0 1 12 9 3 15 13 9 1 10 9 2
15 15 13 15 9 7 9 3 14 13 1 10 0 12 11 2
19 11 11 13 3 0 7 0 1 15 9 7 15 13 15 13 13 15 1 2
11 15 13 3 3 10 9 7 13 1 11 2
16 15 13 15 10 9 15 13 0 1 7 15 13 10 9 9 2
20 15 13 10 9 3 15 13 13 15 9 2 9 7 10 9 1 10 12 11 2
8 10 0 9 13 3 12 9 2
25 0 9 7 9 1 10 9 16 15 13 1 10 9 10 13 1 15 9 7 13 0 1 10 9 2
16 12 9 1 9 7 15 13 10 9 1 10 0 0 12 11 2
39 15 4 13 3 12 9 2 9 2 9 2 7 9 2 1 15 9 7 15 13 14 13 10 9 1 11 7 11 11 11 1 11 11 13 12 1 10 0 2
9 0 2 0 2 7 1 10 0 2
19 15 13 10 15 4 3 13 1 10 9 9 7 11 7 11 13 10 12 2
10 9 1 10 0 9 7 10 0 9 2
2 9 9
13 15 7 15 9 14 9 4 13 1 10 9 9 2
16 15 4 13 1 10 9 7 13 14 13 15 9 1 9 0 2
12 3 15 13 10 9 16 15 13 12 1 15 2
13 15 13 10 0 9 10 13 14 13 1 10 9 2
16 15 13 10 9 7 13 15 1 10 9 10 13 10 10 9 2
23 10 0 9 4 13 3 12 9 7 10 9 13 0 9 1 9 7 0 9 9 1 15 2
7 15 13 3 15 4 13 2
17 15 10 13 1 9 7 10 0 9 4 13 1 9 1 10 9 2
12 10 9 1 1 15 13 1 10 9 1 9 2
4 9 13 3 2
17 10 9 4 13 1 2 3 10 9 1 10 0 9 4 13 1 2
12 0 9 3 10 9 4 13 2 3 10 9 2
6 15 9 13 3 0 2
12 15 13 1 12 10 4 14 13 10 9 9 2
11 9 9 13 3 0 0 1 10 11 11 2
6 15 13 13 10 9 2
13 16 15 13 10 9 2 15 4 14 13 1 15 2
10 9 13 12 5 1 10 9 3 3 2
10 9 13 10 0 9 2 9 3 0 2
7 10 0 15 13 1 9 2
26 15 4 3 13 1 11 2 11 1 11 1 15 12 0 9 7 13 10 9 1 10 9 9 1 11 2
19 15 13 12 3 10 9 13 15 14 13 11 2 15 4 13 9 1 15 2
19 3 3 4 15 13 10 9 1 12 1 10 11 2 15 13 10 9 13 2
59 15 13 1 10 0 9 10 13 15 11 11 1 11 1 9 7 13 15 2 3 15 13 3 2 13 1 15 9 2 15 13 10 9 2 7 9 4 14 13 15 10 0 16 15 13 1 2 2 7 13 15 1 15 9 14 13 10 9 2
23 15 13 3 3 13 3 3 1 1 11 15 13 7 13 15 1 15 9 1 12 10 9 2
17 9 11 1 10 1 15 9 7 13 9 3 1 15 9 10 9 2
44 15 13 1 10 9 2 10 0 9 9 15 4 3 13 7 3 14 13 0 2 10 9 15 13 15 13 10 0 1 15 9 9 1 11 14 9 16 13 1 10 0 0 9 2
11 15 13 15 4 13 10 9 1 10 9 2
2 11 11
3 9 0 2
7 9 7 9 9 14 0 2
40 15 4 13 1 10 9 0 9 2 7 16 15 3 13 10 0 9 1 10 9 2 15 9 9 3 13 1 0 9 7 9 1 10 0 2 3 3 0 9 2
85 15 4 3 13 15 10 0 9 16 15 13 1 9 7 4 13 1 15 2 7 3 15 13 14 13 1 10 2 0 2 0 9 10 13 1 12 9 1 12 9 1 15 0 9 7 15 13 1 16 10 0 9 13 0 1 9 9 2 15 9 13 14 7 13 9 9 9 16 13 1 10 3 0 9 9 1 10 9 2 7 3 13 1 15 2
39 15 13 10 0 2 7 13 10 0 9 1 10 9 9 14 13 1 15 9 1 0 9 2 3 14 13 10 0 9 14 9 15 13 1 7 4 14 13 2
15 15 4 13 9 4 13 15 1 7 3 13 1 10 9 2
40 15 4 3 13 3 3 16 15 13 0 7 15 4 14 13 10 0 9 2 7 4 14 13 3 1 15 7 4 3 14 13 10 9 1 9 7 0 0 9 2
48 13 3 10 0 9 7 10 9 1 10 9 13 1 15 7 15 9 16 15 13 15 13 10 9 9 1 10 9 10 0 3 3 7 10 9 4 3 13 1 7 10 9 13 3 1 10 9 2
45 15 13 14 13 10 9 1 10 9 7 13 15 1 10 9 16 13 1 15 13 2 2 15 4 14 13 15 15 4 14 13 1 2 7 2 15 4 14 13 3 9 4 13 2 2
19 15 13 3 0 14 13 10 9 1 9 3 1 9 1 15 12 9 0 2
26 15 13 1 10 9 16 13 15 10 9 7 3 15 13 3 2 10 9 13 10 0 15 4 3 13 2
10 9 4 13 3 2 3 0 7 0 2
30 15 13 15 13 15 1 9 1 1 15 0 9 1 10 9 1 9 10 13 14 3 3 2 0 2 3 2 0 2 2
34 15 4 3 13 3 1 10 9 7 15 4 13 15 1 10 0 9 9 1 0 0 9 9 7 3 13 15 9 7 13 15 5 12 2
7 10 9 13 12 5 0 2
13 10 0 9 15 13 15 13 9 4 13 15 9 2
11 0 9 2 0 9 2 0 9 2 0 9
27 10 0 9 15 13 3 15 13 1 9 13 16 10 9 9 3 13 1 10 9 7 13 1 10 9 9 2
21 10 9 1 10 0 9 0 14 13 1 9 3 14 13 9 4 13 0 2 6 2
22 15 13 2 15 13 10 9 15 13 1 9 9 2 10 0 9 13 1 10 0 9 2
8 6 2 15 4 13 10 9 2
24 10 9 13 15 9 7 2 13 2 1 15 13 3 0 7 13 10 9 1 9 9 3 3 2
15 15 4 13 0 9 13 1 11 9 9 1 1 10 9 2
25 7 4 14 3 13 16 13 14 13 1 10 9 16 10 9 13 2 7 13 15 11 2 10 9 2
49 16 15 4 13 1 9 2 13 1 10 0 9 7 16 15 13 10 0 9 2 15 4 3 13 1 15 15 13 1 2 10 9 10 13 2 0 2 2 7 3 3 0 13 1 1 10 10 9 2
11 13 15 10 9 7 13 10 9 8 3 2
23 15 13 15 13 3 1 13 11 7 13 11 10 9 1 9 1 10 9 7 3 11 11 2
6 13 15 13 1 11 2
38 15 4 13 1 11 11 1 9 2 0 9 15 13 14 13 10 11 11 7 13 10 9 2 7 13 1 11 2 11 2 11 11 10 9 1 10 9 2
8 15 13 0 9 7 9 9 2
24 15 13 0 0 2 10 9 13 0 2 4 14 4 13 1 1 10 12 0 9 1 10 9 2
29 15 4 13 15 15 4 3 13 2 11 13 9 9 7 10 9 3 10 9 13 3 0 2 0 9 2 13 0 2
15 15 9 13 10 9 9 7 13 0 9 9 7 0 9 2
8 10 9 13 15 15 4 13 2
10 13 15 7 13 2 15 4 13 3 2
18 15 13 10 9 9 1 9 11 11 7 13 10 9 13 1 15 9 2
20 10 0 9 13 15 0 16 10 0 9 14 13 15 0 9 9 1 0 9 2
3 1 11 2
45 15 3 13 10 9 1 14 13 15 2 7 10 0 9 15 13 2 15 13 10 9 16 13 15 9 9 14 13 15 9 7 15 1 10 9 14 13 15 3 3 0 15 9 13 2
7 4 14 13 14 13 3 2
4 2 11 11 2
8 15 13 16 15 13 3 0 2
28 3 1 10 2 16 15 13 1 10 9 15 4 14 13 15 14 13 3 10 9 3 16 15 4 3 13 12 2
25 15 3 4 14 13 15 16 15 4 13 14 13 15 10 2 9 2 14 4 13 14 13 10 9 2
33 15 13 16 10 9 10 9 14 9 13 1 3 13 10 0 9 0 3 15 13 0 16 10 9 4 14 13 10 12 9 1 0 2
14 3 15 4 4 13 10 0 9 7 3 10 13 9 2
37 10 9 4 13 15 16 15 0 9 9 13 1 1 15 9 14 9 16 10 9 4 3 13 1 1 0 9 7 15 13 10 0 9 2 8 2 2
13 1 0 15 4 13 16 10 9 13 0 7 0 2
15 7 3 3 15 13 0 1 15 3 15 4 4 13 3 2
21 6 2 16 13 10 1 10 0 9 15 13 16 10 1 10 0 9 4 13 9 2
13 16 15 13 9 15 4 13 14 13 1 11 11 2
17 15 13 10 3 0 0 9 9 7 1 10 9 15 13 3 0 2
14 15 4 14 13 0 9 10 13 3 0 1 0 9 2
4 0 9 1 11
14 15 3 13 1 11 1 9 7 13 10 3 0 9 2
32 15 13 1 10 0 9 9 3 13 15 9 1 11 7 13 14 13 14 13 10 1 15 9 9 9 4 13 3 7 1 9 2
20 15 4 13 14 13 10 0 9 1 15 13 3 13 13 9 1 10 0 9 2
24 15 13 3 0 14 13 15 9 7 10 9 9 14 13 10 3 0 7 0 9 1 15 9 2
20 15 13 10 9 14 13 3 0 2 3 14 13 3 3 13 1 0 0 9 2
23 1 15 0 9 1 9 9 1 15 0 9 9 15 13 10 9 7 9 14 13 15 9 2
26 15 3 13 15 0 13 1 9 7 13 0 1 10 9 7 9 1 10 9 3 3 1 10 9 15 2
34 15 4 4 13 1 10 9 1 10 9 7 15 4 4 13 16 10 9 4 13 0 1 15 9 1 9 7 11 4 13 15 0 9 2
19 6 10 9 4 13 10 9 7 13 1 11 15 13 10 9 1 0 9 2
25 6 13 15 9 1 10 9 7 9 1 15 0 9 7 0 9 16 15 13 13 10 0 9 0 2
5 0 9 1 11 2
10 9 2 15 13 14 13 1 15 9 2
18 15 13 3 3 0 9 7 13 10 9 14 13 1 15 0 9 9 2
2 0 2
14 15 13 10 9 1 10 0 9 7 3 3 1 9 2
37 6 15 13 1 1 10 9 3 15 4 13 1 10 0 9 1 10 9 15 13 16 15 9 7 15 4 13 14 13 1 15 2 0 2 9 9 2
21 3 3 15 13 15 16 15 13 10 0 0 9 1 10 0 9 3 3 15 13 2
8 15 4 13 3 7 13 3 2
23 16 13 1 10 9 7 13 10 0 9 9 15 13 2 15 13 15 13 1 1 10 9 2
15 15 13 10 9 9 9 7 15 9 13 10 9 9 9 2
2 0 2
12 10 9 13 0 3 16 15 3 13 10 3 2
13 15 13 14 13 10 9 1 10 9 3 13 15 2
36 15 13 0 14 13 16 3 1 10 9 15 4 13 10 9 10 13 0 9 2 0 9 2 7 0 9 2 7 14 13 10 9 16 13 15 2
31 0 9 13 16 3 15 13 10 0 3 13 9 16 15 13 15 4 13 16 10 9 7 9 13 9 1 15 9 7 9 2
3 3 13 2
6 0 9 7 0 9 2
32 15 3 13 9 13 1 15 11 1 10 9 2 7 15 13 12 9 0 3 7 4 13 9 9 3 4 14 13 9 0 3 2
18 15 4 13 1 0 9 1 10 9 7 4 4 13 1 10 0 9 2
19 15 4 13 0 9 1 11 7 11 11 3 15 13 14 13 15 10 9 2
7 10 9 13 0 7 0 2
26 15 13 1 15 15 13 14 13 13 13 15 15 13 4 13 16 15 13 10 9 7 13 0 9 9 2
36 10 9 13 3 0 16 15 15 4 13 7 0 1 13 1 0 9 2 7 15 13 15 10 9 15 13 3 15 13 3 14 13 1 10 9 2
46 3 2 10 9 1 10 9 2 11 13 15 1 14 13 3 15 9 4 13 7 14 13 15 13 16 15 4 3 13 15 1 9 1 10 9 7 13 14 13 15 10 9 1 10 9 2
8 15 13 3 0 3 10 9 2
42 15 13 1 1 10 0 9 3 15 13 7 13 15 9 7 13 3 0 1 9 1 9 9 16 15 13 3 2 7 11 4 13 16 15 3 13 0 3 13 9 3 2
7 15 13 15 9 13 3 2
21 15 9 13 10 0 9 9 9 7 9 9 9 2 3 15 13 3 10 9 9 2
23 15 4 4 13 9 9 1 10 10 9 7 3 13 14 13 10 9 1 11 2 7 11 2
10 15 13 10 9 1 10 9 1 9 2
5 8 2 0 9 2
27 15 13 0 1 9 9 9 9 2 7 13 9 1 0 9 2 15 3 13 16 15 13 10 0 0 9 2
26 8 2 15 3 13 10 9 16 11 13 13 9 7 15 13 3 10 9 14 13 1 15 0 9 9 2
7 3 4 15 13 3 3 2
59 6 15 4 4 13 1 11 1 12 9 2 7 13 12 9 13 15 9 1 11 2 7 15 9 9 2 8 4 13 10 12 9 9 1 9 2 10 4 3 13 15 9 2 9 13 10 9 10 13 9 7 14 13 9 3 3 13 0 2
30 15 13 3 0 16 11 14 0 7 13 9 4 13 10 9 13 14 13 2 7 15 9 4 13 10 9 1 10 9 2
37 3 2 15 4 4 13 16 11 13 10 0 9 14 13 1 2 1 1 15 0 9 7 3 1 3 16 15 13 10 3 0 9 7 10 0 9 2
4 0 9 7 9
18 15 13 11 2 11 13 0 1 10 9 1 15 11 9 12 9 3 2
20 10 0 9 4 13 1 10 9 2 7 15 13 14 3 15 4 13 15 9 2
16 12 9 3 2 9 13 14 13 9 1 10 9 1 15 9 2
9 10 9 13 10 9 1 10 9 2
22 3 2 15 13 14 13 10 9 1 10 9 9 7 3 14 13 10 9 1 10 9 2
6 10 9 4 14 13 2
30 15 0 2 9 9 13 10 9 7 13 1 10 9 2 3 13 10 12 9 3 2 15 3 13 15 9 3 2 2 2
47 15 13 11 2 11 10 0 9 14 13 10 9 9 1 10 9 2 7 4 3 13 3 15 13 16 15 4 14 3 13 14 13 15 1 10 9 9 2 16 15 4 4 13 1 15 9 2
24 6 7 6 2 15 13 10 9 2 10 13 14 4 13 2 9 7 4 14 13 15 10 9 2
15 15 9 3 13 12 1 15 9 7 13 10 9 1 15 2
25 1 10 9 7 9 2 15 13 3 0 14 13 10 9 1 0 0 9 7 0 3 13 9 9 2
17 15 3 13 9 0 1 10 9 2 7 15 3 13 9 14 9 2
7 0 3 2 7 3 10 9
4 11 2 12 2
19 15 4 13 1 10 11 1 10 9 1 0 1 2 1 2 9 9 9 2
32 13 13 1 10 0 9 10 0 9 2 7 13 3 0 14 13 9 1 10 0 9 9 13 14 13 1 10 9 1 12 9 2
17 0 9 4 13 1 10 9 2 1 10 0 9 1 0 9 9 2
19 15 13 12 9 1 15 9 7 9 1 3 12 2 10 9 1 9 9 2
18 1 10 0 9 15 13 12 9 14 13 10 10 9 7 9 15 13 2
13 10 9 7 10 9 9 4 13 1 15 0 9 2
23 15 4 13 1 15 0 9 7 4 4 13 2 10 9 2 13 9 2 7 10 12 9 2
25 9 1 10 9 13 14 13 0 2 7 15 4 3 13 10 9 1 16 3 9 4 13 10 9 2
16 10 9 2 9 9 2 13 0 2 13 9 1 1 10 9 2
37 3 15 13 10 0 9 1 10 3 0 9 1 10 9 1 15 9 3 3 1 9 2 15 13 14 13 10 9 9 10 10 9 14 13 15 1 2
34 10 9 13 0 2 3 10 0 9 0 9 2 7 13 14 13 14 13 2 7 3 0 0 9 13 14 13 15 13 14 13 3 3 2
8 13 0 16 15 15 9 9 13
16 15 13 10 9 13 3 3 0 3 13 1 10 9 1 3 2
6 15 9 13 0 3 2
26 15 10 13 14 13 1 10 9 9 10 13 10 0 12 9 0 15 4 3 3 4 13 1 12 9 2
26 15 13 3 0 1 10 9 7 3 3 4 4 13 15 2 7 10 9 9 15 13 1 13 10 9 2
42 3 2 15 13 15 15 4 14 13 15 16 15 13 10 9 9 2 7 15 13 3 3 0 1 10 9 16 15 13 14 13 13 1 10 9 7 13 15 16 13 3 2
32 15 4 14 13 16 10 9 13 10 0 9 7 15 2 7 15 13 14 13 7 13 1 9 1 12 9 16 15 13 10 9 2
18 1 15 2 15 3 13 14 13 15 9 1 9 7 9 13 10 9 2
25 15 13 0 7 13 15 9 10 15 3 13 10 9 1 7 15 13 1 0 9 7 10 0 9 2
21 1 9 15 13 15 13 11 7 15 13 1 9 15 13 11 2 10 13 14 0 2
49 15 13 2 15 4 14 13 16 15 4 14 13 2 7 16 15 13 14 13 7 13 15 9 1 15 9 2 15 13 10 9 15 4 13 14 13 15 3 9 13 1 10 9 1 10 9 7 9 2
7 10 0 0 15 4 3 13
13 15 13 1 3 10 0 0 9 15 4 3 13 2
4 10 9 13 2
23 15 13 1 15 9 7 16 13 14 13 15 1 2 15 13 15 9 13 1 9 0 14 2
14 15 13 3 12 0 9 16 15 13 14 13 15 3 2
23 15 3 13 15 9 14 9 13 1 7 13 14 13 15 5 12 0 16 15 15 4 13 2
15 15 13 1 10 9 9 7 15 13 15 12 9 9 3 2
16 15 4 13 1 10 9 1 12 9 14 3 13 1 10 9 2
18 3 14 13 16 10 9 9 13 3 3 0 16 13 1 10 0 9 2
16 15 13 0 7 0 2 3 15 13 10 9 15 13 9 1 2
18 15 13 14 13 1 3 12 9 1 15 9 16 10 9 13 3 0 2
33 15 4 14 13 3 15 13 0 14 13 9 9 2 9 9 7 9 9 9 3 3 1 9 9 13 3 0 7 11 11 13 15 2
19 10 0 9 10 13 0 13 10 13 9 7 10 9 9 9 13 3 0 2
7 15 4 3 13 3 3 2
17 11 11 1 11 13 10 12 9 0 1 9 7 9 1 10 9 2
25 15 13 10 9 3 11 11 13 9 12 0 9 1 11 2 15 13 14 13 10 9 1 10 9 2
2 0 9
15 12 1 10 0 9 15 4 3 13 1 10 9 9 9 2
13 15 13 15 9 3 1 10 9 1 10 9 9 2
10 3 12 9 3 2 10 9 13 1 2
23 15 13 15 3 3 14 13 15 13 3 2 7 0 1 10 9 3 10 0 9 13 1 2
31 15 13 3 1 10 0 9 7 15 13 15 3 2 7 10 9 3 15 13 1 10 9 2 10 9 7 9 4 14 13 2
23 3 1 10 0 9 1 12 9 7 10 0 9 1 12 9 2 15 13 10 9 3 3 2
49 3 15 13 15 9 1 10 9 2 15 13 0 2 10 9 2 2 4 15 13 15 4 13 10 9 2 4 15 13 15 4 13 10 9 1 15 0 9 2 4 15 3 13 2 15 13 0 2 2
7 6 2 9 1 10 0 2
13 15 13 3 7 13 15 3 15 13 14 1 9 2
28 15 13 10 9 1 10 9 9 2 7 4 15 13 3 15 13 13 14 13 10 12 9 1 9 1 10 9 2
13 7 15 4 15 13 2 16 15 9 13 10 9 2
22 1 10 9 1 10 9 4 10 9 2 2 15 13 0 2 3 13 1 1 15 9 2
18 15 2 7 9 0 1 15 9 2 4 3 13 1 11 11 11 3 2
16 6 2 16 3 3 10 0 9 15 13 1 10 9 13 1 2
6 4 14 13 10 9 2
21 15 13 1 10 9 9 9 10 15 13 13 1 16 16 15 4 13 14 4 13 2
12 15 13 16 15 4 13 10 9 15 13 1 2
15 15 13 15 4 4 13 3 1 10 12 15 13 14 13 2
13 15 13 15 1 3 15 13 0 7 4 13 12 2
20 3 15 13 1 10 9 7 13 14 13 10 0 9 1 0 15 4 14 13 2
21 15 13 10 0 9 1 9 7 13 15 14 13 13 16 15 13 14 13 10 9 2
19 15 13 10 9 7 10 9 10 4 14 13 7 13 11 1 15 9 3 2
14 10 9 1 10 9 13 3 0 15 4 14 13 15 2
29 15 13 15 15 4 14 13 10 9 15 4 13 7 10 9 4 3 13 15 1 10 9 3 15 4 14 13 15 2
11 15 13 15 4 14 13 15 15 13 1 2
22 15 13 15 14 13 10 0 9 3 7 15 13 15 15 13 14 13 15 1 10 9 2
24 15 13 15 15 13 3 0 15 4 13 9 14 13 15 16 15 4 14 13 7 13 10 9 2
18 15 13 15 4 13 14 13 15 3 7 4 15 3 3 13 10 9 2
22 1 10 9 1 15 9 15 13 15 10 9 4 4 13 7 10 13 10 9 15 13 2
6 4 14 13 10 9 2
19 15 13 3 0 9 10 13 15 9 14 13 14 13 1 1 10 0 9 2
21 15 4 3 13 10 9 1 9 7 3 15 4 13 3 1 10 9 14 0 9 2
31 3 15 3 13 1 11 15 3 13 3 16 15 4 13 15 4 13 0 14 13 10 12 9 9 16 15 13 14 13 3 2
15 15 13 1 1 12 1 10 9 15 13 3 0 7 0 2
17 3 13 1 3 13 0 2 10 9 13 0 7 10 9 13 0 2
15 10 9 9 4 3 13 2 15 4 3 13 7 13 3 2
9 15 13 14 13 10 9 9 3 2
32 3 1 15 0 9 2 15 4 13 1 0 9 7 13 3 14 13 15 9 16 15 4 13 15 4 4 16 15 4 13 3 2
38 10 9 13 3 0 2 13 15 16 3 13 15 9 2 7 3 13 15 14 13 1 3 15 4 13 14 13 9 14 3 13 10 9 16 13 15 9 2
47 15 13 0 14 13 15 7 3 16 13 10 5 12 9 2 10 10 9 9 15 13 15 1 13 15 4 14 13 14 13 16 15 13 9 1 9 2 7 4 13 1 1 10 3 0 9 2
21 15 4 13 16 15 4 4 13 10 9 1 10 9 9 7 10 9 14 0 9 2
4 0 1 9 2
4 15 13 0 2
10 15 4 3 13 10 9 1 10 9 2
17 10 9 7 9 13 14 0 0 14 13 1 10 9 1 10 9 2
11 15 13 0 9 1 10 9 2 11 11 2
5 10 9 9 1 11
8 15 13 0 14 13 10 9 2
13 3 1 1 9 15 13 10 9 7 13 15 9 2
15 3 13 2 3 13 2 14 0 2 7 13 0 9 3 2
33 15 3 13 10 9 9 1 10 9 7 15 13 15 9 9 3 14 13 10 9 16 16 15 4 14 13 1 2 15 4 13 15 2
11 15 13 10 0 9 9 1 11 13 11 2
21 16 15 3 13 9 1 15 9 15 13 2 15 4 13 15 2 15 13 0 2 2
23 15 4 15 13 14 13 2 13 15 4 14 13 15 7 13 3 1 9 3 1 15 9 2
24 15 13 14 13 3 0 7 3 15 13 15 9 9 1 15 0 9 10 13 10 0 9 9 2
22 10 0 9 1 15 13 13 15 13 15 13 3 0 2 15 4 13 14 13 15 9 2
14 5 12 3 15 9 13 3 10 9 13 15 10 9 2
24 11 13 10 0 9 2 13 10 0 9 10 0 9 2 7 15 13 10 9 1 1 10 9 2
7 15 13 10 0 9 3 2
15 15 3 2 13 2 15 1 0 7 15 3 13 1 9 2
6 15 4 3 13 3 2
9 15 13 10 9 9 1 3 11 2
21 15 3 13 15 16 15 13 1 10 9 1 11 7 11 7 16 15 13 3 9 2
9 15 13 15 0 9 1 10 9 2
15 15 13 3 0 1 10 9 16 15 13 10 0 9 3 2
14 3 15 4 14 13 10 0 9 7 15 13 15 3 2
3 0 9 2
3 13 3 2
3 3 0 2
22 13 1 11 11 13 15 0 9 13 1 10 9 2 3 15 4 14 13 15 14 13 2
11 15 13 2 15 13 14 4 13 3 3 2
20 3 2 3 15 13 14 13 15 9 14 13 10 9 15 4 3 13 0 1 2
30 15 13 14 13 1 10 9 2 7 13 15 9 3 15 13 10 9 1 0 16 15 15 13 14 13 10 0 9 13 2
49 13 3 2 11 3 13 15 16 15 13 14 13 3 14 13 10 9 2 15 13 10 9 14 13 16 15 4 13 10 9 2 9 1 1 10 0 2 15 4 13 2 7 15 13 9 14 13 1 2
7 6 2 15 13 9 12 2
19 15 4 14 13 14 13 15 3 2 7 15 4 13 14 13 15 1 15 2
39 3 2 3 16 15 4 13 14 13 16 15 4 13 14 13 10 11 5 12 5 16 13 3 15 11 13 15 14 13 2 15 13 15 13 14 13 15 9 2
33 0 9 2 16 10 4 13 7 13 2 15 13 11 16 15 9 9 4 13 15 1 10 5 0 9 9 1 10 9 1 10 9 2
4 15 13 6 2
48 6 2 3 2 15 4 3 13 1 10 9 9 1 5 12 5 2 10 0 1 11 12 2 12 7 10 10 11 13 14 13 1 10 9 13 2 6 2 15 4 14 13 14 13 10 9 2 2
25 15 4 14 13 14 13 10 9 2 3 2 7 15 13 14 15 15 13 1 9 3 13 10 9 2
13 1 10 9 1 15 0 9 2 15 13 15 1 2
6 9 0 2 0 9 9
13 15 13 3 9 1 10 9 15 13 1 10 9 2
2 3 2
12 16 15 13 15 0 9 16 15 13 1 9 2
4 0 2 0 2
16 6 15 13 3 7 13 3 10 1 15 9 1 10 0 9 2
11 2 15 3 13 15 10 9 3 3 2 2
27 10 9 15 4 13 15 10 9 7 13 15 10 9 3 2 11 2 13 0 7 3 0 2 1 10 9 2
19 3 12 9 2 11 13 10 9 2 3 14 13 1 9 2 16 13 15 2
30 15 3 13 14 13 10 0 9 13 1 10 9 1 10 9 9 9 10 15 4 13 7 10 4 13 14 4 13 3 2
18 10 0 9 13 1 10 9 4 14 13 16 15 3 13 10 9 13 2
19 15 4 13 1 9 2 7 15 13 15 13 10 9 2 9 1 15 9 2
32 15 13 3 1 10 9 11 4 13 1 15 9 2 7 10 9 13 3 14 13 15 7 13 16 15 4 13 9 1 10 9 2
3 15 13 2
3 7 13 2
6 15 3 3 13 15 2
18 15 4 13 14 13 10 0 9 0 9 14 13 3 15 9 4 13 2
15 15 13 13 0 9 2 9 9 7 4 14 13 3 0 2
24 15 4 13 12 9 7 15 3 4 14 13 15 9 2 10 13 14 0 2 15 4 13 2 2
44 9 13 2 15 4 13 0 14 13 10 0 9 1 10 9 9 2 10 15 13 2 7 15 13 14 3 0 7 11 13 9 13 3 2 15 4 13 14 13 14 13 15 13 2
2 0 9
5 13 4 14 13 2
14 15 9 1 11 11 11 4 13 12 1 9 7 9 2
13 16 15 4 13 15 10 0 9 1 9 15 4 2
20 1 11 9 2 12 15 13 9 1 11 11 11 7 13 16 11 14 13 15 2
15 1 12 9 10 9 9 13 1 1 15 9 1 12 9 2
20 15 4 3 13 15 4 4 13 1 10 9 7 10 9 9 15 4 4 13 2
8 10 12 4 13 15 10 9 2
20 15 13 5 12 1 10 9 9 2 10 13 0 7 0 9 1 10 9 9 2
60 1 9 15 13 0 10 0 9 4 13 2 10 9 1 9 13 0 1 10 9 2 10 9 1 9 4 13 10 12 9 0 14 13 10 9 2 10 9 0 9 4 13 1 13 10 9 14 13 1 10 9 2 7 10 9 4 13 10 9 2
7 3 4 15 13 10 9 2
64 16 13 1 11 9 1 11 11 11 2 11 2 10 11 11 11 7 11 11 11 10 0 3 13 15 3 7 13 15 4 13 3 14 13 10 9 7 9 1 9 1 10 0 9 7 1 10 0 9 15 4 4 3 13 7 1 10 0 9 15 4 4 13 2
19 10 9 9 1 11 11 11 13 0 13 3 15 9 14 3 13 1 9 2
10 3 15 13 1 9 13 10 9 9 2
24 15 13 10 9 7 9 1 10 9 13 13 9 9 1 15 9 7 0 13 1 9 14 9 2
16 3 3 15 4 13 14 13 0 9 9 7 0 13 1 9 2
3 0 9 9
27 15 4 13 1 10 9 9 12 9 3 7 1 3 15 4 13 10 0 9 7 4 14 13 1 10 9 2
12 3 2 10 9 9 13 15 14 13 10 9 2
22 10 3 0 9 1 15 3 13 10 11 11 11 7 15 4 13 14 3 13 1 11 2
32 15 3 13 15 7 13 15 1 10 2 0 9 7 3 10 0 9 15 13 2 3 0 2 0 7 3 0 16 13 9 2 2
18 15 13 10 9 3 3 12 9 16 15 3 13 1 10 12 9 9 2
36 15 13 14 13 15 0 9 12 9 7 1 10 0 9 10 9 13 0 3 14 13 15 9 1 15 9 7 3 13 15 16 13 15 0 9 2
29 12 9 1 15 0 9 2 15 13 10 9 1 11 13 15 1 15 9 7 14 13 3 3 3 16 15 13 0 2
20 15 9 13 16 15 13 3 7 13 3 3 16 13 11 1 10 11 2 11 2
18 15 13 16 13 10 9 3 3 16 15 4 14 13 0 13 10 9 2
17 11 3 13 2 16 15 13 3 3 3 4 14 15 13 15 9 2
23 15 13 15 7 13 16 15 4 13 0 14 13 15 7 10 15 13 14 13 13 14 13 2
11 13 15 7 3 3 13 7 13 1 15 2
12 4 14 13 2 15 4 13 9 1 15 2 2
6 2 10 9 13 9 2
10 3 15 13 3 13 3 1 15 0 2
16 11 2 15 4 14 13 15 3 16 13 15 13 1 15 9 2
37 1 15 9 2 13 15 1 15 9 2 15 13 0 1 15 9 16 13 11 13 10 2 0 9 2 3 0 10 0 9 7 0 9 9 15 13 2
7 9 1 9 1 11 11 11
26 15 9 7 15 13 1 11 11 10 9 3 7 4 13 3 10 1 10 0 9 16 15 13 0 9 2
13 6 15 13 15 10 9 14 13 12 10 15 13 2
13 7 15 4 14 3 13 9 1 11 15 13 15 2
39 9 15 4 13 3 4 13 3 0 7 3 13 1 10 0 0 9 1 10 11 11 9 15 4 13 1 2 7 13 15 15 4 13 1 10 9 1 15 2
26 15 3 13 14 13 1 10 0 9 12 9 3 15 13 14 13 10 11 11 11 11 1 1 11 11 2
15 15 13 3 7 13 10 9 9 7 4 14 13 13 3 2
12 15 13 10 0 11 11 11 15 4 3 13 2
10 15 3 13 15 9 9 7 9 9 2
9 7 10 9 15 4 13 13 0 2
9 9 4 3 13 3 7 13 0 2
13 15 9 13 3 0 1 10 9 1 9 15 13 2
11 10 9 13 3 3 3 0 14 13 1 2
12 15 13 3 0 16 13 15 9 3 1 15 2
14 15 4 14 13 14 13 7 13 3 3 1 0 9 2
33 3 9 13 1 10 0 9 3 1 0 7 3 3 9 4 13 3 7 13 15 16 15 13 15 12 9 2 15 4 14 13 15 2
8 7 15 4 13 3 1 0 2
4 11 11 2 11
45 9 15 4 13 1 3 16 9 13 10 9 16 2 10 1 10 0 9 4 13 1 8 9 7 9 2 7 15 4 13 15 16 15 4 14 13 10 9 1 16 13 1 15 9 2
12 15 13 1 11 7 3 13 3 10 9 3 2
7 3 10 9 13 3 0 2
8 16 15 13 15 13 10 0 2
11 7 15 4 14 13 15 1 16 13 3 2
10 11 11 1 11 11 13 14 10 0 9
41 15 13 14 0 1 10 9 1 10 0 9 3 2 7 15 4 13 1 0 9 16 11 11 11 11 13 14 10 9 1 15 9 2 7 13 3 3 0 7 0 2
17 15 4 13 14 13 7 13 15 0 0 9 1 1 0 0 9 2
11 15 13 10 9 9 1 11 12 2 12 2
37 3 15 13 3 15 13 15 11 11 11 2 3 16 15 13 14 13 1 10 9 1 12 9 13 9 2 16 15 4 3 13 15 4 13 1 2 2
16 15 3 13 16 1 12 9 15 2 13 3 3 12 9 2 2
12 12 9 7 3 3 12 9 13 3 0 9 2
23 15 4 14 3 13 15 10 9 14 13 15 4 13 1 10 9 3 2 10 15 4 13 2
14 10 11 11 11 4 14 13 1 9 7 4 4 13 2
9 15 3 3 3 13 15 13 0 2
13 3 13 15 13 0 7 13 1 1 10 9 9 2
28 3 2 3 2 3 15 13 15 13 0 2 3 16 15 13 14 12 5 0 2 2 7 15 4 13 15 13 2
23 15 13 3 0 0 7 4 14 13 14 13 2 7 9 1 10 9 15 13 10 0 9 2
30 15 2 1 1 15 9 2 13 10 9 14 13 10 9 1 15 9 16 15 4 14 3 13 14 13 15 9 16 13 2
32 3 15 11 15 13 1 10 0 9 13 2 15 4 13 0 14 4 13 1 10 9 9 1 15 15 4 13 9 1 15 2 2
5 15 13 15 3 2
64 16 15 13 10 9 15 4 13 1 15 7 13 15 4 13 7 3 13 15 9 2 7 14 13 15 15 4 13 1 3 15 13 9 1 0 9 7 13 15 13 15 15 13 2 3 15 4 14 13 1 15 2 13 1 10 9 2 15 13 10 9 1 15 2
12 15 15 4 13 1 10 0 2 0 9 2 2
16 15 4 13 3 13 11 11 13 1 10 2 0 9 2 9 2
25 15 4 3 13 3 0 14 13 15 12 9 3 2 13 16 15 4 14 3 13 10 9 13 3 2
23 15 4 13 10 9 7 4 13 1 3 0 10 9 13 2 7 10 10 9 1 10 9 2
22 15 13 0 16 11 13 16 15 2 0 2 9 4 14 13 10 0 9 14 13 15 2
39 7 15 4 13 9 1 9 9 15 2 10 9 2 15 4 14 13 3 2 2 7 9 4 13 0 9 7 9 16 15 15 13 3 15 9 13 0 9 2
34 9 15 13 10 9 13 1 10 9 3 2 7 15 13 0 14 13 15 13 0 7 0 14 13 6 16 15 13 15 4 13 10 9 2
35 15 13 2 13 1 15 0 9 2 16 15 13 10 9 1 9 2 3 15 4 4 13 9 3 2 7 4 13 10 9 0 1 0 9 2
46 15 13 15 13 10 9 2 7 16 15 13 10 0 9 2 3 15 13 0 9 16 15 9 4 3 13 1 9 14 13 2 7 15 13 0 1 15 14 13 1 10 9 14 13 15 2
11 7 14 1 10 9 1 0 9 14 9 2
49 15 4 3 13 10 9 1 11 11 2 14 13 15 2 10 4 4 13 15 9 10 9 14 13 7 13 1 11 11 10 9 9 2 13 0 1 10 9 7 3 13 10 9 14 13 1 9 3 2
27 10 9 4 13 14 13 9 3 1 0 9 2 3 13 14 15 0 14 13 15 4 13 15 15 4 13 2
28 15 9 13 3 1 0 2 7 12 1 15 15 13 4 13 10 0 0 1 9 3 15 2 3 3 3 2 2
40 13 10 0 3 0 1 15 9 1 10 9 1 15 2 7 3 4 14 13 1 0 9 13 16 15 4 14 13 14 13 3 2 3 16 15 13 15 0 9 2
3 0 9 3
29 15 13 11 9 2 15 13 3 2 15 4 13 1 9 3 16 13 10 9 7 3 9 13 2 4 15 13 15 2
26 3 15 13 2 15 13 1 10 11 11 9 1 11 11 2 13 1 12 2 4 15 13 1 10 11 2
13 15 13 6 2 11 1 11 11 2 13 11 11 2
23 15 13 7 13 2 6 2 10 11 13 1 11 11 2 7 15 13 1 10 11 2 11 2
11 7 15 13 2 15 13 1 11 1 11 2
39 7 15 13 2 6 2 11 11 11 2 7 15 13 2 6 2 11 13 10 9 2 16 15 13 1 10 11 1 11 15 13 3 0 2 13 11 1 11 2
16 15 13 2 6 2 15 13 1 10 11 11 11 1 11 11 2
21 15 13 2 15 14 13 10 9 2 15 13 14 13 1 9 2 15 13 1 11 2
6 13 11 1 15 9 2
16 15 13 13 2 15 13 1 11 7 11 2 4 15 13 3 2
11 15 13 2 15 13 14 13 10 0 9 2
8 6 2 12 11 11 15 13 2
13 15 13 2 3 15 13 15 15 13 1 11 11 2
54 15 13 10 9 1 10 9 2 15 13 2 15 13 14 13 15 9 2 15 13 2 4 15 13 1 11 7 11 2 15 13 2 15 0 9 2 15 13 12 2 12 2 12 2 12 11 2 13 15 0 2 15 13 2
16 6 15 13 0 2 6 2 15 13 2 13 15 1 9 9 2
5 6 2 15 13 2
19 11 2 1 3 1 11 7 11 6 2 15 13 2 12 9 3 1 15 2
5 15 13 1 11 2
7 15 13 3 3 1 11 2
11 15 13 2 13 15 11 1 1 1 11 2
8 6 2 15 13 3 1 11 2
22 11 2 15 13 2 13 11 11 7 15 13 12 9 3 1 11 7 12 3 1 11 2
19 6 2 15 13 2 3 3 4 15 13 3 2 15 4 14 13 1 11 2
21 6 2 1 0 9 7 9 15 13 1 2 13 10 9 2 7 13 1 11 14 2
12 0 14 13 9 7 14 0 14 13 10 9 2
14 11 13 3 3 3 14 13 15 15 9 3 1 11 2
26 15 13 3 0 2 0 14 13 10 9 7 0 14 13 16 15 14 13 1 9 14 13 13 15 9 2
25 15 9 4 13 3 1 11 7 15 13 15 9 7 13 13 2 9 4 13 1 10 9 2 2 2
20 1 10 9 15 13 12 1 10 9 1 15 9 13 3 10 9 4 13 3 2
19 15 13 15 9 15 13 15 15 4 13 10 9 7 13 15 13 9 1 2
4 15 13 9 2
37 15 3 13 10 9 7 10 9 15 13 1 13 15 4 13 9 3 14 13 1 15 7 4 14 13 3 2 12 9 13 7 13 7 15 13 9 2
37 15 3 13 3 7 4 13 16 9 2 7 9 2 4 13 1 10 9 2 6 1 15 9 2 10 9 13 1 1 10 9 10 13 9 1 9 2
17 15 3 13 3 3 16 14 13 2 15 4 13 1 12 9 2 2
20 6 2 3 15 13 1 5 12 1 9 15 13 15 14 13 1 7 13 0 2
2 6 2
7 15 4 13 1 12 9 2
72 15 13 3 0 1 10 9 2 15 4 13 10 1 12 9 16 15 14 13 3 7 13 10 12 9 10 4 13 2 10 9 13 0 3 14 13 10 9 1 15 7 15 13 3 3 2 7 15 4 14 13 14 13 10 9 14 13 16 15 3 13 10 0 9 7 4 3 13 10 0 9 2
42 3 15 13 16 15 4 14 13 14 13 10 9 14 13 10 9 10 15 13 3 15 4 13 10 9 14 13 9 15 4 13 16 3 15 13 9 16 15 13 15 9 2
3 13 3 2
7 15 13 15 15 13 1 2
15 15 13 3 1 10 9 1 0 9 7 3 15 13 3 2
40 3 10 9 4 3 13 15 4 4 13 15 12 9 2 3 1 15 0 9 9 2 9 7 9 14 13 10 9 15 4 13 1 10 12 2 9 1 15 9 2
14 9 1 9 2 9 9 2 0 9 9 13 0 15 2
21 15 13 10 2 12 2 9 7 13 1 10 0 9 9 12 9 16 15 13 1 2
18 15 3 13 10 12 9 2 10 4 13 2 7 13 1 0 9 9 2
14 15 13 10 9 1 10 5 12 9 2 10 15 13 2
19 10 9 4 13 14 13 1 10 0 9 2 7 15 13 15 1 10 0 2
25 10 9 9 2 10 15 13 1 10 9 2 13 1 0 9 2 13 16 15 13 9 2 3 9 2
18 1 0 9 2 15 4 14 13 1 9 2 7 15 13 9 14 13 2
14 3 1 15 9 10 9 3 2 10 9 13 0 2 2
4 3 10 9 2
32 3 10 9 13 15 9 1 10 9 1 10 9 1 10 9 7 13 15 3 16 15 4 14 4 13 1 12 9 2 10 9 2
5 3 15 13 0 2
23 15 13 1 12 9 2 13 10 9 3 2 7 10 9 1 10 9 1 9 1 15 9 2
31 9 1 10 9 2 9 8 2 16 15 13 10 9 1 10 9 1 15 9 15 4 13 15 16 13 10 9 1 10 9 2
24 16 15 13 15 4 13 10 9 1 15 9 3 1 15 2 15 4 13 15 5 12 1 9 2
11 15 13 10 9 1 10 9 14 13 0 2
20 9 8 2 16 15 13 10 9 9 3 2 15 4 13 15 5 12 1 9 2
42 9 2 16 15 13 10 0 9 2 2 1 12 9 2 15 13 15 5 12 1 10 0 9 2 5 12 1 10 0 9 2 7 1 12 9 15 13 10 0 9 9 2
11 9 8 2 9 13 12 9 1 12 9 2
6 3 3 7 3 3 2
11 16 15 13 3 2 15 4 3 13 1 2
9 2 1 15 2 15 4 14 13 2
6 15 3 13 9 3 2
10 10 10 9 4 13 1 10 9 2 2
20 9 2 0 9 2 9 9 2 7 0 9 9 1 10 9 10 4 14 13 2
17 15 13 10 9 9 1 0 9 7 13 1 10 9 1 0 9 2
4 10 9 9 2
20 9 13 0 2 7 13 10 0 2 0 2 9 2 9 9 10 4 14 13 2
11 9 13 0 1 9 9 10 13 9 9 2
3 10 9 2
15 10 9 13 10 9 1 0 9 9 2 7 3 12 13 2
10 4 14 13 10 9 1 10 12 9 2
11 15 13 3 1 10 9 3 15 13 9 2
3 0 9 2
26 15 4 13 3 16 15 4 13 10 0 9 9 3 1 5 12 2 7 15 4 14 13 15 9 9 2
5 13 1 10 9 2
39 10 0 9 10 4 13 1 10 9 1 11 13 14 13 3 0 9 13 0 9 13 9 16 2 9 2 4 13 14 2 13 2 10 9 2 9 7 9 2
24 10 9 13 2 1 15 7 15 9 9 14 9 2 15 13 10 0 0 9 1 10 0 9 2
11 15 13 10 3 3 7 3 9 2 3 2
17 3 2 10 0 1 10 0 9 13 1 10 0 9 1 10 9 2
34 10 9 9 13 10 0 9 15 4 3 13 13 1 9 1 15 2 15 4 3 3 13 15 13 9 16 15 4 14 13 1 15 2 2
21 16 15 13 3 0 2 15 3 4 14 13 0 9 14 13 16 15 3 13 15 2
14 15 4 13 2 10 9 7 9 13 1 1 10 9 2
47 3 3 2 1 10 12 1 15 15 13 3 2 12 9 1 9 13 15 13 1 0 2 7 13 10 9 1 15 9 2 7 6 2 10 12 9 1 9 4 13 10 12 2 9 9 2 2
11 9 13 3 10 0 2 7 2 0 9 2
24 10 0 9 7 0 9 13 3 3 0 2 0 2 16 10 9 13 3 0 7 5 7 0 2
26 10 9 13 10 12 5 9 1 0 9 1 10 9 1 10 0 2 0 9 15 3 13 1 0 9 2
16 9 13 2 6 2 15 13 0 2 15 4 14 3 13 9 2
8 15 13 15 13 15 10 9 2
11 6 2 6 2 10 9 9 13 3 0 2
23 10 0 9 9 13 3 0 2 7 13 1 9 9 2 3 0 1 10 9 1 10 9 2
14 7 15 2 6 2 15 3 4 14 13 15 15 13 2
35 9 13 0 2 7 9 0 2 7 9 10 4 13 14 13 0 4 13 10 0 9 16 13 15 9 14 13 0 7 0 2 3 3 0 2
41 3 4 15 14 13 1 10 9 13 11 4 13 14 13 0 16 15 9 13 2 7 16 10 0 0 9 13 14 13 2 2 15 4 4 13 10 0 0 0 9 2
38 7 15 4 14 13 3 13 9 0 2 16 3 15 4 3 13 0 2 0 9 3 2 7 0 9 2 0 9 2 0 9 13 7 3 0 9 9 2
21 9 2 3 15 13 1 10 9 2 15 4 13 16 12 7 12 13 15 0 9 2
23 3 15 13 1 12 2 7 13 1 12 2 15 13 10 0 12 7 12 0 9 13 15 2
26 4 15 13 15 4 13 14 13 0 14 13 10 9 3 3 2 7 3 13 3 0 1 15 9 9 2
12 4 13 2 4 14 13 15 9 1 10 9 2
18 1 15 9 10 9 13 15 13 0 14 3 13 1 10 1 10 9 2
33 15 13 16 15 4 13 14 13 3 1 15 7 15 13 3 0 14 13 15 15 4 3 13 1 13 15 14 13 10 1 10 9 2
31 15 13 15 4 13 10 0 9 14 13 3 10 0 10 15 13 4 13 1 1 10 9 2 16 13 10 9 1 3 2 2
23 3 2 16 15 4 13 15 13 1 10 9 2 9 9 7 9 9 13 1 15 0 9 2
16 15 13 15 13 2 0 14 13 15 16 15 13 15 9 2 2
39 6 2 10 9 4 14 13 10 9 2 16 15 13 10 9 15 9 2 16 10 9 13 0 2 3 2 2 7 13 10 9 1 10 9 9 7 9 9 2
7 4 0 9 13 1 15 2
51 15 7 2 8 2 4 14 13 14 13 15 1 15 16 15 4 14 13 15 13 10 9 3 7 8 2 4 13 10 9 15 2 8 13 0 9 14 9 9 7 2 13 10 9 2 1 15 0 9 2 2
10 15 13 10 9 7 2 6 2 3 2
24 10 9 1 9 15 4 13 2 15 13 14 0 7 16 15 13 0 2 15 4 14 13 3 2
6 15 10 9 1 9 2
41 3 1 10 0 2 9 2 2 12 1 10 9 9 13 3 0 13 15 3 0 15 13 16 3 10 9 10 15 13 13 1 12 1 15 9 10 15 4 13 1 2
64 3 2 16 15 3 4 14 13 10 9 1 9 2 9 2 16 15 13 15 10 9 7 9 9 1 10 9 15 4 13 2 15 13 2 3 10 9 2 15 4 13 1 7 13 1 15 9 2 15 13 16 10 9 4 13 3 3 1 10 9 15 13 3 2
19 15 9 2 3 16 15 13 0 2 4 14 13 3 7 13 1 10 9 2
7 13 9 1 2 2 6 2
12 15 4 14 13 3 7 15 4 13 0 2 2
39 16 15 13 14 13 10 2 13 10 9 3 0 15 13 7 13 7 13 15 1 10 9 15 4 3 14 13 2 9 10 4 3 13 15 2 6 2 3 2
8 3 2 4 14 13 15 9 2
13 0 9 1 10 9 13 3 0 7 3 0 9 2
20 14 9 10 13 16 15 13 9 14 13 7 13 9 1 0 9 7 9 9 2
42 15 13 3 3 16 11 11 4 13 0 7 15 4 14 13 15 14 13 15 1 1 10 9 3 3 13 15 1 10 9 15 4 13 1 10 3 0 9 1 15 9 2
3 0 9 2
22 16 3 13 11 11 1 10 9 2 15 13 0 1 10 0 9 13 1 15 11 9 2
14 15 13 15 9 3 1 10 11 14 13 10 13 9 2
80 15 13 3 12 9 1 10 9 9 16 9 13 0 14 13 15 7 4 3 13 14 13 15 9 1 10 9 2 15 13 3 15 15 4 13 14 13 2 7 10 0 9 13 15 10 9 4 1 10 9 13 1 10 9 2 3 15 4 14 13 15 13 3 2 7 15 3 13 10 9 9 2 9 10 10 0 11 13 2 2
24 16 3 2 15 13 14 13 3 1 3 3 12 0 9 16 2 3 2 10 0 13 1 15 2
23 16 15 13 14 13 1 15 9 2 15 4 13 15 13 10 10 9 0 9 13 3 13 2
30 15 4 13 14 13 10 9 1 10 9 9 7 9 9 16 15 4 4 13 1 10 9 7 4 13 15 13 14 0 2
21 16 15 3 13 3 1 15 9 2 15 13 0 7 13 9 3 1 10 9 9 2
8 6 2 12 0 9 2 6 2
23 10 13 11 2 15 13 1 15 9 14 13 3 7 13 10 0 12 9 2 10 13 0 2
23 15 4 14 4 13 3 2 7 15 4 14 13 10 0 9 15 4 13 1 9 3 3 2
14 3 3 2 15 13 1 10 10 9 16 4 13 1 2
23 15 13 10 9 13 2 7 3 13 10 9 16 15 13 3 3 5 12 0 16 15 13 2
31 15 13 15 13 10 0 9 2 7 13 15 2 16 13 7 10 0 9 1 15 9 7 15 9 9 1 3 1 10 9 2
33 3 2 3 15 13 1 10 9 9 2 15 4 13 16 15 13 14 10 0 9 2 7 13 14 3 10 0 9 1 15 9 9 2
24 3 15 13 15 1 1 15 2 1 10 9 15 13 15 3 13 12 1 10 0 9 1 9 2
4 6 2 6 2
10 3 15 13 3 15 0 0 9 13 2
17 15 13 15 4 4 13 1 10 9 2 3 15 13 1 10 9 2
18 1 12 9 3 2 7 12 9 16 15 13 2 15 9 4 3 13 2
31 10 0 9 16 15 13 2 15 4 13 7 13 16 2 15 2 13 15 9 9 2 10 15 4 4 13 1 10 9 2 2
25 3 3 2 15 4 4 13 1 12 9 2 3 15 4 13 14 13 1 7 13 15 10 0 9 2
26 3 3 15 4 14 13 15 3 1 9 2 7 15 3 4 14 13 12 0 9 14 13 1 15 2 2
19 10 0 9 2 10 9 4 13 15 9 9 7 10 0 9 13 14 3 2
53 3 3 2 15 4 14 13 15 3 14 13 1 15 16 3 15 4 14 13 15 9 14 9 9 2 6 2 2 3 15 4 13 14 13 1 11 2 13 1 12 9 3 1 10 9 9 4 15 13 10 9 2 2
22 1 11 15 13 7 3 15 13 10 0 9 2 9 14 13 9 15 13 9 1 15 2
23 3 15 4 4 13 15 1 15 10 9 2 7 15 13 0 15 4 3 13 10 0 9 2
24 10 9 1 10 11 13 3 0 7 15 4 14 13 14 13 10 9 1 9 10 15 4 13 2
26 15 4 3 13 3 3 2 7 3 13 10 0 9 1 10 9 1 9 15 3 13 1 15 9 2 2
