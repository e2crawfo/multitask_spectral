129 17
34 9 9 13 3 3 10 9 0 9 11 11 2 15 10 11 11 13 10 11 11 2 16 11 10 9 9 13 2 3 13 14 0 9 2
17 10 0 9 9 9 1 0 12 12 9 13 10 9 10 9 9 2
25 0 0 9 15 13 2 16 10 9 10 0 0 0 9 13 2 7 3 10 0 9 0 9 13 2
44 10 0 9 3 13 3 10 9 2 16 10 11 11 11 0 9 0 9 3 13 2 16 10 0 12 9 1 3 12 9 13 14 10 0 9 0 2 0 2 9 9 2 9 2
13 10 9 1 10 0 9 12 3 0 9 13 9 2
30 10 9 9 0 9 7 10 11 13 2 15 13 10 0 9 11 0 9 1 0 9 9 7 10 0 9 9 7 9 2
16 11 3 3 12 9 9 13 3 9 2 3 7 0 13 9 2
16 10 0 9 12 9 1 13 10 9 2 7 11 0 9 13 2
11 10 0 12 0 9 7 10 9 9 13 2
48 10 11 11 11 11 2 11 2 9 12 9 13 3 9 9 2 15 13 15 2 16 10 11 10 3 0 9 1 0 9 13 2 16 9 10 9 0 9 13 10 0 0 10 11 11 9 9 2
14 10 9 13 2 16 10 9 10 9 10 9 9 13 2
14 10 15 0 9 3 10 12 9 2 15 10 9 13 2
23 9 3 13 2 11 11 0 9 3 3 13 15 10 11 9 2 7 11 11 3 13 3 2
7 10 9 3 13 13 11 2
30 9 13 10 9 13 2 7 15 13 2 9 3 13 2 7 15 3 13 13 15 2 16 13 3 10 15 0 9 9 2
9 10 11 9 12 9 13 3 9 2
15 10 9 0 13 10 9 9 2 7 0 9 13 10 9 2
6 15 3 13 10 9 2
19 10 0 9 15 13 10 11 2 16 15 13 10 9 7 0 9 0 9 2
10 10 11 0 9 9 0 9 13 3 2
13 10 9 9 3 13 2 7 15 9 13 10 9 2
20 10 0 9 2 11 11 9 2 9 9 1 3 13 9 10 9 0 0 9 2
26 10 0 9 11 10 10 0 12 9 0 9 13 2 15 11 11 9 9 0 9 9 10 11 13 3 2
46 11 11 2 10 9 0 9 9 9 13 2 11 0 9 9 3 13 2 3 13 14 2 16 13 3 10 0 9 9 2 10 0 12 9 9 9 2 10 9 0 9 7 10 9 9 2
32 10 11 11 10 9 3 13 0 9 3 2 16 10 11 1 10 10 9 10 0 0 9 13 13 2 15 7 3 3 13 14 2
14 9 11 13 2 10 9 1 7 0 13 10 9 9 2
24 10 11 9 3 13 2 16 10 9 1 0 9 7 13 9 2 3 0 7 13 10 12 9 2
28 11 1 7 10 9 1 10 9 13 10 3 0 9 2 9 2 7 3 3 10 0 0 0 9 13 10 9 2
27 9 11 15 7 13 2 3 13 9 10 9 9 7 9 2 16 3 13 10 0 13 10 11 0 9 9 2
12 9 1 7 10 9 0 9 13 10 0 9 2
18 0 2 16 0 9 1 0 9 7 13 15 2 13 0 0 9 9 2
24 11 10 9 2 9 2 9 1 3 0 2 0 9 7 10 9 12 9 9 13 10 0 9 2
27 3 15 10 9 13 0 10 9 10 9 2 3 3 10 9 7 13 10 2 9 2 2 7 13 10 9 2
33 10 9 9 3 0 2 7 0 9 3 13 3 7 13 10 9 2 15 2 3 2 3 2 2 10 9 7 13 2 3 13 9 2
13 10 9 0 9 13 10 9 10 9 0 9 9 2
15 10 9 10 9 9 13 3 9 2 13 9 0 9 13 2
14 0 7 0 9 13 2 16 2 15 2 0 13 15 2
25 7 10 0 9 2 7 10 11 11 0 10 9 3 0 9 1 2 16 13 0 9 10 9 9 2
19 15 3 0 2 16 10 9 0 0 9 3 13 2 9 3 13 14 15 2
29 10 9 9 0 9 2 16 9 13 10 2 9 2 2 16 13 15 2 7 15 3 10 10 9 7 10 9 13 2
14 11 9 10 10 0 9 9 3 0 9 1 9 13 2
29 10 9 1 0 9 3 10 9 10 9 0 9 2 10 9 7 10 9 7 13 2 7 3 9 7 13 10 9 2
11 3 3 0 9 0 10 9 1 11 7 2
26 10 0 0 9 10 9 9 13 10 9 9 2 7 9 3 10 9 9 13 2 7 9 13 10 9 2
8 10 11 11 7 13 0 9 2
17 3 10 0 9 9 13 9 2 16 3 10 0 9 7 9 13 2
32 10 9 13 2 16 3 3 7 13 9 2 0 2 2 0 2 9 3 13 10 9 10 9 2 7 0 9 1 0 3 13 2
16 10 0 9 3 13 13 2 16 0 9 12 0 9 13 3 2
9 3 11 11 9 9 9 9 13 2
23 10 9 0 0 9 3 13 0 9 10 9 9 2 13 3 11 11 2 10 11 11 9 2
23 9 1 10 0 0 9 3 13 14 10 9 1 10 9 0 9 2 3 10 0 9 0 2
23 10 0 9 9 15 1 3 13 2 10 0 9 0 12 0 9 13 10 9 9 9 9 2
53 2 3 13 10 15 2 3 13 10 9 7 10 9 2 2 13 9 0 9 11 11 2 15 3 3 10 11 9 10 10 9 13 2 16 10 0 9 3 12 9 2 0 9 9 13 3 10 9 9 10 11 11 2
33 10 0 0 9 0 9 11 11 11 11 0 9 13 3 2 15 7 11 11 11 0 9 13 3 2 12 15 10 9 13 10 9 2
57 2 3 13 15 13 10 11 0 9 9 2 10 9 9 13 2 16 3 13 3 13 2 2 13 11 11 0 0 9 2 10 11 0 9 9 9 10 10 9 3 2 16 3 13 3 15 13 10 0 9 2 3 13 3 3 3 2
23 3 0 2 11 10 11 0 9 2 11 11 1 10 1 10 11 9 13 10 0 9 9 2
37 10 9 0 10 11 0 9 16 3 13 9 10 0 9 9 2 16 10 0 9 13 3 9 1 2 7 10 0 9 9 9 3 13 11 9 9 2
20 11 13 2 2 10 10 9 3 15 13 13 2 3 15 13 10 9 10 9 2
32 7 3 13 2 16 10 9 3 13 0 9 0 9 7 0 0 9 2 16 9 13 10 0 9 2 3 10 9 13 13 2 2
42 11 1 15 10 9 15 2 16 10 2 11 0 9 2 10 0 9 13 13 15 7 9 2 9 9 2 7 10 3 0 11 11 0 0 0 9 2 9 7 13 2 2
18 11 0 9 13 2 16 3 10 11 11 2 7 11 11 0 9 13 2
43 13 10 11 9 2 11 11 10 11 11 0 9 2 15 0 13 10 10 9 2 7 13 10 10 0 9 2 15 10 9 10 9 13 15 2 16 13 10 0 9 0 9 2
27 11 13 2 16 10 11 11 1 2 15 7 10 9 13 9 9 2 3 3 12 0 7 0 0 9 13 2
33 11 11 2 10 11 0 9 9 13 2 10 9 13 2 16 10 11 0 9 3 3 3 13 11 11 9 9 10 0 9 9 13 2
26 15 9 3 13 13 10 9 9 2 16 10 9 9 1 10 0 9 10 9 0 0 9 14 13 13 2
18 11 13 2 16 3 7 13 9 13 2 3 10 0 9 13 10 9 2
43 10 11 0 9 10 11 0 9 0 9 2 9 1 2 13 2 16 10 9 0 11 11 9 13 3 9 11 11 0 9 11 11 2 10 11 9 0 9 2 15 9 13 2
24 11 11 2 10 9 0 9 9 3 13 2 10 0 9 9 3 13 13 10 9 9 0 9 2
21 16 15 3 13 14 2 10 11 13 10 3 9 0 11 11 2 16 3 13 9 2
12 3 15 3 13 2 10 9 3 13 13 9 2
8 0 9 7 13 11 9 1 2
20 11 11 2 10 11 11 11 9 2 13 2 2 16 10 9 0 13 10 9 2
20 3 13 15 1 2 16 15 3 2 11 9 0 2 9 13 12 0 0 9 2
18 9 13 9 10 11 11 11 7 2 0 13 10 9 9 3 0 9 2
15 9 10 9 0 9 7 9 0 9 13 2 0 10 9 2
46 3 9 0 0 0 9 13 11 2 15 10 11 11 0 0 9 10 9 0 9 10 9 7 10 0 9 1 10 2 0 9 2 7 0 13 2 15 15 2 10 9 13 10 9 2 2
23 10 9 9 10 2 10 0 9 0 0 9 13 2 15 10 0 9 10 1 0 9 13 2
24 11 11 1 10 0 9 10 0 11 11 1 0 0 9 15 10 0 9 2 16 13 10 9 2
31 10 9 0 0 9 3 13 2 10 9 13 13 2 16 11 11 9 9 0 2 7 10 9 9 9 11 11 9 9 13 2
26 11 9 1 10 9 9 3 15 13 13 2 16 10 9 10 9 13 10 9 3 9 0 9 9 9 2
26 10 11 9 3 3 13 0 9 2 15 11 11 9 0 9 13 2 3 9 13 3 10 0 9 9 2
58 9 15 13 2 16 10 11 9 2 11 11 9 0 2 9 0 0 9 13 2 15 1 2 16 10 0 11 3 13 10 9 9 0 9 2 10 2 9 10 0 9 2 0 9 9 2 10 9 0 2 0 9 2 11 11 15 13 2
19 10 9 7 13 11 11 2 15 11 9 1 0 9 13 10 9 10 11 2
17 10 0 9 1 15 15 1 13 2 16 10 9 0 9 0 13 2
34 9 10 10 0 9 2 15 10 9 0 2 7 3 3 0 7 3 3 0 2 9 2 13 3 2 11 0 9 0 9 13 0 9 2
23 10 0 9 1 16 10 9 9 10 9 9 13 2 10 0 9 13 10 9 13 9 9 2
14 10 9 9 13 2 16 10 0 9 9 0 9 13 2
26 10 15 0 2 3 10 12 9 0 9 10 9 13 2 16 10 11 0 9 15 10 9 3 13 13 2
28 10 9 15 13 2 16 10 0 9 2 11 11 9 1 10 10 9 3 10 0 9 2 11 11 9 13 3 2
27 11 11 0 9 10 11 0 9 2 3 13 2 16 10 9 0 9 10 15 9 13 3 10 11 0 9 2
22 10 11 0 9 9 13 2 16 13 9 15 1 2 7 10 9 9 9 3 3 13 2
43 10 11 0 0 9 1 3 13 14 10 9 9 0 9 0 2 0 9 10 3 0 9 9 2 3 3 13 2 16 10 0 0 9 9 10 0 9 1 15 7 3 13 2
20 11 11 0 9 2 10 11 11 0 9 9 9 13 2 10 9 0 9 0 2
18 10 9 9 9 13 10 9 9 10 9 2 13 7 13 10 0 9 2
15 13 16 9 2 7 15 3 2 15 13 10 9 0 9 2
6 15 0 9 7 13 2
19 10 0 0 9 9 1 10 0 0 9 9 3 3 13 3 10 9 9 2
10 10 3 0 9 10 9 9 9 13 2
13 10 9 1 10 9 9 10 0 0 9 13 3 2
15 10 9 1 9 9 2 16 13 3 10 0 0 0 9 2
40 0 16 2 16 10 9 9 1 0 0 9 2 7 3 0 9 1 3 13 10 2 7 10 9 3 15 13 2 3 0 3 7 2 16 13 10 0 0 9 2
38 10 11 9 1 10 11 11 13 10 9 9 10 11 11 11 0 9 2 11 11 10 9 1 2 16 10 9 3 0 9 2 7 3 13 4 9 13 2
24 10 9 3 13 14 10 9 9 2 16 10 9 3 12 0 9 13 10 9 1 0 12 1 2
27 11 11 15 0 9 10 9 9 2 10 10 12 0 9 9 9 7 10 3 9 0 9 9 7 9 13 2
17 10 11 3 13 10 9 10 11 11 0 9 0 9 0 0 9 2
27 10 11 7 0 9 13 9 15 9 2 16 10 9 0 9 13 3 10 9 10 9 15 0 0 9 9 2
8 10 0 9 0 9 13 14 2
52 3 0 2 10 11 9 3 13 9 2 16 10 11 11 11 11 11 9 13 3 2 3 10 11 11 3 13 3 10 9 2 15 7 2 16 10 9 9 3 13 13 10 0 9 2 3 10 9 9 13 3 2
23 0 10 12 9 9 13 0 9 10 11 11 0 0 9 3 3 2 12 9 10 11 11 2
24 10 10 0 9 7 0 0 9 9 9 0 2 9 10 0 9 0 9 10 9 1 13 13 2
9 10 9 9 11 11 11 9 13 2
24 10 9 9 13 3 11 11 2 10 9 9 2 15 13 10 3 0 0 0 2 0 9 9 2
25 10 9 3 13 2 15 0 3 13 13 10 9 9 1 2 16 2 9 1 0 2 15 0 2 2
35 11 11 2 10 11 11 9 13 2 10 1 11 11 0 9 10 11 1 0 9 2 7 11 11 2 10 9 9 10 9 0 9 1 13 2
18 10 11 0 0 0 9 2 3 13 0 2 2 16 3 13 10 9 2
21 3 10 10 9 3 2 13 10 9 1 2 2 0 9 13 3 9 10 9 1 2
28 10 9 9 9 13 3 10 9 10 0 0 0 9 2 15 3 10 9 13 10 9 9 2 13 9 11 11 2
45 10 0 9 0 9 3 13 10 0 9 9 2 10 9 1 7 10 10 16 12 12 9 3 0 9 13 14 10 9 2 7 10 0 9 2 9 2 9 0 9 13 13 0 9 2
15 3 10 9 9 9 0 9 3 12 13 0 2 16 3 2
28 10 11 11 9 3 13 2 3 13 10 0 9 0 12 9 2 10 9 0 9 0 9 9 12 9 13 3 2
10 15 7 13 10 9 1 0 9 9 2
16 15 15 13 2 16 10 0 9 0 9 3 13 14 10 9 2
10 15 7 0 9 2 7 9 13 3 2
24 2 10 0 9 10 0 9 10 9 13 10 3 0 0 9 2 2 13 3 10 0 9 9 2
28 11 11 13 2 10 9 9 15 13 2 16 10 9 0 9 12 0 9 13 14 2 7 15 13 10 9 7 2
35 10 9 12 9 1 0 12 0 9 2 7 10 9 7 10 0 9 0 7 0 9 7 3 13 0 10 0 9 13 2 13 10 11 9 2
22 10 9 9 1 12 9 0 2 0 9 13 13 2 15 0 0 7 0 9 13 13 2
15 10 9 9 0 10 0 9 1 13 2 13 3 11 11 2
24 10 11 1 10 9 15 2 16 10 0 9 9 10 0 9 0 12 9 13 10 0 9 1 2
