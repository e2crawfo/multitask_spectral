2002 17
7 1 10 11 13 10 9 2
19 11 11 1 11 13 12 9 14 13 13 9 1 0 9 1 10 11 9 2
29 11 13 11 11 11 1 10 12 2 9 9 1 0 9 1 10 11 11 1 10 11 1 11 2 13 11 11 11 2
1 2
30 11 3 13 11 11 11 11 1 10 12 2 9 9 1 0 9 1 10 11 1 11 11 1 11 2 13 11 11 11 2
18 10 9 1 9 2 9 4 4 13 1 10 9 2 12 2 13 9 2
31 15 4 4 13 9 3 7 10 11 13 10 10 9 2 16 15 13 7 15 13 10 0 9 1 11 2 7 15 13 14 2
16 9 14 9 13 16 11 4 13 15 9 7 15 9 1 9 2
18 0 9 13 9 2 3 15 13 15 4 13 10 9 1 0 0 9 2
9 8 8 8 8 8 8 8 8 2
21 1 10 0 9 1 11 2 9 13 10 9 9 1 10 9 9 2 13 0 9 2
24 10 11 13 3 10 9 1 0 9 1 11 1 10 0 9 2 7 10 9 10 9 13 0 2
20 1 11 2 9 1 9 13 3 1 11 9 3 15 3 13 10 0 0 9 2
29 2 15 13 16 10 11 9 13 10 0 9 1 9 1 15 9 2 16 3 10 9 13 10 0 2 0 9 2 2
12 10 11 9 13 1 10 0 9 2 13 12 2
36 15 13 0 1 15 16 10 9 1 0 11 9 1 10 0 9 4 4 13 3 2 7 3 3 1 9 10 13 0 1 11 9 1 0 11 2
30 11 4 3 13 10 9 9 2 10 9 14 13 10 9 14 9 1 10 2 0 9 1 2 9 15 4 14 13 15 2
27 3 2 15 13 3 10 9 16 10 9 14 13 1 2 7 10 9 9 13 3 0 1 10 9 14 9 2
42 15 13 1 11 11 2 3 3 2 3 3 15 13 10 9 15 13 9 13 2 4 14 13 0 2 2 15 13 10 9 15 0 9 4 13 2 4 14 13 0 2 2
55 15 13 14 3 3 0 10 9 16 15 4 13 2 11 11 4 3 13 10 0 2 9 2 16 10 9 14 9 2 13 9 9 2 10 13 9 12 9 10 9 14 13 9 9 1 15 0 2 13 10 0 2 0 9 2
12 13 10 0 9 2 15 13 10 9 2 3 2
19 15 9 9 1 10 9 1 11 14 9 1 11 2 11 4 13 1 11 2
2 9 2
30 2 11 14 0 9 13 0 0 14 13 1 11 7 14 13 10 12 2 9 9 2 3 16 10 9 1 9 13 0 2
37 10 13 0 9 1 10 13 11 11 1 10 9 13 2 1 1 0 9 1 0 9 0 1 11 2 14 13 10 9 9 2 10 11 4 3 13 2
16 11 14 9 13 10 9 1 0 9 10 4 14 3 4 13 2
16 11 14 9 1 0 11 9 4 3 13 9 9 1 10 9 2
35 16 10 11 7 10 0 9 4 14 13 10 9 14 13 10 9 9 2 9 1 0 0 11 4 13 1 10 13 1 11 11 1 15 9 2
36 3 16 0 0 9 13 0 0 14 13 11 2 11 3 2 10 13 0 2 0 9 13 1 10 0 9 9 1 11 2 11 1 0 0 9 2
21 13 10 9 4 13 10 3 0 9 10 11 11 4 13 1 15 9 1 9 2 2
31 11 13 16 10 0 9 1 0 0 9 1 11 13 11 14 9 1 11 11 11 2 10 0 9 1 11 2 10 9 3 2
30 10 9 1 0 9 1 11 2 12 9 3 1 11 2 2 13 10 9 7 13 0 9 1 10 9 9 1 11 2 2
17 11 2 11 11 2 11 13 16 11 4 13 11 1 10 0 9 2
15 11 9 3 13 1 9 1 10 9 10 13 12 11 0 2
9 1 11 2 15 13 10 0 9 2
35 0 0 9 11 11 2 11 13 10 9 13 2 0 2 7 16 2 10 11 4 13 3 12 9 1 10 11 2 15 1 9 7 9 2 2
34 10 0 11 11 13 10 9 13 2 2 15 13 10 9 1 10 9 1 10 0 9 7 10 9 1 10 9 9 1 10 9 2 2 2
25 10 9 4 3 13 10 0 9 1 10 9 7 4 14 13 9 1 10 9 2 2 10 9 13 2
33 11 13 16 2 0 1 10 11 2 15 13 10 0 9 1 11 2 13 15 9 1 15 1 10 0 9 2 1 10 0 9 2 2
33 1 10 3 0 9 2 10 12 11 4 13 1 9 1 11 2 13 10 9 1 9 9 1 10 9 1 11 7 12 9 1 11 2
55 3 1 10 0 9 1 11 14 9 2 0 9 4 13 16 10 9 4 13 0 1 10 10 3 0 9 16 2 3 1 10 3 0 9 9 7 10 3 0 9 2 10 9 4 13 3 0 16 9 14 13 10 0 9 2
5 15 4 13 3 2
5 15 4 13 1 2
10 3 2 9 13 16 11 4 3 13 2
8 15 13 13 15 2 15 13 2
36 15 15 13 13 16 11 4 13 9 0 1 15 15 4 3 13 2 10 0 9 9 1 10 0 9 2 9 9 2 0 1 10 9 1 9 2
32 9 13 15 10 0 2 0 9 1 9 2 10 0 7 0 9 2 13 9 2 7 10 9 1 9 1 10 13 2 1 9 2
35 10 9 13 16 9 13 1 10 0 9 13 1 10 3 0 15 4 13 2 13 10 9 2 1 2 0 2 9 1 0 2 9 9 9 2
4 10 0 9 2
16 15 13 0 14 13 9 13 1 3 15 9 13 1 15 9 2
34 16 10 9 13 1 10 3 2 13 9 13 2 0 11 9 4 14 13 14 13 11 2 7 11 13 14 3 3 0 1 11 7 11 2
38 16 15 13 14 13 9 16 15 4 13 15 0 9 2 0 9 2 11 13 13 10 0 9 1 15 9 9 1 10 0 13 2 15 2 0 9 9 2
22 13 3 10 0 9 1 9 13 14 13 16 10 0 9 13 10 9 1 10 11 11 2
20 3 11 13 14 13 10 9 7 4 13 9 14 13 15 0 16 13 10 11 2
22 3 2 10 9 13 10 9 1 11 13 0 16 15 15 4 13 1 10 0 0 9 2
5 11 2 11 2 2
28 10 0 9 1 9 1 10 11 13 1 11 1 9 1 10 9 1 0 9 0 11 1 9 1 10 11 11 2
36 2 15 13 10 9 14 13 10 9 1 9 11 13 1 2 2 11 11 2 9 1 10 9 14 2 11 11 2 11 7 10 9 9 2 13 2
33 2 15 4 3 13 9 15 13 1 15 9 2 7 16 15 13 9 1 10 11 15 4 7 13 7 13 1 9 2 2 15 13 2
29 2 16 15 4 14 13 10 9 16 11 4 13 1 10 2 11 11 2 11 2 3 4 10 11 13 1 15 2 2
19 11 13 10 13 9 1 10 9 2 0 9 1 11 14 11 11 11 11 2
24 15 13 16 3 12 9 4 13 1 9 1 0 1 12 9 7 16 0 1 12 13 1 9 2
28 15 13 10 0 12 9 4 4 13 1 11 12 2 16 10 9 4 13 9 1 12 2 12 7 12 9 3 2
17 10 0 0 9 4 3 13 14 13 3 3 0 10 9 11 13 2
14 3 15 13 10 9 1 15 9 2 9 13 14 13 2
19 3 15 0 9 4 13 15 3 13 15 4 13 1 10 9 1 10 9 2
19 11 11 13 1 0 1 11 1 11 2 16 15 4 3 13 9 1 9 2
26 10 11 9 4 13 0 9 1 0 9 2 13 11 11 11 11 2 11 1 10 13 11 1 11 11 2
25 0 9 13 1 1 0 0 0 9 1 11 2 13 10 12 9 0 1 11 2 11 2 7 11 2
23 9 1 9 13 9 1 10 11 9 1 11 7 11 2 3 3 2 13 1 11 2 11 2
13 10 9 7 9 4 13 1 10 11 9 1 11 2
20 9 13 14 13 11 11 11 11 7 11 1 11 11 11 1 9 1 10 9 2
31 11 14 0 9 7 10 9 14 9 7 9 2 1 2 9 4 13 7 9 13 14 13 15 16 10 11 9 4 14 13 2
33 1 0 9 2 11 11 13 0 16 13 15 9 2 13 3 15 0 9 2 3 10 9 13 15 13 0 7 13 0 9 1 15 2
16 10 11 11 13 0 1 11 11 2 7 3 13 9 1 9 2
25 16 11 7 0 9 13 10 9 2 10 9 1 9 4 13 1 13 10 11 1 10 9 14 13 2
17 10 0 11 11 1 10 11 13 0 1 10 0 9 1 10 9 2
34 15 13 16 10 11 11 11 2 10 4 3 4 3 13 16 13 1 10 0 9 2 4 3 13 7 13 15 9 4 13 1 10 9 2
25 10 9 1 9 7 9 1 10 0 0 9 1 11 4 14 13 3 1 0 9 1 10 11 9 2
20 11 11 13 0 1 10 0 9 1 10 11 9 2 7 1 11 7 1 11 2
18 1 10 0 9 1 11 2 13 11 11 10 13 10 9 1 15 11 2
25 2 13 1 10 9 7 4 14 13 3 3 3 7 4 13 14 13 1 10 0 9 1 9 2 2
13 10 0 9 1 11 9 9 10 9 13 0 9 2
31 11 2 11 13 15 2 11 13 15 2 11 13 10 0 9 2 7 10 10 11 13 13 14 13 15 10 10 9 1 9 2
40 1 10 0 0 9 3 4 13 9 1 11 14 0 9 1 9 13 10 9 16 10 9 4 13 1 10 11 11 10 13 1 10 9 1 10 11 11 11 11 2
21 1 10 0 9 2 10 0 9 9 13 15 15 13 9 1 10 0 0 9 9 2
19 0 9 2 0 9 1 11 11 7 11 13 1 10 9 10 10 9 13 2
18 11 3 13 16 15 4 13 7 13 10 0 9 10 9 4 3 13 2
21 11 11 11 13 11 13 4 13 0 0 9 10 0 9 13 14 7 4 14 13 2
26 16 10 9 3 0 2 10 9 13 1 16 15 4 13 7 13 10 9 14 13 10 11 1 0 9 2
14 3 3 15 13 14 13 10 11 2 11 2 7 11 2
16 7 14 3 4 10 12 13 2 7 14 3 13 15 9 0 2
36 10 11 4 3 13 10 0 9 9 1 11 2 7 11 2 10 1 10 9 4 3 3 13 16 15 13 0 9 2 13 3 3 1 0 9 2
24 15 4 13 16 11 13 3 12 0 9 7 7 10 11 7 10 1 15 9 13 10 0 9 2
28 11 11 14 11 11 11 3 13 10 9 1 10 9 1 15 9 7 11 13 14 4 3 13 10 0 9 3 2
14 15 4 13 16 11 11 13 3 3 10 9 0 9 2
19 7 13 16 15 4 13 15 2 13 15 13 15 2 7 15 13 3 0 2
11 10 9 1 11 13 10 9 1 8 8 2
21 0 9 1 10 9 13 9 4 4 13 2 3 1 15 1 0 9 9 1 11 2
23 11 13 9 1 11 2 7 15 13 0 13 16 3 7 3 2 10 9 4 3 13 15 2
9 15 13 1 10 9 1 10 9 2
2 3 2
27 10 11 11 13 1 10 9 9 7 13 10 9 1 11 9 2 0 1 15 13 2 0 2 9 2 2 2
21 3 2 13 0 9 2 10 11 1 11 13 10 9 10 15 13 16 13 11 9 2
2 3 2
13 14 13 1 10 0 2 0 9 2 2 3 3 2
43 3 2 15 4 13 16 15 4 4 3 13 16 10 9 1 0 9 13 0 14 13 1 11 2 13 16 10 9 4 4 13 10 9 1 9 1 3 10 0 12 9 2 2
22 1 0 9 2 10 11 13 3 1 15 0 9 2 13 1 10 9 10 13 3 0 2
10 7 15 4 14 13 15 1 10 9 2
42 15 13 1 10 9 0 9 1 11 3 15 13 11 9 1 9 10 4 13 1 10 9 2 10 9 10 13 3 3 0 1 10 11 2 13 9 10 13 3 1 11 2
9 7 15 4 15 13 1 10 9 2
3 10 9 2
6 15 13 0 2 9 2
22 10 11 2 11 11 11 4 13 11 11 7 11 11 2 13 16 15 13 10 9 9 2
8 3 13 10 9 1 10 9 2
33 11 11 2 12 2 15 1 15 9 13 1 10 13 9 1 10 9 2 13 15 9 1 10 0 9 1 11 4 13 1 11 12 2
19 10 9 13 14 4 13 16 9 9 13 10 9 1 10 9 2 15 13 2
45 2 15 13 1 10 9 7 10 0 9 4 13 7 15 13 3 7 10 10 0 9 4 13 7 15 13 3 10 9 16 15 14 13 3 2 2 11 13 9 1 0 9 1 11 2
16 2 15 13 3 0 9 7 15 13 10 9 3 9 13 15 2
4 10 9 9 2
14 15 13 1 15 9 1 15 9 13 9 2 3 2 2
18 11 13 15 0 9 13 3 5 12 14 13 1 11 1 11 7 11 2
3 0 11 2
28 3 13 10 9 2 4 14 4 13 1 9 10 13 0 9 10 13 0 9 7 3 13 0 14 13 1 9 2
21 9 1 15 3 13 15 13 14 13 3 3 7 13 9 1 9 1 15 0 9 2
46 16 15 13 0 14 13 0 9 1 9 1 10 9 2 10 0 9 1 11 11 14 2 11 11 11 2 9 1 10 11 9 13 3 3 0 14 13 1 2 13 10 0 9 3 2 2
24 1 10 13 10 11 9 1 11 2 12 1 10 9 13 16 16 11 13 10 9 1 15 9 2
18 15 13 12 9 16 15 13 3 11 13 10 9 10 15 4 14 13 2
26 2 9 13 15 2 15 4 13 2 15 13 10 9 1 9 3 3 16 9 4 13 1 10 0 11 2
29 16 15 4 13 1 12 2 15 4 15 9 13 1 15 2 15 4 10 9 13 2 7 10 4 10 0 9 13 2
8 2 10 11 2 15 13 15 2
4 2 9 2 2
20 15 13 10 9 1 15 9 1 10 11 2 3 1 10 2 15 4 14 13 2
6 15 4 3 13 3 2
10 15 3 4 14 13 16 13 10 9 2
13 15 9 13 3 0 3 3 13 14 13 15 9 2
4 2 9 2 2
34 7 1 2 15 13 10 9 1 10 9 1 10 11 11 10 13 10 9 13 1 10 0 9 2 7 15 13 3 3 12 0 9 13 2
19 15 13 10 0 9 1 10 9 13 11 11 13 2 10 11 14 13 2 2
20 15 13 1 9 2 1 10 9 2 1 10 9 13 11 11 1 11 2 11 2
25 15 13 10 9 2 15 7 15 9 11 2 13 2 13 15 7 11 1 15 9 1 11 1 12 2
8 12 9 3 2 15 4 13 2
19 3 15 4 13 10 2 15 13 10 9 2 9 7 15 4 13 0 9 2
4 2 9 2 2
20 2 7 3 15 13 10 9 2 15 13 10 0 9 13 14 13 1 15 9 2
4 2 9 2 2
6 15 13 14 10 9 2
4 2 9 2 2
11 15 13 10 11 9 2 3 1 0 9 2
4 2 9 2 2
13 10 9 4 13 1 15 0 0 9 9 1 9 2
6 11 7 15 13 11 2
9 12 1 10 11 9 13 10 9 2
16 10 9 4 13 1 10 9 13 2 2 10 11 14 13 2 2
3 15 13 2
12 10 9 13 16 13 9 0 1 15 1 9 2
15 15 2 10 15 13 14 13 2 3 3 16 15 3 4 2
4 2 9 2 2
32 2 10 9 2 15 13 12 9 2 12 9 14 13 1 15 13 2 12 1 10 9 4 13 2 15 4 13 10 9 14 13 2
27 7 15 13 15 10 15 9 2 10 15 9 2 13 1 9 10 4 14 13 16 15 13 1 10 11 11 2
5 2 9 2 2 2
7 3 15 13 10 0 9 2
23 7 15 13 14 13 2 4 15 13 16 15 3 13 10 9 13 2 10 11 14 13 2 2
20 15 13 10 9 1 15 2 9 2 2 9 2 13 1 9 11 11 1 12 2
17 15 4 13 0 9 16 11 13 10 0 9 7 5 7 13 11 2
11 15 13 0 16 11 4 13 1 9 9 2
25 15 4 13 11 2 11 2 11 11 2 11 2 11 2 7 9 9 9 11 2 3 3 14 11 2
34 15 13 10 0 9 2 7 15 4 4 13 9 9 10 3 13 16 11 13 3 0 16 13 0 9 1 10 13 9 9 9 1 11 2
10 11 11 13 10 0 9 1 11 11 2
6 15 13 15 1 11 2
26 1 1 11 12 2 12 2 15 9 1 9 13 1 10 11 11 1 11 2 11 1 11 11 2 11 2
40 15 9 1 11 7 10 11 9 4 13 3 0 2 15 4 13 13 3 10 0 9 16 15 4 13 3 2 1 10 0 9 1 0 12 2 12 7 12 9 2
21 15 13 0 0 2 9 1 10 9 1 11 2 10 11 9 7 9 9 1 0 2
7 15 3 13 15 1 11 2
3 6 11 2
23 15 3 13 14 13 10 0 2 9 2 2 1 11 11 11 15 13 15 1 11 10 9 2
6 12 4 13 14 13 2
11 11 11 13 10 9 1 11 12 2 12 2
7 15 7 10 0 2 11 2
23 13 1 10 9 1 11 14 9 9 2 15 13 15 4 13 16 15 4 13 11 3 3 2
17 1 11 2 15 4 3 13 3 3 0 1 10 11 9 7 9 5
3 13 1 11
10 11 13 10 9 1 11 12 2 12 2
13 15 13 14 13 10 9 14 13 11 11 1 11 2
22 11 4 13 12 1 10 3 0 9 1 10 9 1 11 9 1 10 0 0 9 2 2
7 0 14 13 15 1 9 2
33 3 2 9 1 15 4 4 13 1 11 1 10 0 9 2 7 15 13 10 0 9 16 15 13 10 9 14 13 15 13 1 9 2
30 1 10 9 2 13 10 9 13 15 14 13 16 11 4 4 13 10 9 10 9 10 13 10 11 2 11 5 11 9 2
39 16 15 4 14 3 13 10 11 9 11 2 15 4 13 10 0 9 7 13 10 0 9 1 9 16 13 1 11 11 7 11 11 2 1 9 1 11 11 2
19 1 10 9 11 7 11 2 11 2 13 10 0 0 9 1 9 1 12 2
8 15 13 12 9 2 13 9 2
10 10 9 11 13 13 10 0 9 3 2
24 3 12 0 9 2 15 13 14 0 2 3 3 16 15 13 2 16 11 14 2 13 2 11 2
30 15 3 13 9 14 13 15 2 13 15 2 7 13 10 9 1 10 9 2 15 13 15 10 0 0 9 9 13 1 2
75 15 13 0 14 13 16 11 4 13 15 15 4 14 7 13 7 13 10 9 1 10 3 0 0 9 3 3 2 16 13 1 10 13 9 1 11 9 2 15 4 13 10 13 9 1 10 9 2 7 13 2 14 16 15 13 15 13 14 2 16 15 9 4 4 13 1 10 0 9 1 10 11 9 9 2
16 15 13 10 9 1 0 9 9 10 13 0 0 9 9 0 2
8 0 9 1 10 9 1 11 2
5 9 1 10 9 2
8 11 2 15 15 13 13 9 2
23 13 0 9 9 13 10 9 10 0 9 16 13 7 13 10 9 10 0 9 9 4 13 2
25 15 3 13 0 9 1 10 9 16 13 10 0 9 7 13 14 13 10 0 9 9 7 9 9 2
39 10 11 9 14 13 10 9 1 11 11 2 11 14 9 3 12 9 16 10 11 11 11 13 1 1 9 13 14 4 13 1 10 9 1 0 9 1 9 2
32 3 4 10 11 13 1 10 9 3 15 4 13 3 0 11 2 15 13 3 0 1 10 9 1 11 11 2 1 10 11 11 2
33 3 15 13 13 0 0 0 7 0 9 3 2 1 10 9 3 11 9 4 13 1 10 0 9 7 13 14 13 15 9 1 9 2
26 1 10 9 3 10 0 2 0 7 0 9 13 3 0 16 13 2 7 10 11 13 0 14 13 0 2
15 12 9 13 16 10 11 13 10 11 11 16 13 10 11 2
12 11 13 10 9 1 9 1 0 9 7 9 2
15 10 9 1 10 11 1 11 3 13 3 14 13 9 1 2
35 11 2 11 7 11 13 10 11 1 9 2 0 1 15 13 10 0 9 2 10 11 2 7 10 9 1 0 9 2 7 9 1 15 2 2
11 15 3 13 11 11 11 9 1 11 11 2
23 2 3 3 4 10 0 0 11 11 9 4 13 3 14 13 14 13 13 1 10 9 2 2
50 10 9 1 10 11 13 10 9 1 0 9 7 0 9 15 13 14 13 1 10 0 9 2 13 11 2 9 0 9 9 2 10 9 1 9 9 1 11 2 7 3 3 13 10 9 1 1 12 9 2
27 10 11 11 14 15 13 15 1 11 1 11 13 13 10 0 9 7 3 0 2 9 1 0 1 10 11 2
47 11 11 11 9 11 11 2 15 13 0 1 10 11 9 2 13 1 11 12 2 12 2 16 10 0 9 1 10 11 9 1 10 11 11 13 14 2 13 11 2 2 13 1 10 11 11 2
11 15 4 3 13 10 0 9 1 10 11 2
19 7 15 4 14 13 1 1 9 0 3 3 16 15 4 13 1 0 9 2
30 9 1 10 11 13 3 7 13 1 9 14 13 15 1 16 13 15 9 7 13 12 9 9 7 13 3 9 1 11 2
19 15 13 7 0 9 7 4 13 1 0 0 9 10 4 3 4 13 1 2
44 15 13 10 0 0 9 2 8 8 8 8 8 2 9 13 1 9 2 3 9 4 13 1 9 2 2 7 15 13 13 10 9 10 9 16 15 4 14 13 14 13 1 15 2
17 7 3 2 3 3 2 3 9 13 1 9 15 13 1 1 9 2
41 3 15 4 3 3 3 13 3 1 15 2 15 13 3 0 2 13 10 9 9 1 10 11 7 1 10 0 9 1 10 11 11 16 1 11 12 11 13 1 11 2
32 2 10 0 0 0 9 4 13 9 1 10 0 0 9 11 7 13 16 15 4 4 13 10 9 14 2 9 9 2 1 11 2
46 2 15 4 13 7 15 13 15 9 1 9 10 11 11 13 1 14 13 1 11 2 2 0 9 11 11 2 11 13 11 1 10 9 1 11 2 10 9 1 10 0 0 0 9 11 2
14 0 9 2 11 13 16 15 9 4 13 9 1 11 2
43 2 13 2 11 2 13 15 15 9 9 1 11 16 10 9 1 11 7 11 13 10 0 2 2 11 2 11 13 1 10 11 9 9 1 11 2 15 9 9 3 1 11 2
12 15 4 13 16 15 15 13 1 10 9 2 2
41 7 1 11 12 15 0 9 1 11 4 3 13 1 1 12 0 9 1 15 9 2 7 10 11 9 4 13 1 0 9 1 15 9 2 10 13 12 11 9 0 2
16 10 11 13 0 14 13 7 13 2 7 15 13 15 7 3 2
24 15 13 14 3 1 11 7 15 4 4 13 1 15 10 9 16 13 15 10 11 4 4 13 2
20 11 11 1 10 11 11 13 16 10 9 1 10 9 4 4 13 9 8 3 2
8 3 4 15 3 13 1 11 2
15 15 4 14 13 16 11 13 14 13 3 0 7 13 1 2
15 15 3 4 13 10 9 2 3 10 0 4 3 13 3 2
8 11 2 15 13 3 2 6 2
8 9 3 1 0 9 1 9 2
9 15 4 13 11 14 1 3 12 2
3 13 15 13
8 15 4 14 13 15 15 13 2
6 3 4 15 13 1 2
2 11 2
3 13 1 2
15 4 15 13 0 16 15 13 14 10 0 9 15 15 13 2
13 15 4 13 3 9 14 13 0 16 9 13 0 2
16 11 11 13 15 9 9 7 15 7 15 9 4 13 14 13 2
8 11 7 11 4 13 1 15 2
5 13 15 1 12 2
10 15 4 14 13 1 15 1 10 9 2
26 13 15 1 15 9 2 9 1 10 9 1 2 2 7 11 2 15 13 1 0 9 7 13 0 9 2
22 1 9 11 7 15 4 13 16 3 0 15 10 13 16 15 13 1 15 9 0 9 2
4 0 9 2 2
10 15 13 14 13 1 9 2 13 11 2
13 15 4 14 13 3 1 15 7 4 14 13 11 2
10 10 13 9 15 4 13 0 14 13 2
10 15 13 15 13 10 9 7 10 9 2
11 15 13 15 4 13 15 9 13 1 9 2
11 15 13 16 15 13 9 9 15 4 13 2
7 15 4 13 10 9 9 2
20 6 2 15 4 14 13 7 6 15 4 14 13 15 1 1 10 11 11 9 2
11 15 13 15 16 15 13 3 0 7 0 2
13 15 13 9 1 9 15 13 12 7 15 13 15 2
8 3 4 15 13 15 13 0 2
4 4 15 13 2
7 3 4 15 13 10 9 2
7 10 9 13 14 3 0 2
13 4 15 13 15 13 0 1 1 10 11 11 9 2
7 2 11 11 2 2 8 2
3 12 12 9
2 10 2
37 15 13 15 9 2 1 0 9 1 10 11 14 9 16 10 11 4 13 11 11 14 3 13 10 9 14 13 10 9 9 14 13 1 0 9 9 2
36 10 9 1 10 10 9 4 13 13 16 16 15 3 13 9 14 9 1 0 9 3 2 15 13 1 10 9 10 10 0 9 9 4 13 1 2
8 1 0 9 10 9 4 13 2
10 13 15 9 1 3 10 9 4 13 2
46 8 10 11 9 13 14 13 10 0 9 9 1 10 9 16 13 14 13 3 10 7 10 9 4 13 10 9 1 10 9 3 1 13 10 0 9 13 3 0 9 4 13 1 10 9 2
30 15 3 13 10 9 10 3 0 0 9 14 13 15 3 7 3 0 9 4 13 16 13 14 13 16 15 13 0 9 2
6 9 13 3 9 13 2
12 15 4 14 13 3 1 10 9 1 11 3 2
3 15 13 3
2 9 2
26 11 11 11 11 2 11 9 2 9 2 11 2 12 2 9 2 12 2 9 2 12 2 9 2 12 8
5 15 9 9 13 8
5 2 11 2 11 2
12 15 9 13 14 13 10 9 1 11 14 9 2
28 15 4 13 10 9 3 7 3 15 4 13 15 14 13 1 1 15 1 10 9 1 10 9 9 3 10 9 2
8 7 15 4 13 3 13 15 2
16 10 9 13 1 10 13 9 3 7 4 13 0 7 0 9 2
18 16 15 4 13 15 1 9 2 6 13 10 9 3 7 13 10 9 2
11 10 0 9 1 10 9 1 15 4 13 2
8 3 13 15 1 15 9 9 2
13 15 4 13 1 0 9 1 9 14 13 7 13 2
8 15 4 15 13 15 13 0 2
9 6 2 15 13 10 0 0 9 2
8 15 13 15 3 15 13 3 2
7 15 13 15 9 1 9 2
2 8 8
3 12 12 9
20 15 3 13 14 13 15 10 0 9 14 13 15 13 16 15 13 3 1 3 2
37 9 13 15 0 9 1 10 9 3 1 11 2 7 1 10 13 9 2 15 4 13 1 10 0 9 1 9 1 10 9 9 9 1 11 11 11 2
20 15 13 3 3 2 7 15 13 14 13 0 16 15 13 9 13 16 15 13 2
31 15 4 14 13 10 9 9 3 1 15 0 9 2 7 16 15 13 14 13 15 2 15 4 13 3 1 8 7 1 12 2
26 15 13 13 1 10 1 15 1 10 0 12 9 1 11 2 11 2 7 15 13 15 10 1 10 0 2
3 13 9 2
2 11 11
25 9 2 15 13 10 0 9 9 1 11 1 11 11 2 3 3 1 10 11 9 2 13 1 12 2
9 16 15 4 13 15 2 6 13 2
7 8 8 8 1 12 12 9
6 11 2 11 7 11 2
23 3 13 14 13 15 9 1 11 11 9 1 12 5 12 14 13 11 1 11 14 9 9 2
8 15 4 13 11 14 9 11 12
9 15 13 3 16 13 15 10 3 2
2 3 2
1 11
17 11 11 11 11 11 2 11 9 2 12 2 12 9 2 12 2 12
2 11 11
3 12 12 9
15 4 15 4 13 10 9 9 1 9 13 2 9 13 1 2
11 6 13 15 3 1 8 2 13 1 15 2
2 9 2
2 9 2
1 11
10 2 8 2 13 10 13 9 1 12 12
7 15 4 13 15 9 9 2
7 15 0 9 9 13 8 2
18 1 0 9 2 15 9 4 13 1 0 0 9 7 0 9 7 9 2
9 3 13 12 9 2 8 7 8 2
12 16 15 13 10 9 2 6 13 15 1 8 2
1 5
27 2 10 9 13 4 13 3 1 10 9 7 9 1 10 15 4 13 7 4 13 0 7 2 7 0 9 2
34 10 9 2 9 2 9 7 0 9 1 2 7 9 1 10 9 1 9 1 2 10 9 1 9 7 9 0 1 10 13 9 4 13 2
20 16 15 13 15 1 9 2 6 13 10 9 7 13 10 9 1 10 9 2 2
1 5
10 13 6 13 10 11 9 1 11 9 2
23 3 2 15 4 13 10 9 9 2 9 1 10 9 1 10 9 1 9 1 10 9 9 2
1 2
10 4 14 13 14 13 15 1 10 9 2
1 2
3 0 9 2
1 2
1 5
13 11 11 0 9 2 12 0 9 2 12 9 2 8
1 2
2 2 9
2 11 11
3 12 12 9
11 15 13 1 11 11 1 11 13 15 9 2
14 11 13 11 0 13 12 9 15 10 13 3 1 11 2
20 3 2 15 3 13 15 13 10 0 9 2 10 13 0 1 10 3 0 9 2
12 15 13 10 9 1 10 9 1 10 0 9 2
23 15 3 13 16 10 0 12 9 13 10 0 9 3 13 0 9 1 10 13 11 9 9 2
23 11 13 10 0 9 16 13 9 1 10 9 2 15 13 11 4 13 7 4 13 10 9 2
11 11 16 15 4 6 13 9 7 13 3 2
2 9 2
1 11
4 3 15 13 2
12 16 15 13 10 0 9 2 6 13 15 13 2
2 11 11
3 12 12 9
2 8 8
3 12 12 9
5 8 1 12 12 9
27 10 9 13 3 4 13 1 9 10 15 13 14 13 0 2 7 15 4 14 13 16 15 13 0 7 0 2
25 9 13 3 4 4 13 1 10 9 14 13 7 10 9 1 10 9 14 13 10 0 9 13 3 2
11 10 9 13 3 13 3 15 1 10 9 2
34 1 0 2 15 4 13 1 0 9 1 15 1 2 7 13 7 13 1 1 9 1 11 11 7 15 9 2 9 2 9 7 9 2 2
3 12 11 11
26 10 9 13 3 1 10 3 0 9 1 11 11 12 7 15 4 13 3 1 11 11 11 12 7 0 2
12 11 11 11 12 4 4 13 1 0 1 8 2
49 2 13 13 9 2 9 2 2 13 13 9 2 9 2 2 13 13 9 2 9 2 2 13 13 9 2 9 2 2 13 13 9 2 9 2 2 13 13 9 2 9 2 2 13 13 9 2 9 2
2 2 9
2 2 9
2 2 9
2 2 9
2 2 9
2 2 9
2 2 9
2 11 11
3 12 12 9
19 1 7 1 11 12 2 12 10 9 1 9 4 13 1 10 3 13 9 2
15 10 9 13 1 10 0 9 9 9 7 12 9 9 9 2
12 10 9 4 13 1 10 9 2 11 2 11 2
36 1 7 1 11 12 2 12 2 11 11 2 0 9 9 1 11 2 11 2 12 2 12 2 13 7 13 15 16 10 9 4 13 11 2 11 2
52 3 2 15 13 15 16 9 12 1 10 9 2 10 13 1 0 2 9 13 0 1 9 7 0 9 1 10 9 2 4 4 13 16 10 9 10 10 9 4 4 13 1 9 4 7 2 7 13 0 1 9 2
24 15 4 13 14 13 10 9 7 10 4 4 13 1 15 1 10 0 9 7 9 1 9 12 2
12 13 13 10 9 1 10 0 9 1 9 12 2
1 11
11 11 4 13 15 14 13 1 10 0 9 2
2 9 2
3 11 11 11
8 11 2 6 13 10 13 9 2
8 10 0 7 13 9 4 13 2
21 15 13 10 9 13 1 15 9 7 13 10 9 13 9 10 15 4 3 3 13 2
8 15 13 0 14 13 10 9 2
13 13 15 13 16 0 7 15 4 13 3 7 13 2
2 9 2
8 2 11 2 11 2 2 8 2
3 12 12 9
2 11 2
6 15 4 13 1 9 2
4 11 13 0 2
7 15 13 15 1 10 9 2
9 11 13 3 4 13 10 0 9 2
18 15 4 14 13 3 0 2 9 2 15 4 13 1 10 12 9 9 2
6 3 13 15 9 9 2
9 10 9 1 10 9 13 3 0 2
6 4 15 3 13 15 2
6 13 15 13 3 3 2
7 15 0 9 13 0 3 2
9 15 0 9 4 13 1 10 9 2
5 15 13 1 9 2
4 13 1 15 3
1 11
5 3 4 15 13 2
6 4 15 13 10 9 2
6 15 13 0 1 15 2
11 13 3 7 13 1 11 16 15 13 0 2
2 11 11
3 12 12 9
3 11 11 11
2 9 2
5 15 4 3 13 2
7 2 3 13 10 0 9 2
14 10 13 4 13 10 9 1 10 9 9 1 11 9 2
6 9 1 10 15 13 2
6 15 4 13 1 9 2
4 9 9 9 2
8 9 9 12 2 9 2 11 11
11 11 11 2 11 11 2 11 11 2 11 11
8 9 9 12 2 9 2 11 11
11 11 11 2 11 11 2 11 11 2 11 11
4 9 9 9 2
8 9 9 12 2 9 2 11 11
11 11 11 2 11 11 2 11 11 2 11 11
30 13 9 2 9 9 12 2 9 2 11 11 11 11 2 9 2 11 11 2 9 2 11 11 2 9 2 11 11 2 9
16 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11
9 15 13 14 13 9 1 11 11 2
5 15 13 15 13 2
4 3 14 13 2
11 10 9 15 13 3 0 14 13 15 9 2
27 3 13 3 10 13 11 11 9 2 8 7 13 3 1 11 11 7 11 7 13 3 1 1 10 9 9 2
15 10 9 4 13 15 3 1 11 14 11 11 12 9 9 2
16 6 13 2 15 9 13 14 4 13 3 2 15 3 13 9 2
5 10 0 9 9 2
32 9 2 16 15 13 10 9 13 10 9 9 2 6 13 11 11 2 12 2 2 11 11 2 12 2 7 11 11 2 12 2 2
10 15 13 16 7 11 7 11 13 3 2
13 9 9 1 12 2 15 13 9 14 13 10 9 2
20 15 4 14 13 10 0 9 3 15 13 11 7 15 4 13 14 13 1 9 2
14 10 9 4 13 14 13 0 2 11 4 3 13 9 2
2 11 11
3 12 12 9
6 4 15 13 1 9 2
12 3 2 15 13 10 9 1 10 9 10 9 2
7 4 15 13 14 4 13 2
17 1 10 9 2 13 15 3 16 15 4 13 1 12 1 9 9 2
12 15 9 3 13 1 15 2 15 4 15 13 2
9 7 2 15 13 3 0 1 15 2
4 3 13 15 2
6 10 9 1 11 11 2
1 6
2 2 11
7 0 14 13 10 13 0 2
24 15 13 14 13 16 15 13 10 9 13 1 10 9 4 13 15 9 1 1 15 9 0 9 2
12 15 13 14 16 13 10 9 1 9 1 9 2
7 15 13 3 1 10 9 2
3 13 3 2
3 13 9 2
3 13 0 2
6 9 1 15 13 0 2
30 13 3 1 11 1 3 10 9 10 13 10 0 0 16 15 13 15 4 4 13 3 7 3 9 13 15 13 14 13 2
3 13 9 2
23 15 4 14 13 1 15 1 9 7 3 15 13 15 1 10 10 9 13 2 9 13 9 2
10 9 16 13 1 15 14 13 15 1 2
6 15 3 13 13 15 2
10 15 3 13 1 0 9 1 10 9 2
12 15 13 10 0 9 9 1 15 10 13 3 2
6 15 13 3 0 9 2
7 3 4 9 13 1 15 2
5 4 15 13 11 2
5 11 4 13 0 2
8 13 1 3 4 13 3 0 2
14 9 1 3 13 14 13 10 9 0 9 1 0 9 2
14 11 13 0 7 4 13 15 10 3 0 9 1 9 2
4 13 1 9 2
1 11
4 11 11 11 8
1 5
9 13 15 0 9 1 11 11 1 8
17 1 15 15 13 14 1 9 7 13 15 9 14 9 1 15 9 2
7 15 13 3 1 10 9 2
6 13 3 7 13 3 2
1 9
1 11
12 9 15 4 13 3 1 11 1 3 10 9 2
12 11 13 14 13 0 14 13 15 3 1 9 2
9 15 4 3 3 13 3 1 15 2
11 13 15 13 0 9 15 13 11 11 3 2
2 11 11
3 12 12 9
4 1 15 9 2
7 2 13 13 9 2 9 2
3 2 9 2
22 10 9 7 2 7 9 4 13 10 0 9 2 9 9 7 4 3 13 0 7 0 2
36 16 15 13 14 10 13 9 2 15 4 3 13 16 15 4 13 10 9 1 9 2 10 9 2 9 2 9 7 9 1 10 9 4 3 13 2
40 16 15 4 13 10 9 7 2 7 9 1 9 2 6 13 15 3 1 9 7 1 9 2 13 15 3 1 12 12 2 7 3 13 10 9 7 10 15 9 2
3 13 15 2
7 2 9 2 9 2 9 2
11 15 4 13 16 13 15 1 10 9 9 2
16 15 4 3 13 10 9 7 13 15 14 13 15 3 10 9 2
13 3 1 9 9 1 10 9 7 9 1 10 9 2
4 11 11 12 2
18 14 0 16 15 4 13 14 13 12 9 7 12 9 9 1 10 9 2
2 9 2
15 15 4 3 13 1 10 9 13 0 2 0 7 0 9 2
25 15 0 9 4 13 10 9 1 10 0 9 1 10 15 4 13 9 2 9 2 9 7 0 9 2
33 15 4 3 4 13 16 2 0 9 13 3 1 10 9 2 2 7 3 2 16 15 4 14 13 15 1 3 2 15 3 3 4 2
22 1 10 9 3 4 13 2 7 3 15 3 13 0 9 10 15 4 13 14 13 1 2
28 15 4 3 13 14 13 15 9 1 10 9 7 9 10 4 13 15 0 9 7 10 4 13 15 0 9 9 2
64 15 13 15 9 1 15 9 2 7 16 15 13 10 0 9 15 13 0 14 13 15 10 2 9 7 9 2 1 10 10 10 13 15 10 0 9 2 7 13 9 2 15 4 13 16 15 4 4 3 13 1 10 0 2 7 15 13 13 15 3 0 1 9 2
15 15 15 13 14 13 2 9 3 13 14 4 13 15 3 2
7 15 13 10 9 1 15 2
40 15 13 10 0 9 7 10 15 13 1 9 2 1 10 9 2 13 10 9 15 15 4 13 7 1 15 15 4 2 3 2 13 10 9 1 9 13 1 9 2
19 15 13 15 0 9 2 7 15 13 9 1 9 2 14 13 15 0 9 2
23 15 13 10 9 1 2 12 2 9 2 7 10 15 13 13 9 7 2 0 2 9 2 2
18 15 13 14 4 13 1 9 2 10 0 9 7 10 0 9 1 9 2
19 1 9 15 3 4 14 13 14 13 0 1 10 9 1 10 9 7 9 2
20 10 15 13 13 16 2 15 2 14 13 3 1 15 2 7 14 13 15 0 2
2 11 2
17 0 16 3 13 15 1 15 3 2 3 13 14 13 15 11 2 2
14 0 9 13 1 10 0 9 1 10 9 1 10 9 2
9 13 15 13 16 15 13 10 9 2
2 11 2
3 6 11 2
18 4 15 3 13 10 0 9 9 9 10 15 13 1 11 14 9 9 2
10 16 15 13 4 15 13 15 10 9 2
2 9 2
1 11
31 13 4 10 0 9 1 9 0 14 13 10 10 2 9 9 9 1 12 9 2 11 2 1 10 11 11 11 2 0 9 2
32 16 15 4 13 1 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 7 11 2 15 4 13 10 0 9 1 8 2
2 11 2
19 15 13 1 9 1 11 9 1 11 9 7 15 4 14 13 15 9 3 2
19 15 13 14 13 15 1 10 11 9 2 9 2 7 10 9 13 3 0 2
17 13 15 0 16 15 7 9 0 1 10 9 9 13 10 9 9 2
6 15 4 3 13 15 2
3 13 15 2
4 11 11 9 12
8 2 11 2 11 2 2 8 2
3 12 12 9
4 0 9 11 2
19 15 4 13 10 13 9 1 10 9 9 7 0 9 1 15 9 7 9 2
18 15 13 13 10 9 1 10 9 9 9 7 13 9 1 15 1 11 2
43 1 9 2 15 13 9 1 15 9 9 16 10 9 1 10 9 9 1 11 1 2 11 4 13 1 1 9 2 4 15 13 15 4 13 15 1 11 10 15 4 13 1 2
9 3 13 15 0 9 1 10 9 2
10 15 13 3 1 15 9 1 10 9 2
2 9 2
27 11 11 11 11 11 2 11 2 2 11 2 2 12 11 11 9 12 11 2 11 12 9 12 9 12 9 8
11 9 2 4 15 13 9 9 9 10 9 2
19 15 7 9 4 13 3 7 9 1 10 9 13 1 9 9 2 2 2 2
11 3 1 15 9 2 6 13 13 9 9 2
22 1 15 9 2 6 13 15 10 9 14 13 10 9 7 9 15 4 13 13 10 9 2
20 2 13 0 9 2 8 8 8 8 8 8 9 2 2 13 13 9 2 9 2
2 9 2
2 11 11
7 2 8 8 8 8 8 9
13 15 4 13 15 9 1 1 9 9 1 10 9 2
5 15 4 13 15 2
11 15 13 1 10 9 16 13 15 0 9 2
3 0 9 2
2 11 11
18 11 11 2 15 4 13 1 11 11 11 7 1 15 9 1 10 9 2
2 11 11
14 6 13 2 9 2 4 15 13 9 1 11 3 3 2
1 9
1 11
2 11 11
3 13 9 12
2 11 11
17 10 0 9 15 4 13 13 10 9 9 9 1 2 9 1 11 2
10 6 13 15 13 16 15 13 9 0 2
1 11
2 11 11
2 11 2
8 13 4 10 9 1 10 9 2
13 16 15 13 15 13 9 13 1 11 1 9 9 2
11 6 13 15 13 3 15 4 13 14 13 2
3 0 9 2
2 11 11
2 11 11
2 11 2
15 15 4 14 13 10 9 2 0 9 9 2 1 15 9 2
13 10 9 2 0 9 9 2 4 13 1 0 9 2
8 4 15 13 15 15 4 13 2
2 9 2
2 11 11
8 13 13 13 9 12 9 3 2
1 11
2 11 11
2 11 11
6 15 13 0 1 15 2
11 13 3 7 13 1 11 16 15 13 0 2
2 11 11
3 12 12 9
3 13 9 12
2 11 11
2 11 2
20 15 13 0 2 15 4 13 10 0 9 7 13 15 10 9 16 13 9 9 2
3 0 9 2
2 11 11
1 9
2 11 11
2 11 2
11 16 13 2 13 4 10 9 9 1 11 2
15 16 15 4 13 15 13 0 9 13 0 9 1 11 11 2
23 15 13 0 14 13 10 11 9 7 0 9 9 3 2 15 4 13 9 7 9 9 9 2
6 4 15 13 10 9 2
1 11
2 11 11
2 11 11
3 11 11 11
3 12 12 9
4 11 11 2 8
3 12 12 9
2 11 2
17 6 13 13 10 9 9 1 10 9 9 9 1 10 3 13 9 2
8 6 13 9 7 13 1 9 2
1 9
3 11 12 2
2 11 2
14 6 13 10 9 1 10 11 11 11 9 1 15 9 2
9 10 9 4 13 11 12 2 12 2
2 9 2
2 11 11
8 15 4 13 9 1 10 11 2
2 11 11
2 11 2
5 9 1 15 9 2
17 4 15 13 15 10 9 15 13 2 15 4 13 10 9 1 15 2
1 11
3 0 10 2
6 15 9 13 11 11 2
31 15 13 14 13 11 11 1 10 9 1 15 9 2 10 11 16 13 7 11 13 11 11 2 7 15 4 13 15 10 9 2
37 15 4 3 13 10 11 9 9 9 13 0 0 9 13 9 9 9 7 4 13 15 9 2 13 10 0 1 11 11 2 14 13 10 9 9 9 2
22 15 13 11 0 2 0 9 1 12 11 2 12 5 12 11 12 13 3 12 9 9 2
22 3 2 10 9 1 0 0 9 13 14 16 13 1 1 0 9 1 7 9 7 9 2
9 10 9 7 0 9 13 16 13 2
7 9 2 5 12 2 12 2
6 9 2 12 2 12 2
4 9 9 2 12
18 3 15 4 14 13 10 9 9 9 16 10 13 9 13 10 0 9 2
13 15 4 3 13 0 9 7 10 9 13 10 0 2
13 15 4 4 13 16 15 4 13 15 1 10 9 2
3 0 9 2
1 11
16 13 15 0 9 1 11 11 1 8 2 9 2 2 8 2 2
2 11 2
15 6 13 11 11 2 8 12 2 13 10 9 1 10 9 2
1 11
2 11 2
2 9 2
12 15 13 10 0 9 13 10 10 9 15 13 2
1 11
2 11 2
12 9 1 10 9 13 10 0 9 1 15 9 2
32 3 3 2 15 13 1 10 9 16 13 7 15 0 9 9 7 15 9 9 7 4 4 13 10 9 1 10 9 1 10 9 2
20 16 15 4 13 3 1 10 9 15 4 13 0 14 13 10 9 1 10 9 2
50 15 15 4 13 14 13 1 10 9 13 13 10 9 1 11 11 2 15 13 0 1 11 11 7 13 15 14 13 11 14 9 7 13 10 9 1 15 1 10 9 16 15 4 13 14 13 15 1 9 2
19 3 15 13 10 9 9 2 15 4 13 10 9 7 13 15 1 15 9 2
6 13 15 0 1 15 2
6 13 10 13 0 1 15
2 13 9
1 11
2 11 2
8 15 4 13 11 11 1 11 2
14 12 1 10 9 13 16 15 13 0 1 10 9 9 2
12 15 13 3 1 10 3 0 9 2 3 0 2
9 15 4 13 15 1 10 9 9 2
1 11
5 0 11 11 11 2
2 6 2
5 3 4 15 13 2
11 15 13 15 13 10 0 9 3 1 9 2
14 15 13 10 0 9 14 13 1 11 7 15 9 9 2
6 13 15 1 15 9 2
14 15 4 3 13 15 9 7 9 9 3 1 10 9 2
16 3 2 15 13 15 14 13 10 9 1 9 7 9 9 3 2
8 10 9 13 15 15 4 13 2
31 3 2 15 13 10 0 9 16 15 14 13 14 13 15 15 4 13 1 10 9 7 15 15 13 14 3 13 1 1 9 2
15 15 4 13 3 16 13 1 15 3 7 13 10 0 9 2
3 13 15 2
1 2
31 11 11 0 9 7 9 1 9 11 11 1 11 11 1 11 7 11 11 9 9 2 8 8 9 2 12 9 2 13 3 2
1 2
7 2 9 2 9 2 9 2
7 2 9 2 9 2 9 2
1 3
1 11
12 9 11 2 6 2 13 11 7 13 10 9 2
2 11 2
14 15 4 13 14 13 10 9 14 13 1 10 9 9 2
12 11 11 7 11 11 4 13 14 13 3 3 2
12 10 9 1 12 9 7 3 4 13 1 15 2
10 6 13 15 13 10 9 15 4 13 2
3 13 15 2
1 11
2 11 2
18 10 9 13 1 13 9 15 4 13 1 1 10 9 13 10 9 9 2
31 10 9 10 9 9 13 2 10 9 9 1 15 9 9 4 4 13 1 10 13 9 9 10 9 13 9 1 10 9 9 2
25 1 0 2 15 4 13 0 9 13 10 0 9 1 0 9 9 10 9 0 16 13 10 9 9 2
21 15 4 4 13 10 9 13 1 15 12 9 2 12 9 7 9 1 0 9 2 2
19 16 15 4 13 14 13 10 9 1 10 0 9 2 15 4 13 0 9 2
7 6 13 15 13 15 9 2
18 16 15 13 2 15 13 1 10 9 16 13 9 9 1 11 1 11 2
22 1 0 2 15 13 10 9 2 11 11 2 13 1 15 14 13 7 13 1 9 9 2
24 15 4 13 15 9 9 1 10 9 9 2 3 3 0 1 15 2 7 10 0 9 9 9 2
26 16 15 4 13 2 15 4 13 1 10 9 9 1 15 2 15 2 7 11 14 13 1 10 9 9 2
14 6 13 15 13 10 9 7 9 10 13 0 1 15 2
2 9 2
1 11
2 11 2
14 13 15 16 13 1 1 10 9 1 13 9 9 9 2
12 15 13 0 16 10 9 4 4 13 1 9 2
22 3 2 15 3 4 14 13 10 9 4 4 13 14 13 10 9 7 13 3 0 9 2
6 10 9 9 1 12 2
53 11 1 11 11 13 2 10 9 1 10 9 2 7 13 9 9 4 4 13 1 10 13 9 1 11 11 0 9 1 10 11 12 1 10 9 1 9 2 7 0 9 4 4 13 1 9 1 11 11 0 9 2 2
16 4 15 13 15 13 10 9 7 13 1 10 9 1 15 9 2
3 13 15 2
2 11 11
11 13 15 13 3 15 13 10 9 1 11 2
15 15 4 13 14 13 9 1 10 5 12 1 5 12 9 2
17 15 4 13 14 13 10 9 7 10 9 1 10 9 14 4 13 2
15 15 13 15 9 16 10 9 4 4 13 7 13 1 9 2
17 16 15 4 13 9 14 13 1 0 9 3 15 4 13 14 13 2
13 11 13 0 14 13 3 10 9 9 1 10 9 2
19 16 10 9 13 2 15 13 16 15 13 14 13 3 7 13 1 10 9 2
6 3 9 4 13 3 2
1 11
4 9 2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 11
2 11 2
16 15 13 15 10 9 1 12 11 11 11 1 10 11 9 9 2
32 10 9 13 1 3 16 15 13 1 15 14 13 15 13 16 10 11 11 11 11 7 10 9 9 1 11 7 11 4 3 13 2
10 13 15 13 15 15 13 1 10 9 2
13 3 2 13 15 13 1 10 0 9 1 9 9 2
1 11
2 11 2
7 13 10 9 1 10 9 2
15 15 13 14 13 10 9 1 10 11 11 7 11 9 9 2
10 13 15 3 15 9 3 13 10 9 2
7 10 11 9 13 3 0 2
1 11
2 11 2
13 15 13 0 1 10 9 15 4 13 1 10 9 2
9 15 4 13 0 14 13 1 15 2
1 11
13 13 15 13 10 9 7 13 0 14 13 3 3 2
6 13 14 13 15 3 2
3 10 11 11
26 10 15 13 14 13 13 13 1 1 12 0 9 2 0 1 9 2 7 3 13 1 10 9 9 9 2
3 3 0 2
3 9 2 8
3 9 13 2
23 7 15 13 15 13 10 0 9 1 11 11 6 16 10 9 13 0 13 15 15 9 7 9
1 13
3 9 2 8
19 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9
8 10 9 4 13 1 1 11 2
14 15 13 10 9 1 11 7 13 1 9 9 1 11 2
4 13 15 1 2
23 2 2 15 13 10 9 3 3 0 2 3 0 2 3 0 7 3 0 1 10 9 2 2
2 2 11
7 1 9 10 13 1 15 2
4 0 1 9 2
20 13 13 9 9 2 8 7 13 9 9 1 9 2 9 7 10 0 9 9 2
11 0 9 1 9 2 9 9 7 0 9 2
7 1 9 10 13 1 15 2
4 0 1 9 2
31 13 13 9 9 2 8 7 13 9 9 1 9 2 9 7 10 0 9 9 2 0 9 1 9 2 9 9 7 3 9 2
20 13 1 0 9 9 2 9 13 11 11 11 2 10 11 9 2 1 11 9 2
20 1 10 0 9 2 11 2 13 2 15 9 1 10 9 7 13 0 0 9 2
3 10 11 11
8 3 10 9 10 13 1 15 2
4 6 2 6 2
1 5
15 13 11 11 14 11 11 1 10 10 9 7 9 2 2 2
11 11 11 14 11 11 4 13 1 2 2 2
1 9
3 12 9 9
9 5 12 13 3 1 15 11 9 2
23 13 15 0 9 10 4 13 10 9 1 5 12 7 5 12 9 13 3 1 15 11 9 2
15 10 15 13 14 13 13 13 10 9 7 13 15 9 13 2
45 13 15 16 13 15 14 13 1 1 15 0 9 2 3 13 15 9 7 0 9 9 13 16 10 0 9 2 1 10 0 3 0 9 1 11 11 2 13 0 1 9 1 15 9 2
4 13 10 9 2
47 10 9 1 10 9 13 10 9 16 13 9 2 7 13 1 10 11 11 11 2 11 2 2 10 9 12 4 13 0 9 1 9 7 0 9 2 16 0 9 3 0 1 9 1 3 3 2
1 11
4 11 11 11 9
18 3 14 13 15 10 13 11 4 13 10 9 1 9 11 8 13 0 2
31 15 4 3 13 14 13 10 5 12 10 3 3 3 8 4 13 0 16 15 4 13 10 9 1 15 3 3 16 8 0 2
1 9
4 13 15 13 3
1 11
31 15 13 1 10 13 9 2 7 15 4 13 14 13 10 9 1 11 2 16 16 15 4 13 9 7 9 7 0 0 9 2
10 3 6 13 15 15 13 14 7 13 1
12 3 15 13 2 7 15 4 13 0 3 3 2
3 11 11 11
3 9 2 8
52 6 2 0 9 9 13 3 3 0 2 15 4 13 14 13 10 0 9 16 15 13 10 9 15 4 13 14 13 3 7 15 13 1 1 9 3 15 13 10 0 9 3 2 7 15 4 13 10 9 3 6 2
1 13
14 11 15 1 12 13 3 0 14 13 16 15 13 9 2
31 15 4 3 13 10 9 7 13 10 3 0 9 2 7 15 13 10 9 7 3 15 13 3 0 15 13 14 13 10 9 2
19 0 9 1 15 7 4 13 16 15 14 13 10 9 14 13 9 2 0 5
9 9 2 2 11 11 2 2 8 2
3 9 2 9
31 15 4 13 14 13 15 14 13 1 10 9 3 15 4 13 13 9 10 4 14 3 13 2 7 3 13 1 0 0 9 2
22 15 13 10 0 9 1 10 9 9 9 7 10 9 9 2 9 1 10 9 9 9 2
1 8
3 9 2 8
3 11 9 12
22 15 13 10 9 1 11 2 13 1 10 1 15 16 15 13 9 2 15 13 3 0 2
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
1 8
8 6 2 15 13 3 1 11 2
1 13
9 9 2 2 11 11 2 2 8 2
3 9 2 9
34 15 13 10 9 10 13 14 13 0 1 12 1 15 9 1 1 9 2 15 13 10 0 1 12 9 0 0 2 0 9 2 3 0 2
12 15 13 1 9 2 9 9 2 9 2 8 2
17 13 0 9 1 11 7 13 9 2 13 9 1 9 2 3 0 2
8 9 2 2 11 2 2 8 2
3 9 2 9
11 16 15 13 2 10 9 13 15 1 2 2
4 3 3 3 2
8 13 16 15 9 4 13 1 2
12 3 15 4 14 13 14 13 3 15 13 14 2
15 15 4 14 13 10 9 1 10 9 1 2 10 2 9 2
13 9 13 1 10 9 15 13 2 15 13 14 9 2
10 3 10 9 13 10 2 0 2 9 2
1 11
25 15 4 13 1 9 15 4 13 14 13 11 7 11 12 7 13 1 7 1 10 11 2 11 9 2
19 15 13 12 9 3 3 2 7 15 13 0 14 13 2 16 9 13 0 2
15 10 9 4 13 14 13 9 1 11 2 11 2 7 11 2
19 6 13 15 13 16 15 13 0 2 7 16 15 13 10 9 2 6 13 2
13 13 15 3 3 7 15 13 14 13 1 15 3 2
9 9 2 11 11 11 11 2 8 2
24 10 0 0 9 11 11 4 13 14 13 10 11 9 2 1 9 16 3 15 9 4 4 13 2
5 1 0 9 2 8
1 2
7 10 9 4 3 13 0 2
21 15 4 13 10 11 11 11 11 16 15 13 1 15 7 2 9 13 15 1 15 2
17 14 13 2 7 13 16 10 9 4 13 1 15 2 13 1 2 8
3 2 8 2
23 16 15 4 13 9 1 9 16 10 11 9 13 10 9 1 11 2 10 9 4 4 13 2
20 9 9 7 3 11 9 11 11 13 3 1 10 9 1 10 12 2 9 9 2
17 15 13 16 10 9 1 9 9 4 3 3 13 1 10 9 9 2
16 3 0 3 16 11 14 9 4 14 13 1 10 0 12 9 2
1 2
11 13 1 11 11 1 11 11 1 12 12 9
5 6 0 9 9 2
9 10 0 0 9 4 13 15 9 2
17 3 2 11 7 11 13 0 7 10 9 4 4 3 13 1 11 2
35 1 11 0 9 1 10 9 9 1 0 11 1 10 0 9 1 9 11 7 11 2 0 11 7 11 13 3 1 10 0 9 1 0 11 2
20 15 4 13 1 10 0 9 9 1 11 13 12 9 7 13 0 1 12 9 2
49 1 0 0 9 1 10 9 9 1 0 11 1 11 7 11 10 0 11 7 11 13 3 1 10 9 9 1 11 10 4 13 1 9 1 0 9 1 10 9 13 9 1 0 9 2 9 2 8 2
3 11 11 11
10 9 2 2 10 11 11 2 2 8 2
3 9 2 9
9 2 8 8 8 8 8 8 13 2
23 2 9 12 2 12 7 12 1 12 0 9 1 9 7 9 4 13 1 10 11 11 9 2
4 13 10 9 2
6 3 0 1 12 9 2
1 8
29 16 15 13 0 1 2 10 11 11 2 15 4 13 15 16 15 4 13 0 1 12 9 1 0 9 1 10 9 2
8 0 1 15 13 1 0 9 2
7 15 4 3 13 10 9 2
23 10 9 1 10 9 13 16 10 9 4 13 3 15 0 9 7 13 15 13 1 10 9 2
16 10 9 15 4 3 13 9 16 13 10 0 9 1 9 9 2
14 7 16 15 13 15 10 9 2 15 4 13 0 3 2
7 6 13 15 13 9 2 5
1 8
1 9
1 11
8 9 2 2 11 2 2 8 2
18 6 2 6 2 15 13 14 13 9 9 2 9 3 9 1 9 9 2
6 15 13 0 1 15 2
13 0 9 15 13 13 9 14 9 15 13 3 0 2
11 15 4 14 13 13 15 0 7 14 3 2
10 3 3 15 13 3 16 15 13 9 2
30 15 13 0 14 13 1 9 1 9 2 16 15 13 16 15 13 14 9 3 3 1 9 13 9 14 9 13 14 0 5
7 3 15 13 9 7 9 2
10 15 9 13 15 0 9 7 13 15 2
14 3 2 15 13 9 7 13 14 13 9 14 9 5 2
1 8
8 9 2 2 11 2 2 8 2
34 15 9 0 16 9 13 1 9 2 3 15 13 3 1 9 10 0 9 15 13 13 13 1 10 0 0 9 7 9 2 13 10 9 2
7 9 2 11 11 2 8 2
3 9 14 9
18 0 9 7 9 13 1 10 9 10 13 10 9 1 9 1 10 9 2
15 15 13 0 14 13 0 9 1 15 16 15 13 3 3 2
5 0 9 9 1 9
34 10 1 10 9 3 13 0 9 9 16 15 13 1 1 10 1 10 9 1 10 0 9 13 1 10 9 7 9 15 13 1 10 9 2
18 0 9 4 13 1 0 9 1 10 9 14 13 0 9 1 15 9 2
3 0 0 9
18 10 9 1 11 7 11 13 9 1 0 9 1 10 9 1 10 9 2
16 1 10 9 2 15 13 0 9 9 1 15 9 1 0 9 2
25 16 15 4 13 1 10 0 9 1 10 9 2 15 4 13 0 0 9 2 10 4 3 13 15 2
5 0 9 1 2 8
30 0 9 3 15 13 10 0 9 7 9 9 9 10 2 1 10 0 9 9 2 13 1 9 2 9 2 7 9 9 2
39 15 3 13 10 9 1 10 0 9 1 9 14 13 15 1 10 0 9 7 2 3 2 14 13 15 0 1 8 9 15 13 9 1 10 9 7 10 9 2
11 10 9 15 13 15 4 13 10 9 9 2
35 15 13 12 9 2 10 1 10 4 13 1 12 9 10 7 10 9 1 10 13 12 9 13 10 9 16 13 10 9 9 7 9 9 9 2
14 15 13 1 9 1 9 9 7 13 15 4 13 15 2
14 10 9 2 1 1 10 9 9 2 13 0 1 2 2
11 15 13 10 9 1 10 9 4 3 13 2
23 10 9 4 13 15 3 3 16 9 13 0 9 7 10 13 10 0 9 0 9 1 11 2
23 3 15 13 0 14 13 10 9 7 2 16 15 13 10 9 2 13 10 9 1 15 9 2
15 13 15 10 9 3 3 15 13 10 0 9 16 15 13 2
29 15 4 14 13 15 15 13 2 7 1 10 3 0 9 15 4 13 10 0 7 3 0 9 14 13 7 13 9 2
39 15 13 3 0 2 15 3 4 13 0 9 16 3 13 1 9 1 9 2 3 10 9 4 13 15 10 9 7 10 9 7 15 4 14 13 15 0 9 2
24 9 9 13 3 10 0 9 9 2 3 15 13 10 0 9 1 10 9 4 13 10 0 9 2
16 0 9 1 9 15 4 13 1 15 9 7 15 9 13 0 2
13 5 13 1 8 2 0 2 0 2 0 9 9 5
9 10 9 12 9 9 1 10 9 2
3 5 12 9
15 5 12 0 2 0 2 9 0 9 2 0 9 1 9 5
13 5 13 1 8 2 0 2 0 2 0 9 9 5
9 10 9 12 9 9 1 10 9 2
3 5 12 9
15 5 12 0 2 0 2 9 0 9 2 0 9 1 9 5
2 6 2
6 15 9 13 11 11 2
14 15 13 10 0 9 13 1 9 2 1 12 9 9 2
47 15 13 10 9 1 12 9 2 13 10 12 12 9 11 11 2 7 9 1 9 9 2 7 13 1 12 9 1 11 11 2 1 10 9 7 1 9 2 1 2 0 1 11 7 11 11 2
44 3 2 15 4 13 10 9 1 0 9 14 13 9 9 2 1 11 11 2 9 2 10 9 1 9 1 11 11 2 15 4 13 1 9 1 11 2 11 11 2 1 11 12 2
64 15 4 13 9 2 0 9 2 0 9 2 1 9 15 3 13 10 0 9 14 13 15 9 9 2 10 0 9 1 9 13 9 2 9 2 0 7 9 9 9 2 9 2 9 2 9 2 9 2 9 2 12 2 9 2 9 7 9 2 9 2 7 9 2
30 16 15 4 3 13 10 1 10 9 14 13 9 9 2 6 13 15 1 8 7 13 15 13 2 13 15 1 15 9 2
8 13 15 1 15 9 7 9 2
3 0 9 2
2 11 11
35 3 1 10 9 2 1 12 2 14 13 0 2 2 10 11 2 11 9 13 10 9 9 1 10 0 7 0 0 9 1 10 9 1 11 2
25 1 9 16 13 0 9 1 9 1 1 10 0 9 2 10 0 9 13 14 13 10 9 0 9 2
26 7 1 10 0 0 9 2 10 9 9 13 14 13 15 9 4 13 0 2 3 15 13 1 10 9 2
36 11 2 11 13 10 9 1 10 9 7 13 14 13 1 15 9 16 13 15 0 9 1 0 9 2 13 15 4 13 0 9 1 15 0 9 2
45 1 0 9 1 9 2 15 13 1 10 0 9 3 10 9 9 4 3 13 10 9 13 3 10 9 9 14 9 9 7 13 0 1 9 2 10 3 0 2 9 2 13 0 9 2
25 10 9 9 7 9 4 3 3 3 13 14 3 13 0 9 2 3 10 9 4 13 1 0 9 2
13 9 1 10 9 2 4 14 13 11 2 13 11 2
22 3 13 2 11 13 3 1 10 9 16 4 13 1 1 11 1 0 9 2 3 3 2
29 10 11 11 11 11 11 11 11 2 11 2 13 10 9 9 9 1 10 11 11 1 11 11 2 11 2 0 9 2
65 10 9 2 13 1 10 11 11 11 1 11 7 11 11 2 13 11 16 13 10 12 9 9 13 1 1 0 11 11 11 11 9 2 10 11 1 11 11 2 11 2 7 10 11 11 1 11 7 11 11 1 10 11 11 9 1 11 11 2 3 13 1 11 11 2
31 10 0 9 13 16 11 4 14 13 0 0 11 11 9 10 9 1 9 1 0 0 9 9 1 11 11 1 10 12 9 2
37 1 9 1 11 11 1 10 11 11 9 2 0 9 4 4 13 16 15 13 10 0 0 9 9 1 11 11 16 10 9 4 4 13 1 11 9 2
29 3 2 0 9 9 4 13 0 14 13 10 9 1 10 15 13 0 1 10 9 7 4 13 0 2 1 10 9 2
19 2 1 10 9 1 11 11 2 0 9 1 11 11 13 3 0 1 3 2
22 1 0 2 15 13 0 16 11 13 1 12 9 9 2 2 13 11 11 2 11 11 11
28 0 2 9 9 13 11 16 13 11 11 2 3 10 9 12 9 2 13 14 13 9 9 1 10 11 1 11 2
24 11 11 14 0 9 2 0 0 9 1 9 1 11 13 12 9 14 13 1 12 9 1 9 2
20 1 11 2 10 9 1 11 11 11 9 1 11 9 13 12 9 1 12 9 2
27 16 13 10 11 11 9 1 11 2 11 13 9 1 3 12 9 10 9 16 15 13 1 10 11 1 11 2
29 10 11 11 11 11 13 11 13 2 3 0 2 7 4 13 10 0 2 9 9 12 9 1 10 11 2 11 9 2
22 10 9 13 9 9 1 10 11 1 11 3 3 12 2 9 1 11 9 9 4 13 2
16 9 9 13 0 9 16 10 9 14 9 13 0 9 1 9 2
19 1 11 2 11 13 15 12 9 1 9 9 7 11 13 15 12 9 9 2
20 11 13 15 4 13 9 1 15 12 9 11 11 9 7 15 12 9 11 9 2
11 11 11 13 0 9 1 12 0 11 9 2
23 0 9 2 11 13 9 1 11 7 11 7 13 9 1 10 0 9 1 12 9 10 9 2
16 6 13 10 9 3 10 13 0 2 9 1 15 9 7 9 2
3 2 8 2
5 2 11 11 11 2
23 11 4 13 1 0 9 14 13 7 9 7 9 1 10 11 11 11 2 15 13 10 9 2
3 2 2 2
45 2 15 13 14 9 2 0 13 9 9 16 1 10 0 9 13 16 13 3 1 10 11 2 2 13 11 11 2 9 1 11 11 2 12 1 10 9 13 14 13 9 1 10 11 2
21 11 13 16 13 10 9 9 1 12 2 10 3 13 15 1 12 9 1 10 11 2
21 13 10 9 4 13 10 0 9 2 13 10 9 1 10 0 9 13 10 9 9 2
32 16 10 4 13 15 1 10 9 16 10 0 9 14 3 13 10 0 9 2 11 13 0 16 13 1 10 9 1 10 0 9 2
5 2 11 11 11 2
35 1 12 11 2 11 9 11 11 13 10 11 11 11 11 16 10 9 13 14 13 3 5 12 12 1 10 0 9 7 9 9 1 12 9 2
24 2 10 9 1 10 0 9 2 2 2 4 13 0 14 13 0 9 14 13 2 2 11 13 2
32 2 15 13 16 9 2 16 13 1 10 9 2 4 13 3 2 1 10 9 2 2 7 15 4 14 13 15 2 2 11 13 2
14 3 9 4 13 16 11 14 9 4 7 13 7 13 2
46 7 13 3 10 0 9 4 13 0 14 3 13 9 1 10 11 2 1 3 10 9 1 10 9 2 2 15 4 13 1 10 9 16 0 11 13 0 14 8 13 15 0 9 1 9 2
1 2
11 13 1 11 11 1 11 11 1 12 12 9
3 2 8 2
48 3 10 9 13 0 2 10 9 13 2 7 1 10 8 2 13 9 9 2 0 9 11 11 4 13 16 11 13 10 10 9 10 15 13 1 10 12 9 2 10 13 11 11 1 10 9 2 2
7 12 9 13 0 1 0 2
40 16 11 13 1 10 2 9 9 2 15 4 13 0 9 9 7 4 3 3 13 11 2 10 4 3 13 10 0 9 16 13 1 10 11 2 13 10 11 11 2
5 11 9 2 11 11
40 0 0 9 7 10 9 2 9 1 10 0 11 12 2 12 0 9 11 11 13 1 15 0 0 9 9 1 10 11 11 9 1 11 2 11 11 12 2 12 2
17 13 15 1 11 11 14 9 2 11 13 14 13 0 9 1 9 2
18 15 13 16 10 0 9 2 0 2 4 14 13 10 9 9 1 11 2
20 15 4 3 13 9 16 11 13 6 1 3 3 10 9 2 7 1 11 15 2
35 13 15 9 2 11 13 9 1 10 13 11 9 16 15 13 0 14 13 9 1 15 9 7 13 10 9 1 11 14 3 13 11 11 9 2
16 11 3 13 14 13 10 9 1 9 1 0 9 7 15 9 2
28 11 2 10 9 15 16 15 13 9 10 0 0 9 1 11 2 13 10 9 9 2 3 0 7 3 0 2 2
25 4 3 13 10 11 11 7 11 2 15 4 13 16 10 0 0 9 4 13 14 13 10 9 9 2
33 16 11 4 14 13 15 0 9 7 13 10 9 1 11 11 2 3 15 4 14 13 9 1 10 11 11 7 10 11 4 3 13 2
2 11 2
1 2
11 13 1 11 11 1 11 11 1 12 12 9
3 2 8 2
8 2 9 9 2 11 14 11 2
3 2 11 2
25 10 0 0 9 11 4 13 10 9 1 9 9 1 11 1 10 11 11 1 10 9 1 13 9 2
19 1 1 12 9 4 4 13 1 11 2 9 16 15 9 13 1 10 9 2
18 1 9 1 10 9 2 11 13 15 9 16 13 0 9 1 9 9 2
19 13 1 11 11 14 13 2 0 2 9 2 15 0 13 0 9 9 3 2
30 15 13 16 16 11 4 13 3 10 9 1 10 9 2 0 14 13 10 9 10 11 11 11 4 13 1 10 9 9 2
21 11 11 2 11 14 9 13 10 9 9 16 11 13 15 0 9 2 11 11 11 2
26 11 4 13 3 0 1 11 2 16 0 13 10 0 9 9 1 10 9 1 10 9 9 1 0 9 2
26 11 13 10 9 14 13 16 15 13 11 14 13 10 9 2 16 10 0 4 14 4 13 1 11 11 2
4 2 11 11 2
34 2 15 13 14 0 1 11 14 9 1 10 9 7 1 9 1 10 0 9 1 10 11 2 2 13 11 11 2 10 0 11 11 9 2
13 2 7 15 13 16 11 13 15 0 0 9 2 2
3 2 2 2
26 2 10 9 13 14 1 10 0 9 9 7 1 11 14 9 14 13 10 11 14 9 2 2 11 13 2
25 2 11 13 13 1 11 2 16 1 10 9 2 7 10 0 9 4 14 13 9 14 13 15 9 2
11 11 13 14 13 10 11 1 0 9 2 2
24 11 11 4 13 14 13 10 9 9 2 7 13 14 13 10 11 11 2 1 10 0 9 2 2
50 16 11 11 11 13 3 2 11 4 3 13 1 10 9 9 1 10 9 11 13 0 13 11 1 15 0 9 2 16 3 10 0 9 11 4 13 13 13 1 7 13 14 13 9 1 15 9 14 13 2
1 2
11 13 1 11 11 1 11 11 1 12 12 9
9 11 13 10 0 7 10 0 9 2
6 11 13 14 10 9 2
5 11 13 1 11 5
10 3 0 13 10 11 11 1 15 9 2
7 5 12 1 10 11 11 2
1 5
2 5 5
8 10 9 4 15 13 1 11 2
7 0 9 3 3 2 6 2
2 6 2
1 9
9 15 13 11 11 15 13 0 9 3
9 4 15 13 10 9 1 9 9 2
19 2 6 7 15 13 0 1 15 2 16 15 9 4 14 13 15 15 3 2
9 4 15 13 10 9 1 11 11 2
5 15 4 4 13 3
2 6 2
9 15 13 0 3 1 15 0 9 2
5 13 15 15 9 2
12 4 9 14 9 1 11 3 13 3 12 9 2
13 16 15 4 4 13 1 11 3 7 15 13 0 2
1 8
5 13 9 9 9 2
9 15 13 11 14 9 9 1 9 2
21 15 4 13 15 2 15 4 14 13 15 3 3 15 13 15 9 13 3 15 13 9
1 8
7 15 4 15 13 1 11 2
22 9 1 10 9 15 13 1 0 9 1 9 2 9 2 9 2 9 2 9 2 8 2
7 13 13 15 1 0 9 5
9 9 13 1 10 11 9 1 11 2
28 15 4 13 10 11 9 1 10 9 1 11 7 15 13 14 13 1 11 9 13 3 15 4 4 13 1 11 2
7 10 9 1 11 11 9 2
2 10 2
9 15 13 15 13 10 11 11 9 2
15 15 13 15 0 9 10 15 4 3 13 13 10 9 9 2
1 8
17 3 14 13 10 9 9 9 1 0 9 1 9 12 9 1 9 2
13 3 13 10 9 9 1 10 9 10 13 9 9 9
1 8
7 15 13 10 9 9 14 13
14 3 0 9 4 9 9 13 14 13 1 11 1 11 2
9 13 15 12 9 13 11 7 9 2
16 12 1 12 9 16 15 13 0 1 0 15 13 3 12 9 2
3 6 12 9
11 15 13 10 0 11 11 1 11 2 11 2
10 10 11 11 2 11 2 13 10 0 2
8 10 11 11 11 13 3 0 2
12 15 13 14 10 0 9 2 7 13 3 0 2
1 8
2 9 2
5 3 4 11 13 2
14 15 4 13 0 9 1 10 0 9 15 13 15 0 2
5 11 12 2 12 2
12 15 4 13 1 10 9 1 11 12 2 12 2
7 11 4 13 11 12 12 2
9 4 9 0 2 9 13 1 11 2
17 0 9 1 10 9 9 13 1 10 9 2 7 3 6 14 3 2
4 6 2 6 2
10 10 9 1 10 9 9 0 9 13 2
8 3 1 15 15 4 14 13 2
12 15 13 10 0 12 5 9 1 10 11 11 2
6 1 9 11 11 9 2
11 3 1 11 11 2 11 11 2 11 11 2
9 15 13 14 13 3 1 15 9 5
11 3 15 13 12 15 4 13 8 3 15 13
16 15 13 9 1 9 9 13 3 2 15 4 15 13 1 15 2
6 15 13 1 3 0 9
17 15 13 15 1 10 9 9 1 0 9 7 10 0 9 14 9 2
4 13 1 9 2
9 13 15 1 10 0 7 13 15 2
9 13 11 10 0 9 1 10 9 2
7 15 4 13 15 11 1 0
17 15 13 10 9 13 11 2 3 6 2 11 13 14 10 0 9 2
11 15 13 15 9 15 4 13 10 9 15 13
3 6 6 2
6 15 13 10 0 9 2
2 9 2
8 15 14 13 1 11 11 11 2
27 6 3 15 13 1 11 11 11 6 1 10 11 11 7 10 11 11 2 15 13 0 9 14 13 3 3 2
4 6 10 9 2
4 15 13 12 3
5 15 1 9 2 2
6 6 9 9 7 9 2
19 10 1 15 4 15 13 2 11 14 2 11 11 2 11 11 2 11 14 2
2 11 11
19 15 13 16 15 13 1 10 0 9 1 11 14 2 15 9 13 3 3 0
6 11 14 10 0 1 15
11 10 12 15 13 10 3 4 13 11 14 2
12 4 9 13 15 10 9 1 0 9 1 11 2
22 3 15 13 10 9 1 15 3 6 13 15 3 3 16 15 13 9 1 0 9 1 11
23 15 4 14 13 1 9 1 10 9 1 10 9 7 15 4 3 13 9 1 10 9 2 8
13 15 13 10 9 9 1 9 1 11 11 14 11 2
18 15 9 14 9 13 11 9 7 15 4 13 1 11 11 14 1 9 2
23 15 13 0 16 15 15 4 13 2 15 13 9 9 7 15 4 4 13 1 0 0 9 2
3 6 13 2
3 12 2 9
6 9 1 10 11 9 2
19 4 9 13 1 10 11 9 1 15 0 1 11 7 3 3 4 10 11 13
4 10 0 9 2
24 9 13 12 5 12 4 4 13 14 13 3 1 11 14 9 2 15 4 13 15 1 10 9 2
8 11 13 1 11 11 11 9 2
13 15 13 10 9 9 1 9 1 11 11 14 11 2
26 15 4 4 13 1 11 11 14 1 0 11 1 9 7 15 4 13 15 10 9 9 13 1 10 9 2
15 15 13 9 9 7 15 13 15 4 4 13 1 0 9 2
3 6 13 2
3 12 2 9
5 15 4 13 1 8
21 4 15 13 10 9 10 13 10 10 9 9 10 4 3 13 16 10 11 13 15 2
6 13 11 13 9 9 2
39 1 1 10 12 12 13 13 9 1 9 1 10 11 2 12 12 3 13 0 2 7 15 13 9 1 9 10 4 14 4 13 1 15 8 0 9 7 9 2
2 11 2
8 4 15 3 13 10 9 1 2
7 6 15 13 11 15 13 11
1 11
1 11
8 13 15 13 10 0 9 1 2
15 11 13 1 0 2 7 15 13 10 9 10 13 15 13 2
14 15 13 3 3 0 9 1 10 11 1 9 1 11 2
11 15 13 11 13 10 0 9 9 7 9 2
3 15 13 9
10 9 13 10 0 9 1 10 9 9 2
13 3 1 9 9 7 0 9 1 10 9 1 11 2
2 6 2
6 3 15 13 3 3 2
4 12 9 1 9
4 12 9 1 9
5 12 9 1 0 9
8 12 9 1 1 10 9 1 11
4 13 15 10 1
4 3 13 1 15
2 10 9
14 15 13 3 16 13 9 2 3 13 10 9 1 1 15
23 15 13 10 9 1 11 11 11 7 15 13 10 9 1 1 0 7 13 15 4 15 13 2
21 15 4 13 10 9 1 10 9 7 13 15 1 14 13 15 13 15 4 15 13 2
4 13 10 0 9
10 13 15 4 14 13 10 9 7 13 15
18 15 13 0 14 13 13 9 2 3 16 15 4 14 13 15 4 13 2
13 6 6 3 4 15 13 11 11 3 1 11 6 2
4 15 4 14 2
8 15 4 14 13 15 1 11 11
32 15 4 14 7 3 13 10 9 2 10 9 13 0 14 13 10 9 1 15 9 7 11 2 15 4 13 15 0 0 9 2 2
6 11 13 3 1 11 2
4 11 13 0 2
9 13 15 4 14 13 15 3 3 2
22 15 13 1 9 1 9 7 15 13 14 13 1 9 3 15 0 4 15 13 14 13 2
8 9 2 3 9 7 3 9 2
8 15 13 10 9 1 9 9 2
9 15 13 14 0 14 13 9 9 2
11 13 1 15 0 9 2 13 15 15 13 2
14 3 14 2 0 2 9 2 0 9 13 1 10 9 2
1 8
8 13 10 11 10 0 0 9 2
21 15 4 13 10 9 1 9 7 15 13 14 13 16 10 11 13 10 0 0 9 2
3 13 15 2
17 3 2 11 13 16 15 13 10 0 1 0 9 7 9 7 9 2
13 7 9 13 10 0 2 0 2 0 9 0 9 2
6 6 2 15 13 14 2
13 7 15 4 13 10 9 15 13 1 1 10 9 2
6 11 11 7 11 11 2
6 10 12 4 15 13 2
11 15 13 3 3 10 0 9 2 6 13 2
5 13 1 10 11 2
26 15 13 3 0 2 9 12 9 2 11 3 12 2 2 0 9 1 9 7 10 11 3 9 2 12 2
15 10 13 0 12 9 1 0 9 2 3 15 4 14 13 2
14 10 11 13 10 3 0 9 7 10 0 9 12 9 2
7 9 13 1 0 9 9 2
14 15 4 13 1 10 0 9 9 1 15 9 1 11 2
9 4 13 1 10 9 1 0 9 2
6 4 15 13 10 9 2
19 16 15 13 0 16 7 3 15 13 15 9 3 11 4 13 0 14 13 2
4 6 2 3 2
5 3 1 10 9 2
6 13 3 15 4 13 2
15 16 15 13 1 10 11 7 13 1 11 3 15 13 10 9
8 3 4 15 13 9 1 11 2
15 4 10 9 6 13 15 3 15 4 13 10 9 1 11 2
9 13 15 10 9 7 9 6 13 2
6 13 3 0 3 6 2
1 9
6 15 4 3 13 15 2
9 9 15 13 1 10 9 7 0 2
14 3 4 9 13 10 9 1 10 9 1 10 0 9 2
5 15 13 10 9 2
13 13 1 15 9 2 15 4 13 15 10 3 3 2
7 15 4 10 0 9 13 2
12 15 13 10 9 7 15 4 13 1 15 3 2
34 15 4 4 13 3 7 15 13 14 10 0 9 15 13 13 8 8 8 2 7 9 1 15 2 4 9 13 10 9 15 4 13 1 2
10 16 10 9 13 15 13 0 14 13 2
13 13 13 15 7 13 15 1 11 15 4 13 0 2
2 9 2
9 16 15 13 10 9 3 15 13 0
9 9 13 10 9 1 9 1 11 2
28 15 13 15 12 9 9 1 10 0 9 7 4 13 16 9 4 13 15 1 10 0 9 1 11 7 0 0 9
38 15 13 11 11 11 2 10 9 2 15 13 3 1 11 11 2 3 15 4 13 10 0 9 1 10 11 11 2 11 11 2 11 11 2 10 3 0 2
3 11 11 14
6 15 13 3 3 0 3
16 15 4 13 16 15 13 10 9 1 11 11 1 0 9 11 2
20 15 4 13 0 16 13 10 9 1 10 11 11 1 0 9 11 7 1 11 2
7 15 4 4 13 10 9 2
22 10 9 4 13 15 13 15 3 7 15 4 13 9 7 9 2 7 3 3 9 2 2
11 15 4 3 13 10 9 1 0 9 3 2
6 15 4 4 13 7 13
9 6 2 15 4 13 10 9 9 2
4 11 9 9 2
5 3 4 15 13 2
6 16 9 0 4 13 2
5 3 4 15 13 2
7 3 16 15 13 14 13 2
14 7 16 9 0 4 13 2 15 4 15 9 13 1 2
5 15 13 1 11 2
8 15 13 1 10 11 11 9 2
22 10 0 12 4 13 2 9 1 9 2 1 10 0 9 1 10 13 1 11 1 2 8
10 15 4 13 12 16 10 11 11 13 2
6 11 13 3 0 7 0
5 11 11 9 9 2
28 0 9 2 15 13 10 9 13 1 11 2 0 9 2 12 9 1 9 2 15 4 13 16 11 11 13 9 2
1 9
43 15 4 13 13 15 10 9 3 2 15 13 15 4 14 13 15 10 9 1 10 9 2 7 13 15 13 2 13 13 15 14 13 1 10 9 2 7 15 13 9 0 1 15
15 13 2 7 13 2 10 0 9 3 7 13 10 9 3 2
10 10 9 1 9 4 9 1 11 13 2
23 15 4 13 10 9 7 13 14 13 10 9 9 11 9 13 1 9 2 9 2 7 9 2
12 7 15 13 15 0 2 0 9 1 10 9 2
9 6 1 11 9 13 15 0 9 2
11 7 1 10 9 15 13 10 1 15 9 2
14 0 9 2 15 13 2 9 2 9 2 9 2 9 2
6 3 14 13 15 1 2
14 15 13 9 1 13 9 2 9 2 7 0 2 1 9
13 3 4 15 13 14 13 9 9 1 10 9 9 2
2 9 6
16 3 4 9 13 14 13 3 15 13 14 13 10 9 1 9 2
32 3 13 10 9 1 9 3 15 13 10 9 7 13 10 0 9 1 9 9 14 13 15 9 13 14 13 16 13 1 10 9 2
6 13 15 13 1 3 5
8 15 4 13 15 1 16 13 2
24 3 15 13 16 15 13 14 13 1 9 7 15 3 4 14 13 0 16 15 4 14 13 10 9
9 0 9 0 1 11 11 1 11 2
17 1 10 9 9 1 15 9 2 15 4 13 1 10 11 11 11 2
11 1 15 2 15 4 13 0 14 13 9 2
28 13 10 0 9 2 15 4 14 3 13 3 13 0 2 0 2 7 0 1 9 9 2 12 11 11 11 2 2
17 4 9 13 10 9 1 9 1 9 9 3 15 4 14 13 0 2
5 15 4 14 13 2
16 3 16 15 13 10 9 3 2 9 4 13 15 10 0 9 2
9 4 11 11 13 9 16 13 9 2
29 15 13 0 14 13 10 9 1 11 11 2 7 15 4 14 13 13 10 9 16 15 13 12 0 9 1 15 9 2
11 16 15 13 7 13 3 4 15 13 15 2
10 3 4 14 15 13 10 9 7 13 2
47 15 4 14 13 15 13 16 10 9 13 14 0 7 15 4 13 15 3 0 1 10 9 1 10 9 7 16 15 13 10 9 15 9 15 4 3 13 16 3 15 13 10 9 2 9 1 15
7 9 1 11 2 13 6 2
36 15 13 14 13 10 0 9 13 1 15 9 2 1 11 2 1 10 10 9 1 11 4 15 13 9 7 9 16 13 9 2 6 13 2 13 15
24 9 9 13 10 0 9 3 9 9 1 11 7 10 11 1 11 5 10 9 1 11 11 1 11
14 9 1 11 13 10 0 9 1 15 2 10 10 0 2
13 13 11 2 15 13 8 0 7 13 1 10 9 2
13 9 13 0 0 3 16 10 9 4 13 1 11 2
24 15 13 10 0 7 0 9 2 7 15 13 12 9 1 10 9 1 10 9 2 4 15 13 2
15 3 3 14 2 16 15 13 14 10 9 13 1 10 9 2
6 15 13 0 14 13 2
8 9 4 13 0 9 3 3 2
18 3 16 15 13 10 9 7 9 2 15 4 14 4 13 10 12 13 2
17 15 4 13 13 3 10 9 7 13 15 3 1 10 3 0 9 2
23 16 15 13 10 0 9 1 10 9 2 10 13 15 13 0 7 4 13 16 13 1 3 2
3 13 9 2
7 3 4 10 9 13 11 2
32 15 13 14 0 1 10 9 1 10 9 7 15 13 10 9 1 0 9 1 0 7 0 9 1 11 3 15 13 3 10 9 2
30 15 13 9 1 9 13 11 2 15 4 13 10 9 16 15 13 10 9 7 10 9 1 9 15 4 13 1 15 1 2
5 3 13 12 9 2
12 15 13 10 11 1 11 2 3 3 1 11 2
18 15 13 3 10 11 1 11 2 10 9 1 10 3 0 11 11 11 2
10 11 11 13 10 9 3 1 11 11 2
3 9 9 2
62 6 6 15 13 10 9 1 12 9 7 3 15 13 3 11 14 9 7 15 3 13 1 1 15 7 15 4 13 12 1 10 9 15 13 7 12 9 13 1 15 9 9 15 13 15 9 15 13 10 9 7 15 13 10 9 14 9 15 4 15 13 2
5 7 15 13 12 9
13 6 15 4 3 13 3 3 7 13 15 3 15 13
7 15 4 13 1 10 0 9
9 7 1 10 9 15 4 13 10 0
6 3 13 0 9 13 2
5 15 13 3 13 2
5 4 14 13 13 9
2 0 9
7 13 11 11 11 3 0 2
5 13 15 3 0 2
13 16 15 4 13 16 15 13 9 15 13 14 0 2
14 16 15 13 14 0 13 15 0 9 14 13 15 9 2
8 15 4 13 1 11 1 10 9
1 6
2 6 2
12 6 9 1 15 9 13 3 0 1 11 11 2
38 13 9 2 16 15 13 0 9 2 15 4 3 13 1 9 2 15 4 3 13 10 3 15 4 13 0 14 13 1 9 9 2 7 15 13 0 3 2
19 9 2 12 9 2 12 9 7 12 9 2 8 2 1 10 12 9 9 2
13 15 13 14 13 9 1 11 11 15 13 1 11 2
24 15 13 1 11 13 1 11 11 11 12 9 15 13 14 13 0 9 3 3 15 4 13 15 2
7 15 13 0 9 1 9 2
10 15 4 13 1 15 16 15 13 0 2
10 15 4 13 0 9 3 1 10 9 2
35 3 3 16 15 13 10 9 7 13 15 1 9 15 4 14 13 10 9 13 1 15 7 15 9 4 13 9 14 13 16 3 15 13 15 2
29 13 1 11 1 6 12 13 10 9 9 3 13 15 9 13 1 7 13 5 12 1 9 13 10 9 3 1 9 3
9 13 1 11 7 15 4 14 13 2
20 1 15 0 9 1 11 2 15 4 4 13 1 11 16 13 3 1 10 11 2
8 15 4 13 1 11 1 12 9
22 8 2 10 9 1 11 13 10 0 9 10 13 14 3 3 1 10 0 9 1 11 2
14 10 9 15 4 13 3 1 9 3 16 13 10 9 9
27 8 2 15 4 13 14 13 1 10 9 1 10 8 2 3 0 9 2 16 0 2 2 7 10 9 9 9
17 8 2 3 13 10 9 3 15 4 13 0 9 2 9 13 10 9
7 15 13 14 13 15 0 9
12 16 15 4 14 13 15 4 13 10 0 9 2
24 3 4 15 13 9 1 11 11 2 15 4 13 10 0 9 2 7 15 4 14 13 9 6 2
33 15 13 3 1 10 9 2 7 15 4 14 13 12 9 1 11 11 10 13 9 2 3 13 1 9 9 2 0 9 7 9 9 2
16 15 13 16 9 13 3 0 14 13 3 1 10 11 11 9 2
21 7 15 4 13 10 9 2 8 2 3 15 13 10 9 1 9 2 13 9 9 2
13 3 13 10 9 1 10 9 7 13 10 9 9 2
2 6 2
2 6 2
28 15 4 14 13 2 7 15 13 16 15 4 14 13 15 2 4 15 13 16 2 9 13 0 9 1 9 2 6
14 13 15 10 9 1 0 9 0 1 11 7 11 11 2
23 11 11 9 13 3 1 11 2 12 13 1 11 7 11 1 11 11 2 13 1 11 11 2
19 3 1 15 15 13 0 9 10 13 9 1 11 2 12 9 7 11 11 2
6 6 9 9 13 0 2
5 15 13 14 0 2
2 6 2
17 6 9 2 15 4 13 9 1 0 9 9 1 11 1 11 11 2
5 15 13 11 11 2
22 9 2 11 11 2 11 11 11 2 0 0 9 9 3 3 13 1 11 7 11 11 2
21 15 4 13 15 1 11 11 11 2 11 2 12 2 11 11 11 2 11 11 2 8
2 9 2
16 3 4 15 13 9 3 12 2 12 1 15 11 11 12 9 2
32 15 13 9 1 15 9 2 7 15 13 3 1 15 9 2 13 15 10 9 15 4 13 10 9 14 13 10 11 15 13 9 2
56 15 13 14 13 0 14 13 15 1 15 9 2 3 7 3 8 2 15 13 1 10 9 2 7 15 13 3 3 7 2 15 13 15 15 13 3 10 9 16 3 13 3 14 13 12 15 4 13 1 3 3 3 1 10 11 2
42 15 13 14 13 10 11 1 9 2 3 9 2 3 15 13 10 9 10 15 13 1 3 10 13 9 1 9 7 15 4 13 1 15 3 7 15 13 14 13 15 1 15
7 3 13 11 7 11 0 2
3 7 0 2
15 15 4 13 10 9 16 3 11 7 11 13 0 7 0 2
17 15 4 13 1 10 9 1 12 9 7 3 3 15 4 13 9 2
13 15 13 14 13 3 15 13 0 7 0 1 10 9
7 9 7 10 9 1 10 9
5 9 16 13 1 9
4 0 9 1 9
5 15 13 10 9 2
9 9 1 10 11 1 9 7 9 2
6 0 9 1 10 9 2
9 9 1 10 9 1 10 0 9 2
11 4 9 6 13 15 15 13 0 11 2 5
17 0 2 12 13 1 10 9 2 10 0 13 1 10 0 9 9 2
23 0 2 10 4 13 1 9 9 1 10 11 2 3 3 15 10 0 9 9 13 15 2 2
16 15 13 15 9 14 9 7 3 4 15 13 15 2 15 15 2
8 16 15 13 10 9 3 3 2
7 15 9 14 9 13 11 2
15 3 15 13 10 0 0 9 15 13 1 10 9 9 9 2
16 15 13 10 0 9 7 15 4 13 15 1 1 12 9 3 2
21 15 4 10 0 9 13 11 15 13 15 15 16 15 13 10 9 9 1 15 9 2
9 7 15 13 10 9 1 10 9 2
5 15 13 15 2 5
24 15 13 10 0 9 9 10 4 13 11 16 1 10 9 15 3 13 15 9 3 15 13 3 2
17 15 9 4 13 11 16 10 9 15 13 15 13 10 9 11 11 13
11 15 3 13 0 0 9 16 11 11 13 5
12 15 4 15 13 3 10 0 9 9 13 0 2
28 15 0 9 3 13 9 9 7 9 10 1 10 9 13 0 3 15 13 0 15 13 6 14 1 0 9 9 2
5 15 13 3 0 2
10 16 15 13 10 9 15 13 3 0 2
20 16 15 13 10 9 9 7 13 15 1 10 9 7 15 13 9 13 15 1 2
10 16 15 13 14 15 4 13 14 13 2
17 16 15 13 10 9 14 13 10 9 2 10 9 4 3 13 0 2
32 16 15 4 13 10 9 7 15 13 14 1 10 0 9 7 13 7 15 13 15 3 15 15 4 13 15 9 7 3 13 9 2
12 13 15 13 13 9 16 15 4 13 3 0 2
4 16 15 13 2
3 13 15 13
20 15 13 12 9 1 11 11 2 15 13 10 0 9 14 13 1 15 0 9 2
22 15 13 10 9 9 2 9 1 11 11 7 15 9 13 14 13 10 1 10 0 9 2
14 15 4 13 3 1 10 9 10 4 13 3 1 11 2
21 15 13 0 9 15 13 10 0 9 14 13 2 13 16 15 3 13 10 0 9 2
13 2 15 13 1 0 9 7 15 13 0 9 2 2
10 13 1 10 13 3 8 13 3 9 2
33 15 4 13 15 1 10 10 0 9 2 11 11 2 11 2 11 2 8 2 7 15 4 13 3 3 15 13 14 13 0 9 1 2
14 13 1 8 7 13 9 1 3 10 9 1 10 9 2
2 11 9
5 13 10 9 9 2
6 15 13 10 0 9 2
14 13 15 0 14 13 10 9 3 7 1 10 9 9 2
13 0 9 14 13 1 10 9 10 7 10 9 4 13
30 3 2 15 4 14 13 10 9 9 14 13 1 9 1 15 16 15 13 0 14 13 1 10 9 13 9 1 10 9 2
10 15 4 14 13 0 9 1 9 9 2
22 15 4 14 13 14 13 9 1 10 9 15 4 13 7 10 9 15 13 0 1 15 2
23 10 12 9 15 3 13 1 10 9 9 15 4 14 13 10 1 10 9 15 4 13 1 2
32 10 0 9 15 4 13 1 10 9 9 15 13 0 14 13 10 0 1 0 1 15 0 2 7 0 9 16 15 15 4 13 2
11 3 3 15 4 14 13 1 15 3 3 2
7 0 13 13 10 0 9 9
8 15 11 13 2 13 9 3 2
16 6 2 15 13 10 9 7 15 9 13 3 3 0 1 9 2
15 6 0 9 16 15 4 13 2 15 9 13 1 15 9 2
23 15 13 1 15 9 2 7 15 13 3 0 9 1 3 2 15 4 14 13 15 14 13 2
8 15 13 9 1 9 1 3 2
10 9 13 15 9 1 10 9 7 9 2
9 13 15 16 15 13 10 9 9 2
31 15 4 14 13 2 15 3 13 10 9 1 15 9 12 9 3 15 13 3 1 10 9 7 15 13 3 0 1 10 9 2
10 15 4 4 13 9 9 10 0 9 2
11 15 13 0 7 13 10 9 1 1 15 2
15 13 0 15 13 14 0 3 7 13 10 9 1 9 1 2
5 15 4 13 7 13
6 13 13 7 13 13 2
9 4 15 13 10 0 9 9 6 2
15 15 13 10 0 0 9 10 15 9 4 13 15 13 6 13
17 15 13 9 0 0 14 13 9 1 7 9 14 3 13 1 15 9
10 10 9 13 3 0 14 13 9 1 2
13 15 10 13 9 7 9 2 9 2 0 9 8 2
26 10 0 9 4 13 10 9 2 7 15 13 14 13 10 9 3 2 13 15 10 0 9 2 8 8 8
7 13 10 9 13 14 0 2
8 15 4 13 10 9 1 9 2
15 15 13 10 9 1 9 7 15 13 0 7 13 9 1 2
13 16 15 13 0 3 13 1 10 9 9 7 9 2
27 15 4 13 1 10 0 9 0 1 10 9 2 9 2 9 7 9 16 15 13 9 15 4 13 7 13 2
11 9 13 3 10 0 14 13 9 1 3 2
4 0 9 9 2
16 15 4 4 13 10 9 1 11 11 1 10 9 1 9 3 2
24 15 4 13 3 1 10 9 7 15 4 13 16 13 1 15 1 15 9 13 3 15 9 9 2
23 15 13 3 10 3 0 9 7 15 4 14 13 9 3 3 15 13 3 3 10 0 9 2
15 15 3 4 14 13 14 13 15 1 7 13 15 13 0 2
15 13 15 0 16 10 9 1 0 9 14 13 10 0 9 2
7 15 4 0 9 13 0 2
25 0 9 13 10 9 14 13 6 2 10 9 15 13 15 13 14 3 3 0 16 15 13 14 13 2
22 3 14 13 1 15 1 10 0 9 1 9 7 9 2 7 10 0 9 1 15 9 2
8 7 15 13 15 3 1 3 2
13 3 13 0 16 15 13 10 0 9 1 0 9 2
4 9 13 1 15
4 9 13 3 0
4 0 9 7 9
4 0 9 0 9
5 15 13 10 9 2
5 0 9 7 0 9
5 0 9 14 13 2
5 0 0 9 3 2
5 0 9 1 11 2
5 8 0 1 0 9
5 3 8 0 9 2
6 0 2 0 9 9 2
6 0 9 7 0 9 2
6 0 9 1 9 3 2
6 0 2 0 2 0 9
6 10 9 13 1 9 9
6 13 15 4 13 15 1
7 10 9 2 7 0 9 2
7 0 11 9 1 10 9 2
7 10 3 0 2 0 9 2
7 3 13 9 1 0 9 2
8 0 9 7 9 1 10 0 9
8 0 2 13 15 0 1 9 2
8 15 15 13 2 15 4 13 2
8 0 9 0 9 1 10 0 9
9 0 9 9 9 1 10 0 9 2
4 0 9 9 2
5 7 10 0 9 2
9 0 9 2 0 9 7 0 9 2
9 0 9 9 7 9 9 1 9 2
9 10 11 14 11 9 13 3 0 2
5 15 13 10 9 2
5 15 13 10 9 2
6 0 9 2 0 9 2
4 3 10 9 2
1 0
4 9 13 0 2
5 15 13 3 11 2
2 0 9
8 0 9 1 10 9 7 0 15
10 10 1 10 0 9 7 3 0 9 9
6 0 9 7 0 9 2
5 13 15 10 9 2
11 13 9 2 10 0 9 14 13 10 9 2
4 15 13 0 2
8 15 4 14 13 1 9 0 2
4 0 7 0 2
7 0 9 9 13 15 9 2
1 13
4 11 11 13 2
6 11 11 13 15 9 2
3 0 11 2
8 9 16 13 15 9 9 10 5
12 3 0 10 0 7 0 9 13 1 10 9 2
9 10 9 1 9 7 3 0 9 2
4 10 9 14 13
4 11 1 11 2
8 3 15 0 9 1 11 2 11
2 3 0
11 10 9 13 0 2 7 10 9 13 0 2
13 0 7 0 9 1 0 9 9 3 1 10 9 2
13 0 9 1 9 9 2 9 6 2 9 9 6 2
7 15 13 3 0 7 0 2
3 3 0 2
3 0 9 2
6 0 9 13 3 0 2
4 9 13 0 2
4 4 14 13 2
1 11
11 11 11 11 11 11 2 9 1 11 11 2
9 11 11 13 0 9 7 0 9 2
4 3 13 15 2
13 13 1 0 9 10 11 4 13 0 9 1 0 9
14 16 15 4 13 1 0 0 9 2 15 4 14 13 15
1 6
14 4 14 13 0 7 0 2 3 15 4 4 13 0 2
3 0 9 2
12 11 7 11 13 3 0 7 1 9 1 9 2
3 13 10 9
12 15 13 10 0 9 14 13 9 9 9 1 2
6 0 9 7 0 9 2
9 15 13 9 3 7 15 13 10 9
14 0 9 14 13 3 1 10 9 1 9 7 10 9 2
3 0 9 2
7 3 10 9 9 4 13 2
10 5 15 13 10 0 9 1 10 9 2
5 9 14 13 1 2
9 10 9 1 10 9 4 13 0 2
3 10 9 2
5 15 0 0 9 2
12 9 13 0 7 10 9 13 1 10 9 9 2
6 0 9 7 9 9 2
11 0 9 7 9 13 1 9 1 10 9 2
10 0 7 0 1 0 9 7 0 9 2
7 9 3 13 10 9 1 3
6 15 13 10 0 9 2
3 0 9 2
9 3 1 10 2 15 9 13 15 2
1 11
16 10 9 13 0 11 13 10 0 9 9 13 0 7 9 13 0
1 5
17 15 4 3 13 15 1 9 1 9 1 7 13 1 10 0 9 2
2 9 5
16 15 13 1 3 10 0 9 1 12 9 2 13 15 15 13 2
1 11
16 10 9 10 13 0 9 9 2 9 9 2 9 13 9 2 8
13 13 13 2 13 13 11 2 1 11 12 0 9 2
5 6 2 0 9 2
4 9 4 13 2
14 4 13 1 12 11 11 11 2 11 12 2 12 2 12
11 0 9 2 0 1 10 11 11 11 9 2
8 0 9 9 9 2 3 13 2
2 0 2
14 13 10 15 9 2 7 13 15 3 3 15 13 9 2
3 3 13 2
9 9 13 0 2 0 2 7 0 2
4 9 13 0 2
8 13 3 12 9 1 11 11 2
5 0 9 9 7 9
15 15 0 4 4 13 2 2 11 14 11 13 10 0 2 2
11 14 0 2 14 0 2 3 0 9 9 2
10 3 14 13 14 13 10 9 1 3 2
10 3 0 9 1 10 9 1 0 3 2
2 0 2
10 3 0 9 1 10 9 1 0 3 2
5 15 13 10 0 2
7 3 13 1 15 9 9 2
5 15 13 3 0 2
4 13 15 9 2
1 0
8 0 9 13 15 10 0 9 2
6 0 2 0 2 0 2
7 13 10 9 1 15 2 5
2 0 9
11 10 9 13 1 11 9 3 1 11 9 2
8 6 13 10 9 1 15 9 2
3 0 9 2
6 0 9 2 0 9 2
14 9 0 1 10 0 9 9 1 9 2 9 2 9 2
2 0 2
7 15 13 9 13 7 13 2
4 15 13 0 2
6 3 13 7 13 13 2
3 1 11 11
3 0 9 2
19 9 0 0 9 9 2 0 2 0 2 0 2 8 2 13 9 13 3 2
12 5 12 13 9 1 9 14 13 1 10 9 2
6 0 9 9 1 3 2
6 15 13 15 9 3 2
13 15 13 10 9 9 1 15 11 11 10 13 0 2
10 15 3 13 9 2 9 7 9 0 2
23 15 13 10 0 0 9 1 10 11 11 2 15 13 9 15 13 1 0 11 14 13 3 2
24 10 0 9 3 15 13 0 3 15 4 13 10 9 1 9 0 1 9 1 11 15 13 10 0
3 0 9 2
13 15 4 13 15 3 7 4 13 15 1 10 9 2
9 0 9 2 0 9 7 0 9 2
6 15 13 1 1 9 2
6 0 9 2 15 13 2
12 9 4 3 13 1 11 11 11 1 10 9 2
1 0
5 0 9 3 0 2
18 15 13 15 13 0 14 13 9 13 3 3 14 13 9 1 9 9 2
4 14 10 9 9
20 13 3 0 3 15 13 9 2 15 13 10 9 9 2 3 11 10 9 9 2
2 0 9
9 0 0 9 10 15 4 3 13 2
8 9 13 3 0 7 3 0 2
6 9 13 3 3 0 2
2 0 9
10 10 3 3 13 9 1 10 0 9 2
12 10 3 13 7 4 4 13 3 1 10 9 2
1 9
14 15 13 10 9 9 13 3 7 15 13 1 1 9 2
12 15 4 4 13 9 1 15 9 14 0 9 2
4 10 0 9 2
12 11 13 10 9 7 4 3 13 1 10 9 2
11 15 13 14 13 15 14 13 15 9 13 2
13 0 9 2 0 1 10 9 7 0 1 10 9 2
10 10 9 9 9 13 3 0 7 0 2
4 13 0 9 2
3 9 13 2
8 13 1 7 0 9 13 3 2
9 13 10 0 9 13 16 15 13 2
7 13 9 7 13 3 3 2
5 0 9 1 9 2
7 9 13 0 7 3 0 2
15 15 13 12 9 9 3 7 13 15 10 13 1 10 9 2
9 15 13 0 9 1 10 0 9 2
7 15 9 3 3 1 11 2
12 9 13 1 10 0 9 7 9 13 3 0 2
7 15 4 3 13 11 11 2
21 9 13 3 0 2 4 14 13 15 2 7 4 14 13 13 3 1 10 0 9 2
7 0 9 7 3 0 9 2
9 3 0 1 15 12 9 0 9 2
7 0 0 9 9 9 3 2
5 9 10 9 0 2
2 9 0
19 3 3 13 10 9 3 0 7 0 2 7 15 3 4 14 13 10 9 2
7 10 9 13 10 0 9 2
6 15 0 9 14 13 2
23 10 9 13 10 0 2 0 9 2 9 2 0 7 0 9 2 7 10 9 13 0 3 2
3 0 9 9
14 15 13 3 0 1 10 9 9 11 11 11 13 15 2
11 3 15 13 0 14 13 10 9 3 3 2
3 0 9 2
12 15 13 10 0 9 9 15 13 1 11 11 2
2 6 2
9 15 9 7 9 4 14 13 0 2
3 3 13 2
27 0 9 9 9 13 3 0 10 9 9 13 0 9 3 8 13 13 0 0 9 3 7 9 4 13 8 3
9 15 4 3 13 1 10 0 9 2
12 15 4 13 3 12 9 13 1 12 0 9 2
8 15 4 3 13 0 7 0 2
2 0 2
3 0 9 0
6 10 9 3 13 0 2
13 9 9 13 15 9 0 7 0 3 13 11 11 2
5 13 0 3 13 3
4 0 0 9 9
5 0 0 9 9 2
11 11 7 10 9 4 13 3 9 15 13 2
10 10 9 4 13 3 1 10 11 11 2
8 0 9 7 9 1 10 9 2
5 10 10 0 9 2
12 10 9 13 0 7 15 4 13 0 7 0 2
6 15 3 13 10 9 2
11 10 9 13 0 7 3 13 1 0 9 2
8 10 9 13 0 7 13 0 2
5 0 9 7 9 2
8 15 4 13 3 3 7 3 2
7 0 9 7 9 10 13 2
12 15 13 0 1 10 9 10 15 13 1 11 2
12 10 9 13 3 0 7 15 9 13 3 0 2
4 0 9 0 9
12 15 13 3 0 9 7 0 9 14 13 3 2
8 15 13 3 3 14 13 3 2
7 10 0 9 14 13 15 11
3 0 9 9
12 0 9 14 13 10 9 7 13 1 1 9 2
7 0 0 9 7 0 9 2
10 9 13 3 0 9 7 13 0 9 2
2 0 9
21 16 13 10 9 15 0 9 9 13 10 9 4 14 4 13 16 15 4 4 13 2
8 15 4 13 3 13 10 9 2
2 9 13
6 4 14 13 10 9 2
13 15 4 13 15 12 9 3 5 12 3 13 10 2
9 13 3 1 15 9 3 13 15 2
3 13 3 2
2 0 9
30 15 13 10 0 9 0 9 7 13 10 9 16 15 13 10 0 15 13 3 0 9 1 10 11 9 2 9 3 9 2
13 15 13 10 9 9 9 1 11 1 10 9 9 2
9 10 9 4 13 1 10 9 11 2
9 3 15 13 10 9 7 13 15 2
3 0 9 2
1 9
24 3 15 9 13 2 11 13 1 12 9 1 12 9 7 13 15 9 3 7 13 10 0 9 2
8 15 13 15 15 13 9 9 2
5 15 13 0 1 2
29 15 13 0 1 0 2 9 9 2 7 1 9 1 11 11 2 11 2 7 0 9 9 9 1 10 9 2 3 2
3 9 9 2
6 12 9 1 9 9 2
2 0 2
10 4 14 13 15 4 3 4 13 3 2
13 6 2 7 9 9 2 7 9 2 1 10 9 2
2 13 2
7 11 11 1 0 11 14 9
7 11 14 11 13 3 0 2
20 15 9 2 10 9 9 1 11 11 7 11 11 2 13 3 9 1 11 11 2
9 3 2 3 2 0 9 9 9 2
9 13 10 9 3 7 3 16 0 2
11 4 12 5 13 1 9 1 10 0 9 2
7 13 15 11 14 11 11 2
4 10 0 9 2
6 11 11 11 13 0 2
9 3 0 7 3 0 3 1 9 2
7 15 4 13 14 13 9 2
4 9 3 11 2
6 9 13 10 0 9 2
6 11 14 0 9 9 2
14 15 9 13 0 14 13 10 0 12 9 1 12 9 2
15 10 0 9 9 1 9 13 9 1 0 2 9 9 9 2
14 9 2 3 0 1 10 9 9 10 13 14 0 9 2
8 9 2 10 9 13 3 0 2
14 9 13 3 0 2 10 9 1 9 13 9 1 10 9
3 0 9 2
11 15 13 0 1 10 9 0 1 10 9 2
22 15 13 3 0 9 3 1 10 9 2 3 13 2 4 14 13 14 13 15 0 9 9
2 0 9
13 15 13 14 3 10 11 11 11 11 11 4 13 2
20 15 13 2 3 2 1 10 11 11 11 2 10 9 1 10 9 1 10 9 2
24 10 10 0 9 15 13 2 3 0 14 13 7 13 2 10 9 2 10 9 3 10 9 9 2
13 13 1 10 9 13 10 0 9 9 15 4 13 2
2 3 0
34 10 9 1 2 0 9 1 9 2 4 4 3 13 1 2 0 9 1 9 2 3 0 2 0 2 0 2 0 2 7 0 9 9 2
7 0 9 9 1 10 9 2
14 11 4 4 13 1 10 9 1 10 9 9 3 3 2
16 16 15 13 10 9 11 15 4 13 5 12 3 1 9 1 9
4 11 11 13 0
16 15 9 4 4 13 11 11 1 15 9 1 10 0 12 9 2
8 15 4 14 13 1 9 0 2
9 9 1 9 13 3 0 7 0 2
10 13 1 10 9 9 3 1 11 12 2
5 6 10 0 9 2
7 10 9 7 9 13 0 2
15 15 3 13 11 11 16 15 4 13 1 9 1 11 11 2
19 3 2 10 0 9 9 9 13 10 0 9 15 4 13 1 10 11 9 2
7 15 13 0 7 3 0 2
12 15 4 13 10 9 3 1 15 9 2 6 2
4 0 11 11 9
6 15 13 10 0 9 2
8 10 10 0 9 7 0 9 2
8 11 11 11 13 10 0 9 2
4 0 0 9 2
8 13 2 15 16 13 15 9 2
4 0 9 9 2
5 9 13 9 0 2
8 0 16 15 13 1 10 9 2
12 7 3 2 15 4 13 0 16 15 15 13 2
11 13 10 9 2 4 14 13 10 9 9 2
16 11 2 10 9 2 13 3 3 14 13 15 13 0 1 9 2
12 0 7 0 2 3 3 15 9 7 9 9 2
11 15 13 10 11 5 7 3 13 15 9 2
5 3 0 9 9 2
34 15 13 10 9 0 9 13 3 2 7 10 0 13 3 0 2 3 3 1 0 2 15 13 3 14 13 10 9 13 1 1 15 9 2
5 13 15 10 9 2
8 10 9 13 0 7 3 0 2
20 15 13 15 0 9 9 14 13 1 2 7 15 13 10 0 2 9 13 9 2
7 3 3 0 4 15 13 2
24 15 13 10 9 3 7 10 9 13 0 2 3 10 9 13 3 0 0 16 15 13 3 0 2
8 15 4 13 14 13 3 0 2
5 3 0 10 9 2
1 8
2 0 9
5 11 11 13 0 2
15 15 13 10 9 13 7 13 10 0 9 15 4 3 13 2
14 15 13 10 0 0 9 7 15 13 15 1 10 9 2
4 0 9 11 2
33 13 14 13 16 15 13 10 9 15 4 4 13 1 15 9 1 9 2 10 9 15 13 10 9 4 14 3 4 13 0 1 15 2
7 15 4 3 13 3 3 2
6 15 13 10 0 9 2
22 15 4 13 11 11 14 9 3 7 15 13 3 0 16 3 0 7 0 10 9 13 2
13 15 13 10 9 14 13 3 0 7 0 2 13 2
5 13 10 0 9 2
8 10 9 4 14 4 13 3 2
18 9 9 13 9 7 9 1 9 2 3 10 9 13 0 1 10 9 2
7 3 10 0 9 9 3 2
4 15 13 15 2
11 11 13 10 0 9 15 4 3 13 1 2
21 15 13 10 0 9 1 9 7 13 0 14 13 15 9 3 3 1 0 0 9 2
9 15 4 14 4 13 1 15 9 2
6 11 14 11 2 15 9
8 11 14 11 13 3 3 0 2
12 15 13 15 4 13 10 9 1 10 0 9 2
16 3 15 13 3 3 2 3 15 4 13 15 1 9 2 9 2
19 11 11 4 4 13 15 9 1 10 9 9 3 7 15 4 13 3 0 2
19 15 4 3 13 12 0 9 14 13 1 7 15 13 3 0 1 15 9 2
3 3 13 2
2 0 9
13 10 9 13 10 0 0 2 0 2 9 14 13 2
10 11 13 10 0 9 15 13 0 9 2
12 15 9 13 0 7 10 9 1 9 13 0 2
4 4 13 3 2
2 11 2
10 11 11 11 2 9 1 10 15 9 2
15 11 11 11 2 9 16 13 15 10 9 1 10 0 9 2
17 15 13 10 0 9 2 15 9 13 0 7 15 4 13 15 3 2
5 10 0 9 1 11
25 15 13 3 0 14 4 13 11 14 9 9 2 10 10 0 7 0 9 7 10 9 14 13 1 2
6 10 9 13 1 0 2
5 15 3 13 15 5
2 0 9
17 13 1 1 10 9 16 1 1 9 1 9 2 7 15 13 0 2
10 10 9 13 0 7 10 9 13 0 2
16 15 13 10 9 9 9 1 9 2 7 15 13 3 0 15 2
12 0 0 7 3 0 9 1 9 1 0 0 9
8 0 9 1 9 1 0 9 2
17 9 13 3 0 15 13 15 1 10 0 9 7 3 3 10 9 2
7 3 0 16 13 0 9 2
12 10 0 9 1 11 16 13 9 7 9 9 2
18 1 0 9 1 15 1 9 1 15 9 2 9 13 3 7 1 9 2
9 3 0 16 15 13 14 13 9 2
6 0 1 11 3 3 2
14 0 9 14 13 15 13 9 11 11 11 7 11 11 2
21 15 4 13 15 1 9 7 9 2 9 7 15 13 0 7 13 10 9 13 0 2
7 0 9 12 9 1 0 2
3 9 1 11
13 15 13 11 1 15 0 11 1 11 7 11 9 2
9 15 13 3 0 2 0 7 0 2
16 15 13 3 1 10 1 15 9 7 15 13 10 3 0 9 2
7 15 4 4 13 11 3 2
5 12 1 10 0 2
11 11 13 12 1 12 0 9 1 11 11 2
19 15 13 11 11 2 3 1 11 11 2 11 2 7 11 11 3 1 11 2
11 15 4 13 10 0 9 1 9 7 9 2
20 15 13 0 2 0 9 2 15 13 15 13 1 3 2 7 10 9 13 0 2
10 15 13 0 2 7 3 10 0 0 2
8 9 1 9 1 0 9 9 2
10 0 14 13 1 3 1 1 9 9 2
21 15 4 13 15 4 14 13 0 1 10 9 2 7 15 3 4 13 10 0 9 2
18 10 9 9 2 9 13 0 7 13 1 10 0 9 9 1 10 9 2
9 9 13 10 9 0 2 7 0 2
3 13 10 9
3 13 1 2
6 0 2 0 0 9 2
7 10 9 14 13 5 13 2
11 2 0 2 9 1 12 9 4 14 13 2
3 3 0 2
16 13 12 5 1 2 9 2 9 2 1 0 9 4 13 0 2
1 0
3 0 9 2
4 0 9 9 2
5 11 9 9 13 2
5 0 9 2 9 2
3 9 0 2
11 9 0 2 0 2 0 2 7 3 13 2
15 13 10 9 1 10 11 2 10 13 1 10 0 9 2 2
14 9 2 3 0 2 7 3 0 2 7 3 0 9 2
9 9 1 9 13 0 7 3 0 2
16 1 10 9 9 9 2 13 5 13 10 12 0 9 15 13 2
9 4 13 10 9 9 1 9 9 2
3 0 9 9
10 11 11 13 10 0 11 0 9 9 2
15 15 13 13 9 3 7 13 15 13 1 7 13 10 9 2
17 16 15 13 10 9 15 4 13 15 9 2 13 11 11 1 11 11
13 13 1 3 3 2 7 9 13 3 0 7 0 2
8 9 3 0 7 13 3 0 2
8 15 4 13 10 9 1 9 2
20 15 13 15 9 3 7 16 3 3 1 10 9 2 15 4 4 13 3 3 2
7 9 16 13 15 1 10 9
3 0 13 2
11 15 4 14 13 2 15 4 14 13 3 2
28 15 13 0 14 13 10 0 9 2 10 0 9 7 10 9 1 15 0 9 7 15 13 3 1 1 15 0 9
5 0 9 9 1 11
15 16 15 4 13 1 0 0 9 9 2 3 13 3 3 2
8 15 3 13 10 9 9 9 2
3 0 9 2
18 10 9 5 9 2 2 11 11 2 13 10 9 14 13 1 3 3 2
1 11
4 0 0 9 2
16 10 10 0 9 1 10 9 1 10 9 15 4 14 13 15 2
8 0 2 0 9 2 0 9 2
8 3 3 2 10 9 13 0 2
9 15 3 4 4 13 1 0 9 2
6 15 4 13 3 3 2
5 9 1 10 0 9
44 9 1 10 0 9 7 0 9 15 7 15 9 4 13 1 15 0 0 9 2 10 9 1 10 9 13 0 7 10 9 15 4 13 3 8 1 10 9 13 0 2 0 9 9
3 0 3 0
21 10 0 9 15 13 1 3 1 15 9 9 9 15 13 15 4 13 3 10 9 2
24 11 11 13 0 9 2 10 0 9 9 2 7 9 15 13 14 13 15 9 1 0 0 9 2
3 0 9 2
17 15 13 3 0 16 15 3 13 10 0 9 9 1 11 11 11 2
14 3 3 13 14 13 1 11 11 1 10 0 9 9 2
7 7 11 7 11 13 0 2
9 15 4 3 13 15 9 7 9 5
3 0 2 5
20 15 13 10 3 0 9 1 10 9 7 15 13 3 9 1 9 2 0 9 2
27 13 10 12 9 15 13 1 10 11 11 1 10 0 9 10 9 9 9 13 3 10 9 9 9 1 10 9
5 0 9 0 9 2
6 2 10 9 13 0 2
9 15 13 13 3 7 14 4 13 2
18 15 13 3 3 15 13 10 0 9 1 11 7 15 13 10 0 9 2
14 10 9 15 13 3 13 16 10 9 13 3 0 2 2
4 0 9 9 2
12 15 13 3 14 13 10 0 9 1 15 9 2
25 10 12 9 15 13 3 2 15 4 13 13 10 9 2 13 3 10 3 0 9 15 4 3 13 2
10 7 3 15 13 0 9 9 1 11 2
2 0 9
22 10 10 9 14 13 1 0 11 11 1 11 11 1 10 9 1 10 0 9 1 9 2
9 11 11 14 9 9 13 15 9 2
8 10 9 11 13 0 7 0 2
10 13 15 10 9 16 13 11 11 11 2
3 0 9 2
12 15 13 12 1 15 0 9 14 13 1 9 2
31 15 13 10 0 9 1 10 0 9 2 15 13 0 9 14 13 15 1 2 7 15 4 14 3 13 16 15 13 3 0 2
7 7 2 15 13 3 0 2
51 11 13 10 0 9 2 15 4 3 13 0 9 16 3 14 13 15 9 7 9 2 14 13 10 9 10 0 9 2 13 9 7 13 15 4 13 15 2 15 4 13 1 9 15 13 10 0 1 10 0 2
17 16 15 13 3 13 9 1 11 7 11 2 15 13 14 15 9 2
11 10 9 3 13 10 3 0 0 13 9 2
12 15 9 13 0 9 7 10 9 13 3 0 2
11 13 1 10 11 11 1 10 15 9 9 2
36 11 7 11 13 3 0 2 7 3 11 14 13 14 13 1 15 9 2 11 13 3 3 7 13 10 9 7 13 15 11 14 9 4 14 13 2
12 15 13 1 15 3 1 10 9 1 15 9 2
4 15 13 3 0
3 0 7 0
50 13 3 7 13 1 1 3 1 12 9 1 10 3 0 9 15 13 15 4 13 14 4 13 10 9 16 15 13 10 9 7 1 15 9 7 9 2 12 15 13 0 14 13 15 10 0 9 3 3 2
5 13 14 10 9 9
22 15 13 10 9 9 3 7 4 14 13 9 9 7 15 4 13 10 9 9 3 3 2
12 0 15 13 16 15 13 1 15 9 14 13 2
15 13 13 10 9 4 13 9 10 9 1 10 0 9 3 2
7 10 9 13 0 3 3 2
13 10 9 13 15 9 7 3 13 15 15 10 9 2
9 14 0 3 15 13 1 10 12 2
15 15 13 0 1 10 9 2 7 10 9 13 14 3 0 2
10 16 15 13 0 9 2 13 1 11 2
2 3 2
41 9 0 13 15 10 0 0 16 15 13 14 3 12 9 1 10 9 2 10 0 9 13 1 10 9 1 10 9 2 2 7 16 15 10 13 10 0 0 9 9 2
11 7 15 13 14 4 13 1 3 0 9 2
3 0 3 2
15 15 13 1 11 14 10 10 9 7 15 4 3 4 13 2
32 9 9 13 3 0 14 13 16 15 4 14 13 2 10 13 10 9 1 15 1 2 1 10 0 9 1 9 2 7 3 0 2
3 3 0 2
3 0 0 9
5 11 13 0 9 2
15 15 13 3 0 7 13 10 9 14 13 10 9 1 15 2
17 10 9 1 15 9 4 13 3 7 15 13 15 4 13 15 9 2
9 15 13 9 1 0 9 14 13 2
6 15 3 13 15 9 2
3 0 1 11
12 10 9 13 1 3 10 0 15 4 13 1 2
28 15 13 10 11 2 10 9 13 0 1 7 15 4 13 3 0 7 9 10 9 0 1 10 0 9 15 13 2
12 15 13 10 0 9 15 4 13 15 9 9 2
12 13 10 9 3 16 10 9 9 14 4 13 2
12 9 1 10 9 13 3 16 15 13 15 3 2
12 10 9 9 4 13 7 3 10 9 13 0 2
18 9 9 4 14 13 3 13 7 10 13 9 13 10 9 3 16 13 2
10 15 4 13 1 11 1 0 9 3 2
9 15 13 3 3 12 9 10 9 2
10 15 4 3 13 10 9 1 10 9 2
6 15 13 3 3 0 2
7 10 9 4 3 13 0 2
10 11 13 10 0 9 14 13 15 9 2
5 15 13 10 9 2
4 4 14 13 0
20 15 13 14 13 1 10 9 16 15 4 13 1 10 9 1 12 1 15 9 2
2 6 2
9 15 4 14 13 15 15 4 13 2
14 10 0 9 3 13 0 1 15 0 9 14 0 9 2
8 9 13 0 7 9 13 0 2
7 0 9 7 3 0 9 2
5 0 14 13 1 2
34 1 10 0 9 2 15 13 3 0 16 15 4 3 13 2 0 9 2 9 3 3 3 9 13 3 1 0 9 7 9 1 15 9 2
6 3 13 9 2 9 2
3 9 11 2
4 9 15 4 13
15 16 0 15 13 10 9 1 15 16 15 13 3 15 9 2
5 11 11 13 9 2
18 7 15 7 15 9 4 14 13 10 0 9 16 15 13 0 9 3 2
8 10 9 9 13 9 7 9 2
6 15 0 13 15 0 2
9 15 13 14 15 0 0 9 9 2
16 15 13 10 0 9 1 0 9 7 9 15 3 13 9 9 2
12 10 9 13 1 0 9 2 10 9 13 0 2
19 10 9 13 15 0 0 9 1 0 9 9 7 9 1 10 9 7 9 2
3 8 13 2
35 15 13 15 9 14 13 10 9 1 10 9 7 10 9 1 15 9 13 5 12 7 3 15 13 1 9 14 13 15 9 15 13 5 12 2
19 15 13 9 0 7 3 10 9 13 10 9 7 1 15 15 13 14 9 2
7 11 2 15 13 10 0 2
29 10 15 4 13 13 16 11 15 13 10 0 15 4 13 2 3 3 4 10 9 13 10 0 9 16 15 13 15 2
21 15 13 15 1 9 1 11 2 16 15 13 10 9 7 10 9 1 15 13 0 2
4 12 9 9 9
28 15 13 15 11 3 7 15 13 0 16 15 13 0 2 15 13 10 0 9 2 15 13 3 0 1 10 9 2
13 10 9 7 9 13 1 9 7 10 0 13 0 2
12 3 2 15 13 0 9 9 7 10 3 0 9
