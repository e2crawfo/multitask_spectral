200 11
29 1 9 2 0 9 13 4 0 9 16 13 9 15 4 9 4 9 9 1 9 11 7 9 9 1 9 0 9 2
10 1 3 4 15 9 0 1 9 11 2
28 1 11 3 2 9 9 13 16 3 3 4 13 15 0 9 1 11 2 7 16 4 1 15 9 13 1 9 2
8 11 9 13 1 9 9 0 9
19 11 9 13 15 9 1 9 1 0 9 15 4 13 9 0 9 7 9 2
28 11 9 13 15 1 9 2 12 9 2 9 1 0 9 9 7 9 0 1 9 15 4 13 15 9 15 9 2
35 0 4 3 1 12 9 0 9 0 1 9 9 9 1 0 9 2 13 4 1 9 9 0 9 9 9 11 11 3 9 9 0 0 9 2
21 3 12 9 0 1 12 0 0 9 2 0 4 1 9 15 4 13 1 12 9 2
25 16 15 13 0 9 2 9 4 15 13 7 1 15 9 2 13 4 1 9 0 9 9 11 11 2
27 1 9 9 2 9 4 13 1 9 3 12 9 9 2 9 12 9 0 9 7 9 3 1 12 9 9 2
15 9 4 3 13 3 12 0 9 7 3 1 12 9 9 2
20 9 4 3 0 13 15 9 1 9 0 0 9 2 13 15 1 9 0 9 2
15 11 4 1 9 13 16 4 9 9 13 3 12 9 9 2
19 9 4 13 3 9 16 4 1 9 9 9 13 9 1 9 3 12 9 2
31 9 15 4 0 9 13 9 2 7 15 4 0 0 0 9 1 0 12 9 13 4 3 1 9 9 11 15 13 12 9 2
33 1 0 0 9 15 4 0 9 13 0 0 9 2 11 2 2 9 4 13 9 3 12 9 2 7 0 0 9 13 12 9 9 2
11 0 9 3 1 9 13 3 12 9 9 2
12 0 0 9 13 4 9 1 3 12 9 9 2
14 3 12 9 3 9 3 4 0 2 16 4 12 0 2
24 9 4 1 9 13 9 9 9 15 4 13 1 9 2 16 4 15 13 13 3 9 15 9 2
9 15 9 13 13 1 12 9 9 2
45 2 1 12 9 1 11 15 4 1 0 9 0 9 2 9 2 9 1 9 2 9 7 9 1 9 2 9 11 13 4 13 0 9 2 2 13 15 1 9 0 9 0 1 9 2
39 11 4 13 9 2 0 9 2 9 1 9 9 7 9 1 0 9 2 16 4 9 11 1 9 0 9 13 9 1 1 12 9 1 9 9 1 0 9 2
22 9 1 0 9 13 16 4 0 9 1 9 1 0 7 0 0 9 2 13 0 9 2
20 1 9 15 4 13 15 0 9 13 15 0 9 7 9 9 9 7 9 9 2
25 2 9 14 4 9 15 13 9 9 2 2 13 4 1 9 0 9 11 9 1 0 9 11 11 2
27 2 1 15 15 0 0 9 3 13 1 9 7 13 1 9 15 4 3 0 7 13 9 13 0 9 2 2
8 0 0 9 0 9 13 15 9
30 0 0 9 0 9 11 11 13 4 1 9 9 9 16 15 12 13 1 9 0 9 16 4 13 1 9 0 9 9 2
41 0 0 9 0 9 11 11 13 4 1 9 2 12 9 2 16 15 0 13 15 0 9 16 9 9 16 4 9 13 13 9 1 15 0 9 1 9 0 1 9 2
25 2 13 4 15 16 4 15 13 13 0 9 2 2 13 4 1 9 1 0 9 9 11 1 11 2
46 16 3 0 9 0 0 9 2 11 2 2 11 4 0 9 0 9 1 0 0 9 0 1 9 9 2 15 4 9 1 0 9 13 1 15 1 0 9 1 9 12 4 4 0 9 2
22 0 0 9 1 9 11 1 9 1 15 4 9 4 1 9 1 9 9 7 9 9 2
41 15 4 9 1 0 9 13 9 1 15 16 4 9 15 15 4 11 13 16 2 0 9 2 4 13 9 16 13 13 9 0 9 1 9 11 1 11 1 9 12 2
63 9 4 13 7 13 15 0 0 9 11 11 2 15 4 3 13 9 0 9 0 9 1 0 9 2 11 2 2 7 1 15 4 9 13 1 0 9 2 3 4 13 1 9 1 9 0 0 9 1 9 2 0 2 9 2 2 0 1 9 1 9 11 2
46 11 2 15 4 13 16 13 9 1 0 9 7 0 0 9 2 0 4 9 0 7 13 15 1 0 9 2 1 15 4 9 1 11 13 9 1 0 9 2 15 4 1 15 3 0 2
34 0 4 9 0 9 0 9 11 11 7 9 0 0 9 11 11 13 16 4 0 9 9 1 12 4 9 1 11 0 9 9 1 9 2
51 11 2 15 4 3 13 9 0 1 9 1 0 9 2 13 4 16 4 11 13 9 1 0 9 1 11 15 4 0 15 9 9 7 9 0 1 11 11 2 2 9 2 2 3 12 1 0 9 0 9 2
18 3 2 15 7 11 13 4 7 16 4 0 9 9 11 2 11 0 2
33 1 0 15 0 9 13 16 4 1 15 0 9 15 4 13 15 9 4 3 3 13 9 1 9 0 9 0 9 1 2 9 2 2
43 1 9 4 11 11 2 9 0 9 11 2 15 15 3 13 1 9 0 9 1 9 9 11 2 13 9 0 9 11 11 7 13 16 13 9 1 9 0 9 1 0 9 2
36 3 16 15 3 4 0 13 9 2 0 4 9 0 9 1 9 13 16 4 4 9 9 0 1 9 9 9 1 0 9 1 15 15 9 13 2
25 11 4 9 11 7 11 13 2 0 9 7 9 2 2 3 16 1 9 9 13 13 9 1 9 2
25 13 4 7 16 4 1 9 11 13 9 15 15 1 15 13 16 13 9 3 1 9 0 1 15 2
5 11 3 13 1 9
10 0 9 4 13 13 0 9 1 9 2
15 13 14 0 9 2 0 1 3 1 12 9 2 13 9 2
20 0 9 1 11 1 9 2 12 9 2 4 4 0 15 9 1 0 12 9 2
21 0 4 9 1 9 13 9 0 9 2 16 15 4 4 0 16 4 13 15 9 2
21 1 9 4 0 9 1 15 4 14 9 13 3 13 9 13 9 1 0 9 9 2
6 11 4 0 7 0 2
20 1 9 1 0 9 2 3 1 12 15 4 3 13 16 4 13 1 0 9 2
19 2 4 15 14 13 2 2 13 4 11 11 2 12 2 9 0 1 11 2
10 2 3 12 9 13 0 9 1 11 2
14 9 3 13 0 9 2 7 3 15 13 1 9 2 2
38 1 9 16 13 9 7 13 9 2 0 0 9 13 4 0 9 2 9 0 9 2 0 12 9 1 9 9 2 7 9 4 13 9 3 13 1 9 2
24 2 3 4 15 15 13 1 9 2 2 13 4 9 11 11 11 2 12 2 2 9 9 9 2
16 2 3 2 1 9 4 3 12 9 2 7 9 15 4 0 2
18 13 4 13 9 7 9 7 9 9 13 16 4 13 15 15 13 2 2
17 9 1 11 0 4 1 12 0 9 2 0 7 15 0 1 11 2
21 1 9 13 0 9 7 9 15 13 0 9 2 16 0 13 9 1 0 9 11 2
27 2 1 9 9 13 3 0 0 9 9 2 2 13 0 9 9 1 0 9 7 9 9 0 9 11 11 2
21 2 15 4 3 0 1 9 2 3 16 13 13 1 9 9 16 4 13 9 2 2
12 0 9 1 11 3 4 3 0 1 0 9 2
41 2 13 9 15 4 3 4 1 9 7 0 4 1 9 7 4 3 13 15 9 0 1 9 16 4 13 9 0 9 2 2 13 11 11 1 0 9 1 0 9 2
19 2 9 4 3 0 7 3 4 13 0 9 0 0 9 3 1 15 9 2
21 1 15 4 0 9 13 1 0 0 9 2 7 14 7 1 11 2 2 13 4 2
22 7 0 9 13 0 9 2 1 15 7 11 7 0 0 9 13 9 0 9 1 9 2
22 0 9 0 4 9 13 9 15 15 13 0 9 11 7 15 13 9 0 7 0 9 2
41 2 11 4 13 0 0 7 0 9 16 4 15 13 15 9 2 15 9 4 0 3 1 11 2 3 7 1 9 1 9 2 2 13 4 9 11 11 2 11 2 2
28 2 13 15 16 4 9 11 12 9 13 9 1 0 0 9 2 1 15 4 13 9 0 1 9 0 9 2 2
23 3 2 15 4 15 9 3 13 1 9 2 1 15 4 15 3 13 9 7 0 0 9 2
29 2 1 9 13 0 9 7 9 13 4 3 0 1 0 9 2 2 13 4 11 11 2 9 9 1 9 1 9 2
17 3 4 12 9 7 12 0 9 15 15 13 1 12 9 1 9 2
16 1 0 9 9 2 9 1 15 9 13 12 1 12 0 9 2
5 0 9 13 15 9
21 11 11 13 4 9 1 9 9 0 9 1 11 7 11 1 0 9 7 9 11 2
45 0 9 1 11 7 11 2 11 2 11 11 13 4 4 1 9 2 12 9 2 16 4 13 9 15 0 9 1 0 7 9 11 16 15 0 9 13 1 15 9 1 9 1 11 2
30 1 9 9 9 0 9 2 11 2 13 4 1 9 9 15 4 1 9 13 1 9 11 9 0 9 11 2 11 2 2
42 15 9 13 9 15 4 13 9 1 9 9 2 11 2 1 0 9 1 11 7 2 0 9 15 11 13 1 9 1 9 9 1 0 9 2 2 0 4 1 9 11 2
33 11 4 0 1 9 12 9 16 0 9 0 1 9 0 9 0 0 9 15 4 0 9 1 11 15 4 13 1 12 1 12 9 2
21 0 9 2 0 9 0 9 1 9 2 13 0 9 15 15 13 9 9 7 9 2
16 13 13 3 7 0 9 2 16 13 16 13 0 9 1 11 2
53 2 0 4 16 4 3 1 9 1 15 13 13 9 9 9 1 9 11 7 0 9 0 9 16 15 4 11 7 0 9 2 16 15 4 4 9 1 0 9 1 9 2 2 13 4 11 2 13 15 1 9 11 2
27 11 4 3 1 9 9 1 11 1 9 1 9 7 9 7 9 1 9 11 9 1 9 2 13 4 11 2
28 3 3 4 15 13 9 1 9 9 13 4 1 0 9 1 11 7 9 9 16 13 9 2 13 15 1 9 2
15 11 13 9 1 9 0 0 9 11 16 4 13 9 9 2
27 1 0 9 1 11 2 11 3 13 0 9 1 11 11 2 11 2 11 2 11 7 12 0 9 1 11 2
50 9 9 11 0 4 1 3 1 9 1 9 1 12 9 3 4 4 0 2 13 4 0 9 2 3 3 1 9 1 9 3 1 12 9 9 1 15 9 1 12 9 2 15 13 3 1 12 9 9 2
15 9 1 12 13 4 3 9 9 11 1 1 12 9 9 2
45 0 9 9 2 13 15 1 9 0 9 2 2 4 4 0 9 1 9 11 2 9 1 15 11 1 9 13 15 9 1 0 9 2 7 3 15 13 3 1 0 9 1 11 2 2
9 9 7 9 2 11 13 9 1 11
19 11 11 13 4 1 11 16 4 13 9 0 2 0 9 2 15 0 9 2
13 3 15 9 2 9 9 11 11 11 13 15 9 2
20 9 11 11 11 13 1 9 1 0 9 11 11 1 9 1 9 11 1 11 2
22 9 11 11 11 13 4 1 9 2 12 9 2 1 11 9 9 0 2 0 9 2 2
24 9 15 13 1 9 11 7 13 4 9 0 0 9 7 0 9 2 7 3 4 13 9 9 2
24 9 9 11 7 11 11 11 13 4 15 9 1 9 11 2 0 4 1 9 2 12 9 2 2
16 15 0 9 1 9 4 4 1 9 9 0 9 1 12 9 2
32 8 8 8 13 4 1 9 2 12 9 2 16 4 13 12 0 9 7 12 0 9 0 7 0 9 1 0 9 11 7 11 2
20 9 4 9 9 8 8 8 15 4 9 9 9 1 9 1 9 1 9 9 2
28 0 9 2 3 1 9 1 0 0 9 2 11 7 11 11 2 13 4 16 15 11 13 11 1 12 9 3 2
26 16 15 9 13 2 11 7 11 13 4 15 1 3 12 1 12 9 9 2 15 4 13 9 0 9 2
33 9 0 11 7 11 1 11 13 4 12 9 2 1 9 0 9 2 0 9 2 9 7 9 2 1 11 11 2 7 0 0 11 2
12 13 15 16 4 9 9 13 1 0 0 9 2
9 9 9 13 15 1 9 1 0 9
16 9 9 12 9 9 11 15 13 9 13 15 1 0 9 9 2
36 9 9 9 13 4 15 1 9 2 12 9 2 16 4 0 9 1 0 9 15 4 4 0 1 9 12 9 1 12 9 13 3 12 9 9 2
41 9 0 9 2 11 2 2 16 4 0 9 1 9 9 9 1 0 9 4 0 2 13 4 0 9 0 0 9 2 11 2 15 4 13 1 9 1 9 12 9 2
44 1 0 9 1 12 9 9 2 0 9 9 11 0 4 1 3 3 12 9 9 2 16 0 9 9 13 4 0 16 4 15 9 0 9 13 0 7 13 16 9 9 13 0 2
30 3 2 9 9 13 3 13 9 1 9 9 0 0 9 2 11 2 15 3 13 12 9 9 7 15 4 0 9 11 2
40 3 1 9 9 9 1 11 1 9 2 0 9 11 11 2 0 9 2 13 4 9 16 4 0 9 0 1 9 4 1 9 1 9 9 9 15 4 1 9 2
31 2 3 4 15 13 1 9 9 9 11 2 2 13 4 2 3 16 4 9 4 0 2 0 9 2 3 15 12 9 2 2
24 11 4 3 13 9 16 4 12 9 9 4 0 1 9 0 9 9 9 15 4 3 0 9 2
12 2 13 16 4 15 4 0 2 2 13 4 2
31 1 9 9 2 11 3 4 13 9 1 11 7 3 1 0 9 0 9 11 15 15 4 3 3 13 9 9 15 13 9 2
47 16 4 13 16 3 3 4 4 9 1 11 1 15 9 0 9 1 9 2 9 11 1 0 7 0 9 11 11 13 4 16 4 1 12 9 9 13 13 1 15 0 9 1 9 1 11 2
40 2 0 9 1 11 4 16 13 4 12 9 1 12 9 15 11 0 13 15 9 2 16 15 4 15 2 3 2 13 1 9 11 7 11 2 2 13 4 11 2
29 11 4 2 3 2 3 13 1 9 16 9 1 9 4 0 2 3 16 4 0 0 9 1 0 0 9 1 9 2
32 9 9 3 4 13 13 1 9 1 2 9 9 2 15 4 3 15 9 13 11 7 11 1 9 1 15 9 9 1 11 9 2
14 2 15 4 0 16 4 0 0 2 2 13 4 11 2
28 0 0 9 3 15 13 1 9 1 9 7 9 2 9 0 9 1 0 9 7 9 0 9 1 9 1 9 2
10 15 9 13 4 9 0 9 9 9 2
28 2 3 0 13 9 9 2 7 15 4 9 16 15 15 13 2 2 2 13 15 1 9 0 9 9 11 11 2
11 2 4 0 16 4 0 9 0 9 2 2
18 13 15 16 4 9 4 0 1 0 9 9 12 9 9 9 12 9 2
31 1 15 3 4 13 9 9 9 12 9 3 2 1 0 9 11 12 7 12 9 2 3 15 13 9 0 9 1 0 9 2
4 11 11 1 9
13 9 1 12 0 9 1 0 9 13 4 13 9 2
32 1 3 9 0 9 15 4 0 1 0 9 2 0 9 11 11 13 4 1 9 2 12 9 2 9 1 9 15 9 11 11 2
30 11 4 13 1 0 9 16 9 4 1 9 13 1 0 9 2 7 15 13 13 2 15 9 9 15 13 9 9 2 2
21 0 9 9 9 11 11 7 9 1 0 0 9 11 11 3 4 4 0 15 9 2
7 9 4 13 1 15 8 2
17 9 1 0 9 9 11 11 11 7 0 11 11 13 0 9 0 2
23 0 9 13 0 9 1 9 7 2 1 9 9 2 0 12 9 14 4 13 9 13 4 2
36 11 4 13 1 0 9 16 4 13 9 9 7 16 4 15 9 13 1 9 2 7 2 13 4 2 9 13 0 9 7 13 13 1 0 9 2
39 11 9 13 4 1 9 9 1 15 15 13 16 15 9 0 1 9 14 13 1 9 9 2 16 15 13 0 0 0 9 2 15 13 0 7 0 9 2 2
5 9 4 3 13 2
26 11 4 13 15 9 2 15 4 0 1 9 2 16 4 0 1 0 9 2 15 3 13 3 12 9 2
15 9 1 11 13 16 4 0 9 13 9 7 0 0 9 2
37 2 9 15 4 0 11 13 9 1 0 9 2 0 9 7 0 9 2 15 9 14 13 7 12 1 15 9 2 2 13 1 11 9 11 11 11 2
20 11 4 1 9 0 9 2 16 4 9 0 9 2 0 9 2 2 13 4 2
30 2 9 0 9 13 16 11 13 9 1 9 1 11 7 16 13 0 9 9 11 2 15 4 3 13 13 1 0 9 2
26 3 2 13 15 9 13 14 15 13 2 16 4 15 9 1 0 9 7 11 9 0 2 2 13 4 2
12 11 11 1 9 1 0 9 7 9 13 15 2
19 13 16 4 15 9 1 9 13 1 9 9 16 13 9 1 9 0 9 2
13 2 14 13 3 13 16 4 15 9 9 1 9 2
35 3 2 0 9 4 15 15 4 9 0 12 9 1 0 9 9 2 7 15 4 0 9 1 9 11 1 11 2 2 13 4 11 1 11 2
9 11 13 9 2 0 9 2 1 11
9 11 15 13 13 0 9 1 11 2
34 9 0 9 2 9 0 9 11 11 13 4 0 9 9 9 0 11 2 11 2 15 4 13 12 0 0 9 1 11 2 1 11 11 2
21 9 4 13 7 0 9 16 15 13 0 9 7 3 13 1 9 2 13 4 11 2
26 2 0 9 4 4 3 0 9 2 7 0 9 13 15 1 15 2 2 13 4 11 1 15 9 11 2
24 9 0 9 13 4 1 9 1 11 7 11 2 11 2 2 3 15 13 1 0 7 0 9 2
32 2 11 4 4 0 3 16 3 13 7 13 1 0 9 1 0 9 2 2 13 4 1 11 11 11 2 9 9 11 11 11 2
12 2 13 0 9 1 11 2 2 13 4 11 2
12 2 15 9 4 1 0 9 15 0 9 2 2
23 16 15 9 11 1 9 13 1 0 9 11 2 9 1 11 13 13 0 9 11 1 11 2
40 2 13 13 15 9 1 0 11 2 7 3 7 3 2 2 13 0 9 11 11 11 2 15 4 13 9 7 1 0 11 2 3 9 11 16 2 0 9 2 2
33 2 11 4 13 9 2 15 3 13 2 1 9 11 2 7 1 0 9 13 4 3 0 9 1 11 2 2 13 4 11 1 11 2
38 2 0 9 2 9 9 7 9 1 0 2 0 4 9 11 1 11 2 13 4 11 11 2 9 9 8 2 9 2 2 1 9 11 1 0 0 9 2
16 11 13 16 4 11 0 13 9 9 1 15 0 9 7 9 2
38 11 11 2 0 9 1 0 9 7 9 2 3 15 13 16 4 15 2 7 11 13 9 0 0 9 1 0 11 2 11 3 13 3 3 13 1 9 2
28 2 3 4 15 9 13 2 1 0 2 13 0 0 9 2 11 7 11 1 9 2 2 13 4 11 1 11 2
28 2 9 4 15 9 1 11 7 11 2 15 4 9 3 0 2 16 7 9 0 9 2 11 14 13 13 2 2
27 11 2 3 2 13 16 15 11 7 3 13 1 3 0 0 9 1 9 2 7 3 13 9 11 7 11 2
30 2 13 16 4 9 0 9 4 0 1 0 9 15 15 9 13 13 1 9 2 15 3 13 0 9 2 2 13 4 2
7 9 9 0 11 1 9 9
21 9 15 13 0 9 9 1 0 11 2 7 13 0 9 1 9 9 1 0 9 2
33 3 2 1 9 16 4 9 0 9 3 0 2 1 9 0 9 2 2 9 1 0 9 13 4 1 0 9 7 9 0 0 9 2
12 8 8 8 4 13 0 9 7 9 1 9 2
20 13 14 9 9 3 3 12 1 0 9 0 9 1 9 0 11 2 11 2 2
23 0 15 9 1 15 9 13 1 9 11 2 9 0 11 2 2 15 4 3 0 16 9 2
30 3 15 1 9 1 15 0 9 4 13 9 9 2 9 4 9 1 9 9 13 0 9 9 0 9 1 0 12 9 2
19 9 9 0 9 3 4 0 1 0 9 7 0 9 9 1 9 3 9 2
17 0 4 9 16 9 13 0 9 9 9 0 9 2 7 9 9 2
17 3 2 9 13 0 9 7 0 3 0 9 9 2 0 0 9 2
19 3 2 15 3 13 0 9 9 9 7 0 9 9 0 0 9 1 9 2
32 16 4 1 15 0 9 9 3 13 9 2 3 9 9 1 0 9 15 4 13 3 1 0 9 9 2 3 4 13 0 9 2
21 9 0 9 1 11 4 0 2 16 15 4 0 1 3 0 9 0 1 9 11 2
18 11 4 1 9 12 13 16 13 9 0 9 1 12 9 1 9 9 2
23 9 4 13 7 9 9 0 9 1 9 1 12 9 7 9 0 0 0 9 1 0 9 2
29 11 7 11 2 11 2 2 7 11 7 11 11 2 1 15 4 9 9 0 3 2 3 15 13 3 1 3 9 2
8 3 13 1 9 9 0 9 2
33 3 1 0 9 2 9 9 4 1 9 3 4 15 0 4 0 7 0 0 2 1 15 4 13 9 2 0 9 7 0 0 9 2
7 15 15 13 13 0 9 2
29 9 9 11 2 15 4 9 1 12 1 12 2 13 0 9 9 0 9 2 3 0 9 13 4 1 12 7 12 2
19 11 2 7 11 7 11 11 13 4 9 12 1 9 16 4 9 3 0 2
18 9 9 1 9 0 11 3 13 1 9 1 0 9 9 7 9 9 2
10 9 1 15 9 13 4 0 9 9 2
33 11 2 11 2 11 7 11 13 4 16 0 9 9 1 9 9 7 9 2 16 4 11 2 7 11 7 11 11 3 13 0 9 2
10 1 0 9 16 0 9 13 15 11 2
30 1 11 4 2 1 3 0 9 0 1 9 9 7 0 9 9 2 0 9 1 9 0 16 9 9 9 1 0 9 2
10 9 0 9 3 4 12 0 9 9 2
7 3 13 0 9 1 9 2
27 3 2 0 0 0 9 11 13 4 15 0 9 11 8 8 9 8 8 8 2 15 4 9 0 9 11 2
38 1 9 4 9 15 13 11 11 8 2 8 8 7 3 0 0 9 1 0 9 1 12 9 9 13 9 0 9 1 11 2 0 0 9 9 0 9 2
11 0 4 0 9 1 9 12 0 0 9 2
22 13 13 7 9 0 9 1 12 9 0 9 11 8 8 2 15 4 9 1 0 11 2
25 3 4 3 2 9 0 0 9 0 9 2 11 13 0 9 1 15 9 1 9 0 9 1 9 2
