322 11
22 12 0 0 9 11 11 7 11 11 13 3 2 16 11 4 13 1 10 2 9 2 2
12 15 13 2 16 11 9 1 9 13 1 9 2
20 1 15 1 10 9 13 15 2 2 1 10 0 9 13 9 7 0 9 13 2
21 7 16 10 9 4 0 1 14 13 1 9 1 15 2 3 13 10 9 2 15 2
19 1 10 9 13 0 9 9 1 10 9 1 9 7 3 1 0 9 2 2
22 7 15 13 2 2 3 16 15 1 3 13 10 9 1 0 9 2 13 15 1 9 2
12 13 1 9 1 9 4 15 3 13 10 0 2
7 15 13 15 3 3 3 2
10 15 13 3 3 1 9 1 9 9 2
4 9 4 0 2
29 15 13 9 7 13 1 3 1 10 9 1 9 2 15 15 3 4 13 7 3 4 13 1 14 13 0 1 2 2
11 15 13 2 16 9 4 13 9 0 9 2
3 1 11 11
13 9 1 9 1 11 4 3 13 1 9 7 9 2
13 3 4 9 1 10 0 9 13 15 10 0 9 2
28 15 13 9 9 11 11 7 13 2 16 10 0 9 13 3 1 10 9 2 15 9 3 1 9 13 14 13 2
15 11 11 13 1 11 2 3 9 13 1 9 7 0 9 2
20 2 15 4 3 13 15 1 2 16 10 0 4 13 1 11 2 2 13 15 2
18 9 1 11 0 9 2 11 2 2 11 11 2 4 3 13 1 9 2
17 11 4 3 3 13 2 16 9 13 3 3 3 1 9 1 9 2
46 3 13 11 1 10 9 10 9 1 9 7 9 2 3 10 0 1 15 1 9 13 9 1 14 13 9 2 2 15 13 15 2 2 4 9 1 9 1 11 11 7 10 0 0 9 2
21 2 15 4 0 9 2 15 4 13 3 0 10 9 1 9 2 2 13 11 11 2
13 1 0 9 1 12 9 13 0 9 9 1 11 2
4 3 13 9 3
3 1 11 11
8 1 12 13 11 10 0 9 2
28 15 13 9 9 2 7 15 4 3 10 9 2 15 13 15 13 2 16 15 4 4 0 1 9 13 0 9 2
12 15 4 0 9 2 16 11 11 13 1 9 2
16 2 7 3 13 10 0 9 1 10 12 9 2 2 13 15 2
10 12 9 3 13 0 9 9 1 11 2
7 1 0 9 1 12 9 2
20 7 10 9 4 11 11 3 13 15 0 1 14 4 13 10 9 3 1 9 2
22 15 4 3 9 1 7 15 1 9 1 10 0 9 2 15 4 13 9 1 11 9 2
7 12 13 15 1 0 9 2
7 15 13 1 10 9 9 2
5 3 13 15 12 2
9 7 15 13 3 1 10 0 9 2
16 12 2 1 13 9 13 3 3 10 0 9 1 9 1 11 2
8 15 4 0 14 13 0 9 2
9 15 13 2 16 9 4 13 15 2
13 12 2 4 9 13 1 10 7 9 9 1 9 2
15 12 2 15 4 0 2 16 15 4 13 1 9 9 9 2
18 12 2 16 15 4 13 1 9 9 2 3 4 15 3 3 13 3 2
21 12 2 7 13 3 3 0 9 1 9 2 16 15 4 13 9 1 9 1 9 2
29 12 2 16 3 13 10 0 9 2 4 15 3 4 0 1 2 16 15 3 3 13 3 7 13 1 0 9 9 2
13 9 4 3 13 10 9 2 11 11 2 13 9 2
24 2 15 13 2 0 2 2 7 15 4 0 2 16 9 9 7 9 3 4 4 13 1 9 2
46 15 4 3 0 2 15 9 13 1 9 1 10 0 9 2 16 15 4 13 14 13 10 9 2 7 16 15 4 9 1 10 0 9 1 2 15 11 13 7 13 2 2 13 11 11 2
13 2 13 4 3 0 13 2 15 13 3 10 9 2
49 16 15 3 4 13 1 9 2 4 9 4 13 0 2 7 3 4 3 12 0 9 3 4 13 3 3 2 7 15 12 1 9 4 4 13 10 9 2 2 13 11 7 11 2 3 1 9 9 2
25 15 12 13 1 10 0 9 2 15 1 9 4 13 3 2 16 9 7 9 13 14 13 0 9 2
43 3 1 9 1 15 12 13 13 3 1 9 2 13 15 3 1 9 1 2 16 3 4 9 9 3 1 10 9 3 1 10 9 2 1 4 4 3 0 1 10 0 9 2
24 11 7 11 4 0 1 14 13 3 1 0 9 2 16 15 4 3 3 0 1 14 13 15 2
22 7 1 0 15 4 9 15 15 2 2 15 4 3 4 10 0 2 15 4 13 2 2
14 7 9 1 10 9 13 9 1 14 13 1 10 9 2
21 15 4 3 13 9 1 0 9 7 11 0 9 14 13 1 10 9 1 0 9 2
10 15 4 13 9 2 13 11 11 11 2
17 2 9 4 4 0 1 2 16 15 3 4 13 9 3 10 9 2
14 13 9 3 1 9 2 13 15 3 2 2 13 9 2
14 10 0 9 13 3 10 10 0 9 2 13 1 9 2
4 15 13 9 2
6 3 1 11 0 9 2
4 12 13 3 9
10 12 9 4 3 13 9 14 4 9 2
8 10 0 4 13 2 13 9 2
16 3 13 11 2 16 12 9 1 9 13 3 1 10 0 9 2
11 3 13 10 0 9 12 0 9 1 9 2
9 1 14 13 13 9 3 1 12 2
7 15 13 10 9 1 9 2
8 9 4 13 1 10 13 9 2
3 11 11 11
7 10 0 0 9 13 11 2
7 3 13 11 15 1 11 9
35 9 11 11 13 3 10 0 9 1 9 1 12 1 9 1 2 16 3 4 13 9 1 10 10 2 0 0 9 2 9 2 9 7 9 2
18 2 15 13 1 14 13 9 1 9 1 9 1 9 1 10 10 9 2
31 10 0 9 4 13 1 2 16 10 0 9 13 2 16 3 13 10 0 9 7 9 1 9 2 2 13 11 11 1 11 2
35 9 4 1 9 2 15 13 1 9 1 9 2 13 12 9 2 15 13 0 1 9 1 9 1 9 1 12 9 1 9 3 1 12 9 2
23 11 11 13 3 2 16 10 9 1 9 7 9 4 4 3 1 14 13 10 3 0 9 2
2 13 9
31 2 15 13 3 13 1 2 16 9 7 9 4 13 9 1 0 9 2 15 15 4 13 9 7 9 2 2 13 11 11 2
3 13 12 9
27 9 13 1 13 0 9 1 9 1 11 7 11 2 7 9 3 13 9 2 11 2 11 2 11 7 11 2
43 10 12 9 1 9 4 13 12 9 1 9 1 9 2 7 15 13 3 12 9 1 9 10 0 9 2 3 9 13 3 3 2 11 2 11 2 11 2 11 12 7 11 2
17 15 3 4 13 1 9 13 9 3 9 1 1 9 10 0 9 2
21 3 4 15 3 4 13 16 9 4 13 2 16 3 1 9 1 0 9 13 8 2
10 4 15 9 13 9 9 10 0 9 2
22 1 3 14 13 3 0 1 9 2 16 9 1 9 3 4 13 9 1 11 9 9 2
20 4 10 9 1 9 1 9 3 13 14 13 9 8 13 12 9 3 1 9 2
16 3 10 12 3 13 9 1 9 13 1 9 1 10 0 9 2
7 9 13 1 3 12 9 2
13 9 13 3 7 3 1 13 7 0 9 1 9 2
29 2 15 13 14 13 1 10 9 7 13 2 13 15 13 15 1 10 0 9 2 2 13 10 0 9 2 11 11 2
17 1 9 4 15 13 1 9 2 15 13 15 1 9 1 10 9 2
15 10 9 1 9 7 9 13 13 9 1 10 9 1 9 2
9 2 15 13 9 3 1 10 9 2
11 15 13 3 1 9 2 2 13 11 11 2
24 10 10 9 2 2 15 13 14 13 1 0 2 3 0 16 15 4 9 2 9 7 9 2 2
23 12 0 9 4 13 1 9 2 16 15 4 13 10 13 9 2 15 4 13 3 1 9 2
6 3 4 10 9 13 2
36 10 13 9 1 9 11 1 11 13 2 16 0 9 1 9 4 13 14 13 0 9 1 0 9 1 14 13 15 1 14 13 3 1 13 9 2
11 9 12 0 9 13 10 0 9 1 11 2
18 9 12 13 10 0 9 9 1 9 1 14 13 9 7 13 9 3 2
8 9 12 4 11 10 0 9 2
6 2 9 4 3 0 2
5 9 13 3 13 2
13 10 0 9 13 1 9 2 2 13 9 1 11 2
7 2 15 4 4 10 9 2
14 15 4 0 2 16 9 3 4 13 2 16 9 13 2
17 3 3 15 4 13 1 9 2 4 9 3 13 13 7 3 0 2
16 15 4 13 1 2 16 9 4 13 1 10 0 9 1 11 2
17 16 11 13 2 4 15 3 4 13 10 0 1 9 1 9 2 2
3 9 4 0
13 9 12 2 0 9 2 13 9 3 3 1 11 2
10 10 0 9 1 9 2 9 7 9 2
6 2 9 4 13 3 2
6 9 13 3 1 9 2
7 15 4 10 0 9 3 2
24 9 13 10 0 9 1 9 2 2 13 11 11 2 11 11 7 9 1 11 2 9 11 11 2
15 1 10 9 13 10 0 9 9 1 9 1 14 4 0 2
22 10 0 9 4 10 9 9 3 13 2 16 9 4 13 9 1 9 1 9 7 9 2
27 15 13 10 9 13 11 9 2 15 4 13 15 3 13 1 9 2 1 14 13 9 13 1 3 0 9 2
6 7 15 4 3 0 2
11 10 0 9 13 9 2 1 9 2 3 2
5 11 9 1 9 2
12 2 11 4 3 0 1 9 1 10 0 9 2
17 15 13 15 2 16 9 13 3 3 2 16 15 4 13 15 15 2
14 15 4 4 13 3 2 1 15 13 2 7 4 0 2
14 15 13 14 13 1 9 2 7 10 9 4 0 2 2
17 15 4 0 2 16 9 13 14 13 9 3 7 13 1 10 9 2
22 2 15 13 3 1 10 9 7 13 2 16 15 4 3 0 2 9 4 13 9 2 2
12 2 9 13 2 16 10 0 9 13 1 9 2
46 16 15 13 9 1 14 13 2 13 15 2 16 11 9 4 2 13 2 15 1 10 9 2 15 1 10 9 3 4 4 13 1 10 9 2 15 15 3 4 4 13 3 1 9 2 2
28 1 9 1 10 0 1 9 0 0 9 4 11 11 0 1 14 13 2 16 9 3 3 13 14 13 3 3 2
12 2 15 4 13 9 1 11 3 1 0 9 2
28 7 3 1 15 1 9 13 1 9 2 16 15 4 4 13 10 9 3 2 13 15 3 10 0 9 1 9 2
25 16 11 11 13 3 7 13 15 3 1 0 7 15 9 9 2 4 3 0 2 7 3 3 0 2
19 15 4 0 1 2 16 0 9 1 15 4 4 13 9 10 0 9 2 2
2 11 11
14 0 4 13 3 1 11 9 11 11 1 9 1 11 2
4 9 2 11 11
39 1 0 9 2 1 9 1 9 12 7 12 10 0 9 12 2 4 11 11 3 1 9 4 13 10 9 7 13 15 3 1 9 1 14 13 15 1 9 2
23 2 3 4 9 3 13 3 2 2 13 11 9 1 10 13 9 1 11 9 9 1 9 2
12 2 9 1 9 12 13 11 11 3 13 2 2
36 9 11 11 13 15 15 1 9 2 7 1 9 4 15 1 9 13 3 1 2 15 3 4 13 15 3 7 13 2 2 3 4 0 9 2 2
16 3 2 16 3 4 13 10 9 2 15 1 10 9 1 11 2
53 13 1 9 13 9 11 11 2 11 9 2 15 3 1 9 11 11 11 13 9 10 0 9 12 1 11 11 1 10 9 1 9 1 10 9 2 3 2 16 15 4 4 13 15 1 2 16 15 13 11 1 9 2
30 2 10 9 4 13 10 9 3 1 15 2 2 13 10 0 9 1 9 2 7 15 13 1 10 9 1 10 0 9 2
13 9 4 3 3 13 2 7 13 1 10 0 9 2
42 9 2 15 4 13 12 2 4 13 7 13 1 11 9 1 10 0 9 1 2 16 9 4 9 7 10 0 9 1 14 13 1 10 3 2 3 3 7 3 0 2 2
3 1 13 9
23 9 1 9 13 1 9 1 11 9 9 1 0 2 11 2 7 13 15 3 1 10 9 2
14 9 13 2 16 3 1 12 0 4 13 7 13 9 2
30 10 0 2 15 3 4 10 9 2 13 3 1 12 7 0 9 3 1 9 2 15 13 1 9 7 10 0 10 9 2
22 1 14 13 9 13 10 9 10 0 9 1 9 2 16 9 13 1 10 9 1 9 2
29 15 4 3 13 0 9 1 9 1 10 0 9 3 1 11 7 11 2 3 0 9 3 13 3 1 9 1 9 2
36 11 13 9 1 11 1 9 2 7 15 13 2 16 9 9 3 3 10 0 9 13 13 1 9 12 1 12 2 7 1 10 9 1 9 12 2
1 0
34 9 2 15 3 3 4 4 13 15 7 15 0 1 9 2 16 15 13 2 13 1 0 9 2 3 9 9 1 0 9 13 12 9 2
30 0 9 12 9 7 11 11 9 1 0 9 1 11 9 1 9 12 9 2 1 3 4 9 1 0 1 9 10 9 2
1 9
18 0 11 9 1 9 1 16 9 4 0 13 12 9 2 9 12 9 2
8 9 1 0 9 13 12 9 2
17 15 13 0 9 1 9 3 2 3 8 9 1 0 1 0 9 2
16 7 3 13 10 9 9 14 13 1 15 1 9 9 1 11 2
22 0 9 4 11 11 4 13 1 10 9 2 16 9 13 1 11 1 14 13 1 9 2
22 7 3 13 9 3 9 2 1 15 16 11 13 15 9 7 10 0 9 1 0 9 2
17 3 1 16 15 3 4 13 2 3 1 14 13 10 3 0 9 2
13 7 9 13 14 13 1 9 1 9 3 1 9 2
3 13 10 9
23 2 15 13 3 15 2 15 13 2 16 9 13 10 9 2 9 7 13 9 1 10 9 2
27 3 1 14 13 10 0 9 7 13 9 1 0 9 2 13 15 3 10 0 9 9 2 16 15 13 0 2
4 15 13 9 2
10 7 15 4 3 0 2 3 0 2 2
29 11 11 13 10 10 0 9 1 8 9 9 2 2 1 10 9 13 15 10 0 9 2 3 3 4 0 1 9 2
13 2 13 9 2 4 15 3 0 2 2 13 15 2
30 15 13 9 3 2 15 13 10 10 9 2 7 15 13 15 1 9 7 13 2 2 13 9 2 15 13 10 9 2 2
22 15 4 4 12 9 2 16 15 13 10 9 1 10 0 9 1 9 2 11 11 2 2
16 10 9 4 11 11 11 2 13 0 9 12 1 9 9 11 2
75 7 3 13 15 3 10 0 9 1 12 2 3 15 13 10 11 1 2 11 11 2 2 7 9 1 3 11 11 2 11 11 2 11 2 11 11 2 11 11 2 11 11 11 7 11 11 9 11 11 4 3 3 3 13 15 1 9 7 13 3 7 3 1 2 16 11 11 11 13 1 9 3 1 12 2
20 11 11 11 9 1 10 9 1 9 7 3 1 9 4 4 10 0 1 0 2
32 11 11 13 10 3 2 0 9 2 1 11 11 7 9 11 11 7 11 11 1 11 11 4 13 3 7 3 1 1 12 9 2
13 7 15 0 13 2 15 13 9 3 3 1 9 2
14 0 9 4 13 2 13 2 13 7 13 1 15 9 2
7 15 4 10 9 7 9 2
5 10 0 15 4 2
11 1 9 13 3 3 1 10 0 9 9 2
14 9 13 15 1 13 9 2 16 9 13 9 1 15 2
24 3 13 15 15 1 14 13 3 0 9 2 13 9 7 13 9 1 9 1 14 13 1 9 2
27 15 13 3 1 3 3 3 10 0 1 2 13 1 16 9 3 4 13 0 9 1 9 1 1 0 9 2
29 3 13 10 0 9 1 10 0 9 1 10 0 10 0 9 2 7 9 13 3 3 3 14 13 1 10 0 9 2
8 15 4 10 0 9 1 9 2
20 15 15 4 3 15 2 15 3 13 1 2 3 10 7 10 9 1 0 9 2
18 15 4 3 0 9 1 15 9 14 13 2 16 9 3 13 10 9 2
8 7 13 15 13 10 0 9 2
12 0 9 13 3 1 14 13 3 2 13 9 2
26 2 3 13 7 13 9 4 13 9 1 10 0 9 1 9 7 9 1 9 2 2 13 11 11 11 2
45 1 9 7 9 1 9 2 15 13 3 1 9 1 9 7 9 1 2 10 0 9 1 9 2 15 13 3 1 14 13 3 10 0 9 1 10 3 0 2 3 0 7 0 2 2
12 2 15 4 13 10 0 9 1 9 7 9 2
42 10 9 2 3 9 13 15 1 9 1 14 13 3 0 9 2 16 15 3 13 1 9 1 3 14 13 2 15 3 1 9 4 9 7 9 1 9 2 2 13 11 2
10 3 13 3 0 1 0 9 1 9 2
40 15 13 10 0 9 2 2 9 1 11 13 1 10 9 2 15 1 10 13 9 1 10 9 2 10 9 7 10 9 4 13 0 9 7 13 0 9 1 9 2
9 11 11 11 4 3 10 0 9 2
9 7 11 11 2 6 6 6 2 2
36 1 1 10 9 9 1 9 7 0 9 4 10 0 0 11 3 3 3 3 1 10 9 2 11 11 2 12 2 7 9 2 11 7 11 11 2
28 11 13 3 3 9 14 13 3 1 10 9 2 16 11 9 1 10 9 3 13 2 16 15 4 13 1 9 2
10 1 9 13 11 9 3 7 3 9 2
12 2 15 13 2 7 11 9 13 9 1 11 2
24 15 4 3 0 2 15 3 3 13 11 7 13 15 1 0 9 2 2 13 11 11 2 12 2
30 1 0 9 13 9 3 12 9 1 11 9 2 1 14 4 4 13 1 9 1 14 13 2 3 9 4 13 1 9 2
11 7 12 0 9 1 0 9 13 3 9 2
19 7 9 13 10 0 1 11 3 3 10 9 1 10 3 13 9 1 11 2
30 1 9 1 11 11 0 9 1 11 4 9 1 9 13 9 3 1 10 0 9 2 1 9 1 11 4 13 3 1 2
17 15 4 3 13 1 0 9 1 9 1 14 4 4 13 1 9 2
11 15 13 15 2 15 13 1 10 0 9 2
37 15 13 2 9 13 15 3 2 16 15 3 13 14 13 10 9 2 15 3 3 13 0 0 9 1 10 9 2 7 3 13 14 13 3 3 3 2
28 15 4 13 10 0 9 1 3 9 2 9 2 9 2 9 7 9 2 16 15 4 3 13 1 10 0 9 2
32 4 15 0 1 2 16 15 3 3 4 10 0 9 15 13 2 7 1 3 3 3 0 9 9 7 9 2 9 7 9 2 2
3 13 3 3
11 2 10 9 4 3 0 1 9 1 15 2
45 13 3 3 15 13 1 2 15 4 3 3 13 1 14 13 9 1 9 1 15 2 15 3 4 13 15 10 8 0 9 2 3 9 1 15 2 2 13 9 2 15 13 9 3 2
7 2 11 11 4 10 9 2
30 15 4 0 7 0 2 7 16 15 4 9 2 7 15 4 11 11 1 9 2 13 1 9 1 10 11 7 10 11 2
12 15 13 0 9 2 7 9 13 1 0 9 2
11 15 4 3 13 11 7 4 3 13 15 2
17 15 4 3 13 0 9 1 0 2 7 9 13 3 1 9 9 2
25 15 13 3 0 0 9 3 13 1 14 13 9 1 10 0 9 2 2 13 9 9 2 11 11 2
42 1 10 9 2 3 11 13 14 13 2 4 11 11 3 13 1 11 2 2 3 4 15 13 15 1 10 0 9 1 2 16 15 3 13 1 9 1 10 0 0 9 2
2 0 9
11 7 9 11 11 11 4 3 4 10 9 2
10 15 13 0 9 2 4 0 7 0 2
26 15 4 4 10 0 9 1 10 13 0 9 2 15 3 4 13 10 3 0 9 2 2 13 11 11 2
20 3 1 9 13 3 9 2 7 3 13 11 1 9 1 12 9 1 12 9 2
13 1 9 13 11 1 11 11 7 11 11 1 12 2
21 3 13 11 2 11 2 11 2 11 7 13 3 1 9 12 2 11 2 1 11 2
14 10 0 4 11 2 11 2 11 7 11 1 11 11 2
35 15 4 3 13 2 16 11 1 11 11 4 13 10 9 2 3 11 4 13 3 3 1 10 13 9 2 7 9 13 9 7 13 3 9 2
4 0 13 9 2
17 11 13 9 1 12 9 2 7 11 11 13 1 3 12 9 9 2
3 10 0 9
10 9 13 9 1 2 16 15 13 9 2
19 15 13 9 1 14 13 15 1 9 1 10 0 9 3 12 9 1 9 2
18 3 13 11 11 9 2 16 15 13 7 13 3 11 11 7 11 3 2
26 1 9 4 15 4 13 3 1 9 1 15 2 16 15 4 9 2 0 9 7 9 2 15 15 3 2
27 15 4 3 4 3 0 2 16 15 4 13 2 16 9 13 0 9 2 13 15 1 9 1 10 0 9 2
40 16 15 4 13 14 13 15 15 7 15 2 1 9 2 15 3 13 9 1 9 2 9 2 0 9 2 9 2 2 9 2 7 2 15 13 2 15 13 2 2
11 7 15 1 15 4 0 9 0 9 3 2
22 15 13 0 3 9 1 3 14 13 3 7 13 2 16 15 4 13 14 4 0 9 2
32 3 4 3 13 1 9 7 9 2 1 14 13 9 1 14 13 2 10 0 2 3 7 13 15 1 10 0 9 1 10 9 2
5 15 4 3 0 2
34 9 4 1 3 4 3 1 14 13 7 13 1 9 1 10 0 9 1 10 0 9 2 7 0 9 1 16 15 13 3 7 3 13 2
7 2 15 4 10 0 9 2
7 7 15 13 3 3 2 2
15 9 1 11 4 11 11 2 1 3 4 9 1 11 11 2
20 15 4 4 3 1 3 1 11 14 13 2 16 3 11 7 11 4 0 9 2
28 11 0 9 13 1 9 2 11 4 1 9 9 13 11 9 9 2 11 2 1 14 13 15 1 9 1 9 2
10 9 11 11 2 2 15 13 3 3 2
29 7 15 13 3 2 16 15 4 10 0 9 14 13 3 1 9 1 2 7 15 13 3 3 9 3 1 9 2 2
9 15 13 12 9 14 13 10 9 2
19 9 2 15 9 3 13 2 13 2 16 11 1 9 4 13 15 1 11 2
21 10 0 9 13 3 2 3 11 13 3 7 13 1 11 2 16 11 3 13 9 2
22 3 13 11 1 9 1 11 2 3 15 4 13 2 16 3 13 11 1 9 1 11 2
14 3 4 15 13 1 9 2 16 15 3 13 1 9 2
10 7 16 0 4 0 2 13 9 3 2
13 9 1 0 9 1 11 7 11 4 3 3 0 2
49 3 4 3 13 10 0 0 9 3 1 9 1 9 1 12 2 7 1 12 13 15 9 0 9 2 0 9 11 11 2 9 1 10 9 9 2 16 15 3 13 3 1 10 9 1 10 12 9 2
22 3 4 9 3 0 1 10 3 0 9 2 2 15 4 15 1 3 3 3 3 3 2
25 15 13 1 10 9 3 1 10 0 2 0 9 2 3 10 12 9 9 4 13 15 9 14 13 2
13 3 4 0 0 9 7 9 4 10 9 1 9 2
10 15 4 13 0 9 1 10 12 9 2
13 15 4 13 1 9 1 10 13 9 1 0 9 2
21 10 0 4 3 13 1 9 2 16 10 9 4 13 9 1 9 2 2 13 9 2
16 1 10 9 1 9 1 11 4 15 9 13 1 11 1 9 2
17 2 15 13 3 3 2 16 3 13 10 9 2 15 4 13 9 2
27 3 13 15 9 1 9 7 13 13 9 1 9 2 15 4 13 11 9 1 11 9 2 2 13 11 11 2
27 15 13 3 1 11 9 1 10 9 2 15 1 9 1 9 13 0 9 14 13 0 1 12 9 1 9 2
13 9 13 10 9 3 3 2 15 13 1 12 9 2
17 13 3 12 9 2 4 9 13 1 0 9 1 4 15 0 9 2
8 7 3 13 9 1 0 9 2
8 9 4 13 1 9 1 9 2
12 7 9 13 3 9 1 15 1 1 0 9 2
18 11 13 1 10 0 9 1 10 0 9 1 9 2 15 13 1 9 2
27 11 11 2 3 4 13 9 7 13 10 9 1 9 2 4 13 9 3 1 11 11 11 1 9 1 11 2
20 11 2 15 4 15 9 2 12 9 0 7 1 13 9 1 2 0 9 2 2
13 7 15 4 3 10 9 0 9 2 9 7 9 2
14 7 3 4 15 1 3 12 1 11 9 3 0 9 2
18 3 4 15 13 9 7 11 1 9 1 11 11 9 2 9 9 2 2
16 11 11 7 11 11 13 1 10 9 1 14 13 10 0 9 2
22 15 4 4 13 1 14 13 1 9 7 13 14 13 2 3 15 13 16 15 4 9 2
16 7 16 15 13 1 9 2 3 4 15 13 15 3 1 9 2
21 2 6 2 7 15 4 3 13 15 16 15 4 12 9 0 2 2 13 11 11 2
11 2 3 13 15 1 0 9 1 11 9 2
14 15 13 0 9 3 1 10 9 2 2 13 11 11 2
2 0 9
26 2 15 13 16 2 15 13 10 0 9 3 2 2 13 11 7 13 1 9 2 15 4 3 4 0 2
25 11 11 4 12 7 3 1 10 0 9 3 0 1 10 9 1 0 9 2 15 13 15 9 1 2
33 15 4 3 3 0 1 9 2 11 9 4 3 13 0 9 1 9 2 9 2 3 9 2 2 15 1 9 13 1 10 0 9 2
10 3 13 15 10 9 3 3 1 12 2
14 7 9 4 3 2 15 15 4 13 2 0 7 0 2
9 1 9 1 15 13 1 10 9 2
33 2 15 4 3 3 9 2 7 15 13 2 16 9 3 1 9 13 1 9 1 14 13 10 9 2 1 0 9 4 9 13 2 2
9 16 11 13 9 2 4 10 9 2
25 15 4 13 1 12 0 9 1 9 2 3 11 2 3 3 12 1 12 9 13 1 0 1 9 2
25 7 16 15 4 15 2 13 15 3 3 2 16 9 13 15 1 9 1 3 14 4 13 1 9 2
41 2 16 9 3 13 2 3 4 15 13 15 2 2 13 11 11 1 9 1 2 16 9 11 11 11 2 11 2 4 13 14 13 15 15 2 16 9 4 13 9 2
47 3 13 15 3 13 11 0 9 2 11 11 1 9 2 16 9 1 10 0 9 1 9 13 1 9 2 16 2 15 4 3 1 10 9 14 13 2 16 3 4 13 9 1 11 9 2 2
28 11 11 4 1 9 13 9 13 2 16 9 11 4 13 9 2 9 7 9 1 9 1 9 9 1 11 9 2
2 0 9
38 16 11 1 12 9 3 13 0 1 10 9 1 12 9 9 2 4 3 3 13 10 9 1 0 13 9 1 11 9 14 13 0 9 1 4 13 3 2
15 10 0 9 1 11 12 9 7 12 9 4 13 1 9 2
27 12 13 1 9 13 10 9 2 7 0 9 2 0 9 2 9 2 10 9 7 9 13 0 9 1 9 2
24 1 9 13 15 12 13 2 16 9 3 13 1 14 13 2 16 15 13 1 9 1 10 9 2
11 15 13 15 2 15 13 1 2 9 2 2
19 9 12 0 9 13 15 3 2 2 15 13 1 2 16 15 13 10 9 2
12 15 4 10 0 9 2 2 13 2 9 2 2
27 7 1 10 0 9 1 9 9 4 15 0 1 2 16 10 0 4 13 10 9 7 13 10 0 9 3 2
17 2 13 15 9 1 2 16 9 13 13 2 2 13 9 11 11 2
8 9 2 2 3 13 15 15 2
15 15 4 3 3 13 1 15 2 16 3 13 15 1 9 2
23 3 4 10 9 3 13 9 2 7 15 13 3 15 2 16 15 13 1 9 1 11 2 2
24 2 9 2 2 2 15 4 13 1 10 10 9 2 16 15 4 13 1 10 9 1 11 2 2
22 16 9 13 1 11 2 13 9 3 1 10 9 1 2 9 2 1 15 1 10 9 2
17 15 4 13 3 1 10 9 1 14 13 15 2 16 15 4 0 2
