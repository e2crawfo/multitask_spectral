13304 11
11 10 11 1 3 0 9 1 1 12 13 2
7 15 9 11 1 13 4 2
7 15 9 9 12 0 13 2
17 15 12 9 13 7 0 9 9 1 13 1 1 12 9 9 13 2
6 0 9 3 0 13 2
16 15 13 1 12 9 1 9 0 9 1 9 1 0 13 4 2
28 11 11 1 1 0 9 1 9 0 9 1 10 0 9 11 11 1 9 1 13 15 11 11 14 13 4 4 2
10 15 9 7 9 9 1 0 9 13 2
8 15 11 1 0 0 9 13 2
13 0 9 1 15 9 9 7 9 9 1 9 13 2
8 15 9 11 1 9 13 4 2
20 0 9 1 13 10 9 1 9 2 1 1 0 9 15 10 14 0 13 4 2
39 15 1 12 9 9 2 9 9 2 9 9 1 1 9 2 12 9 2 0 7 0 9 2 9 9 2 0 9 1 9 2 0 7 0 9 9 14 13 2
18 15 11 1 1 0 9 9 12 9 1 9 12 9 1 13 4 4 2
19 15 12 0 9 13 15 12 9 1 11 11 1 0 9 1 1 13 4 2
26 15 12 0 9 1 13 7 9 1 15 9 1 12 14 9 13 15 0 9 1 0 9 1 1 13 2
16 7 10 9 1 15 9 7 9 1 0 9 1 13 4 4 2
18 15 9 2 9 9 2 9 7 11 1 9 1 9 14 13 4 4 2
20 15 9 1 9 2 0 2 0 9 2 0 9 7 0 9 1 13 4 4 2
17 15 11 11 1 0 9 1 9 1 0 9 0 13 13 4 4 2
7 9 11 1 0 13 4 2
7 15 11 11 1 0 13 2
26 15 13 4 12 9 13 15 11 1 11 2 11 2 11 7 11 9 1 0 9 9 1 13 4 4 2
18 10 9 14 11 1 13 0 9 12 9 1 12 9 1 13 4 4 2
12 0 9 1 13 9 1 10 9 9 0 13 2
7 15 12 9 1 13 4 2
20 0 9 1 1 15 0 9 1 0 7 0 9 1 13 1 9 13 4 4 2
21 15 11 1 13 10 9 9 12 1 12 7 12 1 12 9 9 1 13 4 4 2
17 15 0 9 1 9 9 13 15 11 11 1 9 1 1 0 13 2
16 15 9 7 9 9 9 13 7 12 11 9 1 9 14 13 2
15 15 11 1 13 10 9 9 12 1 12 1 13 4 4 2
16 9 1 1 0 11 1 0 9 2 9 9 1 9 13 4 2
14 0 9 1 0 9 13 15 9 1 9 13 4 4 2
24 15 15 9 1 9 2 9 2 9 1 9 7 9 1 9 0 9 1 13 7 13 4 4 2
12 11 11 11 11 1 12 9 1 0 13 4 2
12 11 11 11 11 11 11 1 9 14 13 4 2
11 11 11 1 12 9 1 9 1 9 13 2
3 15 13 2
15 11 11 2 11 7 11 1 11 1 1 0 9 9 13 2
10 11 2 11 2 11 9 9 1 13 2
17 11 1 11 7 11 1 9 11 13 1 0 9 11 13 13 4 2
26 11 7 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 1 1 0 9 9 13 2
15 13 1 1 2 11 11 11 11 1 9 7 0 9 13 2
3 15 13 2
10 9 1 15 14 15 15 13 4 4 2
32 11 1 9 9 1 14 9 13 4 4 2 9 15 13 4 13 4 7 15 13 4 4 9 9 1 2 11 1 12 9 1 2
17 15 1 9 7 9 1 9 1 9 1 9 14 13 14 4 4 2
19 11 1 11 11 1 11 9 1 13 4 10 9 0 9 1 9 13 4 2
15 11 2 11 11 1 11 9 11 11 1 1 13 4 4 2
18 15 1 1 9 1 0 9 7 9 13 15 9 1 12 9 13 4 2
10 15 9 11 11 11 1 9 0 13 2
14 9 7 9 1 11 9 1 0 9 13 14 13 4 2
18 11 11 7 9 1 9 7 9 1 9 15 1 9 1 9 13 4 2
19 10 9 9 11 11 11 1 11 11 1 11 1 11 13 1 3 13 4 2
25 15 0 9 1 1 9 1 13 4 9 9 1 9 13 4 7 15 0 9 3 0 9 13 4 2
15 9 1 9 1 10 9 11 11 1 11 11 1 13 4 2
13 3 9 1 13 4 0 9 1 0 9 9 13 2
14 15 12 0 9 11 9 7 11 9 1 1 13 4 2
14 3 15 9 11 11 1 0 9 1 1 1 13 4 2
20 15 0 9 2 3 13 4 9 7 0 9 0 9 1 9 1 9 13 4 2
12 9 1 1 15 11 11 1 13 3 0 13 2
13 15 9 1 1 9 9 1 1 1 13 4 4 2
20 15 9 2 1 1 9 10 13 4 14 13 15 1 15 11 11 13 4 4 2
13 11 9 1 9 1 0 9 15 13 1 13 4 2
9 15 1 0 9 9 13 4 4 2
18 10 9 1 1 10 0 2 0 9 13 15 15 9 1 9 13 4 2
8 15 0 9 1 0 9 13 2
21 15 9 1 0 13 11 1 11 11 13 1 3 15 12 0 9 1 15 13 4 2
11 9 1 9 9 7 9 1 13 4 4 2
13 15 11 1 9 1 9 13 1 1 13 4 4 2
12 15 15 12 0 9 1 1 1 13 4 4 2
12 15 1 0 11 1 0 9 13 4 4 4 2
15 15 9 1 1 0 9 1 9 13 1 1 13 4 4 2
24 10 0 9 1 11 11 1 9 7 11 1 9 1 13 4 11 9 1 9 13 4 4 4 2
29 13 4 4 16 9 1 9 11 9 1 1 9 2 9 9 13 1 9 1 1 11 11 1 10 0 9 13 4 2
16 15 11 1 9 13 15 13 1 1 3 9 13 13 4 4 2
13 10 9 1 9 1 9 1 9 14 13 4 4 2
16 3 9 1 13 9 1 12 9 3 11 1 9 13 13 4 2
21 9 1 1 0 10 9 1 9 11 11 11 1 11 1 0 9 1 1 13 4 2
13 15 9 1 11 0 9 1 9 13 4 4 4 2
30 11 11 2 11 11 11 11 2 11 11 11 2 11 11 11 11 11 11 2 11 11 11 11 7 11 11 14 0 13 2
12 15 9 9 1 9 1 9 13 14 4 4 2
14 11 9 7 15 1 0 9 9 14 9 1 13 4 2
2 15 13
19 12 9 1 11 11 11 15 1 13 15 11 2 11 7 11 1 13 4 2
21 11 2 11 2 11 2 11 7 11 1 0 9 9 1 15 1 13 4 4 4 2
23 11 11 11 2 12 9 2 11 2 11 0 9 1 13 7 11 12 9 1 9 1 13 2
3 15 13 2
14 11 1 13 11 1 1 9 15 13 1 1 0 13 2
10 10 9 15 9 1 9 13 4 4 2
28 0 9 1 3 9 1 0 0 11 11 13 15 13 1 1 12 9 1 9 1 12 9 1 9 13 4 4 2
31 10 9 13 4 7 10 14 9 7 9 1 9 7 9 1 9 13 11 11 9 1 9 1 12 9 0 9 1 13 4 2
18 15 9 1 12 9 9 1 0 9 13 15 11 11 11 11 13 4 2
24 15 9 1 1 9 2 9 2 9 2 9 2 0 9 7 10 9 1 9 0 9 1 13 2
14 9 7 9 1 13 1 1 11 1 12 14 9 13 2
11 10 9 1 9 11 11 1 13 4 4 2
28 9 1 1 9 2 9 2 0 9 2 9 2 9 9 2 9 7 9 1 9 1 14 9 13 4 4 4 2
22 15 1 11 9 9 14 9 1 9 1 9 13 15 9 11 11 11 1 9 13 4 2
9 9 0 9 1 9 14 13 4 2
15 11 11 1 11 11 1 9 11 1 15 1 9 13 4 2
14 3 1 15 9 11 1 9 1 13 9 1 0 13 2
11 11 11 1 11 0 9 11 15 0 13 2
16 11 11 1 11 11 1 12 9 9 13 15 13 1 9 13 2
12 3 1 12 9 1 9 13 11 1 15 13 2
12 11 1 9 1 1 9 1 9 0 13 4 2
12 0 9 1 9 1 0 9 1 0 13 4 2
11 11 1 9 1 11 11 1 15 9 13 2
11 11 11 1 15 13 15 9 1 0 13 2
21 11 11 1 13 1 1 9 1 15 10 9 9 13 15 10 9 11 11 0 13 2
12 15 9 1 1 10 9 9 1 1 13 4 2
20 9 9 11 11 1 11 1 11 1 9 11 11 11 1 10 9 9 1 13 2
12 15 1 15 9 1 9 1 1 0 13 4 2
14 9 1 14 15 11 11 2 11 11 7 11 11 13 2
24 11 11 1 1 7 9 1 9 1 11 11 13 4 4 2 15 15 9 9 1 9 9 13 2
8 15 0 9 1 9 14 13 2
22 9 11 11 7 11 1 9 1 1 0 11 11 11 14 9 1 9 13 13 4 4 2
10 11 11 11 1 14 12 9 1 13 2
17 11 11 11 11 1 13 1 1 12 13 9 7 12 9 0 13 2
17 11 11 1 1 12 9 1 1 9 1 1 10 9 0 13 4 2
18 9 1 14 12 9 1 9 10 9 1 12 9 1 0 13 4 4 2
32 0 12 9 1 10 9 1 9 13 4 11 11 11 1 13 16 9 1 9 3 13 4 4 2 7 9 3 3 14 13 4 2
10 9 1 9 9 1 14 12 9 13 2
11 9 14 0 9 1 9 13 9 13 4 2
11 10 9 11 11 7 11 11 1 13 4 2
15 10 9 9 1 12 9 9 1 0 9 1 13 4 4 2
20 14 3 0 3 0 9 13 15 0 9 7 0 9 1 9 1 13 4 4 2
18 3 14 15 11 11 1 9 1 10 0 9 1 10 0 9 13 4 2
16 15 13 1 3 15 9 14 10 0 9 1 13 1 13 4 2
18 15 10 9 1 15 15 1 9 13 4 4 11 1 10 0 9 1 2
10 10 9 1 9 13 4 11 11 1 2
11 11 11 1 11 1 0 9 13 4 4 2
20 0 9 1 0 10 9 1 15 11 1 9 7 9 12 1 9 13 4 4 2
26 16 15 1 10 14 9 7 9 13 16 9 1 1 15 1 9 1 9 2 9 13 3 0 13 4 2
17 16 0 14 13 4 16 15 1 12 9 3 9 1 1 13 4 2
7 14 13 15 9 13 4 2
11 7 9 1 1 1 0 11 1 9 13 2
10 11 0 9 2 9 2 1 9 13 2
22 10 9 15 9 0 9 2 9 1 0 9 7 9 13 1 9 1 9 1 13 4 2
12 0 9 1 10 9 1 9 14 10 0 13 2
10 0 9 1 1 15 9 1 13 4 2
19 16 15 0 9 2 0 9 7 0 9 1 0 13 16 11 15 9 13 2
22 10 9 1 0 9 15 13 16 15 1 0 9 15 1 9 1 9 1 13 4 4 2
13 15 15 1 0 9 1 9 1 9 14 13 4 2
11 7 9 14 10 9 1 10 0 14 13 2
29 16 15 9 2 9 1 1 9 1 9 1 0 9 1 13 13 4 16 11 1 1 15 13 1 1 10 15 13 2
11 3 14 11 11 11 1 1 12 9 13 2
7 7 15 1 15 9 13 2
22 7 16 7 15 1 9 1 9 7 15 1 13 9 14 11 1 9 1 10 0 13 2
24 15 13 7 9 1 9 13 1 9 13 4 16 15 1 9 11 11 1 10 14 0 13 4 2
12 0 9 1 10 9 1 3 0 9 9 13 2
11 15 9 1 0 11 9 1 13 4 4 2
17 11 9 1 1 9 13 1 11 1 9 1 0 12 11 9 13 2
12 15 11 13 14 14 4 16 13 14 4 4 2
19 16 15 14 0 9 7 9 1 9 13 13 4 16 11 1 9 3 13 2
1 11
14 15 1 9 2 9 10 9 0 9 1 13 4 4 2
20 15 1 9 1 13 4 15 0 13 0 9 1 0 9 9 1 1 0 13 2
20 10 0 2 0 2 0 9 1 15 1 13 4 15 9 1 9 1 13 4 2
15 16 9 1 15 1 9 9 9 1 1 14 9 13 4 2
10 9 1 15 1 9 3 0 13 4 2
23 10 9 1 0 9 1 15 0 9 11 1 9 7 2 9 9 2 1 9 13 9 13 2
10 11 15 1 9 1 9 1 13 4 2
12 11 13 1 3 0 9 1 9 13 14 13 2
24 15 9 1 9 1 9 12 9 0 13 4 15 1 15 11 13 1 1 9 3 10 13 4 2
19 12 9 0 11 11 1 0 9 1 11 1 13 1 9 14 10 0 13 2
11 9 1 0 9 1 12 9 13 4 4 2
12 11 11 1 13 1 1 0 9 1 9 13 2
13 10 9 1 13 1 1 15 0 9 1 13 4 2
13 7 9 1 1 13 1 3 15 10 9 0 13 2
10 7 15 11 1 9 1 0 9 13 2
14 11 13 16 15 15 14 13 16 15 15 14 14 13 2
9 15 14 11 9 1 14 9 13 2
8 7 11 11 11 15 0 13 2
18 9 3 15 12 0 9 13 15 3 1 9 1 9 13 4 4 4 2
32 10 9 1 15 11 1 9 2 11 11 11 2 11 1 9 1 0 9 2 11 1 9 1 13 10 0 9 1 13 4 4 2
18 15 1 12 0 9 1 0 2 0 7 0 9 1 0 9 13 4 2
17 10 9 10 0 7 0 13 16 15 13 1 1 12 9 10 13 2
18 10 9 1 0 9 1 9 1 1 1 12 3 0 9 13 4 4 2
10 9 1 13 4 9 13 14 13 4 2
16 16 15 11 13 13 16 11 9 1 9 13 1 9 3 13 2
23 15 9 13 4 15 9 1 0 9 1 1 2 9 11 1 9 1 14 9 13 4 4 2
21 15 1 14 11 9 1 9 1 9 13 4 0 9 1 3 13 3 0 9 13 2
13 9 1 10 9 1 9 1 1 0 9 13 11 2
11 15 13 13 4 16 9 0 13 4 4 2
16 15 9 1 1 2 9 15 9 1 0 9 9 14 13 4 2
14 3 0 3 15 9 9 1 9 1 14 3 13 4 2
51 0 9 1 13 0 9 13 9 2 0 2 0 9 2 0 9 7 12 9 1 0 9 1 3 9 13 4 10 9 13 14 0 13 4 2 7 11 1 11 9 1 9 1 1 15 15 0 9 14 13 2
24 15 9 1 1 15 10 9 1 1 9 1 0 13 4 9 1 3 1 10 0 13 4 4 2
16 9 15 15 9 13 4 4 2 11 1 0 9 9 11 1 2
19 11 1 9 14 12 12 13 2 7 15 10 9 14 12 12 9 13 4 2
15 9 1 0 9 1 10 9 1 9 1 9 13 4 4 2
12 9 1 9 1 15 11 1 0 0 9 13 2
11 11 1 9 9 1 9 14 13 4 4 2
8 15 1 9 9 10 0 13 2
16 9 1 0 9 13 14 15 1 9 7 9 0 13 4 4 2
14 15 1 0 9 9 10 9 1 12 9 13 4 4 2
9 11 1 3 2 3 9 13 4 2
23 10 9 1 9 13 11 1 12 0 9 1 9 13 4 7 15 9 13 4 2 11 11 2
15 15 1 0 9 9 1 13 10 9 15 1 9 13 4 2
16 9 1 13 14 0 13 4 4 16 15 10 9 15 13 4 2
9 9 1 0 9 0 13 4 4 2
18 15 10 9 1 0 9 1 13 14 13 4 2 7 14 3 13 9 2
9 9 1 1 15 1 10 15 13 2
13 9 1 10 9 1 15 10 9 9 1 13 4 2
20 15 12 0 9 1 15 9 7 9 1 1 13 1 9 1 0 13 4 4 2
11 9 1 1 15 0 0 9 1 9 13 2
10 15 9 7 9 9 0 9 9 13 2
25 10 9 9 1 3 0 9 13 16 15 15 9 1 1 13 0 9 1 9 1 9 13 4 4 2
18 15 15 11 11 11 1 0 0 9 1 9 11 1 3 13 4 4 2
10 15 10 9 0 9 1 13 4 4 2
25 3 11 12 9 9 13 2 7 15 15 12 9 1 9 13 0 9 1 1 0 9 13 4 4 2
12 11 1 9 1 9 13 4 16 0 14 13 2
15 15 9 1 1 10 15 13 2 15 1 12 13 11 11 2
13 15 13 9 9 1 0 2 0 9 1 3 13 2
24 15 15 11 1 9 1 14 3 13 4 4 2 15 11 1 9 1 13 1 15 9 1 13 2
20 15 1 11 11 1 2 11 11 11 2 0 12 9 1 0 9 13 4 4 2
20 10 9 1 11 1 0 9 7 9 9 1 9 1 13 0 9 13 4 4 2
17 15 1 15 10 9 13 1 9 9 9 9 1 10 0 13 4 2
14 10 9 1 10 9 1 0 9 1 9 13 4 4 2
16 10 0 7 0 13 16 11 11 1 11 11 15 0 9 13 2
8 15 10 0 0 9 9 13 2
13 9 7 9 9 1 9 13 9 9 13 4 4 2
13 15 13 15 13 16 15 9 9 1 13 4 4 2
19 11 1 14 12 9 1 9 1 0 13 2 11 1 0 0 11 11 11 2
18 11 1 11 11 7 11 11 1 9 9 1 11 11 11 13 4 4 2
13 10 9 11 11 1 1 0 9 1 9 13 4 2
3 15 13 2
13 11 13 1 1 11 2 11 1 9 3 0 13 2
7 9 15 1 0 9 13 2
12 10 9 9 1 9 10 9 1 13 4 4 2
11 11 11 1 9 15 11 11 13 4 4 2
24 10 9 15 15 0 11 1 11 1 9 1 3 0 0 2 0 7 0 9 1 13 4 4 2
3 15 13 2
14 15 11 1 1 11 7 11 1 0 9 13 4 4 2
12 10 9 1 0 9 1 0 9 13 4 4 2
21 15 1 11 11 11 7 11 11 11 9 2 9 1 14 12 9 1 13 4 4 2
24 15 1 9 1 9 2 9 7 9 1 0 9 13 2 15 15 15 9 1 1 13 4 4 2
3 15 13 2
12 9 1 9 1 11 11 1 0 0 9 13 2
13 15 0 9 9 1 1 0 0 9 9 9 13 2
15 15 15 13 1 3 9 1 9 9 13 4 16 0 13 2
11 16 15 9 0 13 16 10 3 9 13 2
10 0 9 1 9 10 0 13 4 4 2
15 15 1 14 11 1 9 1 13 1 9 14 3 0 13 2
13 16 15 15 9 1 8 13 4 16 15 3 13 2
19 11 2 15 11 14 13 4 4 2 9 2 9 7 0 9 1 9 13 2
13 15 1 3 0 9 15 1 9 1 9 9 13 2
17 15 12 1 12 9 1 9 1 15 1 9 11 1 13 4 4 2
13 15 13 15 9 3 14 9 13 1 1 13 4 2
6 15 11 1 9 13 2
10 15 9 1 3 0 9 1 0 13 2
9 10 9 10 0 9 1 13 4 2
12 16 15 15 13 16 9 1 9 13 14 13 2
16 10 0 9 1 15 9 1 1 9 1 9 12 0 9 13 2
15 15 9 1 11 11 11 0 9 1 1 13 4 4 4 2
10 15 1 9 7 9 13 14 13 4 2
12 15 11 1 3 0 9 2 11 11 2 13 2
14 15 15 0 9 1 13 0 0 9 1 13 4 4 2
9 11 1 9 1 0 9 9 13 2
10 15 9 9 1 9 1 9 0 13 2
15 10 9 1 9 1 0 13 1 1 9 9 13 4 4 2
11 15 9 0 0 13 9 1 0 13 4 2
17 10 9 1 12 9 0 13 1 1 1 15 0 9 13 4 4 2
19 15 1 14 15 10 0 9 13 2 15 15 0 9 1 0 9 13 4 2
11 10 9 11 1 0 9 1 10 0 13 2
15 10 0 9 1 13 1 1 15 11 1 9 13 4 4 2
21 11 0 9 13 2 15 1 15 12 9 9 1 13 11 1 0 9 13 4 4 2
5 15 10 9 13 2
8 15 1 11 11 10 0 13 2
14 11 11 1 15 9 1 0 2 0 9 13 4 4 2
14 10 9 1 0 9 1 13 10 9 13 13 4 4 2
14 9 13 1 3 14 11 11 11 1 9 13 14 13 2
13 11 1 1 15 12 9 1 0 11 13 4 4 2
25 10 9 1 13 15 3 2 11 2 9 1 9 2 13 12 9 16 9 13 2 1 9 13 4 2
18 11 1 9 1 3 1 13 9 1 9 1 0 9 13 14 13 4 2
8 15 11 1 9 13 4 4 2
14 3 14 11 9 1 3 0 9 9 7 9 9 13 2
16 16 15 10 9 1 9 13 4 16 11 11 1 9 3 13 2
12 15 0 9 1 0 9 1 1 13 4 4 2
17 15 1 9 9 1 9 1 8 13 1 1 15 0 9 13 4 2
11 11 1 1 13 0 9 14 13 1 13 2
12 9 9 1 1 10 9 14 12 9 0 13 2
16 10 9 1 9 11 11 1 1 11 11 11 1 1 13 4 2
15 9 1 1 10 9 1 0 2 0 9 1 9 13 4 2
13 15 1 11 2 11 7 11 11 1 9 0 13 2
9 9 9 1 9 9 14 0 13 2
13 7 15 1 0 9 1 9 1 10 9 9 13 2
3 15 13 2
12 11 13 1 0 9 11 1 11 9 1 13 2
12 3 9 1 9 1 9 9 10 0 13 4 2
17 9 1 1 9 1 11 11 1 11 11 1 0 13 4 4 4 2
3 15 13 2
14 15 9 2 9 7 9 9 2 15 3 13 4 4 2
8 15 1 3 0 9 11 13 2
15 7 15 11 7 11 1 15 1 1 0 9 13 4 4 2
26 15 1 15 11 2 11 2 11 7 9 1 15 14 9 1 15 1 1 9 7 9 9 13 4 4 2
3 15 13 2
19 15 9 1 9 1 12 1 12 12 9 1 0 0 7 0 9 0 13 2
16 9 1 1 13 10 0 0 0 9 1 13 12 0 9 13 2
17 7 16 15 9 10 13 16 9 1 1 0 9 7 9 14 13 2
16 15 15 12 12 1 1 12 12 9 1 0 9 13 4 4 2
26 9 10 9 1 0 13 4 16 15 9 1 10 9 1 9 13 4 4 7 15 11 1 15 1 13 2
16 10 9 13 16 11 1 11 11 1 9 1 14 13 4 4 2
23 9 10 0 9 1 13 4 16 9 15 0 13 4 9 1 10 0 9 1 13 4 4 2
19 13 4 4 16 11 1 9 0 9 2 11 11 1 11 11 1 13 4 2
13 15 1 11 1 0 9 9 9 1 0 9 13 2
22 11 1 0 9 1 9 13 10 9 1 9 11 9 1 9 11 1 11 1 13 4 2
13 11 9 1 13 10 0 9 1 12 9 13 4 2
26 9 1 12 9 9 13 2 15 11 11 2 11 11 2 11 11 7 11 11 1 9 1 13 4 4 2
10 10 9 0 9 9 1 0 9 13 2
16 0 9 1 0 7 0 9 1 9 1 9 1 13 4 4 2
7 11 1 10 10 9 13 2
23 15 1 15 12 9 1 10 0 13 2 7 10 0 13 1 3 14 15 9 13 1 13 2
16 10 9 1 9 15 0 9 2 9 2 9 7 0 9 13 2
6 15 9 1 13 4 9
20 10 9 1 9 14 1 9 2 11 11 1 9 7 11 1 9 13 1 13 2
15 9 1 9 1 0 0 9 9 1 9 1 0 13 4 2
14 11 11 1 9 1 11 1 11 11 11 1 13 4 2
29 14 12 9 0 10 9 1 0 0 9 7 9 13 4 9 1 9 1 9 1 13 9 9 1 9 13 4 4 2
22 3 11 1 9 1 0 9 9 1 13 4 16 3 0 9 1 0 9 13 4 4 2
13 10 9 15 0 11 1 9 1 9 1 9 13 2
14 9 1 9 1 15 0 9 1 9 13 14 13 4 2
18 13 4 4 16 9 1 0 0 0 9 12 9 1 1 13 4 4 2
10 15 15 9 1 9 14 13 4 4 2
9 15 1 0 9 15 0 13 4 2
16 11 11 11 1 0 10 0 9 11 1 0 9 1 9 13 2
12 15 11 1 0 9 15 9 9 1 13 4 2
20 10 9 9 1 1 2 9 11 11 1 13 0 9 1 9 14 0 9 13 2
6 15 12 0 9 13 2
8 15 9 1 0 9 0 13 2
18 9 1 13 13 16 10 9 9 11 7 9 11 1 9 9 13 4 2
14 15 1 11 11 7 11 11 11 11 13 1 9 13 2
15 11 1 14 12 9 1 11 9 1 0 9 1 9 13 2
10 10 9 15 11 1 9 13 4 4 2
15 0 9 9 7 0 9 15 1 9 1 12 9 13 4 2
13 9 1 12 9 1 11 1 15 3 0 9 13 2
7 15 1 14 0 9 13 2
9 10 0 9 0 9 1 0 13 2
19 10 9 15 1 9 1 0 9 7 0 9 1 0 9 1 13 4 4 2
18 9 1 1 15 1 11 1 0 9 13 15 15 1 3 0 9 13 2
13 11 1 0 0 9 11 0 9 1 10 0 13 2
9 9 1 15 3 0 9 13 4 2
15 10 9 13 16 15 11 1 1 11 1 15 9 13 4 2
11 10 9 1 11 11 1 9 11 1 13 2
32 10 9 10 9 1 9 13 4 2 10 9 15 1 10 9 14 14 13 4 16 10 9 9 1 1 0 9 1 15 9 13 2
6 9 14 15 13 4 2
23 9 11 1 14 12 9 1 9 1 0 11 9 9 9 1 0 2 0 9 0 13 4 2
29 10 9 14 9 2 9 1 9 1 13 16 9 9 11 1 15 0 9 11 11 1 9 1 11 1 9 13 4 2
15 10 9 7 9 1 14 9 13 2 9 1 0 9 11 2
16 11 9 15 9 1 1 1 9 1 9 1 9 13 4 4 2
18 0 9 1 13 11 1 13 1 3 9 1 10 9 0 13 4 4 2
18 11 1 0 9 1 11 11 7 11 1 9 9 2 3 13 4 4 2
23 0 10 9 1 15 9 13 3 13 4 15 15 0 9 7 9 15 9 1 10 14 13 2
22 10 9 1 9 1 9 1 15 13 1 9 15 9 1 15 1 0 13 4 13 4 2
19 11 1 9 1 9 9 12 9 1 9 12 9 1 14 13 4 4 4 2
10 11 1 9 15 0 9 0 13 4 2
11 11 11 15 1 0 9 1 1 12 13 2
11 15 11 11 1 1 1 14 13 4 4 2
17 0 9 1 0 10 9 1 9 9 1 0 9 13 4 4 4 2
10 15 9 11 9 1 11 1 13 4 2
14 15 14 9 0 9 1 15 9 1 9 13 13 4 2
17 15 1 14 11 11 13 2 15 11 2 11 2 11 13 4 4 2
13 3 9 1 0 9 1 9 14 13 14 13 4 2
26 10 9 11 9 1 0 9 1 0 9 1 13 13 4 2 15 12 9 11 11 1 9 3 13 4 2
30 11 1 14 12 9 1 0 10 9 1 9 9 11 1 15 9 13 4 2 7 15 10 0 2 0 9 13 4 4 2
14 11 1 0 9 1 15 14 12 9 9 1 13 4 2
14 11 9 1 0 3 0 9 1 1 12 13 4 4 2
11 11 1 10 9 1 11 9 1 13 4 2
22 0 9 1 13 11 11 11 1 9 11 11 1 9 1 9 11 9 1 13 4 4 2
15 11 1 1 14 15 9 14 0 14 9 1 13 4 4 2
12 11 11 2 11 2 1 1 14 13 4 4 2
14 0 9 1 0 9 1 9 9 1 0 9 13 11 2
24 9 1 9 11 1 12 9 1 0 11 1 9 11 1 0 0 9 1 3 0 7 0 13 2
21 12 0 0 9 1 0 10 9 1 0 9 1 1 0 11 7 9 14 0 13 2
23 9 9 1 9 1 0 10 9 1 9 11 11 11 1 1 11 11 11 1 13 4 4 2
15 11 0 10 9 1 9 3 0 9 1 13 13 4 4 2
17 13 4 4 16 10 9 1 11 7 15 9 1 9 13 4 4 2
15 3 0 9 11 11 1 9 0 9 9 11 1 13 4 2
22 15 12 0 9 13 16 11 1 9 11 11 2 0 11 2 1 12 9 1 9 13 2
8 11 11 1 12 9 1 13 2
18 0 9 15 13 16 10 9 1 11 1 9 1 1 1 13 4 4 2
20 9 11 11 9 1 9 1 0 13 7 15 9 1 0 9 1 13 4 4 2
11 9 11 11 2 0 9 1 1 0 13 2
19 10 9 1 0 9 1 11 1 12 9 11 7 11 1 9 13 4 4 2
13 10 9 2 0 9 1 0 9 1 1 0 13 2
8 9 1 15 9 14 15 13 2
14 12 9 1 15 0 9 3 9 1 13 4 4 4 2
16 15 15 1 1 9 13 4 10 12 9 11 1 0 9 13 2
12 10 9 9 1 0 0 9 1 0 9 13 2
13 15 14 9 13 4 10 9 11 11 1 13 4 2
12 10 9 0 9 1 0 9 1 9 13 4 2
12 11 1 0 9 9 1 9 13 4 4 4 2
8 15 0 9 9 9 13 4 2
14 11 1 12 14 9 1 13 13 4 12 0 9 13 2
26 13 4 4 16 10 9 9 9 1 13 9 15 13 4 4 2 15 3 1 15 1 13 4 4 4 2
16 9 1 14 1 11 11 11 11 1 9 1 9 13 4 4 2
13 10 9 1 11 1 9 1 13 0 9 0 13 2
25 9 1 0 9 13 2 11 11 1 9 2 11 1 0 9 7 9 1 13 4 9 1 9 14 2
15 11 1 12 9 9 1 0 9 11 2 11 2 0 13 2
14 15 11 11 1 0 9 11 1 13 4 9 0 13 2
15 10 9 1 0 9 1 11 7 11 9 2 9 13 4 2
17 0 9 1 10 9 1 9 1 9 1 11 11 1 0 9 13 2
3 15 13 2
16 3 14 9 14 1 15 14 9 11 1 9 13 4 4 4 2
17 7 3 14 11 1 11 1 1 9 11 13 1 1 0 13 4 2
12 11 1 11 1 11 11 1 9 13 4 4 2
17 10 9 11 1 9 1 9 14 9 1 9 1 1 13 4 4 2
3 15 13 2
10 11 2 11 2 11 9 1 0 13 2
19 15 12 0 14 9 9 14 13 2 7 0 0 9 11 12 9 1 13 2
10 11 1 11 1 9 14 12 9 13 2
15 9 9 1 12 1 12 9 1 9 1 13 4 4 4 2
8 11 1 9 7 9 0 13 2
15 11 0 9 1 14 9 1 10 0 9 1 13 4 4 2
3 15 13 2
9 11 1 13 1 1 10 9 13 2
17 11 11 1 1 1 9 7 9 9 1 13 7 9 1 9 13 2
17 15 1 10 9 9 7 9 13 2 15 9 1 13 4 4 4 2
12 0 9 13 1 1 11 3 0 9 14 13 2
14 15 9 1 13 4 13 1 1 14 12 9 0 13 2
20 12 0 9 13 1 1 11 1 9 1 0 9 13 1 1 9 3 13 4 2
8 0 9 7 9 1 0 13 2
12 11 1 0 9 13 1 1 15 0 9 13 2
6 0 13 4 11 1 9
16 11 1 10 14 9 13 2 10 15 1 9 10 0 9 13 2
15 9 9 1 12 1 12 0 2 0 9 1 0 9 13 2
18 15 1 13 1 0 9 7 9 13 1 1 14 3 0 9 9 13 2
22 11 11 1 14 9 1 1 9 1 15 14 9 14 13 2 7 0 9 3 13 4 2
27 11 1 9 9 1 0 9 1 0 9 1 14 9 13 4 4 2 15 0 9 1 9 14 9 13 4 2
13 11 1 0 0 9 1 11 1 9 9 13 4 2
18 10 9 1 9 15 13 4 7 9 1 0 9 15 1 1 13 4 2
18 10 14 9 10 9 1 9 1 13 4 2 15 15 9 3 13 4 2
14 9 1 1 3 13 1 10 9 15 13 9 13 4 2
24 11 11 1 9 2 9 11 1 9 7 11 1 9 11 1 9 12 1 10 2 14 9 13 2
18 15 13 4 4 16 11 2 11 7 11 11 1 10 9 13 4 4 2
20 10 9 1 9 11 1 11 1 13 7 10 9 11 1 9 1 9 13 4 2
23 15 10 9 1 9 13 11 1 9 9 14 10 15 1 9 1 13 0 9 1 0 13 2
18 10 9 1 13 12 1 9 1 0 7 0 9 10 9 11 13 4 2
9 10 9 1 15 14 13 13 4 2
17 15 9 1 13 13 4 2 16 15 1 15 13 0 9 13 4 2
9 11 1 9 12 9 1 0 13 2
13 0 9 1 9 1 13 12 0 9 13 4 4 2
20 10 9 1 11 11 1 0 9 2 9 3 13 1 9 13 2 13 4 4 2
16 9 1 9 1 9 13 14 0 3 9 13 4 2 0 9 2
13 10 9 1 9 9 1 1 0 12 9 1 13 2
14 9 1 9 1 10 9 1 9 15 9 1 13 4 2
10 15 12 0 2 14 0 9 14 13 2
21 16 10 9 1 15 9 1 9 2 11 1 9 2 13 1 9 0 13 4 4 2
14 15 10 9 1 13 1 9 13 2 11 11 1 1 2
20 9 2 9 7 9 1 9 10 9 1 9 9 11 1 11 11 1 13 4 2
26 11 11 1 9 1 9 1 13 1 3 2 15 9 1 9 1 1 1 15 10 9 1 9 13 4 2
10 10 12 0 9 1 14 12 9 13 2
16 0 9 1 0 9 2 9 1 9 7 0 9 1 13 4 2
7 0 9 1 0 9 13 2
15 10 9 1 1 0 11 9 7 10 0 9 13 4 4 2
17 9 1 1 0 9 1 13 4 11 11 3 14 0 13 4 4 2
13 15 15 13 16 9 1 9 1 9 13 4 4 2
19 11 11 11 11 1 9 11 1 9 10 9 1 9 2 9 1 9 13 2
13 9 9 1 9 1 10 9 1 13 10 13 4 2
18 10 9 1 1 14 12 9 1 2 11 11 2 1 9 13 4 4 2
10 10 9 0 9 9 11 1 0 13 2
21 12 9 7 12 9 0 10 9 1 9 11 11 1 15 0 0 9 1 13 4 2
14 11 11 11 1 9 1 3 10 0 7 0 9 13 2
21 11 11 0 9 1 1 13 10 9 1 1 11 1 9 1 3 0 9 13 4 2
13 11 11 1 11 1 9 13 1 3 12 9 13 2
25 9 1 1 16 11 1 9 11 1 12 9 13 4 4 2 16 15 15 9 1 1 0 13 4 2
37 10 9 1 0 13 1 1 9 11 11 1 11 1 9 10 10 9 11 1 13 16 0 9 1 9 14 14 13 7 11 1 9 14 0 13 4 2
35 9 11 1 9 1 1 15 9 13 2 10 9 9 1 1 0 0 9 1 13 4 9 1 11 1 13 7 15 15 9 1 0 13 4 2
14 11 1 9 1 12 10 0 9 13 2 11 1 9 2
9 9 1 10 9 9 11 1 13 2
21 11 15 15 11 1 9 13 4 7 15 1 15 9 13 9 1 9 13 4 4 2
24 9 9 1 1 1 12 9 9 13 2 15 13 9 1 9 10 3 1 0 13 4 4 4 2
8 9 1 11 0 12 9 13 2
12 10 9 1 9 12 0 2 14 11 11 13 2
20 15 11 1 9 12 11 1 13 4 9 1 0 14 9 1 3 13 4 4 2
17 10 9 1 13 1 9 14 3 0 9 1 1 1 0 13 4 2
9 15 9 1 11 9 13 4 4 2
30 15 0 11 9 1 13 4 7 10 9 13 4 4 2 15 14 10 11 1 13 1 9 3 11 1 9 13 4 4 2
3 15 13 2
13 11 9 1 10 9 1 9 7 9 1 13 4 2
15 11 1 14 12 9 1 9 9 13 15 11 13 4 4 2
7 3 15 9 9 14 13 2
3 15 13 2
13 11 1 11 9 1 1 11 1 9 13 0 13 2
10 10 3 15 1 9 10 0 13 4 2
3 15 13 2
10 11 12 0 2 0 7 0 9 13 2
14 15 3 1 13 1 9 1 1 10 12 9 9 13 2
15 0 9 9 14 9 1 13 1 1 0 9 0 13 4 2
15 11 9 1 9 1 1 15 1 3 0 9 13 2 11 2
16 15 0 9 1 9 13 15 9 12 9 9 1 0 13 4 2
19 15 13 1 9 10 9 1 9 7 9 13 15 9 11 11 1 13 4 2
16 11 1 1 12 9 13 2 15 11 7 11 14 13 4 4 2
15 9 11 9 1 9 13 1 3 10 9 1 9 13 4 2
3 15 13 2
17 11 1 9 10 9 11 11 1 1 11 11 1 9 13 4 4 2
14 11 11 1 9 9 11 7 11 9 1 1 13 4 2
13 11 1 9 11 9 1 9 1 1 13 4 4 2
18 11 1 11 1 1 15 9 13 9 7 9 1 9 1 0 13 4 2
13 11 1 1 15 1 9 3 10 0 13 4 4 2
3 15 13 2
22 11 1 12 9 1 9 9 0 13 1 3 11 0 9 1 11 1 9 9 13 4 2
14 11 1 9 15 9 9 7 0 9 1 13 4 4 2
10 11 0 11 0 3 0 9 9 13 2
17 11 1 15 13 1 1 9 7 9 14 9 1 9 0 13 4 2
3 15 13 2
21 9 1 13 1 1 11 7 15 0 9 1 9 9 2 0 9 7 9 0 13 2
14 11 1 9 1 13 1 3 15 1 0 9 3 13 2
18 9 1 9 9 7 9 1 1 9 9 13 16 9 13 1 9 13 2
46 15 3 0 9 1 9 2 9 2 9 1 1 0 9 1 0 9 1 13 13 4 15 9 1 0 9 1 9 13 1 15 0 9 13 4 4 7 9 2 9 1 9 0 13 4 2
8 15 2 11 11 2 13 4 2
19 11 1 1 14 9 1 13 4 14 12 1 12 9 0 9 1 9 13 2
14 12 9 3 9 1 13 4 0 9 10 9 11 13 2
9 10 9 9 1 3 0 9 13 2
12 9 1 1 10 10 9 1 9 0 13 4 2
18 11 11 11 11 1 13 2 15 9 9 1 12 9 1 9 1 13 2
11 15 1 0 11 11 7 11 11 13 4 2
22 15 10 9 1 9 1 0 12 9 13 15 9 2 9 2 9 7 9 1 9 13 2
21 9 14 11 11 1 0 9 1 9 13 1 3 9 1 15 9 1 9 9 13 2
7 0 9 10 9 11 13 2
7 11 11 12 0 9 13 2
19 9 9 1 1 11 11 1 15 9 14 13 4 7 12 9 9 13 4 2
24 11 1 1 14 0 9 1 13 1 1 15 9 9 13 4 15 12 9 1 9 1 13 4 2
17 0 0 9 15 9 1 14 13 4 7 0 9 9 11 9 13 2
7 0 9 10 9 11 13 2
22 10 9 11 11 1 0 0 9 1 0 13 2 15 9 9 1 14 12 9 1 13 2
18 15 0 14 0 9 13 2 15 1 10 9 1 9 13 4 4 4 2
7 11 11 12 9 0 13 2
10 11 11 0 11 1 3 0 9 13 2
15 9 14 13 1 3 10 9 0 9 15 0 9 11 13 2
11 10 9 12 9 7 10 9 1 13 4 2
20 15 1 11 9 1 9 1 10 0 9 13 2 15 11 11 1 9 13 4 2
11 11 11 11 11 11 1 3 0 9 13 2
8 15 9 13 4 2 9 14 2
8 15 11 1 3 0 9 13 2
13 15 9 1 9 13 9 1 0 9 13 4 4 2
12 10 9 1 9 11 11 1 11 1 13 4 2
16 10 9 1 9 11 1 0 9 13 2 15 9 12 9 13 2
16 9 11 1 1 14 15 9 11 7 11 1 9 14 0 13 2
7 10 9 12 9 0 13 2
18 11 1 11 9 1 9 0 10 9 1 9 1 9 1 13 4 4 2
20 10 9 11 9 1 13 2 7 15 0 11 9 1 9 15 0 13 4 4 2
13 9 1 9 1 12 9 1 0 11 1 9 13 2
13 10 9 1 9 11 11 1 9 11 1 13 4 2
17 9 1 14 12 9 1 11 11 1 9 11 1 15 9 13 4 2
19 10 9 1 12 9 1 11 1 9 13 2 15 10 9 0 13 4 4 2
14 10 9 1 3 0 9 15 13 16 15 0 9 13 2
13 15 9 1 12 12 0 2 0 9 13 4 4 2
7 15 9 13 4 9 14 2
13 10 9 1 9 11 1 9 11 9 1 0 13 2
32 12 9 1 14 0 12 9 1 13 4 13 4 10 9 10 9 1 0 13 16 15 1 10 9 2 9 1 9 13 4 4 2
8 15 11 1 3 0 9 13 2
14 15 12 9 0 2 12 9 0 7 12 9 0 13 2
13 10 9 1 9 11 11 1 9 11 1 13 4 2
17 10 9 11 1 11 9 1 13 4 3 0 9 1 1 12 13 2
11 10 9 1 9 1 12 9 0 11 13 2
21 10 11 1 0 9 1 0 10 9 13 2 15 15 14 9 2 9 13 4 4 2
22 10 9 1 1 15 1 11 11 2 11 11 2 11 11 2 7 11 11 14 0 13 2
9 11 1 1 1 10 9 0 13 2
12 13 4 2 16 10 9 9 9 1 13 4 2
16 15 0 9 1 9 13 1 1 10 9 1 9 13 4 4 2
16 15 14 13 4 4 16 11 9 9 2 9 1 9 13 4 2
22 15 9 13 2 16 0 9 1 13 1 3 14 9 1 9 1 1 9 9 13 4 2
46 9 1 9 1 9 2 15 15 9 1 9 13 2 1 9 15 13 4 15 0 13 1 1 9 9 13 1 1 9 13 4 4 7 0 9 1 13 15 0 9 15 9 13 13 4 2
34 10 9 7 10 9 9 1 9 1 1 9 1 1 0 9 1 9 9 13 16 10 9 1 12 0 0 9 1 9 7 9 14 13 2
45 11 1 0 0 9 1 15 1 12 9 2 11 11 11 2 11 11 2 9 9 2 9 9 2 11 11 2 11 11 2 0 2 0 7 0 9 7 0 7 0 9 13 1 13 2
19 11 11 1 11 1 9 1 9 0 9 2 9 9 9 1 13 4 4 2
12 10 9 1 9 1 9 1 14 0 9 13 2
23 9 9 1 0 9 1 9 1 13 4 4 2 15 11 2 11 7 15 9 13 4 4 2
25 12 9 7 12 1 10 9 1 9 1 1 11 11 11 11 2 11 9 1 3 0 9 9 13 2
13 11 11 1 0 9 13 15 11 9 13 4 4 2
24 12 9 0 0 0 9 7 11 11 11 11 15 9 9 1 9 13 4 2 0 0 9 13 2
25 9 9 1 12 9 0 0 9 1 9 1 9 1 15 9 13 7 11 9 1 9 13 0 13 2
15 11 1 9 11 1 3 0 9 11 11 9 1 0 13 2
11 10 9 9 1 12 9 1 9 1 13 2
18 10 9 9 1 9 11 1 0 13 2 15 9 1 9 1 9 13 2
22 11 1 12 9 1 1 12 13 1 1 1 15 9 9 1 0 9 9 13 4 4 2
20 9 1 1 15 9 11 1 9 1 9 13 2 15 15 10 9 1 9 13 2
15 14 15 9 11 7 9 11 1 15 15 15 9 14 13 2
30 11 14 13 15 9 1 9 13 4 7 15 15 13 16 15 9 1 9 13 4 4 2 15 10 9 9 1 13 4 2
13 0 11 15 9 1 13 4 15 2 15 13 4 2
15 15 9 1 9 15 2 15 13 15 1 9 1 9 13 2
22 11 1 9 11 1 9 9 13 15 9 9 13 7 15 10 9 1 3 10 9 13 2
15 9 1 9 1 14 9 9 1 9 1 0 9 0 13 2
20 9 1 0 9 1 9 13 4 7 9 9 1 9 2 9 9 13 4 4 2
11 9 1 10 9 12 9 0 13 4 4 2
11 0 9 10 9 1 9 1 13 4 4 2
8 10 3 9 1 9 13 4 2
11 10 9 1 2 11 11 2 13 4 4 2
14 11 1 9 10 12 9 1 9 1 9 13 4 4 2
14 13 4 4 16 10 3 9 13 1 9 0 14 13 2
3 15 13 2
10 11 11 1 10 0 9 1 13 4 2
14 15 1 13 1 1 9 2 9 7 0 9 0 13 2
11 11 1 11 2 11 1 9 13 4 4 2
42 11 1 11 11 2 11 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 1 13 4 4 4 2
13 11 7 11 1 11 0 9 1 3 13 4 4 2
17 11 11 2 11 11 7 11 11 1 0 9 15 1 1 0 13 2
3 15 13 2
19 0 9 1 9 1 9 2 9 9 2 9 7 9 9 1 13 4 4 2
3 15 13 2
9 11 1 10 9 1 9 0 13 2
18 9 7 9 9 1 1 0 9 1 9 7 9 9 1 13 4 4 2
17 11 1 0 9 1 1 10 14 9 13 2 15 13 4 4 4 2
14 2 11 11 2 11 1 14 12 9 9 1 0 13 2
10 0 9 1 15 11 9 1 9 13 2
15 15 1 9 7 0 9 9 1 9 1 0 9 13 4 2
15 11 9 1 1 1 9 1 13 15 3 14 0 9 13 2
17 15 9 11 1 9 13 2 15 10 9 9 1 9 13 4 4 2
14 11 9 1 9 13 1 1 9 7 9 9 13 4 2
17 13 4 4 16 0 9 1 15 11 11 9 1 3 0 9 13 2
19 10 9 1 12 9 1 9 13 7 15 11 1 12 9 1 9 1 13 2
12 15 11 1 11 1 12 9 1 9 1 13 2
23 15 9 12 0 9 1 13 4 2 15 11 11 1 11 1 9 13 1 9 1 13 4 2
17 15 1 11 2 11 7 11 10 9 1 9 0 9 1 13 4 2
19 15 1 11 11 14 13 2 15 1 13 1 1 0 9 1 9 13 4 2
14 15 12 0 9 14 13 2 15 0 9 13 4 4 2
7 11 15 1 0 9 13 2
23 10 9 15 9 1 9 1 9 13 4 7 9 1 9 13 15 9 1 1 9 13 4 2
12 9 9 1 1 9 1 9 9 13 4 4 2
34 9 1 9 1 1 10 9 10 0 15 13 4 4 2 16 15 9 9 1 9 1 9 13 4 7 10 9 9 9 1 0 13 4 2
14 11 1 10 9 1 9 1 9 1 9 13 4 4 2
16 9 9 9 13 1 1 1 15 9 1 9 14 13 4 4 2
12 9 0 13 16 9 9 1 14 13 0 13 2
33 11 1 11 1 9 13 11 11 11 11 1 9 1 0 10 9 13 15 15 1 0 9 1 11 1 9 11 11 1 1 9 13 2
23 0 13 16 11 1 14 15 9 1 9 0 13 4 7 15 1 0 9 1 9 13 4 2
13 7 9 1 10 9 1 15 9 1 0 13 4 2
30 16 0 9 1 0 9 1 9 1 9 13 4 7 0 9 1 1 9 1 1 15 9 1 1 15 9 14 13 4 2
15 9 9 1 11 11 1 0 9 11 1 14 9 13 4 2
15 11 1 1 11 1 15 15 0 9 1 13 0 9 13 2
13 10 9 1 11 11 1 14 1 9 9 13 4 2
10 10 9 1 15 9 11 11 13 4 2
19 16 11 1 9 15 1 13 4 15 11 1 9 10 9 1 10 0 13 2
19 15 1 11 1 0 9 1 11 11 11 11 1 9 0 14 9 1 13 2
25 9 1 9 9 1 13 9 1 1 0 9 13 4 4 7 15 15 14 9 1 9 14 13 13 2
32 3 12 0 9 1 1 9 1 9 13 4 11 1 9 9 9 1 15 0 9 11 11 11 1 9 14 13 1 9 13 4 2
15 3 15 10 9 1 0 3 11 11 11 1 13 13 4 2
29 11 1 11 1 12 9 9 1 9 1 1 13 16 15 10 9 1 15 0 9 1 10 9 1 0 14 13 13 2
11 15 3 15 11 1 10 9 13 13 4 2
13 11 1 13 16 15 10 9 11 11 1 8 13 2
22 9 1 9 13 4 11 1 0 9 1 13 13 16 15 3 14 9 1 9 9 13 2
15 0 13 16 11 1 0 12 9 1 9 9 14 13 4 2
17 9 1 10 9 0 9 11 1 13 15 9 9 1 9 1 13 2
32 9 1 9 13 1 12 9 1 13 4 16 9 15 13 4 16 9 9 1 0 11 1 9 1 1 0 9 7 9 3 13 2
34 9 1 1 9 1 9 1 0 9 1 9 9 13 1 9 13 4 2 7 15 11 11 11 1 13 4 1 15 9 1 1 14 13 2
15 9 1 13 4 16 10 9 1 0 9 3 1 13 4 2
36 0 2 0 9 1 13 11 1 12 0 9 9 1 9 1 10 9 1 9 0 13 4 13 16 15 9 1 9 1 9 1 13 1 9 13 2
15 0 13 16 11 11 2 11 1 11 1 0 13 4 4 2
15 10 9 1 0 12 9 1 9 1 9 14 14 13 4 2
25 11 1 15 11 1 9 9 0 13 4 2 7 11 1 10 9 1 15 14 9 14 13 4 4 2
20 11 11 9 1 9 13 4 16 15 10 9 1 9 1 9 9 13 4 4 2
23 11 11 11 1 14 9 1 0 9 1 9 9 14 13 4 1 1 15 9 0 13 4 2
35 0 13 16 9 1 9 1 9 14 13 1 1 11 11 1 9 1 13 4 1 9 12 12 1 0 9 1 14 11 1 9 13 4 4 2
29 11 1 15 9 1 9 9 13 1 11 11 1 11 1 12 9 1 9 1 13 4 11 11 11 1 9 0 13 2
11 10 9 13 1 11 9 1 0 9 13 2
6 10 9 11 1 13 2
26 11 1 9 1 11 1 11 11 1 0 9 1 13 16 9 1 9 1 1 14 15 15 1 13 4 2
16 11 1 11 9 1 11 1 11 11 1 10 9 0 13 4 2
39 9 1 1 11 1 13 16 9 1 1 1 15 15 9 13 4 15 15 10 9 1 15 1 9 14 13 2 16 15 13 13 4 4 16 10 9 8 13 2
11 9 1 12 9 1 9 1 9 13 4 2
22 11 1 13 16 9 1 1 1 15 12 12 0 9 2 14 12 12 9 2 13 4 2
11 15 12 2 12 9 1 11 13 4 4 2
25 15 13 16 15 15 9 9 11 1 11 11 7 11 11 7 11 1 11 1 0 9 13 13 4 2
20 11 1 9 11 11 11 9 9 13 7 11 2 11 1 9 1 1 13 4 2
20 15 13 16 9 1 14 15 15 9 1 14 13 16 9 10 9 1 9 13 2
11 7 2 15 0 9 1 1 15 13 4 2
10 15 9 1 14 0 9 1 0 13 2
38 10 9 1 9 13 4 11 1 0 9 15 15 9 13 9 1 1 13 16 15 9 13 4 4 15 0 9 1 9 1 9 13 4 7 9 13 4 2
27 0 9 1 1 9 0 11 11 11 11 11 1 15 11 11 9 1 9 0 0 9 1 1 9 13 4 2
23 11 1 9 1 0 9 1 13 1 10 9 9 1 12 9 1 0 9 1 0 9 13 2
19 11 11 11 1 11 1 0 9 1 15 0 9 11 11 11 1 9 13 2
14 10 9 1 11 11 11 14 15 9 1 1 0 13 2
15 15 1 10 9 9 7 9 9 1 0 9 14 0 13 2
14 11 11 1 11 1 11 0 11 1 9 13 4 4 2
11 0 9 1 1 15 9 11 13 4 4 2
17 11 1 11 1 11 11 1 11 1 13 11 1 0 9 13 4 2
10 15 1 11 1 9 1 9 9 13 2
11 15 15 12 9 7 12 9 1 9 13 2
14 11 11 1 12 9 13 0 11 11 1 0 9 13 2
20 10 9 9 0 13 4 7 0 9 11 11 0 13 2 1 9 1 13 4 2
17 0 9 2 9 2 11 11 1 9 1 13 1 0 9 9 13 2
19 15 9 13 1 1 15 11 9 1 0 11 9 1 14 12 9 13 4 2
60 10 9 1 0 11 11 11 11 2 0 11 11 11 11 2 11 11 11 11 2 11 11 11 11 2 11 9 11 11 1 9 11 11 7 11 11 2 11 11 1 11 11 11 11 2 11 11 11 7 11 11 11 1 9 11 11 14 0 13 2
21 15 1 10 0 9 7 10 9 1 11 7 11 14 11 1 0 9 1 0 13 2
23 11 11 11 1 11 1 11 11 9 1 9 11 1 9 1 1 12 9 9 1 9 13 2
10 3 1 15 11 11 1 9 13 4 2
27 11 11 1 0 9 1 9 13 1 1 11 11 11 9 9 15 9 11 11 1 1 0 9 1 11 13 2
11 15 9 1 3 11 11 0 9 9 13 2
13 0 13 16 11 1 1 14 11 11 9 1 13 2
13 15 11 1 11 1 1 11 9 1 11 11 13 2
25 11 11 1 9 7 11 11 1 11 11 11 11 1 11 1 12 9 3 11 11 13 1 9 13 2
22 11 7 11 1 0 9 13 4 15 13 16 10 12 9 1 9 1 9 13 4 4 2
54 15 1 14 15 13 16 11 11 9 0 12 9 1 9 0 9 9 1 11 1 9 9 11 11 1 9 13 2 15 14 9 1 0 12 9 1 9 1 9 0 13 4 7 15 9 1 9 13 1 9 1 13 4 2
21 11 1 11 1 15 9 9 1 13 16 11 11 11 7 11 1 0 9 13 4 2
34 15 13 16 11 11 1 1 9 13 4 4 7 15 1 9 13 16 11 11 1 0 9 1 10 0 9 1 9 1 9 13 4 4 2
17 15 1 1 9 1 11 1 9 1 9 12 1 13 12 13 4 2
13 15 1 11 11 1 11 1 9 1 9 13 4 2
28 11 1 13 16 15 15 11 1 0 13 1 1 9 13 4 4 15 11 11 1 0 13 1 9 13 4 4 2
30 11 1 9 9 1 1 1 11 1 13 16 15 11 11 11 1 9 11 11 1 13 4 16 15 11 11 1 9 13 2
21 15 13 16 9 1 13 1 9 1 3 13 1 9 9 10 9 1 9 0 13 2
14 11 1 13 16 11 1 11 0 9 1 1 1 13 2
33 15 1 14 15 9 13 16 9 14 1 11 13 11 1 13 0 11 11 11 0 9 9 1 9 1 1 1 11 9 1 9 13 2
37 9 1 9 13 4 11 1 13 16 15 15 13 11 1 0 13 4 16 15 15 9 13 2 7 15 13 1 3 0 13 16 15 13 14 4 4 2
17 9 1 11 9 11 11 7 9 11 11 7 11 1 14 0 13 2
37 9 1 0 2 0 7 0 9 1 1 11 1 9 11 11 1 11 1 0 0 9 1 0 9 9 1 11 2 11 7 11 1 9 1 0 13 2
15 15 13 16 11 1 11 1 9 9 1 9 12 9 13 2
9 15 9 0 9 1 0 13 4 2
19 15 9 13 16 9 11 11 11 1 9 1 11 11 1 9 1 9 13 2
10 9 1 0 9 13 15 9 13 4 2
19 9 9 1 12 9 3 13 16 9 1 9 10 13 7 9 9 14 13 2
25 11 1 13 16 11 11 11 1 9 1 11 1 9 1 9 1 13 11 1 9 1 9 14 13 2
21 11 11 1 15 1 9 1 0 9 1 9 13 4 9 1 9 13 1 9 13 2
18 9 11 7 9 11 11 11 1 9 13 4 15 0 9 1 0 13 2
11 11 1 13 4 16 10 15 9 14 13 2
24 12 9 1 11 1 9 11 11 7 9 11 11 1 1 0 9 1 9 13 9 1 0 13 2
11 7 9 1 9 1 10 9 1 13 4 2
8 15 9 11 1 9 1 13 2
32 9 1 9 1 13 1 9 9 1 9 1 9 9 1 11 1 9 9 1 12 9 1 9 7 12 12 9 1 9 13 13 2
42 9 11 11 11 1 11 11 1 9 7 0 11 11 11 11 1 11 9 1 1 14 9 1 0 9 11 11 11 1 10 9 1 9 1 9 1 13 9 13 4 4 2
21 15 13 16 12 9 1 3 11 1 11 11 1 9 1 11 13 1 9 1 13 2
11 11 2 11 1 9 1 11 1 9 13 2
21 10 9 1 0 9 7 9 1 13 7 13 1 9 11 11 11 1 9 1 13 2
23 10 9 9 1 9 9 1 9 13 4 4 2 7 9 1 9 9 1 9 1 13 4 2
8 10 9 1 9 15 9 13 2
32 11 1 13 16 9 3 9 1 9 9 13 1 1 9 13 4 4 7 9 9 1 9 1 0 9 1 0 13 9 13 4 2
19 9 14 1 14 9 1 9 9 1 0 9 1 0 13 1 9 13 4 2
10 15 9 1 12 9 1 9 13 4 2
34 15 9 11 11 11 1 9 1 11 11 11 2 11 11 11 2 11 11 11 2 11 11 11 7 11 11 11 1 9 0 9 1 13 2
22 11 11 1 9 1 11 1 11 1 9 13 1 9 1 10 9 1 11 1 9 13 2
19 11 1 13 16 10 9 0 13 2 7 9 1 15 9 14 13 4 4 2
15 11 1 13 16 9 11 1 0 9 1 9 11 9 13 2
21 15 9 1 13 16 9 1 0 9 1 1 0 13 7 9 1 9 1 3 13 2
27 11 11 11 11 11 11 11 11 1 9 11 11 1 15 1 0 9 9 1 9 13 4 9 13 4 4 2
7 11 9 1 9 9 13 2
23 15 13 16 9 1 0 9 1 9 1 9 7 0 9 1 11 1 9 13 4 4 4 2
23 11 1 9 1 0 13 4 11 15 9 1 3 0 9 9 9 1 9 13 4 4 4 2
44 15 13 16 11 11 1 9 11 11 11 1 9 1 9 13 1 9 13 4 4 7 0 9 9 1 2 15 11 1 0 13 4 2 15 9 9 13 1 9 13 4 4 4 2
26 11 1 9 13 16 11 9 11 1 15 9 13 13 4 2 15 11 11 1 15 0 9 14 13 4 2
14 16 11 10 9 1 15 14 9 1 9 13 4 4 2
36 11 1 9 0 11 11 11 1 3 0 9 11 1 11 1 0 9 7 0 9 11 11 1 9 13 16 15 9 9 1 1 9 13 4 4 2
29 11 1 0 9 11 11 1 9 13 14 11 1 11 1 10 9 1 1 9 13 16 9 9 15 9 1 13 4 2
31 10 9 11 1 11 9 11 11 1 9 13 16 15 14 9 1 11 2 11 7 11 1 0 9 1 1 9 13 4 4 2
46 11 1 3 0 9 1 13 16 10 9 1 9 1 9 1 3 10 9 13 2 15 14 9 1 13 4 4 4 7 0 9 9 9 1 9 13 11 2 11 11 1 9 13 4 4 2
22 15 10 9 1 9 1 9 13 16 15 9 11 11 1 9 13 1 15 9 13 4 2
11 11 1 13 16 15 9 1 0 14 13 2
35 11 1 10 9 1 12 0 9 1 9 13 4 7 9 9 9 1 13 4 2 15 12 9 3 0 9 1 9 1 13 4 13 4 4 2
8 9 1 12 1 10 9 13 2
15 7 3 14 15 9 13 15 10 9 12 9 14 13 4 2
23 15 15 9 1 9 1 13 4 16 15 9 1 9 7 9 1 1 0 13 9 13 4 2
27 7 10 9 1 14 9 14 14 13 15 9 1 9 1 13 9 7 9 14 13 1 1 9 13 4 4 2
11 3 9 9 9 1 9 13 4 4 4 2
11 15 9 2 9 7 9 1 9 13 4 2
20 9 9 1 1 10 9 9 1 9 13 4 7 15 9 1 15 9 14 13 2
16 9 11 1 0 11 11 14 10 9 1 9 1 13 14 13 2
11 11 1 12 9 1 12 9 13 4 4 2
22 15 0 11 1 14 15 12 9 1 11 9 1 9 1 0 9 1 9 13 4 4 2
25 15 1 11 11 1 11 11 9 1 12 10 9 1 9 9 1 9 1 9 13 9 13 4 4 2
15 11 1 11 11 1 15 1 12 9 1 9 13 4 4 2
35 15 11 9 1 12 9 1 0 9 1 1 12 0 9 1 0 13 1 1 9 9 1 15 13 12 9 1 14 9 1 9 13 4 4 2
22 0 11 9 1 11 1 12 9 1 11 11 1 11 11 9 1 9 1 13 4 4 2
27 11 11 1 11 1 11 11 1 11 9 1 11 11 9 1 12 0 9 1 0 9 1 9 13 4 4 2
13 15 0 11 1 9 13 1 0 9 1 9 13 2
18 15 10 10 9 13 15 9 1 9 7 15 0 9 1 9 13 4 2
9 15 13 15 15 9 1 10 9 2
14 15 3 0 9 13 15 0 9 9 7 0 0 9 2
19 11 11 11 1 9 1 1 9 1 9 1 9 11 1 10 12 9 13 2
14 7 10 9 1 14 12 9 1 14 13 4 4 4 2
13 15 1 14 14 12 2 12 9 9 14 0 13 2
12 10 9 15 1 9 13 1 9 13 4 4 2
20 0 9 1 12 0 9 0 9 11 11 1 14 12 10 9 1 3 13 4 2
12 15 1 9 11 11 1 9 15 12 9 13 2
12 15 0 12 9 1 9 1 9 13 4 4 2
14 10 12 9 15 9 13 7 15 1 9 9 1 13 2
14 11 11 11 2 11 1 0 9 9 1 0 13 4 2
7 15 15 15 14 14 13 2
17 9 1 10 9 13 2 15 15 9 1 0 13 4 0 9 13 2
21 9 1 9 1 9 9 1 13 10 0 9 1 9 1 13 1 0 13 4 4 2
14 9 13 1 1 15 9 2 9 1 9 13 4 4 2
15 0 9 1 15 9 2 9 1 9 1 9 13 4 4 2
14 15 9 1 13 1 1 14 9 1 9 13 4 4 2
37 10 9 13 4 16 0 9 14 3 14 9 13 4 4 4 7 10 9 1 9 2 9 7 9 1 9 1 9 0 13 4 2 15 0 13 4 2
20 7 0 3 0 9 1 9 9 1 15 9 1 9 1 1 1 9 13 4 2
24 10 0 9 9 14 15 1 15 9 1 9 14 13 4 7 10 15 13 4 9 1 9 1 2
27 11 1 3 0 9 7 0 9 1 11 1 13 4 9 9 11 11 1 0 9 1 9 13 4 4 4 2
16 9 1 15 1 12 12 0 0 9 0 13 1 9 13 4 2
28 10 9 10 9 1 1 0 13 4 4 2 15 11 2 11 7 11 1 9 1 1 1 11 11 1 0 13 2
18 10 9 1 0 13 1 11 1 12 9 1 9 13 1 9 13 4 2
10 10 10 9 15 15 9 0 13 4 2
11 15 11 14 15 0 9 1 13 4 4 2
37 0 9 1 15 13 16 11 1 9 1 0 9 11 1 12 9 0 13 11 11 7 11 1 13 9 1 1 12 0 0 9 0 13 1 9 13 2
9 10 9 1 11 1 14 9 13 2
10 10 9 10 12 9 9 1 13 4 2
8 10 9 1 11 14 0 13 2
21 15 1 11 1 0 9 13 16 15 15 9 1 0 9 1 13 11 1 3 13 2
24 15 1 2 11 1 0 9 7 0 9 1 9 1 12 9 1 0 9 13 1 14 9 13 2
20 11 11 1 11 11 1 1 0 9 1 9 1 11 1 9 0 13 4 4 2
21 11 1 11 9 9 1 0 11 1 11 11 1 10 9 1 0 9 13 4 4 2
19 15 15 9 9 11 1 11 0 13 7 15 1 0 9 11 2 11 13 2
26 11 1 13 13 16 11 11 1 11 9 1 13 4 4 7 15 1 15 0 9 1 9 13 4 4 2
15 11 1 11 1 11 1 0 9 1 0 9 9 13 4 2
18 15 1 14 11 1 15 9 0 13 1 1 11 11 1 9 13 4 2
20 11 1 1 11 1 1 10 0 9 0 13 1 3 11 1 9 13 4 4 2
16 15 13 16 11 1 11 1 9 13 1 1 3 0 9 13 2
31 11 11 11 1 9 9 1 9 1 9 1 11 1 11 1 9 1 13 16 11 1 9 1 9 13 1 15 9 14 13 2
14 11 11 9 13 1 15 9 1 13 4 0 9 13 2
23 15 13 16 9 1 9 2 9 13 1 1 9 1 9 13 1 1 10 15 9 14 13 2
46 9 1 9 2 9 1 0 9 1 0 13 1 1 9 9 1 11 1 9 13 4 11 1 13 16 9 1 3 0 9 1 1 1 13 1 3 11 1 9 13 1 9 0 13 4 2
24 7 11 1 9 0 13 1 1 11 1 11 11 1 9 13 1 1 0 14 13 1 9 13 2
29 11 1 13 16 11 1 11 1 9 1 9 13 15 11 1 13 4 2 7 11 1 15 9 13 11 13 4 4 2
19 9 1 9 1 1 1 15 13 16 15 1 1 9 9 9 1 9 13 2
25 9 1 1 0 9 1 0 9 1 1 1 15 9 13 4 13 16 9 1 1 0 9 13 4 2
28 11 11 11 11 11 2 11 2 11 1 9 11 1 11 1 0 9 7 11 1 0 9 1 13 1 9 13 2
15 11 1 10 9 1 1 15 0 13 1 9 0 13 4 2
32 0 9 1 1 11 11 1 11 1 9 13 4 16 11 11 11 11 11 1 9 9 1 9 1 1 9 1 9 13 4 4 2
28 15 13 2 10 9 1 14 9 13 16 11 1 0 9 1 11 1 9 9 13 1 3 9 1 9 13 4 2
23 9 1 13 16 15 1 3 10 0 9 11 1 0 9 7 11 1 0 9 13 4 4 2
18 15 13 16 16 10 3 9 0 14 13 16 15 10 9 13 4 4 2
16 9 1 13 16 11 1 9 2 9 1 9 1 9 13 4 2
14 10 9 1 11 1 9 1 0 13 1 9 13 4 2
28 15 13 2 15 0 9 0 13 1 1 11 7 11 9 1 9 1 13 7 3 14 15 0 13 1 9 13 2
24 0 13 16 11 11 2 11 2 11 7 11 1 12 9 1 10 0 9 1 9 15 11 13 2
19 11 11 1 9 9 1 1 11 1 0 13 1 10 9 0 13 4 4 2
31 15 1 11 1 9 1 9 13 7 11 1 9 1 9 0 13 1 1 11 1 11 1 15 0 13 1 9 13 4 4 2
25 9 9 1 1 15 10 12 9 9 1 9 7 9 1 0 13 1 14 9 1 9 13 4 4 2
19 11 7 11 1 1 13 9 1 9 11 1 9 1 14 13 4 4 4 2
14 11 1 0 9 9 0 9 1 9 1 13 4 4 2
17 9 15 12 9 1 1 13 9 1 9 1 1 1 13 4 4 2
12 0 9 15 12 0 0 9 14 13 4 4 2
29 10 9 1 9 1 1 11 11 7 11 1 1 0 9 1 9 13 1 0 9 15 9 1 9 1 13 4 4 2
11 15 15 9 9 1 14 13 4 4 4 2
7 15 15 0 9 14 13 2
12 0 9 1 10 9 1 1 0 9 13 4 2
28 11 1 1 10 9 1 9 10 9 1 0 13 4 16 12 9 1 1 10 0 9 1 12 0 9 13 4 2
20 11 1 11 9 1 1 11 1 10 9 11 11 11 11 13 4 11 13 4 2
23 0 11 1 12 0 11 11 1 13 16 11 1 0 12 9 1 9 1 10 9 13 4 2
18 15 9 3 10 13 4 4 16 14 0 9 14 15 9 13 4 4 2
26 16 11 1 9 1 9 11 9 1 0 13 4 4 2 7 9 1 1 1 15 3 14 9 13 4 2
16 0 9 9 1 9 1 9 1 12 0 0 9 13 4 4 2
9 15 9 1 9 1 9 13 4 2
15 3 0 11 11 1 9 1 1 10 9 1 10 9 13 2
24 9 1 9 10 9 1 1 9 1 9 1 15 9 1 13 4 14 16 9 1 9 0 13 2
20 9 7 15 1 9 2 11 11 11 11 1 10 9 15 15 14 13 4 4 2
10 13 4 16 10 9 15 13 4 4 2
4 3 0 9 2
18 16 15 8 13 16 0 0 9 9 1 9 14 9 13 13 4 4 2
19 11 11 11 11 1 11 1 0 9 13 7 9 1 9 9 1 14 13 2
54 11 1 9 9 11 11 1 1 0 9 9 11 11 1 12 9 9 13 7 13 16 15 11 1 10 9 0 13 4 2 15 11 11 1 13 9 7 9 11 11 1 13 1 9 11 11 11 1 11 11 1 13 4 2
25 15 15 13 4 16 15 10 11 11 13 15 0 11 11 11 7 0 11 11 1 9 9 13 4 2
26 16 2 11 11 11 11 1 11 11 1 0 9 1 1 11 11 1 14 10 14 10 9 13 14 4 2
16 16 15 15 11 1 12 9 11 1 12 12 9 1 13 4 2
15 9 15 0 13 4 15 11 11 1 3 9 0 13 4 2
33 15 13 2 3 15 15 12 9 1 11 11 1 12 9 1 9 1 9 1 13 13 4 15 15 9 0 13 1 1 9 13 4 2
7 11 1 12 9 0 13 2
16 15 11 1 0 0 9 1 9 7 13 4 9 13 4 4 2
10 11 11 9 1 9 1 0 0 13 2
10 11 1 3 15 9 10 9 13 4 2
21 9 2 9 1 15 13 16 11 11 1 15 9 9 1 9 1 9 13 4 4 2
27 15 15 13 4 16 11 11 15 13 4 9 9 13 7 10 9 15 11 11 11 11 1 15 9 13 4 2
21 9 13 16 11 1 9 0 13 16 9 9 10 9 14 13 15 15 9 13 4 2
15 11 1 13 16 15 7 11 11 1 9 1 0 9 13 2
7 9 1 9 14 0 13 2
13 11 1 13 16 15 9 9 9 1 13 4 4 2
18 7 11 1 9 1 9 1 1 2 9 9 1 10 9 13 4 4 2
23 11 1 10 9 1 10 9 0 13 2 10 9 1 15 13 16 15 9 10 0 0 13 2
8 7 11 1 9 9 13 4 2
16 10 9 0 9 1 13 4 4 7 15 15 9 14 13 4 2
17 9 9 1 13 13 16 3 10 9 7 9 9 9 1 13 4 2
38 11 16 9 1 11 2 11 13 15 15 9 13 1 10 9 1 9 14 13 14 4 16 9 3 14 13 7 9 7 9 9 1 9 1 9 14 13 2
25 16 16 9 11 11 13 4 16 16 15 9 1 9 14 13 4 16 13 4 16 15 10 9 13 2
22 9 7 9 10 9 1 9 13 4 4 16 0 9 15 9 1 9 7 9 14 13 2
23 9 11 11 1 13 13 16 15 10 9 7 9 9 13 14 15 10 9 9 13 4 4 2
10 15 10 9 10 9 1 14 13 13 2
17 11 1 11 1 9 11 11 11 1 15 9 1 9 13 4 4 2
26 9 1 13 16 11 1 15 9 0 9 1 9 9 13 1 12 9 1 11 11 11 1 13 4 4 2
25 11 1 11 1 11 11 11 1 9 13 15 11 11 1 9 1 0 0 9 1 9 1 9 13 2
54 11 9 1 9 1 1 0 7 0 9 1 0 13 4 11 1 9 9 1 11 1 11 1 11 9 1 11 11 11 2 11 2 1 11 11 11 1 11 1 1 9 9 0 13 7 9 1 0 13 1 9 13 4 2
43 11 11 1 0 11 11 11 11 1 11 1 9 1 1 9 0 13 1 9 1 9 13 4 9 13 4 16 11 9 1 11 9 11 9 1 1 9 1 9 1 9 13 2
24 9 1 13 16 11 1 11 9 1 1 1 15 9 13 4 1 1 1 9 1 9 13 4 2
37 16 11 9 1 11 9 1 15 0 13 0 13 16 9 9 0 13 1 1 11 1 9 1 13 4 4 7 3 15 9 1 15 9 1 13 4 2
27 11 1 11 1 11 11 11 1 9 13 15 11 11 1 9 1 0 0 9 1 1 15 9 1 9 13 2
45 3 2 11 2 11 1 11 1 9 9 1 9 11 11 11 1 9 1 13 16 15 11 9 1 11 11 11 1 11 7 11 1 10 9 1 1 9 1 0 13 1 9 13 4 2
38 15 13 16 9 1 9 13 1 1 0 9 1 11 1 1 9 9 13 7 9 1 11 1 0 9 1 9 1 0 13 1 0 9 13 1 9 13 2
29 15 13 16 11 11 11 7 11 11 11 7 9 9 1 1 9 1 0 9 1 1 9 1 9 13 1 9 13 2
30 9 11 11 1 9 1 11 11 1 0 11 11 11 11 1 11 1 9 1 1 9 0 13 1 9 1 9 13 4 2
19 9 1 9 13 4 16 0 9 11 9 1 1 9 1 9 1 9 13 2
26 11 1 13 16 15 11 1 9 1 9 13 4 2 15 15 9 1 1 9 0 13 1 9 13 4 2
6 15 12 0 9 13 2
18 9 1 0 9 1 0 11 1 9 15 11 1 0 9 1 14 13 2
26 11 1 11 11 1 9 1 11 9 1 1 9 0 9 10 9 13 4 15 0 9 13 1 13 4 2
28 11 9 9 11 1 9 1 11 9 1 13 4 9 1 9 1 9 13 11 1 9 1 9 9 13 4 4 2
30 16 9 1 14 9 1 1 0 11 1 10 9 15 0 13 16 12 9 1 1 9 1 10 9 15 15 9 1 13 2
25 0 9 1 0 10 9 9 1 11 1 1 11 11 11 1 13 4 4 15 0 9 1 1 13 2
18 9 9 1 0 0 9 9 11 1 9 9 1 14 9 13 4 4 2
26 9 1 0 9 1 0 13 4 1 10 9 2 9 9 1 0 9 11 1 1 1 15 13 4 4 2
26 11 9 1 9 1 13 1 9 11 9 1 12 9 9 1 13 4 12 12 9 1 9 0 13 4 2
39 11 2 9 9 1 9 11 11 1 13 13 16 9 1 9 16 9 1 1 13 16 12 9 1 1 9 1 0 9 1 1 15 9 11 11 1 13 4 2
29 15 13 16 11 9 1 0 9 13 9 11 9 1 9 1 9 1 13 4 4 2 16 0 9 1 9 14 13 2
20 0 13 16 9 1 9 1 0 9 13 1 9 1 9 1 10 9 13 4 2
33 15 13 16 11 1 9 11 1 0 2 0 13 1 1 9 9 1 0 0 11 11 1 15 1 11 1 9 13 1 9 13 4 2
23 15 1 1 11 1 11 1 12 12 9 13 10 9 1 11 1 11 1 13 1 1 13 2
22 3 0 7 0 9 1 9 9 0 9 1 9 7 0 9 13 1 9 13 4 4 2
40 11 1 13 16 9 1 1 3 14 9 0 13 4 4 4 7 10 9 1 13 14 11 1 9 1 15 10 9 1 1 0 9 1 1 1 11 11 13 4 2
26 15 13 16 11 11 11 1 12 0 9 13 4 4 4 7 15 1 9 1 9 11 1 14 13 4 2
24 9 1 9 13 1 3 0 13 4 2 16 10 9 15 9 15 9 1 9 13 13 4 4 2
16 15 9 1 12 0 9 13 4 4 2 15 1 9 0 13 2
11 16 0 9 1 1 15 9 1 13 4 2
36 9 1 9 1 13 9 1 13 16 11 2 11 2 11 11 2 11 7 11 11 11 1 9 8 13 1 9 1 9 1 8 13 4 4 4 2
21 9 9 1 13 13 16 11 9 1 0 9 1 1 9 1 9 13 4 4 4 2
27 9 13 4 16 16 11 1 0 9 9 1 13 2 16 15 9 15 0 9 1 9 1 8 13 4 4 2
17 9 1 11 9 9 0 9 2 9 1 9 0 2 0 13 4 2
20 10 9 1 9 13 4 7 9 2 9 9 7 9 2 9 1 9 13 4 2
17 0 9 1 9 9 14 12 12 9 9 13 15 9 9 1 13 2
20 15 15 9 1 0 9 14 14 13 4 7 0 9 1 9 13 4 4 4 2
24 9 7 9 13 4 1 10 9 1 9 0 13 4 16 9 9 9 1 9 0 13 4 4 2
10 9 12 12 9 1 12 9 9 13 2
8 10 9 1 0 9 14 13 2
16 9 9 1 9 1 1 0 12 9 1 9 13 1 9 13 2
14 0 9 1 9 13 4 7 9 1 9 1 9 13 2
10 0 9 12 9 9 13 1 9 13 2
24 9 9 1 12 9 1 13 16 11 7 11 1 9 1 0 0 9 1 1 10 9 13 4 2
12 11 1 14 15 9 1 9 1 9 13 4 2
25 0 2 0 11 2 0 11 2 11 2 11 7 11 1 1 13 0 9 1 1 11 1 9 13 2
12 12 9 1 1 11 1 0 9 13 4 4 2
10 15 9 1 9 1 9 13 4 4 2
15 7 11 1 0 9 1 9 13 4 9 1 0 13 4 2
9 9 9 1 9 0 13 4 4 2
18 9 9 1 1 11 1 0 9 12 7 0 12 9 9 0 13 4 2
11 0 9 1 9 1 0 9 13 4 4 2
18 9 9 1 1 9 1 9 13 1 3 9 1 1 14 9 10 13 2
12 12 2 12 9 1 9 0 13 1 9 13 2
12 9 1 0 9 12 9 7 0 12 9 13 2
12 11 2 11 7 10 0 9 1 9 14 13 2
13 0 9 1 1 9 1 9 9 0 0 13 4 2
15 10 9 1 9 13 9 1 13 4 2 15 9 0 13 2
22 9 7 9 13 1 3 14 11 11 11 11 11 1 14 0 9 1 9 0 13 4 2
11 9 9 1 13 16 15 3 13 4 4 2
24 12 9 1 1 14 9 9 1 13 4 4 2 7 9 9 1 9 1 9 9 0 14 13 2
31 9 13 1 9 1 11 9 7 11 11 11 11 1 13 1 3 13 14 4 4 9 9 1 9 1 11 1 9 13 4 2
32 11 11 11 1 9 7 11 11 9 11 11 1 9 15 9 1 12 9 1 9 1 0 9 1 12 12 9 13 0 13 4 2
26 11 11 11 1 9 13 4 9 9 1 11 7 15 10 9 1 9 1 9 13 1 9 0 13 4 2
9 11 1 9 1 3 0 13 4 2
30 3 11 1 13 1 3 15 0 9 1 9 1 13 11 2 9 1 9 13 1 12 9 1 9 13 9 11 11 13 2
26 12 0 11 9 1 0 13 15 12 9 1 1 11 1 9 1 13 4 4 7 9 1 15 13 4 2
17 16 0 9 1 13 13 16 0 9 1 1 15 10 9 13 4 2
29 12 9 9 1 13 16 11 9 1 9 1 13 4 7 15 3 1 0 12 9 1 11 1 12 9 1 9 13 2
17 15 9 1 0 9 13 7 13 16 15 15 9 1 9 0 13 2
23 0 13 16 9 13 1 9 1 9 1 1 9 9 1 9 1 11 1 11 0 13 4 2
11 15 1 11 1 15 9 0 13 4 4 2
23 9 13 13 4 11 9 9 11 1 14 10 9 13 1 3 3 0 9 1 13 4 4 2
16 11 1 13 4 16 9 9 10 9 1 9 1 13 4 4 2
11 11 1 13 16 9 0 13 4 4 4 2
28 9 9 11 11 11 1 11 11 11 1 9 1 9 1 11 7 15 10 9 1 9 0 13 1 9 13 4 2
42 3 14 13 9 1 1 11 1 0 11 11 11 1 9 11 11 1 13 16 9 13 9 9 1 9 13 7 16 11 1 15 13 4 16 9 9 1 0 9 13 4 2
28 11 1 11 11 1 9 11 11 11 1 13 4 16 11 14 0 9 9 1 13 1 1 0 9 14 13 4 2
16 7 11 11 11 1 9 11 11 1 11 1 3 0 9 13 2
28 0 2 0 9 1 15 9 1 1 9 9 1 9 13 16 9 9 9 1 0 7 0 9 13 1 0 13 2
31 11 11 11 1 9 13 4 0 9 9 11 1 0 9 11 11 1 11 9 12 9 15 1 0 13 1 1 9 13 4 2
33 11 11 1 0 9 7 11 11 11 1 9 11 11 1 9 1 9 13 1 13 11 1 11 1 9 13 1 0 13 4 4 4 2
17 3 11 1 11 1 9 12 9 15 1 0 13 1 9 13 4 2
29 7 2 11 1 9 1 11 1 9 13 4 16 15 9 1 13 1 0 9 1 1 9 9 1 3 14 13 4 2
24 11 1 9 11 7 11 1 13 16 11 11 11 1 1 9 9 12 9 11 1 1 0 13 2
11 15 13 16 11 9 1 13 0 14 13 2
24 0 13 16 11 11 1 9 1 1 1 11 11 1 10 0 9 1 12 14 9 14 13 4 2
14 15 1 14 15 9 1 15 9 1 13 14 14 13 2
16 11 1 11 11 11 1 1 10 9 1 9 0 13 4 4 2
21 9 1 9 13 16 9 1 9 1 9 1 9 2 9 1 11 1 0 9 13 2
35 9 1 9 11 11 11 7 11 11 1 9 1 13 16 11 1 9 1 13 16 9 1 9 2 9 1 13 15 1 0 9 13 4 4 2
13 11 1 13 16 15 15 1 14 0 9 14 13 2
18 14 12 9 1 0 0 9 1 1 12 12 9 1 9 13 4 4 2
17 11 1 13 16 9 1 9 1 12 9 1 12 12 9 13 4 2
12 10 9 9 1 11 11 9 1 0 13 4 2
17 10 9 2 9 11 11 1 9 1 12 2 12 9 1 13 4 2
27 11 1 9 1 13 16 15 10 9 9 1 1 9 1 14 13 2 7 9 1 9 1 15 9 14 13 2
23 11 11 11 11 2 11 11 11 7 9 9 11 11 1 11 1 9 1 11 1 9 13 2
22 11 11 1 15 9 1 13 16 9 1 10 9 11 1 0 9 7 9 1 13 4 2
14 3 2 11 11 1 13 16 11 9 13 1 9 13 2
18 9 13 7 0 13 1 10 9 9 1 1 1 9 7 9 13 4 2
19 11 1 9 9 11 11 11 1 9 1 10 9 1 3 13 1 9 13 2
22 9 1 9 11 11 11 1 9 9 9 1 13 4 9 9 1 0 13 1 9 13 2
25 16 9 1 1 0 9 9 11 11 11 11 7 9 1 1 0 9 9 1 9 0 13 4 4 2
51 9 9 11 11 11 1 11 1 9 1 9 1 1 9 9 11 11 7 11 11 11 1 9 1 0 13 4 1 3 9 13 4 13 16 10 9 9 13 4 4 2 15 9 1 0 14 13 4 4 4 2
35 16 11 1 10 9 1 9 13 16 11 1 9 13 9 9 1 9 1 9 9 11 1 0 9 1 9 1 9 9 13 4 1 9 13 2
33 16 9 9 9 11 11 1 9 1 0 13 1 11 1 11 11 1 9 1 9 1 11 1 13 16 15 10 9 11 1 1 13 2
7 15 13 16 15 0 13 2
7 15 0 9 1 9 13 2
29 11 11 1 11 11 11 1 9 1 13 16 11 1 1 13 15 15 1 9 2 9 13 7 15 0 13 9 13 2
27 15 15 14 13 16 9 9 1 15 14 15 9 1 1 9 13 11 1 0 0 9 0 13 1 9 13 2
52 11 14 0 9 9 1 1 11 11 11 1 0 9 13 1 1 9 13 9 1 11 7 9 9 1 1 9 1 9 13 1 12 9 9 13 1 14 9 13 15 9 9 9 11 11 11 1 13 1 9 13 2
23 11 1 9 1 9 7 11 11 11 1 11 11 11 1 9 1 11 11 1 0 13 4 2
26 9 1 0 7 0 9 1 11 1 9 13 9 1 10 9 1 9 13 4 7 9 9 0 13 4 2
21 10 9 1 0 9 14 13 2 15 9 1 9 13 4 9 1 10 9 0 13 2
37 9 9 1 1 11 7 11 9 1 12 9 14 9 1 9 1 13 9 1 1 10 9 1 0 9 14 13 2 15 9 1 9 1 10 9 13 2
22 11 1 11 2 11 11 2 11 11 7 11 2 11 11 1 1 9 13 1 11 13 2
40 0 9 1 3 9 1 9 0 13 4 3 12 9 1 9 1 11 2 11 2 11 2 11 11 2 11 11 2 11 7 11 1 10 9 1 9 14 0 13 2
32 9 1 1 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 1 9 1 9 1 9 1 14 9 13 2
28 9 9 1 1 3 15 1 0 13 7 9 1 9 1 9 14 13 4 2 7 10 9 1 9 13 4 4 2
18 9 1 9 0 13 4 4 7 10 9 1 9 9 0 13 4 4 2
11 10 9 1 9 1 9 1 9 13 4 2
20 0 9 1 1 9 1 9 11 2 11 2 11 2 11 7 11 1 13 4 2
20 11 7 15 1 1 9 1 9 13 9 13 1 1 9 9 9 9 0 13 2
26 9 9 1 9 9 11 11 1 9 1 9 1 9 13 1 1 9 9 1 9 9 13 4 4 4 2
30 9 1 9 9 9 9 11 11 11 1 9 9 1 0 13 16 9 1 9 0 13 4 4 7 9 13 4 4 4 2
32 15 13 16 10 9 1 9 9 2 9 7 11 11 11 11 11 11 11 11 2 11 2 1 12 9 9 1 0 13 4 4 2
20 0 11 1 1 1 9 1 9 1 1 9 9 1 9 9 1 9 13 4 2
18 11 11 11 1 9 1 11 1 13 4 16 15 15 9 13 4 4 2
10 15 1 14 15 11 1 1 9 13 2
38 9 1 9 9 1 13 16 16 11 0 9 1 0 14 13 4 4 2 16 15 15 9 7 9 0 13 1 1 0 9 1 1 1 9 1 0 13 2
13 15 1 9 1 9 1 9 11 1 0 13 4 2
13 9 14 1 15 1 13 0 9 7 15 13 9 2
19 11 11 2 11 11 11 11 1 11 9 1 9 1 12 12 9 13 4 2
12 11 11 2 11 0 11 1 12 9 13 4 2
12 11 11 2 11 0 11 1 12 9 13 4 2
15 11 11 2 11 11 1 11 9 1 12 12 9 13 4 2
11 11 11 2 11 11 1 12 9 13 4 2
13 11 11 2 11 0 11 1 12 12 9 13 4 2
12 11 11 2 11 0 11 1 12 9 13 4 2
15 11 11 2 11 0 11 7 11 1 12 12 9 13 4 2
14 11 11 2 11 11 1 11 9 1 12 9 13 4 2
17 11 11 2 11 11 1 11 2 11 2 9 1 12 9 13 4 2
14 11 11 2 11 11 11 11 1 12 12 9 13 4 2
14 11 11 2 11 11 11 11 1 12 12 9 13 4 2
12 11 11 2 11 11 11 1 12 9 13 4 2
14 11 11 2 11 0 0 11 1 12 12 9 13 4 2
15 11 11 2 11 11 1 11 9 1 12 12 12 13 4 2
13 11 11 2 11 11 1 12 12 12 9 13 4 2
17 11 11 2 11 11 1 9 9 0 0 9 1 12 12 13 4 2
14 11 11 2 11 11 1 11 1 12 12 9 13 4 2
15 11 11 2 11 11 1 11 9 1 12 12 9 13 4 2
14 11 11 2 11 11 2 11 2 12 12 9 13 4 2
18 11 11 2 11 11 1 11 2 11 1 12 12 12 12 9 13 4 2
43 11 11 1 11 1 11 11 11 1 9 9 7 11 11 11 11 11 7 9 1 1 11 11 11 1 9 1 1 0 11 9 11 11 1 9 1 0 9 13 1 13 4 2
26 9 11 11 11 2 9 11 11 11 7 9 11 11 11 1 9 1 11 1 0 0 9 14 13 4 2
20 9 13 13 4 16 15 0 9 1 1 1 9 13 1 15 9 13 4 4 2
38 15 1 14 9 1 13 4 16 15 0 9 1 1 9 13 4 12 9 9 9 1 0 9 1 11 1 9 0 14 13 2 15 15 9 15 13 4 2
27 15 1 9 1 9 9 1 9 1 9 1 0 12 9 1 0 9 9 13 7 9 1 9 14 13 4 2
31 10 10 9 11 11 1 13 1 13 4 7 9 9 1 9 9 1 10 9 0 9 1 9 1 0 13 1 13 4 4 2
24 9 1 1 1 10 9 9 9 11 11 11 1 1 1 0 9 1 9 1 1 0 13 4 2
34 11 1 0 9 7 9 11 11 1 11 1 9 9 13 1 9 13 4 13 16 10 0 0 9 9 7 0 9 1 9 1 9 13 2
30 9 7 9 1 9 1 0 13 13 11 11 1 9 1 13 16 9 7 0 9 1 9 1 3 9 13 1 9 13 2
12 9 9 10 3 9 1 9 13 1 9 13 2
36 9 9 9 9 1 11 11 1 10 9 1 9 1 11 1 13 16 9 9 9 1 0 9 1 14 10 9 1 0 9 1 9 0 13 4 2
23 15 13 16 9 9 1 9 13 1 1 9 1 10 9 1 9 1 1 0 9 13 4 2
18 15 15 14 13 16 9 11 11 1 12 9 13 1 14 15 9 13 2
26 9 1 11 7 11 9 1 9 1 13 0 9 1 1 11 1 13 9 15 0 9 1 13 4 4 2
34 15 0 9 7 11 1 0 9 11 11 1 0 11 11 1 9 9 11 11 1 0 13 7 13 16 11 1 9 1 1 0 15 13 2
12 13 4 16 15 11 11 14 10 9 1 13 2
24 0 3 11 1 11 1 9 13 1 9 1 13 11 10 9 1 0 9 1 1 13 4 4 2
17 13 9 11 1 11 11 1 9 1 0 13 1 9 14 13 4 2
38 11 11 1 9 11 11 1 11 1 13 16 15 9 11 11 1 9 13 1 1 0 13 2 16 15 11 1 9 13 11 11 1 9 1 9 13 4 2
21 15 15 14 13 4 16 15 15 11 1 13 1 0 13 7 15 15 10 9 13 2
40 0 3 9 9 1 9 0 13 4 16 9 1 0 9 11 11 0 9 1 13 1 1 11 1 11 13 4 4 7 15 1 14 11 11 1 1 0 13 4 2
16 11 11 1 11 13 4 7 15 11 1 0 9 1 13 4 2
17 10 3 9 1 11 1 13 7 15 15 15 9 1 9 14 13 2
19 11 1 0 9 11 11 1 13 4 16 15 11 11 14 10 9 1 13 2
32 15 11 1 3 0 9 13 4 13 16 11 11 14 15 9 1 9 13 7 15 14 13 16 15 13 9 1 15 0 9 13 2
16 11 1 13 16 15 11 7 11 2 9 1 9 13 4 4 2
13 16 11 15 13 4 16 15 1 9 13 4 4 2
30 13 4 4 16 11 1 0 9 1 11 1 1 9 13 4 9 9 1 15 7 15 9 1 9 13 1 9 13 4 2
24 13 4 4 16 11 13 4 16 9 16 9 13 13 4 2 16 15 9 1 3 9 13 4 2
26 9 1 13 13 16 11 1 10 0 9 1 11 11 1 13 4 2 15 13 4 3 9 0 13 4 2
25 10 9 10 9 13 4 2 15 11 11 11 1 9 1 1 9 9 1 0 13 1 13 4 4 2
20 3 9 1 10 9 1 10 9 1 15 9 2 9 14 13 1 13 4 4 2
31 9 1 14 11 1 0 9 9 1 9 1 0 11 11 11 11 1 9 1 0 9 1 10 9 9 13 1 9 13 4 2
26 9 9 11 11 1 9 1 9 13 4 10 9 9 1 9 1 11 1 9 1 9 13 4 4 4 2
23 11 1 13 1 9 9 1 9 1 13 4 11 10 9 9 15 11 1 13 4 4 4 2
37 9 1 1 9 9 7 15 12 9 13 1 1 11 11 13 4 16 11 11 11 11 1 1 9 1 9 9 1 0 7 0 13 1 9 13 4 2
21 9 9 15 14 13 4 16 11 1 10 9 1 0 9 1 12 9 0 13 4 2
17 10 9 1 9 9 1 9 1 1 13 1 9 1 1 1 13 2
39 9 9 1 9 11 11 11 1 13 13 16 9 9 1 10 9 1 9 13 4 16 9 10 9 1 9 1 9 13 4 7 15 9 1 9 0 13 4 2
17 16 9 1 3 13 1 15 14 9 15 15 9 1 14 13 4 2
34 15 13 16 9 14 1 9 9 0 13 1 3 0 9 15 13 16 9 15 9 1 1 0 13 7 15 1 13 1 9 1 9 13 2
33 11 1 15 14 13 13 16 10 9 9 1 1 10 0 9 1 9 0 13 4 4 4 15 9 9 9 0 13 1 9 1 13 2
17 0 9 9 1 11 1 13 0 9 1 14 9 1 9 0 13 2
21 11 7 9 1 0 9 1 9 1 1 12 9 11 1 9 12 9 1 13 4 2
15 16 15 1 9 9 1 9 15 13 12 9 1 0 13 2
15 15 1 15 11 1 0 9 12 9 1 12 9 1 13 2
10 12 9 1 9 12 9 13 4 4 2
12 11 1 9 14 12 12 9 1 14 9 13 2
17 9 9 1 1 9 1 0 9 1 1 11 1 0 9 13 4 2
13 12 9 1 11 1 12 12 9 1 9 13 4 2
30 9 1 0 9 1 13 1 11 11 11 2 11 2 11 11 2 11 11 2 11 2 11 11 7 11 1 0 9 13 2
24 9 1 9 9 1 13 9 9 11 11 11 9 9 1 12 2 12 9 13 1 9 1 13 2
10 12 9 9 1 12 9 9 13 4 2
11 15 9 12 9 1 9 9 1 13 4 2
25 11 1 13 16 11 11 1 9 1 9 9 10 13 1 1 9 1 1 0 9 0 13 4 4 2
29 9 1 9 1 9 1 0 9 12 9 9 9 1 0 13 4 4 2 7 11 11 1 15 0 12 9 9 13 2
10 15 13 16 15 1 12 9 13 4 2
20 11 1 13 16 15 9 1 9 0 13 1 1 0 9 1 13 14 13 4 2
6 15 15 9 13 4 2
12 3 2 12 9 9 1 12 9 9 13 4 2
8 15 9 9 12 9 13 4 2
16 9 12 9 1 9 13 12 9 1 9 12 9 9 1 13 2
36 11 1 13 16 0 11 11 1 9 1 9 9 13 4 7 9 1 0 9 1 13 11 1 9 13 4 4 2 15 1 9 1 9 13 4 2
18 11 1 9 1 13 12 0 9 11 1 11 11 1 13 9 13 4 2
17 0 13 9 1 12 0 11 11 7 12 0 11 11 14 0 13 2
14 11 11 1 11 1 14 10 9 1 0 13 4 4 2
23 10 9 1 9 11 11 11 11 1 9 9 11 11 1 11 11 1 9 11 11 1 13 2
12 10 9 1 11 11 0 12 9 14 0 13 2
20 11 9 11 11 9 1 10 9 12 9 1 9 1 0 9 1 13 4 4 2
13 15 3 1 11 0 11 11 11 1 13 4 4 2
8 15 15 14 12 0 9 13 2
24 11 11 1 15 1 11 11 1 9 0 13 4 1 3 10 9 1 9 1 9 0 13 4 2
21 9 9 11 1 0 9 1 9 1 1 0 13 9 1 1 9 13 1 0 13 2
17 9 1 9 1 0 9 1 9 9 1 9 1 9 13 4 4 2
8 0 9 10 9 0 13 4 2
14 9 9 1 9 1 1 9 9 13 1 1 0 13 2
19 9 9 1 9 1 9 0 13 1 9 9 1 1 1 9 13 4 4 2
21 15 1 10 9 0 9 1 1 13 4 9 1 9 9 1 0 13 4 4 4 2
14 9 1 1 3 0 9 9 9 10 9 1 9 13 2
42 11 11 11 1 13 1 9 1 9 13 16 11 1 11 11 11 1 14 12 0 9 1 0 9 1 9 14 13 16 11 1 14 15 13 4 9 1 9 10 14 13 2
18 16 9 1 13 4 9 1 10 9 1 15 9 2 9 14 13 4 2
11 10 10 0 9 11 1 14 13 4 4 2
19 15 13 1 1 15 13 9 13 16 9 15 1 1 1 15 9 14 13 2
26 9 1 13 13 16 14 9 7 9 1 10 15 9 1 13 4 9 1 1 15 9 14 13 4 4 2
19 9 1 9 11 11 13 4 16 15 9 1 1 15 9 14 13 4 4 2
17 11 1 12 9 10 9 11 11 11 1 1 0 9 13 4 4 2
25 11 11 1 13 13 16 0 10 9 9 1 10 9 1 13 9 1 9 9 1 9 14 13 4 2
22 7 9 1 9 13 4 16 11 11 7 11 1 10 9 1 1 9 1 9 13 4 2
21 9 1 9 1 1 0 9 1 1 1 9 1 9 1 12 9 1 9 13 4 2
11 11 11 11 9 9 1 9 14 13 4 2
18 16 9 1 13 13 16 0 9 13 9 1 9 9 1 9 14 13 2
16 15 9 1 0 9 1 9 1 9 13 13 1 9 14 13 2
14 7 9 9 13 4 16 9 1 9 1 9 13 4 2
29 9 1 1 9 9 9 1 0 9 1 9 1 13 13 16 0 9 13 0 9 1 9 9 1 9 14 13 4 2
27 9 13 4 16 9 1 11 2 0 11 11 2 11 2 11 7 11 1 10 9 1 9 1 9 13 4 2
9 7 9 10 9 1 0 14 13 2
23 10 9 9 14 9 1 13 9 1 9 1 1 11 11 1 0 9 1 9 13 4 4 2
27 9 1 13 13 16 9 1 1 13 9 1 9 1 1 3 9 1 9 1 9 1 13 1 9 14 13 2
26 16 11 11 1 0 9 0 9 7 9 1 1 13 9 1 9 13 1 1 9 1 9 15 13 4 2
17 11 11 1 13 13 16 9 1 9 1 13 4 9 1 9 13 2
19 9 1 1 9 1 9 0 9 1 1 1 12 12 9 1 10 13 4 2
12 7 9 1 9 12 12 9 1 10 13 4 2
21 11 1 11 11 1 11 11 1 11 1 11 9 1 9 13 1 0 9 13 4 2
15 9 1 13 13 16 11 9 7 9 2 9 13 4 4 2
16 9 1 11 11 11 11 15 15 9 1 9 14 13 4 4 2
23 0 9 1 13 1 1 11 16 0 0 9 1 9 13 4 2 16 15 10 0 14 13 2
25 9 9 7 11 1 9 11 11 1 13 16 11 11 11 11 15 9 1 0 9 14 13 4 4 2
26 15 14 9 13 1 3 0 9 11 1 13 4 16 15 0 9 1 9 13 7 9 2 9 0 13 2
22 7 11 11 1 10 9 1 15 9 14 13 11 1 14 15 13 1 13 1 9 13 2
10 3 11 1 9 1 14 11 13 4 2
16 11 1 1 2 9 9 11 1 15 13 1 15 13 13 4 2
20 11 1 9 13 1 1 11 1 9 1 15 14 9 1 13 1 9 0 13 2
33 9 9 1 3 15 9 13 16 11 1 9 1 10 9 1 9 13 4 16 15 15 9 1 9 15 0 9 1 9 13 4 4 2
21 11 1 1 2 11 11 11 1 0 9 1 14 10 9 9 13 1 9 13 4 2
23 9 9 11 11 1 0 9 1 9 1 1 10 9 1 13 1 9 1 9 3 13 4 2
29 11 1 11 11 1 9 13 4 16 15 10 9 1 9 13 1 1 9 2 9 7 0 9 1 1 9 13 4 2
13 0 9 1 1 11 1 11 11 12 9 13 4 2
17 9 1 1 12 9 9 12 9 1 13 12 9 1 13 4 4 2
19 15 1 0 9 1 9 9 13 1 15 10 13 7 12 9 1 0 13 2
18 9 1 1 9 1 9 1 9 13 1 9 13 4 1 9 0 13 2
24 9 1 11 1 9 1 9 10 9 1 11 1 9 1 1 11 1 9 1 9 13 1 13 2
16 16 15 1 9 9 1 9 1 1 9 1 0 9 0 13 2
24 0 10 9 1 9 1 3 0 9 0 13 4 4 7 10 3 9 1 3 0 9 13 4 2
33 9 1 9 13 16 15 9 1 11 1 9 9 1 9 1 9 13 4 4 2 16 11 11 1 1 9 1 9 9 9 9 13 2
15 11 1 11 1 13 1 3 9 1 9 3 9 13 4 2
25 11 1 11 11 1 10 9 1 0 9 13 2 15 0 9 1 0 9 1 9 1 9 13 4 2
17 11 7 3 1 9 1 14 0 9 13 7 15 0 0 9 13 2
24 9 9 1 13 13 16 10 9 1 1 15 11 1 9 1 1 1 13 1 9 13 4 4 2
17 3 9 1 13 13 16 0 0 9 1 11 1 9 1 9 13 2
19 11 1 9 11 11 1 1 11 1 9 1 0 9 9 1 0 9 13 2
34 9 9 1 1 0 12 9 1 1 0 7 0 11 11 2 11 11 2 11 2 0 11 11 7 11 1 10 9 1 9 0 13 4 2
15 0 11 11 1 11 7 11 7 3 1 9 1 9 13 2
20 11 1 1 14 0 9 1 9 13 4 7 11 1 9 13 1 9 13 4 2
9 7 15 3 9 9 1 13 4 2
17 9 9 1 1 11 1 9 9 1 0 0 9 0 0 9 13 2
15 11 11 1 10 9 1 0 0 9 13 1 9 13 4 2
18 10 9 0 9 1 1 2 9 13 1 9 1 9 1 1 13 4 2
29 9 1 9 13 16 10 0 0 9 1 9 1 13 4 16 11 1 0 9 11 2 11 11 1 9 9 13 4 2
18 11 1 3 9 13 4 4 7 0 10 9 1 0 13 1 9 13 2
37 9 1 0 9 9 1 9 1 9 13 4 0 11 7 9 9 9 9 11 11 11 1 11 1 9 9 1 12 9 1 1 0 9 1 9 13 2
27 0 11 1 9 9 1 11 1 11 1 1 15 9 1 9 9 1 0 13 1 1 9 13 1 9 13 2
21 13 4 4 4 16 9 9 0 9 1 9 1 1 1 11 13 4 13 4 4 2
29 12 9 1 10 9 1 0 9 1 1 1 0 11 1 10 9 1 9 9 1 1 1 0 9 13 1 9 13 2
25 11 7 11 1 9 1 0 2 0 13 9 1 9 11 1 9 9 1 11 11 1 13 1 13 2
19 11 11 1 9 1 13 1 12 2 12 9 15 9 1 0 13 4 4 2
16 15 12 9 1 1 11 1 13 1 15 9 1 13 4 4 2
13 15 9 1 9 13 14 15 9 0 13 13 4 2
16 10 9 1 9 9 1 0 10 9 1 9 1 9 13 4 2
34 16 11 1 15 9 1 13 1 9 14 13 14 2 7 15 14 9 13 16 9 1 13 1 9 1 15 9 13 2 13 4 13 4 2
38 11 11 11 1 0 10 9 13 16 15 9 15 13 2 7 15 15 9 13 16 15 9 1 0 13 4 15 15 9 1 13 9 13 14 13 4 4 2
13 10 0 9 1 9 1 9 14 13 4 4 4 2
19 11 11 1 9 11 1 9 1 14 9 1 9 1 9 13 4 4 4 2
8 15 15 9 1 0 9 13 2
25 9 1 1 9 1 3 0 13 4 2 7 9 1 9 1 13 10 9 9 1 9 1 13 4 2
43 9 9 1 9 11 11 1 11 11 1 13 16 12 9 1 1 15 15 9 1 13 1 10 9 13 2 7 10 9 1 9 14 13 16 15 9 15 13 1 1 13 4 2
22 11 1 13 13 16 15 9 11 1 13 4 7 15 11 11 1 1 9 13 4 4 2
15 9 14 13 2 7 12 9 1 9 1 15 3 13 4 2
14 15 13 4 16 0 9 1 13 1 0 9 13 4 2
11 11 1 9 14 15 9 9 13 4 4 2
23 15 13 13 16 15 13 14 14 4 16 12 9 1 15 15 9 13 15 15 9 1 13 2
21 10 9 1 0 13 1 9 13 16 0 9 1 15 15 1 13 1 9 13 4 2
24 11 1 0 9 15 9 1 13 4 7 15 13 4 16 15 14 11 13 15 0 9 1 13 2
46 11 1 9 9 1 11 11 11 11 2 11 2 1 0 9 1 11 1 11 7 0 9 1 1 9 13 1 11 1 0 9 13 4 7 9 1 9 1 9 1 14 13 1 9 13 2
32 15 1 14 9 1 0 9 11 1 11 11 11 7 11 11 11 11 1 1 13 9 1 9 14 0 13 4 1 9 13 4 2
17 15 13 16 15 10 9 1 9 13 1 9 9 1 13 4 4 2
13 0 0 9 1 9 10 9 1 15 14 13 4 2
42 15 10 9 1 14 9 13 16 9 10 9 1 9 1 1 15 9 0 13 1 9 13 4 4 7 10 0 9 13 7 11 7 11 11 1 15 1 1 9 13 4 2
19 3 15 13 4 16 11 1 0 9 7 9 1 10 9 1 15 9 13 2
30 15 10 14 9 13 16 0 9 11 1 11 11 11 7 11 1 11 11 11 1 1 13 9 1 14 9 13 4 4 2
29 11 1 9 11 1 9 1 1 15 9 13 4 16 11 1 11 11 1 1 11 7 11 1 9 13 1 9 13 2
22 12 9 1 9 11 1 13 2 7 10 9 13 15 9 15 1 0 14 13 4 4 2
23 11 9 9 1 0 9 1 0 13 9 9 1 13 1 11 1 9 0 13 4 4 4 2
21 7 11 1 13 13 16 11 1 9 1 9 9 1 1 14 9 13 4 4 4 2
13 1 11 2 15 0 9 0 9 1 9 13 4 2
19 11 11 11 11 1 13 1 9 1 1 9 9 11 11 1 15 9 13 2
19 9 1 1 11 1 13 16 15 15 1 11 1 13 1 0 14 13 4 2
28 11 1 0 11 1 9 1 1 1 11 11 1 13 16 11 1 3 11 7 0 9 1 1 13 9 13 4 2
11 9 1 9 1 1 11 1 9 13 4 2
14 11 3 1 15 11 1 0 13 1 9 1 14 13 2
28 11 1 9 3 13 16 16 11 11 11 0 11 1 9 1 13 1 0 13 16 15 9 1 9 13 4 4 2
30 11 1 11 1 10 9 13 4 14 15 9 1 0 13 1 9 13 16 11 9 1 1 0 2 0 9 13 4 4 2
12 15 15 15 15 10 9 1 9 14 13 4 2
16 11 9 1 1 11 1 1 1 11 1 9 1 0 14 13 2
9 15 2 12 9 1 9 0 13 2
34 3 2 11 1 11 1 0 9 1 14 3 13 4 4 16 11 9 9 1 1 15 0 11 1 9 1 9 13 1 1 0 14 13 2
35 11 1 9 11 11 0 11 11 11 11 11 1 11 11 11 2 11 2 1 9 1 9 13 4 11 9 1 12 0 9 1 0 13 4 2
21 9 1 12 12 9 1 9 9 14 13 4 1 9 1 9 1 0 13 4 4 2
30 16 9 1 9 9 11 11 1 13 16 10 9 1 9 9 1 1 13 4 7 10 9 1 0 9 9 13 4 4 2
25 15 13 16 11 9 1 0 9 9 9 1 1 12 9 1 10 9 1 10 9 1 9 13 4 2
11 3 1 9 9 1 9 0 13 4 4 2
17 15 13 16 9 9 1 1 15 1 10 9 1 9 14 13 4 2
11 10 9 1 9 11 9 1 1 14 13 2
10 15 13 16 15 11 1 1 9 13 2
19 9 9 1 13 16 10 9 1 9 0 13 4 4 4 7 9 0 13 2
18 9 1 1 11 0 11 11 1 9 11 11 0 9 9 1 13 4 2
7 9 1 14 12 9 13 2
21 15 9 9 1 13 14 9 0 13 4 7 15 1 14 3 13 1 9 14 13 2
16 9 1 14 15 9 13 1 13 7 11 3 14 3 14 13 2
22 9 1 13 1 10 0 9 11 11 11 11 1 9 11 0 12 0 11 11 1 13 2
19 11 9 1 1 9 1 9 13 15 14 9 1 11 11 1 9 13 4 2
16 15 11 1 9 11 1 13 2 9 15 9 1 15 9 13 2
5 15 15 15 13 2
6 11 1 15 10 13 2
17 7 11 1 13 4 2 16 15 15 13 16 15 15 9 13 4 2
15 0 13 1 3 15 15 1 12 9 1 1 0 13 4 2
17 10 14 9 1 11 1 13 4 15 9 11 7 9 11 13 4 2
22 15 9 13 1 1 10 9 13 7 15 14 9 11 1 15 9 1 0 14 13 4 2
12 9 11 11 9 9 1 1 11 11 13 4 2
8 15 11 1 9 13 1 13 2
7 7 15 0 9 13 4 2
16 15 15 3 0 13 15 13 16 15 13 4 7 3 13 4 2
17 3 14 15 9 1 3 13 16 15 9 1 15 3 13 13 4 2
10 15 9 11 11 7 0 9 1 13 2
10 9 13 1 9 11 1 9 13 4 2
8 15 12 9 1 9 13 4 2
7 9 9 1 13 4 4 2
11 9 1 14 11 1 9 1 1 13 4 2
16 7 9 9 11 11 11 1 11 7 11 11 1 9 13 4 2
6 7 9 1 13 14 2
11 0 9 15 9 1 9 13 4 4 4 2
12 15 13 4 4 16 15 0 9 9 14 13 2
22 11 11 1 13 2 15 7 11 1 9 0 12 9 1 14 10 9 1 13 4 4 2
24 15 15 9 1 9 13 1 1 15 9 1 1 13 14 4 7 15 9 1 0 9 13 4 2
11 10 13 15 9 1 13 11 3 0 13 2
16 11 1 9 1 14 9 2 3 1 9 1 9 13 4 4 2
11 15 11 1 9 1 9 9 13 4 4 2
13 11 1 9 1 14 9 1 9 1 13 4 4 2
8 0 0 13 4 4 11 11 2
14 9 13 1 11 11 11 1 13 16 11 11 0 13 2
9 15 15 0 2 0 13 4 4 2
17 3 15 9 1 14 13 4 4 7 3 1 15 14 13 4 4 2
25 11 1 13 16 11 1 10 9 13 15 13 14 0 14 7 15 9 1 1 9 1 13 14 4 2
8 0 9 1 9 13 9 11 2
12 9 11 11 1 13 13 11 1 9 0 13 2
13 10 9 11 1 9 1 9 1 9 13 4 4 2
12 7 15 9 1 9 1 1 15 9 13 4 2
24 15 13 16 15 9 1 9 1 0 9 1 13 13 4 4 16 15 0 9 1 1 13 4 2
34 9 9 1 9 1 9 1 9 9 1 9 1 9 13 1 11 11 11 11 11 11 1 9 1 1 9 1 9 1 9 13 4 4 2
13 9 1 9 1 9 13 1 9 14 13 4 4 2
26 11 11 1 9 1 1 11 9 7 9 1 9 9 1 3 1 9 1 0 2 0 9 13 4 4 2
17 9 1 9 1 13 15 1 9 11 11 1 1 15 9 14 13 2
15 9 2 15 0 2 0 12 12 9 13 1 9 13 4 2
18 15 13 4 16 9 1 9 13 4 16 15 9 15 14 9 13 4 2
15 10 9 1 15 9 2 9 7 9 14 9 1 13 4 2
30 15 9 13 4 4 2 15 0 13 9 1 9 1 13 1 1 13 4 4 4 16 15 0 9 1 13 1 13 4 2
26 0 9 1 11 1 13 13 16 11 11 11 1 0 9 1 11 11 13 15 1 9 1 10 14 13 2
45 9 1 9 1 3 9 1 9 2 9 0 13 4 2 3 10 9 7 13 9 1 1 9 1 9 0 9 1 9 1 14 3 13 4 4 7 15 14 15 9 13 9 13 4 2
42 11 1 1 15 9 3 0 13 4 4 7 15 9 1 10 0 9 1 13 1 1 9 13 4 4 7 11 11 1 9 9 9 1 1 9 1 0 9 13 13 4 2
19 11 1 13 16 15 11 1 14 9 1 12 12 9 13 1 9 13 4 2
31 9 9 9 9 11 1 13 16 11 11 1 9 11 11 1 14 9 1 9 1 9 13 1 9 1 9 13 4 4 4 2
21 11 1 14 10 9 1 0 9 13 15 3 9 1 0 13 1 9 13 4 4 2
39 10 9 1 9 1 9 1 9 13 1 9 1 11 1 13 16 10 9 14 9 1 9 13 1 13 4 7 9 1 0 9 1 9 1 14 9 13 4 2
18 11 1 3 13 9 9 1 9 9 7 9 1 9 10 13 4 4 2
14 0 9 13 1 9 9 9 1 9 14 1 0 13 2
42 10 9 1 0 9 1 13 9 9 1 9 15 13 16 9 1 9 9 7 9 1 3 1 13 4 0 9 13 9 13 9 9 1 9 9 9 1 13 4 4 4 2
11 9 9 1 9 14 11 1 13 4 4 2
26 11 1 0 9 1 12 12 9 1 9 14 1 12 12 1 12 12 9 1 1 0 9 13 4 4 2
7 12 14 0 0 9 13 2
26 0 9 11 11 1 11 11 1 1 13 0 9 1 9 13 16 10 9 12 9 1 12 10 9 13 2
14 11 11 11 1 12 9 1 12 9 9 13 4 4 2
15 16 14 9 13 1 12 9 1 9 2 9 13 0 13 2
20 0 12 9 1 9 1 9 1 9 1 9 1 12 9 1 0 13 4 4 2
13 0 9 10 13 16 9 9 1 9 0 13 4 2
9 9 1 1 14 11 1 9 13 2
12 11 11 12 9 1 13 9 9 9 13 4 2
26 15 1 9 9 1 9 1 9 12 12 1 10 13 1 12 12 1 9 1 15 14 0 13 4 4 2
12 15 0 9 1 12 9 9 9 13 4 4 2
19 9 9 9 9 11 11 1 13 16 9 1 1 14 11 1 9 13 4 2
23 11 9 9 1 9 9 11 11 1 13 16 11 11 1 1 1 11 1 1 9 13 4 2
9 9 11 11 1 0 13 4 4 2
25 11 11 11 1 13 13 9 1 1 9 9 11 11 1 13 4 9 1 11 1 3 9 13 4 2
35 9 1 9 11 11 11 1 13 16 10 9 1 13 11 1 9 9 7 11 11 11 1 9 9 1 13 1 9 13 9 13 9 13 4 2
17 15 10 9 15 14 13 4 16 15 9 1 10 0 13 4 4 2
35 0 9 9 11 11 1 0 13 1 15 0 9 1 11 1 13 16 16 15 14 11 1 9 9 1 9 13 16 14 15 9 0 13 4 2
12 7 12 9 1 9 15 0 9 1 9 13 2
51 11 1 0 9 1 15 9 13 4 11 1 11 1 14 9 13 15 14 9 13 16 15 15 9 1 9 9 13 4 4 2 15 15 10 9 1 14 9 13 4 2 15 1 10 9 1 9 13 4 4 2
28 15 13 16 11 11 1 10 9 1 1 9 13 4 4 16 15 9 9 1 10 9 1 9 13 1 13 4 2
29 11 1 13 13 16 11 11 1 12 9 1 9 13 1 9 1 9 10 9 13 4 4 2 15 15 9 14 13 2
9 11 1 15 9 1 9 14 13 2
17 15 13 16 11 1 11 1 9 13 14 16 9 1 9 13 4 2
10 15 11 1 3 9 13 13 4 4 2
12 11 0 9 1 10 10 9 1 10 9 13 2
18 15 13 16 11 11 9 11 11 7 11 11 1 1 14 10 9 13 2
11 7 11 11 10 9 14 13 13 4 4 2
35 15 13 16 11 11 1 9 9 9 3 13 7 11 0 9 1 11 1 10 0 9 1 13 2 15 1 10 9 15 1 0 9 14 13 2
36 11 1 14 9 13 9 9 1 9 13 4 11 1 13 16 10 14 9 9 1 9 1 0 13 1 9 1 13 4 2 15 9 13 4 4 2
18 15 10 9 1 9 15 13 4 4 16 9 9 13 15 9 1 13 2
26 11 1 9 13 4 11 1 13 16 15 15 9 1 9 9 13 4 4 2 3 15 15 9 13 4 2
24 11 9 1 15 11 7 11 1 11 11 11 1 13 15 15 11 1 9 13 1 9 13 4 2
30 11 15 0 13 1 15 9 14 13 4 4 16 15 14 13 7 11 11 11 1 0 0 9 1 1 15 11 3 13 2
17 11 11 1 9 13 4 11 1 10 9 1 15 15 9 14 13 2
40 9 13 1 15 1 9 14 13 4 16 12 9 1 1 1 11 9 1 13 9 13 1 11 1 11 11 11 11 11 1 9 1 14 15 15 14 13 4 4 2
20 10 11 1 15 9 13 7 15 9 1 13 15 9 1 14 13 4 4 4 2
23 13 11 1 9 13 1 9 16 11 1 1 1 15 1 10 9 1 12 9 13 4 4 2
24 12 9 0 9 9 1 9 14 13 4 7 9 13 1 9 1 15 1 15 9 14 13 4 2
22 0 0 9 1 1 11 11 1 13 15 0 9 1 3 14 9 1 9 1 14 13 2
21 13 4 16 11 13 4 16 11 7 11 1 9 9 1 3 15 9 1 1 13 2
7 11 15 3 0 14 13 2
24 0 11 7 11 9 1 15 14 9 15 0 13 15 9 9 1 9 0 9 1 0 13 4 2
9 11 9 1 9 13 0 13 4 2
10 7 15 15 9 10 13 4 4 4 2
15 16 15 1 12 0 9 11 1 11 11 1 13 4 4 2
5 9 13 1 13 9
20 13 4 16 15 1 0 9 12 9 1 0 9 1 1 1 9 9 14 13 2
23 11 1 13 13 16 11 7 11 1 1 1 12 0 9 13 1 9 1 1 1 9 13 2
27 12 9 1 1 1 15 15 1 1 9 13 1 9 7 10 9 1 9 1 13 14 15 9 13 4 4 2
22 11 11 1 9 13 4 16 11 1 9 13 1 9 1 0 9 1 14 12 9 13 2
8 15 1 11 1 9 14 13 2
26 15 12 0 9 13 7 11 1 1 9 9 1 9 10 0 14 13 16 15 9 1 9 13 4 4 2
28 11 11 11 1 0 9 11 11 1 9 11 11 1 15 0 9 11 11 1 9 13 4 15 0 9 13 4 2
20 0 13 16 11 11 1 14 15 0 9 11 11 1 9 13 9 13 4 4 2
10 11 9 1 1 11 1 14 0 13 2
23 11 1 9 11 11 1 9 11 1 9 1 13 16 11 9 1 1 11 1 14 0 13 2
9 11 10 9 1 1 9 1 13 2
25 15 9 1 13 16 15 15 1 9 13 4 15 15 0 13 7 15 1 15 15 14 13 4 4 2
16 11 1 1 15 9 14 13 7 11 1 14 15 9 13 4 2
24 9 1 9 13 1 11 1 9 13 4 7 15 13 16 11 14 11 1 9 1 9 13 4 2
26 11 1 9 1 1 9 13 4 15 13 16 11 1 1 1 14 15 0 13 7 15 9 9 13 4 2
7 11 0 7 0 13 7 2
20 11 1 13 16 11 10 9 1 1 13 15 11 1 9 1 9 14 13 4 2
28 0 13 16 11 1 0 9 11 11 1 11 11 1 9 13 4 4 7 12 9 1 9 1 15 9 13 4 2
30 15 13 16 15 11 1 15 13 4 13 16 11 1 11 1 9 13 4 4 15 15 13 4 11 1 9 1 1 13 2
30 0 9 11 11 1 9 1 1 9 1 13 16 10 9 1 0 9 11 11 1 9 11 11 11 11 1 15 9 13 2
24 11 11 1 0 11 11 1 11 11 7 11 11 1 9 1 9 1 9 1 9 13 4 4 2
10 10 9 11 11 2 11 1 0 13 2
25 11 1 11 11 1 9 1 9 1 0 12 9 1 9 14 13 1 9 13 4 10 9 13 4 2
20 13 4 4 4 16 16 9 1 9 0 13 4 4 16 9 12 9 0 13 2
8 9 0 13 16 9 13 0 2
26 11 11 1 10 9 11 1 9 13 1 0 9 1 9 13 4 1 9 1 9 14 13 1 13 4 2
23 0 13 16 11 7 11 1 1 15 1 9 1 9 13 1 13 12 9 14 13 4 4 2
15 11 1 13 13 16 11 15 10 9 1 1 13 4 4 2
24 3 11 13 4 16 15 12 9 1 11 1 9 1 13 4 4 7 11 15 9 14 13 4 2
22 7 9 1 13 13 16 11 1 10 9 15 9 9 1 9 1 9 1 13 13 4 2
23 9 1 12 9 1 1 0 9 1 1 0 9 1 0 13 1 3 14 12 9 13 4 2
17 10 9 1 0 13 1 1 11 11 11 1 12 9 9 11 13 2
17 2 11 11 2 7 2 0 2 9 9 1 9 13 4 4 4 2
15 10 9 11 1 11 11 11 1 9 9 1 0 13 4 2
23 15 1 11 11 1 12 9 1 13 2 0 9 1 11 10 9 1 13 0 9 13 4 2
28 10 9 1 9 13 16 11 7 11 1 9 1 1 11 11 1 13 1 9 1 10 9 1 9 13 4 4 2
22 7 12 0 9 1 13 13 2 15 11 11 0 15 0 9 1 3 9 13 4 4 2
14 12 9 1 1 9 11 1 14 12 9 15 13 4 2
28 11 11 1 10 9 1 1 0 9 9 1 0 9 1 9 1 9 1 9 13 1 1 9 9 13 4 4 2
16 3 9 9 13 4 10 9 1 9 8 13 9 13 4 4 2
15 15 1 9 9 15 15 9 1 9 9 14 13 4 4 2
31 16 9 9 13 4 4 16 9 1 10 9 1 13 15 9 1 9 14 13 7 11 1 1 1 9 9 13 4 4 4 2
38 15 0 9 1 13 4 16 9 8 13 1 9 1 1 10 9 13 4 4 15 15 13 2 16 10 15 13 4 16 9 9 1 15 0 9 0 13 2
21 10 9 1 11 1 15 0 0 9 9 11 11 1 9 1 9 13 1 9 13 2
13 15 1 9 1 9 14 12 9 13 1 13 4 2
11 7 11 11 1 15 13 1 9 13 4 2
25 16 11 11 1 15 13 1 9 13 4 16 15 11 11 7 11 11 1 9 1 9 13 4 4 2
23 9 15 13 16 11 13 7 13 1 11 1 12 1 1 12 9 11 1 9 11 13 4 2
11 15 0 9 10 9 1 13 9 13 4 2
23 3 11 11 7 11 11 1 11 1 1 9 12 9 13 7 11 11 1 1 0 9 13 2
44 11 11 11 11 0 9 1 9 11 11 1 9 1 9 1 9 9 13 1 9 1 13 4 9 1 9 13 4 12 9 1 9 9 1 13 9 9 13 1 9 0 13 4 2
12 11 1 9 9 1 9 12 9 9 1 13 2
26 7 0 11 11 1 10 9 1 15 9 10 0 9 1 13 12 12 9 9 1 13 1 9 13 4 2
26 15 9 1 9 1 15 10 9 1 9 1 1 1 9 9 1 13 15 9 1 15 9 9 1 13 2
12 9 1 14 11 1 10 9 1 9 0 13 2
15 11 0 10 9 13 15 0 9 1 13 9 9 13 4 2
25 9 11 11 11 1 11 1 10 9 1 0 13 1 1 9 9 1 11 11 11 11 1 13 4 2
20 15 13 16 9 1 9 1 14 11 1 0 9 1 13 15 9 9 13 4 2
28 11 11 11 11 11 11 1 9 11 11 1 0 13 4 9 9 1 1 1 9 9 1 9 1 9 13 4 2
24 9 11 2 11 7 9 1 9 9 1 9 11 11 9 9 1 1 1 0 9 1 9 13 2
24 15 13 16 9 14 1 9 1 10 9 10 9 9 0 13 2 15 9 14 12 12 9 13 2
16 7 15 1 0 13 4 9 1 9 14 12 12 9 13 4 2
42 11 1 13 16 9 9 9 9 2 15 1 15 1 0 9 1 9 13 2 10 9 9 10 9 1 11 11 1 9 1 15 11 1 0 9 7 9 9 1 0 13 2
19 9 1 9 9 1 9 1 9 13 1 12 0 9 1 9 13 13 4 2
13 15 9 1 9 13 4 1 10 9 0 0 13 2
19 15 9 1 11 11 11 11 11 11 7 11 11 11 1 9 13 4 4 2
8 10 9 1 10 14 9 13 2
12 15 3 14 10 9 1 0 9 9 0 13 2
18 11 1 13 16 15 1 0 13 4 9 9 1 9 12 9 9 13 2
9 15 9 15 11 11 1 13 4 2
42 15 9 9 1 9 0 9 2 9 9 9 2 9 9 2 11 1 13 2 9 7 9 1 9 9 9 7 15 1 13 1 9 7 9 1 13 1 13 4 4 4 2
17 9 11 1 13 16 0 9 1 9 1 9 12 9 9 13 4 2
12 10 9 1 15 13 4 4 15 9 13 4 2
17 0 9 15 12 9 1 9 13 1 12 7 12 9 13 4 4 2
12 9 9 1 10 9 12 9 1 13 4 4 2
8 16 15 9 3 0 13 4 2
16 9 11 1 9 1 1 1 9 9 1 0 9 1 0 13 2
22 15 3 0 9 15 13 16 0 9 13 4 7 15 9 1 9 14 3 3 13 4 2
25 11 1 10 0 9 1 9 9 9 1 9 1 1 11 1 11 11 11 11 11 1 11 11 13 2
15 11 7 0 11 11 11 1 1 11 7 11 1 9 13 2
28 9 13 1 3 11 1 9 1 13 16 15 11 11 7 15 1 9 1 1 1 11 1 11 1 9 13 4 2
22 15 13 16 15 0 11 1 13 1 1 0 13 7 15 1 9 13 1 3 14 13 2
20 11 1 13 16 15 0 9 1 9 1 9 13 1 9 1 3 13 4 4 2
16 15 13 16 11 2 11 1 1 10 0 9 1 14 9 13 2
20 13 4 4 4 16 11 14 10 9 1 1 11 1 0 0 9 1 9 13 2
26 3 11 14 9 1 1 9 9 1 9 1 10 13 7 9 1 0 9 1 0 13 1 9 14 13 2
25 11 1 13 4 16 11 1 11 13 4 1 9 1 14 11 1 1 0 9 1 9 0 14 13 2
10 15 0 9 1 12 9 14 14 13 2
17 2 16 2 11 1 11 1 11 9 11 11 11 11 1 9 13 2
17 12 9 1 13 15 9 1 0 9 1 10 9 1 14 9 13 2
30 11 1 11 11 11 11 11 1 12 9 1 9 1 13 16 11 9 1 10 14 9 13 15 11 1 9 1 0 13 2
16 11 1 13 16 10 9 1 15 15 1 9 13 1 0 13 2
34 11 1 13 13 16 12 9 1 1 0 9 7 9 13 1 11 3 14 13 2 7 11 1 9 1 11 15 0 9 1 3 14 13 2
31 3 11 1 11 15 11 13 15 11 1 11 9 1 11 0 9 1 12 9 1 9 13 4 7 12 9 1 0 13 4 2
20 7 11 11 11 11 1 0 9 1 1 0 7 0 9 13 1 9 13 4 2
38 0 13 16 11 1 9 1 11 1 9 11 1 1 1 0 9 9 1 13 4 4 0 9 1 1 15 1 14 12 1 10 9 1 9 13 4 4 2
17 11 1 9 9 1 13 13 4 9 9 1 9 1 9 13 4 2
20 10 9 1 0 9 9 1 1 9 1 13 4 7 9 14 9 9 13 4 2
12 9 1 1 12 9 9 13 3 9 13 4 2
15 9 1 3 1 9 1 9 13 1 9 1 14 3 13 2
10 11 7 9 1 14 9 1 9 13 2
35 10 3 9 1 12 0 9 7 12 9 1 9 1 9 9 13 4 16 3 9 13 4 11 1 9 1 12 9 7 10 9 9 13 4 2
20 9 2 9 7 9 1 12 9 9 1 9 13 16 9 7 9 14 0 13 2
10 9 1 9 9 1 1 14 9 13 2
16 3 1 9 0 13 13 9 14 9 1 9 1 9 13 4 2
12 16 15 15 1 9 1 9 1 9 13 4 2
13 9 1 9 9 9 1 1 0 9 9 1 13 2
14 9 14 12 9 0 9 11 11 3 1 13 4 4 2
11 15 15 0 9 1 1 9 13 1 13 2
10 10 9 1 12 9 1 9 13 4 2
21 11 1 1 10 3 9 1 9 1 1 0 9 1 9 13 7 9 1 9 13 2
13 15 1 12 9 1 14 9 13 9 13 4 4 2
7 11 0 9 13 9 13 2
22 15 0 9 1 1 12 9 9 1 13 7 15 0 9 1 9 1 13 9 1 13 2
13 15 1 9 1 15 9 9 1 15 13 1 13 2
16 11 9 9 1 15 13 16 15 15 9 1 9 13 4 4 2
10 9 0 13 1 3 15 15 9 13 2
11 15 1 15 0 9 1 13 1 13 4 2
30 15 1 9 9 1 9 1 9 13 2 15 9 1 9 1 9 1 9 13 7 9 1 0 9 14 13 1 9 13 2
18 15 1 9 1 12 9 9 1 1 13 7 11 11 1 9 13 4 2
27 10 3 10 9 1 3 0 9 1 9 9 2 11 2 11 11 2 11 2 1 13 4 7 9 13 4 2
15 9 13 14 4 4 16 9 9 9 15 9 1 15 13 2
16 15 9 1 13 13 7 0 9 15 14 13 1 0 14 13 2
9 10 9 1 15 1 9 14 13 2
12 15 1 13 9 9 9 1 9 13 4 4 2
8 10 3 11 1 9 15 13 2
11 9 1 9 1 9 1 9 1 9 13 2
21 9 12 9 9 9 7 9 14 13 16 3 0 9 1 11 13 9 13 1 13 2
15 3 1 11 1 13 4 1 3 9 3 2 3 13 4 2
24 10 9 1 11 11 1 9 13 7 0 9 1 1 0 12 0 9 9 1 9 13 4 4 2
23 9 9 10 9 7 9 1 1 9 1 1 11 11 1 9 9 13 7 9 0 13 4 2
39 11 11 1 9 1 9 1 0 13 4 0 9 9 11 11 11 11 2 11 2 1 9 1 0 9 1 12 9 3 11 11 1 11 11 1 9 13 4 2
31 11 11 11 11 2 11 11 11 11 11 7 11 11 11 1 9 1 13 9 1 11 1 9 1 9 1 9 1 9 13 2
28 9 1 9 13 16 10 9 2 11 11 2 0 13 16 15 9 1 1 14 9 14 1 0 9 14 0 13 2
42 11 11 11 11 1 9 11 11 11 1 13 16 9 0 9 1 12 9 1 13 4 9 1 10 15 9 14 13 4 15 9 7 9 1 0 9 9 1 9 13 4 2
9 11 1 9 1 9 0 13 4 2
35 0 9 1 13 0 9 1 13 4 0 9 9 11 1 9 9 11 1 11 1 0 9 9 12 13 12 9 1 11 11 11 1 9 13 2
15 11 11 11 11 1 0 9 1 1 11 1 9 13 4 2
23 15 13 16 15 11 1 10 9 1 1 1 9 1 9 7 9 1 9 1 9 13 4 2
8 9 9 1 12 9 9 13 2
9 10 9 12 9 1 9 1 13 2
18 12 9 1 13 11 9 1 1 15 0 9 9 1 15 0 9 13 2
18 11 11 11 11 2 11 2 1 1 9 7 0 0 9 13 13 4 2
30 11 9 1 9 13 4 10 9 11 1 9 9 1 9 1 10 9 13 4 2 16 9 1 10 14 10 13 4 4 2
34 10 9 1 13 1 9 9 13 2 9 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 9 11 11 7 11 1 11 11 2
19 9 1 1 9 9 1 9 7 11 7 11 1 9 1 9 14 0 13 2
26 10 9 1 1 9 11 11 7 15 9 9 1 9 9 1 9 7 15 9 1 0 9 1 9 13 2
26 15 9 1 9 1 13 4 9 9 1 11 1 13 1 1 12 0 9 9 11 1 0 13 4 4 2
19 11 11 11 1 9 1 0 0 9 1 1 15 1 9 1 9 9 13 2
12 15 9 1 14 12 9 1 0 9 0 13 2
18 15 1 12 9 1 10 9 9 1 1 0 9 1 1 9 13 4 2
11 15 1 9 1 9 1 9 13 9 13 2
18 0 0 9 9 9 1 9 1 9 1 9 1 9 1 1 13 4 2
14 10 0 9 1 9 9 1 10 9 1 9 13 4 2
23 9 1 11 1 11 11 11 11 1 13 16 11 1 11 1 0 0 9 1 9 13 4 2
28 11 11 1 11 1 13 4 16 11 1 9 11 2 11 9 1 9 9 1 9 13 0 9 1 9 13 4 2
19 15 13 16 9 1 12 9 9 1 12 0 9 1 9 1 9 13 4 2
27 11 11 1 11 11 1 12 9 1 9 9 11 11 1 9 9 13 1 9 1 9 13 1 9 13 4 2
29 11 1 9 0 0 9 11 11 11 1 13 16 9 1 9 11 1 9 1 9 1 9 13 1 9 13 4 4 2
23 11 1 0 11 9 1 11 9 9 1 11 1 13 9 9 1 12 9 1 9 13 4 2
15 9 1 12 9 7 12 9 1 12 9 0 13 4 4 2
20 9 9 1 1 9 1 1 0 9 9 1 1 12 9 1 9 1 9 13 2
22 15 13 16 0 9 1 9 1 9 13 1 3 9 1 9 13 13 1 0 13 4 2
18 0 9 1 9 1 1 11 11 11 11 1 9 13 1 9 0 13 2
13 10 9 1 11 1 0 9 1 0 13 4 4 2
15 9 9 1 1 9 1 9 9 1 15 9 14 13 4 2
34 11 9 1 10 9 0 9 1 13 1 11 1 1 0 9 1 9 13 4 1 9 1 11 11 11 11 1 1 9 0 13 4 4 2
23 11 2 11 11 1 0 9 1 9 9 1 9 1 9 1 9 13 1 9 13 4 4 2
19 9 11 11 11 1 9 1 11 1 9 1 1 9 1 0 13 4 4 2
32 11 1 9 1 0 9 1 9 9 2 9 1 0 9 2 9 9 1 9 2 9 7 9 1 14 9 1 0 13 4 4 2
32 9 1 9 13 4 4 16 9 9 1 0 11 13 4 1 11 1 0 9 1 9 1 13 1 0 9 1 9 0 13 4 2
15 12 0 9 1 11 1 0 9 1 9 13 1 9 13 2
26 11 9 1 9 1 0 0 9 1 1 13 9 1 9 1 11 1 12 0 9 1 0 13 4 4 2
34 11 1 9 9 9 11 11 11 1 13 16 0 9 1 0 9 1 13 9 1 1 1 11 11 11 7 11 11 1 0 13 4 4 2
30 11 1 13 16 11 9 9 1 1 11 1 0 13 4 9 9 11 11 1 13 9 1 1 1 9 1 0 13 4 2
13 15 13 16 9 1 1 1 10 0 9 13 4 2
23 11 11 1 9 1 9 1 13 11 7 11 9 1 9 1 0 9 1 15 9 14 13 2
31 15 12 9 15 9 9 11 1 9 1 10 9 13 4 4 16 15 11 9 1 9 1 9 7 9 1 9 0 13 4 2
9 3 15 10 10 0 9 14 13 2
13 16 10 9 13 15 11 1 1 9 14 13 4 2
26 7 12 9 11 1 9 13 4 4 15 15 0 9 1 9 1 9 7 9 1 1 9 13 4 4 2
24 10 3 11 11 1 13 16 11 11 1 13 12 2 12 9 1 11 11 14 9 13 4 4 2
38 9 11 1 2 9 1 2 9 1 9 1 9 1 0 9 9 1 10 9 10 9 13 4 4 2 15 15 11 11 1 9 13 1 9 9 13 4 2
45 15 0 9 13 16 11 1 13 1 9 2 9 9 1 0 9 1 11 1 10 9 1 3 9 13 4 2 7 9 1 15 13 9 13 1 9 13 16 10 15 9 13 14 14 2
18 3 11 1 9 14 14 13 4 16 9 1 9 10 9 9 13 4 2
15 11 1 9 9 1 2 0 2 11 1 9 13 14 4 2
27 15 1 2 9 1 1 3 0 9 1 1 13 4 1 11 1 13 2 15 15 9 13 1 9 14 13 2
12 7 15 0 13 16 15 9 1 9 13 4 2
19 15 15 14 13 16 0 9 9 1 10 9 13 4 4 2 15 0 13 2
14 11 1 11 1 9 1 9 1 14 9 0 13 4 2
24 15 13 16 11 1 10 9 9 1 1 14 9 9 1 9 9 1 1 2 0 7 0 13 2
8 15 13 1 0 9 13 4 2
8 9 15 9 13 13 4 4 2
38 10 9 1 1 11 9 0 9 1 9 11 11 7 9 9 11 1 1 9 9 1 15 9 7 9 1 1 0 11 11 9 1 9 1 9 13 4 2
21 3 1 15 1 1 11 15 13 9 13 1 9 13 16 10 15 9 13 14 14 2
20 9 1 9 1 11 3 2 3 13 4 16 11 14 15 0 9 13 4 4 2
19 15 13 16 9 1 10 9 7 9 11 11 0 9 9 1 9 13 4 2
19 11 1 9 9 1 1 9 13 4 7 9 15 15 0 13 4 4 4 2
34 0 13 16 11 9 2 9 1 1 0 9 1 1 9 1 0 13 1 11 1 9 13 4 11 11 9 1 1 9 1 9 13 4 2
19 12 0 9 1 9 1 10 9 13 4 7 3 1 0 9 1 13 4 2
35 11 11 1 11 1 9 1 11 1 1 1 9 9 13 1 9 1 1 9 1 9 11 11 1 11 1 9 9 11 11 1 12 9 13 2
32 15 11 1 11 1 11 11 11 1 11 11 11 11 1 0 13 4 10 9 1 9 1 9 1 13 4 1 9 13 4 4 2
47 9 1 11 1 1 1 13 9 1 13 4 4 16 15 11 1 11 11 1 0 2 9 1 9 1 11 7 0 11 11 11 11 11 1 9 13 0 10 0 9 13 15 11 13 4 4 2
35 10 9 1 9 1 11 1 11 1 15 9 1 9 9 1 9 13 4 13 16 9 1 10 9 1 0 7 0 9 2 9 13 4 4 2
15 15 1 0 13 16 10 9 1 9 1 9 1 13 4 2
25 10 3 9 1 11 1 9 9 11 11 11 1 13 16 9 1 12 9 1 9 9 0 14 13 2
21 15 13 16 11 1 9 10 9 1 0 9 0 13 1 1 11 1 9 1 13 2
29 0 13 16 9 7 9 9 1 14 11 1 11 9 1 11 1 13 4 1 9 9 1 9 1 0 9 13 4 2
25 9 1 9 9 13 1 1 9 13 1 0 9 13 4 4 7 15 1 15 11 1 9 13 4 2
41 10 9 0 9 1 0 9 11 1 9 1 0 9 1 9 13 1 12 2 12 12 9 1 9 13 0 9 9 11 11 1 1 10 9 1 9 0 13 1 13 2
21 9 1 0 9 1 9 9 1 9 9 0 13 1 9 13 1 9 14 13 4 2
31 11 1 9 1 9 1 11 9 11 11 1 13 16 9 9 1 9 0 13 1 9 13 0 9 1 9 13 4 4 4 2
26 7 15 10 9 1 0 13 16 11 11 11 11 11 2 11 2 1 15 1 0 9 0 13 4 4 2
48 9 9 1 0 13 4 11 11 1 13 16 11 13 1 15 0 9 10 15 14 13 4 16 15 9 1 12 9 1 16 11 11 1 15 9 0 13 4 7 9 0 13 9 1 0 9 13 2
16 15 13 16 9 0 13 4 2 15 1 15 3 10 9 13 2
36 11 1 13 16 10 10 12 2 12 12 9 15 9 9 1 10 1 9 13 4 2 1 11 11 1 1 9 9 0 13 1 1 9 13 4 2
37 9 9 1 13 10 9 1 1 1 9 13 4 11 11 1 13 16 12 9 7 9 1 12 9 1 1 12 12 9 1 10 1 9 9 13 4 2
27 15 13 16 10 9 0 12 9 1 1 12 9 1 9 9 1 1 12 12 9 1 14 10 1 9 13 2
18 11 1 13 16 10 3 12 12 9 1 10 1 12 9 9 13 4 2
10 10 10 9 9 9 1 13 4 4 2
23 15 13 16 9 9 13 1 12 9 1 12 9 1 12 12 9 1 9 1 9 13 4 2
10 7 10 9 0 9 1 3 10 13 2
33 11 1 0 9 1 9 9 0 13 1 1 9 1 9 13 4 11 1 13 16 15 15 11 11 1 11 11 13 15 8 0 13 2
13 16 3 1 15 15 8 0 13 15 14 13 4 2
14 7 9 1 0 13 1 9 1 15 10 9 13 4 2
18 11 11 11 1 9 9 9 11 11 1 15 9 1 9 13 4 4 2
20 0 0 9 11 1 9 1 9 13 4 9 9 13 1 10 9 13 4 4 2
16 11 1 13 16 15 1 9 9 9 13 1 10 0 9 13 2
20 11 1 13 16 15 9 1 0 13 4 4 16 15 1 9 9 3 0 13 2
16 16 15 10 9 1 9 13 16 15 9 9 1 1 1 13 2
31 11 1 13 16 15 9 1 10 9 1 13 1 1 15 9 1 13 1 9 13 4 7 15 9 1 9 13 4 4 4 2
19 11 1 13 16 15 15 9 1 9 1 9 9 11 11 1 14 9 13 2
12 15 13 16 15 11 1 9 9 1 0 13 2
20 11 1 13 16 15 10 9 1 0 9 1 9 13 7 9 13 4 9 13 2
13 11 1 11 2 11 1 0 9 1 9 13 4 2
22 11 11 11 1 9 9 1 0 9 1 9 13 4 15 9 1 13 4 1 13 4 2
12 15 1 0 13 16 9 9 1 9 13 4 2
15 11 11 1 9 1 11 1 11 11 11 1 9 13 4 2
14 15 9 9 1 9 7 9 1 0 9 1 9 13 2
15 15 0 9 1 0 9 1 1 9 13 4 1 9 13 2
24 0 12 9 1 9 9 1 9 9 12 9 1 13 4 12 9 13 4 1 11 3 0 13 2
43 11 1 13 16 11 1 9 1 10 9 13 4 13 15 1 11 11 1 11 11 11 2 11 2 1 9 9 1 9 1 9 13 4 4 7 10 9 1 9 13 4 4 2
36 11 11 11 11 1 9 1 10 9 9 9 9 1 9 1 13 9 13 7 15 9 13 1 3 14 0 13 0 9 0 13 1 1 9 13 2
21 11 1 10 9 1 0 0 9 1 1 2 11 11 11 2 0 13 1 9 13 2
16 15 9 9 1 9 1 9 13 4 15 0 13 1 9 13 2
12 11 1 9 9 9 1 9 1 14 9 13 2
17 15 13 16 9 2 9 7 0 0 9 1 9 13 1 9 13 2
42 15 13 9 1 0 9 0 13 1 1 11 11 11 11 11 1 9 1 1 2 9 11 11 7 11 11 11 11 11 1 1 0 9 1 15 9 1 9 13 4 4 2
9 15 9 9 1 9 1 9 13 2
12 3 1 11 7 11 1 9 1 13 9 13 2
15 9 1 13 16 9 9 1 9 1 9 10 13 4 4 2
28 15 1 9 1 10 9 2 0 0 9 2 9 1 9 2 9 1 10 9 9 7 9 1 10 9 13 4 2
31 11 9 1 9 13 1 11 11 1 9 1 9 3 13 4 4 7 12 9 15 0 9 1 15 9 1 1 13 4 4 2
18 7 9 1 10 9 1 11 1 12 12 9 1 10 1 9 13 4 2
13 11 1 12 9 1 13 4 12 9 3 13 4 2
17 9 1 9 13 12 0 9 3 14 11 1 0 9 1 9 13 2
14 11 1 1 13 11 9 1 9 1 0 9 13 4 2
22 9 1 0 9 1 12 9 2 9 9 7 9 1 9 2 9 1 9 13 4 4 2
10 9 11 7 11 9 1 9 9 13 2
10 11 1 11 11 11 0 13 4 4 2
22 9 1 0 9 1 1 12 9 1 13 11 9 1 12 12 9 1 9 13 4 4 2
12 12 0 9 9 1 9 1 13 4 4 4 2
16 10 9 1 1 1 9 9 1 13 11 1 1 13 4 4 2
19 11 1 9 1 1 11 9 1 14 11 1 1 12 0 9 13 4 4 2
12 11 9 1 12 9 1 0 9 9 13 4 2
25 11 11 11 11 11 11 1 11 1 11 11 1 13 16 11 1 13 3 9 1 15 9 14 13 2
21 15 15 0 13 4 4 16 11 9 1 9 13 1 1 14 15 9 11 1 13 2
12 11 1 9 1 0 3 11 1 9 11 13 2
8 15 15 15 0 13 4 4 2
14 15 1 12 9 1 9 13 11 1 9 1 13 4 2
24 9 1 12 9 1 11 9 1 11 7 11 11 9 1 12 9 1 12 9 1 13 4 4 2
17 0 11 2 11 11 1 13 12 0 9 1 13 1 9 0 13 2
43 9 1 13 13 16 11 1 9 1 0 9 1 13 4 10 0 9 1 14 13 4 4 4 16 11 1 9 15 0 13 4 4 2 16 10 9 1 9 3 13 4 4 2
9 15 3 9 1 9 13 4 4 2
23 9 9 9 1 13 13 16 10 9 1 9 9 9 13 1 3 14 15 13 4 4 4 2
22 9 1 0 13 9 1 11 1 11 1 1 11 11 11 11 11 1 9 1 9 13 2
9 10 9 1 9 9 2 9 13 2
19 3 11 1 12 12 9 1 14 10 9 7 9 13 1 9 0 13 4 2
22 0 9 1 1 11 11 1 9 9 12 9 1 14 11 1 11 9 1 13 4 4 2
11 3 9 1 9 1 9 13 9 13 4 2
19 15 1 13 4 9 9 1 9 1 9 9 1 13 9 1 0 9 13 2
7 7 10 9 3 13 13 2
9 9 1 15 1 15 9 14 13 2
30 11 9 1 11 9 1 9 9 9 7 9 9 9 1 13 12 0 9 1 1 13 9 1 12 9 1 13 4 4 2
13 13 4 12 9 11 2 11 2 11 1 0 13 2
21 15 1 9 11 1 11 1 13 1 13 2 15 9 11 11 1 1 1 13 4 2
9 0 9 11 1 14 13 4 13 2
10 15 9 11 11 1 1 1 13 4 2
13 9 1 9 9 9 1 9 11 11 0 13 4 2
11 11 1 9 1 12 9 0 9 0 13 2
21 9 1 9 11 11 11 11 2 11 1 12 9 9 1 9 13 1 9 0 13 2
26 9 11 11 11 1 13 9 1 9 1 9 9 9 1 1 0 11 11 11 1 12 9 1 9 13 2
8 15 1 12 9 0 9 13 2
22 15 1 10 9 1 0 9 1 0 9 1 9 1 1 14 12 9 9 0 13 4 2
13 10 9 1 9 1 12 9 1 0 14 13 4 2
60 0 13 4 9 1 11 11 2 15 0 9 1 9 9 13 4 4 1 12 9 2 9 1 12 9 1 12 9 7 12 9 2 12 9 9 9 7 12 9 0 9 1 9 2 15 15 9 1 9 1 9 14 13 4 4 2 0 13 4 2
14 9 1 9 1 9 11 11 11 1 0 13 4 4 2
7 15 9 11 1 9 13 2
40 10 9 9 1 10 9 7 9 13 15 0 9 1 11 11 1 11 11 11 2 11 11 11 11 1 11 11 7 11 11 1 11 11 11 11 1 9 14 13 2
20 11 11 7 11 1 10 9 1 15 15 14 9 1 9 13 1 9 13 4 2
24 11 11 1 9 1 11 1 11 1 11 11 11 11 1 9 13 1 10 9 3 13 4 4 2
46 11 11 1 9 1 1 11 1 12 10 0 9 11 11 11 1 13 4 16 11 1 11 1 9 11 1 11 1 1 0 9 1 1 9 9 7 9 1 9 1 1 1 9 13 4 2
27 0 9 13 1 1 0 9 1 14 9 9 1 9 13 1 9 1 1 11 1 12 10 0 9 13 4 2
29 11 1 1 11 1 0 9 9 11 11 11 1 0 9 1 9 1 1 15 1 12 2 9 2 1 9 13 4 2
39 0 9 11 11 1 12 9 1 9 9 11 1 11 1 9 2 11 11 2 1 13 16 11 1 9 1 9 1 0 9 1 0 9 1 9 0 13 4 2
21 11 1 13 16 11 1 9 1 1 13 1 9 1 11 1 10 9 1 13 4 2
17 11 1 9 1 1 15 9 7 9 13 10 9 1 13 4 4 2
32 15 13 16 11 1 0 9 11 9 13 1 3 15 11 1 3 15 13 2 15 14 15 0 9 1 1 10 9 1 13 4 2
17 0 13 16 11 1 9 1 9 1 9 13 4 7 9 13 4 2
13 11 11 1 9 0 11 11 9 1 9 13 4 2
9 11 1 11 11 1 9 13 4 2
17 11 11 1 9 1 11 11 1 9 1 0 13 1 0 9 13 2
13 15 1 0 9 1 11 11 1 9 1 9 13 2
30 16 11 1 9 1 1 9 1 9 13 4 7 0 9 1 1 12 1 1 12 9 1 11 1 9 1 0 13 4 2
20 0 11 11 11 11 1 9 9 13 16 9 1 11 11 11 1 9 14 13 2
26 9 9 9 1 1 0 9 9 1 11 1 13 16 15 7 9 1 10 0 0 9 1 9 14 13 2
25 15 13 16 16 9 1 9 9 13 4 4 4 7 11 1 0 9 1 9 13 1 9 13 4 2
9 15 0 9 7 9 13 0 13 2
16 9 1 10 9 15 14 9 7 9 1 0 9 14 13 4 2
26 15 13 16 11 9 1 9 14 13 4 7 15 10 9 13 15 15 0 9 9 1 1 14 13 4 2
10 11 11 1 9 1 11 1 9 13 2
22 15 13 16 9 1 9 15 14 9 13 4 7 10 9 1 15 9 0 14 13 4 2
12 9 1 9 9 9 1 14 9 1 9 13 2
14 15 13 16 0 9 1 9 1 0 9 0 14 13 2
23 9 1 9 1 9 1 15 13 16 3 15 11 1 0 9 13 4 7 15 9 13 4 2
12 11 3 0 13 7 9 1 3 0 13 4 2
23 15 13 16 11 1 11 1 9 1 9 13 10 9 0 14 0 0 9 1 9 9 13 2
21 15 13 16 9 1 10 9 0 13 7 9 13 16 11 12 9 3 9 1 13 2
22 11 1 13 16 11 1 9 7 9 1 1 10 9 13 4 2 15 12 0 9 13 2
13 15 3 0 13 7 0 11 1 9 1 0 13 2
20 11 11 11 1 9 13 4 15 13 16 0 9 1 0 9 1 9 13 4 2
18 15 0 13 16 9 1 13 4 14 0 9 1 9 1 9 13 4 2
32 11 1 9 1 9 1 1 0 9 1 9 11 11 11 1 0 13 1 1 11 9 1 15 9 9 1 1 1 13 4 4 2
32 11 1 9 7 0 9 9 11 11 1 9 1 13 4 16 11 1 0 11 1 9 1 9 13 4 4 7 15 11 9 13 2
16 10 9 1 1 11 11 1 12 9 1 0 14 13 4 4 2
34 9 1 9 1 1 11 1 9 9 1 9 13 1 12 0 9 1 1 1 13 4 11 1 9 14 11 9 11 1 11 0 13 4 2
28 9 0 9 1 9 1 1 9 9 9 1 15 11 9 1 9 13 4 4 16 0 9 1 15 0 13 4 2
14 11 15 0 9 1 0 9 10 0 9 1 0 13 2
16 11 11 1 13 9 1 1 11 1 9 1 0 0 11 13 2
37 11 1 9 7 9 1 9 1 9 1 10 0 13 4 11 1 14 12 9 1 12 9 1 0 9 9 1 9 13 15 0 9 1 9 13 4 2
30 11 1 0 9 1 13 9 1 0 9 13 4 10 0 9 1 11 1 0 0 9 1 9 1 10 0 9 13 4 2
21 3 11 1 11 7 11 1 1 13 0 7 9 9 1 0 0 9 9 13 4 2
48 0 9 9 1 9 11 11 1 9 1 9 13 4 13 16 11 7 11 1 1 13 0 2 9 7 0 9 1 10 9 1 13 4 4 16 10 12 9 1 1 3 14 0 0 9 13 4 2
19 15 13 16 11 11 1 15 0 9 1 1 0 9 1 9 13 4 4 2
30 15 1 16 11 7 11 1 9 13 4 16 15 1 11 1 9 14 13 16 16 10 9 0 9 9 1 1 14 13 2
16 15 13 16 0 9 1 11 1 9 3 0 13 4 4 4 2
30 11 0 2 0 2 0 7 0 9 1 3 0 13 4 4 7 11 1 15 15 13 9 1 9 0 9 1 13 4 2
14 15 13 16 11 0 9 1 1 0 9 13 4 4 2
39 15 13 4 1 16 15 0 9 1 9 0 13 2 16 15 13 16 15 13 4 16 11 1 0 0 9 1 9 1 0 9 1 9 15 10 13 4 4 2
17 15 13 16 0 9 1 9 9 1 13 3 9 7 9 13 4 2
34 15 13 16 15 11 1 1 15 0 9 1 15 14 10 9 13 4 4 16 15 15 2 15 1 0 9 1 1 1 9 0 13 4 2
15 15 13 4 16 11 15 9 9 7 9 1 13 9 13 2
17 11 1 13 3 0 9 1 11 1 11 1 12 9 1 13 4 2
32 16 9 1 11 1 9 13 1 15 9 14 13 7 9 1 0 9 13 4 11 1 9 1 9 1 12 9 1 9 13 4 2
38 11 11 7 11 11 1 11 11 1 1 13 9 1 10 9 13 16 12 9 1 3 0 9 13 4 11 1 9 12 1 9 1 13 14 9 13 4 2
17 12 9 13 12 9 13 1 11 11 9 9 9 9 0 13 4 2
15 9 9 11 1 13 7 11 1 3 9 13 1 9 13 2
32 0 10 9 1 1 10 9 1 14 9 11 11 1 9 0 13 7 15 12 9 1 0 9 1 11 1 9 1 0 13 4 2
25 11 11 1 10 0 9 13 7 15 14 12 9 1 0 9 1 11 11 1 9 1 9 13 4 2
33 11 1 1 13 9 11 11 1 9 13 1 3 9 13 7 15 3 13 13 11 11 12 9 13 1 3 14 15 3 13 13 4 2
9 11 1 11 1 14 0 9 13 2
16 15 1 13 11 11 12 9 1 0 9 1 0 0 13 4 2
12 11 12 9 1 0 9 1 11 1 9 13 2
20 15 1 11 11 7 11 11 1 9 1 9 13 1 9 13 7 10 9 13 2
13 11 12 1 11 1 9 1 11 1 9 13 4 2
17 11 11 14 12 9 1 0 9 1 11 1 9 1 0 13 4 2
17 12 9 13 1 3 11 1 11 1 9 1 11 1 9 13 4 2
13 11 11 12 9 1 0 9 1 0 0 13 4 2
11 0 9 1 1 1 11 12 1 0 13 2
28 9 1 13 13 11 1 9 1 0 7 0 9 13 15 9 9 14 14 13 4 4 7 11 1 15 0 13 2
11 10 9 1 11 1 11 1 14 9 13 2
13 12 9 12 9 1 11 1 12 9 13 4 4 2
12 15 1 11 7 11 1 13 9 1 3 13 2
13 11 12 9 1 9 1 11 1 9 1 0 13 2
15 11 1 1 13 9 11 1 11 1 1 13 0 9 13 2
12 11 1 12 9 1 9 1 11 1 0 13 2
18 15 10 14 9 1 11 12 9 1 9 1 11 1 9 1 9 13 2
13 11 12 1 11 1 9 1 11 1 9 13 4 2
18 15 1 13 11 15 9 14 13 4 7 11 1 9 1 0 13 4 2
10 0 9 11 11 1 15 9 13 4 2
26 11 1 0 9 1 1 12 0 9 1 13 16 12 9 1 15 0 9 1 13 1 0 9 13 4 2
18 15 13 16 11 1 1 0 9 1 1 12 0 9 3 14 11 13 2
24 12 9 1 15 2 15 1 0 9 1 9 1 1 15 2 15 9 14 13 1 9 13 4 2
23 15 13 16 11 0 9 9 1 11 1 1 0 7 0 9 13 1 0 9 13 4 4 2
13 11 1 13 16 15 12 9 9 3 14 11 13 2
6 15 0 0 9 13 2
27 15 13 16 3 15 0 9 1 9 1 1 1 14 13 4 2 16 15 15 13 11 1 9 1 9 13 2
19 15 13 16 9 1 0 0 9 1 9 9 7 9 9 1 13 13 4 2
18 11 1 13 1 10 0 0 9 12 9 1 1 13 1 0 9 13 2
18 11 2 11 1 11 9 1 1 11 7 11 1 0 0 9 13 4 2
12 10 0 9 1 12 0 9 1 9 13 4 2
18 11 1 13 16 11 1 1 0 9 13 1 1 10 10 9 13 4 2
18 15 13 16 9 1 9 1 12 9 1 1 0 9 1 9 13 4 2
34 15 13 16 15 11 1 1 9 10 9 0 13 7 15 1 1 15 1 11 1 12 9 1 10 9 1 15 11 1 9 13 4 4 2
17 15 1 14 11 1 9 9 9 9 14 11 1 9 13 4 4 2
17 9 14 1 11 1 1 0 9 1 15 0 9 1 0 13 4 2
25 11 1 11 9 1 12 9 0 9 1 1 0 9 1 9 1 9 2 9 1 9 13 4 4 2
31 3 14 9 0 9 13 2 7 9 1 15 9 13 15 11 11 11 1 0 9 1 10 9 1 1 9 1 9 0 13 2
19 9 1 1 11 1 11 9 1 1 12 9 1 10 9 1 1 9 13 2
16 10 9 3 1 12 9 1 9 13 9 1 9 13 4 4 2
16 9 1 9 13 10 9 1 9 12 1 12 9 13 4 4 2
22 12 0 9 9 1 13 16 10 12 9 1 9 1 9 1 10 9 1 1 9 13 2
29 15 9 1 9 1 10 15 1 15 9 1 13 4 7 3 15 3 1 12 9 1 13 4 15 9 1 9 13 2
11 10 9 1 0 9 1 9 14 13 4 2
23 13 1 15 9 1 9 13 16 16 15 9 13 16 15 7 15 9 1 1 13 4 4 2
11 9 1 0 9 1 9 0 13 4 4 2
44 9 11 1 12 9 1 1 1 9 9 13 1 11 11 11 9 11 1 0 9 1 12 15 13 4 9 1 1 1 3 13 2 15 10 0 9 1 10 9 1 0 13 4 2
15 11 15 9 11 1 13 1 0 9 1 9 1 13 4 2
25 0 11 11 11 11 1 10 9 1 15 1 10 12 9 13 4 2 15 1 14 12 1 9 13 2
34 11 1 0 9 9 11 1 13 2 15 11 1 11 9 9 1 0 11 11 9 1 1 1 15 9 0 13 4 7 15 9 13 4 2
23 11 11 1 11 15 9 13 1 0 13 7 11 1 11 11 11 1 9 15 9 13 4 2
22 0 14 9 15 0 9 13 2 15 11 9 7 11 9 9 1 9 1 15 13 4 2
26 10 9 1 11 15 0 9 11 7 15 0 9 11 11 11 9 1 0 9 11 9 1 13 4 4 2
23 9 1 9 13 1 11 1 9 1 11 11 1 3 9 13 7 11 9 9 1 13 4 2
13 9 1 15 9 1 10 9 1 9 13 4 4 2
14 11 11 1 14 0 9 1 12 0 9 0 13 4 2
13 9 1 12 0 9 1 0 9 1 9 13 4 2
29 9 9 1 9 1 0 13 2 7 9 1 9 0 13 1 15 0 9 13 1 1 0 9 13 1 0 9 13 2
35 0 12 9 1 1 12 9 9 12 9 1 9 9 1 9 13 2 7 12 9 1 11 9 1 12 9 1 9 9 9 0 13 13 4 2
27 9 1 11 11 11 11 1 1 2 0 13 4 9 9 1 11 11 7 9 9 9 1 0 9 1 13 2
20 9 1 13 4 9 1 0 13 4 15 9 1 14 9 1 1 13 4 4 2
37 11 1 13 16 15 9 1 0 9 1 3 13 4 9 13 1 1 0 9 13 2 16 9 1 1 15 9 1 9 14 13 7 0 9 14 13 2
24 9 13 16 12 9 1 9 13 1 9 1 15 0 9 1 0 13 4 15 9 1 13 4 2
22 11 11 11 2 11 1 9 1 9 13 1 1 10 12 12 9 1 9 13 4 4 2
18 15 1 14 9 1 9 1 9 13 1 1 14 0 9 1 9 13 2
24 10 9 1 9 1 9 1 12 9 1 12 9 7 9 1 0 9 1 0 13 4 4 4 2
12 15 13 9 1 1 12 12 9 1 9 13 2
22 11 1 13 16 9 1 1 9 1 10 9 13 4 15 12 9 15 1 10 9 13 2
18 10 9 1 0 9 1 9 1 9 1 9 13 1 9 9 13 4 2
11 14 12 9 1 0 9 1 9 13 4 2
25 9 9 1 9 13 1 1 10 9 11 11 11 11 11 1 12 12 9 1 0 9 13 4 4 2
23 10 9 1 1 11 8 13 9 9 1 9 13 1 9 1 9 12 12 9 0 13 4 2
18 11 1 0 11 11 11 11 1 1 9 13 1 9 9 13 4 4 2
26 15 1 15 9 11 11 11 1 1 9 1 0 13 1 11 11 1 9 15 15 9 1 13 4 4 2
20 9 1 13 13 16 0 9 1 13 10 0 9 1 15 10 9 13 4 4 2
14 11 9 1 1 15 9 1 0 9 1 1 9 13 2
40 9 9 11 11 11 1 13 16 11 11 1 0 9 1 0 0 9 11 1 13 1 9 1 9 13 4 16 10 9 1 9 15 14 15 9 1 1 13 4 2
29 11 1 11 11 1 9 13 4 16 15 15 10 9 13 4 2 15 15 15 9 9 1 13 9 0 15 14 13 2
13 0 11 11 1 9 1 10 9 1 9 13 4 2
22 12 9 1 9 1 11 11 11 1 13 16 11 11 3 10 9 1 9 1 9 13 2
9 15 1 9 10 9 1 9 13 2
25 11 11 11 1 0 9 1 9 13 1 1 11 11 11 11 11 11 11 1 9 11 11 1 13 2
31 11 11 11 11 11 11 1 11 1 11 11 11 1 0 11 11 1 9 1 9 1 13 16 11 11 1 11 1 9 13 2
10 15 11 1 11 1 9 13 4 4 2
20 0 9 1 1 11 2 11 1 11 11 11 11 11 1 15 9 13 4 4 2
16 11 1 11 11 11 11 1 13 1 1 11 1 9 13 4 2
16 11 1 9 11 11 7 9 11 11 9 9 9 1 9 13 2
17 11 1 13 16 9 9 11 11 1 11 11 11 11 11 1 13 2
14 11 1 9 1 9 9 11 11 1 14 9 13 4 2
26 9 1 13 13 16 11 9 9 1 1 0 11 11 11 11 2 11 11 11 7 11 11 1 9 13 2
23 3 9 1 12 9 1 11 1 9 1 13 1 0 9 1 11 9 1 9 1 9 13 2
23 11 1 9 1 11 1 1 1 11 1 0 13 1 11 9 11 11 1 9 1 9 13 2
12 15 1 11 11 1 11 9 1 9 1 13 2
38 15 9 1 0 11 11 11 11 1 11 11 11 7 11 1 1 13 9 1 1 9 1 9 11 1 13 1 1 11 11 1 11 1 9 13 4 4 2
20 11 1 10 9 1 9 13 16 9 9 1 15 9 1 11 1 1 9 13 2
17 15 13 16 12 9 9 1 9 1 1 0 9 1 13 9 13 2
9 9 9 1 1 14 9 0 13 2
24 15 13 16 9 9 1 9 13 1 1 0 9 7 9 1 11 11 1 15 9 14 13 4 2
14 15 13 16 9 9 1 9 1 1 15 11 13 4 2
19 11 1 11 11 11 1 11 13 1 9 1 12 9 1 9 3 0 13 2
25 15 13 16 9 9 1 3 13 7 9 1 9 9 1 9 13 9 1 0 9 9 1 0 13 2
14 15 1 9 9 1 9 9 1 9 1 14 9 13 2
19 15 13 16 9 1 10 0 9 1 9 1 1 0 9 1 9 13 4 2
26 11 11 11 1 11 1 11 9 1 11 1 9 9 1 9 1 13 4 9 1 9 1 9 13 4 2
22 9 1 9 1 9 7 9 9 1 10 9 1 0 9 12 9 1 13 1 13 4 2
22 12 0 9 1 11 11 1 9 0 13 1 3 9 1 10 9 1 9 1 13 4 2
19 12 9 1 11 9 1 11 1 11 11 1 9 9 1 13 1 0 13 2
21 9 1 13 4 16 16 11 1 10 9 0 13 16 15 9 9 1 0 9 13 2
28 0 9 9 1 13 11 1 0 9 11 11 1 9 1 9 13 4 16 15 8 13 1 9 13 4 4 4 2
11 15 10 9 1 9 13 1 9 13 4 2
18 10 9 1 1 13 1 3 11 1 9 9 9 1 9 13 4 4 2
16 11 11 1 11 11 11 11 1 11 1 13 1 9 13 4 2
25 15 13 16 11 1 15 9 1 13 4 16 9 1 9 1 15 15 8 13 1 9 13 4 4 2
9 9 10 9 1 9 13 4 4 2
41 3 9 1 12 0 9 11 11 7 0 9 11 11 1 11 1 9 13 4 13 16 15 0 9 1 0 13 7 10 10 9 9 1 9 1 0 13 1 9 13 2
25 9 1 13 16 0 9 1 9 7 9 1 9 13 1 9 9 1 9 1 9 0 13 4 4 2
13 3 11 11 11 1 11 1 9 1 9 13 4 2
31 9 1 9 9 1 9 11 11 1 10 9 1 9 1 11 1 0 9 1 1 9 0 13 1 9 13 1 9 13 4 2
29 10 9 1 0 9 1 15 9 9 14 13 4 4 7 9 1 10 9 13 4 2 15 1 1 3 9 13 4 2
12 15 10 9 1 0 9 13 1 9 13 4 2
33 15 15 14 13 16 10 9 11 1 9 2 9 1 13 4 4 2 10 9 9 1 9 1 1 11 1 3 9 1 9 13 4 2
17 11 1 13 16 15 9 1 15 9 0 9 1 0 9 14 13 2
22 3 0 9 9 11 11 1 13 16 10 0 9 1 9 9 1 9 1 0 13 4 2
22 9 1 9 13 1 9 13 4 11 1 13 16 9 0 13 1 11 9 1 1 13 2
15 15 1 1 15 15 9 9 11 11 11 1 9 13 4 2
17 0 9 1 9 2 9 1 1 9 1 15 9 1 9 13 4 2
16 10 3 11 1 10 9 1 13 9 1 1 9 13 4 4 2
8 11 1 11 11 1 9 13 2
21 15 13 16 9 9 7 15 9 1 1 0 13 16 15 3 15 9 1 0 13 2
13 9 9 1 9 14 11 11 0 9 1 9 13 2
7 9 1 15 9 15 13 2
6 9 1 15 9 13 2
4 9 15 13 2
17 13 9 1 1 11 11 1 14 11 11 11 1 11 9 13 4 2
17 15 11 11 1 13 16 15 15 9 13 4 7 0 11 13 4 2
9 11 11 0 9 1 1 11 13 2
14 15 1 11 1 9 1 9 1 9 13 4 4 4 2
10 9 1 15 12 0 9 1 9 13 2
16 13 4 4 4 16 3 14 15 0 9 1 1 13 4 4 2
19 11 1 9 1 9 1 0 9 1 9 15 11 1 0 9 1 13 4 2
16 9 9 1 9 13 16 11 9 1 9 9 1 3 15 13 2
10 11 9 11 11 8 0 9 1 13 2
28 11 11 1 15 13 14 10 9 1 15 13 13 16 9 13 1 9 1 9 1 9 1 15 9 0 14 13 2
8 15 9 1 15 9 13 4 2
6 10 9 11 13 4 2
21 9 9 9 1 15 9 9 1 0 13 1 1 11 11 11 11 12 12 9 13 2
32 9 9 1 12 0 9 1 0 9 1 9 1 9 11 11 1 11 1 13 16 9 1 0 9 0 9 11 1 0 13 4 2
30 15 1 11 11 11 11 11 1 13 16 10 9 0 9 13 1 12 9 1 0 13 4 16 9 1 0 13 4 4 2
29 9 1 11 11 1 13 16 9 9 9 0 9 9 1 9 13 1 9 13 7 9 1 15 9 3 10 0 13 2
27 15 13 16 10 9 1 9 1 9 1 0 9 1 9 14 1 9 13 15 9 1 9 1 14 9 13 2
36 11 1 13 16 3 14 9 1 9 13 1 9 7 9 1 9 0 13 7 10 9 1 12 12 9 13 4 15 15 15 9 9 1 0 13 2
29 11 11 11 1 0 9 7 9 9 11 11 1 0 7 0 9 1 9 1 9 9 9 1 15 9 13 4 4 2
25 9 1 13 13 16 15 1 9 0 14 13 4 15 1 15 14 9 1 15 9 14 13 4 4 2
41 9 1 1 10 9 1 9 1 13 9 1 9 1 9 11 11 1 10 9 13 4 16 11 11 1 15 9 1 0 9 13 4 7 10 9 1 9 15 1 13 2
42 9 1 13 13 16 0 9 1 10 9 13 16 9 9 15 15 9 9 13 7 9 1 9 13 1 9 1 9 7 9 1 14 15 1 15 9 13 1 9 13 4 2
29 9 1 9 1 15 14 13 13 16 13 4 4 10 9 1 10 15 14 13 15 12 9 1 0 9 1 13 4 2
9 3 15 9 1 15 9 14 13 2
35 9 1 9 1 13 13 16 9 1 13 9 7 10 9 1 9 1 9 7 9 1 9 14 13 1 10 9 1 15 9 14 13 4 4 2
41 9 1 1 10 0 9 7 9 9 1 11 1 13 9 1 9 13 1 9 1 1 12 9 1 0 9 13 4 15 15 11 11 1 0 9 13 1 9 13 4 2
25 3 1 10 9 1 12 9 9 14 13 4 15 11 7 9 1 0 9 1 1 14 13 4 4 2
17 11 11 7 11 1 9 7 9 1 9 11 1 9 1 9 13 2
13 2 11 7 11 11 1 9 1 9 0 13 4 2
16 10 10 9 13 15 11 11 1 0 9 1 1 3 13 4 2
28 9 9 1 1 0 9 9 1 0 13 11 1 11 1 13 16 0 9 1 11 1 9 1 0 9 13 4 2
21 15 13 13 16 12 9 1 9 9 1 9 11 1 1 9 1 0 9 0 13 2
20 11 1 9 10 9 14 13 16 11 9 1 9 1 9 13 15 14 9 13 2
12 10 9 15 15 9 1 9 1 14 13 4 2
27 1 11 2 15 15 13 16 11 1 9 9 7 9 1 15 9 1 9 1 1 0 9 1 0 13 4 2
33 11 1 1 10 9 1 11 1 0 9 1 9 2 0 9 2 9 7 9 1 9 1 13 4 15 1 9 13 1 9 13 4 2
35 11 1 13 13 16 15 0 13 16 11 1 3 9 1 13 1 9 14 13 7 9 15 14 13 16 15 9 1 14 9 1 9 14 13 2
31 0 11 11 1 0 9 1 9 1 13 16 9 1 15 14 10 9 13 16 0 0 9 1 10 9 1 14 13 4 4 2
20 11 11 1 1 9 13 4 15 13 16 3 9 9 1 13 9 1 9 13 2
19 11 1 13 16 11 1 9 1 12 0 9 0 9 1 3 9 13 4 2
36 15 13 16 0 9 1 9 13 1 3 15 10 9 1 13 4 16 10 9 9 1 0 9 1 9 13 1 1 0 7 0 9 1 9 13 2
13 11 11 7 11 1 11 7 15 9 1 9 13 2
31 15 1 11 7 11 1 11 1 9 1 9 13 16 11 1 13 13 16 15 9 10 9 0 13 16 0 9 0 13 4 2
25 11 1 10 9 1 1 1 15 0 13 4 4 16 11 1 3 14 9 9 0 9 13 4 4 2
24 11 1 13 16 9 1 9 1 1 10 9 13 4 4 16 11 3 14 9 1 1 9 13 2
19 11 1 13 16 15 1 10 9 14 13 4 16 15 9 1 13 4 4 2
7 15 15 9 1 13 4 2
25 15 13 16 11 11 1 9 0 13 7 9 15 13 16 15 15 0 9 1 9 13 4 4 4 2
31 11 1 13 16 15 1 9 7 9 1 0 13 1 9 13 4 7 0 9 15 13 4 4 16 15 0 13 4 4 4 2
37 11 11 11 1 11 11 1 13 9 1 13 9 1 1 11 7 11 0 9 13 4 11 1 11 1 9 9 2 11 2 13 1 9 1 9 13 2
30 11 11 11 1 9 11 11 1 13 16 12 0 9 1 0 11 1 9 1 9 9 9 13 1 1 1 9 13 4 2
26 11 11 1 9 9 11 11 11 1 11 11 1 11 11 11 1 9 11 11 1 10 9 1 9 13 2
16 0 9 1 1 11 12 0 9 1 1 11 1 9 1 13 2
17 7 11 1 1 1 9 1 11 11 11 11 1 9 14 0 13 2
24 11 1 11 1 1 1 9 9 1 1 12 12 9 1 0 9 13 1 9 1 9 13 4 2
32 0 13 16 11 1 11 1 9 9 1 9 1 1 0 11 11 11 1 11 1 12 12 9 1 0 9 13 1 9 13 4 2
32 11 1 9 9 1 12 9 11 1 11 11 2 11 1 11 7 11 1 11 2 11 2 11 1 9 9 13 1 9 13 4 2
20 10 9 1 11 11 11 1 9 9 13 15 9 13 4 7 9 9 13 4 2
24 12 0 9 1 11 1 11 11 11 11 11 11 11 1 1 0 9 1 9 1 0 13 4 2
18 9 11 11 1 11 1 9 9 1 9 11 11 1 0 13 4 4 2
22 11 11 1 11 11 1 15 9 1 13 4 16 9 11 1 9 1 11 1 9 13 2
9 9 9 11 11 1 0 13 4 2
18 15 15 9 1 13 16 11 1 1 0 9 1 15 9 14 13 4 2
33 11 1 9 13 1 12 9 1 11 11 1 11 11 11 11 2 11 2 1 9 1 9 1 1 11 11 1 0 9 1 9 13 2
15 11 11 11 0 9 15 10 9 1 9 1 15 9 13 2
21 10 3 11 1 0 2 0 7 0 9 1 13 4 9 1 9 1 9 13 4 2
20 3 1 0 9 2 9 7 9 1 13 1 0 9 1 9 2 9 13 4 2
25 11 11 1 0 9 1 13 9 13 1 9 0 9 11 11 11 11 1 10 9 1 0 9 13 2
23 0 9 1 10 9 1 11 11 11 2 11 2 1 1 13 4 9 1 15 0 13 4 2
27 16 2 9 1 1 10 9 9 2 9 9 1 9 7 9 9 1 9 1 13 9 1 15 9 0 13 2
20 0 11 9 11 11 1 1 0 9 1 11 11 11 1 9 0 9 13 4 2
21 9 3 9 1 9 2 9 7 9 9 1 9 9 13 1 1 9 13 4 4 2
11 9 1 10 10 9 1 9 13 4 4 2
13 11 1 0 9 9 1 9 13 1 9 13 4 2
26 9 9 1 9 1 9 13 4 15 13 16 0 9 1 9 9 1 15 9 1 9 1 9 14 13 2
9 9 1 1 15 10 9 1 13 2
23 9 9 1 9 13 4 15 13 16 10 9 1 9 1 1 3 10 9 13 4 4 4 2
25 9 9 1 9 13 1 9 1 9 13 4 11 9 1 13 16 10 9 1 9 9 13 4 4 2
9 15 15 9 1 15 9 14 13 2
19 11 1 11 11 1 13 16 9 1 0 9 1 1 15 14 13 4 4 2
20 0 9 1 1 0 9 14 13 7 9 1 9 1 0 9 0 9 1 13 2
15 9 1 9 1 1 15 10 9 1 0 9 1 1 13 2
15 11 9 11 11 14 9 9 13 4 1 9 1 0 13 2
12 15 9 13 16 15 0 9 1 0 9 13 2
9 9 1 1 15 0 9 14 13 2
14 9 1 1 9 9 1 3 10 9 13 4 4 4 2
23 11 11 1 9 9 1 13 9 1 9 9 9 1 14 13 15 1 9 0 13 4 4 2
35 11 11 11 11 7 11 11 11 11 11 11 1 9 1 9 9 11 11 7 11 11 1 9 1 9 9 9 9 1 9 1 1 9 13 2
20 9 1 9 1 9 9 1 11 13 13 1 1 0 9 13 1 9 13 4 2
27 15 1 10 9 1 14 11 13 1 9 13 4 15 10 9 1 1 11 7 11 1 1 11 13 13 4 2
26 11 11 1 9 1 1 9 1 9 10 9 13 4 16 11 1 9 1 11 14 13 1 9 13 4 2
10 10 9 1 9 3 0 13 4 4 2
23 11 11 1 14 10 9 1 9 1 11 1 0 9 1 9 13 1 14 9 13 4 4 2
24 7 9 9 9 1 9 13 16 11 11 1 14 9 0 9 1 14 13 1 14 9 13 4 2
38 16 2 11 11 1 13 1 9 1 9 1 9 1 13 1 1 0 9 1 1 9 1 15 13 1 9 13 16 9 9 1 0 9 0 14 13 4 2
26 0 9 9 1 9 1 9 9 13 13 4 4 7 11 11 1 9 1 9 1 14 9 13 4 4 2
23 7 0 9 13 1 1 9 9 1 11 11 1 9 1 9 1 13 4 9 1 0 13 2
15 9 9 1 9 13 1 14 9 9 1 15 9 14 13 2
15 10 9 11 11 11 11 11 11 1 0 9 1 13 4 2
33 0 9 1 13 4 9 1 13 4 4 16 11 11 11 1 12 13 12 9 1 11 11 11 1 0 9 1 12 9 1 9 13 2
21 12 1 12 9 1 2 9 9 1 0 9 8 13 4 2 15 14 10 9 13 4
22 10 3 9 1 0 9 1 9 7 0 9 1 9 1 1 1 9 0 13 4 4 2
26 3 14 9 9 1 15 0 12 9 11 11 1 9 1 9 1 13 4 9 1 0 13 1 13 4 2
39 9 1 13 4 4 16 2 11 11 1 9 12 1 12 9 1 1 0 9 1 10 9 1 9 1 9 13 16 15 9 1 9 1 9 0 13 4 4 2
23 9 1 9 10 13 1 1 15 13 0 13 4 16 15 9 1 9 13 1 9 14 13 2
22 7 9 1 9 1 3 10 9 2 9 1 13 1 9 2 1 0 13 1 9 13 4
11 9 9 1 9 1 9 1 13 4 4 2
11 9 11 13 1 1 9 9 1 13 4 2
9 9 9 1 13 1 9 13 4 2
13 10 3 0 9 1 9 1 9 13 4 4 4 2
14 0 12 9 1 10 15 13 15 1 9 13 0 13 2
10 9 9 1 9 1 0 9 0 13 2
26 9 1 1 2 9 9 1 10 9 1 9 13 4 16 0 9 1 1 13 9 1 9 3 10 13 2
14 15 9 1 9 13 1 1 3 10 9 1 8 13 4
14 9 9 9 8 13 4 7 9 9 9 1 13 4 2
12 3 9 9 1 9 9 1 9 15 14 13 2
23 9 1 1 2 16 11 11 1 11 9 1 9 9 0 9 2 9 1 12 9 1 13 2
12 10 9 1 9 9 1 3 10 9 14 13 4
21 9 1 1 1 10 9 1 9 13 4 4 16 11 11 1 15 9 13 13 4 2
21 7 11 1 10 9 1 10 10 9 1 1 13 4 4 15 9 14 13 4 4 2
41 9 1 9 1 1 11 11 11 11 1 13 16 0 11 11 11 9 1 9 9 1 10 9 1 0 13 16 9 9 1 9 1 1 3 9 13 4 1 9 13 2
43 10 9 1 11 9 1 9 11 11 1 13 4 9 1 9 1 11 11 1 13 16 9 9 1 0 9 13 1 1 12 9 1 9 9 1 9 0 9 13 1 9 13 2
20 11 11 1 13 16 11 11 1 9 9 1 9 9 1 9 1 13 4 4 2
23 15 13 16 12 9 1 9 9 1 11 7 11 1 9 13 0 9 13 1 13 4 4 2
28 11 11 1 13 16 10 9 9 1 0 9 1 0 9 1 9 11 1 11 2 11 1 1 15 9 14 13 2
23 9 9 1 9 1 1 1 11 1 13 16 11 1 11 1 1 10 9 1 13 4 4 2
40 11 1 9 1 13 0 0 9 1 11 1 13 4 16 15 1 9 11 1 9 1 9 13 4 7 0 9 1 13 4 1 9 1 1 15 13 4 0 13 2
56 15 1 1 9 1 12 9 1 9 1 11 11 11 11 1 13 16 11 9 11 1 11 11 11 7 15 9 1 9 13 4 2 0 9 1 13 4 7 0 9 3 9 13 4 1 9 13 1 3 10 9 13 0 0 13 2
17 11 11 1 13 16 9 11 1 1 9 1 3 9 13 4 4 2
25 15 13 16 9 9 1 15 9 1 9 1 9 7 0 9 1 1 9 13 1 14 9 13 4 2
15 11 11 1 11 11 1 13 4 9 1 9 13 4 4 2
34 11 1 13 16 0 11 11 1 9 7 0 0 9 1 9 9 1 1 15 13 4 9 1 13 4 11 1 11 1 9 14 13 4 2
9 15 1 12 1 12 9 0 13 2
37 11 11 1 0 0 9 1 9 1 13 4 9 9 1 10 0 14 9 1 9 2 9 9 9 0 13 9 1 12 0 0 9 13 1 9 13 2
34 15 1 9 1 11 11 1 9 1 12 9 2 9 9 0 13 4 4 2 7 11 1 13 9 1 10 9 1 3 9 13 4 4 2
30 16 9 1 9 1 13 0 9 9 9 11 11 1 13 13 16 15 0 12 9 1 9 1 0 9 13 9 13 4 2
32 0 9 1 1 1 9 1 13 9 1 0 9 1 9 13 1 3 15 13 16 12 9 1 15 9 1 0 9 0 13 4 2
15 15 13 16 9 9 7 9 1 15 9 9 13 1 13 2
10 15 9 13 1 1 9 14 0 13 2
31 0 13 16 11 11 11 1 1 11 1 1 2 9 11 1 9 11 11 1 0 9 1 1 11 2 11 1 9 13 4 2
24 7 11 11 11 11 7 11 11 11 11 1 9 9 7 9 9 1 9 1 1 13 4 4 2
9 15 1 12 1 12 9 0 13 2
35 11 9 11 11 7 9 9 11 11 1 1 11 11 1 12 9 1 9 13 1 3 11 1 13 16 12 9 1 13 4 1 9 13 4 2
10 11 1 9 13 12 9 9 13 4 2
20 3 2 11 1 11 9 3 10 0 13 2 15 0 9 9 12 1 13 4 2
20 11 1 12 9 1 0 9 1 1 11 1 9 10 9 1 3 0 9 13 2
25 0 9 1 13 16 11 11 11 1 11 1 11 0 11 11 1 9 1 12 9 0 9 13 4 2
21 0 11 9 1 9 2 9 9 1 12 9 1 1 12 9 0 9 1 13 4 2
14 11 1 9 13 9 1 9 13 12 9 9 13 4 2
11 9 1 10 9 0 9 1 14 13 4 2
9 15 9 13 12 9 13 4 4 2
10 15 1 11 11 1 9 12 9 13 2
7 15 9 9 9 12 13 2
15 7 0 9 11 1 11 1 10 9 1 3 10 9 13 2
13 15 0 9 12 9 9 13 15 11 1 12 13 2
13 15 1 1 0 9 1 9 1 0 9 13 4 2
16 9 9 1 9 1 1 10 9 1 9 1 10 9 13 4 2
22 11 9 1 9 0 9 13 4 15 1 12 12 9 1 9 1 14 13 0 13 4 2
11 15 1 9 1 9 1 9 1 9 13 2
19 7 0 9 9 1 9 1 1 9 1 13 7 9 13 14 1 9 13 2
16 9 12 9 11 9 1 12 9 1 14 14 13 4 4 4 2
11 15 9 9 1 14 9 9 1 1 13 2
11 9 1 9 9 9 1 1 13 9 13 2
13 15 1 9 9 1 9 12 9 0 13 4 4 2
44 15 11 1 11 11 11 2 11 2 11 11 11 2 11 2 11 11 2 11 2 11 11 11 2 11 2 11 11 11 2 11 2 11 11 11 7 11 11 2 11 11 0 13 2
20 15 9 12 12 9 13 7 15 15 1 1 3 0 0 9 13 4 4 4 2
19 0 9 9 11 1 11 9 1 10 0 9 1 9 9 1 10 9 13 2
14 0 9 1 9 1 9 1 10 0 9 13 4 4 2
21 15 15 9 7 9 1 1 1 9 13 4 16 15 11 1 10 9 13 4 4 2
31 11 1 11 11 1 9 11 11 1 1 10 0 3 10 9 9 1 11 11 2 11 9 1 9 1 9 13 13 4 4 2
10 10 9 9 1 14 12 9 3 13 2
11 9 15 2 11 11 2 14 13 4 4 2
16 9 12 10 9 1 9 13 4 4 15 15 9 1 1 13 2
14 7 9 1 13 4 4 16 15 12 9 0 13 4 2
14 9 7 15 10 0 9 14 12 12 12 9 0 13 2
8 15 9 1 9 1 9 13 2
15 13 4 4 4 16 10 9 10 9 1 13 1 13 4 2
31 11 9 1 11 1 13 16 10 2 11 11 2 12 12 9 0 13 7 15 1 15 1 13 4 9 1 15 3 0 13 2
17 11 1 11 11 1 9 11 11 1 10 0 9 1 12 9 13 2
21 11 11 2 11 1 1 13 4 9 1 13 1 14 12 12 9 1 9 13 4 2
11 15 0 9 7 9 1 9 1 13 4 2
15 0 9 1 13 4 4 4 16 9 3 0 13 4 4 2
21 11 1 13 16 16 15 9 13 16 15 0 9 1 9 1 2 0 9 2 13 2
15 15 0 9 1 10 0 9 1 0 10 9 13 4 4 2
18 3 11 1 11 11 9 1 12 9 14 1 13 9 1 9 13 4 2
13 15 9 1 12 9 9 1 11 9 1 0 13 2
22 0 13 16 11 1 11 9 9 1 11 9 1 13 1 9 9 1 9 13 4 4 2
29 15 1 14 11 9 1 10 9 1 9 1 9 14 13 4 4 15 9 2 11 7 9 9 1 9 1 13 4 2
9 10 9 1 0 13 4 4 4 2
19 9 1 13 13 16 15 9 1 9 9 1 1 1 0 9 13 4 4 2
16 13 4 4 16 9 1 9 1 9 1 9 9 1 9 13 2
23 9 1 10 9 1 9 1 14 13 4 4 7 9 1 9 1 15 13 4 0 9 13 2
21 9 1 11 2 11 1 0 9 0 13 9 2 9 13 1 9 9 1 13 4 2
26 10 10 9 9 9 1 13 4 15 9 1 11 2 11 1 0 9 1 9 0 13 9 2 9 13 2
20 0 9 1 13 16 10 9 1 11 1 11 11 13 4 11 1 9 13 4 2
15 11 13 15 9 1 9 1 0 9 13 1 9 0 13 2
9 15 1 15 9 2 9 14 13 2
12 10 10 9 11 9 1 11 9 1 13 4 2
20 12 0 9 1 13 16 11 1 9 1 13 1 3 0 9 13 4 4 4 2
12 11 9 9 1 1 0 0 9 1 9 13 2
12 10 9 1 13 9 11 1 9 13 4 4 2
27 11 11 0 12 9 1 9 1 10 9 1 0 9 1 1 1 13 1 9 1 0 11 11 1 0 13 2
15 15 1 11 2 11 1 9 9 1 9 1 0 9 13 2
7 11 11 1 9 0 13 2
20 0 13 16 0 9 12 0 0 9 1 0 9 13 1 9 9 1 13 4 2
27 11 11 0 0 9 1 9 11 1 0 9 13 1 9 0 13 11 1 11 9 1 9 2 9 13 4 2
16 15 1 0 9 13 0 9 1 15 9 13 1 14 9 13 2
13 11 11 1 9 1 9 1 0 9 1 9 13 2
40 11 1 9 2 9 9 7 11 1 9 1 13 4 9 1 9 1 11 1 11 11 11 11 11 1 11 7 15 9 1 0 9 1 9 0 13 1 9 13 2
11 3 11 1 9 15 1 0 9 13 4 2
15 9 13 4 16 9 1 0 0 9 1 9 3 10 13 2
32 11 1 11 11 11 1 1 9 1 9 13 1 11 11 1 1 0 9 13 4 11 1 15 11 1 11 11 11 0 13 4 2
14 9 1 9 1 9 9 1 15 9 1 9 13 4 2
23 11 11 11 1 9 11 11 1 13 16 3 11 1 11 11 1 15 9 1 14 13 4 2
23 11 11 1 13 1 0 9 13 4 4 7 15 1 1 0 11 11 11 11 1 13 4 2
24 9 9 1 9 9 13 1 9 1 10 9 1 3 13 7 15 1 9 13 1 9 13 4 2
14 11 1 13 16 9 15 14 9 1 10 9 14 13 2
22 3 9 1 9 11 11 1 13 4 16 9 1 9 1 13 4 11 1 13 0 13 2
14 11 11 1 13 1 9 14 11 1 14 13 4 4 2
33 11 1 12 0 9 1 13 13 16 11 1 9 1 9 9 1 9 1 1 9 1 0 9 13 7 15 9 9 1 3 9 13 2
27 11 1 13 0 0 9 11 11 0 9 1 9 9 1 13 4 4 16 15 9 1 3 0 9 11 13 2
53 0 13 16 11 1 11 11 1 0 9 11 11 11 1 9 1 9 1 0 9 11 11 0 9 1 1 12 9 1 9 9 13 4 4 7 15 1 0 13 16 9 1 12 9 1 9 9 1 9 14 12 13 2
7 15 3 0 11 11 13 2
12 7 9 9 11 11 1 15 0 9 13 4 2
19 16 11 1 1 11 1 13 16 0 9 1 9 0 13 15 9 13 4 2
18 7 9 1 9 1 1 9 13 1 1 15 11 11 11 0 13 4 2
22 11 1 9 9 11 11 11 1 13 16 11 1 9 1 11 1 9 13 1 13 4 2
26 11 9 1 11 7 15 9 9 1 9 13 16 16 15 9 13 16 10 9 9 9 1 1 9 13 2
11 10 9 9 1 0 11 1 9 13 4 2
36 0 9 15 13 16 10 9 1 14 10 14 9 0 13 11 1 0 11 11 11 1 9 13 4 4 4 7 15 11 11 1 0 9 13 4 2
16 10 9 10 14 9 11 7 15 9 11 1 1 13 4 4 2
11 0 9 11 1 3 15 9 13 4 4 2
13 15 1 11 0 9 1 11 11 1 9 13 4 2
27 11 1 0 13 16 11 1 9 1 13 1 9 13 4 4 7 15 9 13 16 9 1 9 13 4 4 2
16 0 9 13 14 9 9 1 9 1 9 14 0 13 4 4 2
21 0 7 0 9 1 9 9 1 13 4 9 10 9 9 1 9 1 13 4 4 2
25 11 1 0 9 9 11 11 11 0 13 4 2 9 9 1 9 13 1 3 9 1 9 13 4 2
6 9 1 9 3 13 2
14 9 9 1 9 1 1 11 11 11 11 3 0 13 2
16 10 9 1 9 13 4 9 1 9 1 12 9 9 0 13 2
37 16 15 10 9 12 12 9 13 7 15 12 12 9 11 11 11 11 1 9 13 4 16 0 0 9 1 1 15 10 9 12 12 12 12 13 4 2
25 7 9 13 2 15 15 10 9 1 12 9 1 10 1 9 9 1 9 9 1 9 14 13 4 2
24 0 13 16 15 14 9 1 9 13 9 1 9 1 12 9 9 9 1 9 14 13 4 4 2
18 11 11 11 1 1 12 9 1 13 12 11 1 1 9 1 9 13 2
48 9 9 11 11 13 4 2 9 9 1 11 11 11 1 1 14 10 9 1 9 13 9 1 9 1 12 9 9 9 0 13 4 2 15 11 11 11 1 1 9 9 13 1 9 13 4 4 2
20 15 9 13 1 3 9 1 13 4 9 7 10 9 1 9 1 9 13 4 2
12 9 1 9 1 9 13 1 1 15 0 13 2
19 9 1 10 14 10 9 1 13 1 1 11 1 8 13 11 11 11 11 2
30 15 1 9 13 1 9 1 11 11 11 11 1 1 14 9 13 7 9 9 1 9 1 12 9 1 1 9 13 4 2
20 9 1 12 12 1 10 0 9 13 14 11 11 1 1 9 9 0 13 4 2
15 9 0 9 9 1 9 1 9 1 13 8 13 4 4 2
17 10 9 1 9 0 12 12 9 9 13 1 9 14 13 4 4 2
17 0 9 1 10 0 13 1 12 12 1 9 1 0 9 13 4 2
12 0 3 0 9 13 1 9 1 9 14 13 2
13 9 15 1 12 12 9 9 1 1 1 13 4 2
19 9 1 9 13 7 9 9 9 9 1 9 1 15 12 9 9 13 4 2
25 11 11 11 11 11 2 11 1 0 9 1 9 11 1 9 9 1 11 11 11 1 9 1 13 2
24 15 11 11 11 1 1 1 9 13 1 9 1 9 13 4 13 4 16 15 12 0 9 13 2
11 15 9 1 9 13 7 9 1 9 13 2
14 9 1 9 1 13 9 1 11 1 9 0 13 4 2
21 15 10 9 9 7 9 1 9 9 1 1 1 13 4 9 1 13 1 9 13 2
40 9 1 9 13 4 16 10 9 1 9 13 4 4 7 11 1 9 1 0 13 1 13 4 2 16 9 9 1 10 9 1 13 4 4 2 15 1 13 4 2
67 10 9 1 9 1 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 11 2 11 11 11 2 11 11 2 11 11 11 2 11 11 11 2 9 11 11 11 2 11 11 11 7 11 11 14 1 9 13 7 11 1 9 1 9 13 2
26 11 11 11 11 11 11 1 11 11 2 11 2 1 9 1 9 9 11 9 13 1 9 13 4 4 2
20 11 1 11 1 15 11 9 1 1 11 1 9 9 9 13 1 9 13 4 2
21 11 11 1 15 0 9 1 9 13 4 11 1 15 9 13 12 9 1 14 13 2
28 11 1 9 11 11 11 1 13 16 9 9 1 9 1 0 13 4 16 11 15 9 1 9 9 9 14 13 2
13 11 1 15 1 10 9 1 9 9 1 13 4 2
24 11 9 1 1 9 1 9 11 1 9 1 0 9 9 9 11 11 1 11 1 0 13 4 2
25 9 1 9 11 1 0 11 11 11 11 7 11 1 9 11 11 11 1 9 11 1 0 13 4 2
12 11 11 1 15 0 9 9 1 14 9 13 2
27 11 1 9 11 11 1 13 16 9 9 1 0 9 1 1 11 1 11 1 9 1 9 13 4 4 4 2
25 15 0 9 1 9 1 13 0 11 1 13 16 15 11 1 9 13 16 15 9 1 1 9 13 2
34 15 13 16 11 1 9 1 1 14 15 9 11 1 9 0 13 4 2 15 9 11 1 0 11 11 11 11 1 9 1 0 13 4 2
29 11 11 11 11 11 1 12 9 9 1 13 4 4 4 9 11 1 9 11 2 11 1 1 9 1 9 13 4 2
17 9 9 11 11 1 11 1 11 9 1 9 1 9 0 13 4 2
21 9 1 15 13 4 16 11 2 11 11 1 11 1 11 1 9 1 9 9 13 2
17 9 9 9 1 1 9 13 9 1 9 7 0 9 1 9 13 2
28 11 1 13 16 11 1 11 9 1 1 15 11 1 9 1 0 9 1 1 9 1 11 1 11 13 4 4 2
11 15 13 16 15 9 1 9 1 9 13 2
10 9 1 9 9 1 11 13 4 4 2
10 9 1 9 1 1 9 9 0 13 2
23 11 11 1 9 1 11 1 9 1 0 2 0 13 1 1 9 9 1 9 1 9 13 2
37 11 1 9 1 9 1 0 9 1 13 12 9 1 9 7 9 1 0 13 1 9 1 14 12 9 11 2 11 11 1 0 13 9 13 4 4 2
23 9 1 13 13 16 9 1 15 1 12 9 1 11 1 1 9 1 9 1 0 13 4 2
16 9 1 0 2 0 13 1 1 9 1 9 9 1 9 13 2
7 15 12 9 0 13 4 2
10 15 9 11 11 1 1 1 13 4 2
9 15 9 1 1 9 13 4 4 2
42 0 13 16 11 1 11 1 9 9 1 1 0 9 1 13 1 9 13 1 1 13 1 9 1 1 9 11 1 9 1 0 9 1 9 11 11 1 9 13 4 4 2
10 7 15 9 11 11 0 13 4 4 2
7 15 1 15 9 13 4 2
16 11 11 0 0 9 1 11 11 11 1 0 13 1 9 13 2
23 11 1 0 13 1 11 1 9 1 11 11 11 11 1 13 16 9 9 9 1 9 13 2
12 15 0 9 1 13 1 0 9 9 1 13 2
17 11 1 13 16 15 9 15 14 13 16 11 1 15 9 14 13 2
12 11 10 9 1 9 1 0 9 13 4 4 2
28 9 1 9 1 11 1 13 16 11 1 13 13 16 9 9 1 14 9 1 1 1 14 0 14 13 4 4 2
11 15 1 0 9 1 9 13 14 0 13 2
17 9 1 10 9 1 9 1 1 12 2 12 12 9 13 4 4 2
16 0 9 1 9 1 1 11 11 11 1 9 1 0 13 4 2
17 11 1 13 16 0 0 9 1 9 9 1 12 9 13 4 4 2
14 9 1 9 1 9 1 1 14 12 9 13 4 4 2
31 9 9 1 13 10 9 3 11 1 9 9 13 13 4 7 9 1 9 1 9 1 9 13 15 9 13 1 9 13 4 2
16 3 1 9 1 13 16 10 9 1 9 1 0 9 13 4 2
28 11 1 9 13 16 10 9 11 1 11 2 11 1 0 9 1 9 13 4 2 7 11 1 10 9 13 4 2
10 10 9 11 1 10 12 0 9 13 2
13 15 12 0 9 7 9 9 1 12 9 13 4 2
19 7 0 9 15 1 12 0 9 1 12 0 9 7 12 9 9 13 4 2
30 0 9 1 0 9 1 9 1 9 1 1 11 1 11 1 11 1 2 12 0 9 7 9 2 0 13 1 13 4 2
32 9 9 7 0 9 1 0 0 9 1 9 1 1 11 1 9 13 4 1 3 11 10 9 1 9 13 1 0 13 4 4 2
28 12 9 15 2 15 1 15 13 4 9 1 15 9 1 9 1 9 1 13 1 9 13 1 0 13 4 4 2
14 12 9 1 1 12 0 0 0 9 11 1 0 13 2
33 10 9 1 12 9 1 0 0 9 7 0 9 1 9 1 9 1 13 1 9 13 1 0 13 4 12 0 9 2 9 0 13 2
42 9 1 11 1 11 11 11 11 1 1 9 13 1 0 11 11 11 11 11 1 13 16 12 9 1 15 0 9 1 0 13 4 9 1 9 1 0 9 1 9 13 2
31 12 9 1 1 9 1 9 13 4 11 1 13 16 11 1 0 11 11 1 1 11 1 11 11 11 1 9 1 9 13 2
18 11 1 0 9 13 7 15 14 9 1 9 1 9 1 9 14 13 2
34 9 1 1 11 1 0 13 16 15 15 11 1 13 9 1 11 1 0 11 1 9 1 9 9 1 15 9 1 9 1 0 14 13 2
7 9 1 9 13 4 4 2
20 9 1 13 4 4 16 12 9 9 7 9 1 9 13 1 0 13 4 4 2
33 9 1 9 1 9 1 11 1 11 11 1 10 9 1 0 9 0 13 1 13 2 15 9 1 12 9 1 1 9 13 4 4 2
18 12 9 1 0 9 1 9 13 1 1 3 9 1 9 1 9 13 2
20 0 9 1 13 1 1 14 12 9 9 1 9 13 7 9 13 1 0 13 2
28 11 11 1 9 1 9 13 4 11 1 13 16 11 11 1 11 11 11 11 1 15 9 9 1 9 13 4 2
13 7 11 1 11 1 0 13 1 9 14 13 4 2
40 15 1 1 11 11 11 1 1 1 0 9 1 13 4 4 16 11 1 9 1 9 1 1 11 1 15 9 1 9 9 1 0 13 4 7 15 9 13 4 2
17 7 9 1 11 1 9 15 9 9 1 1 14 13 4 4 4 2
35 11 1 10 9 13 4 13 16 11 11 1 11 1 10 10 9 13 4 15 13 1 13 4 16 15 15 9 9 1 1 13 9 13 4 2
31 11 1 13 16 0 9 1 3 1 15 13 13 4 16 11 1 9 1 13 4 9 1 9 7 9 1 9 14 13 4 2
15 11 1 13 16 0 9 1 0 9 1 9 13 4 4 2
23 10 9 1 9 1 11 11 1 11 1 13 11 11 1 11 1 13 4 1 9 13 4 2
22 15 9 13 15 9 1 15 0 9 13 7 9 1 0 13 4 1 15 13 13 4 2
23 9 1 9 1 9 1 15 15 9 9 14 13 4 7 3 0 9 1 9 9 13 4 2
41 15 1 13 9 1 9 13 11 1 11 11 9 1 13 1 11 2 13 4 9 2 15 0 9 1 13 9 1 1 3 2 3 13 4 7 15 12 14 13 4 2
26 13 15 11 11 11 1 9 1 9 13 7 15 9 1 9 1 1 3 12 0 9 13 4 4 4 2
16 11 0 9 1 11 1 11 11 9 1 11 1 13 4 4 2
25 7 0 9 1 15 9 1 0 13 1 9 1 15 9 11 11 11 1 11 9 1 13 4 4 2
14 15 15 9 1 9 12 9 2 9 9 1 13 4 2
12 11 11 1 0 9 1 13 15 9 13 4 2
14 10 3 11 11 15 9 1 1 0 11 13 13 4 2
12 11 15 14 3 11 1 13 1 1 13 4 2
7 10 3 11 0 13 4 2
14 15 9 3 14 11 1 13 15 11 13 0 13 4 2
33 15 11 11 1 15 9 1 9 1 9 13 15 15 0 9 1 9 1 11 1 9 13 3 15 9 11 1 11 11 1 13 4 2
23 11 11 1 15 9 14 13 4 7 15 9 1 10 9 1 9 1 13 1 9 13 4 2
6 9 0 11 13 4 2
10 10 3 11 1 12 9 1 9 13 2
18 9 1 9 13 14 11 15 9 1 9 13 12 9 3 13 4 4 2
36 9 1 3 0 13 1 0 11 15 13 7 9 13 1 1 9 1 1 13 7 15 9 13 1 1 15 9 1 0 13 1 9 13 4 4 2
9 13 15 11 11 11 1 9 13 2
19 9 1 11 11 1 11 1 10 9 1 9 13 7 3 9 13 1 13 2
16 9 1 9 1 1 0 9 0 13 7 11 1 13 13 4 2
31 11 1 15 9 7 9 1 10 9 1 9 13 4 16 15 9 1 13 7 14 13 15 15 9 7 15 9 1 3 13 2
24 12 9 1 9 1 9 13 4 13 4 11 11 1 9 1 15 13 9 13 1 9 13 4 2
12 11 1 12 0 9 11 13 7 15 9 13 2
16 12 9 1 11 11 11 11 1 0 9 11 11 1 9 13 2
19 11 11 11 11 9 1 9 9 13 7 9 11 1 15 9 13 4 4 2
12 15 1 11 11 9 1 1 9 13 4 4 2
16 0 10 9 1 11 1 13 1 15 9 15 9 13 4 4 2
19 9 1 13 1 1 11 11 1 9 1 1 13 10 9 1 13 4 4 2
20 15 9 13 16 15 9 3 13 7 0 9 1 13 1 3 15 10 0 13 2
18 15 13 16 10 0 9 15 13 13 4 7 15 15 0 9 0 13 2
16 15 9 13 16 15 12 9 1 0 15 9 15 3 13 4 2
19 9 11 11 1 13 16 12 0 9 11 11 1 13 1 1 9 13 4 2
14 11 1 13 16 9 1 15 9 13 1 9 13 4 2
24 15 13 16 15 11 11 1 1 1 9 13 4 4 7 9 9 1 15 15 9 11 13 4 2
15 9 1 13 16 9 1 9 9 1 15 14 13 4 4 2
15 0 13 16 11 11 12 9 1 9 1 15 9 9 13 2
22 11 1 13 16 11 11 9 1 1 11 9 11 11 7 11 11 1 14 13 4 4 2
18 15 13 16 11 11 1 10 9 3 1 1 1 9 1 10 9 13 2
9 15 9 13 7 9 14 14 13 2
17 15 0 9 1 9 11 1 9 13 4 2 15 15 9 13 4 2
19 9 1 9 13 7 9 1 1 1 10 9 15 9 3 0 13 4 4 2
36 11 1 13 16 9 1 9 9 1 15 9 7 15 0 9 1 1 1 9 13 1 3 1 10 9 1 9 15 13 1 1 9 13 4 4 2
25 10 0 0 9 14 15 13 1 1 13 7 0 9 1 9 13 2 7 11 11 1 9 13 4 2
55 11 11 1 0 9 9 9 11 11 11 2 0 9 11 11 2 9 9 9 11 11 2 9 11 11 2 9 9 11 2 9 9 11 11 11 2 9 9 11 11 7 11 1 11 11 1 12 9 1 9 9 1 13 4 2
23 11 11 9 1 0 11 11 1 12 9 10 9 1 9 9 13 1 1 0 14 13 4 2
39 11 11 1 11 11 1 11 1 0 0 9 1 11 11 11 11 11 11 1 9 9 9 1 0 9 1 15 2 15 9 1 12 9 1 9 9 9 13 2
15 10 9 9 9 1 1 10 12 9 1 9 13 4 4 2
20 9 9 1 0 9 1 11 11 1 11 1 12 9 1 9 9 1 0 13 2
49 9 9 1 0 9 1 11 1 12 9 1 9 9 13 4 4 7 11 1 0 9 11 11 2 11 11 2 2 9 11 11 11 11 7 9 11 11 11 2 11 11 2 9 1 0 14 13 4 2
38 11 1 9 9 13 1 1 9 1 11 11 11 1 1 11 11 2 9 11 11 2 9 11 2 9 11 11 11 7 9 11 11 11 1 9 0 13 2
22 11 1 9 9 11 11 1 11 1 11 9 1 0 9 9 1 11 1 0 13 4 2
21 15 11 11 2 11 2 7 11 11 1 9 1 0 9 1 1 10 9 13 4 2
26 9 11 1 13 16 9 7 9 2 11 2 11 2 11 2 1 9 7 9 1 15 10 9 13 4 2
20 15 10 9 1 9 0 13 16 15 9 1 14 11 11 1 1 9 13 4 2
15 15 13 16 11 11 1 9 1 14 11 1 9 13 4 2
26 15 9 1 0 9 9 1 9 9 1 0 13 4 13 16 15 13 1 9 1 9 1 9 13 4 2
23 9 9 14 10 9 14 13 2 15 9 1 9 1 9 2 9 7 9 14 0 13 4 2
19 15 15 14 13 16 9 1 9 9 1 10 9 13 1 10 9 13 4 2
22 15 13 16 11 1 9 1 0 11 11 11 1 15 11 11 11 11 1 0 13 4 2
16 7 15 1 15 11 13 1 12 9 1 10 1 9 13 4 2
48 15 13 16 9 1 9 13 4 16 15 15 9 14 13 4 16 15 15 9 9 1 0 9 1 13 13 1 9 1 9 13 16 3 2 3 9 1 9 1 9 9 1 0 9 13 4 4 2
34 11 11 1 9 9 1 9 13 1 1 13 9 1 11 1 11 1 12 9 1 13 0 13 15 1 9 1 13 9 1 1 13 4 2
11 10 3 0 9 1 9 1 9 13 4 2
16 11 7 11 1 1 9 13 14 10 9 0 9 13 13 4 2
13 0 9 1 11 1 12 9 1 0 13 4 4 2
10 13 4 16 9 1 9 14 12 13 2
14 15 9 1 11 7 11 1 11 1 9 13 4 4 2
23 11 1 13 9 1 1 9 9 1 9 1 10 9 13 1 3 11 1 0 9 13 4 2
22 15 1 1 11 9 1 9 9 1 9 11 11 7 11 11 0 9 1 9 1 13 2
19 10 9 11 1 11 11 1 11 11 11 11 1 9 9 1 0 13 4 2
15 11 1 9 14 12 9 11 9 1 11 1 1 0 13 2
35 10 9 1 11 11 7 11 11 1 10 9 13 4 4 16 10 9 1 14 12 9 13 4 2 15 9 9 1 9 13 1 9 1 13 2
41 10 3 11 11 7 11 11 1 9 1 9 9 9 11 1 0 13 16 15 11 9 1 9 13 4 2 16 10 9 1 11 9 1 9 13 14 0 13 4 4 2
16 0 13 16 10 9 11 1 13 1 3 11 1 14 13 4 2
23 11 11 7 11 11 1 13 16 10 3 9 1 14 9 13 4 16 10 9 9 9 13 2
11 9 13 14 9 1 15 1 9 13 4 2
10 10 9 15 9 9 0 13 4 4 2
15 10 3 9 1 13 9 1 9 11 11 1 3 13 4 2
23 15 13 11 11 1 9 13 4 7 9 11 2 11 1 1 11 11 11 1 1 13 4 2
15 9 13 14 10 12 9 15 0 9 13 9 1 13 4 2
28 3 1 11 1 9 1 9 1 13 4 7 11 1 9 13 1 9 1 15 1 11 11 11 1 9 13 4 2
21 9 1 9 13 1 9 9 9 11 11 11 11 13 4 7 0 9 1 9 13 2
23 13 4 16 9 1 1 14 12 9 0 9 13 2 15 15 9 1 9 13 13 4 4 2
8 10 9 1 0 13 4 4 2
14 9 1 9 1 9 1 9 11 7 11 13 4 4 2
13 9 9 1 11 13 0 9 9 1 9 14 13 2
17 13 4 16 11 9 1 9 1 10 9 1 15 9 3 14 13 2
17 11 11 11 2 11 2 9 9 1 9 1 13 9 9 1 13 2
12 15 9 9 1 1 14 0 9 14 13 4 2
29 9 9 1 10 9 13 1 9 0 13 4 4 15 9 9 1 1 14 0 9 1 9 1 1 1 0 13 4 2
16 10 9 9 9 1 9 1 13 1 1 9 13 4 4 4 2
30 11 11 11 1 0 9 1 1 9 1 1 9 13 4 4 9 14 1 12 9 9 1 1 12 9 1 13 4 4 2
13 9 9 1 13 7 10 9 13 14 4 4 4 2
18 15 10 13 1 1 9 2 9 1 9 13 2 7 9 0 14 13 2
14 15 1 9 9 1 0 9 13 1 9 13 4 4 2
22 16 15 0 9 1 9 1 13 9 9 7 0 9 1 9 13 16 9 15 3 13 2
22 11 1 9 1 13 13 16 10 9 1 0 9 1 1 12 0 9 1 9 13 4 2
20 15 9 9 1 9 13 1 13 0 9 1 9 1 9 2 9 0 13 4 2
15 9 1 9 9 9 7 9 9 9 1 9 14 13 4 2
27 11 11 1 11 1 11 1 11 9 1 11 9 1 13 0 9 1 9 1 9 0 13 1 9 13 4 2
21 9 1 9 11 9 1 1 11 1 11 11 1 0 9 9 1 13 1 13 4 2
23 11 1 9 11 11 11 1 1 0 13 4 9 1 9 1 1 9 1 0 9 0 13 2
32 10 9 1 9 11 1 11 9 1 9 12 9 1 9 7 0 2 0 9 2 11 11 11 11 11 2 1 9 0 13 4 2
34 9 1 13 16 0 0 9 1 10 9 1 9 9 9 9 1 9 1 0 13 4 4 7 9 1 1 0 9 1 11 13 4 4 2
19 9 1 13 16 10 9 1 9 1 15 9 9 11 1 9 13 4 4 2
30 11 1 15 9 1 13 16 9 1 9 1 9 11 1 13 4 4 7 15 9 0 9 1 9 1 14 13 4 4 2
26 9 1 9 1 9 9 1 0 9 1 1 11 1 11 11 1 11 11 1 1 12 9 9 9 13 2
18 10 9 11 11 1 9 12 9 9 13 0 9 9 12 9 11 13 2
18 9 1 10 9 11 11 2 11 2 11 2 11 7 11 9 1 13 2
24 9 1 10 9 11 1 11 11 11 1 9 12 9 13 4 0 9 9 12 9 11 11 13 2
24 0 9 1 13 2 13 14 12 9 0 11 11 11 2 11 2 1 9 1 9 13 4 4 2
28 11 7 11 1 11 1 11 9 1 11 11 11 1 9 1 9 1 1 12 0 9 1 9 1 9 13 4 2
13 9 1 0 9 1 10 9 1 11 9 1 13 2
23 11 1 9 1 1 11 1 9 2 9 1 11 1 9 1 9 1 0 9 1 9 13 2
38 9 1 1 0 0 9 1 9 9 11 11 7 9 9 11 11 1 9 13 10 9 1 15 9 1 13 9 1 9 1 9 1 0 13 1 1 13 2
22 3 2 11 11 11 11 11 11 11 11 11 1 9 1 10 9 13 4 1 0 13 2
17 15 13 13 16 9 11 9 1 9 1 9 1 14 13 4 4 2
14 15 1 0 0 7 0 9 9 13 1 0 9 13 2
15 16 2 9 1 11 11 11 1 9 1 9 13 4 4 2
17 9 9 11 11 11 1 14 10 9 1 9 1 9 14 13 4 2
30 0 11 7 11 9 1 0 9 13 1 1 10 9 1 9 1 11 1 0 9 1 11 1 9 13 1 9 13 4 2
24 9 1 0 9 9 16 0 0 7 0 2 9 9 13 4 2 16 11 1 9 13 0 13 2
14 15 13 11 1 11 1 13 1 9 9 13 4 4 2
31 9 1 0 9 11 11 1 13 16 16 11 1 9 9 1 15 9 13 2 16 9 11 11 15 9 13 1 1 0 13 2
12 9 1 1 10 9 1 9 13 4 4 4 2
14 15 13 16 9 9 1 10 9 1 9 13 4 4 2
9 15 1 14 10 9 0 13 4 2
9 7 10 15 1 9 13 4 4 2
12 15 2 15 10 9 1 14 9 13 4 4 2
15 11 1 10 9 1 3 9 13 1 9 0 13 4 4 2
37 9 1 9 13 15 13 11 11 1 9 1 10 9 1 9 1 9 9 1 3 13 4 4 16 15 11 1 1 9 9 13 1 9 1 14 13 2
11 15 1 9 1 9 1 9 13 4 4 2
40 9 1 9 1 9 13 1 1 15 13 9 2 9 9 9 9 11 11 7 0 9 11 11 11 1 12 9 1 0 9 7 9 1 0 9 1 1 9 13 2
13 9 1 9 1 13 11 7 11 1 0 9 13 2
32 11 1 9 3 11 2 11 1 9 13 1 9 1 13 2 3 11 7 11 2 11 2 1 11 1 9 13 1 9 13 4 2
17 16 10 9 1 0 9 1 12 14 9 9 13 1 9 13 4 2
42 0 3 9 1 0 9 1 13 13 16 16 11 1 13 9 1 1 9 9 1 9 13 4 16 12 9 1 9 13 1 1 9 9 9 1 12 12 9 1 9 13 2
25 9 1 13 4 16 0 9 9 1 9 2 9 9 1 9 7 9 9 1 9 1 14 9 13 2
33 15 1 9 1 9 13 16 13 1 9 1 9 9 9 9 9 1 10 9 0 13 4 16 15 0 9 1 9 0 14 13 4 2
28 11 11 1 9 1 9 9 11 11 11 11 2 9 9 11 11 11 7 0 0 9 1 1 9 1 9 13 2
31 11 2 11 11 11 11 11 7 0 9 11 11 11 1 0 11 1 0 0 9 1 9 7 9 1 0 0 9 14 13 2
20 11 0 13 1 3 11 11 1 9 1 13 16 15 15 9 9 1 0 13 2
17 7 15 9 1 0 9 1 1 1 15 14 13 1 9 13 4 2
25 11 9 7 0 9 11 11 1 9 11 1 1 11 1 9 9 9 9 1 9 1 9 13 4 2
8 9 1 15 9 13 4 4 2
16 9 1 11 11 1 10 9 1 1 0 13 1 13 4 4 2
14 15 0 13 7 15 9 1 9 1 13 4 4 4 2
12 15 9 1 1 11 11 13 1 9 13 4 2
20 11 9 1 9 11 11 7 15 9 11 9 14 12 9 9 9 9 9 13 2
9 15 1 12 9 14 9 13 4 2
23 11 1 14 9 1 9 14 13 2 7 15 9 11 1 9 1 13 1 0 9 13 4 2
20 15 9 9 1 0 9 1 9 9 1 9 1 3 1 9 1 0 13 4 2
31 9 9 1 9 9 13 14 11 1 9 11 11 11 1 11 7 11 1 1 1 9 1 9 13 15 9 1 9 13 4 2
31 9 1 11 1 9 9 13 4 9 7 9 1 9 13 16 15 11 7 11 1 0 9 1 9 1 13 1 9 0 13 2
31 9 1 11 7 11 1 9 1 0 9 11 11 2 11 11 11 7 11 11 1 1 11 11 1 0 13 1 9 13 4 2
19 11 11 1 1 1 14 9 11 11 11 1 15 0 13 1 9 13 4 2
11 10 9 1 14 9 11 11 1 9 13 2
21 9 1 13 1 3 11 7 11 1 0 2 0 9 9 1 9 0 13 4 4 2
29 11 1 11 11 11 11 11 1 10 9 1 0 9 1 0 13 1 9 1 11 11 1 0 9 0 13 4 4 2
19 9 1 13 13 16 0 9 0 13 7 15 3 14 9 1 13 4 4 2
17 10 9 1 13 1 1 11 11 1 11 11 1 9 13 4 4 2
23 11 11 11 1 11 11 11 11 11 9 1 9 1 1 11 11 1 1 9 13 13 4 2
19 9 13 4 16 9 1 9 2 9 2 9 14 1 9 1 9 13 4 2
20 9 1 1 2 9 1 9 1 9 13 1 1 9 1 9 1 9 13 4 2
19 9 1 13 4 10 9 1 12 0 9 0 13 1 9 13 4 4 4 2
31 11 11 11 11 11 1 12 9 1 13 16 0 12 9 1 9 1 9 1 9 13 1 9 1 9 1 0 9 13 4 2
23 9 1 9 11 11 1 1 10 9 9 1 12 9 1 1 9 1 14 12 12 9 13 2
13 15 9 13 16 9 1 9 1 12 9 9 13 2
9 0 9 1 9 9 1 9 13 2
11 11 7 11 11 10 9 1 10 3 13 2
46 11 1 13 16 9 1 12 12 9 1 10 0 13 7 15 0 9 1 9 14 13 4 4 4 7 11 11 11 2 11 11 11 11 7 11 11 1 1 9 9 14 9 13 4 4 2
17 15 13 16 10 9 1 12 0 9 0 13 1 9 13 4 4 2
20 11 1 13 16 9 1 9 1 1 9 9 9 1 9 1 9 13 4 4 2
20 15 9 0 13 4 4 7 9 1 0 9 1 15 0 13 4 1 9 13 2
41 15 13 16 9 1 9 1 10 9 1 9 2 9 1 9 2 10 9 1 1 9 2 9 9 2 9 2 9 1 9 7 15 9 1 13 1 9 13 4 4 2
35 11 11 11 11 11 1 1 12 9 1 9 1 1 9 1 12 9 9 15 13 15 0 9 14 13 4 7 12 9 1 13 14 14 4 2
21 12 9 9 1 9 14 15 0 0 9 1 13 4 7 12 9 9 1 9 13 2
17 11 11 11 1 9 1 13 1 3 0 9 1 9 1 9 13 2
22 3 12 9 9 13 9 1 9 1 9 1 9 1 13 1 9 1 9 0 14 13 2
11 9 1 13 9 9 13 7 9 13 4 2
13 9 9 1 11 13 3 2 7 15 9 13 14 2
24 10 11 11 11 1 11 1 9 0 9 13 4 2 15 11 9 9 1 1 3 13 4 4 2
11 10 9 11 11 11 1 14 13 1 13 2
11 0 9 1 9 1 15 14 9 13 4 2
18 11 1 9 1 1 0 9 1 9 9 1 9 1 13 9 1 13 2
17 10 0 9 1 9 1 9 1 9 1 9 9 1 13 13 4 2
29 11 1 9 1 14 1 14 11 11 11 1 9 1 9 0 13 4 4 7 12 9 1 0 9 1 9 13 4 2
22 7 11 9 10 9 1 15 0 9 1 9 13 15 9 1 14 10 9 1 9 13 2
16 3 9 1 0 9 0 13 2 7 9 13 14 9 13 4 2
15 16 9 1 1 9 1 13 1 9 1 9 1 9 13 2
24 11 11 11 11 11 1 9 11 11 1 13 16 2 2 15 1 1 14 9 9 13 4 4 2
16 16 15 14 13 16 9 15 13 16 15 15 13 1 0 13 2
35 15 15 14 13 16 9 1 10 9 3 13 4 2 16 10 9 15 13 4 16 9 9 1 10 9 11 1 3 1 1 9 14 13 4 2
12 7 15 9 1 9 1 13 1 1 9 13 2
9 3 1 10 9 11 1 0 13 2
14 7 0 3 1 0 9 9 1 1 14 13 4 4 2
11 9 1 9 1 1 9 0 13 4 4 2
27 3 14 11 11 1 14 9 13 1 9 2 9 11 11 7 11 1 13 13 16 9 13 9 14 13 4 2
13 9 1 1 2 8 15 14 0 13 1 9 13 2
12 15 9 13 4 4 9 1 9 1 13 1 2
17 11 11 11 1 11 11 15 9 1 1 9 1 1 11 11 13 2
23 11 11 11 1 11 11 1 11 11 1 13 13 16 9 1 0 13 9 1 9 14 13 2
8 9 15 0 13 15 9 13 2
14 0 3 9 1 9 13 1 1 9 1 9 13 4 2
20 9 1 10 9 1 9 9 13 4 4 7 9 1 15 1 13 4 4 4 2
22 11 1 11 11 1 13 0 9 9 1 9 1 9 1 9 1 0 13 1 9 13 2
13 9 1 9 1 1 15 9 13 9 13 4 4 2
13 15 14 9 1 9 1 9 14 13 1 9 13 2
16 9 2 9 1 9 1 1 10 9 1 9 9 13 4 4 2
33 11 1 11 1 1 9 9 13 1 9 13 4 11 1 11 1 12 9 1 0 13 4 16 15 9 0 13 1 9 15 14 13 2
30 11 9 11 11 1 11 1 9 0 13 1 12 9 1 9 13 4 11 1 15 13 16 15 14 9 9 1 1 13 2
23 11 1 11 1 9 1 9 9 1 9 13 4 13 16 15 1 15 1 9 13 4 4 2
10 15 11 9 1 12 0 9 14 13 2
11 15 9 1 9 0 9 1 14 0 13 2
15 15 13 16 0 9 1 9 7 9 1 9 15 13 4 2
31 11 1 13 16 9 1 9 1 13 9 1 15 15 1 11 1 9 14 13 4 7 13 16 9 13 1 15 3 9 13 2
33 11 1 9 1 0 9 1 9 1 11 1 13 16 10 15 9 14 13 16 0 9 1 13 1 9 1 9 1 9 13 4 4 2
27 11 9 1 9 13 4 11 1 13 16 11 0 14 13 16 15 2 9 2 13 2 15 0 0 9 13 2
14 13 4 9 1 9 13 4 7 15 0 9 13 4 2
11 11 11 1 9 1 9 1 9 13 4 2
11 11 2 11 1 0 9 0 13 4 4 2
8 9 1 9 1 9 0 13 2
17 15 10 9 1 14 11 1 9 7 15 9 1 12 9 13 4 2
15 10 15 1 9 9 1 9 1 1 11 13 4 4 4 2
24 15 13 16 11 1 9 2 11 11 2 1 9 13 11 11 9 1 9 1 9 1 0 13 2
18 11 1 9 13 16 11 1 11 1 9 13 4 9 1 9 13 4 2
7 10 15 0 9 14 13 2
10 0 11 1 9 1 9 3 0 13 2
24 9 11 11 11 1 13 13 16 15 15 9 1 9 1 14 12 9 11 13 1 9 13 4 2
18 0 13 16 11 1 0 9 9 11 11 1 9 13 1 9 13 4 2
14 15 13 16 15 0 9 1 0 9 1 0 13 4 2
26 9 11 1 13 16 15 15 9 1 11 11 11 2 11 2 1 9 1 15 9 1 9 14 13 4 2
18 15 11 1 13 16 9 1 12 9 11 13 1 15 9 1 9 13 2
15 15 13 16 11 11 1 9 11 1 10 9 1 13 4 2
22 11 1 9 1 9 1 9 0 13 4 4 14 16 0 11 11 1 9 9 13 4 2
8 9 1 9 11 1 13 4 2
28 3 2 0 9 9 11 11 11 1 9 1 9 2 9 2 9 2 10 9 1 9 2 1 9 9 13 4 2
11 15 15 11 11 1 9 1 13 4 4 2
39 11 11 11 11 1 0 11 11 1 11 1 0 9 1 12 9 1 15 1 1 10 0 9 13 16 10 9 1 15 0 13 4 2 9 13 7 9 13 2
35 12 0 11 11 1 1 1 11 1 9 13 16 15 0 9 1 0 9 11 11 13 7 15 1 11 1 11 7 11 1 9 9 13 4 2
18 15 9 1 9 1 9 13 4 2 15 0 11 11 1 14 0 13 2
29 0 9 1 10 12 9 1 15 9 13 2 15 13 9 9 11 11 2 9 2 7 11 11 11 2 9 9 2 2
25 12 9 1 13 10 9 1 11 11 1 15 9 2 9 7 9 1 0 9 1 1 1 9 13 2
9 9 9 1 15 0 9 1 13 2
15 11 1 9 1 13 16 15 15 12 9 1 9 13 4 2
14 10 3 15 15 9 7 9 1 1 1 0 9 13 2
21 15 15 9 1 1 14 12 9 13 4 2 15 9 11 1 13 1 9 13 4 2
21 0 13 16 11 1 9 1 15 11 1 9 13 4 1 0 9 1 9 13 4 2
27 9 1 9 1 10 0 2 0 0 9 1 10 9 1 13 2 15 11 7 11 12 0 9 13 4 4 2
27 10 9 1 1 11 1 9 14 13 4 15 15 9 1 13 4 2 16 15 11 1 12 9 1 0 13 2
26 15 1 1 0 13 4 9 9 1 1 11 13 4 2 15 15 9 1 1 15 9 0 13 4 4 2
21 11 1 11 1 13 1 9 11 1 15 13 15 11 1 3 12 9 10 9 13 2
19 15 1 11 11 11 11 1 0 9 1 1 14 0 11 11 1 9 13 2
39 7 11 1 0 0 11 11 1 13 13 16 11 1 15 0 9 1 9 1 9 13 4 2 16 11 1 13 13 16 10 9 13 1 1 15 0 13 4 2
20 15 9 1 9 9 1 1 1 14 0 9 1 9 0 2 0 9 13 4 2
35 11 11 11 11 11 1 13 13 16 11 1 10 9 0 13 1 9 13 7 11 11 11 11 11 1 13 13 16 11 1 10 9 14 13 2
20 0 9 11 1 11 11 1 11 1 11 11 1 0 9 1 9 13 4 4 2
12 10 9 1 0 9 11 1 12 10 9 13 2
11 0 9 11 10 11 11 1 13 4 4 2
19 0 9 14 12 2 12 9 1 13 10 0 9 15 9 13 1 0 13 2
30 11 1 12 9 1 11 11 1 11 11 1 13 4 4 7 15 1 15 14 0 9 1 9 1 9 14 13 4 4 2
16 11 7 11 1 1 13 9 1 11 1 12 9 10 13 4 2
28 9 1 15 2 15 1 9 1 0 10 9 7 9 0 13 4 9 1 0 11 11 1 13 1 9 13 4 2
20 12 9 9 1 13 13 1 3 14 15 0 9 13 1 1 13 0 9 13 2
41 12 9 1 13 9 9 9 1 9 1 1 11 1 0 9 9 1 12 9 1 9 7 9 0 13 4 9 1 9 0 13 1 1 0 9 0 13 1 9 13 2
13 9 1 1 10 9 1 9 1 9 13 0 13 2
49 11 11 11 11 11 1 11 11 11 11 11 1 1 12 0 9 9 1 13 16 12 9 15 15 15 14 0 9 1 9 1 3 0 13 7 15 12 9 1 1 15 1 9 1 13 1 9 13 2
16 15 1 1 0 9 11 1 9 9 1 9 1 9 13 4 2
30 11 1 0 9 1 13 4 13 16 12 9 1 9 1 9 0 13 7 9 1 9 13 1 14 3 0 13 4 4 2
12 11 1 0 0 9 1 3 14 0 9 13 2
14 9 1 0 9 1 9 7 9 1 14 9 13 4 2
19 11 1 11 1 11 11 1 12 3 0 9 7 9 1 9 11 1 13 2
12 11 1 14 12 9 1 9 11 1 13 4 2
11 15 0 0 9 1 9 1 13 9 13 2
19 0 9 15 13 16 0 9 1 15 1 1 12 14 9 14 13 4 4 2
27 0 9 1 9 1 11 1 13 16 15 13 1 1 12 9 1 11 11 11 3 14 12 9 1 9 13 2
19 15 1 12 0 0 9 0 13 4 7 9 13 1 1 0 9 13 4 2
20 10 9 1 11 7 11 1 11 11 1 9 0 9 9 13 9 1 9 13 2
13 12 9 9 1 9 1 9 2 9 13 4 4 2
32 12 9 1 9 9 1 10 9 1 9 13 16 0 9 1 9 13 1 9 1 1 9 7 9 1 9 2 9 13 4 4 2
25 12 9 15 1 14 0 13 16 11 1 0 9 11 7 11 1 11 11 11 1 0 9 13 4 2
18 15 1 3 14 12 0 9 1 9 0 9 1 12 9 0 13 13 2
20 15 0 9 14 13 2 7 9 1 15 0 9 1 13 16 15 9 13 4 2
39 15 13 13 0 9 1 2 7 9 9 1 9 1 9 0 14 13 2 15 1 9 7 9 1 1 9 13 7 9 13 1 1 14 0 13 4 4 4 2
12 9 11 9 1 9 1 1 9 13 4 4 2
34 0 9 1 9 13 7 9 13 9 11 7 9 1 13 4 7 11 11 11 1 11 11 1 1 9 0 13 15 9 1 0 13 4 2
9 7 9 1 10 9 3 0 13 2
23 16 15 15 9 7 9 1 9 1 9 13 4 4 16 15 1 15 9 14 13 4 4 2
26 11 1 1 2 9 2 13 1 12 9 13 2 7 9 1 1 10 9 9 1 0 9 13 4 4 2
22 9 7 15 9 1 9 1 15 9 13 4 4 16 9 9 13 15 0 13 4 4 2
23 0 9 15 9 13 1 1 9 1 9 13 4 2 15 15 1 9 1 9 13 4 4 2
14 9 7 9 1 15 9 1 9 13 15 9 14 13 2
23 9 11 7 9 11 11 11 11 1 13 13 16 9 15 9 1 1 9 1 9 13 4 2
20 9 1 9 1 1 12 2 12 9 1 14 11 11 1 9 14 13 4 4 2
36 11 11 1 9 13 4 9 1 0 12 9 9 7 12 9 1 9 13 4 4 7 9 0 13 1 14 9 9 1 0 9 13 4 4 4 2
43 9 1 11 11 7 11 11 1 11 11 2 11 11 2 11 11 2 11 11 7 11 11 1 11 11 11 1 11 11 1 1 12 9 1 9 13 1 9 1 0 13 4 2
11 15 1 11 11 11 1 9 0 13 4 2
23 15 9 9 14 13 16 15 9 1 9 14 13 7 15 9 1 1 1 9 13 4 4 2
18 10 9 1 9 11 11 1 13 4 2 15 9 9 1 9 13 4 2
34 0 9 8 13 11 1 9 2 11 11 11 11 2 1 9 1 9 9 16 9 9 13 1 9 1 13 1 9 1 13 9 0 13 2
11 7 10 9 1 9 1 9 10 13 4 2
30 9 14 1 13 4 12 9 1 1 0 9 1 13 13 16 9 1 0 12 9 1 1 9 1 9 10 13 4 4 2
16 9 1 15 2 9 9 2 16 2 9 9 2 9 13 4 2
47 11 1 11 1 0 2 0 9 1 11 1 9 1 9 1 9 9 13 13 4 16 10 9 9 1 9 9 1 3 10 13 4 2 10 9 14 3 1 1 9 1 10 14 9 13 4 2
19 0 12 9 1 9 1 13 1 9 1 9 1 3 1 1 9 13 4 2
32 9 14 1 13 10 9 1 15 13 4 16 11 1 9 1 1 1 9 1 9 1 12 1 1 12 9 1 1 9 13 4 2
17 9 11 1 13 9 1 1 13 9 1 9 0 9 13 4 4 2
43 11 11 7 11 11 11 11 1 9 1 0 9 11 11 11 1 10 9 1 9 13 4 15 15 9 1 0 9 1 9 1 0 13 1 9 1 9 1 0 13 13 4 2
27 10 2 9 2 1 9 13 9 1 9 13 4 16 0 12 9 1 1 9 1 14 12 9 9 13 4 2
27 16 9 10 9 1 12 9 14 13 16 9 1 10 13 9 0 9 13 7 9 1 1 15 13 4 4 2
28 10 9 1 15 14 13 13 16 9 1 13 1 9 7 0 9 2 9 9 2 13 1 9 1 9 13 4 2
19 9 9 1 10 9 9 13 4 13 4 15 0 9 9 1 13 4 4 2
14 15 14 9 1 9 10 13 1 12 9 13 4 4 2
15 15 13 16 0 9 2 9 1 15 0 9 13 4 4 2
35 0 9 13 0 9 1 9 1 11 15 0 9 1 13 1 9 14 13 4 4 16 11 1 3 0 9 1 11 1 9 1 0 13 4 2
15 9 1 9 2 9 7 9 9 1 3 0 9 13 4 2
21 9 1 1 10 9 1 1 0 7 0 9 12 9 1 14 10 9 1 0 13 2
29 11 11 11 1 13 4 16 9 1 1 11 1 11 2 11 7 11 1 10 9 2 9 7 0 0 9 0 13 2
22 15 1 0 9 1 9 7 9 9 1 9 13 1 1 12 9 1 9 13 4 4 2
12 0 11 1 13 1 1 9 12 13 4 4 2
20 11 9 9 1 14 11 2 11 2 11 7 11 9 1 0 9 13 4 4 2
51 0 9 11 7 11 1 3 13 9 1 1 11 9 1 12 9 15 9 7 9 1 13 4 4 7 9 9 1 3 9 7 9 1 9 1 0 13 4 1 1 12 9 9 9 7 9 9 1 13 4 2
13 9 13 1 3 9 9 3 2 3 0 13 4 2
15 9 9 1 13 1 1 11 11 1 0 13 4 4 4 2
14 9 1 9 1 9 1 1 14 13 1 9 13 4 2
12 0 11 9 1 9 9 0 13 4 4 4 2
23 11 11 11 11 11 1 13 4 16 0 9 1 1 9 1 10 9 0 9 13 4 4 2
12 9 9 1 9 1 14 9 13 4 4 4 2
8 10 9 9 1 13 4 4 2
20 11 11 1 11 1 0 13 1 0 9 1 10 9 1 0 13 4 4 4 2
30 0 9 1 1 11 1 1 1 9 1 9 1 9 14 13 4 2 7 15 1 13 7 0 13 1 15 9 14 13 2
23 11 1 0 9 11 11 1 11 1 13 16 11 11 11 7 11 11 1 9 15 9 13 2
12 0 9 1 9 1 15 9 1 3 13 4 2
33 7 11 11 11 11 1 0 9 1 13 4 9 1 11 1 13 16 9 15 9 1 0 13 2 16 15 0 9 1 0 13 4 2
10 9 1 9 10 9 1 0 13 4 2
20 15 13 16 11 1 11 1 9 9 1 10 9 13 4 2 15 15 1 13 2
20 15 11 9 1 9 10 9 1 9 13 4 7 15 9 1 9 13 4 4 2
18 15 13 16 15 11 1 9 2 9 7 9 1 9 1 14 9 13 2
16 15 11 1 0 2 0 7 12 0 9 1 1 1 0 13 2
9 11 7 11 1 9 15 9 13 2
22 11 1 13 16 11 15 10 0 9 1 1 14 3 13 2 10 9 15 9 13 4 2
11 15 1 15 15 14 13 1 9 13 4 2
17 15 13 16 15 11 11 1 9 9 9 13 1 3 15 9 13 2
14 15 10 9 1 9 13 16 11 1 15 0 9 13 2
15 11 1 1 10 14 9 13 2 15 11 1 0 9 13 2
15 9 1 9 15 9 2 9 7 0 2 0 9 3 13 2
11 15 0 13 16 10 0 9 0 13 4 2
7 15 15 10 9 13 4 2
24 10 9 15 15 13 2 15 15 9 13 4 16 0 10 9 11 0 9 1 9 1 13 4 2
14 15 9 13 16 9 1 0 9 1 9 0 13 4 2
11 15 9 1 1 1 9 0 14 13 4 2
10 9 1 9 1 1 10 0 13 4 2
21 12 9 1 9 1 15 9 13 16 15 9 1 1 14 9 9 1 14 13 4 2
16 7 15 9 0 9 0 13 7 15 0 9 1 0 13 4 2
38 9 11 11 9 1 10 12 9 1 0 13 15 11 11 11 1 9 1 1 9 13 1 1 9 11 1 2 11 11 2 11 11 2 1 1 13 4 2
38 2 11 11 2 11 11 2 1 9 1 11 2 11 11 1 1 11 11 11 1 0 9 1 9 11 11 1 11 1 9 1 13 16 11 9 14 13 2
12 15 9 1 9 1 1 12 9 13 4 4 2
18 11 1 13 16 11 11 1 10 9 1 1 9 14 13 4 4 4 2
25 0 9 15 15 9 9 7 9 1 0 13 4 4 16 15 9 1 15 9 1 1 0 14 13 2
39 0 13 16 11 11 11 1 0 9 13 4 9 1 1 13 4 16 11 1 12 9 1 11 9 12 1 13 15 9 1 9 13 4 10 9 13 4 4 2
11 0 12 9 1 11 11 7 11 11 13 2
16 9 1 0 13 1 3 11 1 9 1 1 9 13 9 13 2
20 11 2 11 11 9 1 12 0 9 7 9 1 10 9 1 1 13 4 4 2
13 11 1 13 16 12 9 1 1 10 9 13 4 2
28 9 1 9 7 15 9 7 0 9 1 9 1 9 1 1 11 11 11 11 2 11 2 0 9 13 4 4 2
18 10 9 1 3 13 4 9 1 11 11 1 9 9 1 9 13 4 2
24 9 1 9 1 9 2 9 9 1 9 2 9 9 7 0 9 1 13 9 1 9 13 4 2
24 11 1 11 11 1 13 1 9 1 10 9 1 0 9 9 7 10 0 9 1 9 13 4 2
11 9 9 12 9 1 9 12 9 1 13 2
27 12 9 9 1 12 9 9 1 9 1 9 13 7 9 12 9 1 12 9 1 0 9 1 9 13 4 2
26 9 1 9 1 9 0 9 1 1 11 11 11 11 1 9 13 7 10 9 1 11 1 9 13 4 2
20 12 12 1 0 7 0 0 9 9 11 11 11 1 0 9 1 13 4 4 2
17 11 11 2 11 7 11 1 9 15 0 12 9 1 13 4 4 2
38 11 11 11 11 1 9 1 11 1 9 13 16 9 13 14 11 1 9 1 0 9 7 11 11 1 13 11 1 9 1 1 13 12 0 9 9 13 2
19 7 11 1 9 1 14 9 9 11 11 1 9 1 0 9 1 13 4 2
24 11 1 13 16 11 1 0 13 1 14 3 9 9 9 13 4 15 15 11 1 9 9 13 2
20 10 0 9 1 9 1 1 11 11 7 11 1 14 11 1 9 13 4 4 2
14 15 13 16 11 1 12 9 9 1 9 1 9 13 2
15 15 1 15 1 11 11 7 11 1 14 10 0 9 13 2
28 0 13 16 11 11 7 11 1 9 1 15 1 1 9 13 1 1 1 12 2 12 12 9 1 9 13 4 2
23 7 11 1 14 15 9 1 9 13 1 1 12 12 1 0 9 13 1 9 13 4 4 2
30 15 1 12 0 9 1 11 2 11 2 1 12 10 0 9 11 11 1 11 1 11 9 1 12 9 1 0 13 4 2
24 11 1 9 9 9 1 9 1 1 11 11 1 9 9 1 12 9 1 0 9 13 4 4 2
24 9 9 1 9 11 11 1 1 9 12 2 12 9 1 1 14 9 9 1 9 13 4 4 2
16 10 9 1 12 9 1 9 1 9 9 1 12 9 13 4 2
20 11 11 0 13 4 1 9 13 1 9 1 12 9 1 9 9 13 4 4 2
20 9 9 11 11 11 1 9 1 12 9 1 9 1 9 9 1 9 13 4 2
29 15 0 13 16 11 1 11 11 11 1 11 11 7 11 11 1 12 9 1 1 9 9 1 0 13 4 4 4 2
40 9 1 9 9 11 11 2 0 9 11 11 7 9 9 11 11 1 9 13 4 16 16 11 15 0 9 1 9 14 13 4 16 15 9 14 0 9 13 4 2
12 11 1 9 1 9 9 11 11 1 9 13 2
28 3 2 12 9 1 9 1 13 4 16 9 9 1 9 13 1 9 1 11 11 1 9 9 9 13 4 4 2
29 0 13 16 9 9 0 13 4 1 9 13 1 0 9 9 1 10 9 1 9 9 1 9 13 1 9 13 4 2
13 9 12 2 12 9 1 1 9 0 13 4 4 2
17 0 9 1 1 11 1 0 9 11 11 1 11 1 9 13 4 2
17 15 11 11 1 11 0 9 1 9 1 14 12 9 0 9 13 2
15 9 1 15 1 13 4 11 10 9 14 15 1 14 13 2
6 11 15 14 9 13 2
10 11 11 1 9 1 12 9 14 13 2
20 0 9 1 13 16 11 11 1 11 1 14 9 15 0 9 14 13 4 4 2
26 11 11 1 0 11 11 1 12 1 10 9 13 4 7 15 15 0 9 1 1 0 9 13 4 4 2
12 10 0 9 1 15 9 1 9 13 4 4 2
20 0 11 1 11 11 11 1 0 13 11 11 1 11 11 11 14 13 4 4 2
9 3 2 11 11 15 9 9 13 2
31 11 11 11 2 11 2 1 0 9 11 11 11 1 13 4 16 11 11 11 1 1 1 15 9 1 0 9 1 13 4 2
29 15 13 16 16 15 9 1 3 9 13 4 4 16 15 11 7 11 1 1 11 1 9 1 0 13 1 9 13 2
19 15 11 9 1 9 13 16 15 9 1 9 1 9 1 14 13 4 4 2
43 11 1 11 1 11 11 1 0 9 9 9 13 1 3 9 1 9 1 11 1 10 9 1 9 13 16 11 11 1 1 11 1 9 1 1 15 9 9 1 9 13 4 2
26 15 13 16 2 15 15 15 1 10 9 1 1 0 13 16 15 15 9 1 3 14 0 14 13 4 2
8 15 9 1 0 9 1 13 4
16 15 3 13 16 2 15 11 1 1 1 14 12 9 13 4 2
34 15 15 11 11 11 1 9 1 1 0 13 4 4 15 15 15 9 13 4 16 11 11 2 11 1 11 1 9 1 11 1 15 13 4
30 15 11 9 1 9 1 9 1 9 1 14 13 1 9 13 4 13 16 10 9 1 11 11 11 1 9 0 14 13 2
27 0 13 16 9 1 9 1 1 11 1 0 9 1 13 4 16 15 11 1 1 9 1 15 9 14 13 2
25 16 2 15 15 14 9 13 16 9 1 9 12 0 9 13 7 15 1 9 13 1 0 13 4 2
17 0 0 9 1 9 1 15 0 9 9 1 9 1 9 9 13 2
13 9 1 0 0 9 1 0 13 9 10 9 13 2
13 10 9 1 11 1 9 1 9 9 13 4 4 2
19 11 1 15 0 9 1 0 12 9 1 9 9 7 0 9 1 9 13 2
24 9 1 0 0 9 1 13 4 0 0 9 9 1 0 12 9 1 1 13 1 9 13 4 2
16 10 9 1 1 10 9 1 11 1 3 12 12 9 13 4 2
22 11 11 1 0 0 9 1 9 1 9 1 9 1 9 13 1 9 1 0 9 13 2
9 15 11 9 11 11 14 9 13 2
36 9 1 1 11 11 11 11 11 1 13 16 11 1 9 1 9 1 13 9 1 13 4 9 1 0 9 1 9 13 1 9 1 9 13 4 2
22 15 13 16 9 0 9 1 0 13 1 1 3 9 1 0 13 1 9 1 14 13 2
13 15 0 9 1 10 9 1 9 13 1 9 13 2
16 11 1 9 14 1 9 0 9 1 9 1 13 1 9 13 2
30 15 9 13 16 0 9 1 0 12 9 1 1 1 10 9 1 0 12 9 1 0 9 1 12 9 1 9 13 4 2
23 15 13 16 11 7 11 11 1 0 9 1 9 13 4 2 7 0 9 1 9 13 4 2
23 11 1 0 9 1 9 1 9 13 4 15 13 16 15 9 9 1 1 0 13 4 4 2
18 15 9 1 1 2 11 11 2 9 1 9 9 9 9 13 4 4 2
15 9 1 0 9 11 1 1 14 11 1 14 9 0 13 2
13 15 0 13 9 15 0 9 1 9 13 4 4 2
15 9 1 11 1 9 1 9 1 0 9 1 13 1 13 2
20 11 1 13 16 9 1 0 9 1 9 1 9 0 9 1 13 14 4 4 2
13 15 13 16 9 1 15 0 9 10 0 13 4 2
24 15 13 16 9 1 0 7 0 9 9 1 13 9 9 1 9 1 9 13 1 13 4 4 2
46 9 1 11 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 11 2 11 11 2 11 2 11 2 11 7 11 1 1 11 11 11 11 7 9 9 1 0 9 0 13 2
34 11 11 11 11 1 10 9 1 9 13 1 3 9 13 4 16 0 9 1 9 0 13 7 15 14 15 1 1 0 9 14 13 4 2
11 10 0 9 1 1 1 9 13 0 13 2
28 9 1 0 9 1 13 9 1 9 13 1 9 13 4 2 16 15 1 10 9 9 1 1 3 14 13 4 2
32 0 9 1 13 1 1 9 13 12 13 4 4 7 11 1 0 9 1 9 1 10 9 13 4 7 15 9 12 13 4 4 2
19 10 9 9 1 9 14 13 4 2 7 9 1 9 1 15 9 13 4 2
34 11 11 1 9 9 2 9 9 2 11 11 11 1 13 16 9 1 9 1 12 9 0 13 4 2 15 9 12 1 12 1 13 4 2
13 11 11 11 11 1 15 9 1 9 1 9 13 2
9 9 9 1 9 13 4 4 4 2
9 15 12 9 9 14 13 4 4 2
15 10 9 2 9 9 7 0 9 0 9 9 13 4 4 2
10 9 9 1 14 0 13 4 4 4 2
23 11 11 11 1 1 12 9 9 9 13 4 4 15 1 12 9 9 15 13 4 4 4 2
17 9 14 11 11 1 9 1 1 9 9 13 1 9 13 4 4 2
36 11 11 1 9 11 11 1 13 16 11 2 11 2 11 7 11 1 9 13 1 9 1 15 11 11 1 9 11 11 1 14 0 13 4 4 2
18 9 13 11 1 11 1 11 11 1 0 9 1 1 1 9 13 4 2
29 9 9 11 1 11 11 1 14 11 11 11 11 1 9 13 9 1 9 13 7 9 9 1 1 1 9 13 4 2
14 11 1 11 11 1 14 9 1 1 1 9 13 4 2
15 9 1 11 11 1 12 9 1 14 0 13 4 4 4 2
32 11 2 11 11 1 11 11 1 11 11 11 7 11 1 0 9 1 1 9 9 1 15 1 9 13 4 1 9 13 4 4 2
15 9 1 1 11 11 1 15 12 10 9 1 0 13 4 2
22 15 1 14 11 11 1 0 9 9 1 9 13 4 9 9 1 9 12 13 4 4 2
16 11 11 11 1 11 1 0 9 1 9 13 1 9 13 4 2
29 9 1 13 13 16 11 11 11 2 11 2 9 0 9 9 1 13 1 1 9 1 9 1 9 1 13 4 4 2
18 11 1 11 9 1 9 7 9 1 0 9 1 1 1 9 13 4 2
22 15 13 13 16 10 9 1 11 1 9 1 9 0 9 1 9 1 0 9 13 4 2
16 9 1 1 2 9 1 9 1 9 1 9 1 9 13 4 2
13 11 1 13 13 16 11 1 0 9 0 13 4 2
10 11 3 0 9 1 9 13 4 4 2
36 11 9 11 11 1 1 2 11 2 11 11 2 11 1 11 9 11 11 1 9 1 9 1 9 1 9 7 9 1 0 9 1 9 13 4 2
18 11 1 9 1 0 11 1 15 14 9 1 10 9 1 9 14 13 2
13 3 2 11 1 10 9 1 15 9 0 13 4 2
23 15 13 16 15 12 0 2 0 9 1 9 13 7 9 1 9 1 11 1 0 9 13 2
15 11 1 11 1 15 9 1 9 1 9 1 9 13 4 2
20 11 9 1 13 16 0 9 9 1 0 13 1 1 11 1 10 9 13 4 2
10 15 11 1 0 13 9 1 0 13 2
18 15 11 9 1 9 1 9 9 1 0 13 9 1 0 9 13 4 2
33 11 1 0 9 1 9 1 12 9 9 7 11 11 11 1 12 9 9 9 1 9 1 9 0 9 9 1 13 1 0 9 13 2
21 11 9 1 13 13 16 9 9 1 1 11 11 1 14 9 9 1 9 13 4 2
18 15 10 9 1 10 9 13 7 15 9 9 1 9 1 1 1 13 2
11 11 1 10 9 0 9 1 9 13 4 2
12 7 15 15 0 9 1 0 9 13 4 4 2
17 11 1 9 1 9 1 9 1 1 1 15 9 1 0 13 4 2
13 11 1 10 9 1 9 1 9 1 14 9 13 2
14 15 13 16 10 9 1 11 9 1 9 13 4 4 2
16 7 15 1 1 15 9 10 9 1 9 1 9 13 4 4 2
32 9 1 13 13 16 0 9 9 1 0 13 1 1 10 9 1 9 1 9 13 1 9 1 9 7 0 9 1 9 13 4 2
30 11 7 11 1 9 0 9 1 9 13 1 3 11 11 11 1 9 13 16 9 9 7 9 1 1 10 0 9 13 2
15 15 13 16 9 10 0 9 1 0 10 9 1 9 13 2
22 15 15 13 1 3 9 9 1 11 11 1 1 3 12 12 9 13 1 9 13 4 2
13 9 15 11 1 1 12 12 9 1 9 13 4 2
20 11 1 13 16 15 11 7 11 1 9 1 9 13 15 9 1 1 9 13 2
21 11 1 13 16 9 1 0 9 0 11 11 1 9 7 9 1 10 9 9 13 2
24 11 1 13 16 11 1 11 11 11 11 1 10 0 9 1 1 12 12 12 9 0 13 4 2
25 15 1 11 11 11 11 1 9 1 1 13 4 9 1 0 9 1 12 2 12 12 9 13 4 2
38 15 1 11 1 11 9 1 11 1 11 11 1 9 7 0 9 1 9 1 1 11 11 1 13 2 2 10 9 13 4 4 15 0 14 13 4 4 2
22 7 2 9 10 9 1 0 9 1 3 9 9 13 1 1 10 9 1 9 13 2 2
40 11 7 11 1 9 0 9 1 12 0 9 1 0 9 11 1 11 11 1 13 16 11 7 11 1 0 9 1 3 2 9 9 2 13 1 1 9 13 4 2
14 0 13 16 11 1 9 1 9 1 12 9 13 4 2
22 11 1 15 9 0 9 1 9 9 1 1 1 0 12 12 9 9 1 9 14 13 2
15 15 1 15 11 9 1 11 7 11 9 9 1 14 13 2
23 15 15 9 1 15 15 15 13 4 9 1 9 7 9 14 1 9 1 9 1 9 13 2
29 11 1 9 9 1 0 9 1 13 1 3 11 1 9 13 16 10 9 1 0 13 4 9 1 9 0 9 13 2
37 11 11 1 11 1 0 9 1 9 13 4 9 1 9 1 9 13 4 13 2 2 15 15 15 9 13 13 4 16 15 15 10 9 1 9 13 2
29 11 7 11 1 11 1 9 1 12 9 1 9 1 1 14 9 9 1 9 2 9 1 14 12 9 1 9 13 2
22 15 1 11 11 1 9 1 12 0 9 13 4 16 16 11 1 9 1 0 9 13 2
35 11 11 11 11 7 11 1 11 11 11 1 9 1 9 9 1 13 12 9 1 11 1 11 1 9 11 11 7 9 11 11 1 9 13 2
17 9 1 10 12 9 1 12 9 1 1 0 9 13 1 9 13 2
19 15 12 9 1 1 9 9 1 1 14 9 7 9 14 1 14 9 13 2
28 10 12 9 1 1 11 2 11 11 1 1 1 13 4 1 11 1 1 11 1 9 9 9 1 10 9 13 2
23 11 1 1 10 0 9 9 9 13 1 1 12 9 1 9 9 1 9 13 1 9 13 2
20 12 9 1 10 9 9 9 1 1 12 9 1 11 11 1 1 14 9 13 2
19 9 9 1 0 10 9 1 11 9 1 1 11 15 9 14 9 13 13 2
26 10 9 1 11 1 11 11 11 11 1 13 16 11 1 9 1 0 9 0 9 1 9 13 4 4 2
17 0 0 11 1 1 10 0 9 1 13 4 0 11 1 9 13 2
30 9 9 11 11 1 15 0 9 1 11 1 9 9 2 9 9 2 1 9 13 0 15 9 1 3 9 13 4 4 2
38 9 9 1 11 1 10 9 1 9 13 4 13 16 0 9 10 9 1 9 13 4 16 11 1 11 11 1 12 9 9 1 0 9 1 9 13 4 2
17 10 9 1 1 14 15 9 1 1 15 9 11 1 1 13 4 2
34 9 9 1 9 9 1 12 0 9 1 13 16 2 15 10 9 1 0 9 13 16 11 1 9 1 1 15 9 11 1 1 13 4 2
8 11 1 15 0 9 13 4 2
35 2 9 1 1 2 9 9 1 13 9 1 13 4 4 16 11 1 11 1 11 11 1 12 9 1 9 1 1 12 9 1 9 13 4 2
61 0 13 16 9 1 1 11 11 1 11 2 11 11 11 1 11 1 0 2 0 2 9 1 9 13 1 3 11 11 1 11 1 3 0 9 11 11 1 11 1 1 9 0 13 7 11 2 11 11 11 2 1 10 9 1 1 9 14 9 13 2
17 9 9 1 9 11 11 11 1 9 9 9 1 14 3 13 4 2
20 9 1 9 13 16 9 9 1 9 11 11 11 11 1 9 1 13 4 4 2
32 16 2 10 9 1 9 1 1 9 9 11 7 9 2 3 1 9 1 11 1 0 2 0 2 9 1 9 13 1 13 4 2
21 10 9 13 16 11 1 15 11 1 9 13 0 9 1 0 9 1 13 4 4 2
26 9 1 9 9 1 9 13 4 0 9 9 1 9 13 1 9 7 9 1 9 1 9 13 4 4 2
20 9 1 9 9 1 13 4 16 10 14 10 0 12 9 1 9 14 13 4 2
12 15 11 11 1 9 1 9 1 9 13 4 2
16 15 1 14 9 9 1 9 1 9 1 9 1 9 13 4 2
17 11 11 11 11 1 11 1 13 2 9 9 14 13 4 4 4 2
26 9 9 1 9 1 9 13 4 16 9 9 1 9 1 9 1 0 9 9 1 9 1 13 4 4 2
21 11 1 13 16 0 9 1 0 9 1 9 10 9 12 9 14 9 1 13 4 2
46 13 4 4 4 16 11 1 15 0 7 0 9 1 10 13 1 9 1 15 1 9 13 4 4 2 7 11 11 1 13 1 9 9 1 1 1 15 1 1 15 9 14 13 4 4 2
18 11 1 13 16 15 0 9 13 16 9 9 1 1 9 1 9 13 2
34 9 9 11 11 1 13 16 9 9 9 7 9 1 9 1 9 1 1 14 13 2 7 15 13 4 16 10 9 9 1 14 13 4 2
22 12 9 15 14 13 4 4 4 16 9 9 1 9 1 9 1 0 9 14 13 13 2
16 11 11 1 0 9 9 7 9 1 9 1 9 13 4 4 2
17 15 1 15 1 0 9 1 9 1 12 9 1 9 13 4 4 2
21 15 9 7 9 1 9 1 3 12 9 7 12 9 1 9 0 13 4 4 4 2
21 9 9 3 9 9 1 9 1 9 13 4 4 16 9 1 10 9 14 13 4 2
15 11 1 11 11 1 15 1 1 11 1 9 14 13 4 2
43 16 0 9 1 13 1 9 1 9 3 10 9 1 14 13 4 2 7 0 9 9 3 9 0 13 4 4 7 15 13 4 16 9 14 13 1 15 0 9 13 4 4 2
24 11 1 11 11 11 11 1 12 0 11 11 1 11 1 9 1 0 11 1 1 1 9 13 2
14 15 1 12 10 9 1 14 9 7 9 1 9 13 2
12 0 12 9 1 15 9 1 0 0 11 13 2
22 11 11 11 1 9 13 1 12 9 1 9 12 9 11 1 9 9 1 9 13 4 2
47 15 1 11 11 11 11 2 11 2 1 9 11 11 11 2 11 11 2 11 2 1 9 11 11 11 2 9 9 11 11 11 11 2 9 9 11 11 11 1 14 9 9 1 9 13 4 2
9 10 15 1 9 9 13 4 4 2
22 0 12 9 1 14 12 0 9 1 14 11 1 9 1 9 13 1 9 0 13 4 2
14 15 1 10 9 11 11 11 7 11 11 1 0 13 2
18 3 14 11 1 9 9 1 9 13 2 15 9 1 9 9 13 4 2
7 15 9 1 9 13 4 2
16 9 13 1 3 0 11 1 15 12 0 9 11 1 9 13 2
11 9 1 10 0 9 1 9 13 9 13 2
11 10 9 1 11 1 9 11 14 0 13 2
17 15 12 9 7 12 9 1 14 10 9 9 9 1 9 0 13 2
11 11 1 1 9 1 9 13 0 14 13 2
24 15 0 9 13 15 11 1 12 9 9 1 12 9 1 9 9 9 1 0 14 13 4 4 2
12 10 9 13 2 11 11 11 7 11 11 11 2
33 9 1 9 15 13 15 11 1 9 10 0 9 13 4 16 11 1 12 0 9 11 11 11 7 11 11 11 1 9 14 13 4 2
19 11 1 12 0 9 1 13 16 11 1 1 9 1 9 13 0 14 13 2
36 11 1 9 1 14 9 1 2 9 2 7 2 9 2 1 9 1 9 14 13 4 2 16 15 9 9 1 9 1 15 0 9 13 4 4 2
14 11 11 10 9 1 2 9 2 1 9 13 4 4 2
52 0 9 2 11 11 11 2 1 0 12 9 1 13 4 4 16 9 9 1 1 9 11 1 11 1 1 1 9 1 0 13 4 9 1 0 7 0 9 1 1 9 1 9 1 9 13 1 9 13 4 4 2
31 15 1 10 9 1 13 1 12 1 12 9 1 1 9 1 9 7 9 1 9 13 1 1 0 13 1 9 13 4 4 2
37 2 9 2 9 1 1 0 9 1 9 7 9 1 9 13 4 4 16 15 9 2 0 9 7 9 1 1 1 9 13 1 15 9 1 14 13 2
28 11 1 0 9 11 2 11 1 9 13 4 9 1 13 16 14 12 12 9 9 9 1 9 9 13 4 4 2
18 7 12 12 9 9 14 1 13 12 12 9 1 9 0 13 4 4 2
11 10 9 1 10 9 12 12 9 13 4 2
32 11 11 1 1 11 11 11 9 11 1 11 1 1 0 9 1 9 1 14 9 2 9 7 9 1 1 10 14 9 13 4 2
30 11 1 12 9 1 11 1 9 13 13 16 11 11 1 11 11 2 11 1 1 9 0 13 1 9 0 7 0 13 2
6 15 3 0 13 4 2
41 11 1 11 1 13 9 11 11 1 9 1 13 4 16 10 9 1 12 12 9 1 1 1 0 9 1 9 9 0 13 1 1 9 1 15 9 14 13 4 4 2
33 15 13 16 11 11 1 11 11 2 11 1 9 1 13 4 11 11 11 1 12 12 9 1 10 1 9 1 1 11 13 0 13 2
29 9 1 11 1 0 11 11 11 1 0 9 1 15 11 1 9 2 9 7 9 1 9 1 13 1 1 9 13 2
12 0 9 1 9 1 10 9 1 9 13 4 2
20 11 11 11 11 1 1 1 9 9 11 11 1 9 11 11 1 9 13 4 2
32 11 11 11 11 2 11 11 11 2 11 11 11 1 9 11 11 2 15 9 11 7 9 11 11 1 14 9 1 9 0 13 2
31 11 11 11 11 2 11 11 11 11 11 2 11 11 11 11 11 7 9 9 1 9 11 11 11 14 10 9 1 0 13 2
16 0 11 9 1 9 13 11 1 11 11 11 9 9 1 13 2
17 15 1 9 11 11 2 11 11 2 11 11 7 10 0 9 13 2
33 11 1 9 12 9 9 1 9 1 13 1 3 14 12 10 0 9 1 9 13 4 15 0 9 1 9 1 9 1 1 9 13 2
21 9 7 0 9 1 13 9 11 1 9 13 1 3 9 9 13 1 0 13 4 2
15 15 2 15 1 9 13 1 1 9 1 9 3 13 4 2
10 0 9 11 1 9 1 3 9 13 2
12 10 9 1 15 0 9 1 9 1 9 13 2
15 11 1 13 11 1 9 1 9 13 0 9 1 9 13 2
23 11 1 9 11 1 14 12 9 12 9 9 7 9 13 4 15 9 1 9 1 9 13 2
10 11 1 9 1 14 9 1 9 13 2
18 0 9 1 9 13 1 1 11 1 9 1 9 9 1 9 13 4 2
10 10 9 1 9 1 0 9 14 13 2
9 11 1 9 1 9 1 9 13 2
29 11 11 1 1 12 9 1 13 9 1 9 7 9 1 9 13 1 1 0 9 1 0 9 1 0 9 13 4 2
23 9 1 11 1 9 9 9 1 11 1 10 9 13 4 9 11 1 1 1 0 13 4 2
29 11 1 15 3 0 7 9 1 1 13 4 13 16 15 11 9 1 10 9 1 1 11 9 11 11 1 9 13 2
13 11 1 13 16 11 11 9 7 9 1 9 13 2
23 15 11 11 1 9 13 16 11 11 9 1 15 11 7 11 1 9 1 1 3 14 13 2
31 11 1 0 9 1 0 9 11 11 1 11 1 9 9 9 11 11 1 13 16 15 11 1 9 0 13 1 0 9 13 2
17 9 1 9 1 1 11 11 1 9 1 9 9 12 9 0 13 2
26 10 9 11 2 11 1 11 11 11 1 9 1 0 0 13 1 9 9 1 9 1 9 13 4 4 2
33 0 13 16 11 11 2 11 1 9 1 1 11 1 11 11 1 11 13 1 11 11 1 9 1 1 9 1 12 9 13 4 4 2
10 10 9 1 11 1 9 0 13 4 2
21 7 11 1 11 1 11 11 11 9 1 11 1 9 13 1 9 1 9 13 4 2
12 9 1 12 1 1 12 9 0 13 4 4 2
12 0 12 9 15 15 9 9 1 1 13 4 2
38 11 1 11 11 9 1 11 1 9 3 13 1 9 13 4 7 11 1 9 1 9 1 9 9 1 15 13 13 4 16 9 9 0 13 1 0 13 2
29 11 11 11 1 9 1 11 11 1 0 9 1 15 9 13 1 3 11 11 15 0 9 0 13 1 9 1 13 2
26 11 2 11 1 9 0 13 1 3 9 1 9 13 4 16 15 11 11 1 9 9 13 4 4 4 2
25 0 0 9 1 13 13 16 0 9 1 10 9 1 14 9 13 4 15 9 9 1 1 0 13 2
21 9 9 11 11 11 1 14 10 9 11 2 11 11 11 11 1 12 9 13 4 2
34 15 11 1 13 4 16 0 9 1 9 10 9 1 0 13 4 10 9 1 11 11 11 11 2 11 2 1 9 1 0 13 4 4 2
18 15 13 16 11 7 11 11 11 2 11 2 10 9 1 13 4 4 2
15 11 11 11 1 1 9 9 1 9 9 1 1 9 13 2
28 15 0 11 11 11 11 1 9 9 1 13 16 9 11 11 11 11 1 0 9 0 13 1 9 13 4 4 2
30 11 11 11 11 1 14 12 9 9 1 13 16 0 0 9 1 10 9 13 4 4 2 15 0 9 1 0 13 4 2
16 9 1 15 14 14 13 4 7 15 1 14 14 13 4 4 2
37 3 9 1 10 9 0 9 1 1 1 10 9 1 10 13 16 11 9 1 13 11 11 1 11 1 9 1 1 1 0 9 1 15 9 14 13 2
23 11 7 11 11 1 14 9 13 16 11 9 1 11 1 11 11 1 9 9 13 4 4 2
13 15 1 13 4 9 1 0 9 1 9 13 4 2
24 10 9 1 0 11 7 11 1 0 9 1 13 13 16 9 1 0 9 1 0 13 4 4 2
15 15 15 14 13 4 4 16 11 1 9 9 13 4 4 2
28 11 11 11 11 11 1 0 9 1 13 4 16 9 1 1 1 0 9 1 9 9 1 9 13 4 4 4 2
42 9 1 13 13 16 9 15 9 13 4 16 11 1 9 1 9 1 15 0 9 1 1 9 1 0 9 1 9 13 7 9 1 1 9 14 13 1 9 9 13 4 2
32 10 9 1 9 1 10 9 13 15 15 9 13 7 10 9 1 1 10 9 13 4 15 1 1 13 4 4 16 9 13 4 2
18 9 9 1 12 9 13 4 4 15 11 11 1 1 9 13 4 4 2
16 11 1 1 11 9 1 9 1 1 1 9 14 13 4 4 2
33 11 1 13 13 16 11 1 12 9 11 1 1 13 4 2 15 11 2 11 9 1 11 11 7 11 1 1 11 11 11 0 13 2
9 15 15 14 11 1 1 9 13 2
28 9 1 11 1 10 9 9 9 13 4 2 14 10 9 11 11 1 12 0 9 1 10 10 0 9 13 4 2
12 10 0 9 9 7 9 2 12 1 13 4 2
10 9 1 9 10 9 1 13 4 4 2
20 9 1 10 9 7 11 1 10 9 1 9 1 13 9 2 9 13 4 4 2
28 10 3 9 1 10 9 1 9 13 4 1 9 13 4 2 15 9 13 12 0 2 0 9 1 13 4 4 2
19 10 9 1 9 1 9 13 4 2 9 1 15 9 3 14 13 4 4 2
21 0 9 7 9 9 1 9 14 1 10 9 1 0 11 1 15 9 13 4 4 2
23 9 1 11 2 11 2 11 7 11 1 10 14 12 9 9 1 9 1 13 9 13 4 2
26 9 1 9 13 16 9 1 13 4 9 15 14 15 9 1 11 1 13 4 7 0 9 1 0 13 2
27 9 9 1 1 11 1 9 14 0 13 4 4 7 15 1 15 9 1 9 0 9 1 3 14 13 4 2
23 11 1 9 9 1 9 9 11 1 0 11 11 1 9 9 1 9 1 0 9 13 4 2
21 9 9 15 9 2 9 1 9 1 13 14 15 9 1 13 1 9 13 4 4 2
27 9 11 1 12 9 1 9 13 4 13 16 10 9 1 9 13 2 15 15 14 0 9 13 13 4 4 2
22 9 1 9 1 9 13 4 16 0 9 15 13 1 7 13 1 1 9 9 1 13 2
27 15 1 9 0 9 1 1 10 10 9 9 1 9 0 13 4 4 4 2 15 9 1 1 9 13 4 2
12 9 1 13 13 16 15 10 9 13 4 4 2
24 11 11 1 9 9 7 11 1 12 12 1 11 0 9 1 9 1 9 3 13 1 9 13 2
32 10 0 9 10 9 1 3 0 9 11 11 2 9 9 2 7 11 11 1 3 13 1 9 9 1 9 13 1 9 1 13 2
30 0 0 0 9 1 13 16 9 1 1 10 9 1 0 11 2 11 11 1 10 9 10 9 1 9 1 0 13 4 2
11 10 9 1 9 13 1 3 10 9 13 2
10 7 15 15 3 14 0 9 13 4 2
24 11 2 11 1 10 9 1 0 9 2 9 1 1 15 9 0 9 1 1 12 9 9 13 2
11 15 2 11 11 2 1 9 13 4 4 2
30 11 1 9 1 1 9 9 1 10 9 1 9 9 1 15 2 15 1 14 15 9 2 9 1 9 2 9 13 4 2
28 11 1 9 9 9 1 13 7 15 1 9 1 9 13 11 11 11 1 13 9 1 9 3 0 13 4 4 2
20 11 11 1 1 1 11 1 13 9 1 1 11 1 0 11 1 13 4 4 2
25 9 13 4 4 16 0 9 1 13 4 9 1 1 0 9 1 9 1 14 15 9 1 13 4 2
18 15 9 0 9 9 1 12 2 12 9 1 0 9 9 11 1 13 2
24 9 1 13 4 4 16 9 1 11 1 9 1 9 1 1 11 11 1 9 13 4 4 4 2
13 11 1 14 11 1 15 9 1 0 13 4 4 2
25 15 13 16 15 11 1 12 10 9 1 13 2 13 4 4 15 1 11 3 9 7 9 13 4 2
13 15 1 9 1 14 11 1 13 1 9 13 4 2
42 0 13 16 10 9 1 9 1 10 9 14 13 4 16 11 1 11 1 13 4 4 4 7 15 11 1 11 9 1 14 3 0 13 4 16 11 11 15 9 13 4 2
18 10 9 1 11 7 11 1 0 9 1 15 1 1 9 14 13 4 2
19 11 7 11 1 1 0 9 1 11 1 9 1 12 0 9 0 13 4 2
11 11 11 1 15 9 12 7 12 13 4 2
10 15 9 11 1 0 9 1 1 13 2
15 9 1 15 9 1 9 2 9 1 9 1 9 14 13 2
23 15 11 1 15 9 1 13 0 9 1 1 11 11 1 12 12 9 0 13 4 4 4 2
17 9 13 4 4 4 16 9 1 9 12 12 1 9 13 4 4 2
28 11 1 11 9 0 9 9 1 11 11 1 1 9 13 1 3 11 11 1 0 9 1 12 9 0 13 4 2
12 15 1 0 12 9 1 12 9 0 13 4 2
25 15 13 16 11 1 0 13 4 9 1 9 1 9 11 11 1 12 1 1 12 1 13 4 4 2
14 0 13 16 9 9 13 9 1 9 12 13 4 4 2
17 15 9 11 1 1 11 7 11 9 1 1 9 1 1 0 13 2
18 12 9 1 11 11 1 13 9 1 9 11 11 1 12 13 4 4 2
14 11 1 0 9 9 1 11 1 1 11 11 1 13 2
13 11 11 1 9 9 1 9 1 9 13 4 4 2
9 15 1 9 1 9 13 4 4 2
23 9 1 1 9 1 1 9 0 9 0 13 4 4 15 15 0 9 14 13 4 4 4 2
30 11 1 11 1 9 9 11 11 1 15 12 9 9 1 13 16 11 9 9 9 1 1 11 1 0 9 9 13 4 2
23 15 13 16 11 11 1 9 13 13 4 2 16 15 13 13 16 11 1 15 9 13 4 2
29 11 1 13 16 11 11 1 0 9 13 7 15 9 9 1 9 1 13 11 2 11 1 9 1 9 1 9 13 2
30 9 9 1 15 13 4 1 16 15 10 9 1 11 11 2 11 1 9 2 9 13 2 15 15 13 1 9 13 4 2
19 10 9 1 15 13 16 11 2 11 1 10 9 9 1 1 0 14 13 2
47 16 15 13 16 11 9 14 1 9 1 13 0 15 9 1 9 13 2 15 11 1 15 14 10 9 13 1 9 13 4 15 9 1 15 0 9 1 1 1 14 13 1 9 13 4 4 2
18 15 13 16 15 15 9 1 1 0 0 9 1 9 13 4 4 4 2
39 15 1 2 11 11 11 11 11 1 0 9 15 11 9 1 1 10 9 0 11 11 11 11 1 1 13 4 7 15 1 9 1 9 0 13 1 13 4 2
18 9 9 1 13 9 9 1 13 4 9 1 9 13 12 13 4 4 2
35 15 13 16 15 11 1 11 1 9 11 11 1 1 3 9 1 13 7 9 1 3 11 13 1 1 15 0 9 13 1 9 13 4 4 2
19 16 2 9 1 9 13 4 16 9 1 11 9 1 11 13 4 4 4 2
28 11 1 13 16 11 1 9 1 10 9 1 0 13 4 4 1 3 9 1 0 9 7 9 1 13 4 4 2
20 9 1 9 1 9 13 1 1 15 13 16 15 1 1 3 1 9 13 4 2
10 3 9 1 11 13 14 0 9 13 2
15 10 9 1 12 9 1 0 13 1 14 9 13 4 4 2
20 11 1 11 11 11 11 11 11 1 1 2 9 1 12 9 1 9 0 13 2
15 9 1 0 9 1 9 1 13 15 9 13 4 4 4 2
30 11 1 0 9 1 9 11 11 11 11 11 2 11 1 13 4 16 10 0 9 3 13 4 15 1 14 9 13 4 2
17 9 1 9 11 11 1 13 16 9 1 9 1 10 9 0 13 2
19 11 11 11 11 11 11 1 9 1 12 0 9 1 9 13 1 13 4 2
11 10 9 1 9 1 9 13 4 4 4 2
29 11 11 11 1 11 11 11 11 11 2 11 2 1 13 15 9 0 9 1 9 1 0 13 1 0 13 4 4 2
15 0 9 1 9 7 0 9 9 1 14 0 9 13 4 2
19 11 11 11 7 11 11 1 14 12 9 13 9 1 1 10 9 13 4 2
27 11 9 1 9 1 13 16 9 11 1 9 1 1 13 9 13 1 9 1 12 0 9 9 13 13 4 2
19 12 9 1 9 11 11 11 11 1 11 1 1 11 1 9 13 4 4 2
25 9 1 10 9 1 13 1 9 9 1 0 9 1 15 14 9 9 13 1 9 13 1 3 13 2
45 11 7 11 11 1 9 1 1 9 1 9 1 13 16 11 11 11 1 13 4 16 15 11 1 11 11 11 11 11 2 11 2 1 1 12 0 0 9 13 1 3 14 9 13 2
14 10 0 9 0 9 7 11 1 9 1 0 9 13 2
20 15 13 16 11 1 0 9 1 9 13 1 1 11 10 9 11 1 9 13 2
22 15 1 11 1 9 9 1 11 11 11 11 1 10 9 1 9 0 13 1 13 4 2
15 10 9 9 1 11 1 9 11 1 9 13 1 9 13 2
29 16 9 9 1 0 9 1 13 1 9 13 4 11 11 1 10 9 1 15 14 9 1 9 13 1 9 13 4 2
26 11 1 9 13 1 11 11 1 9 9 1 9 11 11 11 1 13 16 9 1 0 13 4 4 4 2
32 7 15 10 9 1 1 10 0 9 1 15 0 9 1 0 13 1 0 13 15 11 1 9 1 9 7 9 1 9 13 4 2
13 15 13 16 9 1 9 11 1 9 1 0 13 2
33 11 2 11 11 11 1 9 0 13 1 1 11 1 11 11 11 11 15 9 1 1 11 1 9 9 1 9 1 9 13 4 4 2
12 15 3 9 11 11 11 1 12 9 1 13 2
18 11 1 1 1 14 9 1 1 9 1 10 9 13 4 1 9 13 2
33 11 2 11 1 1 0 9 11 11 1 13 11 11 1 10 9 14 0 13 16 11 11 1 12 9 9 1 1 11 1 9 13 2
11 7 15 9 15 1 11 1 14 13 4 2
15 9 15 1 9 13 4 4 16 9 15 9 1 14 13 2
31 11 1 9 1 0 9 1 1 11 1 1 11 0 13 4 3 0 13 4 4 7 9 1 0 11 1 9 3 10 13 2
22 9 1 9 9 1 9 1 0 9 14 13 1 0 9 11 1 9 14 13 14 13 2
22 9 9 2 9 7 15 0 0 9 1 0 9 1 1 11 11 11 11 13 4 4 2
7 7 11 15 0 14 13 2
29 11 16 11 1 11 1 9 1 9 13 4 16 15 15 0 9 1 9 13 4 15 15 10 9 1 9 13 4 2
27 0 9 15 13 16 11 11 11 11 11 11 7 11 2 11 11 11 1 11 1 14 0 13 1 9 13 2
9 10 9 9 9 1 13 4 4 2
38 11 9 11 11 7 11 1 11 11 1 1 9 13 1 9 1 11 11 1 13 9 9 1 1 11 11 1 1 9 9 1 9 1 9 13 4 4 2
30 3 14 2 9 1 1 0 7 0 9 9 1 0 2 0 13 1 3 11 1 9 1 10 0 9 1 0 13 4 2
30 12 9 1 1 0 9 9 13 7 0 12 9 1 1 15 9 14 13 4 16 15 0 13 1 9 1 13 4 4 2
42 9 9 1 9 1 1 11 15 9 13 4 4 16 0 0 9 1 1 10 9 1 9 1 1 15 9 9 1 0 2 0 13 1 9 1 0 9 14 13 4 4 2
41 10 9 1 11 1 1 14 15 0 13 4 4 4 16 9 7 9 9 1 9 0 13 1 1 15 9 9 1 9 1 0 9 13 7 15 1 9 9 0 13 2
40 11 11 11 2 11 2 1 0 9 7 9 1 9 11 11 7 15 9 1 1 9 1 0 2 0 9 1 9 1 9 9 11 11 1 9 1 9 13 4 2
19 15 13 4 16 11 1 10 9 9 1 2 0 2 0 9 1 13 4 2
20 11 1 9 13 4 16 9 1 9 1 13 1 1 9 15 14 13 4 4 2
36 11 1 11 11 1 9 1 12 9 1 15 13 16 11 1 0 9 9 1 10 9 10 9 1 13 4 16 9 1 9 1 9 10 0 13 2
18 15 13 16 11 1 13 4 9 1 1 11 1 0 9 1 13 4 2
15 15 13 16 9 1 13 1 1 9 9 14 13 4 4 2
30 9 9 1 0 9 11 11 11 1 13 16 11 11 11 11 13 4 4 16 15 11 1 9 1 9 14 13 13 4 2
19 7 15 1 9 1 9 9 1 0 0 11 11 1 9 1 0 13 4 2
35 11 11 11 11 11 1 9 11 1 13 16 16 11 11 1 1 1 15 9 14 13 4 2 3 15 11 11 1 0 9 1 13 4 4 2
51 3 11 1 11 11 11 7 11 11 11 1 9 11 11 11 7 11 11 1 11 1 12 0 9 1 13 16 0 0 9 1 13 1 1 11 11 2 11 2 1 9 11 11 1 0 9 1 1 0 13 2
17 15 11 9 1 1 9 1 13 1 14 0 9 0 14 13 4 2
12 9 14 1 14 12 11 9 11 1 0 13 2
25 9 1 9 9 1 1 11 9 1 9 13 4 1 9 1 11 7 11 1 9 1 1 9 13 2
23 11 11 1 12 9 1 14 9 1 9 1 12 9 1 13 12 9 13 1 9 13 4 2
28 9 1 11 11 1 9 11 11 11 1 13 16 9 1 9 1 9 7 9 1 1 15 9 14 13 4 4 2
18 11 1 11 2 11 2 7 11 1 0 9 1 9 1 15 9 13 2
19 7 2 11 2 11 11 2 11 7 0 9 1 11 1 9 1 9 13 2
24 9 9 1 0 3 9 9 1 9 1 1 13 4 11 11 11 11 11 1 9 0 13 4 2
26 16 2 0 9 1 9 11 11 11 1 9 13 4 12 9 1 9 1 9 13 13 1 9 13 4 2
13 2 0 9 2 1 9 0 9 1 13 4 4 2
10 9 1 14 10 9 9 13 4 4 2
10 15 1 9 13 1 10 15 13 4 2
9 15 9 0 2 8 9 1 13 2
21 0 9 1 12 9 10 9 9 1 1 0 9 1 9 9 1 9 13 4 4 2
10 15 9 13 1 15 2 8 9 13 2
7 9 0 9 13 4 4 2
17 10 9 9 1 12 9 1 12 12 1 9 1 9 13 4 4 2
12 9 2 9 1 9 1 0 0 9 0 13 2
7 15 9 0 9 1 13 2
11 9 13 14 14 15 1 9 14 13 4 2
17 9 9 1 9 13 1 9 1 9 7 9 1 14 0 9 13 2
9 9 1 14 15 13 4 4 4 2
11 10 9 10 9 9 1 9 1 13 4 2
13 9 1 15 9 2 9 7 9 9 12 13 4 2
13 11 1 12 0 9 0 12 9 1 9 1 13 2
14 15 1 9 1 11 1 12 9 1 9 13 4 4 2
7 15 9 1 0 9 13 2
6 10 9 1 9 13 2
6 15 14 12 9 13 2
9 10 9 12 9 15 1 13 4 2
8 9 1 1 15 9 14 13 2
12 12 9 13 0 9 1 9 9 13 4 4 2
7 9 9 1 9 13 4 2
10 15 1 15 0 9 1 13 4 4 2
18 15 11 9 1 11 9 1 12 9 1 12 12 1 9 13 4 4 2
13 12 9 1 15 12 12 1 9 1 9 13 4 2
19 10 9 11 2 11 2 11 2 11 2 11 14 9 1 0 9 0 13 2
7 12 9 9 13 13 4 2
6 10 3 9 13 4 2
14 15 1 9 9 9 1 14 12 9 9 9 13 4 2
11 3 15 12 9 1 1 0 9 13 4 2
10 15 15 15 9 1 14 13 4 4 2
15 12 0 9 15 0 9 1 13 10 9 1 0 13 4 2
8 15 9 1 12 9 14 13 2
13 0 9 1 13 1 1 15 10 9 1 13 4 2
17 9 1 1 12 9 15 15 9 1 13 0 9 1 13 4 4 2
10 10 3 15 9 1 9 13 4 4 2
21 9 0 13 1 3 9 9 1 9 1 9 13 4 15 9 15 13 0 13 4 2
24 15 1 14 10 9 1 9 9 13 4 4 2 15 9 2 8 14 9 1 0 13 4 4 2
11 9 1 9 1 14 10 9 13 4 4 2
16 10 0 9 15 13 2 15 10 9 13 9 1 9 13 4 2
28 3 2 8 0 9 15 0 9 13 9 13 4 4 2 16 15 9 1 9 1 9 2 9 13 13 4 4 2
9 9 13 1 9 14 15 13 4 2
7 10 9 14 15 0 13 2
13 0 9 1 9 13 16 10 9 15 9 13 4 2
17 10 9 1 9 10 3 1 13 16 9 9 13 1 14 13 4 2
12 3 0 9 1 10 9 3 15 9 13 4 2
6 9 1 14 13 4 2
26 0 9 15 13 16 9 1 0 9 9 1 9 13 1 1 15 9 1 1 9 13 13 14 4 4 2
20 9 1 12 9 7 12 0 9 1 1 9 1 9 11 1 13 4 4 4 2
17 10 9 1 9 1 14 12 9 9 1 9 13 4 1 9 13 2
17 12 9 1 13 0 9 1 1 15 3 0 9 13 4 4 4 2
24 9 1 11 2 11 11 2 11 2 11 7 9 9 9 11 1 15 9 1 9 13 4 4 2
10 10 9 11 11 1 0 13 4 4 2
11 9 1 9 1 9 11 11 1 13 4 2
30 16 10 9 1 11 11 11 1 9 1 15 0 9 14 13 4 4 4 2 7 11 1 0 9 1 13 4 4 4 2
18 3 11 1 10 12 9 7 12 11 1 12 0 9 13 4 4 4 2
18 0 9 11 7 9 9 1 1 10 9 1 9 14 3 13 4 4 2
24 0 13 16 11 11 1 1 1 11 7 9 9 1 0 0 9 13 11 1 15 9 13 4 2
15 3 11 1 11 11 11 0 9 1 1 1 13 4 4 2
25 9 9 1 11 11 1 15 9 14 13 4 4 2 7 9 1 9 11 1 14 13 4 4 4 2
15 9 9 1 12 9 7 9 11 11 11 1 10 9 13 2
26 3 0 9 11 11 11 1 14 10 9 1 9 13 4 13 16 10 9 0 9 1 1 0 14 13 2
29 11 1 9 1 9 1 0 13 4 11 11 9 11 11 1 11 1 13 16 11 11 13 16 9 1 13 4 4 2
24 15 1 14 15 13 16 0 9 9 1 9 1 11 11 11 1 9 1 0 14 13 4 4 2
35 9 1 9 1 11 1 13 16 16 15 13 4 16 9 1 13 4 9 1 9 1 14 13 2 16 15 0 9 1 9 1 9 13 4 2
23 15 13 16 11 11 15 14 11 1 15 14 9 13 4 4 7 15 15 14 0 14 13 2
54 9 1 13 1 11 11 1 0 9 1 1 1 13 4 1 11 1 13 16 15 15 1 1 15 9 14 13 2 7 0 9 1 15 13 13 16 16 9 13 16 15 11 1 13 4 4 7 15 15 14 0 14 13 2
22 15 11 1 10 9 1 0 13 4 16 11 11 9 9 1 9 1 9 13 4 4 2
25 15 1 14 15 13 16 10 9 14 0 14 13 2 16 0 9 1 9 9 1 11 14 13 4 2
25 16 2 15 13 4 16 11 11 1 11 9 1 0 15 14 11 1 9 1 1 9 14 13 4 2
32 11 1 13 16 11 11 11 11 11 1 15 11 1 9 1 1 1 9 13 4 4 2 7 15 0 9 1 9 14 13 4 2
28 3 9 1 9 1 13 9 1 0 13 1 1 9 1 10 9 1 8 13 4 15 9 9 9 1 13 4 2
26 10 9 13 16 11 9 11 11 3 2 8 9 13 4 7 11 11 11 1 9 9 1 9 14 13 2
14 11 11 11 11 1 10 9 1 9 0 13 4 4 2
12 9 9 9 9 9 9 1 13 4 4 4 2
12 9 1 9 1 9 1 1 12 9 13 4 2
15 9 11 10 9 1 15 1 9 1 0 0 13 4 4 2
10 9 13 7 9 1 13 4 9 8 2
17 9 1 9 1 1 11 1 15 13 9 13 15 15 0 13 4 2
12 9 9 1 1 13 9 9 1 9 14 13 2
12 11 11 11 1 14 9 13 7 9 14 13 2
12 9 9 9 11 11 11 1 9 14 0 13 2
13 3 1 12 9 1 9 1 9 1 13 3 13 2
31 11 11 11 11 1 11 1 9 1 13 10 9 1 9 1 13 4 11 11 11 1 9 11 11 11 1 9 1 9 13 2
16 9 11 1 9 0 13 9 9 9 9 9 1 13 4 4 2
13 9 1 0 9 1 14 9 1 9 13 4 4 2
23 16 9 1 15 0 9 14 13 4 15 15 9 7 9 1 9 1 9 14 13 4 4 2
19 0 9 1 9 14 13 4 15 9 8 13 4 1 9 0 13 4 4 2
39 11 11 11 11 1 0 0 9 1 1 11 11 1 11 1 9 1 9 1 1 9 1 9 1 9 9 11 11 11 1 9 1 10 9 1 9 13 4 2
16 3 9 1 9 13 1 9 13 4 15 9 11 1 14 13 2
14 9 1 9 13 4 15 9 1 9 1 9 0 13 2
7 3 9 1 9 13 4 2
6 15 12 9 14 13 2
9 11 1 9 0 9 1 13 4 2
12 11 1 9 12 12 9 11 1 9 13 4 2
11 3 1 11 1 15 1 3 14 13 4 2
11 3 1 9 1 15 9 9 1 14 13 2
17 9 9 9 11 11 11 14 9 9 1 1 9 1 1 13 4 2
15 9 1 13 9 1 11 1 9 1 9 1 9 13 4 2
12 15 9 1 1 9 1 0 13 4 4 4 2
13 9 1 0 9 1 11 1 10 9 0 13 4 2
13 9 0 13 4 15 9 1 14 15 9 14 13 2
17 9 9 1 0 9 1 14 11 1 9 1 13 1 9 14 13 2
11 11 1 9 1 9 14 11 1 14 13 2
11 0 9 13 1 1 11 1 15 9 13 2
31 15 1 11 1 9 1 9 1 13 1 14 9 13 4 7 3 1 11 11 11 1 9 1 9 1 1 9 1 9 13 2
15 9 1 9 1 11 1 9 1 13 13 1 9 9 13 2
25 9 1 11 1 9 13 4 4 7 10 9 1 9 1 13 9 9 1 1 1 3 13 4 4 2
34 11 1 9 13 4 9 9 1 1 9 9 11 11 1 11 1 13 16 15 11 9 1 11 1 11 11 11 7 0 9 1 9 13 2
18 11 9 1 10 0 0 9 1 0 9 9 9 1 1 9 13 4 2
18 9 1 13 4 12 0 9 1 9 11 1 9 9 11 11 11 13 2
17 9 1 1 9 11 11 1 9 13 7 15 11 9 1 9 13 2
36 9 1 0 0 11 9 11 11 11 1 13 16 9 1 9 1 1 1 0 9 1 15 14 13 4 4 7 15 11 9 1 9 13 4 4 2
13 11 9 1 14 12 9 11 1 13 1 9 13 2
12 11 1 13 16 11 9 1 11 11 0 13 2
15 10 9 9 1 3 10 0 11 11 11 1 14 9 13 2
17 15 13 16 15 11 9 1 1 1 11 1 9 1 14 9 13 2
44 11 1 0 9 1 9 1 9 1 1 1 13 4 1 15 13 16 11 15 14 9 9 1 1 0 13 16 9 9 7 9 1 9 1 9 1 15 3 10 14 13 4 4 2
25 3 11 11 11 1 9 13 4 16 11 7 11 1 1 1 0 9 9 0 9 1 14 0 13 2
24 9 1 11 1 1 11 1 11 11 11 7 11 11 11 11 11 1 14 9 13 1 9 13 2
18 15 1 11 11 1 11 11 1 12 0 9 1 11 1 9 13 4 2
26 0 9 1 15 14 0 13 16 9 11 12 9 9 1 13 7 9 1 0 9 1 1 9 9 13 2
22 0 9 1 0 9 2 9 7 9 9 1 0 9 1 11 1 15 9 1 9 13 2
22 10 3 11 1 0 2 0 9 1 12 9 1 9 13 4 7 12 9 0 13 4 2
26 9 11 1 11 9 1 9 9 9 1 9 1 13 13 9 1 12 0 11 11 1 9 13 4 4 2
11 10 9 1 12 9 1 0 13 4 4 2
28 11 2 11 7 11 1 9 1 9 9 1 10 2 10 9 13 2 7 9 1 9 1 15 9 14 13 4 2
56 15 9 1 0 9 0 9 1 13 4 4 2 9 9 1 9 1 9 9 13 4 4 2 9 1 9 0 2 0 9 1 13 4 4 7 9 1 9 1 9 1 9 13 4 15 15 1 0 9 1 9 10 0 14 13 2
15 9 1 12 9 1 12 1 13 14 9 1 0 9 13 2
6 9 9 1 13 4 2
13 9 2 9 1 9 1 13 9 1 10 9 13 2
17 15 13 16 12 9 1 11 1 9 1 9 13 15 9 13 4 2
22 11 7 11 1 12 0 9 1 1 11 1 15 9 9 1 9 1 9 2 9 13 2
21 9 1 9 1 1 12 9 1 15 2 15 1 9 9 1 9 13 1 9 13 2
25 9 1 1 12 9 10 9 11 1 0 9 1 15 2 15 1 9 9 1 9 2 9 13 4 2
42 9 9 1 0 9 1 1 11 7 11 1 1 11 11 2 11 1 13 9 1 11 11 1 1 12 9 1 9 1 15 15 1 9 9 1 9 1 9 2 9 13 2
34 11 1 11 11 1 11 11 1 9 11 11 11 1 11 1 9 9 7 9 1 9 11 1 0 9 1 0 0 9 11 11 1 13 2
22 11 11 1 11 1 1 1 11 11 1 0 9 1 0 9 11 11 1 9 13 4 2
16 9 1 15 14 13 4 4 16 9 1 15 9 1 9 13 2
23 3 9 1 9 9 9 9 1 0 13 4 4 7 15 0 9 1 0 9 13 4 4 2
24 0 9 1 11 7 11 1 3 11 7 11 1 9 9 13 1 0 9 1 9 13 4 4 2
36 0 9 11 1 11 1 11 11 11 1 11 9 1 1 0 0 9 1 12 9 1 0 9 1 9 1 9 9 13 1 9 1 9 13 4 2
57 11 7 11 1 9 9 13 1 9 1 9 15 13 16 11 15 1 15 0 9 1 0 13 1 0 14 13 4 2 7 11 1 15 9 1 9 9 0 13 4 4 7 9 9 13 1 1 15 11 11 1 9 13 1 9 13 2
9 9 1 9 1 9 13 1 13 2
20 9 1 9 12 9 9 11 11 11 1 12 9 1 9 11 1 13 4 4 2
19 7 9 1 9 12 9 9 11 11 11 0 9 9 1 9 13 4 4 2
13 11 11 11 11 14 15 9 1 9 1 9 13 2
15 9 1 0 9 1 1 11 11 1 9 13 4 4 4 2
16 9 13 7 0 9 9 1 1 10 9 1 9 13 4 4 2
26 11 1 11 1 1 1 12 0 9 9 1 11 1 9 7 0 9 13 1 9 1 0 13 4 4 2
15 11 1 11 1 9 1 13 4 9 0 13 1 13 4 2
10 11 11 1 15 9 11 1 13 4 2
35 11 1 13 16 11 11 1 10 9 1 9 13 1 9 13 4 4 7 9 11 7 11 11 11 11 1 13 4 9 0 13 1 13 4 2
18 11 7 11 11 11 11 11 11 11 2 11 2 1 0 9 9 13 2
20 15 13 16 11 1 0 10 9 1 10 9 1 10 9 11 1 1 13 4 2
16 11 1 13 4 4 4 16 15 15 10 9 1 0 14 13 2
35 11 11 11 1 9 1 1 0 13 4 12 9 7 9 1 9 1 0 12 0 9 10 9 1 0 13 4 4 2 15 9 13 0 13 2
25 15 1 11 11 11 1 11 1 9 9 9 1 1 0 9 7 9 13 1 1 9 1 9 13 2
31 11 1 13 4 11 1 13 16 15 15 13 9 13 16 11 11 11 1 15 15 9 0 13 4 9 1 9 1 13 4 2
12 11 11 1 13 11 11 1 15 9 0 13 2
14 15 1 9 1 11 7 15 0 9 11 13 4 4 2
19 9 9 11 11 11 1 13 16 11 1 11 7 15 9 9 11 13 4 2
9 9 1 9 9 1 9 13 4 2
18 11 11 1 13 9 1 9 15 13 15 11 1 0 13 1 9 13 2
8 10 10 9 1 9 9 13 2
8 9 9 1 9 1 9 13 2
19 0 13 16 11 1 0 11 1 11 2 11 2 11 1 11 1 9 13 2
10 9 1 12 9 1 9 1 9 13 2
18 9 1 1 11 1 11 11 11 9 9 7 11 11 11 1 9 13 2
15 11 1 11 11 9 1 9 1 9 3 0 13 4 4 2
28 0 9 1 9 1 0 9 1 12 9 1 9 13 4 7 12 1 10 9 1 9 1 9 13 4 4 4 2
23 10 9 1 11 1 9 1 11 7 11 9 1 1 0 0 9 1 9 0 13 4 4 2
31 0 13 16 11 1 10 9 1 13 9 1 12 1 10 9 1 9 13 4 4 7 12 12 1 10 9 0 13 4 4 2
13 15 14 15 1 10 9 9 1 9 13 4 4 2
13 12 9 1 1 9 1 12 9 13 4 4 4 2
27 12 0 9 9 1 13 16 9 9 11 1 1 0 12 9 1 11 9 1 12 9 1 9 0 13 4 2
9 15 1 12 9 0 13 4 4 2
49 11 1 3 0 9 1 9 11 11 1 9 0 13 2 3 15 11 11 11 1 14 12 9 1 15 9 11 11 1 9 1 9 1 13 1 9 1 13 11 1 11 11 11 1 1 0 9 13 2
11 0 11 1 12 9 1 15 9 14 13 2
18 9 9 14 11 11 13 4 7 0 9 1 11 1 9 1 9 13 2
26 9 1 2 11 9 15 9 1 13 2 7 2 11 1 9 1 9 0 14 13 2 1 9 13 4 2
14 15 1 11 1 9 1 12 9 14 11 1 13 4 2
21 15 11 1 9 1 11 11 14 11 1 0 13 1 9 0 13 1 9 13 4 2
38 11 11 1 14 11 1 9 1 9 1 9 13 4 7 11 1 9 1 9 9 11 11 11 1 11 1 0 13 11 11 1 0 13 1 9 13 4 2
16 0 13 16 9 11 11 1 9 11 11 11 11 1 9 13 2
22 15 9 11 11 1 11 1 10 9 13 2 15 15 9 9 1 13 9 13 4 4 2
11 11 1 11 1 11 11 11 11 9 13 2
11 9 1 1 9 1 0 9 13 4 4 2
19 0 7 0 9 1 10 0 9 9 1 9 13 1 1 11 13 4 4 2
10 15 12 11 11 9 9 14 0 13 2
24 11 11 11 11 11 11 7 11 11 11 1 10 0 2 0 9 12 0 9 9 1 9 13 2
17 11 1 11 11 11 11 11 11 1 9 1 15 9 13 4 4 2
15 10 9 0 0 9 1 9 9 1 9 0 13 4 4 2
7 11 11 1 15 9 13 2
18 0 2 0 9 7 11 11 9 11 11 9 1 9 9 1 0 13 2
18 9 1 1 12 11 11 11 9 7 12 11 11 9 9 1 9 13 2
14 15 1 12 9 1 12 0 2 0 9 15 9 13 2
17 9 1 0 9 1 13 14 12 12 9 1 9 13 1 9 13 2
15 9 1 1 15 9 13 1 9 11 1 1 0 14 13 2
26 12 9 3 9 7 9 1 0 13 11 1 12 9 1 15 0 9 1 14 12 9 1 1 13 4 2
10 0 9 1 1 10 9 0 13 4 2
11 9 1 13 1 9 1 15 9 14 13 2
34 9 1 9 1 12 9 1 11 9 1 11 11 1 9 2 9 1 13 1 11 11 0 9 1 9 1 0 13 15 9 1 13 4 2
17 15 15 9 1 13 4 4 15 15 9 1 15 9 13 4 4 2
10 15 1 9 1 9 15 1 13 4 2
20 9 9 1 1 1 9 13 1 11 3 2 3 9 1 9 13 14 13 4 2
22 12 9 1 9 13 1 0 10 9 1 0 9 11 1 15 0 9 1 9 13 4 2
17 15 15 9 12 0 9 1 9 11 11 1 12 9 1 13 4 2
24 0 13 16 11 1 0 9 1 12 12 9 1 12 9 1 9 11 1 9 0 13 4 4 2
18 9 9 1 12 0 9 1 1 10 9 1 9 9 13 4 4 4 2
12 16 15 10 9 1 9 13 1 9 13 4 2
13 9 1 1 0 11 11 1 9 0 13 4 4 2
14 16 15 14 15 9 1 1 0 9 13 4 4 4 2
16 11 11 1 9 1 1 15 9 1 9 13 1 9 14 13 2
6 15 15 10 9 13 2
14 9 1 12 9 1 14 0 9 9 1 9 1 13 2
13 3 15 9 9 9 2 9 2 1 13 4 4 2
21 9 1 13 13 16 15 9 1 0 9 1 13 1 1 1 3 14 9 13 4 2
11 0 13 16 11 11 0 9 1 0 13 2
11 10 9 1 0 9 1 9 13 4 4 2
19 9 1 1 11 15 9 1 2 9 1 9 7 9 1 9 13 4 4 2
18 9 1 13 16 10 9 1 9 9 0 13 7 15 9 13 4 4 2
24 9 15 1 9 13 1 13 0 14 13 4 15 1 15 9 1 9 13 1 9 14 13 4 2
36 16 15 12 2 12 9 1 9 1 9 13 1 9 13 4 4 7 0 9 0 13 1 3 15 0 9 7 9 1 9 1 14 9 13 4 2
14 15 15 9 1 1 0 9 7 9 13 4 4 4 2
24 9 9 1 13 13 16 9 1 0 9 1 9 1 1 1 9 13 1 1 9 13 4 4 2
20 9 1 9 1 9 7 15 0 9 1 1 15 9 1 13 1 9 14 13 2
10 15 1 14 15 9 1 13 4 4 2
28 15 0 9 1 9 1 10 13 1 1 9 1 11 1 11 9 1 12 10 9 9 9 13 1 9 13 4 2
16 15 1 0 9 7 0 9 1 9 1 9 14 13 4 4 2
34 11 9 11 11 1 11 11 1 0 9 1 12 9 9 1 10 9 13 4 13 16 12 0 9 7 9 1 1 9 13 4 4 4 2
17 0 9 1 12 10 0 9 1 1 9 1 0 9 13 4 4 2
12 15 9 13 4 1 9 1 9 14 0 13 2
32 15 13 16 9 1 0 9 1 9 1 9 1 1 13 4 1 2 11 11 11 11 2 2 11 2 1 9 13 4 4 4 2
11 15 13 16 9 12 11 13 13 4 4 2
26 10 9 1 11 1 9 13 4 4 7 9 13 16 0 12 9 1 1 15 9 1 0 13 4 4 2
21 15 13 16 0 9 1 9 9 2 11 11 2 1 11 9 1 13 1 0 13 2
16 16 11 15 1 0 13 4 16 15 0 9 14 13 4 4 2
26 15 15 14 13 16 9 1 3 14 15 9 2 9 9 0 13 15 15 9 1 1 11 0 13 4 2
37 15 13 16 11 1 13 1 9 2 9 9 11 11 1 1 1 13 4 7 10 3 11 9 1 0 9 2 9 9 1 9 9 14 9 1 13 2
21 9 11 1 9 1 9 1 0 9 1 9 1 9 13 4 15 9 1 9 13 2
15 15 13 16 10 9 1 9 9 1 0 7 0 9 13 2
20 15 15 13 10 0 9 1 13 4 4 2 7 15 9 8 13 9 13 4 2
12 9 11 1 13 16 9 1 15 9 14 13 2
33 7 15 16 9 1 13 9 13 2 15 9 1 1 1 12 2 12 0 9 2 9 0 13 4 4 4 16 3 10 9 14 13 2
22 0 13 16 10 9 1 9 1 9 9 1 10 0 9 1 0 9 8 13 4 4 2
33 9 1 9 1 1 9 9 9 1 9 13 4 7 3 1 15 9 1 9 1 12 0 9 1 0 13 1 9 13 4 4 4 2
23 9 11 1 15 14 13 16 9 1 0 0 9 1 9 1 12 9 1 0 13 4 4 2
53 15 9 11 11 11 1 1 9 9 1 1 0 9 1 9 1 9 13 4 0 2 0 11 11 11 11 11 11 11 1 0 13 4 4 16 3 9 1 0 9 16 11 7 9 1 9 13 1 15 9 14 13 2
48 11 1 11 1 15 11 9 11 11 1 9 13 7 15 0 13 16 9 9 1 0 7 0 9 1 9 1 0 9 13 4 7 11 7 9 1 9 1 15 9 1 9 1 14 13 4 4 2
23 16 11 1 10 9 1 9 1 0 9 0 13 1 9 1 9 1 14 9 13 4 4 2
25 11 1 13 16 11 7 9 1 0 9 1 9 0 7 0 9 1 9 1 9 1 14 13 4 2
30 11 1 1 11 1 0 9 1 0 9 1 9 1 0 9 1 1 0 9 1 9 9 1 9 1 1 1 9 13 2
34 10 9 1 15 0 13 16 9 0 9 1 9 1 9 1 13 4 3 11 7 9 1 9 1 15 9 1 9 13 14 13 4 4 2
33 15 15 14 0 13 16 0 9 1 9 1 1 1 9 9 9 1 13 0 9 1 9 14 10 9 1 3 13 4 14 13 4 2
30 15 1 11 1 9 9 1 9 7 15 9 9 1 13 0 9 1 9 1 9 9 11 11 1 14 9 2 9 13 2
44 11 1 13 16 9 1 10 9 1 9 9 1 9 13 4 1 1 9 9 9 11 2 11 2 11 7 11 1 11 2 11 2 11 1 1 12 12 9 1 9 13 4 4 2
20 7 0 9 9 1 0 9 1 1 10 9 1 12 12 9 1 9 13 4 2
24 10 9 10 9 1 11 1 10 9 9 1 13 4 12 12 9 1 9 1 1 13 4 4 2
27 9 9 9 1 1 15 3 10 9 9 1 12 9 7 9 1 14 12 9 14 9 1 9 13 4 4 2
15 9 11 11 1 9 1 13 1 15 12 9 1 9 13 2
28 15 13 4 15 3 0 9 9 9 2 11 11 11 11 2 2 11 2 11 2 1 9 1 9 13 4 4 2
28 15 9 1 12 9 14 15 9 13 4 15 14 11 1 0 13 1 3 1 0 9 9 1 9 0 14 13 2
14 0 13 16 15 15 9 9 1 12 9 13 4 4 2
24 11 11 1 9 9 9 11 11 1 13 16 15 11 7 11 1 11 2 11 1 9 13 4 2
14 11 1 10 9 1 1 2 11 2 1 9 13 4 2
23 11 1 13 16 16 10 9 9 1 9 9 1 12 9 13 4 16 9 11 11 1 13 2
15 7 16 9 1 12 9 9 13 1 15 11 11 1 13 2
12 11 1 13 16 10 9 1 11 0 13 4 2
8 15 3 15 9 1 9 13 2
13 10 9 15 9 1 9 1 9 14 13 4 4 2
16 11 11 1 11 1 11 11 11 1 9 1 3 0 13 4 2
15 7 15 1 14 15 13 16 9 1 15 9 13 4 4 2
23 9 1 0 9 11 11 1 11 1 9 1 9 13 4 13 16 11 1 9 3 0 13 2
22 7 15 13 2 11 1 15 1 12 0 9 9 7 0 9 13 2 9 1 9 13 2
28 11 1 9 11 11 11 11 1 11 1 9 1 13 16 0 9 1 0 9 1 1 0 9 14 13 4 4 2
27 15 13 16 0 9 1 15 9 1 9 1 0 13 4 16 9 1 15 1 0 9 13 1 9 14 13 2
14 9 1 15 14 12 9 13 7 9 15 1 0 13 2
30 15 13 4 4 16 15 9 1 9 1 11 1 9 1 1 0 9 1 9 0 9 1 1 0 0 9 13 4 4 2
43 9 9 1 11 1 0 0 9 9 9 9 11 11 11 11 1 11 9 1 13 9 1 9 1 0 9 13 4 12 9 1 0 9 1 9 13 7 9 1 0 13 4 2
26 11 1 11 1 9 13 9 9 1 15 9 1 9 13 7 0 9 1 9 9 13 1 0 13 4 2
45 11 9 1 0 13 9 9 1 13 9 1 9 1 9 9 1 9 9 9 11 11 11 1 9 1 12 0 11 11 11 2 11 2 1 9 9 11 11 11 11 1 15 9 13 2
22 0 11 1 11 9 1 12 12 9 9 7 12 9 1 9 1 9 13 13 4 4 2
28 11 1 9 1 9 7 9 1 9 1 9 1 0 13 1 11 1 9 1 1 13 9 1 11 13 4 4 2
31 11 9 1 10 9 10 0 9 7 9 1 0 9 1 9 13 1 1 9 7 9 1 9 13 7 15 13 4 13 4 2
30 15 1 2 11 9 0 11 1 10 9 1 12 9 1 12 9 1 9 13 4 7 15 9 1 0 13 4 4 4 2
6 3 9 15 1 13 2
23 7 15 10 9 1 9 13 16 0 9 1 1 11 1 9 12 9 1 9 1 13 4 2
36 11 11 1 9 1 11 11 1 11 11 1 0 12 9 11 11 11 1 1 11 11 1 9 13 1 10 9 12 9 1 9 13 1 9 13 2
20 9 1 13 16 11 11 1 1 9 9 1 9 12 2 12 9 1 13 4 2
24 12 12 1 10 9 1 11 11 1 9 1 3 0 0 0 9 1 1 1 13 4 4 4 2
20 10 9 1 0 9 9 13 1 11 1 11 2 11 1 9 13 9 13 4 2
21 11 12 9 1 1 9 1 9 11 2 11 1 9 9 1 9 9 11 1 13 2
17 11 11 1 11 11 11 1 12 12 9 9 9 9 9 13 4 2
15 15 1 9 9 11 1 0 9 1 9 13 1 9 13 2
22 9 1 13 13 16 11 1 15 9 0 9 0 11 11 11 11 2 11 2 1 13 2
21 11 11 1 15 11 0 11 7 11 9 9 1 1 12 12 9 9 13 1 13 2
17 15 9 14 12 11 11 11 1 12 0 9 1 9 1 13 4 2
11 3 10 0 9 11 11 1 1 14 13 2
16 9 0 0 9 11 11 1 13 13 4 9 1 9 13 4 2
21 11 1 0 9 1 13 13 9 1 1 10 9 1 0 0 9 1 13 4 4 2
17 11 1 15 10 9 9 7 11 1 9 9 1 13 9 13 4 2
30 16 9 1 9 2 9 13 1 11 1 0 9 1 11 11 1 11 11 1 13 4 16 11 11 1 11 1 9 13 2
13 3 10 9 1 15 14 12 0 9 9 13 4 2
22 15 13 9 1 1 9 13 1 0 2 0 9 9 7 0 9 1 1 1 0 9 2
10 10 9 9 1 9 13 4 4 4 2
30 11 11 11 2 11 11 11 11 2 11 2 1 9 9 1 13 4 16 10 9 1 10 9 9 1 0 13 4 4 2
16 9 1 9 9 2 9 9 2 1 9 9 11 1 13 4 2
17 15 1 9 7 9 1 9 9 1 1 0 9 1 9 13 4 2
12 15 1 11 11 1 1 14 9 8 13 4 2
15 7 2 10 10 9 1 1 9 13 1 9 13 4 4 2
23 9 1 9 8 13 1 3 15 12 9 1 1 12 1 12 9 1 1 9 13 4 4 2
18 9 1 10 9 1 13 1 1 9 9 9 1 0 13 4 4 4 2
10 15 9 9 9 1 9 13 4 4 2
21 15 9 1 9 9 0 9 1 7 14 9 9 1 3 14 0 13 4 4 4 2
15 9 1 10 9 9 1 1 9 9 1 9 13 4 4 2
16 15 15 13 4 4 4 16 9 9 9 1 9 14 13 4 2
27 11 1 9 9 11 11 11 1 13 13 16 13 1 12 2 12 9 1 10 9 9 1 0 13 4 4 2
14 9 13 16 15 9 2 9 3 1 1 10 0 13 2
30 15 9 1 1 9 14 1 9 14 12 12 9 8 13 4 7 2 10 9 1 1 10 9 12 12 1 13 4 4 2
48 11 9 1 9 1 9 1 0 9 1 3 13 1 1 9 11 11 1 0 0 9 1 11 11 11 7 11 11 2 11 1 11 11 15 1 13 4 7 9 1 1 0 9 2 9 13 4 2
24 9 15 13 15 11 1 0 9 1 10 9 1 9 13 16 9 1 15 13 1 14 13 4 2
20 9 14 15 1 10 9 13 4 16 15 2 15 1 13 1 0 14 14 13 2
19 15 1 0 9 11 11 7 11 11 11 1 9 1 0 13 1 9 13 2
8 9 11 1 14 9 1 13 2
38 11 1 0 9 11 11 1 11 0 11 11 1 11 1 0 9 1 9 1 2 0 13 2 1 1 15 7 12 0 9 1 1 11 0 13 4 4 2
50 11 2 11 11 2 11 11 1 11 1 15 9 13 4 13 16 11 2 11 11 1 9 11 11 11 2 11 11 11 11 1 9 9 11 11 7 12 9 1 1 11 11 11 1 11 0 13 4 4 2
53 11 1 13 16 11 11 11 2 11 2 1 11 11 2 9 2 2 11 2 11 11 2 0 9 2 7 11 2 0 9 1 0 9 1 1 1 9 2 1 0 9 1 1 10 9 1 1 9 0 13 4 4 2
46 15 15 14 13 16 0 9 1 10 9 3 13 4 16 11 15 11 1 9 13 14 13 4 2 16 9 9 2 9 9 7 0 0 9 1 9 1 15 1 15 9 1 15 9 13 2
29 0 13 16 11 1 9 9 1 1 1 11 1 1 2 9 2 9 13 1 11 11 10 9 1 9 13 4 4 2
9 11 11 10 9 11 1 9 13 2
14 15 13 16 10 0 9 1 0 9 13 4 4 4 2
30 11 9 1 0 9 1 11 11 9 1 1 0 9 1 1 11 9 11 1 11 11 9 1 0 9 11 1 13 4 2
23 13 4 9 9 1 14 0 12 9 1 9 1 13 4 4 2 15 15 9 13 4 4 2
20 11 11 9 1 10 9 1 11 2 11 7 11 9 1 10 9 1 9 13 2
17 11 1 1 9 2 9 2 9 7 0 9 9 1 12 9 13 2
28 0 9 1 9 9 11 11 1 9 9 1 13 16 13 4 9 11 14 11 11 1 9 11 1 13 1 13 2
18 11 9 1 0 13 9 13 1 0 11 11 9 1 11 0 9 13 2
22 11 11 1 9 1 9 9 1 13 4 1 3 11 1 9 1 11 9 1 9 13 2
25 11 11 1 12 9 1 1 13 11 1 0 11 1 12 9 1 9 13 0 9 1 9 13 4 2
40 10 9 1 9 1 1 0 9 1 9 1 11 11 1 11 11 1 12 9 1 1 11 11 1 13 4 7 9 1 12 9 11 7 11 1 0 13 4 4 2
23 0 9 1 15 1 11 1 9 13 2 16 9 1 9 13 9 1 9 15 13 4 4 2
27 0 9 1 9 11 11 1 13 16 9 1 9 11 11 1 9 13 4 16 11 1 11 1 13 4 4 2
18 9 3 9 11 11 2 11 11 7 11 11 1 9 1 13 11 13 2
17 11 1 11 1 11 11 9 1 12 9 1 13 4 1 9 13 2
9 10 9 9 9 9 1 13 4 2
21 0 9 1 9 1 11 11 1 9 9 11 11 1 1 13 4 9 1 9 13 2
14 9 1 11 1 9 1 1 13 15 15 9 13 4 2
16 9 1 1 1 9 1 13 4 9 1 11 1 9 13 4 2
28 9 9 11 11 1 13 16 11 10 9 1 13 4 15 11 2 11 2 1 0 11 9 1 12 9 13 4 2
10 11 15 1 9 1 9 1 9 13 2
13 11 1 13 16 11 1 9 9 9 13 13 4 2
18 9 1 13 1 0 9 7 12 9 1 9 1 9 13 4 4 4 2
12 11 11 1 9 1 14 9 1 15 13 4 2
17 9 1 11 1 9 7 9 1 12 9 1 12 9 0 13 4 2
28 11 9 1 11 11 1 9 0 13 0 9 11 11 1 1 0 9 1 0 13 1 15 15 9 1 0 13 2
16 9 9 1 13 16 9 1 9 1 0 13 1 9 14 13 2
49 9 11 11 11 2 9 11 11 7 9 11 11 1 9 1 11 1 9 1 9 12 9 1 1 13 4 7 11 9 1 9 1 9 13 1 9 1 0 9 1 0 9 0 13 1 9 13 4 2
23 9 1 11 1 1 9 0 13 1 11 9 1 13 4 2 9 2 1 14 9 13 4 2
42 11 11 1 9 9 1 1 0 9 1 0 13 4 4 16 2 9 2 11 1 1 2 1 3 13 1 15 9 14 13 2 16 15 9 1 9 13 1 9 14 13 2
14 10 9 1 3 13 9 1 0 9 1 0 13 4 2
10 16 10 9 9 1 11 1 0 13 2
38 11 9 1 11 1 1 0 9 1 9 1 0 13 1 9 13 4 9 1 0 9 11 11 1 0 9 1 10 9 1 3 9 13 1 13 4 4 2
18 11 9 1 15 9 1 13 16 9 0 9 1 9 1 13 4 4 2
17 11 9 1 15 0 9 1 13 4 16 9 9 1 9 14 13 2
42 0 13 16 11 11 11 1 11 9 1 11 7 12 9 1 1 9 0 13 4 7 11 11 11 1 11 2 11 2 11 2 11 7 0 9 1 1 9 13 4 4 2
20 11 1 11 11 1 9 1 9 13 7 0 0 9 0 13 15 9 14 13 2
29 9 9 1 9 7 9 1 9 13 1 1 11 1 9 1 11 1 11 1 12 9 1 1 15 9 0 13 4 2
25 11 1 11 9 1 9 1 1 0 7 0 9 13 1 1 12 0 9 2 9 1 9 13 4 2
13 7 11 11 1 9 1 0 9 3 14 9 13 2
57 0 11 7 11 1 9 11 11 11 1 9 1 11 0 9 1 12 9 1 13 9 1 1 9 1 11 1 9 11 11 1 9 1 13 16 10 9 1 11 9 1 0 9 14 13 1 1 15 12 0 9 9 1 9 13 4 2
8 11 1 15 0 9 0 13 2
35 11 1 0 9 11 11 11 1 1 2 9 1 15 9 1 9 13 16 15 1 0 9 1 1 9 1 9 14 13 1 9 14 13 4 2
20 9 1 9 1 9 13 1 1 11 1 3 10 11 9 1 9 13 4 4 2
20 9 1 9 1 9 1 9 13 1 1 11 1 11 1 10 9 1 9 13 2
23 10 9 1 9 1 9 0 13 13 4 16 15 9 1 9 1 1 9 1 9 0 13 2
15 11 1 9 1 9 1 9 10 9 1 1 9 13 4 2
22 11 9 11 11 11 1 13 16 11 11 1 9 0 13 1 15 0 9 14 13 4 2
18 11 1 12 9 1 9 1 9 7 11 9 1 9 1 9 13 4 2
7 7 10 9 14 0 13 2
14 9 1 1 1 9 1 9 1 15 9 14 13 4 2
29 11 1 9 1 0 13 4 11 1 13 16 3 1 11 9 1 1 11 14 12 9 1 11 1 9 13 4 4 2
26 11 1 9 1 9 1 0 9 1 13 4 4 16 9 1 9 1 1 0 9 15 3 0 14 13 2
22 0 9 1 9 1 0 9 13 4 7 15 10 9 1 13 1 1 10 9 0 13 2
18 11 9 1 9 1 0 9 1 11 11 11 1 14 9 13 4 4 2
29 9 1 13 4 4 16 11 10 0 13 4 4 16 0 9 1 0 9 1 13 15 1 14 15 9 13 0 13 2
43 11 1 1 11 1 11 11 1 0 9 1 0 13 4 1 3 0 9 9 1 9 13 4 0 9 1 12 0 9 1 9 1 13 0 9 1 9 13 1 9 13 4 2
39 12 9 1 11 1 12 9 9 1 0 9 1 1 9 13 1 3 11 1 11 1 13 4 9 9 1 0 9 1 12 9 9 1 9 1 0 13 4 2
34 15 1 11 1 9 1 9 1 1 9 1 9 13 4 4 2 7 0 7 0 9 1 9 1 1 13 1 9 9 1 13 4 4 2
17 0 9 1 0 13 1 1 9 1 10 12 9 1 9 0 13 2
34 3 11 1 11 11 11 1 13 16 11 7 11 1 1 1 9 1 0 13 1 3 15 1 1 11 1 9 1 13 15 9 14 13 2
17 15 13 16 15 10 9 13 2 15 15 15 15 1 13 4 4 2
24 15 13 16 9 10 15 14 9 14 13 2 15 1 10 15 9 13 2 15 15 1 0 13 2
26 11 1 11 11 11 1 13 16 11 1 9 0 9 1 9 1 13 9 2 9 7 9 0 13 4 2
48 11 1 9 1 0 9 1 12 9 1 1 1 9 1 0 13 1 9 1 9 13 1 9 13 4 4 2 7 10 14 9 1 13 13 16 9 1 9 1 1 9 13 1 15 9 14 13 2
33 9 1 9 13 1 9 9 9 11 11 1 13 16 15 13 13 16 9 0 13 4 4 7 12 0 9 1 9 0 13 4 4 2
22 9 1 11 1 13 16 9 9 13 1 3 15 1 9 1 7 3 0 9 13 4 2
27 15 1 14 9 1 0 9 1 1 9 9 13 1 15 9 1 9 13 1 13 9 3 13 1 9 13 2
46 11 11 11 11 1 9 1 1 11 1 13 16 14 12 2 12 9 1 0 9 9 1 0 9 1 13 4 7 15 9 1 9 13 4 16 15 15 9 1 15 0 9 14 13 4 2
23 15 13 16 10 9 0 14 13 16 9 9 0 9 1 1 13 1 15 9 1 9 13 2
16 15 13 16 11 11 11 11 11 0 13 16 12 9 9 13 2
21 15 13 16 9 9 1 0 9 1 9 1 1 15 1 15 9 14 13 4 4 2
26 11 11 11 11 10 9 11 1 1 0 9 1 9 1 1 12 12 12 9 13 1 9 13 13 4 2
22 7 9 9 1 0 13 4 4 16 15 11 1 9 1 9 13 1 15 9 14 13 2
21 9 1 11 1 0 11 11 11 11 1 11 1 9 1 9 13 1 9 13 4 2
15 9 9 9 1 11 1 15 13 9 1 10 9 13 4 2
22 9 1 9 9 1 0 9 1 13 4 1 11 9 1 9 1 14 0 9 13 4 2
26 9 1 0 9 1 13 4 4 16 9 9 1 0 9 1 13 1 9 1 9 1 3 9 13 4 2
35 9 1 1 11 11 1 9 13 4 11 1 9 7 9 9 11 11 1 13 16 9 1 13 4 0 9 1 9 13 4 1 9 13 4 2
16 10 9 1 9 13 1 1 9 11 9 9 1 9 13 4 2
22 9 11 9 7 11 9 9 1 0 9 1 9 13 1 0 15 9 11 9 1 13 2
17 11 7 11 1 9 3 11 11 7 11 11 11 1 10 9 13 2
8 9 0 9 13 1 9 13 2
14 9 1 11 7 11 9 1 9 1 9 14 13 4 2
15 11 1 1 9 9 1 0 9 1 13 12 0 9 13 2
7 15 15 15 9 14 13 2
23 15 13 16 9 1 9 1 9 1 11 7 11 9 9 1 9 1 9 1 14 9 13 2
18 7 15 1 9 11 7 11 9 9 1 0 9 1 1 13 4 4 2
18 9 11 1 9 1 1 9 1 9 13 1 1 9 14 1 9 13 2
15 11 1 9 1 1 12 0 9 9 1 14 9 13 4 2
26 9 14 1 12 9 9 1 9 13 9 1 1 11 11 11 11 1 11 11 2 11 1 9 13 4 2
21 14 12 9 13 9 1 0 9 1 12 9 1 1 12 0 11 1 0 13 4 2
13 11 1 11 11 0 12 9 1 14 9 13 4 2
16 11 1 13 16 9 1 1 1 15 9 1 14 14 13 4 2
16 9 1 10 0 9 11 1 9 9 1 11 9 9 9 13 2
18 14 12 0 9 1 9 1 9 1 0 9 1 9 1 9 9 13 2
10 10 9 1 1 9 1 9 13 4 2
22 9 1 9 13 4 9 15 9 7 9 1 9 1 9 1 9 1 1 1 0 13 2
22 9 1 13 1 12 9 1 11 11 11 11 7 11 11 11 11 11 11 14 0 13 2
13 11 7 11 3 0 7 0 0 9 0 13 4 2
16 12 9 1 9 13 4 1 3 9 11 7 11 1 13 4 2
24 9 1 10 9 1 10 12 9 1 0 9 1 9 1 1 15 2 15 1 9 1 13 4 2
21 12 9 12 9 0 2 0 9 1 11 1 11 11 2 11 11 11 1 9 13 2
13 11 1 15 0 9 7 9 13 9 1 9 13 2
22 9 2 9 7 9 1 9 13 1 11 11 1 1 9 13 7 0 9 1 0 13 2
20 15 9 1 1 9 13 2 9 1 1 9 13 7 13 14 15 0 13 4 2
10 9 9 11 11 9 9 13 4 4 2
11 11 1 9 1 10 9 9 1 9 13 2
12 11 1 13 16 9 1 15 9 9 0 13 2
12 9 1 14 15 9 1 9 1 0 13 4 2
25 11 1 14 15 1 13 16 9 1 1 16 15 3 10 9 15 9 1 13 4 16 15 13 9 2
31 11 11 1 1 9 13 1 9 15 13 2 15 13 4 1 11 1 13 16 12 9 15 11 1 9 1 9 13 4 4 2
19 3 11 1 9 11 11 15 1 13 7 15 15 9 9 13 1 9 13 2
7 15 15 10 9 0 13 2
8 15 10 9 15 9 13 4 2
19 15 1 11 1 11 1 15 1 0 10 9 13 15 11 1 0 13 4 2
19 11 1 13 16 15 1 8 9 0 9 1 3 14 0 13 13 4 4 2
13 10 9 1 11 11 1 1 15 9 14 13 4 2
8 10 9 9 1 1 1 13 2
14 11 1 13 16 15 9 14 9 1 0 13 4 4 2
20 15 0 9 13 16 0 9 13 1 1 15 15 9 1 0 14 13 4 4 2
15 11 1 13 16 9 13 1 3 14 15 9 13 9 13 2
15 11 1 13 16 11 1 9 1 1 15 9 10 13 4 2
18 15 0 9 11 11 11 1 9 1 10 9 9 1 9 2 9 13 2
14 15 11 14 1 9 1 9 1 9 1 9 13 4 2
26 11 1 13 16 15 15 15 11 2 11 2 11 7 0 9 1 13 4 15 9 9 1 13 14 13 2
26 15 9 1 13 4 13 16 15 12 9 15 9 9 11 11 1 15 1 9 1 9 13 1 13 4 2
23 0 0 9 1 9 13 1 3 11 13 9 1 9 9 15 9 11 9 11 11 1 13 2
27 11 1 0 9 1 0 11 9 1 1 9 13 4 4 7 11 9 15 14 0 9 0 13 1 13 4 2
18 11 11 1 1 1 11 1 11 1 9 1 9 13 4 1 9 13 2
15 11 9 1 1 11 9 7 15 0 9 9 14 0 13 2
43 11 9 1 1 9 11 11 2 11 11 11 2 11 11 2 9 11 7 11 11 1 9 0 9 1 3 9 1 13 3 11 1 11 11 11 1 9 14 9 1 13 4 2
10 15 9 11 1 0 9 1 14 13 2
20 11 1 9 9 13 1 3 15 11 1 1 11 1 9 0 9 13 4 4 2
23 11 9 11 11 1 9 9 7 9 1 1 1 0 13 15 9 1 14 13 4 4 4 2
33 7 11 0 9 1 0 12 9 1 11 9 1 9 1 13 9 11 1 9 1 1 0 9 13 15 9 9 1 13 1 9 13 2
18 11 9 1 9 1 9 1 13 1 9 11 1 0 9 1 13 4 2
19 11 9 1 12 0 9 1 0 9 1 0 13 1 9 14 9 14 13 2
28 16 0 13 4 4 12 9 9 1 11 9 1 9 13 4 1 9 14 9 9 1 0 9 1 13 4 4 2
30 11 1 1 0 13 4 11 11 11 11 2 11 11 7 11 11 1 9 14 12 12 9 9 9 11 11 1 9 13 2
7 15 14 10 9 1 13 2
32 9 1 9 1 11 1 9 7 12 9 1 1 12 11 11 1 13 16 15 9 1 9 1 0 9 9 9 1 13 4 4 2
12 11 1 11 15 13 10 9 11 11 14 13 2
15 3 11 7 11 9 1 9 11 1 14 11 1 13 4 2
25 9 1 13 16 11 9 1 9 11 11 1 9 11 11 1 9 1 9 9 11 11 1 9 13 2
16 9 1 10 10 9 1 11 1 9 13 4 1 9 13 4 2
7 7 15 9 14 13 4 2
19 11 9 1 9 12 9 3 9 1 0 9 1 9 9 1 13 4 4 2
34 13 4 4 4 16 11 0 9 9 9 11 11 1 1 15 0 13 1 13 4 4 16 9 1 11 1 9 1 9 1 0 9 13 2
11 3 9 1 1 10 9 1 9 13 4 2
12 11 11 1 1 9 13 0 14 13 4 4 2
18 11 9 1 9 13 16 11 11 11 1 0 9 1 0 0 9 13 2
12 3 11 11 1 1 10 9 1 9 0 13 2
19 15 13 13 16 9 9 1 15 9 1 14 13 4 1 15 10 9 13 2
15 15 11 1 9 14 13 7 15 1 15 9 14 13 4 2
29 9 1 1 16 9 1 15 9 1 9 13 4 4 2 16 9 1 0 9 1 15 10 9 1 9 14 13 4 2
14 9 1 9 1 15 9 13 1 9 1 10 9 13 2
13 9 13 1 15 15 9 1 9 13 1 9 13 2
22 11 11 1 13 13 9 1 9 13 1 9 1 1 1 9 1 13 1 9 13 4 2
20 11 11 11 11 1 13 13 16 15 14 9 1 9 14 13 1 0 9 13 2
17 15 14 13 13 16 9 9 1 9 9 1 13 1 9 13 4 2
40 10 9 1 0 11 1 0 9 11 11 7 11 11 1 13 16 9 9 1 10 9 11 11 1 12 9 13 15 0 13 1 1 15 0 10 9 1 0 13 2
19 9 1 9 13 1 0 9 1 1 15 12 9 1 9 9 13 4 4 2
15 9 1 9 1 9 9 0 13 1 9 9 13 4 4 2
31 10 9 1 11 11 11 1 9 11 11 11 11 11 11 2 11 2 1 0 9 9 1 9 9 1 9 9 13 4 4 2
7 9 9 12 9 1 13 2
23 16 10 9 1 9 9 1 9 13 4 16 15 10 9 1 9 1 11 1 0 9 13 2
21 9 9 1 9 13 1 9 1 9 1 9 9 1 13 2 15 9 1 13 13 2
23 9 9 1 9 1 1 1 9 11 7 9 11 9 11 11 11 11 1 9 11 13 4 2
10 9 15 9 1 9 1 9 9 13 2
16 11 11 11 1 0 9 11 11 11 14 15 1 9 1 13 2
28 9 11 1 0 9 11 11 1 11 1 0 9 1 10 9 13 7 13 14 13 15 9 0 9 1 13 4 2
16 9 1 9 15 1 13 15 15 9 1 1 9 9 13 4 2
12 0 9 1 9 1 14 10 3 9 14 13 2
29 12 9 1 11 11 11 1 0 9 11 11 11 1 15 9 7 9 1 9 1 15 9 9 13 1 9 9 13 2
31 11 11 11 11 1 9 1 0 13 9 1 14 15 0 9 13 7 0 9 9 1 9 1 9 9 9 9 9 13 4 2
7 10 9 1 0 9 13 2
23 15 1 0 13 9 1 9 9 1 9 13 4 0 9 11 1 12 9 9 1 13 4 2
13 10 9 1 9 11 1 0 9 0 13 4 4 2
12 9 11 1 15 11 11 11 1 1 13 4 2
13 15 9 9 1 11 11 1 1 0 9 9 13 2
42 9 9 9 1 1 9 1 15 1 11 7 11 2 11 2 2 11 11 11 2 11 2 2 11 11 2 11 2 7 11 11 2 11 2 9 9 0 13 4 4 4 2
19 11 0 9 1 15 11 11 11 11 1 10 9 9 7 9 13 1 13 2
22 11 1 11 1 0 9 0 11 11 1 1 0 9 9 1 1 9 1 9 13 4 2
33 11 11 1 12 0 9 11 2 11 11 7 11 1 1 9 9 9 11 11 11 1 9 1 12 2 12 0 9 1 9 13 4 2
9 10 9 9 7 9 1 9 13 2
22 15 9 11 1 9 1 13 9 7 9 7 9 9 1 9 9 1 10 9 1 13 2
20 13 4 4 16 11 11 11 11 1 9 9 11 1 1 15 1 1 9 13 2
23 0 13 16 11 11 1 10 9 1 0 9 13 4 2 7 15 15 0 9 14 13 4 2
29 9 1 1 9 9 11 11 11 1 9 1 11 11 11 11 1 9 1 0 9 1 0 9 13 1 9 13 4 2
14 10 9 11 11 1 12 9 1 12 9 1 9 13 2
9 10 12 14 9 1 9 11 13 2
15 9 15 9 7 9 0 13 1 1 3 9 13 4 4 2
16 11 1 0 9 1 9 13 1 9 1 9 1 0 13 4 2
27 11 11 1 11 1 0 9 1 12 9 1 13 7 12 9 1 10 9 1 0 13 1 9 14 13 4 2
19 11 1 11 1 9 2 9 13 1 3 9 1 0 9 3 13 4 4 2
10 14 15 9 9 12 12 13 4 4 2
23 9 1 12 12 9 0 0 9 1 12 9 9 1 15 14 12 12 9 9 13 4 4 2
13 9 1 9 1 9 14 11 1 9 13 4 4 2
18 10 9 1 9 1 9 1 9 14 1 14 9 13 1 9 13 4 2
33 11 11 1 9 7 9 1 9 13 4 11 11 11 11 1 11 1 13 2 9 1 9 1 10 15 13 9 1 9 13 0 13 2
16 9 1 12 9 1 9 9 9 1 9 9 1 13 4 4 2
19 9 1 9 7 9 1 9 7 9 1 9 9 9 1 13 4 4 4 2
26 11 1 11 1 11 11 1 9 13 1 3 15 11 1 11 9 1 9 13 1 9 0 13 4 4 2
38 11 1 11 1 11 1 11 1 9 1 13 4 4 2 7 10 9 1 11 1 9 13 4 1 1 11 1 9 1 9 9 1 9 13 4 4 4 2
15 11 1 9 1 9 13 4 1 11 1 0 9 13 4 2
28 11 1 11 1 1 9 13 13 1 11 1 9 11 1 9 14 13 4 2 7 15 11 11 11 13 4 4 2
23 11 9 11 11 1 13 1 11 1 9 11 11 1 11 1 14 15 11 1 13 4 4 2
28 11 1 11 1 9 1 9 1 9 1 9 1 1 9 11 1 9 1 9 0 13 12 0 9 13 4 4 2
36 11 7 11 15 10 9 1 13 4 4 16 11 1 12 9 11 11 15 9 9 13 1 9 13 4 16 15 15 9 14 15 9 0 13 4 2
46 15 1 1 9 1 0 13 4 16 11 1 11 1 12 9 1 1 14 9 1 12 7 11 1 12 7 11 1 12 9 1 9 11 1 12 9 1 13 4 4 15 14 12 13 4 2
10 10 9 11 1 12 1 10 13 4 2
15 15 1 14 15 9 1 3 0 9 13 1 3 13 4 2
36 9 1 1 10 9 1 0 0 9 1 0 9 13 1 11 7 11 11 1 14 9 13 4 4 4 7 10 9 11 11 1 0 13 4 4 2
13 11 1 13 11 11 14 10 9 1 13 4 4 2
22 11 1 9 1 9 0 13 1 3 11 11 1 1 14 3 9 1 9 13 4 4 2
47 11 1 9 1 0 13 4 4 16 11 1 10 9 0 13 4 4 16 15 11 7 11 1 14 12 9 1 9 13 1 9 13 4 4 2 15 11 1 10 9 1 1 0 13 4 4 2
26 7 2 0 9 1 1 0 11 11 15 2 0 9 2 1 0 9 13 1 15 9 14 13 4 4 2
18 9 1 9 1 11 1 15 7 12 9 1 1 9 0 13 4 4 2
30 3 11 11 1 11 11 1 9 9 1 1 9 1 9 1 9 1 13 4 11 1 9 1 3 13 1 9 13 4 2
13 15 9 1 0 9 1 15 0 13 1 13 4 2
34 10 9 1 1 9 1 11 1 11 1 11 11 9 1 9 1 9 9 11 11 7 0 11 11 11 11 1 9 1 9 13 4 4 2
35 15 1 11 1 9 7 9 9 9 1 0 9 1 9 1 1 9 1 1 11 9 11 11 11 1 1 14 9 1 9 13 4 4 4 2
10 12 9 11 7 11 14 13 4 4 2
12 7 11 9 15 14 9 1 9 1 3 13 2
28 11 1 9 1 15 11 9 9 11 2 11 2 11 2 11 8 13 4 7 9 1 9 0 13 1 9 13 2
60 11 1 0 0 9 11 11 1 11 9 11 11 11 1 9 1 9 7 10 9 9 1 9 1 9 7 9 13 1 9 1 11 9 2 15 9 11 11 7 11 1 11 1 9 9 9 9 11 14 11 11 11 1 1 0 9 0 13 4 2
26 3 11 1 13 13 16 9 1 9 7 9 1 9 1 1 9 7 0 9 1 0 9 13 4 4 2
27 9 9 9 11 11 11 11 1 13 16 11 11 11 1 9 11 11 1 3 9 1 0 13 4 4 4 2
15 11 11 1 15 1 15 9 9 9 1 0 14 13 4 2
40 11 1 11 9 1 11 9 1 0 9 1 11 11 2 15 9 11 11 2 0 9 9 11 11 2 0 9 11 11 7 11 9 11 11 1 0 13 4 4 2
35 11 1 9 11 11 1 13 16 11 11 7 0 9 9 1 1 11 11 1 0 9 1 13 1 9 13 1 9 1 9 0 13 4 4 2
19 9 1 11 11 1 0 9 1 11 9 0 9 1 0 2 0 13 4 2
11 9 9 9 1 13 2 8 4 13 4 2
12 15 9 1 9 12 9 9 1 1 13 4 2
15 13 1 12 9 1 1 9 1 0 9 13 1 9 13 2
13 9 1 1 13 1 0 9 1 9 0 13 4 2
17 0 9 1 9 1 9 2 9 9 13 4 15 9 9 0 13 2
29 11 1 13 9 1 1 9 1 10 9 1 11 1 3 13 9 1 9 1 9 1 1 13 9 1 10 9 13 2
20 9 1 9 13 16 9 1 9 9 14 13 1 1 9 1 10 9 13 4 2
12 9 1 13 1 1 14 0 9 14 13 4 2
21 11 11 1 0 9 1 9 7 0 7 0 9 1 9 1 9 1 9 13 4 2
11 11 7 15 1 1 9 1 3 9 13 2
16 11 1 9 3 13 0 9 1 9 1 9 1 0 13 4 2
22 9 9 1 12 9 1 1 0 9 1 11 1 9 1 10 9 1 9 14 13 4 2
10 10 11 1 9 0 7 11 11 13 2
20 11 1 14 9 1 11 7 11 1 1 10 9 1 9 13 9 13 4 4 2
28 15 11 11 11 1 13 9 1 9 1 11 7 11 1 1 13 10 9 1 9 1 15 3 13 9 13 4 2
21 9 9 12 12 9 1 1 11 7 0 11 1 0 9 1 0 9 9 13 4 2
24 11 11 2 11 2 11 7 11 11 1 10 0 2 0 9 1 14 9 13 1 9 13 4 2
12 9 9 1 1 0 12 9 1 9 0 13 2
6 15 9 1 9 13 2
14 11 1 9 9 1 1 9 1 9 12 9 9 13 2
22 7 0 9 13 1 1 1 9 1 9 12 9 9 3 13 12 9 9 1 13 4 2
18 0 9 1 1 9 1 14 12 9 14 9 1 9 1 9 13 4 2
17 16 15 15 1 15 9 2 9 1 9 1 9 14 13 4 4 2
22 9 7 9 1 9 11 11 1 9 1 9 11 1 11 7 11 0 9 1 13 4 2
29 11 1 0 9 11 1 9 13 3 12 0 9 9 1 12 9 1 9 13 4 7 12 1 10 9 0 13 4 2
21 11 11 11 11 11 1 11 11 1 11 11 11 1 11 1 0 9 1 9 13 2
8 11 11 1 11 13 4 4 2
15 11 1 13 9 9 1 11 9 7 11 9 1 13 4 2
23 11 9 9 9 1 0 9 11 11 1 13 16 0 9 12 9 1 11 9 9 1 13 2
14 10 9 1 12 9 13 4 7 12 9 0 13 4 2
26 9 1 10 9 10 9 13 16 10 14 9 1 11 7 0 11 1 1 13 1 9 9 13 4 4 2
27 9 1 10 9 1 9 14 13 2 15 11 1 11 11 9 1 11 13 1 1 9 1 9 13 4 4 2
29 9 1 1 9 9 1 1 13 9 10 0 13 16 9 9 1 9 2 9 9 7 9 9 0 9 0 13 4 2
10 10 9 1 9 1 9 14 13 4 2
31 10 9 1 0 12 9 1 13 16 9 1 1 9 1 9 9 13 4 4 7 0 9 1 9 1 9 9 13 4 4 2
12 15 10 9 1 14 0 9 11 9 1 13 2
19 10 9 1 12 9 1 9 1 14 9 13 4 7 12 9 0 13 4 2
14 9 1 1 3 1 12 9 1 9 1 9 13 4 2
26 15 10 9 1 9 1 1 11 1 9 11 11 11 1 9 1 12 0 9 9 1 9 13 4 4 2
46 9 1 1 0 9 1 0 11 1 12 9 1 9 1 11 9 1 11 11 11 1 11 0 9 1 9 12 9 9 13 12 9 1 13 4 7 12 9 1 0 9 1 0 13 4 2
21 14 10 9 10 9 1 11 1 9 1 9 13 12 9 1 9 1 9 13 4 2
28 9 1 12 0 9 1 11 1 9 1 11 1 11 13 4 12 9 1 9 13 7 12 9 1 0 13 4 2
26 9 1 11 9 1 12 9 9 1 9 13 9 1 12 9 1 13 4 7 12 9 1 0 13 4 2
35 12 0 9 1 9 1 11 9 1 11 9 9 1 10 9 1 9 9 0 9 9 13 12 9 1 13 4 7 0 9 1 0 13 4 2
11 10 9 1 12 1 10 9 0 13 4 2
19 10 9 1 11 1 9 1 9 1 9 13 9 0 12 9 1 13 4 2
22 9 1 11 11 9 1 11 1 9 1 9 1 9 13 11 1 12 9 1 13 4 2
12 10 9 12 9 1 13 1 9 13 4 4 2
31 11 1 0 9 1 9 11 11 2 11 11 1 11 1 14 9 14 9 9 9 13 4 7 0 3 11 1 9 13 4 2
32 11 11 11 1 11 2 11 11 2 11 11 11 2 1 13 9 9 7 0 9 9 1 3 15 9 13 1 9 13 4 4 2
11 9 9 1 9 1 11 1 14 9 13 2
38 9 11 11 7 9 11 11 1 9 1 1 11 11 11 1 13 9 1 9 9 1 9 0 13 9 1 9 13 1 9 1 9 13 1 9 13 4 2
25 9 1 13 4 4 16 9 0 14 13 7 9 1 15 0 13 4 13 1 9 0 13 4 4 2
22 7 9 1 9 1 0 9 1 9 13 4 2 7 9 1 9 13 1 9 13 4 2
16 15 9 9 9 1 9 1 10 0 9 1 13 1 13 4 2
30 9 9 1 10 9 1 1 9 9 1 9 1 9 1 9 1 14 13 1 9 13 4 7 9 15 13 1 0 13 2
11 15 9 9 1 9 10 13 13 4 4 2
7 15 1 9 1 13 4 2
12 11 1 14 11 11 2 11 1 9 0 13 2
21 9 1 9 2 9 9 11 11 7 11 11 1 9 1 1 9 13 9 0 13 2
32 15 13 13 16 9 9 9 1 9 13 0 12 9 1 9 1 9 13 4 7 15 13 1 1 15 1 9 1 9 14 13 2
9 10 9 1 14 9 9 1 13 2
38 9 9 10 9 1 9 9 1 14 0 13 2 15 10 9 1 13 13 16 13 1 12 9 1 9 9 13 4 4 15 1 10 9 1 0 9 13 2
21 9 11 11 1 13 13 16 11 11 9 9 9 1 0 9 13 9 13 4 4 2
25 9 1 11 1 13 4 0 9 11 11 14 11 1 12 9 1 9 9 1 9 1 0 13 4 2
14 9 1 9 13 16 15 14 0 9 1 0 13 4 2
18 0 9 11 11 11 2 11 2 7 11 2 11 2 1 13 4 4 2
8 15 9 11 11 1 13 4 2
11 9 1 15 9 13 0 9 0 13 4 2
22 13 4 9 1 9 11 1 9 9 1 13 9 9 1 9 1 14 9 13 4 4 2
22 9 1 11 1 11 11 11 1 9 1 9 1 9 7 9 13 1 9 9 13 4 2
17 9 11 11 1 13 16 9 1 10 9 1 0 9 13 4 4 2
18 11 0 11 11 11 1 9 1 11 11 1 12 9 1 9 13 4 2
5 11 15 0 13 2
10 15 9 1 9 9 1 13 4 4 2
17 9 9 1 13 16 0 9 11 2 11 1 11 9 1 9 13 2
18 15 10 9 1 13 4 2 10 9 1 11 1 9 11 14 13 4 2
10 10 9 15 9 11 1 14 13 4 2
14 11 2 11 1 0 0 13 1 3 11 11 13 4 2
9 11 15 15 9 13 9 13 4 2
11 15 12 9 1 1 9 9 1 13 4 2
17 15 1 11 9 1 14 9 1 13 11 7 11 1 9 13 4 2
32 11 1 9 1 13 16 15 10 9 1 11 11 11 1 9 1 1 0 11 9 13 4 4 2 15 15 9 1 13 13 4 2
27 10 9 1 11 9 1 15 1 9 1 14 13 4 2 7 11 7 15 12 9 11 9 1 9 14 13 2
6 11 13 11 13 4 2
13 15 15 9 13 4 7 15 1 15 11 13 4 2
19 11 1 1 11 1 9 9 1 9 0 13 7 15 1 15 11 13 4 2
11 9 1 9 13 1 11 1 15 11 13 2
8 11 13 1 1 15 11 13 2
15 15 11 1 9 1 15 11 1 9 13 7 11 13 4 2
17 11 1 15 11 1 9 13 7 2 11 1 0 9 1 13 4 2
18 15 1 11 11 1 0 9 11 11 11 15 11 1 1 11 13 4 2
41 11 1 9 13 16 11 1 11 1 9 1 11 1 11 13 1 15 12 9 2 9 2 12 11 2 12 2 12 9 11 2 9 2 9 9 7 0 9 13 4 2
11 11 1 12 9 1 15 9 9 13 4 2
14 10 9 15 11 1 14 12 9 1 9 13 4 4 2
23 11 11 1 11 1 11 7 9 9 1 9 1 0 9 13 1 9 1 9 13 1 13 2
26 9 1 0 9 1 9 13 4 13 16 9 1 15 10 14 10 9 1 9 1 9 13 4 4 4 2
39 9 11 11 11 7 9 11 11 11 1 13 16 11 11 1 11 11 1 1 9 1 9 13 4 4 16 15 9 1 9 1 9 1 9 13 1 9 13 2
39 9 1 13 16 15 13 4 16 15 10 0 9 13 4 4 15 9 7 11 11 1 11 11 1 9 1 0 13 1 1 9 1 9 13 1 9 13 4 2
26 11 11 1 11 11 1 11 11 1 0 9 1 1 11 1 9 1 9 1 1 9 1 10 9 13 2
17 9 1 9 1 12 9 9 1 9 9 13 1 9 13 4 4 2
10 9 1 9 1 9 1 9 13 4 2
27 13 16 9 1 11 11 1 1 9 1 9 1 9 1 13 7 9 1 9 9 1 13 1 9 13 4 2
30 3 10 9 1 14 9 13 16 9 1 0 9 1 13 9 1 1 0 0 9 7 0 9 1 9 1 9 13 4 2
31 10 9 11 11 1 1 9 1 0 0 9 9 9 1 13 4 4 16 10 9 1 15 9 1 1 0 14 13 4 4 2
15 7 15 9 1 9 1 1 15 0 9 1 10 14 13 2
18 15 15 9 1 9 13 16 15 10 9 1 0 13 1 1 9 13 2
24 9 1 13 16 10 0 9 13 16 9 1 9 9 9 1 9 1 9 1 13 4 4 4 2
10 10 0 9 1 9 9 13 4 4 2
26 11 11 11 1 9 11 11 1 9 1 1 11 9 13 1 9 1 12 9 3 9 1 9 13 4 2
28 11 1 15 13 16 16 0 11 11 13 16 10 9 1 13 1 9 1 15 12 9 3 15 9 13 4 4 2
30 0 13 16 11 9 1 1 9 1 12 9 1 9 1 9 13 11 9 13 1 9 13 4 7 9 14 13 4 4 2
20 11 2 11 1 11 9 1 9 1 11 1 12 9 1 9 13 9 13 4 2
27 0 9 1 1 9 11 11 1 11 9 0 15 9 1 13 13 4 7 9 13 1 3 15 9 13 4 2
15 9 1 11 1 9 0 13 15 9 1 1 13 4 4 2
18 3 9 1 11 9 1 11 1 9 1 12 9 1 9 1 9 13 2
14 0 9 1 13 16 9 1 13 1 15 0 14 13 2
19 9 1 13 16 9 1 11 1 3 0 11 11 1 1 9 1 9 13 2
13 10 9 1 9 9 7 9 1 0 9 13 4 2
15 9 9 1 9 1 11 12 3 10 0 9 13 4 4 2
28 15 13 4 4 4 16 13 1 3 9 1 9 13 4 1 9 1 9 13 1 9 1 9 1 9 13 4 2
16 10 9 1 9 1 1 9 1 9 1 14 3 9 13 4 2
18 9 1 9 1 9 13 1 1 11 11 11 11 9 11 1 13 4 2
17 9 1 9 1 9 13 1 1 1 9 0 13 1 9 13 4 2
22 7 0 9 1 10 9 0 13 4 16 9 1 10 9 9 1 10 0 13 1 13 2
18 11 11 1 11 11 1 12 9 1 10 9 1 9 13 10 9 13 2
65 2 11 11 11 11 11 11 11 11 2 1 13 4 4 16 9 1 11 2 11 2 2 11 2 1 13 4 4 16 15 14 0 9 1 15 9 1 12 9 1 1 14 9 1 13 4 4 4 2 7 10 9 1 1 9 1 0 9 1 0 14 13 4 4 2
29 15 1 9 1 9 1 9 1 9 14 10 9 13 4 4 2 15 9 1 1 0 0 9 1 0 13 4 4 2
17 9 1 9 11 11 11 1 11 11 11 11 1 9 1 13 4 2
43 9 1 15 13 4 4 16 15 9 1 2 9 2 9 13 1 3 15 9 1 9 1 13 4 4 4 2 7 15 1 1 9 1 9 13 1 3 14 9 0 13 4 2
11 16 10 0 9 1 10 9 13 4 4 2
31 15 15 0 13 4 16 9 9 1 9 1 13 4 4 2 7 0 3 9 15 9 1 9 1 9 13 1 9 13 4 2
28 9 1 13 4 4 16 10 9 9 9 1 12 12 9 13 4 2 15 1 12 12 9 1 9 9 13 4 2
25 16 9 1 10 9 1 0 9 1 0 13 4 4 16 9 1 9 1 9 1 13 4 4 4 2
20 11 1 10 9 12 12 9 1 14 12 9 9 9 1 9 1 9 13 4 2
19 0 9 1 9 1 0 9 1 9 1 9 9 1 9 1 13 4 4 2
17 10 9 13 16 0 9 1 15 11 1 1 13 9 13 4 4 2
12 13 4 4 16 11 0 9 1 0 9 13 2
29 11 2 11 7 11 1 0 9 13 4 16 15 9 9 1 9 1 9 13 0 9 1 1 15 9 13 4 4 2
12 11 14 3 14 10 9 1 9 13 4 4 2
22 0 9 1 13 16 10 9 1 11 11 1 13 4 16 15 9 9 1 9 14 13 2
15 0 9 15 14 9 1 13 12 9 1 9 13 4 4 2
18 11 1 9 11 11 1 11 1 12 0 9 11 1 9 13 4 4 2
18 10 9 1 1 11 9 9 9 1 9 1 9 13 1 0 9 13 2
14 15 11 1 9 13 4 4 16 9 1 11 13 4 2
13 9 1 13 16 0 0 9 1 9 1 9 13 2
12 10 9 9 9 9 1 9 1 9 13 4 2
17 9 9 1 9 1 11 1 9 1 9 1 9 13 14 4 4 2
19 11 1 9 1 1 11 7 11 1 9 1 12 9 9 1 9 13 4 2
12 11 1 10 9 10 9 9 13 4 4 4 2
14 0 11 11 11 11 1 0 9 11 1 9 13 4 2
10 11 11 1 11 1 9 1 13 4 2
17 11 1 11 1 9 13 1 1 9 9 1 9 14 13 4 4 2
31 11 1 9 1 1 12 9 14 9 13 4 2 15 12 9 1 9 2 9 7 9 1 1 9 0 13 1 9 13 4 2
26 11 11 1 11 1 0 13 4 16 3 0 9 1 11 9 1 9 7 9 1 9 13 4 4 4 2
11 7 11 1 9 1 0 9 1 9 13 2
36 9 11 11 11 1 9 1 9 1 0 9 11 11 1 11 9 1 9 1 13 4 9 1 13 4 4 12 9 1 9 9 1 1 1 13 2
23 9 1 9 1 10 9 11 9 1 1 1 13 9 9 11 11 11 1 13 1 9 13 2
33 11 1 9 13 16 11 1 9 9 1 0 9 1 9 0 13 7 15 9 13 1 1 1 12 9 2 9 0 13 4 4 4 2
28 11 1 9 13 16 0 9 1 9 13 1 1 9 11 1 9 1 13 0 9 2 9 1 9 13 4 4 2
23 11 11 11 11 1 9 1 0 9 1 3 13 1 13 1 9 1 1 1 9 13 4 2
27 11 1 13 4 16 11 9 1 11 9 1 9 1 1 0 9 1 9 0 9 1 13 4 0 9 13 2
19 15 11 9 1 10 9 1 9 13 2 15 0 9 1 0 13 4 4 2
37 11 9 11 11 1 13 16 11 11 7 15 9 10 9 1 9 10 3 13 4 4 7 15 1 11 7 11 9 1 9 13 4 9 1 9 13 2
35 11 1 10 9 1 9 13 16 11 11 1 0 9 11 11 11 1 9 9 9 1 13 4 14 15 9 13 1 1 10 9 0 13 4 2
19 15 10 9 1 9 0 13 1 3 11 11 1 0 9 1 9 13 4 2
40 11 1 13 16 0 9 1 9 9 9 10 9 1 9 13 16 9 1 11 9 1 1 9 7 9 1 9 1 0 13 4 9 1 9 1 9 9 13 4 2
49 10 9 10 9 1 13 4 4 16 11 9 1 0 9 9 1 13 4 4 4 7 10 9 1 9 13 4 4 4 16 11 9 1 9 11 11 11 1 10 0 9 1 12 9 1 13 4 4 2
14 10 9 1 1 0 9 1 9 14 13 4 4 4 2
70 15 1 9 11 11 11 1 9 1 12 0 9 1 9 13 7 15 10 9 1 9 13 1 1 13 13 16 2 11 11 1 11 11 11 2 11 1 9 15 13 2 15 1 10 9 0 15 13 2 7 10 9 1 9 1 9 1 9 1 10 9 9 13 2 15 15 1 0 13 2
33 11 11 2 11 2 1 11 11 11 11 1 13 16 9 11 1 11 11 1 0 9 11 11 1 9 1 1 3 9 13 4 4 2
20 11 1 11 1 12 9 1 9 1 13 16 11 1 9 1 9 0 13 4 2
28 15 13 16 16 3 9 13 1 13 9 13 4 2 16 15 0 9 13 16 9 11 1 9 1 1 9 13 2
12 15 15 9 14 13 16 15 9 1 9 13 2
33 9 1 3 13 1 9 1 9 1 1 1 13 4 1 15 13 16 11 11 1 11 1 11 1 14 13 1 10 0 9 13 4 2
36 11 11 15 0 9 1 9 1 0 13 4 2 7 15 15 9 1 0 13 4 16 15 3 9 13 7 11 1 0 13 7 15 1 9 13 2
48 0 9 1 9 1 3 9 13 4 0 13 7 0 0 9 1 11 11 1 1 1 10 9 1 3 13 1 9 1 15 13 16 9 1 0 9 1 1 1 15 10 13 1 9 1 14 13 2
20 11 1 13 16 15 12 9 13 4 4 16 9 13 4 16 9 1 9 13 2
12 15 13 16 15 1 1 9 9 3 9 13 2
26 15 13 16 11 11 1 1 10 15 9 14 13 2 15 15 0 9 1 9 13 1 1 0 13 4 2
18 9 1 9 0 9 1 0 13 4 4 7 15 3 1 0 13 4 2
11 15 15 9 14 13 16 9 3 10 13 2
20 11 11 11 7 0 9 11 11 12 9 3 12 9 1 3 9 13 4 4 2
16 9 9 1 1 15 1 9 9 1 0 9 14 13 4 4 2
18 11 9 9 3 11 11 1 9 9 1 0 13 1 9 13 4 4 2
19 9 9 1 9 13 16 11 1 1 9 1 9 1 1 13 4 4 4 2
15 7 9 9 1 11 1 0 9 9 1 13 0 14 13 2
17 9 9 1 1 11 9 11 11 13 4 16 11 1 15 9 13 2
17 15 1 15 15 15 1 11 11 1 9 9 1 13 4 14 13 2
15 11 11 11 1 11 1 10 9 1 0 13 1 9 13 2
14 15 1 11 11 11 1 1 9 1 9 13 4 4 2
15 11 9 11 11 1 12 0 9 1 0 13 1 9 13 2
19 10 9 1 11 11 2 9 9 11 11 7 11 1 0 9 14 0 13 2
12 15 1 11 9 10 0 9 1 14 0 13 2
24 11 2 11 1 11 9 1 9 1 9 1 11 1 9 1 9 13 1 12 9 1 13 4 2
16 9 1 9 9 1 1 9 1 1 9 1 9 13 4 4 2
9 10 9 11 11 1 9 1 13 2
21 9 1 13 16 11 9 1 11 9 1 9 9 1 1 9 9 13 4 4 4 2
15 10 3 12 9 1 13 9 1 9 1 9 9 13 4 2
14 0 9 1 9 1 15 9 1 9 1 9 14 13 2
23 0 9 1 1 9 1 0 9 1 9 13 1 9 9 1 12 9 1 0 9 13 4 2
31 0 9 1 13 16 9 1 9 1 3 2 3 9 1 9 13 2 7 15 15 13 1 9 13 4 7 3 9 13 4 2
24 9 1 15 9 1 9 14 13 15 9 1 13 9 1 10 9 1 15 9 1 9 14 13 2
22 9 1 9 13 1 1 9 1 0 9 1 9 14 13 4 2 7 9 9 13 4 2
15 15 1 9 1 9 1 9 13 7 12 9 1 13 4 2
19 15 9 1 9 7 15 9 1 1 1 15 9 1 9 14 13 4 4 2
19 11 1 11 11 1 9 13 1 9 13 14 10 10 9 0 13 4 4 2
25 9 1 10 9 1 11 2 11 2 7 11 1 9 1 1 9 1 11 13 1 9 13 4 4 2
14 7 9 9 1 9 9 13 11 1 15 9 13 4 2
21 15 1 14 15 1 9 13 10 10 9 9 1 9 11 1 9 1 3 13 4 2
23 0 9 9 11 11 1 13 16 10 10 0 9 1 9 1 9 11 13 4 11 13 4 2
10 15 1 10 9 9 1 1 11 13 2
15 15 1 14 12 9 9 13 1 9 9 1 1 11 13 2
29 11 9 9 1 9 10 9 1 1 9 1 9 14 13 15 1 0 9 9 11 11 7 11 11 9 9 1 13 2
36 1 11 2 15 10 9 1 9 13 1 1 9 9 1 14 13 4 16 15 15 1 13 11 11 13 1 9 1 9 13 1 1 15 13 4 2
27 0 13 16 9 9 1 11 1 11 13 1 13 14 10 14 10 12 9 0 9 9 1 1 3 13 4 2
27 10 9 1 12 0 2 0 9 13 4 4 7 10 9 1 15 13 1 0 9 1 9 15 1 14 13 2
33 11 1 0 9 13 4 1 9 1 9 13 4 11 11 1 11 1 10 9 1 12 9 1 9 1 0 13 1 9 0 13 4 2
25 10 9 1 0 9 1 9 1 1 0 9 7 11 11 1 0 11 11 11 1 9 0 13 4 2
22 11 11 1 1 11 1 10 9 1 11 1 0 11 11 1 9 1 14 0 9 13 2
34 16 3 1 11 11 1 0 9 1 11 9 11 11 1 15 0 0 9 1 13 16 11 9 1 11 1 9 1 15 15 14 13 13 2
17 11 11 1 13 16 11 11 1 9 9 1 1 9 1 9 13 2
13 9 1 13 4 9 11 1 14 0 13 4 4 2
30 15 1 9 1 11 1 11 11 2 11 1 9 1 0 9 11 11 1 9 0 13 1 3 9 1 9 0 13 4 2
44 7 0 11 11 11 11 1 9 13 7 11 11 11 1 9 1 1 1 3 13 1 9 1 9 1 9 9 11 11 1 13 16 10 9 1 15 0 9 13 1 3 9 13 2
15 16 9 1 13 16 15 13 1 9 13 16 15 15 13 2
14 16 0 9 1 13 4 16 15 13 1 9 14 13 2
46 16 15 9 0 13 1 3 14 11 1 9 13 16 15 11 1 0 11 11 7 11 9 1 9 1 11 7 11 1 9 1 11 1 11 9 1 11 11 11 11 9 1 9 0 13 2
27 15 11 11 9 1 1 1 13 4 9 1 1 9 1 13 16 15 0 9 11 1 1 0 14 13 13 2
43 11 11 11 1 9 11 11 1 10 9 1 9 13 4 4 16 11 2 11 7 9 9 1 11 11 1 9 1 11 1 9 1 9 1 0 9 1 13 1 9 13 4 2
42 9 9 1 10 9 1 11 1 0 9 11 11 0 13 16 11 7 9 1 11 1 9 13 4 0 9 1 9 13 4 14 2 11 11 11 1 9 13 1 9 13 2
22 11 1 11 1 14 9 1 9 1 9 14 13 4 15 9 9 1 10 9 13 4 2
44 3 1 11 11 1 9 13 4 11 9 11 11 1 13 16 11 9 9 1 12 9 1 9 1 0 13 4 4 7 10 9 10 0 13 16 9 1 15 14 0 9 13 4 2
51 0 9 1 9 0 13 1 11 11 1 9 1 9 1 9 1 13 9 13 1 3 11 1 9 9 9 11 11 11 1 13 16 16 9 1 0 9 15 9 1 9 13 4 16 9 15 9 13 4 4 2
29 15 11 1 0 12 9 1 15 13 16 9 1 12 9 9 2 9 7 9 1 9 1 9 1 1 9 13 4 2
18 15 16 15 14 15 9 1 1 13 4 16 9 15 9 13 4 4 2
25 15 13 16 15 9 1 9 13 16 15 15 0 13 16 9 1 0 9 9 1 9 1 1 13 2
47 9 7 9 1 1 9 1 0 9 13 4 9 11 1 13 16 9 1 12 9 1 15 9 1 9 0 9 1 13 4 7 9 1 10 9 1 9 1 1 15 2 15 1 0 13 4 2
32 9 13 1 9 1 9 1 9 9 1 13 16 0 9 7 9 1 9 1 9 1 0 9 1 12 0 9 1 9 13 4 2
14 15 9 1 13 1 9 1 9 1 14 0 9 13 2
35 15 1 1 9 13 4 15 13 16 11 1 14 12 9 9 0 9 1 8 13 4 4 2 15 1 12 9 9 1 9 0 13 4 4 2
24 9 9 1 0 13 4 9 7 0 9 1 9 1 1 15 0 9 14 13 4 1 9 13 2
18 15 13 16 11 11 11 1 9 14 15 0 9 1 9 13 4 4 2
19 9 11 1 9 13 16 0 9 1 11 11 1 9 3 14 0 13 4 2
12 10 9 9 9 1 15 0 13 1 0 13 2
36 10 9 1 9 11 1 9 1 3 9 13 4 11 11 1 11 11 11 1 9 1 9 1 9 9 13 1 1 12 12 9 13 1 9 13 2
16 11 1 13 16 0 9 1 10 9 12 12 9 13 4 4 2
32 9 1 11 11 11 1 9 9 1 10 9 1 9 0 13 16 9 7 9 15 2 15 1 0 13 7 15 9 13 0 13 2
29 9 9 1 9 9 1 9 7 9 1 9 13 1 1 11 7 9 1 11 11 11 11 1 9 1 14 9 13 2
37 15 9 1 11 1 13 16 9 9 1 0 2 0 12 12 9 1 0 13 4 1 9 13 4 4 2 15 1 12 12 9 0 14 13 4 4 2
13 15 9 1 1 0 13 9 1 13 1 9 13 2
37 15 0 9 11 1 11 1 9 7 9 9 13 1 13 13 9 1 1 9 1 0 9 1 13 1 1 9 1 9 7 9 9 1 9 13 4 2
11 9 1 9 9 1 13 1 9 13 4 2
19 16 9 1 1 9 11 11 7 12 9 11 11 1 10 9 0 13 4 2
11 11 11 1 1 11 1 1 10 9 13 2
13 7 11 13 1 1 15 9 14 9 13 13 4 2
14 10 11 1 11 7 11 15 2 15 9 13 4 4 2
10 10 9 0 9 0 13 4 4 4 2
18 7 9 1 9 12 1 12 9 1 11 1 9 13 1 9 13 4 2
25 10 9 0 9 1 9 11 1 11 1 9 13 4 7 9 11 1 11 9 1 13 9 13 4 2
17 11 1 11 11 13 0 10 9 1 9 1 3 13 1 13 4 2
8 10 9 1 1 9 14 13 2
23 9 9 11 11 11 1 13 16 9 13 4 9 1 13 1 1 9 1 3 9 13 4 2
10 15 1 9 13 1 9 13 4 4 2
26 9 1 9 13 14 9 9 1 13 4 7 15 9 1 7 9 2 3 13 2 15 9 1 13 4 2
21 15 1 9 1 9 1 0 9 1 12 9 11 1 13 7 11 1 9 9 13 2
15 9 1 1 9 1 11 1 9 1 0 9 13 4 4 2
17 9 13 1 3 15 0 9 9 13 4 15 9 14 13 4 4 2
33 10 3 11 11 1 0 11 11 11 1 11 1 12 9 1 13 16 11 1 9 13 13 1 1 10 9 9 2 9 1 9 13 2
14 11 3 10 11 1 9 1 10 9 9 13 4 4 2
20 7 9 15 13 16 15 1 9 13 4 7 9 1 9 14 9 1 13 4 2
36 2 9 2 9 1 9 13 1 1 1 9 13 1 9 1 11 1 11 1 11 11 11 11 1 9 11 1 11 1 9 1 3 3 13 4 2
10 11 1 10 9 9 1 1 1 13 2
31 9 1 13 9 1 1 11 9 9 1 1 13 1 11 7 11 9 1 9 1 1 9 13 1 1 11 1 9 13 4 2
24 10 9 1 8 13 1 1 9 1 11 11 11 11 1 12 12 9 1 9 1 9 13 4 2
12 10 12 9 1 11 1 9 1 9 13 4 2
21 9 1 9 9 1 12 12 13 1 1 11 9 1 12 12 9 1 9 0 13 2
21 9 9 1 9 1 9 13 4 1 9 11 1 11 9 1 11 1 13 4 4 2
23 9 13 1 3 11 1 11 9 1 12 0 9 1 9 13 11 1 14 11 0 13 4 2
21 13 4 4 16 11 9 1 14 11 1 9 11 11 1 9 9 1 13 4 4 2
19 11 9 14 9 1 9 9 1 12 12 1 9 1 9 13 13 4 4 2
36 0 0 9 1 1 14 12 12 9 11 11 0 9 1 9 1 9 8 13 1 9 1 12 9 1 9 11 1 9 13 12 12 9 13 4 2
32 0 9 1 12 12 9 3 14 9 1 13 2 15 3 1 0 11 1 9 1 9 1 10 9 9 13 9 1 0 13 4 2
27 10 9 11 1 12 0 9 1 9 1 11 2 11 0 9 1 9 13 2 15 1 12 12 9 0 13 2
25 10 9 11 1 9 9 1 9 1 13 10 9 11 11 1 9 9 0 13 15 9 13 4 4 2
19 9 1 13 14 9 1 0 3 9 1 0 9 1 0 13 1 9 13 2
36 9 1 9 1 3 3 13 1 3 10 9 1 14 9 9 9 1 13 2 15 9 1 9 13 1 3 9 13 1 9 1 9 8 13 4 2
10 9 9 1 14 15 1 13 4 4 2
32 15 9 9 1 11 1 11 1 9 1 0 13 2 14 10 9 15 9 1 12 0 9 1 0 9 1 12 12 9 0 13 2
13 9 1 9 1 1 9 1 9 7 9 0 13 2
19 9 13 4 1 11 1 9 0 13 4 9 1 1 15 9 1 0 13 2
14 13 4 4 16 9 1 9 1 14 11 13 4 4 2
16 9 13 4 1 11 1 9 11 0 9 1 9 1 0 13 2
23 11 11 11 11 1 0 9 13 9 1 9 13 11 11 1 11 9 1 0 13 4 4 2
11 15 9 1 11 13 1 9 13 4 4 2
21 3 1 15 9 13 4 2 7 9 1 11 1 9 13 4 16 15 9 14 13 2
12 3 1 15 9 9 9 9 1 0 13 4 2
22 0 11 11 1 9 9 11 11 1 13 16 11 9 1 9 13 1 9 13 4 4 2
26 0 13 16 11 1 11 9 1 9 9 9 1 11 11 1 9 13 4 2 15 9 1 0 13 4 2
23 9 1 9 1 9 13 1 13 9 1 1 11 1 11 1 9 1 0 13 1 9 13 2
20 0 13 16 11 2 11 11 11 1 9 9 11 11 1 9 13 4 4 4 2
29 10 9 1 12 9 1 13 9 1 1 12 0 9 9 11 11 2 11 11 7 11 11 15 9 1 13 4 4 2
17 15 9 12 9 3 13 4 7 11 7 10 9 1 9 13 4 2
21 9 1 1 2 11 1 15 9 14 13 4 4 4 2 16 15 9 14 13 4 2
21 11 11 9 1 11 11 1 9 10 0 13 2 16 9 1 9 15 1 13 4 2
5 9 9 1 13 2
33 9 1 15 9 13 2 15 11 15 13 4 13 4 4 16 15 9 13 14 14 2 16 15 9 1 15 9 13 7 13 4 4 2
22 11 1 13 1 9 0 13 4 4 2 15 1 11 11 9 1 10 9 0 13 4 2
12 15 11 1 9 7 9 1 3 9 13 4 2
20 3 11 1 9 11 11 11 1 13 16 15 9 1 15 14 0 14 13 4 2
12 15 13 16 10 9 9 13 11 13 4 4 2
19 15 10 9 11 1 1 11 11 11 1 9 1 1 1 15 9 14 13 2
19 9 9 1 1 2 11 1 11 11 1 9 1 11 9 1 9 1 13 2
28 15 15 9 1 11 1 11 11 11 11 11 11 11 1 11 13 1 1 11 11 1 9 9 13 13 4 4 2
15 10 3 0 9 1 1 11 11 1 9 1 15 13 4 2
27 11 11 1 9 1 13 16 11 9 1 11 1 1 9 0 13 4 2 15 9 1 15 0 13 4 4 2
10 11 1 9 9 1 9 13 4 4 2
5 9 1 9 14 13
23 11 9 1 11 1 12 9 0 13 13 16 10 9 1 11 1 0 13 1 9 14 13 2
29 15 1 11 11 11 0 13 1 9 14 15 0 13 4 16 15 11 11 9 9 1 9 1 1 11 1 0 13 2
12 11 9 1 13 16 15 15 9 14 13 4 2
23 10 9 1 11 9 1 13 4 4 16 15 11 1 9 1 0 13 1 1 1 0 13 2
22 9 1 13 4 4 16 16 11 9 13 13 4 16 15 11 9 1 0 13 4 4 2
13 13 9 13 4 16 10 9 10 9 13 4 4 2
29 16 15 9 14 11 13 1 14 13 2 16 15 14 10 9 1 15 13 2 15 11 1 0 9 9 1 13 4 2
15 15 14 10 9 1 13 2 15 15 9 1 0 9 13 2
6 11 7 11 13 1 9
20 0 3 10 9 11 13 2 15 1 11 1 0 9 9 1 9 13 4 4 2
32 15 10 9 1 11 11 11 1 9 1 9 13 2 15 15 13 4 16 15 9 1 13 4 15 9 13 9 1 9 13 4 2
7 15 1 15 9 11 13 2
10 11 1 11 1 9 7 11 11 13 2
13 11 1 9 1 14 11 11 1 9 13 4 4 2
26 10 9 15 1 13 9 11 1 13 13 4 2 7 9 1 9 1 13 4 10 9 9 1 13 4 2
7 15 1 10 9 11 13 2
8 11 11 1 14 15 15 13 2
22 15 9 9 11 11 1 9 1 3 9 13 2 7 15 9 2 9 13 1 9 13 2
10 15 15 11 7 11 13 1 9 13 2
16 12 9 0 11 1 10 9 11 1 15 0 9 14 13 4 2
22 10 9 11 1 11 9 1 1 0 9 1 9 13 2 15 0 0 9 1 9 13 2
29 9 1 1 10 9 1 15 9 1 9 13 4 9 14 0 14 13 2 7 15 0 13 9 13 7 9 13 4 2
13 10 9 11 9 1 9 7 11 11 13 14 13 2
18 10 3 9 9 7 9 1 9 0 9 1 15 1 9 13 4 4 2
40 9 9 1 12 9 1 2 11 11 2 1 13 16 11 1 15 0 9 1 9 13 4 4 4 7 9 2 9 1 15 9 1 9 1 0 13 4 4 4 2
21 3 11 1 11 1 9 9 1 9 13 1 9 1 12 9 1 0 13 4 4 2
25 11 11 1 3 0 9 9 11 11 11 1 9 1 11 1 12 9 1 0 9 1 9 13 4 2
18 10 0 9 1 0 9 0 13 4 7 15 9 1 15 9 14 13 2
15 9 1 9 2 9 1 9 15 0 9 1 13 4 4 2
16 11 1 11 7 11 1 14 9 1 0 13 15 0 9 13 2
10 0 9 1 11 11 11 1 9 13 2
15 0 9 1 1 12 0 9 1 9 11 9 13 4 4 2
19 11 1 15 0 9 1 13 4 16 9 1 9 9 7 11 11 1 13 2
22 16 15 15 0 9 1 9 0 14 13 4 7 10 9 11 11 1 0 13 4 4 2
14 11 1 11 11 11 1 9 1 0 13 1 9 13 2
13 9 1 9 1 11 1 9 1 9 13 4 4 2
20 11 11 1 15 9 0 13 4 11 1 12 9 1 0 9 1 9 13 4 2
7 11 11 1 10 9 13 2
19 11 1 9 1 1 10 9 1 14 12 9 1 9 1 9 13 4 4 2
22 11 11 11 11 11 11 1 9 0 13 4 13 16 15 9 1 9 1 10 0 13 2
12 9 1 12 0 9 7 12 9 13 4 4 2
14 15 15 0 9 9 7 9 1 9 1 1 9 13 2
22 15 10 9 1 9 1 1 0 9 7 9 7 9 1 0 0 9 1 1 9 13 2
22 11 11 11 11 1 13 16 15 9 1 9 2 9 2 9 7 0 9 1 9 13 2
20 15 9 1 15 12 10 0 9 13 4 4 15 0 9 1 15 9 13 4 2
27 11 11 11 1 15 9 9 1 13 16 15 0 9 1 9 13 15 0 9 1 1 11 11 1 9 13 2
18 15 0 12 9 1 10 9 9 13 4 4 15 9 1 0 9 13 2
20 15 10 9 11 11 1 9 1 9 13 2 15 15 9 1 9 1 13 4 2
16 15 9 1 9 1 13 10 9 1 0 9 1 14 9 13 2
7 15 0 9 1 0 13 2
18 11 9 11 11 1 14 9 1 9 1 9 0 9 1 9 13 4 2
8 9 9 1 9 10 9 13 2
21 11 0 11 11 11 1 9 9 9 11 9 1 0 9 1 9 13 11 11 13 2
15 15 11 9 1 0 0 9 1 1 9 1 10 9 13 2
9 15 9 1 9 1 0 9 13 2
15 9 1 13 16 0 9 15 9 9 1 1 13 4 4 2
16 10 3 11 11 1 9 1 0 9 1 1 9 13 4 4 2
11 15 0 9 3 0 9 1 13 4 4 2
12 15 9 1 9 2 9 1 9 13 4 4 2
22 0 9 1 1 9 1 13 0 9 9 2 9 2 9 2 0 9 7 14 9 13 2
17 15 11 1 11 11 11 11 2 11 11 11 7 15 9 0 13 2
13 10 9 1 9 1 9 13 15 1 0 13 4 2
32 11 11 1 11 11 11 1 9 11 1 10 0 9 0 13 4 15 9 1 15 14 9 13 4 7 13 1 15 13 4 4 2
15 11 11 9 1 10 9 11 1 11 1 9 1 0 13 2
30 9 1 1 13 1 0 9 1 1 14 0 9 13 4 9 1 0 13 1 9 14 0 10 9 1 10 13 4 4 2
30 7 11 11 11 11 11 11 2 11 2 1 9 1 13 13 16 11 11 1 1 10 9 1 9 13 10 0 13 4 2
28 15 1 15 3 0 13 4 16 11 2 11 1 9 11 11 1 13 4 11 11 11 11 11 1 9 8 13 2
15 9 13 1 10 0 9 1 1 1 10 9 15 1 13 2
16 10 9 1 9 1 15 9 1 9 1 9 0 13 4 4 2
42 11 1 0 9 11 11 11 1 11 1 9 1 13 9 1 13 16 15 9 1 1 14 14 13 4 16 12 0 9 13 4 16 15 15 1 1 10 9 13 4 4 2
10 7 14 13 16 9 1 9 13 4 2
28 11 13 4 16 3 10 13 16 14 12 9 9 1 14 9 1 9 13 4 0 13 1 9 0 13 14 4 2
17 16 15 9 13 4 4 16 15 15 9 1 9 1 3 14 13 2
20 11 1 10 9 1 0 9 1 11 1 9 9 1 9 1 1 0 13 4 2
16 15 1 9 13 11 1 0 10 9 1 1 10 9 13 4 2
27 11 1 9 9 1 9 1 9 13 1 12 9 13 4 16 9 9 1 1 10 9 15 10 0 14 13 2
24 9 1 9 1 13 4 9 9 1 9 1 13 4 9 9 9 16 9 1 9 13 4 4 2
26 11 9 13 4 16 11 11 11 1 1 9 13 1 1 1 1 0 9 0 13 9 1 1 0 13 2
26 11 1 9 11 11 11 7 11 11 11 1 11 11 11 1 11 11 1 10 9 1 1 9 13 4 2
14 0 9 2 11 11 11 2 1 10 0 9 13 4 2
48 9 1 1 15 0 9 9 11 1 11 1 11 0 9 2 11 11 11 11 2 1 9 13 15 15 15 11 9 1 0 9 1 9 9 13 1 9 7 15 9 2 9 1 1 1 9 13 2
22 15 1 11 7 11 2 11 2 11 1 10 0 9 1 13 2 9 1 14 9 13 2
32 9 1 1 11 11 11 11 1 0 9 7 11 11 11 1 9 11 1 11 1 9 1 11 11 2 11 1 0 13 4 4 2
29 11 1 0 9 1 14 15 9 1 9 1 1 9 13 4 2 7 13 9 1 15 9 9 1 9 13 4 4 2
31 11 11 11 11 1 1 1 13 10 9 1 13 4 16 11 2 11 7 0 9 1 11 11 11 1 10 9 1 9 13 2
14 11 0 11 11 1 9 1 9 1 9 1 0 13 2
19 9 1 0 13 4 1 3 1 15 9 11 2 11 2 11 13 4 4 2
38 9 1 13 4 16 11 11 1 11 11 1 9 9 1 13 4 7 11 1 11 1 11 2 11 1 0 9 1 1 9 13 1 1 14 13 4 4 2
45 2 11 11 11 2 1 13 16 11 1 10 0 9 1 1 1 13 4 4 4 2 15 13 13 16 11 1 9 13 4 7 15 14 15 1 14 13 4 10 0 9 1 13 4 2
11 15 15 11 7 0 9 1 9 13 4 2
31 0 11 11 11 7 11 1 11 11 11 1 1 11 2 11 11 1 14 12 9 1 0 9 13 1 9 0 13 4 4 2
21 13 4 4 16 12 9 1 0 9 10 0 9 1 9 0 13 1 1 3 13 2
41 9 1 1 9 1 1 1 0 9 13 1 1 11 9 1 0 11 1 11 1 0 9 11 11 11 11 1 9 7 0 9 9 9 1 9 11 11 1 9 13 2
15 16 10 9 1 1 9 7 9 1 9 15 14 13 4 2
14 7 9 1 13 13 16 10 9 11 1 13 4 4 2
25 11 9 1 12 0 9 1 13 16 11 7 11 1 1 0 9 1 0 9 0 14 13 4 4 2
18 11 11 9 11 11 1 1 2 9 0 0 9 1 14 13 13 4 2
21 11 11 1 10 9 1 15 9 14 13 7 10 9 1 14 9 13 4 4 4 2
32 9 1 13 16 3 0 11 9 1 14 11 1 1 9 9 1 9 1 9 13 4 7 9 9 10 9 1 3 13 4 4 2
21 9 1 15 14 13 4 16 11 11 11 11 11 1 9 1 14 9 13 4 4 2
15 16 15 10 9 1 11 9 1 15 0 9 14 13 4 2
26 11 9 1 1 13 4 9 9 1 9 0 13 4 10 9 1 13 16 9 0 9 1 13 4 4 2
18 12 9 1 1 9 0 13 7 3 14 15 0 9 3 13 4 4 2
24 12 12 0 9 9 13 1 1 11 13 4 0 9 9 1 9 9 1 1 1 13 4 4 2
43 11 11 11 11 2 11 2 1 11 1 11 11 11 1 1 1 9 1 9 14 13 4 1 3 11 11 14 11 11 1 1 13 1 10 9 1 9 0 13 1 9 13 2
22 12 0 9 9 1 10 9 15 12 9 1 1 1 9 1 9 13 1 3 13 4 2
31 11 1 9 9 11 11 1 9 1 9 2 9 7 9 0 13 1 0 9 1 15 13 9 1 1 9 1 10 9 13 2
32 15 13 16 9 1 9 13 1 11 11 11 2 11 2 1 9 7 15 9 9 1 13 9 1 1 9 1 10 9 13 4 2
22 9 1 0 13 16 10 9 12 9 1 1 9 1 9 13 1 0 13 4 4 4 2
11 9 1 9 11 1 9 11 11 1 13 2
15 9 1 1 1 9 11 11 11 9 1 0 14 13 4 2
19 0 13 16 11 1 11 11 1 0 9 1 1 11 1 0 13 4 4 2
36 15 1 11 1 9 1 9 9 9 1 0 9 11 11 1 0 9 11 11 1 13 11 11 11 1 9 1 0 13 1 9 14 13 4 4 2
12 16 11 1 0 9 1 3 9 0 13 4 2
15 15 9 1 13 4 9 1 9 1 9 14 13 4 4 2
18 9 10 0 9 1 1 12 9 1 9 13 1 9 3 14 9 13 2
31 15 1 1 9 1 13 16 9 11 11 11 11 1 12 9 7 11 11 11 1 12 9 9 13 1 9 3 13 4 4 2
27 15 1 14 12 0 9 15 9 13 4 1 9 13 15 13 11 11 2 11 11 11 11 7 11 11 11 2
21 10 9 1 9 13 4 1 9 1 3 14 0 9 1 9 9 1 1 13 4 2
14 0 9 1 9 13 13 4 9 9 9 9 1 13 2
28 9 1 1 12 9 9 1 9 0 9 1 9 1 13 4 7 0 9 1 0 9 1 9 1 9 13 4 2
21 11 11 1 9 1 1 10 9 1 9 1 9 15 14 12 9 14 13 4 4 2
12 9 1 10 9 1 9 10 9 1 13 4 2
12 7 11 11 11 1 9 1 9 12 9 13 2
6 15 9 12 12 13 2
15 11 11 1 10 9 1 12 9 9 13 1 9 13 4 2
21 11 1 12 9 9 13 1 3 10 9 1 9 1 9 12 1 13 12 13 4 2
17 10 9 1 12 9 9 13 1 9 1 12 12 1 9 0 13 2
25 9 11 2 11 1 1 9 1 0 9 1 9 1 13 12 1 12 12 9 13 1 9 13 4 2
26 15 1 14 11 11 1 0 12 9 1 0 9 1 9 13 12 1 12 12 9 13 1 9 13 4 2
45 12 0 9 1 9 13 15 9 13 4 1 9 1 11 1 11 7 11 9 1 11 1 9 1 9 1 0 13 4 0 11 11 1 9 1 9 13 4 1 9 1 0 13 4 2
34 9 11 11 7 9 11 11 11 1 9 1 15 12 9 1 9 1 13 16 15 15 15 9 9 14 13 16 9 1 1 9 13 4 2
24 9 0 13 4 4 16 9 1 9 7 0 9 1 9 1 1 9 13 1 3 15 9 13 2
31 9 11 11 0 0 9 1 13 1 12 0 9 11 11 14 11 11 11 11 1 15 9 11 11 1 9 13 1 1 13 2
8 11 1 9 9 1 13 4 2
14 13 1 3 11 10 9 1 15 9 11 1 13 13 2
20 9 9 1 11 1 9 14 13 1 9 1 1 15 13 2 7 15 14 13 2
15 3 1 11 1 9 0 11 1 9 1 0 9 1 13 2
14 9 1 9 9 1 0 13 7 15 9 1 9 13 2
6 9 1 14 9 13 2
19 9 1 14 12 9 11 11 1 13 16 15 9 1 11 1 1 13 4 2
14 9 1 11 1 9 1 9 13 2 7 15 14 13 2
16 3 1 9 1 9 11 11 1 11 1 9 1 1 0 13 2
23 9 9 1 13 16 9 1 1 9 13 4 7 10 9 13 4 1 1 15 9 13 4 2
22 11 1 9 9 9 1 9 0 13 4 1 11 1 11 11 11 1 9 1 9 13 2
11 9 1 1 11 1 9 1 9 0 13 2
20 9 1 11 1 9 1 13 16 9 1 15 9 1 0 14 9 13 4 4 2
14 0 9 1 14 13 1 15 1 0 9 13 4 4 2
20 15 1 15 9 9 1 1 13 7 10 9 1 9 1 9 13 0 14 13 2
25 11 9 1 9 1 13 16 9 1 9 11 11 0 9 13 7 15 9 1 9 1 1 13 4 2
7 15 1 9 0 13 4 2
28 12 9 1 9 13 1 3 9 1 9 1 0 9 1 9 1 0 13 4 9 1 9 13 4 1 9 13 2
28 11 11 11 11 1 1 11 11 11 1 0 9 1 9 0 13 15 1 11 2 11 1 9 1 9 13 4 2
14 11 1 9 9 1 9 1 15 9 14 13 4 4 2
38 9 1 11 11 1 9 1 9 1 11 1 13 16 10 9 1 0 12 9 1 9 1 9 13 4 7 11 2 11 1 1 15 9 0 13 4 4 2
28 9 1 9 1 9 10 13 1 1 9 1 9 1 9 13 4 7 15 9 13 4 4 15 9 13 4 4 2
28 15 13 4 1 16 15 11 1 0 9 1 9 9 13 4 11 1 13 16 15 14 9 15 15 9 14 13 2
15 7 15 9 1 1 11 1 9 1 9 13 4 4 4 2
26 11 11 11 11 1 13 16 9 1 9 1 0 9 1 13 1 9 13 1 9 1 15 9 14 13 2
37 15 13 16 0 12 9 1 1 14 12 12 9 1 9 1 9 13 4 7 9 13 1 0 9 15 13 15 15 9 1 12 9 0 13 4 4 2
35 9 1 9 1 1 11 11 11 11 1 13 4 9 1 9 1 11 1 13 16 9 1 9 1 13 1 9 3 0 13 7 9 0 13 2
7 9 1 9 14 10 13 2
17 10 9 1 9 13 1 1 9 1 1 9 1 15 9 14 13 2
17 15 15 0 9 1 13 1 9 13 4 9 1 1 0 14 13 2
29 15 13 16 11 1 13 1 15 9 1 9 13 4 16 15 12 9 9 1 13 15 1 0 9 0 13 4 4 2
29 11 1 11 11 1 9 1 9 1 11 1 13 16 9 10 9 1 9 1 1 11 11 11 1 9 1 9 13 2
23 15 13 16 9 1 9 1 9 1 3 13 1 1 14 9 0 9 9 9 13 4 4 2
40 11 1 9 13 16 15 11 11 11 11 1 9 7 11 1 0 9 11 11 1 11 1 9 1 1 9 13 16 15 1 0 9 1 9 1 9 13 4 4 2
20 11 9 1 1 9 9 11 1 9 9 1 1 11 11 1 9 1 9 13 2
14 0 13 16 11 1 11 1 9 13 9 9 13 4 2
8 15 11 9 1 13 4 4 2
15 9 1 1 11 1 9 13 0 9 1 9 1 0 13 2
25 15 1 1 9 1 9 13 4 16 11 1 11 11 11 1 9 1 11 1 0 9 0 13 4 2
15 10 9 1 1 15 11 11 1 1 11 1 13 4 4 2
11 15 0 9 1 9 13 16 15 9 13 2
17 11 1 11 11 11 7 11 11 1 0 9 1 1 9 13 4 2
31 9 1 13 16 11 1 11 11 1 9 1 0 13 4 13 4 16 15 1 11 1 11 9 1 13 15 9 14 13 4 2
10 7 10 9 1 11 11 1 9 13 2
23 0 9 1 1 11 1 12 9 1 9 13 1 3 11 1 11 1 9 1 13 4 4 2
16 9 1 2 15 11 0 13 4 1 9 1 15 9 13 4 2
9 15 9 15 11 11 1 0 13 2
36 9 9 9 11 11 1 13 16 11 11 1 9 1 1 9 9 1 0 13 0 9 1 0 9 7 2 9 9 9 2 1 1 3 0 13 2
21 15 0 13 16 9 9 1 15 9 1 10 9 1 9 1 0 9 13 4 4 2
38 0 9 2 11 11 11 2 1 13 4 12 9 1 15 13 16 11 1 11 11 9 1 9 1 12 9 1 0 9 1 0 13 1 9 13 4 4 2
42 9 9 9 7 9 9 9 1 9 1 9 1 9 1 15 9 13 4 13 16 9 13 4 4 4 7 15 9 1 9 1 9 1 15 9 10 9 1 0 13 4 2
18 15 13 16 9 2 11 11 11 2 15 9 9 9 1 0 9 13 2
16 9 9 1 13 16 15 11 11 11 1 9 9 13 4 4 2
15 15 1 9 13 1 9 13 1 9 1 9 13 4 4 2
29 16 2 15 13 16 0 9 10 9 1 0 9 0 13 7 15 9 13 16 3 14 10 9 1 9 9 13 4 2
29 9 9 1 13 16 0 9 9 1 9 1 15 9 13 4 4 7 0 9 1 12 9 9 1 0 9 1 13 2
32 15 13 16 15 12 0 9 7 9 2 11 11 11 1 11 11 2 2 2 11 11 11 11 11 2 7 11 11 11 0 13 2
25 11 1 12 9 0 11 9 1 13 9 7 9 1 0 9 1 9 1 1 0 9 1 13 4 2
19 15 13 13 16 15 10 9 1 11 7 11 1 1 0 9 10 0 13 2
15 15 15 13 13 4 16 11 9 1 1 3 0 15 13 2
13 0 9 11 7 11 11 1 11 1 1 0 13 2
14 11 11 1 10 9 13 15 1 11 1 9 13 4 2
19 10 9 12 9 7 12 9 1 0 13 12 9 1 11 9 1 13 4 2
12 15 9 13 11 1 9 7 9 1 3 13 2
11 0 9 1 11 1 0 9 1 0 13 2
31 15 11 1 1 0 13 1 3 9 1 9 13 4 13 16 11 1 13 0 0 9 1 15 9 9 1 10 0 13 4 2
8 0 11 9 11 1 9 13 2
17 15 0 13 16 9 10 9 1 9 13 4 15 1 0 13 4 2
28 11 1 11 1 9 9 7 9 13 1 10 12 9 15 10 0 9 1 1 12 9 1 13 15 9 13 13 2
29 11 1 0 11 1 13 16 15 15 15 0 11 9 1 1 1 9 13 4 2 15 15 9 9 1 13 4 4 2
14 15 15 15 9 1 10 9 7 9 1 13 13 4 2
22 15 10 9 1 1 10 9 11 2 11 2 11 2 11 2 11 7 11 1 13 13 2
9 10 10 9 1 0 9 13 4 2
18 11 1 13 16 11 1 15 9 1 13 1 15 9 0 13 4 4 2
41 11 11 11 11 1 11 1 9 1 0 13 16 11 11 11 1 11 11 11 11 11 11 1 1 1 0 0 9 1 13 1 1 9 9 1 10 0 9 0 13 2
27 11 1 9 1 9 1 13 11 7 9 1 9 9 1 9 1 13 16 9 9 1 0 9 9 13 13 2
24 16 15 15 13 1 0 13 4 2 16 15 9 9 1 0 9 1 0 9 13 1 9 13 2
14 15 1 14 0 9 1 1 14 9 13 4 4 4 2
18 15 13 16 0 9 1 10 9 9 13 2 15 10 9 7 9 13 2
25 9 1 9 1 9 1 13 4 15 12 10 9 13 4 2 15 15 9 7 9 1 10 13 4 2
11 12 10 9 15 15 1 14 9 14 13 2
20 11 1 12 0 12 11 0 9 9 1 9 1 0 9 13 1 9 1 13 2
16 11 0 11 1 11 9 1 11 11 9 1 9 13 4 4 2
8 11 3 10 9 1 9 13 2
15 11 1 13 16 15 11 1 9 1 10 9 1 9 13 2
16 15 1 15 3 0 9 13 2 7 15 11 1 0 9 13 2
22 15 11 0 13 2 7 15 13 4 16 10 9 1 11 7 11 9 1 9 0 13 2
15 15 9 1 11 11 1 9 13 1 1 9 13 4 4 2
15 15 13 16 10 0 9 1 15 9 13 1 1 0 13 2
27 11 11 9 1 11 9 1 13 1 11 1 13 16 10 9 1 9 14 15 10 0 9 1 13 13 4 2
20 15 15 9 13 1 9 13 4 15 10 9 1 9 1 9 1 9 13 4 2
14 11 1 11 0 13 1 9 9 1 15 1 14 13 2
24 11 1 0 9 1 9 13 1 11 1 9 1 14 1 9 13 4 4 16 15 9 0 13 2
14 15 13 16 15 9 1 3 9 2 9 14 13 4 2
17 11 1 15 9 13 4 2 7 15 1 15 11 0 13 4 4 2
11 15 11 11 11 1 1 9 13 4 4 2
20 11 1 0 9 9 11 11 11 15 9 1 1 9 1 9 1 13 4 4 2
20 11 1 15 12 12 0 9 9 1 9 1 9 1 12 12 9 9 13 4 2
47 9 1 0 13 4 12 9 1 13 4 4 16 11 1 10 9 9 1 11 2 11 1 11 2 11 1 9 1 11 11 1 15 14 0 9 1 9 9 1 1 1 3 10 9 13 4 2
24 0 13 16 11 1 9 9 1 13 0 2 0 9 1 9 9 11 11 1 9 1 13 4 2
9 11 11 11 11 11 1 9 13 2
19 10 9 12 9 1 11 11 2 11 2 11 1 9 9 1 1 12 13 2
15 11 1 13 4 9 1 9 1 10 9 1 0 13 4 2
20 11 9 1 1 11 1 11 2 11 2 11 11 1 9 14 12 9 9 13 2
30 15 15 1 1 11 11 1 9 11 11 11 1 13 4 15 15 13 16 15 10 9 1 1 1 0 9 13 4 4 2
17 2 11 2 9 1 1 15 10 9 1 9 1 10 9 13 4 2
20 15 1 14 15 14 9 9 1 13 1 9 9 1 3 10 9 9 13 4 2
16 11 2 11 1 11 2 11 1 1 15 12 9 9 9 13 2
11 15 1 9 1 12 12 9 9 13 4 2
19 11 11 11 11 11 15 9 9 1 9 13 1 9 1 11 1 1 13 2
24 15 14 11 2 11 1 12 0 9 13 4 2 7 15 10 9 1 12 12 9 14 9 13 2
12 11 1 11 9 1 12 12 9 9 13 4 2
21 11 11 1 9 13 1 9 9 1 0 9 1 13 4 9 1 9 13 4 4 2
15 9 1 9 1 9 13 11 1 0 9 1 13 4 4 2
12 15 10 14 10 9 9 1 1 9 13 4 2
15 10 9 1 9 11 1 11 11 1 1 1 13 4 4 2
32 0 9 9 1 9 13 1 9 9 1 0 9 13 4 1 9 1 1 1 12 9 1 0 9 7 9 1 1 9 13 4 2
19 15 1 9 1 0 9 1 13 9 1 9 1 13 1 9 13 4 4 2
17 11 1 11 1 0 9 9 1 12 1 10 9 13 4 4 4 2
23 0 9 9 7 9 1 13 13 16 11 11 11 11 15 9 1 0 13 1 13 4 4 2
19 3 14 11 1 9 9 14 13 2 7 10 9 9 14 15 9 1 13 2
16 9 1 13 13 16 9 9 1 9 13 1 9 13 4 4 2
20 3 14 11 1 15 9 9 14 13 2 7 9 9 14 10 9 13 4 4 2
10 15 9 1 14 9 14 13 4 4 2
15 9 9 0 7 0 0 9 1 9 1 9 13 4 4 2
28 9 2 9 2 9 9 11 11 1 0 9 1 9 2 11 2 11 11 2 1 9 9 1 1 9 13 4 2
11 9 9 1 9 1 10 9 1 9 13 2
17 15 10 9 11 11 11 1 13 4 1 9 1 9 1 0 13 2
18 10 9 9 9 11 11 1 0 12 9 1 14 9 1 9 13 4 2
17 10 9 1 9 1 13 4 1 9 1 9 9 1 9 13 4 2
22 0 2 0 9 9 11 11 1 9 2 11 11 11 2 1 14 9 9 1 9 13 2
10 15 15 9 9 1 13 4 4 4 2
42 11 1 11 11 11 11 1 9 2 11 11 11 2 1 3 9 1 13 16 10 9 1 0 9 13 4 4 2 10 9 1 0 9 0 9 2 9 9 1 9 13 2
15 15 13 16 9 9 9 9 1 9 1 0 13 4 4 2
21 11 1 15 9 1 12 9 1 9 13 1 13 4 4 2 15 15 9 13 4 2
21 0 10 9 9 1 13 13 16 9 9 1 14 9 9 13 1 9 13 4 4 2
12 9 1 9 1 9 13 15 9 13 4 4 2
19 0 9 1 9 2 9 9 1 12 0 9 1 9 1 9 13 4 4 2
36 11 11 11 11 11 11 1 11 1 9 1 12 0 9 1 13 16 9 1 12 9 12 0 9 9 9 1 9 1 9 1 9 1 13 13 2
23 10 9 1 0 9 1 0 9 1 0 2 0 7 0 9 1 9 1 9 1 9 13 2
25 11 11 11 11 11 1 13 16 11 2 11 2 11 7 11 11 9 3 0 9 1 13 4 4 2
21 9 1 9 13 1 3 9 1 1 1 9 1 9 1 1 9 0 13 4 4 2
22 15 13 16 3 0 9 1 9 1 1 11 1 9 0 9 1 1 1 13 4 4 2
31 11 11 11 11 11 1 13 16 9 0 9 1 9 0 13 1 9 7 9 1 0 7 0 0 9 2 9 13 4 4 2
28 15 13 16 16 10 9 0 9 1 0 13 1 9 13 4 4 2 16 9 15 1 0 9 13 1 9 13 2
35 12 0 9 1 9 1 11 1 13 16 9 1 0 9 1 12 0 9 0 13 7 9 1 9 1 0 0 0 9 0 13 1 9 13 2
36 15 13 16 10 9 1 9 1 13 4 12 9 7 12 0 0 9 1 10 13 4 0 9 1 9 1 1 1 12 9 9 0 13 4 4 2
32 11 11 11 1 9 11 11 1 0 10 9 1 0 13 4 4 15 0 11 11 11 11 1 9 13 4 1 9 13 4 4 2
28 9 1 13 16 11 9 1 1 1 9 1 13 4 9 1 9 1 11 1 9 13 4 1 15 9 14 13 2
18 16 15 15 9 13 16 11 11 2 11 1 9 1 9 15 1 13 2
29 11 1 9 0 13 4 9 1 13 16 0 11 11 11 11 1 11 1 13 9 1 9 1 1 13 4 4 4 2
42 0 13 16 11 1 9 1 1 9 1 13 4 16 15 11 1 10 9 13 15 9 1 1 0 9 1 1 9 13 4 4 7 9 1 9 1 9 14 13 4 4 2
16 9 1 11 1 14 9 13 4 1 11 1 9 1 13 4 2
14 9 1 15 11 11 1 9 13 15 1 15 9 13 2
10 15 0 9 1 13 1 1 13 4 2
19 9 13 1 3 11 1 10 9 1 9 13 16 9 1 0 9 15 13 2
11 7 2 15 15 13 16 9 15 1 13 2
52 11 1 0 13 16 15 10 9 1 1 15 14 15 9 0 14 13 2 16 11 11 2 11 1 15 14 12 9 0 13 4 15 15 9 1 9 13 1 9 13 4 4 16 10 9 11 11 1 0 13 4 2
29 11 1 3 13 16 15 11 11 2 11 2 11 11 2 11 7 11 11 2 11 1 11 11 1 9 0 13 4 2
13 15 9 1 1 12 9 1 9 14 0 13 4 2
34 15 10 14 9 13 16 11 11 11 1 9 1 11 11 2 11 1 11 9 1 0 13 4 9 1 1 1 14 15 15 9 14 13 2
14 7 2 15 15 9 13 16 9 1 9 15 1 13 2
27 9 1 1 11 1 0 9 14 9 13 4 4 7 9 11 11 1 13 4 10 9 1 15 9 14 13 2
19 12 3 0 9 1 11 11 1 9 1 9 9 1 11 1 9 13 4 2
18 10 9 11 11 1 0 13 7 15 1 9 1 0 0 9 9 13 2
22 9 1 0 9 1 12 9 1 0 7 9 9 1 1 9 9 1 14 9 13 4 2
38 9 1 13 9 1 0 9 7 0 9 1 9 13 1 9 0 13 1 9 13 1 12 9 1 9 1 9 9 1 9 13 4 15 9 0 13 4 2
29 0 9 7 9 1 0 9 11 11 1 11 9 1 9 9 9 1 13 4 9 9 1 11 11 1 9 13 4 2
40 11 1 9 11 11 7 9 11 11 11 1 9 1 11 11 1 10 9 1 13 4 15 13 4 4 16 9 9 1 9 13 1 9 15 0 9 14 0 13 2
39 9 1 10 9 13 4 16 9 9 9 1 1 1 9 1 9 13 4 4 7 9 1 1 9 9 9 1 14 9 13 4 2 15 0 9 0 13 4 2
33 9 1 13 16 16 9 9 1 0 14 13 4 16 15 0 14 13 4 7 16 15 0 13 4 4 16 15 1 0 14 13 4 2
32 9 1 0 9 1 0 13 11 1 15 9 1 13 16 13 9 1 9 9 1 0 9 1 9 1 0 9 1 9 13 4 2
30 11 9 1 9 9 1 9 1 11 1 9 13 3 14 9 9 13 1 1 9 9 13 13 9 1 9 13 4 4 2
10 0 9 11 1 14 15 9 13 4 2
27 11 1 13 16 9 9 1 1 10 9 1 9 13 1 9 0 13 14 0 9 1 0 9 1 9 13 2
23 9 1 9 13 16 9 1 0 9 1 9 0 9 1 9 7 9 9 9 1 9 13 2
19 0 13 16 9 1 0 9 1 1 10 14 10 12 0 9 14 0 13 2
21 10 9 15 14 9 1 9 14 13 7 15 12 9 1 1 10 9 0 13 4 2
17 9 1 10 12 9 1 1 12 12 10 0 9 8 13 4 4 2
19 15 11 1 11 11 11 11 11 1 9 1 0 2 0 9 13 4 4 2
31 11 11 11 1 9 11 11 1 2 11 1 0 2 0 9 13 4 4 2 9 9 1 1 11 11 1 9 13 4 4 2
22 10 9 1 9 1 1 11 1 15 11 1 11 1 13 4 2 15 11 0 13 4 2
12 11 14 13 16 11 1 12 9 9 13 4 2
29 9 1 1 11 1 10 9 3 13 4 4 4 16 11 3 14 11 1 1 10 9 0 13 4 16 15 13 4 2
9 11 1 9 11 1 9 14 13 2
10 11 1 11 1 9 14 9 14 13 2
22 11 1 13 4 16 11 15 0 9 1 13 9 1 9 13 1 15 1 0 13 4 2
25 11 11 11 1 3 0 11 13 4 1 11 1 11 11 11 11 7 11 11 11 1 15 9 13 2
17 11 1 9 0 13 16 13 1 9 1 11 7 0 9 10 13 2
19 15 1 14 15 13 16 9 7 9 1 13 1 15 9 1 9 13 4 2
10 15 11 1 11 13 1 9 14 13 2
36 9 9 1 11 11 11 11 11 11 1 9 7 11 1 9 1 1 1 13 4 16 15 9 13 16 15 0 9 1 15 0 9 10 0 13 2
22 11 1 12 9 1 1 9 1 10 0 9 13 1 1 0 9 13 1 14 9 13 2
27 15 1 14 15 0 11 1 11 13 1 9 13 7 13 16 15 0 9 1 13 1 9 1 9 0 13 2
24 11 11 1 11 9 1 12 9 1 12 9 1 9 13 4 13 1 9 3 0 13 4 4 2
21 9 9 1 11 1 13 4 16 15 9 1 9 13 4 13 1 15 9 14 13 2
16 10 9 1 9 1 12 9 1 9 1 1 11 11 13 4 2
33 11 11 11 1 9 11 11 11 1 11 1 10 9 1 9 13 16 11 11 1 11 11 13 9 1 9 13 4 13 1 13 4 2
13 15 13 16 11 1 9 13 15 9 14 13 4 2
43 9 1 9 9 11 11 1 13 16 10 9 1 11 1 13 4 16 15 9 1 1 9 13 4 13 16 0 13 7 16 11 9 14 13 13 4 16 15 15 9 14 13 2
28 11 1 11 11 1 11 11 11 11 1 13 4 16 9 9 13 4 16 9 9 1 7 0 9 1 9 13 2
21 16 11 1 9 1 9 1 15 13 13 16 10 9 1 15 9 14 13 4 4 2
45 9 9 1 0 9 13 1 9 13 1 12 9 2 11 11 2 11 11 1 10 0 9 1 9 1 9 1 11 7 11 1 9 1 9 1 1 15 9 3 13 1 0 13 4 2
8 11 11 1 11 14 0 13 2
28 11 2 11 2 11 7 11 1 10 11 11 1 0 9 9 7 9 9 1 1 10 9 1 9 0 13 4 2
17 9 1 15 1 11 11 11 11 1 9 1 9 1 9 0 13 2
17 10 9 1 9 13 16 11 1 0 9 1 10 9 0 13 4 2
33 11 11 9 7 11 7 11 1 9 1 11 11 11 2 11 2 1 3 11 1 0 12 9 1 15 1 9 3 14 13 4 4 2
16 11 9 9 1 0 9 1 9 1 9 1 9 13 4 4 2
15 9 11 11 11 1 9 11 11 1 9 1 13 4 4 2
22 15 11 11 9 1 13 16 11 1 15 0 9 14 13 2 15 1 9 13 4 4 2
28 9 1 1 11 1 9 1 13 16 15 12 9 1 11 11 1 1 15 9 9 1 14 13 1 9 13 4 2
34 15 13 16 0 11 1 11 11 1 9 9 1 0 9 1 1 0 13 4 4 15 1 0 9 9 1 15 1 15 9 13 13 4 2
38 11 11 1 9 1 13 16 11 1 9 1 1 15 9 11 11 1 9 1 1 14 13 4 4 2 7 15 15 15 0 13 1 9 14 13 4 4 2
8 11 1 11 1 9 0 13 2
12 11 1 9 1 1 15 9 1 0 14 13 2
24 11 1 13 2 15 13 16 12 9 1 9 1 1 9 1 13 1 1 9 2 9 0 13 2
28 11 11 11 1 0 2 0 9 9 11 11 1 9 1 0 0 9 1 9 1 1 12 9 1 9 13 4 2
25 9 9 1 0 9 1 13 1 0 9 1 9 13 7 12 9 1 1 9 1 15 9 13 4 2
13 0 9 1 12 9 1 9 1 9 13 4 4 2
11 11 11 9 1 9 9 1 9 14 13 2
9 9 11 11 11 1 1 9 13 2
35 11 2 11 11 11 9 1 9 9 1 9 1 0 9 9 13 2 0 9 1 9 13 2 11 11 7 0 9 14 10 0 9 13 4 2
11 15 15 9 1 9 13 0 13 4 4 2
10 9 1 10 9 1 9 15 13 4 2
41 0 9 1 9 1 11 1 9 1 1 9 11 11 11 1 10 9 9 1 0 13 4 15 9 9 1 9 11 11 1 15 9 1 9 13 4 15 10 9 13 2
16 7 9 11 11 11 1 3 2 3 13 1 15 9 13 4 2
13 11 1 13 16 15 9 9 1 11 1 9 13 2
18 11 1 9 1 9 1 12 9 1 1 9 9 9 13 13 4 4 2
27 0 13 16 11 11 1 11 11 1 9 2 11 11 2 1 9 9 1 13 9 9 1 9 1 9 13 2
9 9 1 14 12 9 13 4 4 2
23 11 11 11 11 11 2 11 2 1 3 0 9 9 1 9 9 14 13 1 9 13 4 2
26 15 1 11 1 9 1 11 2 11 1 1 9 1 0 9 9 12 9 14 9 13 1 9 13 4 2
15 7 9 7 9 1 9 9 1 9 1 9 13 4 4 2
21 0 9 1 1 11 1 11 9 1 1 9 1 0 9 9 1 9 13 4 4 2
37 15 1 9 1 0 9 9 0 12 9 1 1 14 12 9 14 9 13 4 4 7 9 7 9 1 0 9 9 1 0 9 1 9 13 4 4 2
37 9 1 1 11 1 13 13 16 9 1 9 0 13 4 1 11 7 11 1 9 1 9 0 9 1 1 0 13 7 15 9 1 1 0 0 13 2
27 0 13 16 10 12 9 1 9 1 9 13 1 1 0 9 1 0 9 1 1 9 10 3 13 4 4 2
44 11 11 1 0 9 9 2 11 2 1 13 4 9 1 0 13 1 1 0 9 1 11 2 11 1 9 1 11 11 1 12 12 12 9 1 0 0 9 13 1 9 13 4 2
24 16 2 11 11 2 9 1 9 1 9 1 9 13 1 3 14 9 13 4 1 9 1 13 2
24 7 2 9 1 9 1 1 11 11 11 11 0 9 1 0 9 13 4 1 9 1 14 13 2
21 11 1 3 10 9 10 9 1 13 16 9 1 9 13 1 0 9 1 9 13 2
24 9 1 9 1 13 4 11 11 11 1 9 1 9 13 1 0 9 1 14 9 13 4 4 2
18 15 1 3 1 13 4 4 9 1 1 0 9 1 9 0 13 4 2
10 11 1 1 11 11 9 1 9 13 2
37 9 1 0 9 1 0 9 15 9 2 9 9 1 13 2 7 15 9 10 9 9 1 13 4 2 15 0 11 9 1 15 9 1 0 13 4 2
10 15 15 1 12 9 9 13 4 4 2
23 0 2 0 12 0 11 1 13 16 9 1 10 9 1 13 9 1 1 13 1 13 4 2
19 11 10 9 1 1 12 13 15 9 1 9 1 9 1 9 13 4 4 2
7 15 12 9 14 0 13 2
21 15 14 15 0 9 0 14 13 4 4 16 9 1 15 9 1 9 13 4 4 2
30 11 1 13 16 15 9 1 13 13 16 9 9 1 1 15 12 9 13 2 7 9 1 1 9 1 9 15 10 13 2
9 9 1 1 15 15 9 14 13 2
12 9 1 9 13 9 1 9 1 13 4 4 2
36 15 3 2 8 9 1 9 1 3 13 1 9 13 4 4 2 16 16 15 14 9 0 9 1 13 4 16 0 9 13 7 15 9 0 13 2
18 0 12 9 1 9 7 9 1 9 1 0 13 7 13 1 9 13 2
8 9 1 9 1 13 4 4 2
19 15 1 15 1 9 1 9 13 4 4 2 7 15 1 3 13 4 4 2
10 11 1 13 16 15 15 13 4 4 2
8 10 9 1 9 13 4 4 2
15 15 15 13 4 7 13 4 4 16 15 9 15 13 4 2
11 15 15 15 9 1 13 7 15 9 13 2
22 9 1 12 9 14 13 2 7 11 1 15 9 13 4 1 9 1 1 1 14 13 2
15 15 13 16 9 1 9 1 9 13 1 9 14 13 4 2
12 9 1 12 9 13 16 15 9 13 4 4 2
20 15 1 15 9 1 1 0 13 4 7 3 13 1 1 9 2 9 13 4 2
18 15 1 9 1 9 1 1 9 13 7 15 1 15 9 1 13 4 2
12 11 1 13 16 9 15 1 11 13 4 4 2
17 15 13 13 16 15 11 1 0 9 1 9 1 9 13 4 4 2
17 15 13 4 4 16 9 1 9 1 1 14 15 15 0 13 4 2
9 0 9 1 9 11 0 13 4 2
13 9 1 9 10 0 13 7 9 3 13 4 4 2
17 9 1 14 12 9 2 11 2 12 0 9 1 9 1 13 4 2
9 9 13 4 9 1 1 13 4 2
14 12 9 1 15 15 1 3 1 9 1 13 1 13 2
10 15 1 0 9 13 7 9 13 4 2
20 11 1 13 16 15 15 9 9 1 13 4 13 4 7 15 9 9 1 13 2
14 9 3 13 1 15 13 16 15 9 15 13 4 4 2
6 15 9 13 4 4 2
18 15 1 12 9 15 9 13 4 4 2 7 9 15 3 13 4 4 2
11 11 1 3 12 9 1 9 13 4 4 2
22 0 0 9 1 9 3 3 0 9 1 13 4 4 2 7 15 14 9 13 4 4 2
14 9 1 9 9 1 13 7 9 1 3 13 4 4 2
18 15 1 12 12 12 12 1 10 9 1 0 9 1 13 4 4 4 2
13 12 9 0 9 0 11 11 14 13 4 4 4 2
11 11 11 11 1 14 11 13 1 9 13 2
26 11 2 11 11 11 1 13 9 1 0 9 1 13 1 3 9 1 0 9 1 9 9 13 4 4 2
34 9 1 0 9 1 9 9 9 11 11 1 1 0 9 1 1 1 9 1 9 9 7 9 1 1 0 13 9 1 9 13 4 4 2
30 11 1 0 13 4 0 9 1 1 11 11 1 13 9 9 1 1 12 9 0 13 7 12 9 1 9 13 4 4 2
9 0 11 9 1 12 9 0 13 2
26 11 1 9 9 1 13 12 9 1 13 16 15 9 1 9 1 1 15 9 1 9 13 4 4 4 2
22 15 11 11 1 0 9 1 12 9 1 9 11 1 13 4 9 9 1 13 4 4 2
17 9 1 9 1 0 13 4 9 1 1 9 3 1 0 14 13 2
9 0 9 9 9 1 13 4 4 2
13 15 9 9 1 9 1 13 4 9 13 4 4 2
9 13 1 9 1 14 0 9 13 2
9 0 9 1 15 0 9 13 4 2
19 9 9 13 11 1 12 9 9 1 9 11 11 1 13 2 9 0 13 2
16 15 9 1 9 1 9 1 13 4 4 7 3 13 4 4 2
16 15 9 7 9 14 1 1 15 9 13 1 9 13 4 4 2
17 16 10 9 1 13 13 16 15 9 1 9 14 13 4 4 4 2
29 11 1 0 9 11 11 1 11 11 1 0 9 11 11 1 13 16 10 9 10 9 1 13 1 9 13 13 4 2
36 9 9 1 9 13 1 9 13 4 11 9 11 1 13 4 4 7 15 1 11 2 11 7 11 1 9 1 9 13 1 9 1 13 4 4 2
20 9 9 1 9 1 14 9 1 1 11 11 11 1 9 1 9 14 13 4 2
17 3 11 9 9 1 1 14 9 1 9 9 1 9 13 4 4 2
12 11 9 9 1 10 14 9 1 9 13 4 2
30 11 1 11 11 2 11 1 9 13 9 7 11 1 11 9 1 9 9 1 1 11 1 9 14 0 9 13 4 4 2
24 7 9 1 12 9 13 1 3 14 0 9 7 9 9 15 9 1 9 13 1 13 4 4 2
29 9 9 11 2 11 2 11 2 11 2 11 2 11 11 7 11 11 11 1 9 13 15 9 1 9 13 4 4 2
18 9 1 13 13 16 11 2 11 14 15 9 1 9 1 13 4 4 2
9 15 1 10 9 13 4 4 4 2
23 9 9 1 13 13 16 11 1 11 1 12 0 9 13 1 11 9 1 0 9 13 4 2
18 11 1 11 11 1 9 13 1 11 11 14 15 1 9 13 4 4 2
50 11 11 13 4 1 3 11 1 15 0 9 13 15 15 12 9 0 9 1 3 13 4 16 9 1 13 9 1 9 9 13 4 4 7 10 9 1 11 9 13 15 3 11 1 9 1 9 13 4 2
18 11 9 1 10 9 13 15 11 2 11 1 9 1 9 13 4 4 2
28 9 1 13 13 16 11 1 1 9 13 1 11 0 10 9 13 15 15 0 9 1 9 1 9 13 4 4 2
19 9 9 1 12 9 9 1 9 1 11 13 10 9 1 9 13 4 4 2
28 11 2 11 1 1 9 13 1 9 1 9 13 4 4 4 16 11 1 10 15 9 1 15 9 13 7 14 2
24 0 9 15 11 1 14 11 2 11 1 9 9 1 13 10 9 1 9 13 1 13 4 4 2
20 11 11 11 1 9 9 1 9 9 0 9 1 9 9 9 1 13 4 4 2
33 9 9 9 0 9 13 13 4 4 2 7 9 1 9 14 1 11 1 14 10 15 9 14 13 2 15 9 9 0 9 13 4 2
18 11 11 11 11 11 9 13 4 16 15 1 10 9 14 13 4 4 2
19 7 3 14 9 9 1 1 10 9 1 12 9 9 1 9 13 4 4 2
12 10 9 1 0 0 9 1 9 14 13 4 2
18 7 15 10 9 9 13 4 1 1 15 9 9 13 1 9 13 4 2
13 0 13 16 9 9 0 9 1 9 13 4 4 2
11 11 1 12 9 9 1 9 9 13 4 2
20 11 1 12 9 9 15 14 15 9 1 9 9 0 9 1 9 13 4 4 2
11 10 9 1 9 3 9 1 9 13 4 2
11 10 9 1 11 11 11 9 14 13 4 2
12 10 9 1 0 9 0 9 3 0 13 4 2
16 9 9 1 10 9 0 13 1 15 0 9 1 9 10 13 2
14 9 9 1 9 0 9 1 1 14 13 4 4 4 2
14 9 1 15 1 12 12 9 9 9 13 4 4 4 2
8 7 10 15 15 0 9 13 2
11 0 9 1 1 9 9 15 14 0 13 2
19 11 1 1 9 1 11 11 11 9 1 9 9 9 1 9 13 4 4 2
12 7 10 9 9 9 1 9 9 1 1 13 2
6 15 9 0 13 4 2
10 9 15 0 13 1 9 13 4 4 2
17 0 13 16 9 9 9 1 9 1 11 1 9 1 0 9 13 2
16 11 1 11 11 11 12 9 1 9 1 11 9 11 11 13 2
25 15 0 9 1 1 0 7 0 9 1 1 2 9 11 1 0 9 9 1 14 9 2 9 13 2
13 11 15 13 1 3 11 1 11 11 11 1 13 2
15 12 9 1 0 7 0 9 1 9 1 9 1 9 13 2
23 9 1 1 2 0 11 1 11 11 1 11 1 1 13 4 9 9 1 1 1 9 13 2
19 12 9 1 13 16 9 1 9 1 11 2 11 9 1 0 9 13 4 2
22 15 1 14 12 9 1 9 7 9 1 9 1 9 1 9 1 1 1 14 9 13 2
46 9 1 1 11 1 1 1 11 11 11 11 7 11 1 11 1 9 11 11 0 13 7 11 11 1 1 11 11 11 11 2 9 9 11 11 11 7 11 1 11 1 9 11 11 13 2
19 15 9 1 1 11 11 11 11 11 11 11 7 11 9 11 11 1 13 2
18 3 1 9 1 9 11 11 11 7 0 11 11 11 11 1 9 13 2
18 0 13 16 11 9 13 1 3 11 1 11 1 15 0 11 9 13 2
11 15 1 15 0 9 11 1 11 13 4 2
29 9 9 11 11 1 11 1 9 13 16 11 11 1 9 7 15 1 9 9 11 1 9 1 0 13 4 4 4 2
13 11 11 1 11 1 0 0 9 1 9 13 4 2
43 10 9 9 15 11 1 9 2 9 11 11 11 1 9 1 13 15 11 1 13 16 15 11 11 11 1 9 13 4 7 15 15 13 4 16 11 1 15 0 13 4 4 2
19 11 11 1 9 1 9 9 1 1 0 9 1 15 13 9 0 13 4 2
14 15 9 1 10 12 9 1 1 14 9 0 13 4 2
25 11 9 1 13 16 11 11 11 1 9 1 9 13 1 11 11 1 9 1 9 1 0 13 4 2
12 15 10 9 11 11 1 9 1 14 13 4 2
27 11 1 12 9 1 0 9 9 13 1 1 11 11 11 2 11 2 1 11 1 11 9 1 0 13 4 2
31 11 1 9 1 9 13 4 11 1 9 11 11 1 13 16 10 9 11 1 9 1 11 1 9 13 1 9 13 4 4 2
24 11 1 11 11 1 9 13 4 11 1 13 16 15 9 12 1 12 9 1 13 14 1 13 2
10 10 9 9 9 1 1 0 14 13 2
22 11 1 13 16 10 9 1 14 9 13 16 11 9 1 1 15 9 1 3 13 4 2
27 11 1 13 16 15 11 1 0 11 1 9 1 15 9 14 13 7 3 15 0 9 13 1 0 14 13 2
21 11 1 13 16 15 13 4 16 11 11 1 12 0 9 7 9 1 9 0 13 2
15 15 13 4 1 16 11 1 11 1 11 1 9 15 13 2
15 11 1 13 16 15 15 9 1 9 1 9 1 13 4 2
28 11 1 11 11 1 11 1 0 13 4 11 11 11 2 11 2 1 9 1 0 7 9 1 9 9 13 4 2
13 11 1 13 16 10 9 9 1 0 9 9 13 2
18 15 15 9 1 9 1 10 9 13 1 13 4 15 0 9 13 4 2
46 11 11 2 11 2 1 0 9 1 9 9 7 9 1 9 13 4 1 9 1 1 1 11 1 13 16 9 1 14 0 7 9 1 9 1 0 9 1 9 1 1 9 1 9 13 2
12 15 9 1 9 1 9 1 15 9 14 13 2
20 7 11 1 9 1 9 1 1 11 11 11 9 13 4 1 9 1 9 13 2
22 11 9 9 1 9 9 7 9 0 13 0 9 7 9 1 9 1 9 1 1 13 2
23 11 11 2 11 11 11 11 11 11 11 11 1 11 1 15 12 9 9 1 10 9 13 2
30 15 13 16 10 9 1 1 11 11 11 11 11 3 0 9 13 2 15 0 10 9 1 9 1 10 9 1 9 13 2
37 9 7 9 9 1 0 0 9 1 9 11 11 1 13 16 10 9 7 9 1 10 9 7 9 2 9 2 9 2 9 9 1 9 14 9 13 2
13 10 3 13 1 9 9 1 10 9 1 0 13 2
25 11 11 1 9 1 9 9 1 9 1 13 4 11 1 0 11 1 1 9 14 0 13 4 4 2
24 15 11 1 15 9 1 9 13 4 11 11 1 9 13 16 15 11 1 11 9 1 9 13 2
40 7 9 1 11 11 1 11 11 11 1 9 13 4 16 11 11 11 1 9 13 4 16 11 11 11 11 1 0 9 1 9 1 9 1 9 2 9 13 4 2
12 11 1 10 9 1 11 1 12 9 13 4 2
22 9 15 9 13 16 11 1 9 3 0 13 4 16 11 9 1 9 0 14 13 4 2
42 11 9 11 11 1 15 9 1 9 1 9 1 1 9 1 13 16 11 1 9 1 9 1 9 0 13 15 0 9 1 1 0 9 11 11 1 11 13 4 4 4 2
26 9 9 1 9 0 13 1 1 9 13 1 9 1 11 1 13 16 9 1 0 13 1 13 4 4 2
13 15 0 7 0 9 0 9 1 9 0 13 4 2
24 11 1 11 1 1 1 13 4 1 15 13 16 16 15 15 9 1 9 13 4 16 9 13 2
36 11 1 11 1 13 11 9 9 1 11 1 0 9 9 13 7 9 1 9 1 1 15 12 9 1 0 9 11 11 1 14 13 4 4 4 2
14 11 1 9 14 13 1 1 1 9 1 15 9 13 2
24 11 1 11 11 11 1 9 13 4 13 4 16 11 9 1 9 12 9 1 1 13 4 4 2
32 11 9 1 1 1 15 0 11 11 11 1 9 1 0 13 4 13 16 10 9 1 11 1 1 11 1 10 9 13 4 4 2
25 11 1 13 4 16 11 9 1 11 1 1 13 4 12 0 9 1 14 10 0 9 13 4 4 2
25 11 1 11 11 11 11 1 0 9 9 1 13 4 16 11 9 1 9 1 15 15 9 14 13 2
8 11 15 1 9 13 4 4 2
18 11 1 2 0 9 2 11 2 1 1 12 9 1 10 9 13 4 2
32 11 11 1 15 9 1 1 1 11 1 13 16 15 11 9 1 9 1 1 11 1 1 15 9 9 13 1 1 14 13 4 2
28 15 13 16 11 9 1 9 1 9 1 9 1 9 1 14 12 9 9 13 1 0 9 1 3 14 13 4 2
27 0 11 11 11 11 11 1 9 1 1 1 13 4 9 1 11 1 13 16 15 15 1 15 9 14 13 2
12 10 9 11 1 0 9 11 11 11 1 13 2
18 11 1 9 13 16 0 11 11 11 9 1 0 9 13 1 0 13 2
23 11 1 0 9 13 1 1 1 15 13 16 10 9 1 9 15 9 0 14 13 13 4 2
28 11 1 13 16 15 15 15 14 13 16 11 1 15 9 13 7 15 14 14 13 16 15 15 9 15 14 13 2
22 11 1 13 16 16 0 9 7 11 11 1 15 9 13 4 16 11 14 3 14 13 2
13 11 1 13 16 15 15 0 9 1 9 14 13 2
20 15 9 13 13 16 15 11 1 15 9 1 0 9 1 9 1 0 9 13 2
22 9 1 13 0 9 2 11 7 11 2 1 9 11 11 1 9 7 9 1 9 13 2
35 12 0 11 7 11 1 9 11 1 13 16 16 9 13 4 4 16 10 9 1 0 13 4 4 4 16 15 9 1 15 13 4 4 4 2
35 11 1 0 2 0 9 9 11 11 1 10 9 13 16 10 12 9 1 9 1 1 0 13 4 4 4 2 11 1 9 10 13 4 4 2
15 11 1 10 12 9 1 11 9 1 11 0 9 13 4 2
17 15 13 16 11 9 15 1 11 1 1 9 1 9 13 13 4 2
23 16 15 15 0 2 0 13 16 15 11 7 11 1 10 0 9 1 0 13 13 4 4 2
12 11 1 9 11 9 9 1 1 9 13 4 2
15 11 1 13 16 15 9 1 9 13 4 16 9 0 13 2
11 15 15 9 1 9 1 14 0 13 4 2
19 11 11 1 9 9 11 11 11 11 11 1 1 15 9 0 13 13 14 2
26 15 13 16 16 0 9 11 7 11 1 3 13 1 0 13 4 16 15 3 0 9 11 11 1 13 2
17 15 0 9 15 14 13 16 10 0 9 1 12 9 9 13 4 2
25 16 11 11 9 1 9 9 13 1 1 3 14 13 16 15 10 12 9 1 9 15 13 4 4 2
31 15 13 16 15 14 9 1 10 14 13 16 15 1 12 9 1 13 4 11 1 15 10 12 9 1 9 1 9 13 4 2
26 15 9 13 16 12 9 10 9 1 9 1 9 13 7 9 0 9 1 15 2 15 1 0 13 4 2
34 11 9 1 11 11 1 11 7 11 1 12 0 9 13 4 15 13 4 4 16 11 1 0 9 1 11 11 1 9 13 4 4 4 2
25 3 1 9 1 13 4 4 16 9 9 1 0 13 1 9 0 9 1 1 13 4 9 1 13 2
11 10 9 11 11 2 11 1 9 1 13 2
19 11 1 0 9 1 0 13 1 1 15 14 9 9 1 9 1 9 13 2
29 7 11 7 11 1 13 4 0 9 1 1 11 1 0 9 1 0 9 1 9 1 1 14 0 13 4 4 4 2
29 10 9 1 11 1 11 11 11 11 1 14 13 4 16 9 9 1 9 1 9 11 1 0 9 1 1 13 4 2
14 10 9 1 9 9 9 1 10 9 1 14 13 4 2
20 11 1 0 9 1 9 1 9 9 1 9 1 9 13 1 9 3 10 13 2
29 16 11 11 11 1 11 1 14 9 9 1 0 13 4 11 1 9 9 1 10 10 9 1 13 1 9 13 4 2
14 15 14 13 1 15 11 1 9 9 1 9 13 4 2
14 9 1 9 1 9 1 9 1 0 9 0 3 13 2
19 15 1 0 9 1 9 7 11 11 1 10 9 1 3 10 9 13 4 2
15 11 11 1 14 0 9 1 9 1 3 10 9 13 4 2
16 11 9 1 1 9 7 11 11 1 9 9 1 9 13 4 2
18 7 10 9 11 11 1 9 13 1 1 9 1 9 9 13 4 4 2
16 15 1 0 0 9 1 14 12 12 9 9 1 9 13 4 2
15 15 3 10 9 11 1 13 4 7 11 0 9 1 13 2
22 11 11 11 1 9 1 1 11 11 1 15 1 14 12 12 9 9 1 9 13 4 2
10 15 15 9 1 13 4 10 10 13 2
13 10 9 11 1 12 12 9 9 1 9 13 4 2
28 0 9 1 0 9 1 15 1 12 12 9 9 1 9 13 4 4 2 15 0 9 1 1 1 3 0 13 2
14 11 11 11 14 12 12 9 9 1 9 13 4 4 2
14 7 9 9 1 12 12 9 14 9 1 9 13 4 2
13 15 1 9 9 9 1 12 12 9 9 13 4 2
14 9 1 1 0 9 1 9 1 11 9 0 3 13 2
14 15 15 1 12 12 9 1 10 9 1 9 13 4 2
16 7 11 1 12 12 9 9 9 1 0 9 1 13 4 4 2
15 15 1 11 11 1 10 9 1 12 12 9 9 13 4 2
24 13 1 9 15 13 16 9 1 9 1 9 1 9 9 1 9 13 1 9 14 3 14 13 2
16 10 9 15 1 12 12 9 1 10 9 1 9 13 4 4 2
15 7 9 1 0 9 9 1 9 15 9 14 0 13 4 2
13 0 0 9 1 9 9 1 12 12 9 9 13 2
31 11 11 11 11 1 10 9 9 13 4 15 0 9 11 11 1 11 11 11 11 11 2 11 2 1 9 1 0 9 13 2
19 15 9 13 4 11 1 9 11 11 11 1 10 9 1 9 9 9 13 2
27 11 1 11 9 2 11 11 11 11 1 2 9 1 15 9 13 4 0 11 1 0 9 1 9 13 4 2
12 15 13 16 9 1 9 10 0 7 0 13 2
30 16 15 3 10 9 0 13 13 4 7 9 1 11 11 1 0 9 1 13 13 4 16 15 10 0 9 13 14 4 2
13 11 1 13 2 15 14 12 9 1 9 14 13 2
7 15 12 12 0 9 13 2
34 11 1 9 1 9 0 13 4 9 11 1 13 16 11 15 12 9 2 12 9 9 7 12 12 11 1 1 9 9 9 13 4 4 2
21 10 9 10 9 1 9 13 16 15 0 9 0 7 0 9 1 9 13 4 4 2
13 15 13 16 11 9 1 12 0 9 1 1 13 2
8 15 9 14 1 9 0 13 2
36 11 1 15 9 1 9 1 9 9 1 9 13 4 1 11 11 1 9 1 9 13 4 16 15 0 9 1 9 1 13 0 9 1 9 13 2
14 9 9 1 9 13 2 7 9 14 15 1 9 13 2
28 15 13 16 9 1 10 9 12 9 11 1 9 1 13 4 4 2 7 10 9 1 10 9 14 13 4 4 2
10 9 15 13 16 15 9 1 9 13 2
31 11 2 11 1 9 1 9 2 9 1 0 9 13 4 1 1 9 1 9 1 0 9 1 9 13 1 0 9 13 4 2
16 9 1 0 12 9 1 0 9 1 9 1 0 9 13 4 2
17 0 9 1 1 9 1 0 9 1 12 9 1 1 9 13 4 2
21 11 11 1 9 1 3 12 0 9 13 4 3 10 9 14 12 0 9 13 4 2
24 9 1 1 3 9 11 1 0 9 1 12 9 13 4 4 3 11 1 12 9 13 4 4 2
15 9 1 9 1 0 9 2 9 7 9 1 9 0 13 2
19 9 11 1 9 1 12 9 0 0 9 13 4 7 12 9 13 4 4 2
12 9 1 9 1 9 1 1 14 0 9 13 2
36 9 1 11 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 2 11 2 11 2 11 1 10 9 1 13 1 9 0 13 2
13 9 1 9 1 3 0 9 11 11 1 13 4 2
17 10 9 1 1 10 0 9 1 15 12 0 9 1 9 13 4 2
15 9 11 1 1 12 0 7 12 0 9 9 1 13 4 2
10 7 10 9 10 9 12 7 12 13 2
16 9 11 1 12 0 7 12 0 9 9 1 9 13 4 4 2
19 9 1 9 2 9 1 0 9 13 1 1 9 1 9 1 9 0 13 2
34 9 11 1 9 1 1 9 1 3 12 9 7 9 13 4 4 3 10 9 10 9 13 12 1 13 7 9 11 1 10 9 12 13 2
17 0 9 1 1 14 0 0 9 1 12 9 1 1 9 13 4 2
35 11 11 1 11 11 11 11 1 11 7 11 11 1 9 9 1 9 13 1 3 15 11 1 11 11 1 14 11 1 1 9 13 4 4 2
14 15 14 9 13 4 16 11 15 9 9 13 4 4 2
15 11 1 11 11 11 11 1 9 9 1 11 1 9 13 2
35 15 1 12 9 0 13 11 1 11 1 13 16 2 15 15 1 10 9 1 0 13 1 13 4 16 15 0 13 16 11 15 9 1 13 4
58 2 15 13 16 15 7 11 11 1 10 9 1 0 9 0 13 4 4 16 0 9 1 9 9 1 1 11 1 9 13 15 10 9 1 3 0 9 13 4 4 7 15 2 9 2 1 9 13 1 1 0 9 1 0 9 13 4 2
20 16 2 9 1 11 1 15 14 13 4 16 11 1 3 15 9 13 4 4 2
15 11 1 10 0 9 9 1 0 13 1 7 0 13 4 2
30 15 3 13 16 15 13 10 14 9 13 4 4 16 11 11 15 0 9 1 9 13 1 10 9 1 3 13 4 4 2
28 11 1 13 16 2 15 3 14 0 7 0 9 13 15 9 1 0 13 1 9 7 13 1 9 1 3 9 13
28 15 10 9 0 13 4 16 16 15 11 11 1 1 13 4 4 16 15 15 14 0 9 1 1 13 4 4 2
27 11 11 7 15 0 9 11 11 1 1 0 9 1 13 13 4 9 1 0 13 1 9 13 4 4 4 2
35 13 4 4 4 16 12 9 1 1 9 1 0 9 0 13 4 4 4 7 9 13 16 0 12 9 1 1 15 0 9 9 13 4 4 2
13 9 1 9 12 2 12 9 1 13 4 4 4 2
20 16 9 1 9 1 9 7 0 9 0 13 1 12 9 1 9 13 4 4 2
15 0 9 1 1 9 11 1 13 9 1 9 13 4 4 2
36 9 1 13 13 16 9 1 9 9 1 0 9 1 13 13 10 3 0 9 1 13 1 9 1 0 12 9 1 1 9 9 1 9 13 4 2
39 11 11 1 13 4 4 4 16 11 11 15 9 1 13 2 15 13 9 1 9 13 2 7 9 1 9 13 4 16 10 9 11 1 9 1 13 4 4 2
18 3 15 11 11 7 11 11 14 13 4 4 2 15 9 11 11 13 2
56 12 9 1 1 10 9 1 0 9 13 4 2 15 1 0 10 9 1 11 11 1 10 0 9 9 13 4 2 15 0 9 11 1 13 4 7 0 9 11 11 11 2 11 2 7 11 11 11 1 11 1 0 9 0 13 2
23 9 1 3 0 9 9 1 9 1 1 13 4 4 9 1 11 11 11 11 1 9 13 2
27 0 9 15 13 4 16 11 9 9 1 1 13 4 4 7 0 9 1 9 1 9 13 1 9 14 13 2
26 11 1 13 16 12 9 9 2 9 1 15 9 13 4 4 7 15 15 9 3 13 1 9 13 4 2
12 15 13 4 16 3 14 15 15 9 13 4 2
21 11 11 1 1 9 9 1 9 14 10 9 1 13 9 1 0 9 13 4 4 2
17 9 1 1 12 9 1 13 9 1 13 1 9 1 9 13 4 2
24 16 2 9 1 15 14 13 13 16 9 1 9 1 11 7 11 1 1 0 9 14 13 4 2
24 7 9 1 0 9 13 4 1 3 10 9 1 0 9 1 1 11 9 1 9 13 4 4 2
41 11 11 11 1 0 9 11 11 7 0 9 11 11 1 15 15 1 13 4 9 2 9 1 9 1 1 11 11 1 0 0 0 9 11 1 15 9 9 13 4 2
11 9 1 11 1 10 9 1 9 13 4 2
26 0 9 1 9 9 9 9 9 1 9 1 10 9 1 11 9 1 9 9 11 11 11 14 0 13 2
18 9 1 12 9 1 9 1 9 15 1 0 13 1 1 9 13 4 2
22 9 1 9 12 9 1 15 9 13 4 16 11 7 11 1 3 9 15 13 4 4 2
39 9 1 2 0 2 13 4 9 11 11 7 11 11 11 1 9 1 0 9 1 9 9 1 11 9 1 9 9 1 15 9 1 9 13 1 9 13 4 2
20 15 0 9 1 0 11 1 9 7 11 1 9 1 9 1 9 13 1 13 2
25 9 13 1 3 9 9 1 9 9 11 11 11 1 9 13 7 11 1 10 9 1 1 13 4 2
41 0 13 16 11 9 2 9 1 15 9 1 3 13 4 7 15 0 9 1 15 9 13 4 16 11 1 15 1 9 13 7 11 11 11 1 9 1 13 9 13 2
28 11 1 9 1 9 13 16 11 1 0 11 7 11 9 1 9 13 1 1 11 1 0 9 13 1 9 13 2
27 10 9 9 13 1 12 9 1 11 1 11 9 1 15 9 1 12 0 9 13 15 12 9 0 13 4 2
24 7 9 9 9 1 9 1 10 9 1 11 2 11 11 1 12 11 0 13 0 9 13 4 2
6 15 9 12 9 13 2
11 9 1 13 13 16 15 15 9 14 13 2
12 11 11 11 11 11 1 9 1 11 0 13 2
21 9 1 10 9 1 9 9 1 13 1 3 15 12 9 1 9 1 9 13 4 2
38 12 0 9 1 12 9 1 13 4 16 9 9 9 9 1 12 9 9 1 9 0 13 4 4 4 7 16 15 9 13 4 16 15 9 1 9 13 2
26 11 11 2 11 11 11 2 11 11 7 11 11 11 1 1 1 0 10 9 1 15 1 9 14 13 2
30 10 3 11 11 1 11 11 1 9 1 9 1 9 1 9 9 9 0 13 4 7 10 9 1 12 9 0 13 4 2
11 15 11 11 1 12 0 9 9 0 13 2
26 11 9 1 11 9 1 9 9 12 12 9 12 9 9 1 1 13 11 9 1 12 9 0 13 4 2
10 10 9 12 9 1 9 13 4 4 2
27 0 9 1 13 16 15 1 9 12 12 9 11 9 1 11 1 12 9 1 9 1 9 12 11 0 13 2
16 9 9 1 13 10 9 1 9 3 12 9 7 12 9 13 2
8 9 9 1 15 8 13 4 2
18 9 7 11 9 1 10 12 9 11 2 11 11 11 1 9 1 13 2
9 15 1 12 9 11 1 0 13 2
26 0 9 11 7 11 1 1 9 9 1 12 9 14 9 9 1 10 9 11 1 10 9 1 9 13 2
27 11 1 13 9 1 13 4 4 16 11 1 11 13 1 9 1 9 1 12 9 1 9 13 4 4 4 2
15 15 11 11 11 7 11 11 11 1 12 0 9 0 13 2
16 11 9 9 1 11 1 3 13 1 9 3 0 13 4 4 2
21 11 1 9 13 4 16 15 11 11 11 2 11 2 1 10 9 1 1 9 13 2
17 11 1 3 9 13 1 9 1 11 1 1 15 9 14 13 4 2
17 3 0 9 1 1 11 9 11 11 3 14 11 11 1 9 13 2
29 11 9 7 11 1 9 11 11 1 13 4 16 11 11 15 1 13 7 9 1 2 3 1 15 9 14 13 4 2
15 11 1 3 9 13 1 15 10 9 1 1 11 9 13 2
37 11 1 11 1 15 13 4 11 1 0 9 1 9 13 4 16 15 0 9 1 1 15 9 14 13 2 7 11 1 10 9 1 0 13 4 4 2
9 15 14 9 1 10 9 14 13 2
17 15 11 9 11 11 1 11 1 9 1 15 3 0 9 13 4 2
11 15 9 11 1 10 9 1 0 14 13 2
21 15 13 13 16 9 11 1 3 1 9 13 4 4 2 7 11 9 1 0 13 2
16 11 16 3 13 9 13 4 16 15 9 1 3 13 4 4 2
17 11 11 1 13 16 9 9 1 1 11 1 0 9 9 13 4 2
16 15 1 2 9 0 9 0 13 1 14 9 13 4 4 4 2
9 16 11 1 15 1 10 9 13 2
37 15 13 4 1 16 15 11 1 9 1 10 9 0 13 4 4 2 11 1 13 16 11 9 1 13 1 3 11 9 11 11 12 9 15 9 13 2
18 2 11 2 1 10 9 9 1 1 9 11 1 9 15 2 14 13 2
15 11 11 1 9 9 1 9 1 15 12 9 1 13 4 2
8 15 1 10 9 7 9 13 2
11 15 9 9 1 3 0 9 1 13 4 2
10 12 9 1 14 12 9 13 4 4 2
11 15 13 0 9 1 12 9 13 4 4 2
30 9 2 9 2 9 2 9 7 0 2 9 9 15 0 13 4 7 9 13 9 1 9 15 9 1 1 9 13 4 2
16 15 1 10 14 9 1 15 9 1 1 11 11 11 0 13 2
17 9 9 1 9 1 14 13 4 2 7 15 15 0 9 14 13 2
14 2 9 2 1 12 9 10 9 9 1 1 0 13 2
10 9 1 9 1 3 9 0 13 4 2
16 12 9 1 13 9 1 0 11 1 12 9 1 9 13 4 2
10 9 1 11 7 11 9 3 0 13 2
9 15 11 7 11 9 14 0 13 2
10 11 1 12 1 10 9 1 9 13 2
12 9 9 1 13 1 10 9 0 13 4 4 2
11 15 14 13 0 9 15 1 15 1 13 2
11 9 1 9 13 15 9 1 8 13 4 2
23 12 9 9 1 9 14 1 9 1 9 13 4 2 7 9 1 9 9 1 14 13 4 2
12 9 9 1 9 1 9 9 0 13 4 4 2
23 9 1 1 9 1 1 1 3 12 9 9 2 12 9 9 7 12 9 9 13 4 4 2
17 9 14 1 9 1 1 9 1 13 4 9 14 13 4 4 4 2
18 9 1 15 9 9 11 1 11 7 11 1 9 1 14 9 13 4 2
28 9 14 1 12 12 0 9 1 1 9 13 1 9 13 1 9 1 9 9 1 9 1 1 1 13 4 4 2
23 9 1 1 9 13 7 0 9 1 9 1 1 9 1 12 12 1 9 1 9 13 4 2
16 9 1 11 1 11 7 11 1 14 9 9 1 9 13 4 2
28 9 1 9 1 11 11 1 9 9 9 9 11 11 1 9 1 10 9 11 13 9 1 9 1 13 4 4 2
13 11 1 9 11 1 1 10 9 1 0 0 13 2
32 11 1 1 0 9 9 9 1 15 3 12 9 1 9 0 13 2 3 15 11 11 11 1 1 1 12 0 9 9 13 4 2
19 9 1 14 0 9 13 4 11 1 0 9 1 1 0 9 0 9 13 2
36 11 1 9 3 9 13 4 11 1 12 9 1 12 9 1 1 12 9 1 12 9 1 12 13 2 15 11 1 1 11 1 3 0 9 13 2
17 9 9 9 11 1 15 9 1 12 9 7 12 0 9 14 13 2
9 15 1 15 0 9 12 9 13 2
18 9 1 13 13 11 1 0 9 12 9 1 12 9 13 8 13 4 2
16 11 1 11 1 13 4 0 9 9 9 12 9 1 13 4 2
18 10 9 1 11 1 9 9 1 12 2 12 1 9 0 13 4 4 2
21 9 11 11 1 9 12 0 11 1 9 13 4 15 0 13 0 9 1 13 13 2
10 15 1 10 15 13 15 9 13 4 2
25 11 2 11 1 0 9 2 0 9 7 9 1 1 0 9 1 11 0 9 1 9 13 13 4 2
36 11 1 1 3 1 1 9 14 11 11 1 9 13 7 14 12 9 1 12 9 7 12 9 1 9 1 12 9 13 0 9 1 9 13 4 2
13 0 9 1 1 12 9 1 12 9 1 9 13 2
14 11 1 15 0 9 1 14 12 9 1 9 0 13 2
16 9 11 2 11 2 11 1 9 1 15 9 11 11 1 13 2
10 10 3 11 9 9 1 13 4 4 2
28 14 12 9 1 15 15 9 0 13 15 9 1 0 12 9 1 15 13 4 9 1 9 1 9 1 9 13 2
23 9 11 11 12 9 3 9 1 0 14 13 7 12 9 13 11 1 9 1 8 13 4 2
32 11 1 3 13 13 9 9 11 11 1 13 4 9 1 9 1 9 13 7 0 9 9 1 9 1 13 1 0 9 0 13 2
14 0 9 1 12 9 1 12 9 1 12 9 13 4 2
10 11 1 12 9 1 15 9 0 13 2
26 11 1 9 1 0 9 1 11 1 3 9 13 7 12 9 7 12 9 1 9 1 12 9 13 4 2
30 15 1 9 13 9 1 0 9 13 1 3 0 13 4 11 0 9 1 11 11 1 9 1 11 11 1 9 13 4 2
16 11 1 11 1 1 12 9 1 0 0 9 1 14 13 4 2
23 15 1 10 9 11 11 2 11 2 11 2 7 11 11 2 11 2 11 2 1 9 13 2
10 11 11 1 9 11 1 10 0 13 2
20 16 2 9 1 9 1 11 1 15 9 13 2 15 15 9 1 14 13 4 2
26 11 11 11 2 11 2 1 11 1 11 11 1 13 9 1 1 12 9 9 1 9 1 9 13 4 2
45 12 12 9 9 1 0 11 2 11 11 1 1 9 9 9 1 9 1 1 0 9 1 9 9 1 1 9 2 9 13 1 11 11 1 1 0 9 13 1 9 14 13 4 4 2
12 11 11 11 11 11 1 11 1 11 0 13 2
23 9 13 4 4 4 16 15 11 1 11 1 9 1 0 9 1 9 1 13 1 9 13 2
19 11 1 11 11 11 11 11 1 1 9 1 1 15 10 9 1 9 13 2
13 11 1 11 11 1 11 11 1 0 9 1 13 2
25 11 1 9 9 1 9 13 1 9 1 11 15 9 1 0 9 9 1 9 1 13 1 9 13 2
21 9 1 10 9 13 4 13 16 9 0 9 1 9 9 1 1 13 1 9 13 2
13 11 11 1 3 12 12 9 9 1 9 13 4 2
12 11 2 11 9 1 15 1 15 9 14 13 2
16 15 0 9 1 9 7 9 1 11 1 9 1 0 13 4 2
22 15 13 16 11 0 9 1 9 9 9 1 9 13 4 4 7 0 11 13 4 4 2
25 9 1 11 9 1 9 1 11 13 4 4 4 7 15 1 9 7 9 1 11 13 4 4 4 2
19 9 1 11 1 12 9 1 9 1 1 12 9 9 13 1 9 13 4 2
28 11 11 1 9 1 1 11 1 0 9 1 9 9 1 1 11 7 11 1 3 13 1 9 1 14 9 13 2
25 9 1 13 16 11 11 2 11 2 11 9 1 9 7 11 1 15 9 1 9 1 9 14 13 2
26 11 11 11 1 11 9 11 11 1 12 9 1 9 11 1 15 1 9 14 13 4 1 9 13 4 2
24 11 1 9 11 11 1 9 1 9 0 13 11 1 9 13 4 1 9 13 1 9 13 4 2
36 11 11 1 9 1 9 11 11 1 11 1 9 0 13 4 15 9 13 16 15 9 1 0 9 1 14 15 9 1 9 1 1 14 13 4 2
34 0 13 16 11 1 11 1 11 1 9 11 11 1 9 13 4 7 15 12 9 1 14 9 1 9 13 4 7 9 9 1 13 4 2
26 15 10 14 9 13 4 16 11 1 9 1 9 1 9 13 1 1 1 11 1 12 12 9 13 4 2
27 11 11 1 15 9 1 13 4 16 15 10 9 13 4 16 11 11 1 13 11 13 1 9 13 4 4 2
8 15 1 15 9 14 13 4 2
25 11 1 15 9 1 15 14 13 4 16 10 9 1 9 1 13 15 0 9 1 9 0 13 4 2
16 15 0 13 1 3 11 1 9 9 1 15 9 14 13 4 2
19 10 9 1 9 1 11 7 11 11 11 2 11 2 1 9 0 13 4 2
46 11 1 9 1 0 9 11 11 1 13 15 15 13 4 16 11 1 0 9 1 15 0 9 1 9 9 0 13 4 7 15 9 1 9 1 9 1 1 1 11 11 1 9 0 13 2
17 11 1 13 16 15 11 11 1 13 9 1 9 1 1 13 4 2
32 11 11 1 9 11 11 1 11 1 15 13 16 11 1 11 1 9 1 9 9 1 1 11 11 1 1 10 9 1 9 13 2
23 15 13 16 15 15 13 16 11 1 11 1 10 0 9 7 11 1 10 11 0 9 13 2
46 11 11 1 9 11 11 1 0 9 1 13 9 1 13 16 11 15 0 0 9 1 1 10 9 1 9 1 13 4 4 15 15 9 9 13 1 1 9 1 9 13 9 13 4 4 2
28 11 1 11 1 11 1 9 9 9 1 9 1 9 1 13 16 15 9 13 4 16 11 1 3 9 13 4 2
20 7 15 9 1 9 15 0 13 4 4 7 9 1 9 1 9 13 4 4 2
13 11 1 13 16 11 1 11 1 1 10 0 13 2
13 11 1 0 9 13 7 11 1 1 0 9 13 2
19 11 11 11 2 11 2 1 0 0 9 1 12 0 9 9 13 4 4 2
26 15 3 0 13 11 9 9 1 9 1 9 1 9 1 13 1 9 1 15 9 13 1 9 14 13 2
35 11 1 9 1 10 0 9 10 9 1 13 4 15 15 15 0 9 11 1 0 0 9 1 1 13 1 1 3 2 3 9 13 4 4 2
27 11 9 11 11 11 1 13 9 9 9 1 9 1 1 11 1 9 1 13 0 9 1 1 14 0 13 2
22 15 12 9 1 0 9 1 11 1 11 7 15 0 9 1 9 1 9 1 0 13 2
35 0 9 1 15 11 1 0 9 16 9 1 11 1 0 9 11 11 11 1 9 1 9 1 0 9 1 1 1 9 13 1 1 13 4 2
28 9 1 9 1 9 9 1 13 4 1 11 1 9 1 1 14 11 11 1 9 14 1 9 1 9 9 13 2
20 15 9 1 11 1 13 16 9 9 1 13 10 9 1 1 10 0 9 13 2
18 10 9 1 0 9 1 9 9 1 0 13 4 9 9 14 0 13 2
21 11 1 10 9 1 11 1 9 1 12 9 1 1 12 9 1 13 1 9 13 2
20 10 9 1 11 1 13 0 9 2 0 2 0 9 7 9 1 9 0 13 2
30 9 1 11 11 11 7 11 1 9 1 11 2 11 1 0 9 13 1 11 11 1 13 1 9 14 14 13 4 4 2
23 9 1 9 1 11 9 9 1 1 9 1 9 1 10 12 9 9 1 13 4 4 4 2
31 11 9 11 11 1 15 10 0 9 1 13 1 1 1 13 4 15 15 9 13 16 15 15 10 9 1 0 14 13 4 2
10 10 9 1 0 9 14 13 4 4 2
26 11 1 11 11 11 11 1 11 1 11 11 11 11 1 0 9 1 11 1 9 1 0 9 13 4 2
22 15 1 14 15 11 1 9 2 9 7 9 1 9 1 0 13 1 9 14 13 4 2
18 11 7 11 1 0 9 1 9 1 1 12 0 9 1 9 13 4 2
33 11 1 12 9 1 9 1 13 11 1 13 16 11 1 12 9 1 15 9 1 1 9 13 4 7 15 15 15 9 13 13 4 2
34 15 1 14 15 13 16 11 1 11 11 1 9 13 16 11 1 0 9 11 1 11 1 9 1 1 9 7 9 9 1 9 13 4 2
46 11 11 11 1 1 9 1 1 11 1 15 12 9 9 1 13 16 11 11 11 11 1 3 10 0 13 7 0 9 1 9 2 9 7 15 9 1 1 11 1 15 9 13 4 4 2
25 15 13 16 11 11 1 0 13 4 7 9 1 9 1 0 13 4 11 11 1 9 13 4 4 2
31 13 4 4 4 16 15 1 11 11 7 11 1 9 1 1 12 9 1 0 9 1 1 2 9 0 9 1 0 9 13 2
23 9 1 1 12 9 1 9 1 12 9 1 12 9 1 9 13 7 12 0 9 0 13 2
29 9 9 1 11 1 9 13 16 11 1 0 12 9 1 15 9 1 1 9 13 4 4 7 15 9 13 13 4 2
20 11 1 13 16 16 15 15 13 4 2 16 15 1 11 1 11 11 0 13 2
21 15 1 14 15 13 16 11 11 11 1 1 15 9 1 11 1 1 0 9 13 2
32 15 1 14 15 13 16 11 1 11 11 1 9 13 16 11 1 0 9 11 1 9 1 1 9 7 9 9 1 9 13 4 2
36 16 11 1 10 9 1 11 7 11 1 3 15 9 0 14 13 4 7 0 9 1 1 1 14 15 10 9 1 9 1 0 14 13 4 4 2
29 15 13 16 11 1 0 9 1 11 11 11 1 9 1 15 9 9 1 9 7 9 9 1 9 1 9 13 4 2
40 11 11 11 11 2 11 2 1 11 1 13 16 11 2 11 11 11 1 15 12 9 1 13 1 1 11 1 11 11 11 1 0 13 15 2 0 9 2 13 2
13 12 9 1 1 9 0 9 1 9 13 4 4 2
33 7 16 11 11 11 1 11 11 1 0 0 11 2 11 12 0 9 1 13 1 9 13 4 16 15 15 9 13 1 1 0 13 2
39 11 1 9 11 11 1 13 16 16 11 7 11 1 1 15 9 1 13 1 1 11 1 11 1 9 1 9 14 13 2 16 14 12 0 9 1 13 4 2
29 7 16 15 9 13 4 16 10 9 11 11 7 11 1 13 4 16 15 2 9 11 2 15 9 1 13 13 4 2
12 15 13 16 0 11 1 0 9 0 13 4 2
17 11 1 9 11 11 11 1 11 1 13 16 15 11 1 11 13 2
18 15 15 0 13 9 13 2 7 9 9 1 9 7 11 11 13 4 2
16 3 11 1 11 1 0 13 1 9 1 9 11 1 13 4 2
27 11 1 13 9 1 13 4 4 16 11 11 13 12 9 1 1 9 1 15 12 9 1 13 1 0 13 2
24 11 1 13 15 15 1 1 15 9 9 14 13 4 2 15 11 1 11 13 1 9 13 4 2
14 10 9 1 11 11 11 1 1 1 9 14 13 4 2
35 3 2 11 1 11 9 1 9 1 9 1 13 16 9 1 11 1 0 9 1 1 15 11 2 11 7 11 7 11 9 1 0 13 4 2
13 16 11 1 11 15 13 4 16 15 0 9 13 2
26 9 1 1 11 9 1 9 0 13 1 9 1 11 1 13 16 15 15 1 1 15 9 14 13 4 2
17 7 10 9 1 9 1 9 13 4 16 15 0 9 0 13 4 2
19 15 13 16 15 14 12 9 1 1 9 1 9 1 12 9 1 0 13 2
23 15 13 16 9 1 1 9 1 1 1 9 1 1 9 1 9 14 14 13 4 13 4 2
24 11 1 13 16 11 1 10 9 1 1 13 1 9 2 9 7 9 1 1 0 9 13 4 2
17 11 11 11 11 11 1 0 9 1 9 12 13 1 9 13 4 2
16 15 9 1 9 13 1 9 13 4 9 1 9 1 9 13 2
26 9 9 1 11 11 11 11 1 11 11 11 11 7 11 11 11 11 2 11 2 1 9 9 13 4 2
23 10 9 1 11 11 1 13 16 9 1 12 9 1 9 1 15 9 13 9 0 13 4 2
18 9 1 0 9 14 9 1 15 9 13 9 0 13 10 9 13 4 2
27 11 11 1 13 16 16 11 9 9 1 13 9 1 3 14 13 4 16 9 1 15 1 9 13 4 4 2
20 15 0 13 16 2 15 14 9 1 0 9 9 1 9 9 1 14 13 4 2
23 15 1 0 3 9 15 1 0 9 1 9 1 10 13 7 15 1 9 1 14 9 13 2
17 15 13 16 9 14 13 1 10 9 14 13 7 15 9 13 4 2
31 0 9 1 9 1 9 12 9 13 1 11 11 13 4 11 11 1 13 16 9 1 9 0 9 1 13 4 14 9 13 2
26 15 9 1 9 1 9 13 7 13 16 11 11 1 10 9 1 9 1 9 1 9 1 9 13 4 2
27 11 9 11 1 13 7 0 2 0 9 1 9 1 9 1 1 11 9 1 9 1 15 9 1 9 13 2
40 12 9 0 9 7 12 9 1 9 13 1 3 11 1 13 9 1 3 0 7 3 0 9 9 9 2 11 11 2 1 9 3 11 1 11 11 1 13 4 2
15 10 9 1 9 1 13 9 1 12 9 1 0 9 13 2
12 9 1 9 11 11 1 11 11 1 13 4 2
30 9 9 1 3 0 9 1 15 9 0 13 4 10 9 1 9 1 11 1 11 11 1 9 11 1 11 11 1 13 2
26 16 12 14 9 9 1 9 9 1 9 13 4 4 7 15 1 1 9 11 16 11 11 1 13 4 2
14 9 1 1 9 1 9 1 0 9 1 13 4 4 2
14 9 1 1 9 1 3 13 4 12 9 1 0 9 2
19 11 9 9 1 9 1 3 13 1 1 11 11 1 11 1 0 9 13 2
31 9 1 9 1 9 13 4 16 15 11 1 0 9 1 9 0 13 16 10 9 1 9 13 1 1 14 0 13 4 4 2
47 9 0 9 9 11 11 7 9 11 11 11 1 9 1 11 11 11 2 11 2 1 11 9 1 12 0 9 1 9 1 1 13 2 2 9 13 1 1 9 9 13 1 9 14 13 4 4
21 9 1 9 9 9 1 9 13 4 16 15 9 1 1 0 9 9 3 9 13 2
55 9 1 9 1 1 0 9 2 9 2 11 1 9 13 16 15 9 9 1 9 13 16 15 12 9 1 1 2 11 11 1 2 0 9 1 9 0 13 7 15 9 9 9 1 13 4 16 10 9 1 0 13 4 4 2
19 9 1 10 9 1 14 9 13 4 2 15 1 9 9 1 9 0 13 2
21 9 1 13 16 0 9 1 0 13 1 9 1 0 7 0 9 13 1 9 13 2
31 15 1 14 9 1 9 1 0 9 9 11 11 11 1 13 4 16 15 11 11 1 0 7 0 9 13 1 1 9 13 2
31 9 1 1 9 11 1 13 16 9 1 12 12 10 9 0 13 2 15 1 9 9 7 9 9 1 9 0 13 4 4 2
28 11 1 9 1 9 9 0 13 1 1 9 1 9 13 2 7 9 1 15 14 11 11 1 14 9 13 4 2
21 11 1 15 9 1 9 1 1 9 1 9 7 15 9 1 1 14 9 13 4 2
35 9 9 1 1 11 11 11 2 11 11 11 2 11 2 7 11 11 11 1 9 1 1 11 1 12 7 11 1 12 9 0 13 4 4 2
19 10 9 11 2 11 11 7 11 11 1 0 9 1 1 9 13 4 4 2
42 11 11 11 2 11 2 1 9 1 1 0 9 9 1 0 13 1 9 1 1 12 9 1 0 13 1 3 9 14 1 9 1 14 12 12 9 11 1 3 13 4 2
16 7 2 9 1 10 9 1 1 9 1 9 1 9 0 13 2
18 10 2 10 9 15 9 1 13 4 2 15 14 0 9 13 13 4 2
7 15 9 14 3 0 13 2
22 10 9 1 9 11 1 1 1 9 1 1 12 1 12 9 10 9 1 13 4 4 2
16 9 1 0 0 9 1 9 14 14 12 1 12 9 10 13 2
28 9 9 10 9 1 0 13 16 15 14 0 9 1 9 1 1 9 7 0 0 9 1 1 10 9 13 4 2
16 11 11 11 1 9 3 12 9 13 15 13 12 9 13 4 2
14 11 11 1 9 14 12 9 1 13 12 9 13 4 2
13 11 11 1 14 9 12 1 13 12 9 13 4 2
24 11 11 11 1 0 9 1 13 1 1 9 0 9 13 0 9 13 1 9 1 13 4 4 2
13 0 9 1 9 7 9 1 9 13 1 9 13 2
30 11 1 14 10 9 1 15 9 13 4 4 2 7 11 9 1 3 1 9 13 4 11 7 11 1 15 9 13 4 2
33 11 11 11 1 11 1 9 1 1 2 11 9 11 11 1 13 16 9 10 9 1 9 1 9 7 9 1 9 13 1 9 13 2
24 15 10 9 9 1 13 16 15 15 9 9 1 0 13 7 3 14 3 10 9 1 8 13 2
24 7 9 1 9 9 11 1 13 16 9 1 0 9 1 0 9 1 9 9 1 0 13 4 2
14 9 1 13 16 0 9 1 0 13 1 10 9 13 2
24 11 11 11 11 11 10 9 1 9 2 9 1 1 11 1 0 2 0 9 1 9 1 13 2
36 11 1 9 1 1 1 9 0 13 4 13 16 0 7 9 9 1 9 13 4 1 13 9 1 0 9 1 0 9 1 1 13 4 4 4 2
37 11 11 11 2 11 2 2 11 7 11 1 9 1 1 13 9 1 1 11 11 11 1 1 11 11 11 11 7 0 9 11 11 11 14 0 13 2
27 9 1 1 10 9 1 14 13 16 9 9 1 1 10 9 9 1 9 12 1 12 12 1 13 4 4 2
14 15 10 0 9 1 3 14 0 13 4 1 9 13 2
24 9 1 13 16 9 1 10 9 1 0 13 16 15 0 9 1 14 9 1 9 1 9 13 2
27 9 1 11 9 1 9 11 11 1 13 7 11 1 9 1 11 11 2 11 11 11 7 11 11 0 13 2
14 9 1 1 1 11 11 11 1 1 12 9 13 4 2
16 0 9 1 9 7 9 9 1 12 9 9 13 1 9 13 2
20 0 9 1 9 1 12 9 9 7 9 9 9 1 12 9 13 1 9 13 2
21 0 9 1 9 9 7 9 9 1 12 9 9 9 1 1 0 13 1 9 13 2
24 0 9 9 9 1 13 4 4 15 10 0 9 1 1 9 9 1 12 9 9 13 0 13 2
33 9 1 9 1 9 1 3 1 1 13 1 9 1 1 11 11 9 1 9 1 9 1 9 13 7 9 13 1 9 13 4 4 2
28 11 11 11 11 11 1 13 16 0 9 1 9 1 13 11 1 13 9 7 9 9 1 9 9 9 13 4 2
31 9 1 11 1 11 11 1 0 9 1 13 13 9 1 9 9 13 4 11 1 13 16 9 15 1 1 10 0 9 13 2
16 15 10 9 15 1 9 1 13 9 1 9 14 9 1 13 2
25 15 13 16 11 1 9 1 9 1 13 9 1 1 15 1 9 1 0 9 1 12 9 0 13 2
25 15 12 9 9 1 13 7 12 9 7 12 9 9 1 1 1 13 4 7 12 12 9 0 13 2
16 11 1 13 16 9 1 9 1 9 1 13 9 13 4 4 2
8 11 1 15 13 4 0 13 2
11 15 13 16 9 9 1 10 0 9 13 2
23 9 9 1 9 11 11 1 11 1 13 16 11 1 11 1 9 1 0 9 13 4 4 2
18 15 13 4 16 11 1 0 9 10 9 1 10 9 1 9 13 4 2
18 0 9 0 9 1 9 1 11 1 9 1 0 11 1 9 13 4 2
12 10 9 1 9 1 11 11 1 13 4 4 2
17 15 1 11 11 1 0 9 1 9 1 11 1 9 1 9 13 2
36 11 11 1 9 1 9 11 9 1 0 9 1 15 9 1 13 1 14 15 14 13 2 7 15 3 13 16 11 1 11 1 9 13 4 4 2
9 15 11 11 1 9 1 9 13 2
22 0 13 16 11 9 1 0 9 1 11 1 9 13 4 16 15 11 1 14 13 4 2
25 15 11 1 11 9 9 9 1 9 1 9 7 0 9 1 9 1 14 11 1 1 9 13 4 2
15 0 9 1 10 9 1 11 1 9 1 9 13 4 4 2
21 2 11 11 2 13 9 1 9 1 9 13 1 9 1 9 1 9 9 13 4 2
20 15 1 0 9 0 9 1 9 15 9 7 0 9 1 11 1 9 13 4 2
21 7 2 9 7 9 1 1 13 4 1 9 1 11 1 9 3 1 1 0 13 2
38 11 11 11 1 9 1 13 9 1 9 1 0 9 2 11 11 11 2 9 7 0 9 7 9 1 0 9 1 9 13 1 9 1 14 9 13 4 2
20 9 1 9 9 1 0 0 9 1 9 9 1 2 9 11 2 1 13 4 2
21 15 1 9 9 9 1 11 11 11 2 11 2 1 13 13 9 0 13 13 4 2
35 9 1 9 1 1 11 11 11 11 11 11 11 11 1 9 1 13 16 9 1 0 2 11 11 11 2 11 11 1 9 1 9 13 4 2
23 0 9 1 9 7 9 1 1 13 4 1 15 14 9 1 11 1 9 14 13 4 4 2
22 10 9 9 2 9 2 9 7 9 1 9 7 15 14 9 1 11 0 13 0 13 2
24 10 9 1 11 1 9 1 0 13 4 11 1 9 1 9 1 0 9 13 1 9 13 4 2
15 15 1 1 11 1 9 1 9 1 0 9 0 13 4 2
15 15 1 14 13 4 16 10 9 1 9 1 9 13 4 2
21 11 11 1 0 9 9 1 15 9 1 11 11 11 2 11 1 0 9 13 4 2
10 11 11 11 1 15 0 13 4 4 2
25 15 1 10 9 1 1 0 9 2 0 9 7 0 9 1 11 1 9 1 9 13 4 4 4 2
21 11 11 1 13 16 9 1 0 0 9 1 0 0 11 9 1 9 13 4 4 2
12 11 1 1 10 9 13 1 11 0 9 13 2
20 15 1 0 13 4 0 9 2 9 1 1 14 0 0 9 1 0 13 4 2
37 9 14 1 13 9 1 9 13 1 9 1 1 11 11 11 11 11 11 3 14 9 1 9 1 9 13 1 1 11 2 11 11 11 11 9 13 2
40 11 1 9 9 9 9 11 11 1 13 16 15 9 14 1 9 1 1 15 9 1 9 13 1 1 9 9 1 1 3 14 11 11 11 11 11 11 9 13 2
18 11 1 13 16 9 8 8 13 4 7 9 9 9 1 1 13 4 2
11 15 1 12 9 7 12 9 9 13 4 2
12 15 1 9 1 9 9 1 9 14 13 4 2
31 15 13 16 9 15 9 9 1 13 7 9 9 1 1 9 12 9 9 1 1 9 2 9 1 1 14 9 13 4 4 2
32 11 2 11 1 13 9 1 1 1 0 13 4 2 9 2 1 9 7 9 1 9 13 4 4 16 15 9 1 9 14 13 2
24 11 7 11 1 13 10 9 11 2 11 2 11 2 11 11 2 1 9 11 1 1 1 13 2
11 15 9 14 1 11 1 0 13 4 4 2
16 15 1 11 1 9 7 11 1 9 1 9 13 1 9 13 2
18 9 1 11 7 11 9 1 9 1 9 14 13 1 1 13 4 4 2
13 15 13 4 4 16 0 9 9 11 1 14 13 2
25 15 15 14 9 13 4 4 16 15 0 9 1 15 9 13 4 7 9 1 1 15 9 13 4 2
23 15 9 9 1 9 1 13 4 7 15 13 4 4 16 10 9 1 15 0 9 13 4 2
22 9 9 7 9 1 13 1 14 9 13 4 4 7 9 13 4 1 9 13 4 4 2
18 2 11 11 2 1 11 9 1 11 1 15 12 0 9 1 9 13 2
20 9 11 11 7 15 9 11 11 1 0 9 2 9 1 1 9 1 9 13 2
26 10 9 1 0 2 11 11 2 9 1 9 1 1 11 2 11 1 0 9 1 14 9 1 9 13 2
14 11 2 2 11 11 2 1 9 9 1 0 9 13 2
19 11 11 11 1 11 1 9 13 9 9 1 10 9 10 9 0 13 4 2
37 11 1 1 11 11 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 7 11 1 14 9 0 13 4 2
22 9 9 9 1 12 12 1 10 9 1 9 10 9 2 11 11 2 1 9 13 4 2
16 15 1 11 1 2 11 11 2 1 9 11 1 13 13 4 2
21 10 0 9 1 1 14 12 9 1 14 10 9 11 1 3 0 9 13 4 4 2
20 0 9 9 1 0 9 14 15 10 9 1 3 10 9 1 9 0 13 4 2
34 9 11 11 1 1 11 1 9 9 13 1 3 2 11 11 2 15 0 3 9 13 1 3 14 1 0 3 9 1 9 1 14 13 2
21 15 15 13 9 13 4 4 16 12 10 9 14 13 15 9 1 9 0 13 4 2
18 15 10 9 13 16 3 1 10 10 9 14 10 9 1 13 4 4 2
17 10 9 7 10 9 1 2 10 9 2 10 15 1 13 4 4 2
14 15 9 1 13 1 10 9 1 9 1 9 13 4 2
17 16 15 1 9 1 9 13 16 15 14 9 1 13 1 14 13 2
22 9 13 2 9 9 13 4 2 9 7 9 9 2 15 14 0 13 2 13 4 4 2
15 10 9 1 12 2 12 9 1 9 15 9 1 13 4 2
13 0 9 9 1 14 0 2 0 9 1 13 4 2
15 9 9 1 1 9 2 9 1 10 10 9 13 4 4 2
9 11 9 1 1 9 9 13 4 2
17 11 2 11 9 1 11 1 12 9 1 11 1 1 11 9 13 2
12 15 1 13 9 9 1 14 9 11 9 13 2
16 10 9 1 13 14 9 2 9 7 9 1 9 13 4 4 2
8 10 9 1 0 9 9 13 2
15 9 9 1 9 9 13 1 1 15 9 9 11 9 13 2
16 14 12 9 1 15 1 9 9 1 13 1 9 1 0 13 2
14 15 9 1 13 1 10 9 1 9 1 0 13 4 2
11 15 10 0 9 1 10 9 1 13 4 2
13 15 15 0 9 1 1 15 9 2 9 14 13 2
17 9 1 14 13 2 15 9 1 1 15 14 9 9 14 13 4 2
23 9 9 11 11 11 1 1 11 1 1 11 1 14 10 9 1 9 1 9 13 4 4 2
18 11 2 11 7 11 9 1 0 9 1 10 9 1 1 9 13 4 2
12 9 9 10 9 1 9 13 1 9 1 13 2
18 12 9 1 1 11 11 9 9 13 11 11 11 11 9 1 11 13 2
17 15 13 4 16 3 9 14 9 9 13 3 9 13 0 13 4 2
24 9 1 11 11 11 11 11 1 9 1 11 1 12 0 9 1 9 1 9 9 13 4 4 2
34 0 3 11 11 11 11 11 11 1 11 11 11 1 9 1 11 1 12 10 9 9 9 11 11 11 1 9 9 1 9 0 13 4 2
18 11 1 11 1 9 9 11 11 1 9 1 0 9 1 0 13 4 2
25 11 1 11 1 10 0 9 1 9 9 0 13 15 12 9 1 9 9 1 11 9 1 13 4 2
20 11 1 15 9 11 13 4 4 4 4 2 15 15 0 9 1 0 13 4 2
19 11 1 15 11 0 0 9 1 11 1 8 0 9 1 0 13 4 4 2
12 15 1 9 7 9 1 12 0 9 0 13 2
15 11 9 15 1 12 0 2 0 9 9 0 13 4 4 2
36 0 3 12 9 1 9 1 9 13 4 11 11 11 11 11 11 11 1 9 11 11 11 11 11 11 1 11 11 11 1 9 1 9 13 4 2
14 15 1 11 1 9 0 13 15 11 1 1 13 4 2
21 11 1 11 1 11 1 9 1 10 14 9 1 15 9 11 1 1 13 4 4 2
14 11 0 9 1 11 9 1 9 13 1 0 9 13 2
19 15 1 11 11 11 1 11 11 7 11 9 11 11 14 9 13 4 4 2
46 11 1 9 1 11 11 1 11 2 15 9 7 11 1 11 9 11 11 2 11 9 1 9 11 11 2 9 9 11 11 7 11 9 11 11 1 1 0 2 0 9 9 0 13 4 2
18 11 1 15 9 11 11 1 0 9 1 9 9 1 13 1 9 13 2
22 0 14 9 11 11 1 15 9 1 9 1 9 0 13 4 2 15 0 13 4 4 2
36 0 13 16 11 11 1 15 9 9 11 1 9 1 1 10 9 0 13 4 4 2 15 15 9 2 9 1 9 7 9 13 3 13 4 4 2
32 0 2 0 9 0 13 1 12 9 1 9 1 11 1 9 1 1 11 1 15 9 1 9 13 4 7 0 9 9 14 13 2
26 11 11 1 11 11 11 1 11 7 11 1 0 0 9 1 13 15 11 1 9 1 3 13 4 4 2
36 10 9 9 1 11 2 11 11 11 1 0 9 1 12 9 1 13 4 1 11 1 15 9 1 2 0 9 2 9 13 1 3 13 4 4 2
21 0 9 1 13 16 11 11 11 1 0 10 9 1 15 9 0 14 13 4 4 2
29 16 15 13 4 4 4 16 11 1 9 3 13 1 3 11 11 1 9 1 9 1 9 13 1 15 0 13 4 2
27 10 9 1 9 1 12 9 1 9 13 4 11 11 11 2 11 2 1 9 7 15 9 1 9 13 4 2
31 9 1 13 13 16 9 1 0 0 9 1 9 13 1 3 11 10 9 1 9 13 1 1 3 10 9 0 13 13 4 2
15 11 1 15 9 9 13 4 15 2 0 9 2 13 4 2
26 15 9 1 9 13 4 4 7 15 13 4 16 9 9 13 1 3 10 9 1 9 13 1 9 13 2
19 15 13 16 15 1 11 1 9 1 12 9 1 11 1 9 13 4 4 2
15 7 15 11 1 0 9 2 9 1 1 9 0 13 4 2
29 11 1 9 11 1 9 1 9 0 9 11 1 9 13 4 7 15 0 9 1 0 13 1 9 13 4 4 4 2
12 11 1 0 9 1 9 1 1 13 4 4 2
47 9 9 9 11 11 1 11 11 11 1 0 9 11 11 11 2 11 11 11 1 9 11 11 11 7 11 9 11 11 11 1 1 10 9 1 3 10 9 13 1 3 10 9 13 4 4 2
42 11 9 11 11 1 1 0 9 1 9 1 9 0 13 4 11 1 11 11 11 1 13 16 10 9 9 1 9 14 13 4 2 15 0 9 1 9 13 1 13 4 2
26 11 1 11 1 9 1 15 12 0 9 1 13 16 0 9 1 15 9 1 1 1 9 14 13 4 2
49 11 1 11 2 11 9 11 11 7 11 9 11 11 1 0 9 1 9 9 9 9 13 4 11 1 9 13 16 11 1 15 9 9 13 1 1 9 1 9 1 9 13 4 2 15 11 9 13 2
25 11 1 11 1 9 13 16 11 1 11 2 11 1 12 9 1 9 1 1 9 9 13 4 4 2
24 9 1 9 1 9 1 9 13 7 0 9 1 12 9 1 9 1 1 1 9 13 4 4 2
32 11 9 1 11 11 1 13 1 9 9 1 1 11 1 11 9 9 11 11 11 7 0 9 1 9 1 9 1 9 1 13 2
32 11 11 7 11 11 11 11 2 11 2 1 9 1 11 11 1 11 11 1 11 1 12 9 1 13 1 9 1 9 13 4 2
18 9 1 11 1 0 11 11 11 1 9 1 0 9 13 1 9 13 2
42 11 9 1 11 11 1 9 9 9 2 11 2 0 13 9 1 11 11 1 9 1 9 13 4 13 4 16 9 11 7 11 1 11 11 1 9 1 0 9 13 4 2
7 15 13 4 3 0 13 2
29 11 1 13 4 4 16 11 7 11 1 9 1 1 10 9 3 13 4 16 9 11 1 10 3 1 13 4 4 2
15 11 1 1 9 1 9 1 9 2 9 2 13 4 4 2
25 11 7 11 10 9 11 1 0 9 9 1 13 2 15 15 0 9 1 1 9 1 13 4 4 2
12 9 1 14 0 9 11 1 13 1 9 13 2
27 11 1 9 1 13 4 16 11 11 1 9 9 1 0 13 4 11 11 1 11 1 11 1 9 13 4 2
18 15 11 11 9 1 0 12 9 1 9 1 9 1 1 13 4 4 2
16 16 12 9 1 0 9 9 1 11 7 11 1 9 14 13 2
27 7 15 11 10 9 1 9 1 9 13 4 4 15 9 13 16 9 1 11 11 9 1 0 9 13 4 2
16 11 11 1 9 0 11 1 11 1 10 9 1 0 9 13 2
18 15 10 0 11 13 15 11 1 9 1 13 1 3 9 13 4 4 2
29 11 1 9 1 13 16 11 11 11 1 11 1 11 1 10 12 9 13 2 15 0 3 11 1 14 9 13 4 2
40 15 0 11 1 1 11 14 11 2 11 14 11 2 11 14 11 2 11 14 11 2 11 14 11 2 11 14 11 2 11 14 11 7 9 11 14 11 0 13 2
51 0 9 11 1 9 1 1 1 11 1 13 4 16 11 1 11 11 11 1 11 11 1 9 1 1 15 10 9 0 13 4 15 10 9 1 11 2 11 7 11 1 11 1 9 13 1 0 9 13 4 2
17 11 11 11 11 2 11 2 9 11 11 1 15 9 13 4 4 2
33 15 13 16 16 9 12 0 9 2 11 2 1 15 0 9 1 13 1 0 14 13 16 3 15 0 9 11 1 0 9 13 4 2
39 11 11 1 15 9 0 13 4 11 11 11 11 1 9 9 11 1 15 11 1 9 9 1 13 16 11 1 0 9 1 1 1 0 13 9 1 9 13 2
11 15 11 1 9 1 13 1 0 9 13 2
13 11 1 9 1 11 11 2 11 2 1 9 13 2
10 15 1 11 1 9 9 9 9 13 2
19 15 13 16 16 11 7 11 0 9 13 4 4 16 11 15 14 13 4 2
26 15 13 16 0 9 11 1 11 1 11 11 1 11 1 9 13 4 4 7 15 9 1 13 4 4 2
19 16 11 7 9 9 15 9 14 13 4 16 0 13 16 15 11 1 13 2
32 0 13 16 11 11 1 11 11 1 11 11 11 1 9 1 13 4 16 11 9 1 9 0 13 1 3 14 15 0 9 13 2
19 0 13 16 11 1 11 11 1 9 1 1 11 11 1 9 1 13 4 2
8 11 1 9 11 1 13 4 2
16 10 9 10 9 7 11 1 9 9 11 11 1 1 13 4 2
23 10 9 1 13 4 4 11 1 0 11 11 7 10 0 9 11 11 1 9 11 11 11 2
29 11 1 9 13 16 11 11 1 14 0 13 16 10 9 10 0 9 1 13 2 7 15 9 1 9 13 4 4 2
31 11 11 11 1 13 16 15 11 1 10 0 9 1 1 1 9 13 4 4 2 15 11 1 9 1 9 11 1 13 4 2
15 16 11 11 3 2 3 0 13 4 16 15 15 9 13 2
17 15 13 16 9 13 1 15 10 0 9 1 9 1 9 13 4 2
28 15 9 13 16 15 0 9 15 10 9 1 10 9 1 9 13 4 15 11 11 1 10 9 1 9 13 4 2
12 11 11 10 9 1 9 1 9 13 14 13 2
20 15 13 16 11 1 15 9 9 1 13 4 7 10 0 9 1 9 13 4 2
15 15 13 16 9 1 10 9 1 9 1 0 9 13 4 2
18 11 1 13 16 0 9 1 10 9 1 9 1 9 13 1 9 13 2
40 3 15 9 1 0 9 13 1 13 4 7 9 1 9 13 4 16 10 9 15 13 2 15 11 1 9 1 0 9 12 12 9 1 15 9 1 13 4 4 2
31 9 14 1 11 1 9 13 4 16 0 9 1 0 9 1 15 9 1 12 12 9 1 11 2 11 9 1 9 13 4 2
13 15 9 13 4 16 10 9 11 1 13 4 4 2
16 11 1 9 13 16 10 0 9 15 14 11 1 13 4 4 2
11 15 0 9 1 0 9 1 0 13 4 2
15 0 13 16 11 11 11 1 9 1 0 9 13 4 4 2
22 15 13 16 10 9 1 15 10 9 13 4 2 15 9 0 9 1 9 1 13 4 2
21 3 10 9 13 16 11 11 1 10 9 1 9 1 9 13 1 9 13 4 4 2
24 11 1 0 9 11 11 1 9 1 1 11 11 1 11 1 15 11 11 11 1 1 0 13 2
17 9 1 15 0 9 1 9 0 12 9 10 13 1 9 13 4 2
26 11 11 11 1 11 1 9 13 1 12 9 1 11 11 1 12 9 1 1 0 9 1 13 4 4 2
19 15 1 11 9 1 11 1 9 9 9 11 11 11 1 1 0 13 4 2
16 15 9 1 15 9 1 9 11 11 1 13 1 9 0 13 2
35 9 1 9 1 13 16 11 1 15 9 14 13 4 2 7 9 9 1 9 1 1 9 1 9 1 15 0 13 1 15 1 0 9 13 2
40 9 1 9 11 11 11 1 1 9 9 11 1 1 1 9 14 13 1 1 1 3 1 9 1 1 9 1 13 1 1 12 9 9 13 1 9 13 4 4 2
48 11 1 0 9 1 9 1 3 13 7 11 1 9 9 9 1 9 13 1 9 1 0 13 1 9 13 4 9 11 11 1 13 16 0 9 1 15 15 9 1 2 9 2 13 4 4 4 2
22 15 9 1 9 13 4 16 15 9 7 10 9 1 0 9 1 9 13 0 13 4 2
46 11 1 11 11 11 1 9 11 11 1 12 9 1 0 13 4 11 1 13 16 11 11 1 9 13 2 11 1 9 9 9 1 9 13 7 9 9 13 1 9 1 0 13 4 4 2
35 15 13 16 15 0 9 1 9 1 3 13 4 4 7 0 9 15 9 1 9 13 4 4 7 0 9 1 15 15 9 13 4 4 4 2
25 11 1 13 16 9 1 15 9 1 9 1 9 13 4 4 4 2 15 15 15 1 13 4 4 2
16 13 1 14 9 13 7 15 13 4 4 15 14 9 14 13 2
30 15 0 9 1 9 13 16 15 10 9 1 9 13 7 0 9 7 9 1 9 13 1 9 1 9 13 0 13 4 2
41 2 11 11 2 1 0 9 1 15 15 13 4 0 13 4 4 16 3 15 9 2 9 7 9 1 9 1 9 13 1 9 7 9 1 9 14 13 1 9 13 2
18 15 15 9 14 13 7 9 1 9 13 1 15 9 1 9 14 13 2
18 11 11 11 2 11 2 1 9 11 11 1 9 1 3 13 4 4 2
24 11 1 13 4 16 11 11 10 9 1 11 1 1 13 4 9 1 1 9 0 13 4 4 2
14 7 9 1 3 0 13 4 1 15 3 9 13 4 2
18 9 1 13 13 16 11 11 1 9 1 11 9 1 0 13 0 13 2
11 9 15 11 1 9 1 9 13 4 4 2
16 11 1 9 13 4 16 9 11 9 1 13 4 13 4 4 2
16 12 9 1 9 1 10 9 1 12 9 13 4 4 4 4 2
15 0 3 11 11 1 12 9 0 9 1 1 13 4 4 2
10 11 9 1 9 13 4 13 4 4 2
16 11 1 9 10 9 1 9 9 1 1 1 13 4 4 4 2
21 11 1 13 4 16 11 9 1 9 0 9 1 10 7 9 1 9 1 10 13 2
19 11 9 11 11 11 1 11 9 1 11 11 1 9 1 9 0 13 4 2
19 15 13 16 9 1 9 13 11 9 0 9 1 13 1 9 13 4 4 2
14 15 13 16 9 1 10 9 9 1 1 13 4 4 2
27 15 13 16 11 2 11 7 11 1 9 1 9 13 1 9 3 14 11 1 9 1 0 9 1 9 13 2
31 11 11 1 11 11 11 1 9 1 9 13 1 12 0 9 9 9 11 7 11 2 11 1 9 1 11 1 0 13 4 2
27 9 9 1 15 9 1 12 9 1 9 9 9 1 15 9 1 13 4 9 1 9 9 13 1 13 4 2
22 11 11 1 13 13 16 9 1 15 13 1 0 9 13 16 15 15 9 13 4 4 2
62 11 11 11 7 11 11 2 11 11 11 11 1 1 1 0 0 9 9 1 0 13 4 9 9 11 11 11 2 9 11 11 11 7 11 11 11 1 9 1 12 9 1 9 9 1 9 13 1 13 16 15 10 9 1 15 9 1 9 13 4 4 2
18 15 1 14 11 11 1 9 9 1 9 1 12 9 1 13 4 4 2
45 12 9 1 1 1 15 9 0 9 11 11 7 11 11 1 15 13 16 9 1 15 0 13 4 4 4 2 9 1 9 1 10 9 13 4 4 7 15 0 9 1 3 10 13 2
22 15 1 9 1 13 16 15 14 9 9 14 13 16 9 1 9 10 9 1 13 4 2
39 9 9 1 9 1 11 11 1 10 12 9 7 0 10 9 9 9 1 9 7 9 1 9 7 9 1 9 1 9 7 15 9 1 9 13 1 13 4 2
31 11 11 1 13 13 16 9 9 1 1 13 4 9 9 1 13 7 15 9 9 1 10 9 0 7 0 9 14 13 4 2
15 9 1 12 9 1 11 11 11 1 9 13 1 13 4 2
38 9 1 13 13 16 16 15 1 9 1 9 13 4 1 9 1 9 1 0 15 9 1 9 14 13 4 4 2 16 15 11 11 1 9 13 4 4 2
19 15 13 16 9 9 1 9 13 1 9 7 9 1 9 1 9 13 4 2
24 15 15 9 1 13 16 9 1 9 1 0 9 9 1 9 1 0 9 1 9 1 9 13 2
30 9 1 9 1 13 16 15 15 9 1 13 4 4 16 9 9 1 9 13 4 9 1 9 1 9 1 9 13 4 2
11 11 11 11 0 9 1 9 1 11 13 2
18 15 1 12 9 15 3 0 9 1 9 15 2 15 1 9 1 13 2
28 11 1 0 9 11 11 11 1 11 1 11 1 13 16 11 11 11 0 9 1 9 1 11 13 1 0 13 2
36 11 1 9 9 11 11 11 11 1 1 9 1 9 1 1 13 16 11 11 1 12 9 1 11 1 13 1 1 9 13 1 9 13 4 4 2
34 11 1 9 1 0 11 9 1 9 13 11 1 11 11 11 1 14 11 1 9 13 11 11 11 13 1 1 1 14 9 2 9 13 2
11 11 11 1 3 14 15 9 13 13 4 2
23 11 1 13 16 11 1 0 9 13 4 1 1 11 11 1 9 1 10 9 13 4 4 2
10 7 15 1 15 9 14 13 4 4 2
14 3 11 10 9 1 1 11 0 11 11 13 4 4 2
20 16 15 13 16 11 9 1 13 14 0 9 1 13 1 0 9 14 0 13 2
15 15 13 16 0 9 14 9 9 1 3 13 1 0 13 2
38 11 7 11 11 1 11 1 12 9 1 1 11 11 11 2 11 2 1 9 1 0 9 9 9 7 0 0 9 1 9 1 9 1 9 2 9 13 2
28 9 1 12 0 0 9 1 11 11 11 11 7 11 11 11 1 9 1 12 9 9 0 13 1 9 13 4 2
38 15 1 14 12 9 1 11 11 1 11 11 11 1 11 11 1 9 13 4 11 11 1 0 9 9 9 1 9 1 1 0 9 13 1 14 9 13 2
45 11 11 11 11 11 11 7 11 11 1 11 11 11 11 11 1 0 9 1 0 9 1 9 1 12 9 1 9 9 7 0 0 9 1 9 1 9 1 9 1 9 2 9 13 2
36 9 1 1 12 9 1 0 9 1 9 13 1 1 11 7 11 11 1 1 11 11 11 2 11 2 1 3 0 13 1 9 1 14 9 13 2
28 9 1 11 1 9 13 4 13 16 11 7 11 11 1 1 11 11 9 1 13 10 9 1 9 1 9 13 2
50 15 9 13 4 13 16 11 11 11 2 11 1 0 9 1 9 1 0 13 2 15 1 9 1 9 1 0 9 1 0 9 1 1 1 0 13 4 4 7 11 11 10 9 1 11 1 1 9 13 2
24 0 9 1 9 13 1 1 11 11 11 1 11 1 9 1 0 13 4 1 9 1 9 13 2
13 15 1 11 1 0 0 0 9 1 9 9 13 2
33 10 9 1 9 9 11 11 11 1 13 16 9 1 10 9 1 0 9 1 13 4 4 1 3 14 9 1 9 1 9 13 4 2
23 0 9 1 0 13 1 9 12 9 1 0 13 7 10 9 1 12 12 9 1 9 13 2
29 10 9 1 9 9 1 11 11 11 1 13 16 9 9 1 9 1 10 9 1 15 10 9 1 9 13 4 4 2
16 10 0 9 1 9 1 9 9 1 9 1 13 4 4 4 2
17 7 0 9 10 9 1 0 9 1 9 13 1 0 14 13 4 2
20 10 9 1 9 9 11 11 11 7 11 11 11 11 11 11 11 11 0 13 2
18 10 9 1 9 11 11 11 1 9 11 11 11 1 12 9 13 13 2
14 9 11 1 9 1 14 10 9 1 9 13 4 4 2
14 11 7 11 1 13 0 9 1 11 9 9 1 13 2
20 15 9 3 13 4 4 7 15 1 14 11 1 9 1 9 13 4 4 4 2
17 9 1 9 1 11 9 1 13 9 9 1 9 0 13 4 4 2
12 9 1 10 9 1 9 1 9 13 4 4 2
11 11 9 1 12 9 14 0 13 4 4 2
27 11 1 11 11 11 1 9 1 9 1 13 9 1 1 12 9 1 14 13 4 4 2 7 12 0 13 2
15 11 9 9 1 13 12 9 1 14 9 14 13 4 4 2
18 9 1 9 1 1 1 11 11 1 12 9 1 13 4 1 9 13 2
10 11 11 1 11 7 11 9 1 13 2
21 11 9 1 9 1 12 9 9 2 9 2 9 2 9 1 9 0 13 4 4 2
29 11 9 13 9 11 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 14 12 9 1 9 13 4 4 2
30 11 11 11 1 11 7 11 11 1 9 11 11 7 15 9 11 2 11 7 12 0 9 11 9 9 1 13 4 4 2
8 15 1 1 15 9 14 13 2
38 11 1 12 9 11 2 11 7 11 11 9 1 9 1 9 13 1 1 9 11 11 1 1 13 4 4 16 9 1 10 9 13 1 1 1 13 4 2
25 9 1 11 7 11 1 3 13 4 7 0 9 1 13 1 12 0 11 1 10 9 14 13 4 2
31 9 11 11 11 1 9 11 2 11 2 11 2 11 2 11 7 11 11 1 13 16 9 1 1 9 1 0 9 13 4 2
11 11 11 1 0 9 1 14 9 13 4 2
12 15 9 1 9 1 14 12 9 1 9 13 2
22 9 13 7 9 13 1 0 7 0 11 11 7 11 11 11 1 0 13 4 4 4 2
14 11 11 1 9 1 11 9 1 1 13 4 4 4 2
30 9 1 10 9 1 9 13 1 11 11 11 11 11 1 12 9 9 9 9 1 12 9 9 1 9 0 13 4 4 2
15 11 9 1 9 1 11 11 1 10 9 0 13 4 4 2
30 11 11 11 1 11 1 13 16 0 9 1 9 1 9 1 9 13 1 1 9 9 1 2 9 1 2 9 13 4 2
15 15 15 14 13 16 0 9 1 9 1 13 14 4 4 2
17 11 1 9 1 9 13 4 13 16 9 9 9 1 10 0 13 2
29 11 1 13 0 9 1 1 11 1 11 1 9 13 16 15 0 9 1 15 9 1 11 0 9 1 9 14 13 2
17 15 13 16 9 1 13 1 1 11 11 1 12 0 9 13 4 2
27 13 9 1 11 11 1 13 16 10 9 0 14 13 7 9 9 1 9 13 1 9 1 9 13 4 4 2
28 15 13 16 9 1 13 9 7 9 1 9 1 9 1 1 9 13 4 7 3 14 15 1 9 13 4 4 2
34 11 9 1 9 13 4 11 11 1 9 13 1 9 1 0 13 4 11 1 13 16 15 9 9 13 1 9 1 9 14 13 4 4 2
20 12 9 1 9 1 11 13 11 11 11 15 12 9 9 1 0 13 4 4 2
24 0 9 1 9 1 9 1 15 13 16 9 9 10 9 1 2 9 1 2 9 13 4 4 2
28 11 1 13 16 10 9 1 15 11 11 11 11 11 1 9 1 9 9 1 0 9 1 9 13 1 13 4 2
30 9 9 1 9 1 9 1 9 1 11 1 13 16 15 15 14 14 13 4 2 16 15 15 0 9 13 4 4 4 2
28 11 1 9 1 13 0 9 1 1 11 1 13 16 10 0 9 1 11 1 9 13 1 9 1 15 0 13 2
17 11 1 13 16 15 0 9 1 10 9 11 1 9 1 13 4 2
27 15 13 16 15 9 13 16 15 14 0 9 9 15 9 1 10 9 1 9 1 9 13 1 9 14 13 2
27 11 11 1 9 13 1 9 1 0 13 4 11 1 13 16 12 9 1 9 1 9 15 9 14 13 4 2
11 9 1 12 9 9 13 1 9 13 4 2
17 7 10 9 1 15 9 14 13 16 15 1 14 9 9 13 4 2
17 15 13 15 13 0 13 16 9 9 1 9 1 9 13 4 4 2
20 11 11 1 13 16 11 11 1 9 1 11 9 1 11 1 0 9 13 4 2
15 15 10 9 1 0 13 16 15 9 1 12 9 9 13 2
29 11 11 1 9 9 1 13 1 0 9 9 1 11 1 11 1 13 1 1 0 12 0 9 11 1 0 13 4 2
24 10 9 11 1 11 1 11 7 11 1 1 9 13 4 0 9 1 1 9 13 4 4 4 2
28 11 11 1 9 1 1 11 9 11 1 1 12 9 9 13 4 1 1 11 1 11 13 1 9 0 13 4 2
11 15 0 9 9 11 1 11 14 13 4 2
18 3 2 11 1 11 1 1 13 4 1 12 0 9 1 0 13 4 2
24 15 13 16 11 2 11 11 0 13 1 3 9 1 0 9 1 14 13 14 9 13 4 4 2
14 0 9 9 1 11 13 1 13 9 1 9 13 4 2
24 0 9 9 1 11 9 1 1 11 11 11 1 13 4 12 9 1 1 12 0 13 4 4 2
14 14 12 12 9 14 11 2 11 7 11 1 13 4 2
35 11 1 11 11 11 2 11 2 11 11 11 1 13 16 11 1 11 1 1 9 13 1 11 1 9 13 1 1 0 9 1 0 13 4 2
23 11 1 1 11 1 11 2 11 11 11 1 14 13 4 1 3 2 0 2 9 13 4 2
36 12 0 9 1 1 11 9 11 1 1 11 11 7 11 9 1 1 12 9 9 1 9 1 13 4 1 1 11 2 11 9 0 13 4 4 2
16 10 9 1 12 9 1 9 13 4 7 12 9 0 13 4 2
17 9 1 9 7 9 1 13 1 1 10 9 1 9 13 4 4 2
23 0 13 16 11 11 1 0 9 1 9 1 1 11 7 11 9 9 1 0 9 13 4 2
9 15 1 0 9 9 13 4 4 2
20 9 9 1 9 1 1 11 11 11 1 15 9 1 0 9 1 9 13 4 2
16 9 9 11 11 11 1 11 1 12 0 0 0 9 0 13 2
15 15 12 0 9 1 1 12 9 1 14 9 13 4 4 2
12 12 9 0 9 7 9 1 14 9 13 4 2
21 0 11 9 11 11 2 11 11 7 11 11 11 1 9 1 9 9 13 4 4 2
13 3 11 11 7 11 11 1 9 9 13 4 4 2
11 11 11 1 11 11 1 9 13 4 4 2
35 0 11 9 7 0 0 9 11 11 1 11 1 9 0 13 4 13 16 9 1 10 9 1 10 9 1 9 1 0 9 1 9 13 4 2
18 0 11 11 11 11 1 9 11 11 1 9 9 1 9 13 4 4 2
19 11 11 1 9 11 11 11 1 9 7 9 9 1 9 0 13 4 4 2
15 11 11 1 9 9 1 13 9 1 9 1 13 4 4 2
11 11 11 9 1 9 1 9 1 3 13 2
14 11 1 0 9 7 0 9 9 1 3 0 13 4 2
14 0 0 9 11 11 1 11 11 1 9 13 4 4 2
10 3 11 11 1 9 1 9 13 4 2
12 11 1 11 11 1 0 9 0 13 4 4 2
13 11 1 9 1 10 9 1 0 9 0 13 4 2
16 3 9 9 11 11 1 9 11 9 9 1 13 4 4 4 2
14 11 11 11 1 9 9 1 0 9 13 4 4 4 2
38 0 9 1 11 11 1 1 11 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 7 11 11 13 2
32 3 0 9 9 1 15 1 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 7 11 11 1 14 0 13 4 4 2
29 12 11 9 1 9 1 9 9 1 12 9 1 0 9 1 9 13 4 11 1 9 9 1 12 0 9 0 13 2
17 10 9 1 15 0 11 11 1 11 11 11 11 11 1 1 13 2
36 11 9 9 1 9 12 1 12 13 1 13 9 1 15 0 9 13 1 1 12 11 2 11 11 11 2 1 9 1 15 12 9 1 9 13 2
13 15 0 9 1 1 9 13 1 14 9 0 13 2
14 7 9 1 1 1 3 15 9 13 1 9 13 4 2
46 10 9 1 1 11 2 11 2 9 11 11 1 15 9 1 13 16 0 9 1 12 9 1 12 9 0 13 4 15 1 11 11 1 11 11 11 11 1 9 1 9 2 9 13 4 2
22 10 9 1 3 12 11 1 9 1 1 14 9 13 7 0 13 1 1 0 13 4 2
21 11 1 9 7 9 9 1 9 1 1 1 15 9 1 9 13 1 9 13 4 2
35 16 11 1 1 2 9 0 11 1 9 1 14 15 14 0 13 16 0 9 9 10 9 1 9 13 7 14 15 9 1 12 9 14 13 2
22 11 1 13 16 10 9 1 9 13 1 1 10 11 1 9 1 9 11 11 1 13 2
38 9 1 11 11 1 9 11 1 1 2 11 1 11 11 2 11 1 11 11 2 11 1 11 11 2 11 1 11 11 7 11 1 11 11 11 0 13 2
29 11 11 1 0 9 1 9 2 11 2 1 9 1 0 9 1 9 9 2 9 2 1 9 13 1 9 13 4 2
15 7 15 1 3 9 1 9 13 1 12 9 0 13 4 2
17 0 9 1 13 16 11 11 11 1 0 9 1 12 9 13 4 2
9 9 10 9 1 0 9 9 13 2
30 16 15 13 16 0 9 1 9 9 1 9 1 14 10 11 1 0 13 4 15 14 13 4 9 1 13 1 0 13 2
15 16 9 10 9 1 1 15 0 9 0 14 13 4 4 2
47 9 10 9 0 11 14 11 11 2 11 11 11 11 11 2 11 11 11 7 11 11 11 11 11 1 9 9 1 0 9 1 9 14 13 1 11 11 1 9 1 13 1 9 13 4 4 2
26 9 1 13 16 12 0 9 1 11 9 1 9 1 9 1 9 9 1 1 11 9 1 13 4 4 2
35 11 1 11 11 11 1 10 9 0 13 16 11 1 0 0 12 9 9 1 9 1 11 11 11 11 11 11 1 0 9 11 1 13 4 2
46 0 13 16 9 11 1 0 11 11 11 11 1 9 9 1 9 1 1 11 11 1 13 4 7 11 1 13 4 10 9 1 1 11 11 11 1 9 11 1 12 9 9 0 13 4 2
28 9 1 12 0 9 1 9 1 15 0 9 9 13 1 1 13 1 9 13 4 15 9 1 1 13 4 4 2
28 11 1 10 0 9 1 9 1 1 0 9 11 11 11 1 13 16 11 11 1 0 0 9 1 9 13 4 2
29 11 1 10 9 1 3 0 13 4 9 1 13 16 15 9 9 1 11 1 9 1 10 9 1 0 9 13 4 2
24 15 13 16 15 14 0 9 1 9 1 9 7 15 9 1 13 1 9 13 9 1 1 13 2
21 15 11 11 11 1 10 9 1 0 9 1 1 11 11 11 1 9 0 13 4 2
30 11 11 11 11 11 11 1 13 16 0 11 11 11 1 9 9 13 1 9 13 1 9 1 9 9 1 15 9 13 2
23 15 9 0 12 9 9 1 9 9 0 11 11 11 1 11 1 0 12 9 1 0 13 2
23 11 1 13 16 15 13 4 16 11 1 11 11 1 11 13 9 9 13 1 9 13 4 2
14 7 9 10 9 1 9 13 1 3 14 15 9 13 2
15 15 10 0 9 0 11 2 11 11 1 0 13 9 13 2
14 15 9 1 1 11 11 1 9 1 0 9 13 4 2
14 0 9 15 10 0 9 1 9 1 9 1 0 13 2
20 12 0 11 11 1 9 1 9 1 9 13 7 10 9 15 12 9 1 13 2
29 0 9 10 9 1 1 13 4 4 4 15 11 1 9 9 13 11 11 11 13 4 4 7 15 3 11 14 13 2
7 0 9 0 13 4 4 2
14 10 9 1 9 1 9 1 9 14 13 4 4 4 2
10 9 1 9 2 9 13 4 4 4 2
14 15 1 14 9 1 9 7 9 14 13 4 4 4 2
22 9 1 0 9 13 4 4 7 10 9 1 9 1 13 1 14 0 9 13 4 4 2
27 11 11 1 9 1 9 1 9 13 4 10 9 1 9 13 4 13 16 15 15 1 0 9 13 4 4 2
15 15 9 15 12 9 1 1 12 9 1 9 13 4 4 2
23 11 1 15 15 9 1 9 13 1 9 13 15 11 1 0 9 1 1 12 9 9 13 2
18 11 1 13 16 15 15 9 11 1 9 1 15 9 14 13 13 4 2
24 11 13 4 16 9 1 15 9 11 11 11 1 9 11 11 9 1 9 1 11 13 4 4 2
9 15 9 9 1 9 13 4 4 2
13 11 1 9 1 11 11 11 1 11 13 13 4 2
12 15 11 1 9 11 11 11 1 13 4 4 2
12 11 1 9 1 1 15 9 11 0 14 13 2
11 11 1 0 2 9 1 10 9 0 13 2
14 11 1 13 16 15 0 9 15 9 7 9 1 13 2
11 10 9 1 9 13 15 0 13 4 4 2
20 11 11 11 11 1 13 4 16 11 9 11 11 1 0 13 1 1 0 13 2
16 15 13 16 10 9 9 1 11 11 11 1 12 9 14 13 2
21 11 11 1 0 11 9 1 9 1 13 7 0 9 1 9 1 1 0 13 4 2
26 11 11 1 9 1 9 1 11 11 1 13 16 11 11 0 13 1 1 15 15 9 9 0 14 13 2
15 15 13 16 9 1 9 1 1 10 9 1 0 13 4 2
14 11 11 11 1 9 1 9 1 0 13 11 13 4 2
38 11 1 9 9 1 11 1 9 1 1 1 13 4 9 1 9 1 11 1 13 16 15 1 11 11 11 11 1 15 1 9 1 1 10 9 13 4 2
21 10 9 1 11 11 11 9 13 7 3 1 10 9 1 9 13 4 1 9 13 2
12 15 1 0 9 9 7 9 1 9 13 4 2
26 11 11 1 9 1 11 11 1 9 7 11 11 1 9 1 1 1 2 15 9 13 4 0 14 13 2
23 15 15 9 14 13 16 11 11 1 0 9 1 11 1 9 7 9 1 9 13 4 4 2
23 11 1 10 9 9 9 13 4 2 15 1 10 9 14 13 16 0 9 10 9 1 13 2
12 16 2 0 9 10 9 1 0 9 14 13 2
38 16 2 15 14 9 1 9 7 9 1 9 1 13 4 1 9 1 1 1 9 13 2 15 10 9 1 9 14 13 4 16 9 9 1 0 14 13 2
11 11 1 9 9 7 9 1 0 9 13 2
12 7 2 15 9 1 9 15 15 1 0 13 2
18 14 9 1 1 15 0 14 13 16 15 15 9 1 9 1 13 13 2
28 11 11 1 9 1 9 1 1 0 13 7 9 1 9 1 11 11 1 1 9 13 1 15 14 0 14 13 2
17 9 1 9 1 9 1 10 14 10 12 9 1 9 13 4 4 2
17 7 2 9 1 11 1 9 1 10 14 10 12 9 1 9 13 2
12 0 9 1 9 1 9 1 0 9 13 4 2
27 15 2 16 9 13 4 4 4 16 9 1 12 9 1 1 12 2 12 14 10 9 1 9 13 4 4 2
10 11 1 1 11 11 1 9 0 13 2
11 7 2 0 9 1 9 13 1 9 13 2
12 11 2 11 11 1 1 9 11 13 4 4 2
21 7 2 11 1 0 9 1 9 1 9 1 3 9 1 1 14 13 4 4 4 2
17 15 12 2 12 9 1 9 9 1 9 13 1 1 13 0 13 2
18 11 13 4 9 1 1 9 2 9 9 7 9 1 0 9 13 4 2
7 9 1 9 0 9 13 2
7 9 1 9 14 13 4 2
14 0 9 1 13 1 1 9 1 9 14 13 4 4 2
18 9 1 1 10 9 1 10 9 0 13 4 2 15 9 1 14 13 2
35 15 1 10 9 10 9 1 0 7 0 9 1 9 13 4 4 15 7 14 0 9 14 13 7 14 15 15 9 1 13 9 13 4 4 2
22 11 1 9 1 11 11 11 1 9 1 1 13 10 9 0 13 2 15 3 0 13 2
15 10 9 1 9 1 13 13 1 9 0 9 1 14 13 2
20 15 1 2 0 9 1 14 13 1 9 13 16 15 1 0 9 1 13 4 2
11 9 1 9 13 1 1 0 9 14 13 2
24 0 9 1 1 0 9 7 0 9 1 1 1 9 15 0 9 1 9 14 13 4 4 4 2
12 3 2 10 9 1 3 9 13 1 9 13 2
19 3 2 9 2 9 1 0 9 1 9 9 1 1 9 1 1 13 4 2
16 9 1 0 13 4 9 7 9 1 1 3 0 9 13 4 2
24 11 1 9 1 12 9 15 14 9 13 4 4 16 9 1 0 9 8 13 1 9 14 13 2
9 16 2 15 0 9 0 13 4 2
21 11 1 0 11 11 7 11 11 1 10 9 13 2 9 1 10 0 9 14 13 2
21 0 11 11 11 11 1 0 9 1 11 1 11 11 11 1 9 1 0 9 13 2
22 11 1 9 7 11 1 0 11 11 11 11 1 15 9 9 9 1 13 9 0 13 2
21 11 1 1 1 11 1 9 1 11 2 11 7 11 11 1 9 9 0 13 4 2
37 11 1 9 13 1 1 0 11 11 11 2 11 11 1 9 11 11 11 2 11 1 9 11 11 11 7 9 9 11 11 1 10 0 9 0 13 2
24 11 1 11 1 9 1 9 1 1 15 9 1 13 11 7 11 9 1 1 0 9 0 13 2
45 15 1 10 9 1 1 13 4 2 15 9 1 13 9 1 1 13 7 15 9 1 9 14 13 4 1 0 11 2 11 11 11 11 3 11 1 9 13 9 1 0 9 1 13 2
31 0 9 1 1 9 1 9 1 0 9 1 9 13 1 1 15 11 11 11 14 9 9 15 0 9 1 11 13 4 4 2
25 15 1 0 2 0 13 4 1 0 13 4 11 1 11 9 11 9 11 11 1 1 15 9 13 2
15 16 15 9 1 1 1 3 15 14 13 1 9 13 4 2
25 7 9 1 13 13 16 11 1 11 1 9 1 9 1 11 11 1 13 4 0 9 1 9 13 2
39 11 1 0 9 1 1 2 15 11 11 1 1 9 1 9 1 15 9 1 3 9 13 4 1 9 13 4 11 1 9 1 1 0 9 1 14 9 13 2
28 15 9 13 16 15 9 9 1 9 1 12 9 9 1 9 13 4 15 9 1 9 0 13 1 9 14 13 2
34 9 1 1 2 11 1 9 1 11 1 9 9 1 15 9 1 13 1 9 1 9 13 1 1 13 4 9 1 9 1 14 9 13 2
28 11 9 1 9 13 16 11 1 15 13 1 15 0 9 1 9 13 7 10 0 9 1 3 9 14 13 4 2
40 16 11 15 1 9 1 1 15 14 13 1 13 4 4 7 15 0 9 1 13 13 16 16 9 1 15 14 13 16 9 13 1 9 1 9 14 13 4 4 2
26 0 13 16 10 9 1 11 1 11 1 11 11 2 11 11 7 11 11 1 1 14 15 9 13 4 2
13 16 15 9 11 11 1 9 9 9 13 4 4 2
29 9 1 1 15 9 0 13 7 0 9 1 9 1 9 1 9 13 1 1 11 11 11 14 11 9 11 13 4 2
28 9 1 15 11 11 1 15 0 9 11 11 2 11 11 2 11 11 7 11 11 1 1 9 2 9 13 4 2
16 15 11 11 1 1 9 1 15 0 9 1 9 14 13 4 2
20 10 9 1 1 11 11 11 11 1 0 9 9 1 12 9 9 1 0 13 2
29 10 9 11 1 9 2 9 1 12 1 12 12 9 1 13 4 15 9 1 14 9 1 8 13 1 9 13 4 2
13 15 1 9 1 9 0 9 1 9 1 13 4 2
23 10 14 9 1 13 9 1 13 4 12 0 9 14 9 13 9 1 1 1 13 4 4 2
21 9 1 9 10 9 1 0 0 9 1 0 0 9 9 1 9 1 3 13 4 2
16 14 10 9 1 10 9 10 9 1 9 1 9 13 4 4 2
28 10 9 1 10 9 1 9 1 9 3 13 1 1 15 1 9 1 9 0 13 1 13 9 9 1 13 4 2
18 15 1 9 13 1 1 11 11 1 9 9 1 12 9 13 4 4 2
47 9 9 1 9 1 13 1 9 7 15 1 13 9 1 9 1 9 13 1 1 12 9 1 11 1 11 11 1 9 9 11 11 11 1 9 1 12 0 12 0 0 9 9 0 13 4 2
23 15 12 9 1 1 10 9 1 10 9 1 13 9 1 9 1 9 1 9 13 4 4 2
19 10 9 1 15 1 13 14 12 9 1 10 9 3 13 15 13 4 4 2
52 9 1 13 9 13 4 16 9 1 15 9 1 10 9 1 9 13 4 16 9 1 0 9 1 10 0 9 1 10 9 0 13 2 15 9 9 1 14 9 1 14 0 0 9 1 8 13 1 9 13 4 2
29 10 9 1 9 9 2 9 1 0 9 1 9 13 4 15 8 13 1 1 12 1 12 12 9 1 13 4 4 2
20 10 0 9 9 1 1 15 13 9 1 0 9 13 1 1 9 1 13 4 2
24 9 13 4 16 10 9 1 9 9 9 12 7 12 9 1 10 0 0 9 1 9 1 13 2
26 10 9 11 0 7 0 9 1 10 9 1 9 1 9 1 13 10 9 1 15 10 9 13 4 4 2
45 10 9 1 9 1 9 14 1 11 11 1 9 9 11 11 11 1 9 9 11 11 1 9 1 9 1 13 4 13 4 2 15 0 13 4 9 11 9 13 4 11 13 4 4 2
38 15 1 11 11 11 11 1 9 11 7 9 11 7 11 11 1 9 11 11 11 1 10 9 1 10 0 9 1 9 13 1 9 1 13 4 4 4 2
32 10 9 1 9 9 1 1 10 0 9 1 9 3 13 4 4 2 15 1 9 1 9 0 13 1 13 9 14 13 4 4 2
22 10 9 1 11 11 1 10 0 0 9 1 13 1 9 1 1 15 9 13 4 4 2
44 9 9 1 9 11 1 1 9 11 11 11 2 9 11 2 9 11 11 2 9 11 11 11 2 9 11 11 11 2 9 11 11 11 7 9 11 11 11 1 12 9 0 13 2
29 11 1 15 1 9 14 14 14 13 4 2 7 11 1 9 11 1 9 1 9 1 9 11 11 1 3 9 13 2
22 9 1 9 7 0 9 1 1 11 1 15 9 2 11 11 2 1 10 9 8 13 2
21 11 11 1 11 1 9 11 11 1 1 1 0 9 1 1 15 9 14 9 13 2
10 11 1 13 14 9 14 9 13 4 2
15 9 12 12 9 9 8 13 1 3 9 1 9 13 4 2
25 15 1 11 11 7 0 9 1 9 1 1 9 7 11 11 1 9 1 9 13 1 9 13 4 2
26 0 9 1 9 1 0 9 1 13 9 1 1 1 13 0 9 9 1 3 15 1 0 13 4 4 2
9 16 0 9 1 1 9 0 13 2
9 9 1 9 14 3 1 10 13 2
11 11 1 14 15 13 1 1 0 14 13 2
29 9 13 1 1 11 1 9 13 1 0 9 1 11 1 9 11 11 9 15 13 7 14 12 12 9 1 9 13 2
8 15 11 1 1 9 14 13 2
19 0 9 7 15 9 1 9 1 14 11 1 3 1 13 1 9 0 13 2
39 9 0 13 1 11 11 1 1 11 7 11 9 1 9 13 4 7 2 11 11 2 1 11 11 1 9 13 4 11 11 1 0 9 9 1 14 13 4 2
20 11 11 1 1 11 1 9 13 7 9 1 9 1 11 1 9 1 9 13 2
20 9 9 1 9 1 1 1 9 13 4 4 14 12 9 0 9 1 13 4 2
10 9 1 14 12 9 1 15 9 13 2
17 11 1 1 2 11 11 2 15 1 14 12 9 0 13 4 4 2
13 11 1 1 9 1 9 11 7 11 1 13 4 2
11 15 1 9 11 1 12 9 3 11 13 2
8 15 12 9 1 9 13 4 2
30 3 14 15 9 1 9 12 9 1 13 4 2 7 9 1 11 7 11 1 9 10 13 12 1 12 9 1 14 13 2
10 11 11 1 15 9 1 1 9 13 2
22 11 1 3 0 12 9 1 13 7 9 1 1 9 13 7 9 1 9 13 1 13 2
20 11 2 11 9 1 9 1 1 15 9 1 13 10 9 13 9 13 4 4 2
24 11 2 11 9 1 9 1 1 9 13 9 9 1 9 1 3 1 9 14 13 4 4 4 2
31 11 2 11 2 11 11 2 11 9 3 14 11 1 0 13 4 11 1 11 9 1 1 1 11 9 15 3 13 4 4 2
28 15 1 11 9 1 12 9 15 9 1 1 0 13 4 2 15 1 12 1 9 7 0 1 9 13 4 4 2
31 9 9 9 1 9 10 9 1 9 13 7 3 13 1 10 9 1 13 4 2 7 3 1 9 1 0 9 15 9 13 2
46 16 11 11 1 13 4 2 15 0 9 1 11 9 15 9 1 13 4 4 2 15 10 9 1 9 1 0 9 16 11 11 1 13 13 4 2 7 9 9 10 9 1 13 4 4 2
28 9 1 11 9 8 13 1 3 14 11 1 9 15 3 13 4 4 7 11 1 9 9 15 1 13 4 4 2
31 16 9 1 11 14 13 4 2 15 9 11 1 12 9 13 2 7 9 11 9 1 9 10 9 1 14 15 9 13 4 2
26 0 10 9 1 15 9 1 9 0 13 9 1 13 1 1 15 9 1 15 1 13 1 9 13 4 2
13 10 9 1 9 1 9 1 0 9 13 4 4 2
21 3 16 9 11 9 1 13 16 9 9 1 9 15 9 1 1 15 0 13 4 2
24 11 9 1 13 14 11 11 1 9 9 9 1 1 9 1 15 9 1 9 1 13 13 4 2
31 15 0 9 13 16 10 9 1 9 1 15 9 1 0 9 1 9 13 4 2 10 9 9 1 15 9 14 13 4 4 2
24 7 9 13 1 3 2 9 10 9 0 13 4 7 9 1 9 11 9 1 9 14 13 4 2
16 11 1 11 1 13 9 14 10 9 1 12 9 1 9 13 2
20 16 9 9 10 9 1 9 1 1 14 13 4 16 3 10 9 14 13 4 2
49 12 9 1 12 9 9 1 9 1 1 9 1 9 13 4 9 11 1 13 4 16 16 0 0 9 3 11 2 11 7 11 11 9 1 9 13 1 9 1 9 13 16 15 3 0 13 4 4 2
35 11 1 9 9 11 11 1 13 16 16 15 15 1 1 0 9 1 13 4 4 16 15 9 1 12 9 14 12 9 9 13 1 0 13 2
21 11 1 13 16 15 10 9 1 9 13 7 10 9 1 1 15 14 13 4 4 2
28 0 3 11 11 1 13 4 16 16 15 9 13 1 9 1 9 13 4 4 16 15 15 13 1 1 0 13 2
37 9 9 1 9 0 0 9 11 1 0 0 2 11 2 1 9 1 13 16 16 11 1 9 9 1 9 1 9 13 16 9 1 15 0 9 13 2
11 11 1 13 16 11 11 15 0 9 13 2
21 15 14 15 1 13 16 16 15 15 15 9 13 16 9 9 14 0 13 4 4 2
17 15 15 0 13 16 16 15 15 13 4 16 15 9 1 9 13 2
14 11 1 10 9 9 1 0 9 1 0 13 4 4 2
26 11 13 4 16 9 0 9 11 1 9 1 1 9 13 4 2 15 11 1 9 1 0 13 4 4 2
12 11 1 12 9 7 9 1 9 13 4 4 2
10 9 15 9 1 1 1 9 13 4 2
29 11 9 1 0 13 1 1 11 11 11 11 2 11 2 9 1 14 0 13 4 2 15 1 10 9 9 13 4 2
31 15 13 13 16 16 9 1 0 9 1 11 1 15 9 15 9 1 1 11 13 4 4 2 16 9 1 9 13 4 4 2
30 0 13 16 0 9 9 2 11 11 11 11 0 0 9 1 11 11 1 12 9 1 12 9 9 1 9 13 4 4 2
13 11 1 11 11 11 11 0 9 11 1 9 13 2
17 15 15 12 0 9 1 9 13 1 3 14 0 9 1 9 13 2
9 10 9 11 1 12 9 1 13 2
22 9 1 1 11 11 7 11 11 1 11 1 11 9 1 9 9 1 9 1 9 13 2
18 11 1 0 9 9 11 2 11 2 11 2 11 2 11 7 11 13 2
32 11 11 11 1 9 11 11 1 13 16 0 9 9 0 9 1 13 2 7 15 1 1 15 9 1 0 9 14 13 4 4 2
14 15 9 9 1 9 1 10 13 1 9 1 9 13 2
28 10 9 1 0 9 1 11 11 1 14 11 2 11 11 1 12 9 1 9 9 7 11 11 1 0 9 13 2
24 11 1 13 16 11 7 0 11 11 11 11 1 11 2 11 11 1 11 1 13 1 9 13 2
23 11 1 11 11 13 1 3 0 0 9 1 15 9 1 0 9 1 9 9 13 4 4 2
29 11 2 11 11 2 11 2 7 11 11 11 11 11 1 1 11 11 11 1 9 11 11 11 1 0 13 4 4 2
26 0 3 11 7 11 9 14 11 1 9 13 4 4 16 11 11 0 9 1 11 1 9 14 13 4 2
23 11 1 9 9 11 11 1 13 13 1 10 9 0 13 16 15 14 15 9 1 0 13 2
13 7 11 11 9 1 15 13 15 9 14 13 4 2
12 7 15 13 10 0 13 16 11 11 13 4 2
20 11 11 1 9 13 15 11 1 9 13 4 4 16 15 11 1 9 1 13 2
15 0 15 10 9 1 9 13 7 12 9 13 11 13 4 2
19 15 9 13 16 9 1 9 0 13 1 3 14 11 11 0 11 13 4 2
26 15 9 13 16 11 1 9 9 13 1 3 9 9 1 9 9 1 13 16 11 11 0 11 13 4 2
31 7 11 11 1 13 13 16 0 9 1 0 13 14 0 9 9 1 0 13 4 4 7 0 9 9 1 1 13 4 4 2
16 15 1 11 11 1 0 11 13 4 0 9 1 0 14 13 2
12 11 15 10 9 1 14 13 4 1 0 13 2
27 11 1 3 14 13 1 1 13 13 16 11 11 1 15 9 1 9 0 13 1 1 15 9 13 4 4 2
21 11 11 7 11 9 14 10 9 1 0 13 16 11 1 9 1 11 1 9 13 2
9 11 11 1 9 1 13 4 4 2
20 12 11 11 1 9 13 4 7 0 11 11 1 11 15 9 13 1 9 13 2
27 10 9 13 16 11 11 11 11 1 1 15 13 4 4 16 15 0 9 1 9 13 7 0 9 1 13 2
17 11 7 11 9 1 13 13 16 11 11 1 10 13 13 0 13 2
19 11 11 1 15 15 12 9 1 9 1 1 1 11 1 15 9 13 4 2
32 11 1 12 9 1 11 1 11 11 1 9 1 9 13 4 13 16 12 9 1 9 9 1 12 9 9 1 9 0 13 4 2
19 11 11 1 15 1 15 9 13 15 0 0 9 1 9 1 0 13 4 2
13 7 9 14 1 15 9 9 1 9 1 13 4 2
19 15 2 11 11 1 0 9 15 9 1 9 13 15 11 9 14 13 4 2
14 11 2 11 11 11 1 15 11 1 9 13 4 4 2
17 15 9 1 13 13 16 11 11 1 11 0 9 1 9 13 4 2
10 15 11 9 7 15 9 1 9 13 2
18 11 1 13 13 16 10 9 1 15 9 13 14 16 15 0 14 13 2
10 11 3 1 9 1 9 13 4 4 2
18 15 9 1 13 13 16 15 1 11 0 9 1 11 1 13 0 13 2
21 15 1 3 3 14 11 9 11 1 0 9 1 9 9 13 1 9 13 4 4 2
34 11 1 9 11 1 11 11 0 11 11 11 1 9 1 12 9 1 11 1 12 9 2 12 9 7 0 9 1 9 9 0 13 4 2
27 9 9 1 1 11 11 1 11 11 11 1 9 9 0 13 4 4 7 15 11 1 1 1 14 13 4 2
10 3 9 10 9 1 9 13 4 4 2
31 9 1 13 16 9 1 9 1 1 9 13 4 15 15 9 1 13 12 9 13 15 9 1 1 11 11 13 4 4 4 2
10 9 1 13 9 1 11 1 9 13 2
17 9 1 0 0 9 1 15 9 13 15 13 16 15 0 14 13 2
48 11 11 11 1 9 1 13 13 16 16 10 9 1 11 1 1 1 14 13 4 4 7 9 1 11 1 9 0 13 15 9 13 16 10 9 10 9 13 4 4 15 11 1 9 9 1 13 2
31 11 1 9 9 11 11 11 1 13 2 16 10 9 1 9 13 1 9 1 9 1 1 1 15 9 1 9 13 9 13 2
16 7 15 0 13 16 11 1 14 9 9 13 9 13 4 4 2
22 0 0 9 1 0 13 9 1 9 1 1 0 9 9 1 1 12 12 9 13 4 2
30 11 1 9 1 0 9 1 13 4 11 9 9 1 9 1 9 1 9 9 1 14 12 12 9 13 1 9 13 4 2
18 10 9 1 11 9 9 1 0 9 1 12 2 12 12 9 13 4 2
21 11 11 11 1 1 10 9 1 0 9 1 13 1 1 9 0 13 4 4 4 2
25 11 9 1 11 11 11 2 11 2 1 1 10 9 9 1 9 13 4 2 11 11 15 9 13 2
17 11 1 9 1 9 1 11 9 9 1 12 9 0 13 4 4 2
17 10 9 1 9 1 11 11 11 1 0 9 1 11 13 4 4 2
27 11 1 9 1 13 4 4 0 9 13 4 1 0 13 1 11 11 1 11 1 9 9 1 0 9 13 2
23 9 1 9 13 16 9 9 1 1 12 9 1 1 11 11 11 11 11 1 9 9 13 2
5 15 9 14 13 2
25 11 11 1 9 1 1 12 9 9 0 13 4 2 15 1 12 9 0 9 11 11 1 14 13 2
18 15 1 15 10 9 10 9 1 13 4 15 11 11 1 13 13 4 2
30 0 9 1 13 16 9 1 9 1 9 14 1 14 11 11 11 2 11 2 1 11 0 3 0 11 11 1 9 13 2
21 11 1 13 4 9 1 1 11 11 1 9 1 12 9 7 10 9 0 13 4 2
34 11 9 11 11 11 1 11 11 1 0 9 1 1 10 9 1 9 13 4 15 11 1 11 11 11 1 9 11 11 1 13 13 4 2
36 0 9 9 11 11 7 9 11 11 11 1 12 0 9 1 11 0 11 11 1 0 9 9 9 1 9 1 11 1 9 13 1 9 13 4 2
41 11 11 11 1 0 12 9 9 1 9 13 4 9 1 9 1 9 9 2 9 9 2 9 9 7 11 9 1 9 1 9 1 3 9 9 13 1 9 13 4 2
27 15 1 14 9 1 9 1 10 9 1 9 13 4 1 1 10 9 3 14 0 13 1 9 14 13 4 2
37 9 1 9 1 0 9 1 13 4 9 1 1 1 9 1 1 1 13 4 9 1 9 0 13 4 13 16 9 1 9 9 1 15 9 14 13 2
10 9 1 0 9 0 9 13 4 4 2
37 15 1 14 9 1 11 2 11 2 11 2 11 2 7 11 9 1 9 1 1 11 0 13 1 1 9 9 1 11 11 1 9 13 1 13 4 2
19 12 9 7 12 9 13 1 1 11 11 1 11 1 9 13 14 4 4 2
20 11 11 11 1 11 1 12 7 11 1 12 9 1 0 13 1 9 13 4 2
17 15 1 14 9 1 10 9 11 9 1 9 13 12 13 4 4 2
46 11 7 11 1 9 1 9 13 4 16 16 10 9 13 1 9 1 9 3 9 13 1 13 16 11 2 11 1 9 9 13 4 4 2 16 9 1 3 10 9 9 1 1 13 4 2
14 11 11 1 0 9 12 9 11 1 9 1 13 4 2
15 16 10 9 12 0 9 13 4 15 11 11 0 14 13 2
13 16 0 9 1 13 1 9 15 10 13 4 4 2
12 0 9 14 0 9 9 1 1 3 13 4 2
16 15 11 11 1 13 1 9 1 9 0 9 0 13 4 4 2
39 11 9 1 9 7 11 9 9 11 11 1 1 11 1 11 9 1 13 0 9 1 9 13 2 16 0 12 2 12 9 1 9 9 9 0 13 4 4 2
17 15 1 1 9 1 0 9 0 11 11 1 0 9 1 13 4 2
23 10 9 1 9 1 11 2 11 2 11 7 11 1 11 1 12 2 12 9 13 4 4 2
10 11 1 0 9 12 9 0 13 4 2
20 9 11 1 1 15 1 9 14 1 11 1 10 12 0 9 9 1 13 4 2
13 11 1 11 9 1 11 1 12 9 3 13 4 2
14 10 0 9 11 2 11 11 1 9 1 13 4 4 2
11 15 10 9 1 11 11 11 11 13 4 2
18 10 9 11 2 11 11 1 9 13 1 1 0 9 1 13 4 4 2
33 3 10 9 13 4 4 4 2 15 12 9 1 11 2 11 2 11 2 11 7 11 2 11 9 1 13 1 0 13 4 4 4 2
20 7 15 15 9 0 13 4 4 16 11 2 11 11 1 0 9 0 14 13 2
17 0 13 16 11 1 9 1 11 0 13 4 1 9 13 4 4 2
23 9 11 1 1 10 12 0 9 1 0 9 1 9 1 13 9 13 0 9 1 9 13 2
11 15 1 9 9 1 9 14 13 4 4 2
15 10 9 10 0 9 1 14 11 1 9 9 13 4 4 2
12 15 15 12 10 9 1 14 9 13 4 4 2
15 11 1 11 11 11 11 1 10 0 9 1 9 13 4 2
22 11 1 13 16 11 1 0 9 13 9 9 1 9 13 1 9 3 9 13 4 4 2
15 11 1 11 1 0 9 9 11 11 1 14 10 9 13 2
20 11 11 1 1 0 9 1 9 1 1 15 9 0 9 14 13 4 4 4 2
14 15 12 9 1 10 9 13 4 1 9 13 4 4 2
20 10 9 1 13 1 9 13 4 4 2 10 9 1 9 7 9 9 0 13 2
20 9 9 1 13 16 9 1 9 0 9 1 12 9 13 4 1 9 10 13 2
15 9 1 1 9 1 0 9 1 1 9 13 4 4 4 2
14 9 1 0 12 9 1 9 15 14 0 13 4 4 2
28 11 1 0 9 1 1 9 7 10 0 9 1 9 3 9 13 4 4 7 9 1 9 1 9 13 4 4 2
25 9 2 9 9 1 12 0 9 9 1 0 9 1 9 1 1 3 2 3 14 0 13 4 4 2
11 11 11 11 1 0 3 9 1 9 13 2
16 9 1 13 9 1 0 9 1 0 9 13 7 15 14 13 2
17 15 10 14 9 1 11 11 7 11 11 1 14 10 9 13 4 2
31 11 11 1 13 4 16 9 13 9 0 9 7 0 9 1 9 13 2 10 9 1 15 0 9 1 15 14 13 4 4 2
16 9 9 1 13 16 9 1 9 9 11 11 9 1 14 13 2
14 9 1 14 12 12 9 1 0 9 1 9 13 4 2
13 15 9 1 13 4 10 9 1 13 4 4 4 2
11 0 9 1 15 9 1 13 4 4 4 2
35 9 1 9 1 13 13 4 9 1 11 1 13 16 11 11 1 10 0 9 10 0 13 16 15 9 1 9 1 1 14 8 14 13 4 2
28 11 11 11 7 0 11 11 11 1 1 11 1 11 1 11 11 11 11 1 13 9 3 9 1 14 0 13 2
22 16 2 12 9 1 9 2 11 11 7 11 11 1 0 9 1 9 1 14 9 13 2
10 12 9 0 2 0 9 1 11 13 2
12 9 1 1 11 1 15 10 14 0 9 13 2
15 11 1 13 16 10 9 0 9 1 1 12 0 9 13 2
24 3 1 11 1 15 11 9 1 9 1 11 1 1 11 11 1 12 0 9 9 1 0 13 2
25 12 9 1 9 1 0 9 1 0 9 9 13 4 13 16 15 15 14 9 1 15 9 14 13 2
27 11 1 13 16 2 9 1 15 9 14 13 2 9 1 15 9 14 13 7 15 15 14 9 1 9 14 13
15 9 1 10 9 9 13 15 0 9 1 13 1 13 4 2
12 15 13 16 15 9 1 9 1 0 13 4 2
9 10 9 11 1 0 13 4 4 2
13 10 0 9 1 15 14 9 1 9 14 13 4 2
11 11 1 13 16 10 9 9 1 1 13 2
19 9 1 11 2 11 7 11 1 13 9 1 13 4 0 9 9 14 13 2
28 11 1 9 1 9 0 13 4 11 1 13 16 9 1 13 1 1 10 3 1 9 7 0 9 1 9 13 2
27 9 1 1 12 9 1 11 11 11 11 1 11 1 0 9 2 9 9 7 0 9 9 1 14 9 13 2
23 11 1 13 16 12 9 1 0 9 7 9 1 9 13 1 1 12 0 0 9 13 4 2
20 11 11 1 11 11 1 9 9 1 9 1 14 9 13 1 0 13 4 4 2
16 15 1 12 9 9 9 0 13 1 1 0 9 1 9 13 2
28 11 1 13 16 11 7 11 9 9 2 9 1 0 9 1 9 7 0 9 9 1 9 1 14 13 9 13 2
15 12 9 1 9 9 1 0 12 9 1 14 9 13 4 2
21 11 1 11 1 1 0 7 0 9 2 9 1 1 12 12 9 1 9 13 4 2
15 11 2 11 11 11 1 9 13 4 11 1 10 9 13 2
26 11 11 11 1 11 1 11 1 0 11 11 11 1 9 1 0 9 1 13 9 2 9 1 9 13 2
12 11 1 11 1 9 9 7 11 1 9 13 2
23 3 10 0 9 13 15 0 11 1 11 1 0 11 1 9 1 10 9 1 9 13 4 2
32 11 1 9 2 9 1 13 16 11 11 1 9 1 9 1 9 9 1 9 1 13 4 4 2 15 9 1 15 0 9 13 2
13 11 1 13 16 15 11 1 9 1 9 13 4 2
16 15 12 0 0 9 1 9 1 9 0 13 1 10 9 13 2
16 11 1 11 1 9 7 11 1 9 1 1 15 9 0 13 2
22 11 1 11 1 11 11 2 11 11 2 11 11 1 10 0 9 13 1 9 13 4 2
15 15 11 11 11 11 2 11 11 7 11 11 14 0 13 2
29 10 0 9 9 1 9 11 1 1 0 9 13 1 0 11 11 11 11 1 9 1 9 13 1 1 13 4 4 2
31 0 9 1 12 0 9 1 13 16 11 9 1 3 13 4 0 2 0 9 1 0 9 3 14 13 1 9 13 4 4 2
16 13 1 10 9 1 12 9 1 1 10 3 13 1 9 13 2
23 11 11 11 11 11 11 13 4 4 7 0 11 11 9 11 11 11 14 11 13 4 4 2
31 9 1 13 16 12 0 0 0 9 9 1 9 14 1 0 9 9 1 1 11 11 2 11 11 11 11 1 9 13 4 2
14 15 1 11 1 11 11 11 1 0 9 13 4 4 2
27 15 13 16 11 1 12 0 0 9 1 9 1 9 1 13 0 9 1 11 11 7 9 1 1 9 13 2
20 15 9 13 16 15 0 9 7 9 2 9 9 1 9 1 9 0 13 4 2
18 16 15 12 14 9 1 9 0 9 1 0 13 1 1 10 0 13 2
41 9 1 13 16 0 0 9 1 12 9 1 9 1 1 0 9 1 0 9 13 1 9 13 4 11 1 11 1 9 9 1 12 0 9 9 13 1 9 13 4 2
45 11 11 1 9 1 0 9 1 9 2 9 7 0 0 9 1 9 1 14 0 13 1 9 0 13 1 9 1 0 9 1 13 16 11 11 1 11 11 1 11 1 9 13 4 2
28 0 9 1 11 11 1 9 1 9 9 1 9 1 10 12 9 1 9 13 1 11 11 1 8 13 4 4 2
42 9 1 13 4 9 1 13 4 4 16 10 9 7 9 9 1 0 9 2 9 9 1 0 9 2 9 9 7 0 9 1 1 0 9 1 1 9 9 13 4 4 2
28 9 1 9 11 11 1 13 16 11 15 3 11 11 1 0 9 14 13 15 1 15 0 9 13 1 9 13 2
16 16 11 1 9 1 1 9 1 0 9 1 10 9 13 4 2
17 11 11 11 11 11 2 11 2 1 0 9 1 9 13 4 4 2
23 9 1 9 9 7 11 11 11 2 11 2 1 11 0 13 1 14 9 13 4 4 4 2
28 11 11 11 1 9 11 11 1 13 4 16 9 9 1 0 9 1 1 9 11 1 9 1 9 1 0 13 2
37 0 9 9 11 1 11 1 0 9 1 0 13 4 11 1 13 16 11 1 0 9 1 1 0 9 1 9 1 15 9 1 15 9 13 4 4 2
20 9 1 9 9 7 11 1 11 0 13 7 9 1 1 15 12 0 9 13 2
21 16 15 11 1 9 14 1 0 13 4 9 1 15 13 1 15 9 9 14 13 2
39 15 13 16 11 1 0 9 1 0 13 4 4 16 9 1 13 1 14 9 1 9 13 4 4 7 15 15 14 9 1 11 1 1 15 9 14 13 4 2
36 11 1 13 16 11 1 1 14 10 9 1 9 13 4 4 15 9 15 9 1 9 1 0 9 7 9 1 13 9 1 9 1 9 13 4 2
38 15 13 16 11 0 13 1 3 9 1 9 1 10 10 9 1 9 1 9 13 2 15 1 9 13 1 13 1 1 9 9 1 9 1 13 4 4 2
24 15 13 16 10 9 1 9 1 9 1 9 1 13 1 1 11 11 1 11 1 0 13 4 2
17 15 13 16 15 9 15 14 13 16 11 1 3 9 14 13 4 2
10 9 10 9 1 9 1 1 0 13 2
11 9 1 0 13 4 1 15 3 13 4 2
45 15 13 4 1 16 15 9 1 0 0 9 15 15 15 9 1 13 1 1 13 4 2 11 1 9 1 3 13 4 4 2 15 13 16 11 1 1 14 0 9 1 13 4 4 2
23 9 11 2 11 1 1 11 11 11 2 11 2 8 13 1 0 9 11 11 2 11 13 2
11 10 9 0 9 1 1 0 13 4 4 2
13 11 11 1 10 9 1 0 9 0 13 4 4 2
14 10 9 1 9 11 11 7 11 1 9 1 0 13 2
25 11 11 11 1 1 9 1 15 9 9 1 1 0 9 1 1 13 4 0 9 1 9 13 4 2
113 9 1 9 9 1 9 12 12 7 15 9 1 9 1 9 2 9 9 9 1 12 12 9 7 15 9 1 9 1 9 2 12 12 9 7 15 9 1 9 9 9 1 9 1 9 2 15 9 1 9 7 9 1 9 1 12 12 9 7 15 9 1 9 1 9 2 15 9 1 11 1 12 12 9 7 15 9 1 9 2 12 12 9 7 15 9 1 0 9 1 9 2 9 7 12 12 7 15 9 1 11 9 9 1 9 1 9 11 1 1 13 4 2
23 0 13 16 11 11 11 1 1 11 11 11 1 12 0 9 11 11 1 9 13 4 4 2
20 10 9 1 1 0 9 0 9 1 0 9 1 0 9 1 9 9 1 13 2
21 10 9 0 9 1 11 11 1 9 1 1 11 7 11 11 11 1 1 13 4 2
14 11 11 11 10 9 1 9 13 11 11 1 13 4 2
18 15 9 1 9 1 9 1 0 13 14 0 9 1 1 0 14 13 2
35 11 7 11 1 1 11 11 11 11 2 11 2 1 14 10 9 1 9 2 9 1 0 9 9 1 10 9 9 13 1 9 13 4 4 2
8 10 9 11 11 1 0 13 2
36 11 1 9 7 0 9 11 11 11 1 11 1 13 16 9 1 15 9 9 1 9 1 1 9 9 1 9 9 1 12 9 1 9 13 4 2
22 15 13 16 15 13 0 13 4 4 16 9 1 9 1 0 9 12 9 13 4 4 2
20 10 9 1 9 1 10 9 1 9 9 1 0 9 9 12 9 13 4 4 2
31 0 3 11 11 1 9 9 9 11 11 1 13 16 9 9 1 0 9 0 9 9 1 9 1 15 14 13 4 4 4 2
21 15 13 16 9 9 1 9 9 1 14 12 1 12 9 1 9 13 4 4 4 2
20 16 2 13 4 4 16 9 9 7 9 9 1 0 9 1 9 14 13 4 2
22 15 13 16 0 9 1 9 1 9 9 1 13 1 1 9 1 1 15 9 14 13 2
35 0 13 16 11 11 1 9 9 1 0 9 1 9 1 11 7 11 11 9 13 4 1 3 11 11 1 9 9 1 9 9 13 4 4 2
12 9 9 1 9 9 13 1 11 3 14 13 2
21 11 11 11 10 9 13 15 1 9 1 11 1 1 0 0 9 1 9 13 4 2
37 0 9 1 9 2 11 2 1 9 9 1 9 1 1 1 9 15 2 9 2 9 2 9 2 0 13 1 12 9 1 1 1 9 13 4 4 2
26 9 9 9 1 9 11 11 1 13 16 11 9 1 1 10 9 9 1 15 9 1 12 9 13 4 2
22 16 2 0 9 1 9 1 9 7 0 9 1 14 10 9 1 14 9 9 13 4 2
24 15 9 1 1 1 10 9 2 9 2 9 2 9 2 1 9 1 1 0 9 1 9 13 2
11 15 15 11 9 12 9 1 13 4 4 2
16 9 1 9 9 1 9 1 1 9 1 0 9 14 13 4 2
55 9 11 11 1 13 2 2 15 15 1 15 13 1 13 14 4 4 4 16 9 9 1 0 13 4 9 0 9 9 0 13 4 4 16 9 12 10 9 1 0 0 13 4 2 15 15 9 7 0 9 1 9 13 4 4
31 11 11 1 0 9 7 11 11 11 1 9 11 1 11 11 1 13 9 1 9 1 11 11 1 9 1 0 13 4 4 2
18 3 1 11 1 9 9 1 15 11 11 1 0 9 1 13 4 4 2
32 11 1 9 1 1 9 1 13 16 11 11 11 1 11 11 2 11 2 2 11 2 1 1 1 9 1 9 14 13 4 4 2
31 15 13 16 9 1 11 11 1 1 9 13 1 9 13 2 7 15 11 2 11 2 2 11 2 1 14 9 14 13 4 2
21 0 13 16 9 1 10 9 1 9 1 0 9 9 11 11 1 0 13 4 4 2
39 9 1 9 1 1 1 0 0 9 11 11 1 10 9 1 0 13 4 16 9 9 7 9 9 1 11 11 11 1 11 11 1 1 9 13 1 14 13 2
18 9 1 1 11 1 11 1 0 9 11 11 1 9 1 9 14 13 2
23 11 1 13 16 11 11 1 9 1 11 11 1 9 1 10 9 1 0 14 13 4 4 2
22 7 2 9 1 9 9 1 1 1 0 0 9 11 11 11 11 1 9 1 13 4 2
18 11 1 13 16 11 11 1 9 1 11 11 1 9 1 9 13 4 2
26 9 1 13 16 0 9 1 15 15 0 14 13 4 16 9 1 9 1 0 9 0 9 7 9 13 2
28 9 1 9 1 9 1 9 13 4 13 16 9 9 1 1 9 15 14 9 1 11 1 9 1 13 13 4 2
34 9 1 13 16 9 9 1 0 9 1 11 1 9 1 13 9 14 0 13 15 9 13 4 16 9 15 15 14 9 0 13 13 4 2
19 9 1 1 11 1 13 16 9 9 1 1 9 1 1 0 0 9 13 2
12 15 9 2 9 11 1 0 9 14 0 13 2
29 9 9 1 1 12 9 1 0 9 14 13 15 15 9 13 4 16 9 1 9 1 1 15 9 1 13 4 4 2
29 12 9 1 13 4 16 9 1 10 9 1 11 1 13 4 16 16 15 15 13 4 16 15 1 9 14 0 13 2
13 11 1 13 16 11 1 10 9 0 9 1 13 2
6 15 9 13 4 4 2
31 9 1 10 9 1 14 9 13 16 9 9 1 10 9 9 1 14 9 13 4 15 1 9 7 9 1 1 9 13 4 2
20 15 1 12 10 9 1 9 14 13 2 15 9 1 10 9 1 13 4 4 2
32 9 1 15 1 14 9 13 16 10 14 10 12 9 1 9 1 9 13 4 7 15 9 13 1 1 9 1 9 13 4 4 2
29 9 1 1 9 1 12 9 15 1 13 2 16 9 9 1 9 13 14 14 4 16 9 9 1 1 9 13 4 2
30 9 11 1 13 16 11 11 1 0 9 1 9 1 13 10 9 1 13 7 14 13 1 15 9 0 14 13 4 4 2
36 11 9 11 1 0 9 1 9 7 9 1 9 1 13 9 14 1 13 0 9 1 1 15 11 1 0 9 0 9 13 1 9 13 4 4 2
11 9 1 15 11 7 0 9 1 9 13 2
37 10 9 1 11 13 0 11 11 11 11 1 13 16 15 9 13 16 10 9 9 1 9 1 1 0 9 7 9 1 9 1 15 9 1 9 13 2
18 0 9 1 13 4 10 9 1 1 12 9 1 9 1 13 4 4 2
19 11 1 0 9 1 12 9 7 12 0 9 1 12 9 1 0 13 4 2
15 9 9 1 9 7 9 13 9 1 1 9 13 4 4 2
36 11 1 11 11 11 11 11 11 1 11 1 10 9 1 9 13 4 13 16 9 9 1 1 0 9 1 11 1 13 4 9 15 0 9 13 2
36 0 3 0 11 11 11 11 1 11 1 11 11 11 11 11 1 9 1 1 13 2 2 15 9 13 16 15 9 1 12 9 1 9 13 4 2
7 15 9 1 9 13 2 2
21 9 1 11 11 1 9 1 9 1 1 15 15 14 11 9 1 0 11 9 13 2
26 15 15 13 4 16 15 15 11 1 0 9 0 13 4 1 9 13 4 2 15 15 10 9 13 4 2
24 12 9 1 9 1 11 13 0 11 11 1 9 13 16 9 1 0 9 1 0 9 0 13 2
22 15 1 11 11 1 11 1 13 16 9 11 1 9 1 11 1 9 10 13 4 4 2
17 11 11 1 11 1 0 9 9 1 13 4 9 1 9 14 13 2
19 0 13 16 11 9 1 9 1 1 9 9 9 1 9 13 4 4 4 2
38 9 1 12 0 9 9 1 9 0 13 1 9 13 4 4 2 7 11 1 9 1 11 11 11 11 2 11 2 1 9 9 15 14 0 9 0 13 2
9 10 9 0 9 9 9 1 13 2
24 11 1 3 0 9 1 1 12 11 11 11 1 11 1 0 9 12 9 1 9 13 0 13 2
32 2 11 2 2 2 11 11 11 2 7 0 9 2 11 11 11 2 1 9 12 0 11 1 11 1 9 9 1 13 4 4 2
8 16 3 1 15 13 4 4 2
25 15 1 9 1 9 13 1 11 9 12 0 9 1 1 9 7 9 1 1 3 2 3 13 4 2
11 12 9 1 11 1 0 0 9 1 13 2
43 12 9 1 9 1 10 3 0 9 1 12 9 1 9 1 9 1 9 1 9 13 13 1 1 9 14 1 9 9 7 9 1 10 9 0 13 16 9 1 9 13 4 2
13 15 0 9 13 2 15 0 9 1 15 9 13 2
8 0 9 1 9 1 9 13 2
28 11 2 11 7 11 1 1 10 9 3 11 11 2 11 1 13 7 15 1 0 9 1 14 3 10 9 13 2
12 16 11 1 9 13 9 1 9 0 13 4 2
29 11 2 11 2 11 7 11 1 14 9 1 9 1 1 11 1 9 1 0 9 1 9 9 1 15 14 13 4 2
27 9 1 14 12 9 1 11 1 9 1 9 1 9 13 7 3 3 2 3 15 9 1 13 4 13 13 2
32 11 1 1 0 0 9 2 11 2 11 2 11 7 11 1 0 9 1 9 1 15 2 15 9 1 10 0 9 1 9 13 2
17 11 1 10 9 1 13 1 1 11 1 9 1 12 9 13 4 2
15 7 9 13 9 1 15 7 9 1 9 1 9 13 4 2
9 15 1 9 1 9 10 14 13 2
12 9 1 9 0 13 15 15 9 13 0 13 2
36 0 9 1 9 7 11 11 11 1 8 11 11 1 13 16 0 9 1 1 15 9 13 4 7 0 9 1 13 1 10 9 1 9 13 4 2
35 10 9 1 0 9 11 11 11 1 13 16 9 14 1 9 1 13 4 9 1 9 1 9 1 11 1 0 9 1 9 13 1 9 13 2
20 10 9 1 10 9 1 14 8 13 4 2 15 0 9 1 13 4 4 4 2
20 15 13 16 10 9 1 9 9 7 11 1 1 9 13 1 1 14 13 4 2
18 9 1 1 11 2 11 2 11 7 11 1 9 0 9 1 13 4 2
11 9 7 9 14 15 13 1 3 14 13 2
25 16 9 1 0 9 1 10 9 1 14 13 1 9 13 4 2 7 10 9 1 15 3 14 13 2
37 0 9 1 10 9 9 9 1 14 1 13 7 16 11 3 0 13 15 15 9 1 9 1 13 14 4 7 15 9 1 9 1 1 9 13 4 2
14 0 13 16 15 1 12 9 10 9 8 13 4 4 2
10 10 9 12 9 1 12 9 13 4 2
21 12 9 1 11 1 11 1 9 13 4 2 7 12 9 1 11 1 9 13 4 2
32 11 11 11 2 11 2 1 9 9 1 9 1 10 12 9 1 1 13 9 1 11 1 11 11 11 11 1 0 13 4 4 2
32 3 9 1 15 1 1 9 13 4 4 2 7 13 4 4 16 9 9 9 14 13 10 9 1 9 13 1 9 13 4 4 2
23 10 9 1 0 9 1 9 1 9 1 9 7 10 9 1 9 1 9 13 4 4 4 2
34 13 4 4 4 16 10 9 13 1 3 15 9 1 9 14 0 13 2 10 9 1 9 1 10 9 1 9 0 13 1 9 13 4 2
13 9 1 9 1 14 10 9 1 9 13 4 4 2
29 7 10 9 1 9 13 4 4 16 9 9 1 9 0 13 1 9 1 9 9 9 14 13 1 0 13 4 4 2
13 0 9 1 1 9 9 1 9 13 4 4 4 2
23 10 9 14 13 4 4 16 9 9 1 12 0 9 13 1 11 11 1 9 0 14 13 2
31 0 13 16 11 11 1 11 9 1 1 9 1 1 11 11 1 15 9 13 4 16 10 12 9 1 12 0 9 13 4 2
22 10 12 9 9 1 9 1 11 9 11 11 11 11 1 9 11 11 11 1 9 13 2
24 14 12 9 13 9 1 9 1 9 1 11 11 1 11 1 13 9 1 13 9 1 0 13 2
22 9 1 1 13 1 3 10 9 1 9 1 1 13 9 1 9 13 1 3 9 13 2
13 15 14 15 13 13 16 15 10 9 1 0 13 2
18 15 15 15 9 9 1 9 1 9 1 13 4 1 9 1 0 13 2
17 15 1 11 11 1 10 9 1 0 9 1 15 9 13 4 4 2
61 9 1 9 1 1 9 1 9 1 11 2 11 1 9 11 11 2 11 2 11 1 9 11 11 2 11 2 11 1 9 11 11 2 11 2 11 1 9 11 11 2 11 2 11 1 9 11 11 11 7 11 2 11 1 9 11 11 11 0 13 2
23 0 9 1 9 1 11 1 9 1 9 1 11 1 9 1 12 9 1 9 1 9 13 2
7 9 1 14 10 9 13 2
9 9 1 1 9 9 14 13 4 2
25 3 9 1 9 9 1 1 9 14 1 1 9 0 13 4 4 3 9 1 12 9 15 13 4 2
25 10 9 1 13 1 1 11 11 11 1 9 1 9 11 11 1 14 9 13 7 15 9 14 13 2
10 9 0 9 1 9 1 13 4 4 2
41 11 11 11 11 11 1 13 13 11 9 11 11 11 1 0 9 1 13 16 10 9 1 9 15 1 0 9 1 14 13 15 1 0 9 9 1 13 14 4 4 2
9 15 11 11 7 11 11 0 13 2
10 15 1 11 9 14 9 1 13 4 2
16 11 9 9 13 4 4 2 9 9 2 9 9 2 9 13 2
16 11 1 1 1 9 1 9 11 11 7 11 11 13 4 4 2
22 9 1 1 9 11 11 1 11 9 1 13 16 15 11 11 1 13 1 9 13 4 2
22 7 9 9 0 13 7 9 1 9 0 14 13 7 11 1 9 1 9 9 13 4 2
17 11 1 1 1 11 11 11 1 13 9 13 4 7 9 0 13 2
16 10 3 11 1 9 11 11 13 2 13 4 9 13 4 4 2
33 11 9 1 10 9 1 9 1 1 9 1 9 0 14 13 15 11 11 3 13 7 9 1 9 1 1 13 15 9 1 9 13 2
8 15 1 9 9 1 0 13 2
16 15 1 9 3 13 7 9 9 1 1 3 0 13 4 4 2
14 9 2 9 1 1 9 3 9 1 9 14 13 4 2
34 9 1 2 11 11 11 1 13 9 9 1 9 13 1 2 9 1 1 9 11 11 11 1 9 1 9 9 14 1 1 0 13 4 2
21 9 9 9 1 9 15 9 13 15 9 1 0 9 1 9 9 13 1 1 13 2
39 11 1 1 1 15 11 11 1 9 9 13 1 9 13 15 9 1 9 13 9 13 4 16 9 1 9 15 1 9 13 4 15 1 9 0 13 4 4 2
28 15 9 13 16 9 9 9 11 11 1 13 1 9 14 13 4 2 15 15 10 9 11 1 1 13 13 4 2
27 15 15 9 1 11 1 13 3 9 9 1 9 13 4 7 15 1 14 9 1 9 3 13 4 4 4 2
38 11 11 1 13 16 15 15 9 1 13 15 9 9 11 11 1 9 9 1 13 4 4 2 7 9 0 9 9 1 13 1 9 14 14 13 4 4 2
22 11 11 3 15 9 13 4 16 9 1 11 1 13 4 7 15 9 9 1 9 13 2
9 0 9 1 14 9 9 13 4 2
8 11 11 3 9 13 4 4 2
26 0 9 1 15 9 1 9 1 9 13 15 11 1 13 16 15 9 13 16 9 1 9 15 13 4 2
17 15 13 13 16 16 15 9 14 13 16 9 1 9 3 14 13 2
13 11 1 11 11 11 11 11 1 9 11 11 13 2
18 11 11 11 1 3 11 0 13 1 3 15 11 1 0 9 9 13 2
28 11 1 15 11 11 11 11 1 9 1 1 11 1 1 1 11 1 9 1 9 1 9 13 4 1 9 13 2
12 15 1 15 11 11 11 11 11 1 14 13 2
11 15 11 11 11 1 14 13 1 9 13 2
24 0 9 1 9 1 11 0 10 9 13 15 9 1 0 9 1 13 9 9 0 13 4 4 2
15 0 0 11 11 14 9 1 9 1 9 13 9 13 4 2
13 9 1 15 9 1 9 7 3 1 0 9 13 2
16 9 1 9 1 15 9 2 9 2 9 7 9 1 9 13 2
31 11 11 1 9 1 9 2 9 2 9 1 9 2 15 1 1 9 7 9 1 9 1 9 10 0 9 1 0 13 4 2
20 15 1 9 1 9 1 15 9 1 9 2 9 7 13 4 0 9 13 4 2
11 9 1 9 1 9 9 13 7 0 13 2
14 9 1 9 1 15 9 1 0 2 0 2 9 13 2
8 9 7 9 10 14 10 13 2
33 0 9 2 15 11 1 9 1 0 13 15 9 2 9 2 9 1 9 7 9 1 9 2 9 2 9 7 9 1 0 9 13 2
36 15 1 0 9 1 9 7 9 1 9 2 9 1 9 2 11 11 7 11 9 1 9 2 0 0 9 7 3 1 3 13 4 0 9 13 2
12 9 1 9 1 1 11 9 13 9 13 4 2
8 11 1 9 14 10 9 13 2
11 9 7 9 1 9 10 9 1 13 4 2
11 9 1 0 9 7 9 1 9 14 13 2
15 9 9 1 14 9 1 9 1 9 1 14 9 13 4 2
23 11 1 9 13 1 15 0 9 15 13 4 2 15 0 9 0 9 1 13 4 4 4 2
14 11 11 9 9 1 14 9 1 10 9 13 4 4 2
26 9 1 3 0 9 9 1 9 1 9 1 1 12 9 1 9 11 1 9 13 1 9 13 4 4 2
32 11 1 12 0 9 1 0 9 1 1 11 1 9 1 13 14 12 9 9 2 9 1 9 1 1 9 1 9 13 4 4 2
17 10 9 1 15 9 9 1 14 12 9 1 1 9 1 13 4 2
24 11 11 11 11 11 1 1 9 2 9 1 1 1 11 1 0 9 1 9 0 13 4 4 2
32 11 11 11 11 1 9 11 11 1 1 0 10 9 1 1 9 1 13 4 9 9 1 10 9 9 1 0 9 0 13 4 2
36 11 1 1 11 7 11 1 1 12 9 0 11 1 13 1 1 9 14 12 13 2 7 15 10 9 1 10 9 9 1 10 9 13 4 4 2
27 11 11 1 13 0 9 11 11 1 11 1 9 13 4 13 16 15 9 1 15 3 13 9 1 9 13 2
9 1 15 2 15 15 9 14 13 2
17 10 9 11 1 15 9 1 11 1 13 9 1 0 13 4 13 2
34 15 1 15 9 1 15 9 1 14 13 4 1 9 14 13 2 15 1 9 11 11 7 11 1 9 11 11 1 1 0 9 14 13 2
19 11 1 13 16 15 9 1 13 9 1 9 15 9 1 9 9 14 13 2
18 15 15 10 9 14 13 2 15 15 15 7 9 1 15 9 13 4 2
25 15 15 9 1 14 13 1 9 13 4 13 16 11 2 11 7 11 1 14 9 9 1 13 4 2
12 15 2 15 1 15 9 13 1 9 13 4 2
25 11 1 13 16 11 12 0 9 13 2 15 9 11 11 2 11 11 11 7 11 11 1 13 4 2
20 15 0 9 1 13 9 1 0 9 1 13 16 15 10 9 9 13 4 4 2
8 15 10 0 9 1 9 13 2
15 10 9 1 9 13 1 1 15 15 15 1 0 13 4 2
14 11 11 1 9 11 11 1 14 9 1 0 9 13 2
18 11 11 1 1 2 15 0 9 11 11 11 7 0 9 1 9 13 2
12 10 0 9 1 9 13 1 15 9 13 4 2
12 7 3 15 9 11 1 15 9 1 1 13 2
24 9 1 9 1 13 9 1 1 1 15 13 13 16 9 1 9 1 15 9 1 10 9 13 2
22 10 9 15 9 1 13 4 2 15 1 3 12 11 11 0 11 9 1 1 13 4 2
25 7 2 9 1 1 15 1 13 16 15 11 11 1 9 11 11 1 13 1 14 15 13 4 4 2
14 11 9 1 1 9 14 11 11 1 13 1 14 13 2
12 7 11 11 15 10 9 1 9 1 14 13 2
13 11 11 11 12 9 3 9 1 9 13 4 4 2
24 15 15 15 14 9 9 13 13 4 4 2 16 15 0 9 15 9 1 9 13 4 4 4 2
19 11 1 11 11 11 11 1 11 1 11 11 1 9 1 9 1 9 13 2
19 15 1 11 1 11 11 9 1 9 13 4 4 16 9 1 9 13 4 2
22 0 9 1 13 4 4 4 16 11 1 10 9 13 11 1 0 9 1 9 13 4 2
24 11 11 1 1 1 11 10 9 0 14 13 4 4 2 15 10 9 1 13 9 1 13 4 2
15 13 4 4 15 15 9 1 0 9 1 8 0 9 13 2
9 9 1 11 9 11 1 13 4 2
12 11 9 1 11 1 13 7 9 1 9 13 2
26 15 9 1 0 13 4 15 3 11 11 11 1 9 13 7 15 13 1 11 11 1 13 1 0 13 2
7 15 0 9 14 13 4 2
16 11 9 14 11 1 11 9 1 9 13 1 9 13 4 4 2
17 15 11 11 1 11 2 11 9 1 1 14 15 9 13 4 4 2
24 11 9 1 10 2 9 2 1 0 11 1 11 9 1 11 1 9 1 13 1 9 13 4 2
16 11 1 13 11 1 9 1 9 1 10 9 2 9 13 4 2
22 9 15 1 13 4 16 11 11 11 1 12 9 1 11 1 15 9 13 13 4 4 2
6 15 13 9 0 13 2
20 15 1 11 11 9 1 13 4 2 15 9 11 11 11 11 1 13 13 4 2
18 15 1 9 15 13 4 16 11 1 1 11 9 12 13 4 4 4 2
18 7 11 11 11 1 10 9 13 4 11 11 11 11 1 10 9 13 2
14 11 1 9 1 11 11 1 14 9 1 9 13 4 2
23 11 11 11 1 11 2 11 1 0 9 9 1 11 1 10 0 9 1 0 9 13 4 2
15 15 13 13 16 11 11 1 10 9 12 10 0 9 13 2
51 11 1 11 1 9 11 11 1 11 11 11 11 1 0 11 1 12 9 13 4 9 13 4 16 15 10 9 1 9 13 4 11 11 1 12 9 0 0 2 0 0 9 1 3 9 13 9 1 0 13 2
26 15 13 13 16 12 9 0 10 9 10 9 1 11 1 11 11 1 1 11 7 11 1 13 4 4 2
16 10 9 12 9 13 4 4 15 1 12 9 15 14 0 13 2
20 11 2 11 1 0 9 1 9 1 10 9 1 0 14 14 13 4 4 4 2
42 0 9 2 9 7 0 9 1 12 0 9 11 11 11 1 13 16 11 1 0 0 9 1 0 9 1 9 7 9 9 7 9 1 9 0 9 1 1 13 4 4 2
20 3 11 1 9 13 4 11 7 0 0 9 1 10 9 1 9 14 14 13 2
31 11 1 13 16 0 9 1 0 11 11 1 11 11 11 1 1 11 11 1 11 11 2 11 1 14 0 13 4 4 4 2
21 11 7 11 11 1 1 13 10 9 1 9 1 1 0 9 1 0 13 4 4 2
19 15 13 16 10 9 1 13 4 9 12 9 1 12 9 1 0 13 4 2
19 11 1 1 13 9 11 9 1 0 11 7 11 9 1 9 9 13 4 2
30 15 13 16 11 1 9 1 1 11 7 11 9 1 14 11 11 1 0 13 1 11 1 10 9 1 9 13 4 4 2
9 15 15 3 14 9 13 4 4 2
27 11 1 13 16 11 1 15 0 9 11 11 1 9 13 4 2 10 9 11 1 15 0 13 4 4 4 2
29 11 11 1 11 1 3 9 13 1 9 1 0 13 4 11 1 13 16 15 10 9 1 9 13 1 15 9 13 2
12 11 11 1 11 1 9 1 3 14 13 4 2
20 11 11 11 1 1 11 11 1 9 13 1 9 1 9 1 9 13 4 4 2
22 9 9 1 13 13 16 11 11 1 11 1 1 11 11 1 9 12 9 1 13 4 2
19 16 0 9 1 13 4 16 9 1 13 1 1 10 9 13 4 4 4 2
25 11 1 9 9 9 1 0 9 1 13 1 3 15 9 2 9 1 13 1 9 1 13 4 4 2
33 11 11 1 11 11 11 11 1 1 11 11 1 9 1 9 12 9 13 1 9 1 9 1 0 9 1 13 1 9 1 9 13 2
23 11 11 11 1 0 9 9 11 11 1 10 9 1 9 9 9 1 13 1 9 13 4 2
23 15 13 16 11 1 9 1 9 9 13 4 7 9 11 11 1 1 0 9 1 13 4 2
14 9 13 1 1 1 15 13 16 15 12 0 9 13 2
11 7 9 1 9 1 15 9 0 9 13 2
8 9 10 10 0 13 4 4 2
9 10 9 9 1 0 9 1 13 2
13 10 9 1 9 12 1 12 11 11 1 1 13 2
16 11 1 10 9 1 15 9 1 9 1 9 1 9 13 4 2
32 11 1 13 16 9 9 1 1 13 1 9 1 9 1 9 9 1 1 9 1 10 1 13 1 1 15 15 10 9 14 13 2
9 11 1 10 9 1 0 9 13 2
12 15 15 14 13 16 10 9 15 1 13 4 2
13 11 1 11 11 1 9 1 12 9 0 13 4 2
19 0 9 15 0 13 4 15 11 11 11 9 1 9 1 0 13 4 4 2
18 9 1 9 1 11 1 9 9 1 9 9 1 9 9 13 4 4 2
18 10 9 9 14 15 1 0 9 13 4 7 0 15 0 9 13 4 2
16 10 9 1 13 13 16 10 9 1 9 1 14 15 13 4 2
12 10 9 9 15 1 9 13 9 13 13 4 2
37 9 1 0 9 11 11 11 11 2 11 2 1 13 13 16 15 0 14 14 16 0 7 0 9 1 13 1 9 1 1 9 1 9 1 0 13 2
9 15 13 4 16 9 1 9 13 2
41 11 0 10 9 1 9 11 11 11 13 4 16 9 1 13 16 15 0 2 0 7 0 9 1 9 1 9 13 10 9 1 9 1 13 1 9 1 0 9 13 2
7 15 15 1 1 0 13 2
13 15 12 9 7 9 9 1 1 15 14 13 4 2
18 16 15 1 13 4 4 16 15 9 7 9 1 15 9 14 13 4 2
29 0 13 16 0 11 1 11 11 11 1 9 1 13 9 1 1 9 3 11 11 1 9 9 0 9 13 4 4 2
30 9 1 15 13 0 9 13 1 13 16 3 1 9 1 9 1 0 9 1 10 0 9 1 9 13 1 9 15 13 2
28 10 9 9 15 1 0 9 13 4 16 10 9 1 1 9 1 12 2 12 9 1 9 1 0 9 13 4 2
23 10 12 9 1 9 13 1 11 13 1 9 13 4 10 9 1 15 9 1 9 13 4 2
22 11 11 11 9 13 4 13 4 16 10 9 1 9 9 1 9 1 14 0 13 4 2
11 15 9 1 1 13 1 15 9 14 13 2
9 9 9 1 0 9 1 9 13 2
35 11 11 11 11 11 2 11 2 1 9 11 11 11 2 15 9 1 0 9 1 9 13 4 2 1 9 9 1 1 0 9 1 0 13 2
9 9 1 14 9 15 0 14 13 2
13 15 1 10 0 9 7 9 1 14 9 13 4 2
11 15 1 14 9 9 1 14 9 13 4 2
10 7 10 15 0 9 9 1 9 13 2
8 15 15 9 13 1 14 13 2
20 11 1 0 9 11 11 1 13 13 16 10 9 14 0 9 9 1 14 13 2
24 10 9 1 9 10 9 7 9 1 1 13 4 2 10 9 1 10 9 1 0 9 13 4 2
14 15 0 9 1 9 13 1 1 15 9 13 4 4 2
19 15 9 1 1 9 13 13 4 16 9 1 10 9 15 9 1 0 13 2
13 9 15 14 13 16 15 0 9 1 1 9 13 2
18 15 9 13 16 15 9 14 13 4 15 9 9 9 13 4 4 4 2
28 11 11 11 1 9 11 11 11 1 14 9 13 16 9 10 9 7 0 9 1 9 13 10 9 1 9 13 2
22 7 11 9 11 11 11 14 10 9 1 9 9 1 9 1 9 13 1 13 4 4 2
49 10 9 1 1 16 11 11 9 11 11 1 11 1 9 1 11 9 1 9 1 9 1 13 1 13 4 2 11 1 9 13 4 16 15 11 3 13 13 4 7 15 1 10 9 1 13 13 4 2
29 11 1 12 0 9 1 9 1 9 9 0 13 4 11 11 9 11 11 1 13 16 15 9 13 16 15 15 13 2
21 15 11 1 10 9 1 13 13 4 15 15 9 9 1 9 13 1 9 13 4 2
27 9 1 11 0 9 1 15 13 1 9 1 9 13 4 1 1 1 13 4 9 1 11 1 10 9 13 2
13 15 0 9 11 1 11 1 9 1 0 13 4 2
25 2 11 11 11 2 0 9 1 9 1 1 11 11 11 1 11 1 11 0 9 1 13 1 13 2
12 15 13 13 16 9 15 0 9 13 4 4 2
22 9 7 0 9 1 0 10 9 9 9 9 1 13 9 1 0 9 13 13 4 4 2
20 10 9 1 0 13 4 9 1 3 2 3 13 1 9 1 9 13 4 4 2
18 0 9 1 15 15 13 1 3 15 15 0 9 1 9 9 13 4 2
18 15 1 15 9 1 9 13 7 11 11 11 15 10 9 13 13 4 2
7 11 1 3 0 9 13 2
14 15 11 1 9 14 11 1 11 11 0 13 4 4 2
19 15 9 1 9 0 13 16 11 9 1 13 9 1 0 9 13 13 4 2
24 15 14 0 9 15 13 16 15 9 1 15 9 7 9 1 15 9 1 1 1 13 13 4 2
13 3 15 10 14 10 9 9 1 9 13 13 4 2
20 11 11 9 11 1 9 1 13 14 9 1 13 9 1 0 9 9 13 4 2
9 15 9 1 9 1 0 9 13 2
12 9 1 12 9 15 14 9 1 9 13 4 2
19 3 10 9 9 1 15 11 2 11 7 0 0 9 14 9 13 4 4 2
18 11 11 1 9 13 4 12 9 13 4 16 10 9 0 9 13 4 2
12 9 9 1 9 9 13 7 13 1 0 13 2
18 10 3 9 13 7 3 3 10 3 1 13 7 3 1 0 13 4 2
13 15 1 9 0 13 2 15 15 1 9 14 13 2
19 9 1 13 16 10 14 9 1 9 13 9 13 4 7 15 9 13 4 2
23 15 9 13 13 2 7 10 15 15 10 9 1 13 16 9 1 1 15 9 14 14 13 2
27 9 1 0 13 12 9 1 13 15 13 4 16 16 15 0 9 1 9 1 13 9 1 13 4 4 4 2
22 10 14 9 7 15 9 1 9 0 9 1 9 1 13 7 15 9 13 4 4 4 2
12 0 10 9 1 12 9 1 13 4 4 4 2
16 3 10 14 9 13 4 16 10 9 15 0 9 1 13 4 2
8 11 1 9 1 3 9 13 2
18 9 9 1 0 0 9 1 11 1 13 16 9 1 15 1 9 13 2
22 9 9 1 1 0 13 1 11 11 1 9 13 16 0 11 9 9 1 9 13 4 2
26 9 1 13 4 9 1 9 1 9 13 4 11 1 13 16 9 1 10 9 1 0 9 15 1 13 2
15 15 15 14 9 13 16 15 9 1 10 0 9 13 4 2
23 15 13 16 9 1 13 4 9 1 9 1 11 11 11 1 12 12 9 1 9 13 4 2
19 11 0 9 1 13 11 9 14 13 7 15 1 9 1 9 1 9 13 2
17 11 11 1 12 9 1 0 9 1 9 0 11 11 1 9 13 2
24 11 1 13 9 11 1 15 13 16 0 9 9 14 13 1 12 0 9 1 10 9 0 13 2
11 15 10 14 9 11 1 13 14 13 4 2
8 15 0 9 1 9 10 13 2
21 15 13 16 0 12 9 1 15 10 15 13 4 2 15 15 9 1 9 13 4 2
21 9 1 9 13 11 11 9 13 11 1 15 9 1 11 1 13 1 9 13 4 2
7 15 15 15 14 13 13 2
5 15 9 14 13 2
13 10 9 1 9 1 9 9 1 3 13 4 4 2
30 11 1 11 7 11 15 3 0 13 4 4 7 9 11 1 11 9 9 1 9 13 4 2 7 15 9 0 14 13 2
14 16 15 1 1 10 9 1 9 3 0 13 4 4 2
19 15 0 9 12 9 9 8 13 4 2 15 0 9 1 12 9 3 13 2
21 11 11 2 11 2 11 2 11 7 11 11 1 10 9 9 7 9 1 0 13 2
15 10 9 11 7 11 1 10 9 1 9 13 1 9 13 2
21 9 11 1 9 14 12 9 11 9 1 9 1 1 13 4 1 9 13 4 4 2
14 9 9 1 13 16 9 1 1 1 15 9 14 13 2
28 9 9 1 12 9 1 13 16 11 1 9 0 9 12 9 9 8 13 4 15 10 9 1 1 1 0 13 2
10 15 0 9 12 9 9 8 13 4 2
60 9 1 1 0 13 1 9 1 11 1 11 1 1 13 1 11 9 2 11 1 11 1 1 13 1 11 9 2 11 1 11 1 1 13 1 11 9 2 11 1 11 1 1 13 1 11 11 9 7 11 1 11 1 1 13 1 11 9 13 2
36 9 9 1 0 12 9 1 11 1 10 9 1 0 9 7 11 7 11 1 10 9 1 0 9 7 9 1 1 9 13 1 9 0 13 4 2
27 9 1 11 1 11 11 11 2 11 2 0 13 1 1 11 11 1 12 9 1 9 13 1 9 13 4 2
39 11 11 11 11 11 1 9 11 11 1 11 1 12 9 1 0 9 1 1 9 1 13 16 15 0 11 1 11 11 1 11 11 1 12 9 1 9 13 2
10 10 3 9 9 1 10 9 0 13 2
28 9 1 10 9 13 4 11 0 13 1 9 13 15 9 9 1 10 0 9 9 1 14 0 13 1 9 13 2
16 15 13 16 15 15 14 9 1 13 7 11 1 9 14 13 2
17 16 15 9 0 14 13 16 9 1 1 0 9 9 13 4 4 2
14 15 13 16 9 10 9 9 1 11 11 1 9 13 2
19 11 2 11 1 11 1 13 9 1 11 11 11 1 15 9 14 13 4 2
21 15 1 1 12 9 1 13 16 9 1 9 1 1 9 14 15 9 1 0 13 2
24 11 11 11 11 1 9 9 9 9 11 11 1 13 16 9 1 9 1 15 9 14 13 4 2
16 9 1 1 11 11 1 9 1 1 9 12 9 13 4 4 2
9 9 0 9 1 9 13 4 4 2
18 15 13 16 9 1 1 15 1 12 12 9 1 9 1 9 13 4 2
22 9 9 11 11 1 11 1 13 0 9 1 13 4 9 1 1 0 9 0 13 4 2
39 11 1 9 1 9 11 11 11 7 9 9 1 9 9 11 11 1 0 2 0 13 4 9 1 11 1 9 1 13 9 7 9 1 0 9 0 13 4 2
28 11 1 11 1 9 7 9 1 1 1 9 0 13 4 13 4 16 9 1 10 9 1 0 9 15 1 13 2
32 9 9 9 1 0 9 1 1 11 1 13 9 9 1 13 4 2 15 0 9 13 16 11 1 9 3 13 10 9 1 9 13
11 11 11 11 15 9 1 1 13 4 4 2
12 15 0 9 1 9 1 9 1 13 4 4 2
20 10 9 1 0 9 1 9 1 9 9 1 13 1 14 9 9 13 4 4 2
22 9 1 9 13 16 12 9 1 1 10 9 0 13 4 4 7 9 9 1 13 4 2
57 0 9 1 9 1 9 2 9 2 9 7 0 9 1 1 0 13 7 15 14 13 1 9 7 9 1 9 1 1 9 1 9 1 11 11 11 2 9 9 2 9 9 9 9 2 9 2 9 7 0 0 9 1 9 13 4 2
18 10 9 1 9 14 13 2 15 11 11 11 1 10 9 13 4 4 2
30 10 3 10 9 14 13 16 10 9 1 9 9 1 14 13 4 4 7 15 9 14 13 7 9 13 1 10 9 13 2
17 10 3 9 9 1 9 13 7 9 1 15 13 1 9 13 4 2
15 10 9 1 1 0 0 9 1 14 9 1 13 4 4 2
45 9 1 1 9 1 9 1 10 9 1 9 1 1 13 1 9 7 0 9 0 13 4 2 7 0 2 0 9 1 1 11 1 13 0 15 14 9 1 9 9 1 1 13 4 2
28 11 11 1 11 11 1 0 9 1 9 9 0 13 4 4 2 3 15 1 11 1 14 12 9 0 13 4 2
26 10 9 1 1 15 14 9 9 13 4 16 3 10 9 1 10 9 1 9 9 1 14 13 4 4 2
47 11 1 13 4 16 11 2 11 1 11 11 11 1 9 3 13 1 1 13 9 1 9 1 12 9 1 1 13 4 9 9 1 0 9 1 9 14 13 2 7 15 0 9 13 4 4 2
31 11 1 9 9 1 9 11 11 1 11 1 12 9 1 13 16 9 9 1 11 1 9 0 9 1 14 15 9 14 13 2
17 15 13 16 12 9 0 9 13 1 9 13 1 9 13 4 4 2
16 15 9 13 7 9 13 1 9 1 1 0 9 1 13 4 2
40 15 13 16 15 0 9 1 11 1 14 9 13 4 4 16 10 9 9 1 1 15 14 13 4 4 16 0 9 7 9 1 11 11 0 9 14 13 4 4 2
25 12 9 1 9 1 15 13 16 9 1 10 9 1 13 15 9 13 7 15 15 0 9 14 13 2
17 15 9 1 15 11 1 1 13 4 7 15 15 0 13 4 4 2
28 15 13 16 11 1 11 1 14 15 0 13 4 16 0 9 1 9 14 13 1 11 11 1 1 15 13 4 2
19 15 13 16 9 1 13 9 1 9 1 9 1 13 14 15 0 9 13 2
27 0 0 9 1 9 9 1 9 1 9 13 1 1 11 1 11 9 1 0 9 9 1 9 13 4 4 2
15 9 1 9 1 9 9 1 14 12 9 1 1 13 4 2
14 9 1 3 0 0 13 1 12 9 1 13 4 4 2
38 9 1 9 9 9 11 11 1 11 1 13 16 14 12 9 9 1 0 0 9 1 10 9 1 9 1 9 1 1 0 0 9 1 9 13 4 4 2
26 11 1 13 16 9 1 13 4 9 1 9 13 1 1 10 9 1 0 9 9 1 9 13 4 4 2
18 15 15 14 13 16 10 9 1 9 1 9 3 10 0 13 4 4 2
21 2 15 9 1 0 9 13 7 10 9 1 9 1 9 1 9 14 13 4 4 2
32 9 1 9 1 9 1 3 14 0 13 1 1 0 9 1 3 0 9 1 13 4 7 10 9 1 10 14 10 12 9 13 4
30 11 1 12 9 1 9 0 12 0 9 1 14 12 0 2 0 9 1 9 1 12 9 7 9 1 12 9 0 13 2
31 0 13 16 11 11 1 13 0 0 9 1 10 9 1 14 12 9 13 4 4 7 12 9 0 0 9 1 9 13 4 2
31 11 1 13 16 15 15 14 9 1 13 1 10 9 1 9 13 4 4 7 9 9 11 11 1 9 1 3 14 0 13 2
23 15 3 13 16 16 15 0 9 1 9 13 2 15 15 13 1 1 9 1 9 13 4 2
25 0 9 1 11 11 11 1 11 1 11 11 11 1 1 11 1 9 1 9 13 1 9 13 4 2
31 2 11 11 11 11 11 2 1 13 13 16 11 11 1 11 1 9 13 1 1 0 11 1 3 0 9 1 9 13 4 2
25 11 1 11 0 11 11 11 1 11 1 13 11 11 1 1 10 9 1 9 13 1 9 13 4 2
18 15 0 11 1 14 11 11 1 10 9 1 9 13 1 9 13 4 2
37 11 1 11 1 11 9 1 1 11 9 1 13 9 1 9 13 4 0 11 11 11 11 1 13 16 15 14 9 11 1 9 1 9 14 13 4 2
13 9 1 1 1 11 1 9 11 1 1 0 13 2
21 15 13 16 11 9 1 9 10 9 13 4 4 15 0 9 11 11 1 9 13 2
26 11 1 13 4 4 9 9 1 9 13 4 15 13 16 10 9 9 11 1 1 0 9 13 4 4 2
28 0 11 11 1 13 16 9 9 1 9 0 13 1 3 0 9 9 1 1 15 9 0 9 1 13 4 4 2
21 10 9 11 1 0 9 7 9 1 9 1 13 1 10 9 1 9 13 4 4 2
14 1 11 2 11 1 1 14 11 1 0 9 13 4 2
9 7 11 1 9 15 10 3 13 2
19 15 2 11 1 11 1 9 1 1 10 9 1 9 1 1 13 4 4 2
23 0 9 9 11 11 11 1 13 13 16 11 11 1 9 1 9 1 9 9 1 13 4 2
16 11 1 11 1 11 11 1 1 9 13 1 1 9 13 4 2
15 16 2 11 11 15 11 1 1 9 1 9 13 4 4 2
30 11 1 13 16 11 1 9 10 12 0 9 1 0 13 15 11 7 11 1 9 1 1 11 1 9 1 1 13 4 2
16 7 3 1 11 11 1 10 9 1 9 13 1 9 13 4 2
19 11 1 9 1 9 13 4 15 13 16 11 1 9 1 9 1 13 4 2
12 11 11 10 9 11 1 1 9 13 4 4 2
12 15 9 1 11 1 1 0 0 13 4 4 2
23 10 9 1 9 9 11 11 1 13 16 15 9 11 1 1 3 0 9 13 4 4 4 2
16 7 15 11 2 11 9 2 9 1 9 1 9 13 4 4 2
23 11 11 1 13 16 11 11 11 1 1 1 0 9 1 15 14 13 1 1 0 14 13 2
22 16 15 13 4 16 11 1 1 1 15 14 9 15 11 1 9 1 9 13 4 4 2
12 7 9 1 11 1 9 1 9 14 13 4 2
16 11 1 11 1 9 1 1 14 15 9 11 1 13 4 4 2
26 11 11 1 11 1 9 9 13 1 9 1 0 13 1 3 15 15 9 1 9 9 1 9 13 4 2
32 11 11 1 9 13 16 0 9 9 7 11 11 1 13 4 4 10 0 9 1 1 9 1 9 1 0 9 1 9 0 13 2
13 10 9 11 1 11 11 11 11 11 11 1 13 2
18 15 13 16 11 2 11 1 9 1 12 12 9 9 1 9 13 4 2
12 15 9 9 1 12 12 9 9 1 9 13 2
22 0 9 1 0 9 9 7 0 9 1 9 1 13 4 11 1 1 0 9 0 13 2
17 10 9 11 11 1 1 9 9 1 1 12 12 9 9 0 13 2
16 7 9 9 1 1 12 12 9 9 11 11 1 1 13 4 2
26 15 0 13 16 11 11 1 0 9 1 15 1 15 14 9 1 1 9 1 9 1 9 14 13 4 2
16 11 1 13 16 0 9 1 9 1 9 11 11 1 13 4 2
40 9 9 1 3 13 1 9 1 0 13 4 1 9 1 9 1 9 13 1 9 1 13 10 9 1 15 13 16 9 1 15 1 1 3 15 9 14 13 4 2
24 11 9 1 11 9 1 11 9 1 12 9 11 11 14 11 1 9 1 9 9 1 13 4 2
15 11 1 9 1 15 9 9 13 12 12 9 1 9 13 2
16 9 1 9 13 1 3 1 11 1 9 1 9 9 1 13 2
13 9 1 9 1 9 0 13 9 9 13 4 4 2
16 0 13 16 11 1 9 9 9 11 11 0 9 1 0 13 2
8 15 10 9 11 1 0 13 2
23 0 9 1 11 1 11 9 1 13 1 11 11 1 9 7 0 9 11 1 14 13 4 2
19 11 11 1 0 9 11 14 11 11 1 11 9 1 11 11 1 9 13 2
17 15 11 1 9 13 13 4 2 7 15 1 1 13 9 14 13 2
17 15 9 0 14 13 4 7 9 12 9 9 13 1 9 13 4 2
23 11 1 9 1 15 15 13 9 14 13 15 11 1 15 9 1 15 9 11 9 1 13 2
13 9 1 9 1 9 1 9 1 9 0 13 4 2
31 9 1 1 11 9 14 12 9 11 1 11 0 9 1 9 1 9 13 15 9 1 9 13 4 12 12 9 1 9 13 2
17 9 1 13 16 16 9 14 13 16 2 15 14 2 13 4 4 2
16 9 1 9 11 2 11 2 1 3 13 1 1 13 4 4 2
18 9 13 1 3 9 1 9 1 9 1 9 1 9 1 13 4 4 2
33 13 4 4 16 11 1 10 9 1 9 1 9 13 15 9 9 13 4 4 2 7 15 10 9 14 13 15 9 1 9 13 4 2
33 11 0 9 1 9 13 1 13 4 4 4 16 15 1 9 9 1 11 1 13 4 7 14 10 9 1 15 9 1 14 9 13 2
19 9 1 9 13 11 1 10 9 15 9 9 0 9 1 0 13 4 4 2
15 10 9 1 11 11 1 9 11 11 1 14 13 4 4 2
23 10 9 1 9 2 3 10 9 1 9 14 13 4 7 15 1 15 9 14 13 4 4 2
14 9 0 9 1 0 13 1 1 0 9 13 4 4 2
22 11 2 11 1 1 9 1 9 13 4 11 11 11 1 11 1 9 9 13 4 4 2
13 10 9 1 14 12 9 1 15 9 0 14 13 2
30 9 1 9 13 1 9 1 9 12 9 1 0 13 4 4 2 7 15 1 11 11 10 9 1 9 0 13 4 4 2
15 0 13 16 15 14 9 1 1 9 1 9 0 13 4 2
18 9 1 0 13 1 9 1 13 9 1 13 1 9 9 1 13 4 2
21 9 1 1 16 15 9 1 9 13 4 16 15 15 1 9 1 14 0 13 4 2
20 9 1 12 9 1 1 9 1 10 0 9 11 11 1 0 9 1 0 13 2
31 9 1 13 16 11 1 11 1 9 13 1 10 9 1 9 1 9 11 11 1 0 13 4 2 7 15 1 14 13 4 2
46 12 9 1 1 13 9 1 1 11 1 11 7 11 1 11 1 13 1 10 9 1 12 2 12 9 1 11 2 11 7 11 2 11 1 12 9 1 9 9 2 9 1 9 13 4 2
11 0 9 1 10 9 11 1 9 1 13 2
21 15 9 11 11 11 1 0 13 4 2 10 9 15 11 1 11 1 14 13 4 2
29 9 1 13 13 16 10 9 1 11 11 1 10 9 0 14 13 4 4 4 2 7 15 9 1 9 14 13 4 2
39 0 9 1 13 13 16 16 15 10 9 14 12 2 12 9 1 13 2 7 12 9 1 9 1 9 13 1 1 12 9 1 14 10 0 7 9 13 4 2
27 11 11 11 11 1 1 1 11 11 1 0 9 0 13 1 11 1 9 1 11 11 1 0 9 13 4 2
19 15 9 13 4 16 11 9 11 9 11 11 1 9 1 9 13 4 4 2
19 11 1 9 1 1 13 9 1 1 15 11 11 11 11 1 9 9 13 2
16 11 1 11 1 13 16 10 9 1 15 0 9 13 4 4 2
14 9 9 1 13 9 1 11 11 1 11 1 13 4 2
16 15 1 11 11 1 11 11 1 9 9 13 1 9 13 4 2
13 9 1 0 9 1 10 9 11 11 1 9 13 2
7 15 1 9 1 9 13 2
17 11 11 1 9 9 1 0 9 13 7 11 11 1 9 13 4 2
11 11 1 0 9 1 9 1 9 13 4 2
40 15 1 9 1 15 9 1 13 16 9 1 1 11 1 15 9 0 13 4 4 4 7 9 9 14 9 13 4 4 2 15 15 9 0 13 1 9 14 13 2
28 9 1 13 16 9 1 9 1 10 9 13 4 4 16 15 10 9 1 9 13 7 15 1 9 13 13 4 2
56 9 11 11 11 7 9 11 11 11 1 9 1 9 9 7 11 11 1 9 1 9 1 9 1 0 11 11 1 13 4 9 1 13 1 9 13 1 9 1 10 9 1 13 1 3 15 3 1 9 1 9 13 9 1 13 2
27 11 11 1 1 1 0 9 11 11 1 13 16 9 13 4 4 16 9 9 1 1 14 13 4 4 4 2
42 9 9 1 1 1 9 11 11 1 13 16 12 9 9 9 9 13 4 16 9 1 11 2 11 11 11 1 1 11 11 1 15 14 9 9 9 1 9 14 13 4 2
50 9 0 9 1 13 4 1 9 13 2 0 9 1 1 9 13 1 9 7 0 9 11 11 1 1 1 0 9 11 11 1 13 16 0 9 1 1 0 9 9 1 9 0 13 0 9 1 1 13 2
20 0 9 11 1 1 1 0 9 11 11 11 1 13 16 9 9 0 13 4 2
33 9 1 10 9 1 13 1 3 15 3 1 9 1 9 13 9 13 4 11 1 12 9 1 1 13 1 9 1 1 9 0 13 2
9 11 1 9 9 1 9 13 4 2
46 0 9 1 1 9 1 1 9 1 10 9 1 9 13 1 9 0 13 7 11 11 11 1 9 13 9 1 10 9 1 9 13 1 9 13 4 14 9 13 1 9 13 4 4 4 2
22 11 1 10 9 9 1 9 1 9 0 13 1 0 9 1 9 1 0 13 4 4 2
16 10 9 1 9 11 9 1 9 1 9 0 13 1 13 4 2
19 11 1 9 9 1 9 13 1 9 7 9 1 0 9 0 13 4 4 2
13 11 11 11 1 9 14 10 9 1 13 4 4 2
37 9 1 11 2 11 11 1 9 1 10 9 11 11 1 9 1 9 7 9 1 10 12 9 1 0 13 2 15 10 9 1 13 9 14 0 13 2
18 9 1 15 9 1 12 12 9 1 9 1 11 2 11 11 13 4 2
16 10 9 11 1 13 9 1 9 1 9 13 1 13 4 4 2
18 9 1 9 1 1 11 1 13 9 1 9 1 9 3 10 13 4 2
10 15 1 10 9 9 1 10 0 13 2
7 9 7 9 15 9 13 2
18 9 1 1 3 10 9 1 10 9 12 9 9 9 1 9 0 13 2
13 11 1 13 9 1 9 14 9 14 12 9 13 2
21 3 11 11 1 14 15 9 9 1 11 1 13 9 1 9 13 1 9 13 4 2
31 9 1 1 11 11 1 12 9 11 11 11 11 11 1 12 0 9 9 1 9 1 10 9 1 9 13 1 9 13 4 2
17 15 1 14 11 11 1 11 1 9 1 9 14 9 13 4 4 2
16 11 9 9 1 1 12 9 9 1 11 1 9 13 4 4 2
17 0 9 11 9 9 1 1 12 9 9 1 11 1 9 13 4 2
17 9 1 13 13 16 10 9 9 7 9 1 0 9 13 4 4 2
16 11 11 1 9 1 11 1 14 12 9 0 13 1 9 13 2
28 15 1 9 1 0 13 4 4 4 7 16 15 15 0 2 0 13 16 14 12 9 1 10 9 0 13 4 2
16 11 11 1 1 14 10 9 1 0 9 1 9 9 13 4 2
13 11 11 9 1 9 1 10 9 1 9 13 4 2
28 9 1 9 7 9 9 1 9 11 11 1 9 13 16 10 9 14 11 11 1 1 9 14 1 0 13 4 2
15 11 1 13 16 10 9 0 12 9 1 13 0 13 4 2
15 14 12 2 12 9 9 1 1 10 9 1 9 13 4 2
20 9 9 0 13 1 9 9 1 0 2 0 9 9 11 11 1 13 4 4 2
20 11 11 11 2 11 11 11 11 7 11 11 11 1 9 1 9 13 4 4 2
13 3 1 15 0 2 0 0 9 1 14 9 13 2
12 15 11 11 7 11 11 1 9 14 0 13 2
16 9 9 1 9 13 16 15 11 11 11 1 1 14 9 13 2
20 0 13 16 10 9 14 12 12 9 11 11 11 1 13 9 1 9 13 4 2
13 15 11 1 3 0 9 1 1 12 13 4 4 2
12 11 1 9 1 0 9 1 9 11 1 13 2
24 11 11 1 13 0 9 1 9 1 1 15 9 14 9 9 1 15 0 9 1 9 14 13 2
17 0 9 9 11 1 9 9 1 1 14 15 1 0 13 4 4 2
16 10 9 15 3 1 1 9 1 9 1 9 14 14 13 4 2
12 11 1 10 12 12 9 15 9 1 9 13 2
23 0 9 1 1 13 1 9 1 9 9 1 12 9 1 1 12 9 1 9 1 9 13 2
22 9 1 12 9 9 1 0 7 0 9 1 1 11 11 1 12 9 1 0 13 4 2
58 11 1 9 1 10 0 9 1 9 1 9 13 2 15 11 11 11 2 11 2 1 9 7 11 9 1 9 11 11 2 12 9 11 13 4 7 0 11 2 11 2 9 11 11 11 2 11 11 11 11 7 11 11 11 11 0 13 2
14 9 1 15 9 9 1 0 9 1 0 9 13 4 2
10 9 1 0 9 1 9 0 14 13 2
19 9 1 9 0 13 2 9 9 1 9 0 13 7 9 12 0 9 13 2
10 9 1 0 9 1 9 1 9 13 2
12 9 1 11 7 11 9 1 14 10 9 13 2
24 0 9 1 9 2 11 2 1 11 9 1 9 9 1 9 1 13 1 9 13 4 4 4 2
43 9 1 9 14 1 11 1 12 9 9 1 9 1 13 9 1 0 9 0 13 4 1 3 11 1 12 9 9 1 9 1 1 9 1 1 1 14 9 1 9 13 4 2
20 11 9 11 11 1 11 1 9 1 12 9 9 1 9 1 11 1 13 4 2
39 11 1 9 1 9 9 1 15 12 10 9 13 15 11 1 11 11 11 11 11 1 11 11 1 1 13 1 15 14 9 1 9 1 9 1 0 13 4 2
17 11 1 9 1 9 1 9 1 1 7 3 1 9 13 4 4 2
21 15 1 11 9 1 9 1 9 9 1 9 13 1 3 10 9 13 4 4 4 2
23 0 13 16 9 1 11 1 9 1 12 9 9 1 9 9 1 1 0 9 0 13 4 2
37 11 1 12 9 9 1 1 11 11 1 11 11 1 13 4 9 1 9 1 11 11 11 11 11 1 11 1 9 1 9 1 1 15 9 0 13 2
12 11 1 9 13 16 11 9 13 1 9 13 2
20 0 13 16 11 11 11 2 11 1 11 1 9 12 9 13 12 12 9 13 2
11 9 1 11 1 9 1 12 9 9 13 2
26 11 11 11 1 12 9 0 9 1 9 1 0 9 1 11 11 11 2 11 2 1 0 13 13 4 2
20 11 11 1 9 13 16 11 1 9 11 11 11 1 0 13 1 1 13 4 2
19 7 11 1 0 9 1 1 11 11 1 1 9 1 9 0 13 4 4 2
16 9 1 11 9 1 9 1 9 1 9 1 1 10 9 13 2
32 9 1 9 13 16 11 9 1 9 1 9 0 9 1 13 4 2 15 0 9 9 1 9 13 4 4 7 11 1 0 13 2
21 15 1 9 1 9 13 16 11 9 1 9 1 11 9 1 9 1 9 10 13 2
29 10 9 11 9 1 9 1 9 9 1 9 1 1 7 3 1 13 9 1 1 15 9 1 3 10 14 9 13 2
31 11 11 11 11 11 11 1 11 1 0 11 11 11 11 1 0 9 13 4 11 1 1 0 9 1 10 9 1 9 13 2
28 10 3 11 1 10 9 9 1 9 13 15 13 4 4 16 0 9 9 11 11 1 11 1 0 9 13 4 2
51 11 11 1 11 11 1 9 11 11 1 11 1 9 1 13 16 11 11 9 9 11 0 13 15 15 11 7 11 1 0 9 1 9 1 9 1 1 2 9 9 9 1 0 7 0 9 1 14 9 13 2
16 10 9 1 9 9 0 11 11 11 1 11 11 1 9 13 2
21 11 11 1 11 11 1 11 1 0 11 11 11 1 0 9 1 11 1 9 13 2
7 15 1 11 11 11 13 2
6 11 1 15 11 13 2
12 15 15 9 0 11 11 11 11 1 13 4 2
34 11 9 2 11 11 2 1 9 13 4 16 11 0 9 11 11 1 1 11 11 13 7 15 11 1 9 13 11 11 1 9 13 4 2
47 15 1 0 11 11 11 11 1 11 1 0 9 11 11 1 9 1 1 11 1 13 16 11 1 11 1 13 1 9 9 1 11 1 13 4 9 1 9 1 9 13 1 15 10 9 13 2
26 11 1 11 1 11 11 11 1 11 2 11 9 9 1 15 12 9 1 13 1 1 9 13 4 4 2
27 11 1 9 9 15 9 13 4 13 16 11 11 1 9 13 1 1 11 1 9 1 1 1 9 13 4 2
12 7 15 15 1 1 15 9 14 13 4 4 2
19 11 1 11 1 9 13 1 10 9 1 15 12 9 13 1 9 13 4 2
9 11 11 11 11 1 9 14 13 2
29 11 1 11 1 11 11 11 11 11 1 9 1 9 1 13 16 11 1 13 4 9 11 0 0 9 1 1 13 2
23 11 1 13 16 15 11 1 0 13 4 16 15 15 11 13 7 10 9 1 13 9 13 2
14 10 9 1 11 7 11 9 15 15 1 9 1 13 2
24 15 13 16 16 11 1 11 10 9 1 15 12 9 13 11 13 13 4 16 15 15 9 13 2
21 16 11 11 1 9 1 13 4 16 15 9 13 11 13 1 11 1 0 11 13 2
22 15 1 11 1 11 1 0 11 11 11 11 12 9 1 1 12 9 13 11 13 4 2
23 11 9 1 11 9 1 1 13 4 9 9 13 1 9 3 0 13 9 1 13 4 4 2
29 9 1 9 11 11 1 9 11 1 12 9 11 7 11 11 1 0 2 8 13 4 9 2 9 9 13 4 4 2
29 0 13 16 11 9 1 9 7 11 11 1 9 11 11 11 1 11 9 1 9 13 9 13 1 10 9 13 4 2
32 11 1 9 1 1 11 9 1 12 2 8 9 13 1 1 9 11 7 11 7 15 9 1 14 0 2 8 9 13 4 4 2
18 15 13 4 4 4 16 11 1 11 9 1 9 12 12 9 13 4 2
29 9 1 1 15 9 1 11 1 13 4 16 9 1 0 9 1 9 13 1 3 15 9 1 14 9 13 4 4 2
32 13 4 4 4 16 11 1 9 13 4 16 12 9 1 9 1 0 9 11 11 11 2 11 2 7 11 11 11 13 4 4 2
14 7 9 1 9 1 11 11 7 9 1 0 9 13 2
33 15 1 11 1 9 13 11 9 1 1 15 0 9 13 7 15 1 15 0 14 13 16 11 7 11 1 1 15 11 1 0 13 2
17 10 9 1 1 12 9 1 1 15 14 15 13 1 0 14 13 2
18 11 1 9 1 1 11 9 1 1 1 15 14 9 3 14 13 4 2
40 15 1 9 1 9 1 9 13 2 9 1 1 11 1 11 7 11 11 1 9 1 9 1 12 2 8 9 7 0 12 9 9 11 1 13 1 9 13 4 2
25 11 1 13 4 0 9 1 1 12 9 1 9 1 9 1 9 1 9 1 10 2 8 9 13 2
15 15 9 1 0 9 1 12 0 9 1 1 9 0 13 2
25 11 1 13 4 9 1 9 1 1 10 9 1 9 1 11 13 15 9 1 0 9 13 4 4 2
19 11 9 1 9 1 9 1 9 1 9 1 1 9 1 0 9 13 4 2
18 15 11 7 11 1 15 2 8 9 1 9 1 0 9 0 13 4 2
7 15 1 11 1 9 13 2
12 9 1 11 11 1 9 12 12 9 13 4 2
16 0 9 9 1 12 9 1 11 1 9 12 12 9 13 4 2
14 10 9 9 1 3 0 9 9 7 9 0 13 4 2
30 7 11 1 15 0 9 0 13 1 1 15 12 12 9 1 9 13 7 15 1 14 10 9 9 1 9 13 9 13 2
27 11 11 1 11 11 11 1 13 9 1 0 13 4 11 11 11 11 11 9 13 1 0 9 13 4 4 2
33 11 11 11 11 11 1 11 11 1 11 9 1 10 9 1 9 13 13 4 4 7 10 9 1 13 15 1 9 0 13 4 4 2
22 12 9 14 15 1 13 13 16 10 9 1 9 11 11 1 14 15 13 4 4 4 2
12 10 10 9 13 15 11 11 1 10 0 13 2
17 0 9 10 9 1 13 14 13 15 10 9 1 0 13 4 4 2
28 10 0 9 1 9 1 9 15 13 16 0 13 1 1 15 1 10 9 1 10 9 1 0 14 13 4 4 2
17 15 11 11 14 0 13 15 1 14 12 9 10 9 1 0 13 2
22 15 14 15 0 13 4 4 16 11 11 11 1 11 11 1 14 10 9 1 9 13 2
25 11 11 11 1 9 1 1 11 9 1 11 11 1 9 1 9 13 4 15 1 9 14 0 13 2
11 3 10 9 1 9 11 1 13 4 4 2
17 15 9 13 4 15 11 11 1 10 9 1 9 13 4 4 4 2
17 0 9 1 9 1 13 10 9 1 0 9 1 13 4 4 4 2
14 16 9 15 1 1 15 1 1 9 13 1 13 4 2
38 9 1 9 1 13 13 16 16 11 1 9 13 1 9 13 16 11 1 12 9 1 1 11 11 1 12 9 1 14 10 9 1 15 0 13 4 4 2
12 9 9 1 9 1 13 14 0 13 4 4 2
14 11 11 1 10 9 1 12 9 1 0 13 4 4 2
33 10 9 13 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
27 9 1 1 9 1 9 1 1 11 11 1 9 2 9 9 2 1 9 1 9 9 1 9 13 4 4 2
11 15 1 11 11 11 1 14 9 13 4 2
31 11 11 1 11 1 9 1 9 1 1 9 2 9 13 9 1 9 1 9 13 7 11 1 10 9 0 9 13 4 4 2
13 11 11 1 0 11 11 9 1 9 1 0 13 2
21 9 1 9 1 9 11 11 1 11 11 1 11 1 1 9 13 1 9 13 4 2
16 15 13 13 2 2 11 11 1 9 1 9 3 0 13 4 4
34 9 1 9 1 15 9 9 13 4 16 15 1 3 10 9 11 11 1 0 9 1 14 13 4 7 9 3 11 1 9 13 4 4 2
22 11 7 11 1 11 1 0 9 9 13 7 11 11 1 9 1 9 13 4 4 4 2
26 11 11 7 0 11 11 1 1 3 15 15 9 1 9 1 9 13 1 1 0 9 1 9 14 13 2
17 11 10 9 1 0 9 1 9 1 0 13 1 9 13 4 4 2
36 11 11 11 11 2 11 2 1 9 11 11 11 1 1 12 9 1 1 11 11 11 11 2 11 2 9 1 11 2 11 11 0 13 4 4 2
11 16 9 9 13 1 3 15 9 14 13 2
18 11 1 1 11 0 0 9 9 1 1 1 15 9 14 13 4 4 2
23 11 11 1 15 11 11 11 11 9 13 1 3 9 1 11 1 0 9 1 13 4 4 2
21 11 1 1 9 9 1 1 9 9 1 9 7 15 9 1 0 0 9 13 4 2
8 7 15 0 9 14 13 4 2
15 15 13 16 11 11 2 11 12 9 1 1 0 13 4 2
12 15 9 9 1 15 1 13 4 1 0 13 2
32 11 1 13 16 0 9 12 9 2 9 2 9 1 9 13 4 15 9 9 1 0 13 1 0 9 1 9 13 1 9 13 2
30 15 13 16 15 0 9 9 11 7 11 7 0 11 11 2 11 1 11 0 9 9 1 9 1 0 9 0 13 4 2
19 11 1 13 16 0 2 11 11 11 2 11 1 1 9 1 9 0 13 2
12 10 9 1 9 1 9 1 9 1 9 13 2
24 3 10 9 1 1 11 10 9 1 14 9 13 4 4 16 9 1 9 1 0 13 4 4 2
14 11 11 11 11 1 11 1 12 0 9 1 0 13 2
11 0 12 9 1 15 10 0 9 9 13 2
17 10 3 11 0 0 9 1 11 11 11 1 15 9 1 3 13 2
24 15 11 2 11 11 1 14 9 13 2 15 0 9 1 0 9 1 0 9 13 1 9 13 2
26 9 1 1 11 11 1 11 2 11 7 11 11 1 9 1 1 0 0 9 1 9 13 1 9 13 2
23 0 2 0 11 1 12 9 1 9 11 11 7 11 1 0 0 9 1 9 13 4 4 2
24 11 11 1 13 1 11 2 11 7 3 11 11 1 13 1 11 11 11 1 11 1 9 13 2
28 11 11 11 1 11 1 10 12 9 9 7 11 1 1 11 2 11 2 11 11 2 11 7 11 14 0 13 2
15 10 9 1 9 1 0 9 1 13 1 9 14 0 13 2
24 11 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 0 13 2
21 2 11 11 11 2 1 9 1 1 0 0 9 1 0 13 1 9 13 4 4 2
16 0 9 11 1 0 2 0 9 1 9 1 9 13 4 4 2
13 11 1 11 1 14 10 9 9 1 0 13 4 2
12 3 1 11 7 11 1 14 15 0 13 4 2
26 11 1 9 1 13 1 0 11 2 11 11 1 12 9 12 0 9 9 1 9 0 13 1 9 13 2
17 0 12 9 1 11 2 11 9 1 0 12 9 1 9 13 4 2
19 11 1 0 9 1 13 4 11 1 1 1 9 9 14 13 4 4 4 2
43 11 11 11 11 11 1 11 1 9 1 12 0 9 1 13 16 11 1 11 9 1 9 7 9 0 13 1 3 15 1 9 1 13 4 9 9 1 3 9 13 4 4 2
25 11 1 13 16 11 11 1 0 9 1 9 7 0 9 1 1 10 0 9 13 1 1 0 13 2
37 12 0 9 1 9 1 11 0 0 9 1 1 1 0 9 1 9 13 4 15 13 16 11 1 14 12 0 0 9 0 13 2 15 12 9 13 2
30 11 11 11 11 11 11 1 13 16 11 1 0 9 1 9 9 9 9 1 0 13 1 1 15 0 9 14 13 4 2
45 9 9 1 10 9 9 13 4 1 9 1 1 1 15 13 16 9 9 1 13 4 9 1 9 13 1 9 1 0 9 0 13 2 7 10 9 9 13 4 1 15 9 14 13 2
29 15 13 16 11 14 9 1 9 1 1 9 9 1 0 9 0 13 1 1 11 11 1 10 9 9 13 4 4 2
26 11 1 13 13 16 9 9 1 9 1 9 7 15 9 1 0 9 7 9 1 3 9 13 4 4 2
41 11 11 11 1 13 16 11 11 1 11 7 11 1 1 0 9 1 9 1 1 9 9 0 13 1 9 1 11 7 11 1 9 9 9 1 12 9 13 4 4 2
32 11 7 11 11 1 1 11 1 9 9 1 9 1 1 11 1 0 11 11 1 9 1 1 11 1 12 9 1 9 13 4 2
24 9 1 10 9 1 9 1 0 9 1 9 7 0 9 1 9 1 9 13 1 1 13 4 2
34 9 9 1 9 1 1 11 1 0 13 4 12 9 1 9 13 4 9 9 11 11 11 7 9 11 11 11 1 11 1 10 9 13 2
30 9 9 11 11 11 1 9 1 13 16 9 1 9 1 1 1 15 9 1 9 13 4 7 10 9 1 9 13 4 2
26 9 1 13 16 9 1 10 9 1 9 3 1 0 13 7 9 1 9 1 10 9 1 0 13 13 2
29 9 1 1 1 11 1 9 13 4 0 9 11 11 11 1 13 16 0 0 9 1 9 9 1 14 13 4 4 2
31 15 13 16 9 1 0 7 9 1 0 9 7 0 9 1 0 9 1 9 1 13 11 11 1 15 9 1 0 13 4 2
36 15 15 14 9 13 16 0 9 1 11 11 11 11 7 10 9 9 1 0 13 4 4 2 16 10 9 1 0 9 1 1 1 0 9 13 2
34 9 1 1 1 11 7 11 11 1 9 13 1 9 1 11 11 1 12 9 1 9 13 2 15 1 10 9 1 10 9 13 4 4 2
12 15 13 16 10 9 1 0 9 13 4 4 2
37 11 11 1 11 11 7 11 1 11 7 11 11 1 1 12 0 9 0 13 10 9 1 15 12 9 9 9 15 9 1 13 4 1 9 13 4 2
22 9 13 4 13 4 0 9 1 12 9 0 13 4 7 12 9 0 9 1 0 13 2
21 11 9 1 10 9 11 1 10 9 13 15 11 11 1 12 9 9 13 4 4 2
28 0 9 1 13 16 11 11 1 9 9 11 9 1 11 11 11 11 1 13 4 4 2 10 9 0 9 13 2
12 9 13 14 9 1 3 9 13 9 13 4 2
10 9 1 12 9 9 1 14 13 4 2
8 0 9 1 14 9 13 4 2
18 15 1 15 0 14 13 16 10 9 1 10 9 13 4 7 0 13 2
23 0 13 16 11 9 15 12 9 1 0 9 1 9 13 4 1 3 9 10 13 4 4 2
21 10 9 1 13 4 0 9 1 9 11 1 9 14 11 1 9 1 9 13 4 2
26 11 1 9 9 9 11 11 11 1 13 16 11 1 9 9 11 9 1 10 9 1 9 1 9 13 2
15 7 9 1 15 0 9 1 9 1 15 9 14 13 4 2
41 10 9 1 1 0 9 1 13 4 9 7 9 1 9 1 0 13 4 4 4 7 15 9 1 12 9 2 11 2 11 2 11 7 11 1 3 9 13 4 4 2
23 10 9 1 11 1 11 9 1 9 13 4 10 14 10 12 0 9 1 9 13 4 4 2
20 9 9 1 13 16 15 9 15 14 0 9 1 9 13 1 1 9 1 13 2
19 11 11 11 11 2 11 2 1 11 11 1 11 1 0 9 13 4 4 2
18 15 0 9 7 9 13 1 9 1 9 1 13 1 9 13 4 4 2
20 0 13 16 11 9 7 15 1 11 11 10 9 1 9 1 9 13 4 4 2
13 3 11 2 11 11 11 1 9 9 1 0 13 2
20 11 11 2 11 2 1 0 9 11 11 1 12 9 1 9 9 1 13 4 2
13 9 1 10 9 9 11 15 9 1 13 4 4 2
18 11 1 11 1 9 0 13 1 1 0 9 1 9 1 0 13 4 2
17 11 1 11 1 0 9 1 9 1 0 9 1 9 9 13 4 2
19 9 9 1 1 9 0 13 1 1 15 11 1 0 2 8 9 13 4 2
34 15 13 16 15 9 13 16 11 11 1 11 11 1 15 15 9 9 13 15 15 9 9 1 10 9 11 1 13 1 0 13 4 4 2
8 9 10 9 9 13 4 4 2
13 15 9 1 9 9 9 7 9 9 13 4 4 2
15 15 13 16 11 1 9 1 1 9 1 9 9 13 4 2
18 15 0 9 1 0 13 1 1 9 1 9 13 1 1 0 13 4 2
15 11 1 9 13 1 1 15 9 9 1 3 9 13 4 2
27 9 9 1 9 13 4 15 13 16 9 1 9 1 15 9 1 3 13 7 9 11 11 1 0 9 13 2
14 9 10 9 0 9 9 1 0 13 1 13 4 4 2
53 11 1 11 11 11 11 1 0 13 1 9 1 13 4 0 9 9 1 0 11 11 11 11 1 11 1 13 4 16 11 11 1 9 1 11 9 13 1 1 11 3 2 11 9 2 1 1 1 9 13 4 4 2
32 11 9 9 1 9 11 11 1 1 15 9 9 1 15 9 1 13 16 11 1 0 11 0 13 1 1 11 1 9 13 4 2
15 11 9 1 0 9 1 9 1 1 11 1 11 11 13 2
37 15 9 9 1 1 15 11 11 1 9 1 9 1 1 0 9 1 9 1 0 9 9 9 1 9 1 11 11 1 9 1 9 1 0 9 13 2
27 11 11 11 11 2 11 2 1 0 9 11 11 1 9 1 10 9 1 9 13 1 9 13 4 4 4 2
7 10 9 11 1 13 4 2
13 11 1 11 11 11 9 1 9 13 1 9 13 2
21 11 9 1 1 9 1 0 9 1 15 1 1 15 9 13 4 1 9 0 13 2
28 0 9 1 9 13 1 1 9 2 9 1 9 13 1 3 11 11 11 11 1 9 7 9 1 9 13 4 2
12 9 1 0 9 1 11 11 1 0 9 13 2
22 11 1 9 9 1 13 16 9 11 1 12 9 9 9 9 1 0 13 13 4 4 2
22 15 1 9 7 9 1 9 1 13 10 0 9 13 2 15 9 3 10 13 4 4 2
23 11 1 13 16 9 1 9 9 1 0 13 1 3 15 9 1 0 9 1 13 4 4 2
15 15 13 2 2 10 9 1 15 9 1 9 7 9 13 2
18 10 9 8 0 13 7 15 15 1 3 7 9 1 1 9 13 13 4
31 11 10 9 1 0 9 0 13 16 9 7 9 1 0 9 9 1 0 13 7 15 9 1 9 1 13 10 0 14 13 2
17 7 11 7 11 11 11 10 15 14 9 1 0 9 13 4 4 2
26 0 13 16 11 11 11 11 1 1 11 11 1 9 1 0 9 10 13 9 1 9 1 13 4 4 2
5 9 1 9 13 2
27 15 1 0 2 0 9 1 9 1 9 1 13 7 9 9 0 9 1 9 13 1 1 15 9 14 13 2
31 11 1 13 16 10 10 9 9 7 9 1 1 0 9 1 0 13 7 10 9 1 10 9 1 0 9 3 13 4 4 2
20 15 1 1 10 9 1 11 11 1 11 11 11 1 1 9 9 13 4 4 2
18 7 10 9 9 3 13 7 0 9 1 0 13 1 9 13 4 4 2
22 12 9 1 1 11 1 10 12 12 9 13 2 15 10 13 12 12 12 9 0 13 2
8 10 9 9 9 1 0 13 2
12 15 1 11 1 9 10 9 1 13 0 13 2
19 11 1 13 4 16 9 2 9 1 13 4 1 9 1 9 14 13 4 2
13 15 13 16 9 9 1 9 13 4 1 9 13 2
23 16 11 11 1 10 9 13 4 4 16 15 9 0 13 7 15 14 15 9 13 4 4 2
14 15 13 16 9 7 9 1 9 9 13 4 4 4 2
23 15 9 2 9 7 9 1 9 1 9 13 1 0 9 1 9 1 9 3 13 4 4 2
11 9 1 1 9 1 10 9 1 9 13 2
34 9 1 11 11 1 11 11 11 11 1 9 1 0 9 1 0 9 1 9 1 12 9 1 13 16 9 1 1 9 1 15 12 13 2
25 10 9 1 9 1 10 9 1 0 9 1 13 4 0 9 1 12 9 1 9 13 9 13 4 2
22 9 7 9 1 9 1 9 13 4 0 13 0 9 1 9 7 9 1 0 13 4 2
46 10 9 1 11 1 13 11 1 0 9 1 9 13 1 11 1 9 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 1 9 13 0 13 4 2
21 12 9 11 11 2 11 11 11 7 11 11 1 14 15 9 1 1 0 13 4 2
21 15 9 13 4 4 16 9 1 1 12 0 9 0 13 2 15 10 9 9 13 2
29 11 1 10 9 1 1 10 9 1 0 9 13 1 9 13 15 9 1 9 13 4 7 0 9 1 9 13 4 2
18 11 11 1 9 11 11 1 13 16 9 9 1 9 1 0 9 13 2
18 9 9 15 13 1 13 16 9 1 9 1 0 9 1 15 13 4 2
11 10 9 1 0 9 11 11 0 9 13 2
14 9 1 11 1 0 9 11 11 11 11 14 0 13 2
19 11 1 9 13 13 11 11 1 0 9 11 11 1 9 1 0 13 4 2
14 11 11 1 11 11 11 11 11 1 1 0 13 4 2
12 11 1 9 1 10 9 9 0 13 4 4 2
13 10 9 15 11 1 0 12 0 9 1 13 4 2
14 16 2 15 11 1 10 9 1 9 9 0 14 13 2
31 9 1 9 13 1 1 11 1 9 1 9 9 1 13 4 2 7 15 15 14 13 7 11 11 1 9 1 0 13 4 2
20 11 11 1 9 1 9 13 1 3 11 11 11 0 11 1 9 14 13 4 2
9 15 15 9 10 11 9 1 13 2
13 11 9 9 11 11 11 1 13 1 9 1 13 2
21 10 9 9 9 1 9 1 1 15 3 13 4 7 9 9 1 1 0 13 4 2
14 11 11 11 1 1 13 1 9 9 1 15 13 4 2
9 9 1 1 11 11 1 9 13 2
16 9 1 1 2 11 11 11 11 11 1 11 9 1 9 13 2
20 11 1 15 11 2 11 9 1 12 9 1 0 9 7 12 9 13 4 4 2
15 15 1 15 9 1 9 1 12 9 1 12 12 9 13 2
13 10 3 15 9 11 1 11 9 11 11 1 13 2
21 11 1 11 11 1 10 0 0 9 1 1 9 1 9 13 1 1 11 13 4 2
25 15 11 11 1 1 2 11 11 2 9 1 15 7 0 9 1 12 9 1 9 1 9 13 4 2
27 11 1 9 13 1 3 15 12 9 1 11 2 11 1 9 13 4 2 7 11 1 15 0 13 4 4 2
20 10 9 1 9 1 13 1 3 11 9 1 15 12 12 9 13 11 13 4 2
15 11 11 10 9 11 1 11 7 11 1 0 9 1 13 2
11 10 9 1 15 11 1 11 1 13 4 2
21 9 11 1 10 9 1 9 1 13 4 2 15 15 9 13 1 1 11 13 4 2
10 9 1 1 11 1 9 3 0 13 2
12 15 9 1 0 9 13 1 9 3 13 4 2
13 9 1 1 9 1 9 13 2 15 0 9 13 2
12 11 1 9 1 0 12 9 1 9 13 4 2
33 0 9 1 9 9 1 9 13 2 15 15 1 0 9 12 9 3 13 4 12 9 9 1 13 4 2 7 0 9 12 9 13 2
15 3 11 1 9 1 1 9 13 2 15 10 9 13 4 2
12 11 2 11 11 11 9 0 9 14 0 13 2
10 14 12 12 9 9 1 13 4 4 2
11 15 0 9 9 1 9 1 13 4 4 2
19 15 9 1 13 14 12 12 9 1 9 1 3 1 9 1 9 13 4 2
18 11 11 1 14 11 2 11 7 11 9 1 0 9 1 13 4 4 2
20 9 1 10 9 1 9 1 9 1 9 1 15 1 9 1 10 9 13 4 2
16 11 2 11 7 11 2 11 9 1 0 9 1 13 4 4 2
13 11 2 11 7 11 1 9 0 9 12 9 13 2
16 11 1 11 1 0 12 9 1 9 13 1 9 13 4 4 2
16 9 1 0 9 9 1 12 9 0 9 1 0 13 4 4 2
16 11 1 1 11 9 7 11 9 1 3 10 12 9 9 13 2
21 0 12 9 1 15 0 9 1 1 1 0 9 12 1 12 9 3 13 4 4 2
16 9 9 1 15 0 12 9 1 9 2 9 1 9 13 4 2
10 11 1 9 3 10 12 9 9 13 2
36 11 11 1 11 1 0 11 11 11 1 9 1 0 9 11 11 1 9 13 1 9 1 9 1 9 13 1 1 12 0 9 1 9 13 4 2
15 9 1 13 16 0 9 12 9 1 1 15 9 9 13 2
13 9 1 13 16 0 9 1 13 4 9 0 13 2
14 9 1 9 9 1 9 1 9 13 1 9 13 4 2
26 9 1 15 14 13 16 15 9 13 4 16 11 9 1 0 13 4 4 7 11 15 9 13 4 4 2
40 10 9 1 9 13 4 9 11 11 7 9 11 11 11 1 9 1 13 16 9 9 11 9 1 9 9 9 1 15 14 9 1 10 9 1 9 13 4 4 2
25 9 1 13 16 15 9 13 10 0 13 16 15 9 13 4 4 7 10 0 9 1 9 15 13 2
34 0 13 16 9 14 1 11 11 1 9 1 12 9 0 13 13 4 16 15 15 0 9 13 7 15 1 0 9 1 15 9 14 13 2
16 11 11 1 1 1 13 4 16 9 11 1 0 13 4 4 2
30 0 13 16 11 11 1 11 11 1 9 13 4 16 15 1 9 13 9 13 4 4 7 11 1 9 1 9 13 4 2
21 7 9 1 12 12 2 12 12 9 2 1 9 13 9 15 9 1 0 13 4 2
26 9 2 9 1 1 9 9 1 13 4 9 1 12 9 1 9 1 13 10 0 9 1 15 9 13 2
8 9 11 11 1 12 9 13 2
21 7 9 1 9 2 11 1 9 2 11 11 2 12 0 2 1 3 14 13 4 2
15 11 11 12 9 1 12 13 9 1 12 9 1 13 4 2
30 0 9 1 9 12 0 9 9 1 9 13 4 9 1 13 0 9 1 12 9 1 9 13 12 0 9 1 9 13 2
16 12 9 1 0 10 9 11 1 11 11 9 1 13 4 4 2
17 9 9 1 13 16 15 1 0 9 9 2 11 2 1 15 13 2
19 15 13 16 10 0 9 1 12 9 1 13 11 11 1 12 9 13 4 2
19 15 1 12 9 1 9 1 1 13 4 7 15 12 9 1 0 13 13 2
22 9 1 13 1 3 15 0 9 1 9 13 2 15 11 11 11 9 1 0 13 4 2
10 9 1 13 9 1 9 1 15 13 2
13 11 11 13 4 15 9 7 9 13 4 4 4 2
27 11 11 11 1 13 13 9 1 1 11 9 11 11 3 11 11 11 2 11 2 1 9 9 14 13 13 2
14 15 15 10 9 9 1 0 9 1 14 13 4 4 2
24 9 9 1 10 9 1 1 14 9 1 11 1 9 1 9 1 0 14 13 1 9 13 4 2
22 9 1 1 10 9 14 9 1 13 4 4 16 10 9 1 15 9 1 14 13 4 2
25 11 11 11 1 9 1 11 9 11 11 1 9 9 0 13 1 3 11 11 9 1 9 1 13 2
26 11 1 12 9 3 9 1 9 13 7 11 11 1 11 1 9 9 7 9 1 9 1 9 13 4 2
7 7 9 15 1 0 13 2
15 9 1 9 13 16 11 11 11 11 1 9 1 13 4 2
15 15 9 1 13 1 1 11 11 1 15 9 1 9 13 2
17 11 11 11 1 9 1 11 3 9 1 9 13 1 9 1 13 2
18 9 0 9 1 9 0 13 1 9 1 9 1 11 1 0 14 13 2
14 16 2 9 11 11 1 12 9 3 9 14 13 4 2
24 9 1 0 9 1 1 2 11 1 9 9 1 9 1 1 11 9 3 10 9 1 14 13 2
13 7 9 1 10 9 15 10 9 1 0 14 13 2
22 9 9 1 9 13 16 11 11 1 11 1 9 14 13 1 9 1 9 10 13 4 2
11 9 1 10 9 11 3 0 9 9 13 2
8 15 2 15 10 9 13 4 2
12 7 11 11 15 1 9 1 3 13 13 4 2
15 15 2 15 11 1 9 9 3 14 13 1 9 13 4 2
15 11 1 0 9 7 9 1 9 11 11 11 1 11 13 2
12 15 15 1 13 12 12 9 1 9 1 9 2
22 10 9 15 15 11 11 11 11 11 1 9 13 1 3 11 11 1 0 9 1 13 2
24 15 9 1 9 1 2 11 11 2 1 9 1 9 13 4 13 16 10 15 14 9 14 13 2
21 15 1 14 15 0 0 9 1 15 10 9 1 9 13 7 9 1 9 9 13 2
18 10 3 15 9 9 1 9 1 1 12 12 9 13 1 14 9 13 2
19 0 9 1 13 9 7 9 1 1 9 9 1 10 9 3 14 9 13 2
20 15 13 16 11 11 11 2 11 7 11 1 9 9 1 1 1 0 13 4 2
14 11 11 11 11 11 1 9 9 1 0 9 13 13 2
35 15 9 13 16 11 11 11 7 11 11 11 7 11 11 11 11 1 1 1 12 9 1 1 11 1 0 10 9 1 12 12 9 9 13 2
9 12 12 9 1 9 1 9 13 2
13 9 1 11 11 11 11 1 9 1 0 9 13 2
48 11 9 9 1 11 11 11 11 11 11 1 9 13 1 3 15 0 9 1 11 1 13 16 10 9 15 1 14 11 1 9 1 14 13 4 7 15 11 1 9 14 10 9 1 9 13 4 2
35 9 1 9 7 9 1 0 9 13 4 15 13 16 3 14 11 11 2 11 1 1 1 9 1 0 9 13 1 1 11 1 9 13 4 2
26 9 1 9 1 13 9 1 9 13 4 15 13 16 10 9 1 9 13 1 1 15 1 9 13 4 2
21 9 1 0 9 11 11 11 1 9 9 1 1 12 12 1 9 11 1 9 13 2
23 15 1 11 11 11 1 11 7 11 1 11 11 13 2 15 15 9 1 1 9 9 13 2
7 15 1 11 9 9 13 2
27 11 1 0 9 11 11 11 1 11 11 11 2 11 2 1 0 0 13 4 15 9 13 1 9 13 4 2
19 15 13 16 11 11 1 9 1 1 11 1 12 2 11 2 1 9 13 2
7 11 1 15 9 14 13 2
17 11 1 11 1 9 9 1 9 1 9 1 11 1 0 9 13 2
12 0 13 16 11 9 11 11 11 1 9 13 2
22 7 11 11 11 0 9 1 15 10 9 1 1 9 1 9 1 14 9 13 4 4 2
27 11 1 9 1 11 9 1 9 1 13 1 3 11 11 11 1 9 13 1 1 11 1 9 13 4 4 2
24 0 9 11 11 11 1 1 11 1 0 9 11 11 1 14 11 1 0 13 1 9 13 4 2
38 11 9 9 11 11 11 11 11 2 11 2 1 0 11 11 1 0 9 9 1 9 13 1 12 9 1 11 1 10 9 1 9 13 1 9 13 4 2
27 15 13 13 16 11 7 11 9 1 16 9 13 15 9 14 13 16 9 9 1 9 1 15 0 13 4 2
29 11 1 9 11 1 9 11 11 1 0 9 1 13 9 2 9 1 1 11 7 11 1 15 9 1 9 13 4 2
16 15 14 13 1 15 15 9 9 1 9 1 3 14 9 13 2
15 15 1 0 9 1 15 1 0 10 9 1 13 1 13 2
46 12 0 0 9 1 9 13 4 11 11 11 1 0 9 7 15 11 11 11 1 9 11 11 1 13 16 11 1 11 7 9 1 1 9 9 1 0 13 4 16 15 12 0 9 13 2
20 11 1 9 1 9 13 4 11 1 13 16 9 1 15 1 0 9 13 4 2
32 0 13 16 11 11 1 11 9 1 12 9 1 9 1 9 13 11 13 1 3 0 11 1 11 1 1 9 1 9 13 4 2
15 11 11 11 11 11 1 9 11 1 9 9 1 9 13 2
22 3 11 1 12 9 1 13 16 9 1 1 9 9 14 15 9 1 9 13 4 4 2
13 11 7 9 9 1 10 9 1 0 9 13 4 2
30 11 11 1 0 11 11 11 1 9 1 11 1 3 14 9 13 2 3 15 9 1 14 9 1 9 13 9 13 4 2
30 9 1 11 11 1 9 1 0 9 13 1 11 11 1 0 13 1 15 0 9 1 1 14 15 15 9 13 14 14 2
17 11 11 11 1 9 1 1 14 15 15 1 1 3 0 11 13 2
41 11 1 2 11 11 2 1 13 16 11 11 1 9 2 15 12 12 9 0 13 2 1 1 16 9 1 0 9 1 9 13 4 16 15 9 9 1 0 9 13 2
19 9 11 11 1 11 11 2 11 11 0 9 1 12 9 9 14 13 4 2
19 10 9 1 1 11 11 1 9 1 9 13 1 9 1 3 9 13 4 2
39 9 14 1 11 1 9 11 11 1 9 1 0 13 7 11 11 1 0 9 1 13 4 1 11 9 1 1 13 1 9 15 0 9 1 14 14 13 4 2
17 11 11 11 1 15 0 0 9 1 9 10 9 1 10 14 13 2
32 11 11 2 11 11 11 2 11 11 11 7 11 11 1 10 9 1 1 0 11 11 1 15 1 13 9 1 9 1 9 13 2
25 11 11 11 11 11 11 1 10 0 9 9 1 11 11 11 1 9 1 0 13 1 9 13 4 2
20 15 13 16 0 9 1 13 4 9 7 9 1 9 1 0 14 13 4 4 2
19 11 11 1 9 9 9 9 7 0 9 9 1 9 1 0 13 4 4 2
35 12 0 9 1 11 1 13 16 10 9 7 0 9 1 15 0 13 4 16 11 11 11 11 11 1 1 9 1 9 1 1 9 13 4 2
24 16 15 14 13 4 4 16 10 9 1 1 9 13 4 15 10 9 1 9 14 13 4 4 2
22 15 13 16 10 9 1 1 9 1 9 13 4 16 9 9 1 0 9 1 0 13 2
20 11 1 13 16 9 1 0 9 13 4 4 7 15 1 0 13 1 9 13 2
29 0 9 1 9 1 9 1 9 13 4 13 16 15 9 1 3 9 14 13 7 11 1 9 0 9 1 1 13 2
27 10 9 1 9 1 9 1 9 9 11 11 11 1 9 11 11 11 11 1 9 1 0 9 1 9 13 2
17 15 13 9 10 9 1 9 1 9 13 9 1 9 13 13 4 2
11 7 15 15 9 1 0 14 13 4 4 2
27 11 9 11 11 11 1 11 11 1 13 0 9 1 9 13 4 9 1 9 9 13 4 1 9 13 4 2
16 15 13 11 9 15 14 9 1 0 9 1 9 14 13 4 2
13 15 13 13 10 9 9 9 1 0 9 13 4 2
34 9 9 1 13 13 16 11 1 9 1 0 9 1 9 7 0 9 1 9 1 13 4 15 9 1 9 7 9 1 15 9 14 13 2
40 9 1 9 9 11 11 11 1 9 11 11 11 7 11 1 9 9 11 11 11 1 0 9 11 11 1 11 1 13 16 11 9 1 9 1 1 0 14 13 2
20 7 11 1 11 1 9 1 13 4 9 1 9 7 15 9 1 9 14 13 2
27 10 9 1 0 9 7 0 9 1 9 1 9 7 9 9 1 9 1 9 13 9 1 1 9 13 4 2
31 11 11 1 13 16 15 1 11 1 11 1 9 13 4 2 15 1 9 14 1 14 12 12 1 10 9 9 13 4 4 2
15 15 13 16 0 9 9 9 1 9 13 1 9 1 13 2
18 11 1 9 1 11 11 11 7 0 0 9 1 9 1 9 13 4 2
12 11 1 11 1 9 1 9 13 1 9 13 2
21 15 11 1 9 13 16 15 11 9 1 9 1 9 13 1 1 9 13 4 4 2
13 11 1 11 9 9 1 9 1 3 0 9 13 2
17 15 1 11 14 10 9 1 1 9 1 0 9 13 4 4 4 2
18 12 0 9 1 1 11 1 12 9 1 10 9 11 9 1 13 4 2
41 15 1 12 1 10 0 9 11 1 11 2 11 9 1 9 9 1 1 9 1 13 4 4 7 12 1 10 9 11 1 11 1 9 1 9 9 1 9 13 4 2
20 15 1 11 2 11 2 11 0 0 9 1 12 1 1 12 9 11 1 13 2
16 11 1 12 0 9 9 10 9 1 9 1 9 13 4 4 2
8 15 1 12 11 11 1 13 2
25 9 1 1 11 1 14 11 2 11 2 11 1 0 9 1 12 1 10 0 9 9 13 4 4 2
13 9 7 0 9 10 9 1 9 1 1 13 4 2
18 3 11 1 11 9 14 9 1 9 1 12 0 9 13 4 4 4 2
21 15 9 1 9 1 11 1 12 1 10 9 11 1 9 9 1 9 13 4 4 2
38 15 12 11 2 11 2 11 2 12 11 11 11 2 12 11 11 2 12 11 2 12 11 2 11 7 12 11 2 11 2 11 0 0 9 1 9 13 2
31 9 1 0 0 9 13 4 1 9 1 0 9 13 4 11 7 11 2 11 1 12 9 9 1 9 13 1 9 13 4 2
42 11 1 11 11 11 11 1 0 9 1 13 16 9 1 13 10 9 1 13 0 2 0 9 1 1 9 13 4 16 10 9 1 9 1 9 1 9 1 9 13 4 2
22 11 7 11 2 11 1 1 11 2 11 2 11 7 11 1 14 0 9 13 4 4 2
42 9 1 9 1 9 13 4 16 15 9 1 1 9 1 9 1 9 1 13 16 2 2 11 11 11 11 1 9 9 1 9 9 1 9 1 1 9 1 9 13 4 2
13 9 9 1 10 9 1 9 14 13 1 9 13 4
22 9 1 13 16 11 11 11 2 11 2 11 1 1 9 1 10 9 0 13 4 4 2
44 11 1 11 11 1 9 1 9 1 12 9 1 11 1 0 9 11 11 1 15 9 13 4 10 9 1 9 13 4 16 15 9 11 11 1 10 9 1 9 1 9 13 4 2
21 11 11 11 1 0 9 11 1 9 1 11 1 11 11 13 1 9 1 9 13 2
18 11 1 13 16 15 10 9 1 11 9 9 9 1 15 14 13 13 2
17 15 1 1 15 10 9 15 13 13 15 15 9 1 13 4 4 2
27 15 13 16 0 11 11 11 11 12 9 1 15 1 11 13 13 15 15 9 1 9 1 9 13 4 4 2
20 16 11 1 15 0 9 1 14 13 16 9 1 15 10 9 1 15 13 4 2
26 11 11 9 1 9 1 9 1 0 11 1 0 13 1 1 1 13 4 12 9 1 9 13 4 4 2
23 0 13 16 15 0 13 1 1 9 1 10 9 1 11 11 11 1 12 9 0 13 4 2
46 15 1 14 11 1 11 9 1 9 1 0 9 1 13 1 9 1 0 13 4 13 16 0 9 9 1 9 9 7 9 1 0 9 1 9 13 1 9 1 0 9 1 9 13 4 2
41 9 11 9 1 9 11 2 11 2 11 2 11 1 9 1 9 1 9 13 4 0 11 9 1 13 16 11 1 9 1 0 13 1 1 11 2 11 9 0 13 2
24 15 12 9 1 1 9 2 9 2 9 7 0 9 13 1 15 9 1 13 0 9 0 13 2
15 11 1 9 1 11 1 9 13 1 9 13 1 9 13 2
25 11 1 13 16 11 9 1 0 9 1 13 4 4 7 9 1 1 9 1 0 9 9 1 13 2
8 7 11 9 10 15 0 13 2
15 11 1 9 1 0 9 1 9 1 1 15 14 13 4 2
26 11 1 15 14 13 16 11 1 15 10 11 11 11 9 13 4 15 11 11 1 9 1 9 14 13 2
28 15 13 16 0 9 1 9 1 9 13 1 9 1 9 1 1 1 9 13 1 3 14 11 15 9 0 13 2
31 11 11 11 11 1 11 1 13 16 11 1 1 11 1 9 1 0 9 13 7 15 11 1 1 9 1 15 9 14 13 2
15 15 1 11 1 0 9 1 0 9 13 4 1 9 13 2
34 2 11 11 11 11 2 0 9 1 11 11 11 11 1 9 1 13 16 11 11 11 1 9 1 14 11 1 11 1 15 9 13 4 2
9 15 15 1 15 9 7 9 13 2
14 7 15 11 1 1 15 9 1 15 0 9 14 13 2
44 15 1 11 11 1 0 2 11 11 11 11 2 9 1 15 9 13 4 11 1 13 16 11 1 0 11 11 11 11 13 4 16 0 9 2 9 2 13 9 1 1 0 13 2
17 15 9 13 13 16 15 9 1 3 0 9 1 9 1 9 13 2
25 11 1 13 16 15 10 14 9 1 9 13 15 11 1 11 11 11 1 15 11 11 1 1 13 2
14 15 13 16 11 14 1 11 1 12 0 9 9 13 2
9 15 0 9 1 9 1 3 13 2
9 15 15 11 10 0 13 4 4 2
31 9 1 1 0 9 1 13 4 9 1 9 0 13 4 0 11 11 11 11 1 13 16 15 9 1 1 0 13 4 4 2
36 11 11 11 1 9 9 1 9 1 11 9 1 0 12 9 1 0 9 1 0 13 4 11 1 13 16 15 15 1 14 0 9 1 13 4 2
14 11 1 13 16 15 9 1 1 9 1 13 4 4 2
14 15 9 1 9 13 15 0 9 1 1 13 4 4 2
26 11 1 11 1 9 13 4 13 16 10 9 12 9 1 9 13 16 15 15 0 9 1 9 13 4 2
19 11 1 13 16 15 13 1 9 13 16 0 9 1 9 15 13 4 4 2
12 15 13 16 15 14 9 9 1 9 14 13 2
18 11 1 9 13 4 13 16 0 9 1 9 9 1 1 0 9 13 2
15 9 1 9 13 1 9 11 1 3 14 13 4 4 4 2
11 11 11 1 11 13 9 15 13 4 4 2
26 9 9 1 0 9 1 9 13 4 16 0 11 11 1 15 1 13 1 15 9 9 14 13 4 4 2
22 15 1 11 11 1 0 12 9 1 0 9 1 9 0 13 1 9 0 13 4 4 2
31 9 9 1 1 11 11 1 9 1 0 13 1 3 11 1 9 1 9 1 9 1 1 10 9 9 0 14 13 4 4 2
24 9 1 1 10 9 11 1 0 9 1 11 1 0 13 1 0 0 9 1 9 13 4 4 2
27 15 11 11 1 9 12 1 12 9 9 1 1 13 4 4 15 12 9 1 13 1 9 13 4 4 4 2
38 9 1 11 2 11 11 1 1 13 9 1 9 1 1 1 13 4 16 0 9 1 14 11 2 11 2 11 7 11 1 14 9 1 10 9 13 4 2
20 7 11 2 11 11 2 11 2 11 11 7 11 1 0 0 9 13 4 4 2
27 9 1 1 0 11 11 1 15 1 12 9 9 13 4 7 10 9 1 0 9 12 9 14 13 4 4 2
13 16 15 1 15 9 1 12 9 10 9 13 4 2
22 10 9 0 11 11 1 12 9 1 1 15 1 12 9 9 13 15 12 9 10 13 2
17 11 1 12 9 1 1 1 12 9 9 13 15 12 9 10 13 2
27 9 1 1 1 0 11 1 0 9 1 12 9 1 1 1 12 9 9 13 4 4 15 12 9 10 13 2
13 7 0 11 1 9 1 12 9 10 9 13 4 2
21 15 1 11 1 12 9 1 1 12 9 9 13 4 15 9 1 12 9 10 13 2
25 11 2 11 7 11 1 12 9 1 1 15 1 12 9 9 13 4 15 9 1 12 9 10 13 2
29 11 11 11 11 11 11 11 1 10 9 1 9 13 4 16 9 11 9 1 9 9 1 9 1 9 13 4 4 2
24 15 13 16 15 15 13 4 16 10 0 9 1 1 9 13 4 15 9 1 9 13 4 4 2
25 9 1 10 9 1 9 13 4 1 11 11 1 13 16 9 9 9 1 3 1 9 13 4 4 2
6 15 12 0 9 13 2
14 15 13 16 9 9 15 0 13 4 15 15 13 4 2
11 7 15 9 1 15 9 14 13 4 4 2
43 11 11 1 10 9 9 1 9 13 4 1 1 1 13 4 1 11 1 13 16 9 1 15 1 1 15 13 13 10 9 1 13 7 9 1 10 9 13 15 15 13 4 2
34 11 11 11 1 0 9 1 9 13 1 9 13 1 9 13 4 1 1 1 13 4 1 11 11 1 13 16 15 0 7 0 14 13 2
12 16 15 1 15 1 15 9 14 14 14 13 2
28 11 0 9 1 9 1 11 11 1 11 1 12 9 13 4 4 15 9 9 11 11 9 1 9 1 9 13 2
29 9 9 1 13 1 9 1 9 1 1 9 1 9 1 9 1 1 0 9 2 9 2 9 1 9 14 0 13 2
18 9 1 9 1 9 13 4 16 15 9 7 9 1 1 9 13 13 2
12 10 9 1 0 11 11 11 11 14 0 13 2
10 10 12 9 1 11 1 9 9 13 2
20 9 9 1 9 13 1 1 9 13 16 0 9 1 14 9 1 9 13 4 2
36 15 1 11 1 9 1 13 1 9 1 9 11 1 10 9 1 3 1 9 1 9 13 4 15 9 1 0 9 1 9 1 0 13 4 4 2
16 11 0 9 3 11 2 11 7 11 11 1 9 9 1 13 2
15 16 15 9 13 4 4 2 7 15 0 14 13 4 4 2
19 15 9 9 1 15 10 9 0 13 1 13 15 15 1 0 9 13 4 2
24 11 11 1 9 1 11 11 9 1 1 9 9 7 9 1 1 9 1 9 1 14 9 13 2
48 3 1 9 1 9 13 4 16 11 0 9 11 0 14 13 2 7 15 15 0 13 12 2 12 9 13 4 4 7 15 1 9 1 0 9 15 13 2 15 14 9 1 0 13 1 9 13 2
26 16 11 11 1 9 1 9 1 13 4 16 14 9 9 1 15 0 13 1 1 9 9 13 4 4 2
17 11 1 11 1 11 1 9 1 11 1 0 9 13 1 9 13 2
30 9 1 13 16 9 1 9 9 1 1 15 9 7 0 0 9 1 11 9 13 1 9 1 11 1 9 1 9 13 2
33 11 1 0 9 11 11 11 1 15 12 9 9 1 13 16 15 13 13 4 16 9 1 9 9 1 1 11 1 10 9 13 4 2
19 15 15 14 13 4 16 15 15 10 9 1 11 9 1 9 0 13 4 2
48 9 1 0 9 1 11 13 1 11 1 9 1 13 13 4 9 1 9 1 11 1 13 16 16 15 15 9 13 4 7 15 1 11 9 1 11 9 1 9 13 0 13 2 16 15 0 13 2
19 10 9 1 11 1 11 1 11 1 9 1 0 9 13 1 9 14 13 2
16 11 11 1 11 11 11 1 13 13 16 11 9 1 9 13 2
16 11 1 0 9 1 13 16 15 15 15 0 9 13 4 4 2
12 16 15 13 2 16 9 1 15 0 13 4 2
34 9 1 9 1 9 1 12 0 9 10 9 13 2 15 11 1 11 1 12 0 9 1 13 16 15 3 14 12 9 1 11 1 13 2
17 15 12 9 13 2 15 9 1 11 1 0 9 1 13 4 4 2
19 11 11 1 13 4 16 9 9 1 9 13 1 12 9 14 15 0 13 2
25 3 2 11 1 11 1 12 9 1 12 9 13 4 2 15 9 1 11 11 1 9 14 0 13 2
19 12 9 1 1 11 1 13 4 9 9 9 1 9 1 10 9 13 4 2
18 11 1 15 14 9 13 16 9 1 13 1 1 15 0 9 13 4 2
28 9 1 0 9 11 1 10 9 1 1 11 1 0 13 4 16 9 9 1 9 13 14 0 9 14 13 4 2
32 15 9 1 1 3 0 9 15 13 16 15 11 9 13 1 9 13 14 9 1 13 4 7 14 15 9 13 1 9 13 4 2
41 11 7 11 1 1 9 7 0 9 1 9 13 1 1 13 10 9 1 0 9 1 11 1 10 9 1 9 13 16 15 0 9 1 0 9 1 9 13 4 4 2
30 0 9 1 0 9 9 11 11 1 9 1 15 13 12 0 9 1 9 13 16 11 1 9 1 15 9 14 13 4 2
12 9 9 9 11 11 1 0 9 1 9 13 2
19 0 9 1 13 16 9 1 13 1 1 15 1 1 15 9 14 13 4 2
18 16 11 1 9 9 1 9 1 15 9 1 11 1 0 13 4 4 2
15 12 9 1 0 9 1 9 13 1 9 1 14 9 13 2
21 0 9 1 9 9 9 11 11 7 0 9 1 9 9 9 9 11 11 1 13 2
19 9 13 4 4 16 11 11 1 0 9 0 9 1 9 13 1 9 13 2
20 0 13 16 0 12 9 1 11 2 11 1 1 12 12 9 1 9 13 4 2
13 12 9 1 9 1 9 1 1 15 3 10 13 2
33 11 11 11 1 12 0 9 1 13 4 16 9 1 9 1 1 9 2 9 1 15 9 1 9 1 1 9 1 9 13 0 13 2
17 15 15 1 13 7 0 13 1 1 14 3 9 1 9 13 4 2
16 10 9 9 2 9 7 9 1 10 0 9 1 14 0 13 2
17 9 1 11 11 9 1 9 1 9 1 9 1 1 10 9 13 2
28 9 1 11 1 9 1 11 1 11 11 11 9 1 15 9 1 9 1 9 13 1 13 4 1 9 13 4 2
20 10 9 15 0 9 9 1 13 4 7 15 9 2 9 9 9 13 4 4 2
31 3 11 11 11 1 12 9 9 1 10 9 11 1 0 11 11 11 11 1 9 11 1 12 9 1 9 1 13 4 4 2
17 11 11 11 1 11 1 0 11 11 1 11 1 10 9 13 4 2
27 9 1 1 11 1 11 11 2 11 1 12 9 13 15 10 9 1 14 15 9 1 1 1 0 13 4 2
31 11 1 9 9 1 9 0 13 7 9 1 10 9 1 0 11 11 11 1 9 11 9 1 1 10 9 1 9 0 13 2
29 10 9 11 10 9 1 1 10 9 1 9 13 4 7 10 9 1 1 1 15 14 9 13 1 15 9 13 4 2
16 15 1 9 1 10 9 1 9 1 12 9 9 1 13 4 2
21 11 11 2 11 1 15 10 9 1 0 11 11 1 1 9 11 11 1 13 4 2
21 7 15 15 9 1 1 9 2 9 1 1 13 15 15 9 1 0 13 4 4 2
13 9 1 10 9 1 9 1 1 0 13 4 4 2
31 11 1 0 9 1 12 9 1 14 11 11 11 7 11 2 11 2 11 11 1 13 4 1 9 1 1 9 0 13 4 2
12 0 9 1 12 0 9 1 10 9 13 4 2
29 0 9 1 13 16 11 1 0 9 12 0 9 9 1 13 9 9 9 1 11 11 1 14 9 13 1 9 13 2
6 15 12 0 9 13 2
17 9 9 11 11 1 13 16 11 11 1 0 9 11 1 0 13 2
20 15 0 9 1 9 1 9 13 4 7 3 3 9 1 1 9 14 13 4 2
10 11 11 1 0 9 9 1 9 13 2
24 11 1 13 16 15 0 9 1 14 13 4 4 16 9 1 9 11 7 11 14 13 4 4 2
31 7 0 9 1 1 0 9 1 9 1 13 4 10 9 13 4 4 16 9 1 9 10 0 9 1 9 1 13 4 4 2
38 11 1 11 11 11 1 9 1 1 11 1 10 0 9 1 15 9 0 13 7 0 9 1 13 4 2 15 9 14 1 9 1 9 15 1 13 4 2
20 11 1 14 0 9 1 1 1 13 1 1 9 1 3 0 9 1 13 4 2
29 9 1 13 4 16 0 9 1 12 10 9 9 1 13 4 2 15 0 13 7 15 3 13 1 0 9 9 13 2
38 2 11 11 11 2 1 9 1 13 4 9 1 13 1 9 13 4 16 3 11 11 11 1 9 1 9 7 9 9 9 1 0 9 15 13 4 4 2
32 9 1 0 9 1 1 9 1 9 2 9 7 9 0 9 2 0 9 7 15 0 9 1 1 1 13 1 0 9 13 4 2
17 9 14 1 0 9 9 1 0 9 1 12 9 1 13 4 4 2
54 0 11 16 0 0 9 2 9 1 9 2 0 11 16 0 0 9 7 0 9 1 9 2 0 9 1 11 16 0 0 9 7 0 9 1 9 7 0 9 1 11 16 0 0 9 2 9 1 9 1 13 4 4 2
40 9 9 1 1 11 9 1 9 1 9 11 1 12 9 2 11 1 12 9 2 11 11 1 12 9 2 11 1 12 9 7 11 7 11 1 12 9 13 4 2
31 11 9 1 1 12 9 9 1 13 13 16 11 0 9 1 10 9 1 11 1 3 13 4 7 11 1 3 0 9 13 2
40 14 12 9 9 10 9 1 0 13 16 11 9 13 1 1 3 0 9 13 7 12 9 9 1 9 13 16 9 0 9 1 1 11 1 11 9 9 1 13 2
27 12 9 11 1 13 13 16 0 12 9 1 11 11 9 13 1 1 13 1 9 1 9 13 1 0 13 2
22 10 12 9 9 1 13 13 16 11 14 0 9 1 15 0 9 1 13 1 0 13 2
20 12 9 9 10 9 1 0 13 16 11 1 13 4 9 1 9 1 9 13 2
28 0 9 1 11 1 9 9 13 1 9 13 4 10 9 9 2 9 9 7 9 9 1 3 10 0 13 4 2
21 11 11 11 1 9 11 11 1 15 1 12 0 9 9 1 9 1 1 9 13 2
14 11 11 1 13 16 9 1 10 9 9 0 13 4 2
9 15 9 9 1 1 9 13 4 2
11 11 1 15 11 2 11 9 1 0 13 2
21 15 13 16 9 1 9 7 9 1 9 1 1 15 9 1 10 15 14 13 4 2
17 15 3 15 13 4 16 9 1 14 9 1 0 9 14 13 4 2
13 10 9 1 9 1 9 1 13 1 9 13 4 2
17 15 15 1 12 9 1 0 11 11 11 1 9 1 1 9 13 2
12 10 9 9 1 9 0 11 1 13 4 4 2
14 11 11 1 15 1 0 9 1 0 9 1 0 13 2
16 15 13 16 11 7 11 1 0 9 1 15 0 13 4 4 2
11 15 15 1 15 10 0 9 14 13 4 2
9 15 1 9 3 0 7 0 13 2
8 15 9 1 15 9 14 13 2
15 15 13 4 16 0 11 1 11 2 11 1 9 13 4 2
15 11 11 11 1 11 11 1 11 11 11 1 9 13 4 2
8 15 14 12 9 9 13 4 2
16 10 9 9 12 0 9 9 1 3 0 9 1 1 12 13 2
9 10 9 9 12 9 1 0 13 2
11 10 9 9 1 13 9 1 13 4 4 2
21 9 2 9 7 0 9 13 11 11 1 15 1 9 9 1 1 14 12 9 13 2
13 9 1 15 10 9 1 9 1 1 1 9 13 2
11 15 1 15 9 9 1 9 1 9 13 2
12 15 12 9 0 9 9 1 1 13 9 13 2
13 15 9 1 13 4 9 1 0 9 13 4 4 2
18 11 11 15 9 11 11 1 1 11 2 11 1 12 0 9 1 13 2
31 0 9 1 11 11 1 13 4 1 9 1 11 11 1 10 9 13 2 15 11 1 11 9 10 9 1 9 13 4 4 2
52 9 9 11 11 1 9 1 9 9 15 9 13 1 0 9 13 16 11 11 1 11 7 15 9 11 14 1 9 7 15 9 13 1 11 1 0 9 2 9 2 1 15 11 11 1 15 9 1 9 13 4 2
17 10 9 1 9 1 1 9 11 11 11 1 9 11 1 11 13 2
14 15 15 10 9 1 1 11 9 1 0 9 1 13 2
14 16 0 9 1 9 1 13 15 9 0 13 4 4 2
30 11 1 9 9 11 11 1 9 1 13 16 11 9 1 15 13 7 9 1 9 13 1 13 4 15 15 13 4 4 2
26 0 13 4 11 1 9 2 9 9 11 11 11 7 9 11 11 7 11 11 1 14 15 13 4 4 2
8 10 9 9 9 1 9 13 2
18 10 9 0 13 4 9 11 11 1 9 1 11 1 13 11 13 4 2
20 0 13 16 11 1 12 0 9 9 11 7 11 11 1 1 0 13 4 4 2
17 11 9 9 1 0 9 1 0 11 1 11 1 9 1 14 13 2
28 13 4 4 16 15 15 11 1 0 13 11 11 1 9 11 11 1 11 1 9 1 1 11 1 9 13 4 2
11 9 11 15 0 11 11 1 9 14 13 2
21 10 9 9 1 9 1 11 7 15 9 11 14 11 1 11 9 1 13 13 4 2
32 0 13 16 11 1 11 11 11 1 11 2 11 11 1 11 9 1 9 1 12 0 9 1 13 10 9 1 15 13 4 4 2
18 11 11 11 1 3 13 4 16 0 9 1 9 1 15 9 14 13 2
15 9 1 14 1 9 7 9 1 12 2 9 2 13 4 2
10 10 9 11 2 11 7 11 1 13 2
13 16 2 9 3 14 13 4 15 1 0 13 4 2
27 9 1 9 1 13 1 1 9 1 1 9 1 1 3 14 2 9 2 1 9 14 0 13 4 4 4 2
18 9 1 1 12 9 1 9 1 12 9 1 10 9 1 9 13 4 2
27 2 9 9 2 0 13 1 9 1 13 11 11 11 11 11 11 1 2 9 2 1 9 0 13 4 4 2
20 12 9 1 10 9 1 0 13 1 9 1 0 9 9 1 0 9 13 4 2
25 9 9 1 9 1 9 1 9 1 9 1 1 9 7 9 1 1 1 0 13 1 9 13 4 2
24 9 9 1 13 13 16 9 1 1 2 9 9 13 4 2 15 1 1 9 0 13 4 4 2
12 7 9 2 9 1 9 9 1 1 13 4 2
24 7 2 9 0 9 1 9 10 14 9 1 9 7 9 1 9 1 1 1 0 13 4 4 2
13 10 9 1 15 14 9 9 1 0 13 4 4 2
15 9 1 10 12 9 13 2 15 9 9 1 9 12 13 2
14 9 1 11 1 13 1 9 1 10 9 1 13 4 2
20 9 1 10 9 16 0 13 4 4 16 9 9 13 1 9 1 9 0 13 2
22 9 1 9 1 10 9 14 13 4 16 9 13 14 2 9 1 0 9 0 13 4 2
12 9 1 15 14 9 1 0 14 13 4 4 2
17 15 9 1 9 13 7 15 10 9 1 15 9 1 0 13 4 2
12 10 9 9 15 9 1 9 0 13 4 4 2
7 15 11 3 9 14 13 2
35 9 1 9 9 11 11 1 13 13 16 2 9 2 0 13 4 1 9 1 9 10 9 1 13 4 7 9 1 0 9 1 9 0 13 2
36 9 1 12 0 9 1 13 13 16 9 1 0 9 1 13 1 1 9 9 1 9 1 9 13 1 3 9 1 9 13 1 9 13 4 4 2
19 15 1 9 10 0 9 1 2 9 9 2 13 1 14 9 13 4 4 2
24 9 1 9 1 14 9 13 1 9 13 4 4 7 2 10 9 9 1 10 9 1 9 13 2
32 0 9 11 1 13 9 1 9 1 14 2 9 9 2 1 9 13 4 7 10 9 1 9 1 1 1 15 9 14 13 4 2
18 9 1 9 9 1 9 13 16 11 1 9 1 9 1 9 13 4 2
25 0 9 1 9 0 13 1 3 14 11 1 9 9 9 11 11 11 11 1 9 1 13 4 4 2
12 11 0 9 15 11 11 1 9 1 13 4 2
16 9 1 9 13 1 1 11 1 12 14 9 8 14 13 4 2
33 15 0 12 1 1 1 11 1 11 2 11 11 1 13 4 7 9 1 0 9 0 9 11 0 13 1 1 9 1 14 13 4 2
20 11 1 11 1 11 11 1 1 9 9 1 15 15 0 9 0 13 4 4 2
21 11 11 11 11 1 0 11 13 1 9 13 13 9 1 9 1 9 14 13 4 2
29 0 9 12 9 1 13 1 11 1 0 9 14 0 9 1 13 4 7 0 9 1 15 9 9 2 9 13 13 2
43 9 1 0 11 11 11 11 11 1 0 9 1 9 13 9 1 0 9 13 1 11 1 0 9 1 0 9 1 11 1 9 9 13 9 12 2 12 1 15 9 13 4 2
18 0 9 1 14 11 1 0 9 13 4 12 2 12 1 9 13 4 2
26 7 15 1 9 1 9 0 13 1 9 1 15 10 0 9 13 4 7 0 9 1 9 1 9 13 2
21 0 9 1 15 15 9 1 3 12 11 11 13 15 9 1 9 9 1 13 4 2
18 0 9 1 14 11 15 1 9 14 13 4 7 3 15 9 13 4 2
15 10 9 1 13 16 11 9 1 1 15 9 13 4 4 2
25 7 0 9 1 15 0 9 1 9 1 12 0 9 7 9 9 13 4 9 1 9 1 13 4 2
39 15 1 14 0 9 11 12 2 12 1 0 9 13 1 0 13 7 11 1 3 12 9 0 13 15 9 1 0 14 13 4 7 0 9 1 9 13 4 2
13 11 10 9 1 9 1 0 13 1 1 13 4 2
14 0 9 13 1 1 9 15 9 9 13 13 4 4 2
18 7 15 15 0 9 11 1 13 1 11 11 1 9 0 13 4 4 2
12 15 13 16 15 15 15 9 9 13 14 13 2
8 3 15 15 9 1 0 13 2
19 11 7 11 1 9 9 1 11 1 11 7 11 11 1 9 13 4 4 2
14 11 11 11 15 11 11 1 9 1 9 1 9 13 2
26 9 9 11 11 11 1 11 1 9 1 0 9 1 9 1 13 16 11 11 1 9 13 3 0 13 2
11 9 1 9 1 9 0 13 4 4 4 2
17 15 9 1 9 1 0 11 11 11 1 11 11 1 1 1 13 2
17 11 11 1 13 16 11 11 1 1 1 13 1 10 14 9 13 2
8 15 1 3 14 9 13 4 2
7 11 15 9 1 0 13 2
19 15 13 16 11 11 7 11 1 9 1 9 1 1 1 9 13 0 13 2
8 11 1 9 9 13 4 4 2
14 11 11 1 15 9 14 14 13 7 15 13 0 13 2
15 11 1 10 9 1 11 11 1 9 0 7 0 12 13 2
21 9 1 9 15 13 16 0 9 1 9 1 1 9 1 9 1 13 1 9 13 2
32 9 1 9 1 3 14 0 13 1 1 11 15 13 15 9 13 16 9 1 9 1 0 9 1 9 1 15 10 9 13 4 2
10 15 15 9 1 0 13 1 9 13 2
10 15 1 10 9 1 9 9 14 13 2
23 11 11 1 9 1 13 9 7 9 1 9 1 9 0 9 1 0 7 0 9 1 13 2
34 11 1 11 11 11 1 9 11 11 1 13 4 16 0 9 1 9 14 13 1 15 11 11 11 1 1 0 9 1 9 0 13 4 2
25 9 1 0 9 1 9 1 0 9 1 12 9 1 13 1 1 1 9 1 0 9 13 4 4 2
23 10 9 1 11 11 1 9 11 11 1 11 11 11 11 2 11 2 1 0 13 4 4 2
27 11 1 13 16 12 9 1 9 13 4 1 1 15 9 14 13 1 15 0 9 9 1 9 13 13 4 2
17 0 9 1 1 0 9 1 0 9 1 13 1 9 13 4 4 2
17 0 9 1 9 1 11 1 11 11 1 9 1 0 13 4 4 2
22 11 1 1 11 11 11 11 1 0 13 7 11 1 9 1 1 11 1 9 14 13 2
22 11 1 11 1 0 9 1 15 15 0 9 9 13 1 0 11 9 1 9 13 4 2
15 9 1 13 4 1 10 9 12 9 1 9 13 4 4 2
16 11 1 10 9 1 9 11 1 11 9 1 13 4 4 4 2
35 11 2 11 11 11 1 3 13 4 1 3 0 11 11 11 1 13 16 15 15 9 1 9 9 1 1 2 9 1 9 2 1 1 13 2
19 15 13 16 9 1 9 7 9 1 0 9 0 13 9 1 9 13 4 2
28 11 1 9 13 14 11 1 13 16 10 9 9 1 9 7 9 1 0 9 1 13 1 0 9 1 0 13 2
19 9 1 9 13 4 1 9 7 15 9 15 13 4 2 15 14 13 4 2
37 11 1 10 9 9 1 9 11 1 14 13 16 12 9 1 1 9 9 1 9 12 0 9 1 13 4 1 13 13 9 1 11 9 0 14 13 2
16 11 1 10 9 1 9 11 1 11 9 1 13 4 4 4 2
7 7 0 9 0 14 13 2
32 11 11 11 2 11 2 1 9 11 11 1 11 1 13 16 11 11 16 11 11 1 1 9 9 13 4 16 15 15 9 13 2
38 11 1 0 9 1 9 1 9 13 1 9 13 4 11 11 1 0 11 1 13 16 9 1 1 1 10 9 1 12 0 9 2 9 0 13 4 4 2
15 15 13 16 11 9 1 9 1 12 0 9 1 9 13 2
24 11 1 13 16 0 9 1 15 0 13 4 16 11 1 9 1 9 1 15 0 9 14 13 2
37 15 1 10 15 14 9 13 2 15 13 13 16 9 1 9 1 0 13 1 9 13 2 7 15 14 10 9 1 12 0 9 13 1 9 13 4 2
18 0 13 16 11 10 9 9 2 9 9 1 9 13 11 13 4 4 2
15 15 11 11 11 1 9 1 12 9 9 1 14 0 13 2
45 10 9 1 11 11 1 9 1 9 13 4 11 1 13 16 11 1 1 11 1 9 0 9 1 0 14 13 2 16 11 1 15 1 15 9 9 7 9 9 1 14 9 13 4 2
20 11 1 13 16 15 14 11 0 9 13 2 15 1 0 9 0 13 4 4 2
36 15 1 14 11 1 9 13 4 13 16 16 11 11 3 11 1 9 13 4 1 9 1 9 1 9 9 13 4 2 16 15 15 14 9 13 2
23 0 9 2 11 11 2 1 9 1 9 13 1 1 0 9 1 11 11 11 1 9 13 2
51 11 11 11 11 11 1 11 11 1 9 0 13 10 9 1 9 7 10 9 15 1 10 9 0 13 2 15 9 1 15 1 1 1 9 13 1 9 13 4 15 1 14 9 1 0 9 0 14 13 4 2
23 15 1 11 11 1 0 9 1 9 1 10 9 1 11 11 1 9 1 1 13 4 4 2
15 11 11 1 13 9 9 1 11 9 11 1 9 13 4 2
11 10 9 1 12 9 1 9 13 4 4 2
20 9 9 1 9 1 9 0 13 9 9 1 0 9 1 10 9 1 9 13 2
26 9 9 11 11 1 13 16 9 9 11 11 11 1 9 1 9 9 15 13 7 9 1 9 9 13 2
22 11 11 1 9 1 9 9 1 1 9 9 1 10 9 1 11 9 1 9 13 4 2
11 11 11 9 1 10 9 1 9 13 4 2
14 0 9 9 11 11 1 11 9 1 9 1 9 13 2
19 11 11 1 9 11 11 1 9 9 7 9 1 9 1 10 9 0 13 2
23 11 9 11 11 1 14 9 1 13 9 1 0 13 4 9 1 1 1 10 9 13 4 2
17 11 15 11 11 11 1 13 0 9 1 9 1 13 14 4 4 2
42 15 14 11 1 0 9 1 12 0 14 9 1 13 4 1 11 11 1 10 0 9 1 9 1 9 2 9 13 4 7 9 9 1 3 0 9 1 9 1 13 4 2
24 11 1 10 9 9 1 11 11 1 1 11 11 2 0 11 11 7 0 10 0 9 13 4 2
29 10 14 9 1 10 9 2 9 9 11 1 9 1 13 13 4 15 10 9 1 9 1 13 1 9 13 4 4 2
8 3 15 9 1 13 4 4 2
15 3 1 9 13 16 9 9 1 0 9 1 13 4 4 2
13 9 9 1 13 0 9 1 1 15 0 9 13 2
28 9 1 13 4 9 1 13 9 0 13 16 9 9 1 9 9 1 9 1 0 9 1 9 9 1 9 13 2
15 9 1 0 9 1 14 12 9 10 9 1 9 13 4 2
12 7 2 9 9 1 9 1 0 13 4 4 2
17 9 1 9 1 12 9 14 9 1 9 1 9 13 4 4 4 2
20 11 11 1 9 9 1 9 1 0 13 4 9 1 10 9 9 1 13 4 2
21 10 9 1 1 9 1 0 9 14 13 1 9 1 9 1 14 9 13 4 4 2
24 0 9 9 1 11 11 9 1 9 1 9 14 9 12 9 7 12 9 14 9 0 13 4 2
22 7 9 1 9 9 1 15 9 13 7 9 1 9 1 1 9 1 10 9 13 4 2
15 15 1 9 7 9 13 1 1 9 14 9 9 1 13 2
29 16 2 9 1 9 1 9 13 14 10 9 1 9 1 12 9 1 1 12 9 14 9 1 9 13 9 13 4 2
15 15 1 9 9 1 9 1 9 12 9 14 9 13 4 2
32 9 9 1 9 11 11 11 11 1 9 9 1 9 11 11 1 13 13 16 0 12 9 1 9 9 3 0 9 13 4 4 2
13 9 1 11 11 1 9 9 1 9 10 13 4 2
10 16 10 9 3 0 9 13 4 4 2
18 0 9 1 9 1 9 12 9 14 9 1 13 12 9 13 4 4 2
15 9 1 1 0 9 1 10 9 12 12 9 1 9 13 2
24 15 1 11 1 10 9 1 9 1 9 10 13 1 1 0 9 1 9 1 9 13 4 4 2
18 9 9 1 9 11 11 1 13 13 9 9 1 9 9 3 10 13 2
8 16 0 9 1 9 0 13 2
9 9 9 1 9 1 9 13 4 2
16 0 10 9 1 9 9 1 12 1 12 9 1 9 13 4 2
17 11 1 9 13 16 13 1 9 1 9 9 1 0 9 0 13 2
28 11 11 1 9 9 1 9 1 0 11 11 11 11 1 13 4 16 1 9 1 15 9 1 15 9 14 13 2
24 11 1 0 13 2 15 0 9 1 9 13 4 7 15 15 15 9 1 13 4 1 1 13 4
28 15 15 14 13 16 12 9 1 1 11 11 1 15 0 9 11 11 13 11 1 9 13 11 13 1 1 13 2
14 15 13 16 15 9 1 9 1 10 9 1 9 13 2
33 11 1 11 1 9 1 9 13 4 11 1 13 16 2 9 9 1 9 14 9 13 7 10 9 1 9 1 15 9 14 13 4 4
20 15 10 9 1 15 9 14 13 16 9 1 10 9 1 9 3 13 4 4 2
19 15 3 13 16 9 9 11 11 1 14 10 9 1 9 1 9 13 4 2
14 11 1 9 13 16 15 0 9 1 0 9 0 13 2
30 15 3 13 16 0 11 11 11 11 1 10 0 9 1 15 9 1 13 4 7 15 9 1 9 13 1 1 13 4 2
37 16 2 15 15 15 13 4 16 15 15 0 9 9 1 11 9 1 13 4 15 15 13 16 15 1 9 15 1 13 15 1 15 9 1 13 4 2
16 11 1 13 16 15 9 1 0 9 1 1 3 9 1 13 2
14 15 15 11 9 9 9 1 9 13 1 1 13 4 2
20 11 1 9 0 11 11 11 2 11 2 1 9 9 9 13 1 9 13 4 2
22 15 1 11 9 9 1 9 1 1 11 1 12 12 9 1 9 1 9 13 4 4 2
30 11 1 11 11 11 1 15 11 11 1 0 0 0 9 1 9 13 1 1 13 4 9 1 11 1 9 13 4 4 2
25 11 1 11 11 11 1 13 4 9 1 11 11 11 1 11 1 9 9 9 13 1 9 13 4 2
35 11 1 13 9 1 11 1 13 4 16 11 0 0 9 1 11 9 9 9 13 1 9 13 7 10 9 1 15 11 1 9 1 9 13 2
32 11 9 11 11 11 1 11 1 13 16 11 11 11 1 13 4 9 1 11 9 1 1 1 9 1 9 1 9 1 9 13 2
20 9 9 9 11 11 11 1 1 10 9 1 0 7 9 1 9 1 9 13 2
15 15 13 16 9 1 9 2 9 1 12 0 9 0 13 2
16 15 1 0 9 1 9 1 0 9 1 12 0 9 13 4 2
13 11 1 9 13 16 11 11 9 0 14 13 4 2
32 11 9 1 13 16 11 9 1 0 13 4 16 11 11 1 0 9 13 1 3 15 9 1 9 13 1 10 0 9 15 13 2
33 11 11 11 11 1 1 1 0 12 9 1 0 13 4 15 13 16 9 0 13 1 3 14 11 11 1 9 9 13 4 4 4 2
16 15 13 13 16 10 9 1 10 9 15 1 13 4 4 4 2
41 15 9 13 4 13 16 11 11 11 1 13 16 11 11 1 1 9 0 14 13 7 15 9 13 16 12 9 9 0 13 4 1 3 15 9 9 0 13 4 4 2
26 11 1 9 13 16 11 11 11 11 11 7 11 11 1 15 1 1 1 0 2 0 9 13 4 4 2
33 11 1 11 2 11 9 9 1 14 12 9 1 12 9 9 1 9 1 9 13 12 12 9 1 9 1 9 1 12 9 13 4 2
21 10 9 1 9 13 14 11 9 1 3 11 7 11 11 9 1 9 1 0 13 2
21 11 9 1 10 9 2 9 7 11 1 9 13 1 9 9 1 9 1 9 13 2
21 15 1 11 9 11 11 1 9 1 13 4 7 9 1 9 1 13 1 0 13 2
19 11 2 11 2 11 2 1 11 11 11 1 11 11 1 9 1 9 13 2
10 9 1 11 9 1 1 1 0 13 2
10 9 1 1 9 15 9 1 0 13 2
17 11 1 13 16 11 9 12 9 14 12 0 9 15 9 1 13 2
17 9 1 15 9 2 9 7 9 1 13 12 9 1 0 13 4 2
9 11 1 1 9 1 9 13 4 2
9 9 15 1 11 11 13 13 4 2
17 15 11 11 1 9 1 9 1 13 15 9 1 13 9 13 4 2
17 9 9 1 12 9 1 13 12 9 1 10 9 1 9 13 4 2
15 15 1 9 12 9 1 9 12 9 1 13 0 13 4 2
15 9 11 1 13 16 9 1 1 9 7 9 14 9 13 2
6 15 9 14 12 13 2
24 11 1 9 15 9 15 9 2 9 13 14 12 9 9 1 9 9 1 9 11 11 1 13 2
10 9 1 9 1 10 9 1 0 13 2
10 9 11 11 1 9 1 15 9 13 2
13 15 1 9 1 10 9 7 9 1 0 13 4 2
18 9 1 9 1 9 13 1 1 11 7 11 11 1 9 1 9 13 2
23 11 2 11 9 1 9 1 9 1 9 1 11 1 11 11 7 11 1 1 9 0 13 2
11 9 1 15 14 9 1 9 0 13 4 2
14 7 9 11 11 1 13 13 16 10 9 9 1 13 2
16 9 1 1 9 13 13 4 9 1 9 14 12 12 9 13 2
14 9 1 9 1 11 11 1 10 0 9 1 9 13 2
35 0 11 11 11 11 1 15 9 1 11 1 10 2 0 2 9 1 9 13 11 1 11 9 1 11 1 9 1 9 13 1 9 13 4 2
31 15 13 13 16 10 9 1 0 9 1 14 11 9 11 11 1 9 1 9 1 10 9 13 15 1 9 1 9 13 4 2
46 15 11 9 1 0 9 13 7 11 11 7 11 11 1 1 9 13 4 11 1 9 13 16 10 11 9 7 11 1 10 0 9 1 0 9 1 15 11 13 1 9 1 9 13 4 2
41 11 11 11 1 15 9 2 11 11 11 11 11 2 1 13 4 16 9 1 11 11 1 0 9 1 10 0 9 1 14 11 9 1 1 11 1 9 0 13 4 2
23 7 3 15 0 9 14 13 1 11 1 11 11 11 1 14 11 9 1 1 9 13 4 2
31 15 0 9 1 13 9 1 11 1 13 16 11 1 11 9 1 15 9 10 11 9 1 9 2 9 1 1 0 13 4 2
13 15 10 9 13 15 9 9 1 14 0 9 13 2
37 15 13 16 11 1 9 1 1 15 11 1 15 13 1 9 13 16 15 9 9 1 10 0 9 1 9 13 4 15 11 1 15 1 13 0 13 2
23 11 11 1 0 9 1 15 9 13 16 9 1 11 1 3 11 1 9 1 9 13 4 2
25 10 9 14 12 9 1 9 1 2 9 2 1 2 9 2 7 14 0 2 9 2 1 0 13 2
55 11 1 11 11 1 1 1 11 1 13 1 1 9 9 1 9 13 1 11 1 13 16 16 11 1 15 9 14 13 1 9 11 1 3 14 13 4 16 11 11 9 1 1 11 1 15 0 9 1 11 1 9 13 4 2
20 9 0 9 13 16 11 7 11 11 12 14 9 1 1 11 1 9 14 13 2
21 13 9 1 9 1 11 1 0 9 9 7 9 1 0 13 1 9 13 4 4 2
20 11 11 11 11 1 11 1 13 16 15 1 0 9 1 9 8 10 13 4 2
23 15 1 14 11 11 1 13 16 11 1 11 1 9 9 1 0 9 1 14 9 13 4 2
24 15 13 16 11 11 11 1 9 1 0 9 10 9 1 9 1 7 14 11 1 13 4 4 2
9 0 9 9 10 0 7 0 13 2
17 9 1 1 15 9 1 0 7 0 13 9 1 9 1 13 4 2
20 10 9 1 13 1 1 9 9 9 7 9 0 13 1 10 9 1 9 13 2
49 9 9 1 9 9 7 0 9 9 1 9 1 9 1 9 13 4 11 11 1 13 16 9 1 9 13 16 11 11 11 1 9 1 0 9 3 10 9 1 9 1 7 14 11 1 13 4 4 2
25 15 1 14 9 9 1 9 1 0 9 1 0 9 1 9 1 0 13 1 1 1 15 9 13 2
32 11 11 1 9 1 15 13 13 4 16 11 1 0 9 1 9 9 1 1 0 13 1 1 0 9 1 0 9 15 13 4 2
20 11 11 11 1 13 16 11 1 11 1 9 9 1 0 9 1 9 13 4 2
12 0 9 1 13 1 9 1 12 9 9 13 2
28 15 13 16 9 10 9 1 9 13 4 4 7 15 1 15 14 9 11 1 11 9 0 13 1 3 13 4 2
19 11 1 11 11 11 1 13 4 16 11 1 9 1 11 0 9 14 13 2
17 15 13 16 11 9 1 9 1 1 12 9 1 0 9 13 4 2
37 11 11 11 1 9 1 1 12 9 1 11 1 11 1 11 9 1 9 1 1 9 9 1 0 9 1 1 1 9 13 1 9 1 14 9 13 2
37 15 13 16 11 9 1 9 1 9 1 0 9 1 1 1 0 9 13 4 4 7 10 9 1 11 1 15 14 0 9 1 11 14 0 9 13 2
39 12 0 9 9 1 11 1 1 1 13 4 16 12 9 1 9 2 9 7 9 1 1 11 9 1 9 13 4 4 15 11 1 9 1 15 1 0 13 2
16 15 13 16 16 11 9 13 4 16 15 1 11 14 0 13 2
8 10 9 15 14 0 14 13 2
23 9 14 1 9 13 11 2 11 9 9 1 11 1 0 9 0 13 1 12 0 9 13 2
48 16 2 10 9 1 11 11 11 1 11 9 2 0 2 11 11 2 11 11 11 1 11 11 11 2 11 2 11 11 11 2 11 2 1 9 11 11 7 11 11 11 1 11 9 1 9 13 2
20 11 1 11 11 9 13 1 9 1 11 11 1 0 15 9 0 13 4 4 2
10 16 10 9 9 1 0 9 13 4 2
17 9 9 1 9 1 11 2 11 1 9 13 1 9 13 4 4 2
34 9 1 11 9 11 11 11 1 9 1 13 16 3 15 15 13 4 16 9 9 1 11 1 11 1 9 13 1 15 9 13 4 4 2
23 11 1 13 16 11 11 1 11 1 9 0 9 1 10 9 1 0 9 1 1 1 13 2
13 9 1 10 9 9 1 10 9 9 2 9 13 2
26 11 2 11 2 1 9 11 11 7 11 11 1 11 1 10 0 9 11 1 9 2 9 1 9 13 2
36 11 9 11 11 11 1 2 9 1 9 2 1 9 13 4 11 1 13 16 9 1 9 15 7 11 1 0 9 1 15 1 15 0 14 13 2
29 0 11 11 1 9 1 10 9 1 9 1 9 13 4 0 11 9 1 9 1 9 11 1 9 1 14 13 4 2
28 11 11 11 11 11 11 11 11 1 13 16 9 10 9 1 9 13 1 1 15 11 11 11 1 9 9 13 2
14 10 9 15 11 1 14 13 7 11 1 0 14 13 2
13 15 13 16 9 1 3 14 9 13 4 0 13 2
19 9 1 13 1 10 9 1 9 1 1 0 13 16 9 9 1 9 13 2
23 15 9 1 13 16 9 1 9 1 13 4 4 4 16 10 9 1 9 1 1 9 13 2
17 15 13 16 9 1 13 1 1 9 9 1 0 7 0 9 13 2
8 15 1 12 1 9 13 4 2
26 15 1 9 9 11 1 13 16 11 1 0 11 11 7 11 1 10 9 1 15 0 9 13 4 4 2
14 10 9 1 9 0 12 9 1 10 9 1 0 13 2
21 0 11 11 11 1 15 1 12 9 9 13 4 4 7 12 1 9 13 4 4 2
10 10 9 1 9 0 14 13 4 4 2
14 9 1 10 9 1 9 1 1 15 9 0 13 4 2
16 15 13 16 10 9 1 13 0 9 9 1 9 1 14 13 2
14 16 15 13 16 9 0 12 9 1 3 14 13 4 2
15 15 11 1 11 9 1 1 15 1 14 0 9 13 4 2
30 10 0 9 1 1 11 11 11 11 15 9 0 14 13 13 10 9 9 1 9 11 1 9 1 0 9 13 13 4 2
13 11 1 11 1 9 1 14 0 9 10 0 13 2
16 11 7 11 1 9 1 1 0 9 0 9 1 0 13 4 2
21 15 1 0 9 0 9 1 1 13 15 2 15 1 9 13 1 9 1 9 13 2
17 11 1 0 9 1 1 16 0 9 13 4 16 3 9 0 13 2
25 9 9 1 0 9 9 1 3 13 1 9 13 1 11 11 11 11 11 1 9 1 10 0 13 2
32 9 1 9 9 11 11 1 1 2 15 3 14 0 9 1 9 1 13 10 9 1 15 9 13 16 3 10 9 14 13 4 2
10 15 0 9 1 9 1 0 13 4 2
30 11 9 1 10 3 1 13 1 11 11 13 4 16 11 7 15 0 9 1 13 1 9 1 0 9 1 9 14 13 2
14 9 1 10 9 1 15 2 15 1 9 0 13 4 2
20 7 11 1 10 9 11 1 11 1 1 9 13 15 11 1 0 13 0 13 2
18 14 10 9 1 9 9 1 9 15 2 15 1 1 9 13 4 4 2
9 15 1 0 9 1 9 0 13 2
16 11 0 9 1 9 1 13 1 1 9 1 9 13 13 4 2
33 15 13 16 9 1 13 1 9 1 14 16 11 1 0 9 1 10 9 13 16 0 9 12 9 1 9 13 1 1 0 13 4 2
12 11 1 11 1 9 1 0 9 10 0 13 2
29 11 1 9 1 0 13 4 15 13 13 16 15 9 1 14 11 11 11 1 11 1 9 13 1 1 13 4 4 2
16 11 11 1 0 9 11 11 11 15 1 11 1 0 13 4 2
19 15 13 13 16 9 1 0 13 1 9 13 1 9 1 10 9 13 4 2
10 15 15 9 1 14 0 9 13 4 2
10 11 1 15 13 15 9 1 9 13 2
54 11 9 1 11 1 11 9 1 9 1 9 1 10 9 1 9 1 9 13 7 9 1 9 7 9 1 0 9 13 1 1 9 1 1 15 9 1 9 13 1 1 9 13 1 9 1 11 11 1 0 9 13 4 2
48 9 9 11 11 11 7 9 11 11 11 1 9 1 9 9 1 9 1 10 9 1 9 9 13 7 9 9 0 13 1 1 11 1 1 1 13 4 1 9 1 9 1 9 13 1 13 4 2
19 9 1 0 9 11 11 11 11 11 11 11 11 1 9 1 10 9 13 2
17 11 11 1 0 9 11 11 1 11 1 11 11 11 1 9 13 2
12 15 9 11 11 11 1 11 1 10 9 13 2
29 11 9 1 10 9 11 1 9 1 9 0 13 7 11 11 11 1 9 13 1 1 9 13 1 0 13 4 4 2
35 9 1 11 1 11 9 1 3 15 9 1 0 7 0 9 1 11 9 1 9 1 1 11 7 11 11 11 13 1 9 13 1 9 13 2
19 15 11 1 9 1 1 15 9 1 11 11 11 1 13 1 9 14 13 2
19 11 1 9 1 1 9 1 13 16 11 13 1 15 11 1 13 13 4 2
25 15 13 2 11 1 15 15 9 1 9 1 11 11 1 9 12 9 11 1 13 1 9 13 4 2
15 11 11 11 1 9 1 15 15 15 0 9 14 13 4 2
42 15 13 16 15 12 9 1 9 1 13 15 15 13 1 9 13 4 16 9 9 1 11 1 9 1 0 13 14 11 9 1 0 2 0 7 0 9 14 13 4 4 2
15 11 1 9 9 13 1 10 9 1 15 9 1 9 13 2
33 15 13 16 15 13 4 16 11 1 9 13 1 9 1 0 13 1 1 15 11 11 11 7 11 11 1 9 1 14 0 13 4 2
26 0 13 16 10 0 9 1 9 9 1 9 9 1 9 0 10 9 1 13 12 1 12 13 4 4 2
32 15 15 11 1 11 11 11 2 9 11 11 11 1 11 11 2 11 11 11 1 11 11 7 11 11 11 1 11 11 0 13 2
22 16 11 11 15 0 13 4 4 16 11 1 11 1 9 13 1 9 14 0 13 4 2
21 16 11 1 9 11 11 11 1 13 4 16 15 3 14 9 3 13 1 9 13 2
20 15 13 4 16 11 11 13 1 9 1 9 12 2 12 9 1 13 4 4 2
25 11 11 3 14 10 9 1 9 13 13 4 4 2 15 3 9 1 9 1 9 9 1 13 4 2
20 9 1 13 13 16 9 9 3 15 15 9 1 9 9 7 9 1 9 13 2
28 10 9 9 1 1 10 9 1 3 9 1 9 1 9 3 13 4 7 15 1 9 9 11 1 0 13 4 2
22 7 9 9 13 1 3 9 1 0 9 1 9 13 4 10 9 11 11 13 4 4 2
27 7 9 9 10 9 14 13 16 9 1 10 9 9 1 0 13 7 9 0 13 1 3 15 1 15 13 2
21 11 9 1 11 11 2 11 7 11 1 10 9 1 9 1 9 1 9 13 4 2
34 9 1 9 1 1 10 11 9 1 1 9 14 1 14 12 12 9 11 2 12 12 9 11 7 12 12 9 11 9 1 0 13 4 2
16 16 9 1 11 1 10 9 1 1 9 1 10 9 13 4 2
32 11 11 1 12 0 9 1 1 9 9 15 1 1 14 13 16 9 1 1 10 9 11 11 1 0 13 15 9 1 15 13 2
19 15 13 13 16 3 9 10 9 1 9 13 4 7 15 9 10 13 4 2
25 15 11 11 15 10 9 1 10 9 13 4 4 16 9 1 0 9 1 0 9 1 9 13 4 2
28 15 13 13 16 9 9 13 1 3 14 9 1 10 9 13 4 4 16 15 0 9 1 9 14 13 4 4 2
14 11 11 11 1 10 9 1 9 13 1 1 13 4 2
18 9 1 13 13 16 9 9 9 1 9 7 9 1 9 1 9 13 2
14 9 1 9 13 2 15 1 15 9 9 1 9 13 2
37 11 1 11 11 11 1 13 16 9 1 9 1 9 0 13 9 0 13 1 1 11 7 9 9 0 0 9 11 1 0 9 13 1 9 1 13 2
15 15 15 0 7 0 9 1 9 13 1 9 1 14 13 2
14 7 15 1 0 9 1 9 13 1 15 9 14 13 2
15 11 1 13 16 15 11 11 1 14 10 9 13 4 4 2
19 11 11 1 0 13 4 4 16 9 1 1 9 1 9 3 13 4 4 2
26 11 1 11 1 12 9 1 9 1 13 1 9 1 15 9 0 13 1 1 9 13 1 9 13 4 2
9 14 11 1 10 9 1 9 13 2
23 15 0 9 13 16 0 9 10 9 1 9 1 1 10 9 14 9 1 14 13 4 4 2
58 11 11 1 11 11 1 13 4 9 1 11 2 11 11 11 11 11 1 9 0 0 9 1 13 9 1 1 9 2 9 1 9 1 10 9 1 10 9 13 16 15 0 9 14 12 12 9 13 15 0 9 1 9 1 14 10 13 2
13 15 9 1 9 1 1 14 0 9 0 14 13 2
47 0 0 9 9 13 4 11 11 11 1 11 1 9 1 9 7 9 1 9 13 4 13 16 9 1 9 1 9 1 1 3 12 2 12 12 9 0 13 4 15 15 1 9 9 13 4 2
20 11 1 11 11 1 13 16 14 12 2 12 9 9 14 0 9 1 0 13 2
21 10 9 11 1 1 15 9 1 9 13 4 4 15 0 9 1 9 13 4 4 2
29 15 13 16 9 1 9 13 1 1 12 12 9 1 9 13 4 4 7 10 9 1 14 9 14 13 4 4 4 2
22 11 1 11 11 1 10 9 1 0 9 13 4 13 16 3 9 1 15 9 13 4 2
22 9 1 9 9 1 1 0 13 7 15 0 14 13 16 15 15 9 13 1 9 13 2
29 15 13 16 9 13 4 7 15 15 14 13 4 16 9 9 1 1 9 1 0 9 12 9 1 3 13 4 4 2
9 15 3 10 9 1 9 13 4 2
22 11 11 1 9 13 16 12 12 9 9 1 9 15 9 1 9 1 9 15 13 4 2
25 9 1 9 13 1 9 1 9 3 1 15 13 4 4 16 15 9 1 1 9 9 14 13 4 2
21 11 11 1 13 16 11 11 1 1 15 15 0 9 1 13 1 1 9 14 13 2
39 11 1 11 11 11 11 1 9 13 4 16 11 1 11 11 1 9 1 11 1 14 0 9 9 7 0 9 1 0 0 9 2 9 2 1 9 13 4 2
17 15 9 2 9 9 9 2 0 13 1 9 1 9 14 9 13 2
27 11 11 1 11 1 12 9 1 11 11 11 2 11 2 1 0 9 1 15 1 9 1 0 13 4 4 2
18 15 13 16 11 1 0 9 1 1 15 13 4 4 2 15 14 13 2
28 11 1 13 16 11 1 0 0 9 1 0 13 4 7 11 1 0 9 9 10 9 1 9 1 9 13 4 2
25 15 13 16 11 1 1 11 1 14 9 1 13 4 7 15 1 9 9 13 1 9 13 4 4 2
25 9 1 9 1 14 11 1 11 11 1 9 1 0 12 9 9 1 12 9 9 1 9 13 4 2
20 10 9 12 0 9 11 11 1 13 4 4 7 15 12 9 1 0 13 4 2
14 15 13 16 9 1 11 11 11 1 9 13 4 4 2
11 15 1 11 9 1 12 9 14 13 4 2
11 15 1 1 11 9 1 9 13 4 4 2
23 9 9 1 9 1 13 7 0 9 1 0 13 1 1 9 1 0 9 1 9 13 4 2
13 15 9 7 9 9 1 9 1 0 13 4 4 2
41 11 1 13 16 11 11 1 0 0 0 9 1 1 1 15 1 11 1 0 9 1 9 1 1 12 9 0 13 4 2 15 9 1 12 12 12 9 1 9 13 2
34 15 1 11 11 11 1 9 11 11 11 1 11 1 9 13 4 11 1 9 1 11 1 14 9 9 13 7 11 0 13 1 9 13 2
24 15 11 0 13 1 9 1 11 1 0 9 1 9 13 16 15 10 9 1 9 13 15 13 2
27 9 11 11 11 1 11 1 0 9 9 7 15 1 9 1 1 12 12 12 9 1 0 9 1 9 13 2
20 9 7 9 1 0 9 1 1 1 9 9 9 11 1 11 1 9 13 4 2
19 9 9 1 9 14 1 12 9 1 1 15 12 9 1 9 0 13 4 2
13 9 1 13 13 16 11 1 11 1 9 13 4 2
14 15 9 9 1 10 9 13 16 15 9 9 1 13 2
17 11 11 1 11 9 1 15 9 1 1 1 9 13 1 13 4 2
16 11 11 11 11 11 11 11 1 12 9 1 9 1 11 13 2
27 9 2 9 1 15 9 1 1 11 11 11 2 11 2 11 11 11 11 2 0 9 7 0 9 0 13 2
9 11 9 2 9 1 3 9 13 2
39 15 9 1 1 11 1 11 11 1 1 11 11 11 1 0 9 1 1 9 13 11 11 1 13 9 1 1 9 7 9 1 0 9 1 9 1 9 13 2
19 3 1 15 11 11 0 9 1 0 2 0 9 11 11 11 1 9 13 2
24 15 11 1 11 11 1 11 11 11 11 11 11 1 11 11 9 1 9 9 1 14 9 13 2
16 11 1 11 11 11 1 9 9 1 0 9 1 14 9 13 2
16 10 9 1 11 11 11 11 11 7 11 11 11 14 0 13 2
9 11 11 9 9 11 11 13 4 2
32 11 11 1 9 1 11 1 12 9 1 9 13 9 7 11 1 0 9 1 9 1 15 1 1 3 0 9 1 9 13 4 2
14 15 0 9 1 9 9 7 9 2 9 14 0 13 2
15 15 10 9 13 15 13 15 9 1 9 1 9 13 4 2
18 9 1 15 9 1 10 0 9 1 9 1 9 13 4 9 13 4 2
21 10 9 1 9 1 12 9 9 1 12 9 7 9 9 1 0 13 4 4 4 2
30 9 1 9 11 11 11 1 13 16 9 0 13 4 9 1 10 9 15 13 4 15 15 9 1 1 0 13 4 4 2
22 11 1 0 12 9 1 12 0 0 9 1 9 9 7 12 0 0 9 9 13 4 2
16 15 1 2 3 0 9 1 0 9 2 9 1 9 14 13 2
31 15 0 9 1 12 9 1 12 9 2 12 1 12 9 2 12 1 12 9 7 9 1 12 1 12 9 0 13 4 4 2
17 9 1 13 16 10 9 11 11 1 14 9 1 13 4 4 4 2
24 11 1 1 10 9 9 7 9 11 11 1 11 11 9 1 11 1 0 9 9 1 13 4 2
23 10 9 1 15 11 11 9 1 0 9 1 9 9 7 12 0 9 1 0 13 4 4 2
18 15 1 10 9 1 9 1 9 13 15 9 9 1 14 9 13 4 2
30 12 9 1 9 1 15 13 16 9 9 15 1 13 4 13 7 15 9 12 9 1 14 11 11 1 15 13 4 4 2
10 15 9 0 13 4 9 9 1 13 2
39 15 11 1 13 4 16 12 9 9 1 3 10 9 2 9 1 9 13 4 4 2 15 9 1 9 1 9 13 16 9 1 9 9 1 9 13 4 4 2
28 12 9 1 9 1 9 13 1 13 9 1 1 15 9 13 1 1 11 13 4 9 1 0 11 13 4 4 2
36 9 9 11 2 11 1 9 11 11 1 15 0 9 11 11 1 9 1 1 1 9 13 15 15 14 9 13 9 1 0 11 1 1 13 4 2
27 9 1 10 9 1 15 14 9 1 9 14 13 7 9 14 12 9 9 11 11 11 11 11 1 13 4 2
27 9 1 1 2 9 1 0 0 9 1 9 1 10 9 1 3 9 13 16 15 12 9 13 1 9 13 2
11 9 1 11 1 9 12 9 9 13 4 2
20 9 1 9 11 11 7 9 11 11 1 9 9 1 0 9 1 9 0 13 2
32 0 13 16 0 11 11 1 14 12 9 1 9 13 1 1 11 11 1 11 1 11 13 4 12 9 1 11 1 13 4 4 2
33 11 7 11 1 11 2 11 1 9 9 1 9 1 1 0 9 9 13 1 9 1 11 1 11 1 9 9 1 0 9 13 4 2
37 9 9 1 11 1 11 9 1 9 1 0 9 11 9 11 11 7 0 9 11 11 1 9 1 9 14 13 1 9 1 9 11 11 1 13 4 2
32 9 9 9 9 9 9 11 11 1 9 1 9 1 1 1 15 9 1 13 4 9 1 9 13 4 7 9 1 9 13 4 2
34 12 9 1 11 1 10 12 9 9 13 15 11 7 11 11 1 9 9 1 15 9 1 9 13 7 9 13 4 9 1 1 9 13 2
13 15 10 9 13 15 15 0 13 9 1 13 4 2
20 10 9 1 1 9 2 9 13 14 4 15 9 7 9 15 1 13 4 4 2
36 15 12 9 13 4 16 15 14 15 9 13 4 15 12 9 1 9 9 1 1 11 1 9 13 1 10 9 1 9 13 1 9 13 4 4 2
14 15 10 9 13 4 15 15 9 1 9 13 4 4 2
24 15 0 9 13 0 9 1 9 11 11 1 0 13 9 13 16 11 7 11 1 9 13 4 2
27 15 9 13 0 13 11 1 9 1 3 9 13 13 0 9 1 10 0 13 16 15 9 1 6 13 4 2
16 9 11 1 15 11 1 15 1 13 7 3 9 13 1 13 2
17 10 3 10 0 9 1 12 9 9 1 9 13 15 0 13 4 2
12 11 1 15 3 9 13 7 15 9 1 13 2
19 15 9 1 9 3 13 15 0 9 1 0 0 9 1 9 1 15 13 2
14 11 1 13 16 10 9 1 15 9 1 9 13 4 2
38 10 0 9 1 9 13 4 10 9 1 1 10 9 15 10 9 0 2 0 9 15 1 0 9 11 11 1 9 13 4 15 3 1 9 9 14 13 2
17 11 1 9 15 12 9 1 9 13 7 0 9 9 1 13 4 2
40 11 11 1 0 9 1 0 9 13 4 13 16 11 2 11 1 10 9 1 9 9 1 9 13 4 7 10 9 15 13 1 9 13 15 1 9 1 13 4 2
45 11 1 9 1 9 2 12 9 1 9 7 0 9 1 9 1 9 13 1 9 1 11 1 13 16 15 14 15 0 13 13 4 16 9 1 9 13 1 9 15 9 14 13 4 2
25 11 9 1 9 11 1 11 11 1 9 9 13 1 9 1 13 16 15 15 15 9 14 13 4 2
6 9 3 3 9 13 2
18 3 2 9 1 1 10 9 1 9 1 9 11 1 14 13 4 4 2
26 15 1 14 0 11 9 1 14 11 2 11 1 10 9 1 9 13 11 1 9 1 14 3 13 4 2
25 16 15 10 9 14 13 16 11 1 9 1 11 9 1 9 1 9 1 9 1 9 0 14 13 2
24 11 11 1 13 16 11 9 11 9 1 12 0 9 13 11 11 7 9 1 9 1 9 13 2
14 10 14 9 10 9 1 9 13 13 15 9 13 4 2
29 12 0 9 1 9 1 15 13 16 9 9 1 0 9 1 0 13 1 1 9 1 14 15 1 0 9 13 4 2
25 15 13 16 9 9 9 1 0 9 1 0 13 1 1 14 12 9 9 13 1 9 13 4 4 2
46 11 11 11 11 1 11 11 1 9 13 4 11 7 11 1 12 0 9 1 1 3 11 1 9 13 1 9 13 3 11 1 12 9 1 1 13 4 9 9 1 9 1 9 13 4 2
18 0 9 1 1 15 0 11 11 1 12 9 1 15 0 11 9 13 2
17 15 9 1 1 1 11 11 11 11 1 0 9 1 9 13 4 2
16 15 1 11 1 0 11 11 11 11 1 11 1 9 13 4 2
7 10 9 11 11 11 13 2
18 11 11 15 9 1 0 9 1 11 1 11 1 0 9 1 11 13 2
15 11 1 15 11 11 11 7 11 11 11 1 1 9 13 2
12 12 9 1 1 9 1 9 0 9 13 4 2
28 3 1 15 10 9 11 1 1 0 13 4 15 15 15 1 11 11 11 11 11 1 0 9 1 1 9 13 2
25 11 11 1 13 1 1 11 1 11 11 1 9 13 1 9 1 11 1 11 1 15 9 13 4 2
13 11 1 13 13 16 11 1 10 9 0 14 13 2
23 15 11 1 11 1 0 9 1 1 1 13 4 15 15 13 16 15 0 9 1 9 13 2
19 11 1 3 13 4 13 16 12 9 1 10 9 1 9 1 9 13 4 2
26 11 2 11 1 1 0 9 1 10 9 1 15 9 13 1 9 13 15 13 11 2 11 0 9 9 2
15 11 1 13 16 11 9 0 9 11 9 1 9 1 13 2
20 15 1 1 14 10 9 15 14 15 9 1 12 9 1 1 9 13 4 4 2
15 15 13 16 12 9 1 1 8 10 9 3 15 14 13 2
30 11 11 11 11 11 11 1 11 1 11 1 11 9 0 13 4 11 1 1 1 14 15 9 13 4 1 9 13 4 2
18 7 11 11 11 2 11 2 1 10 9 1 9 13 1 9 13 4 2
11 11 1 9 15 1 11 14 13 4 4 2
20 9 9 11 1 11 1 11 1 1 15 9 15 9 11 11 1 1 13 4 2
15 15 9 14 1 9 1 0 9 1 1 1 13 4 4 2
12 11 11 1 10 9 11 11 1 9 1 13 2
50 11 11 1 9 11 11 1 11 1 9 13 4 13 16 11 0 11 2 15 13 9 7 9 15 12 9 1 13 4 2 15 11 9 13 7 15 0 13 16 11 11 11 1 1 14 15 9 13 4 2
22 16 11 1 15 9 1 15 14 13 16 11 1 9 1 1 1 9 3 1 13 4 2
9 15 15 9 15 0 14 13 4 2
42 15 9 1 9 9 9 2 11 2 1 9 13 16 15 11 7 9 9 1 0 9 7 11 11 11 11 11 1 9 1 9 13 10 11 9 11 1 9 9 0 13 2
18 0 0 11 1 9 11 1 10 9 1 11 1 9 1 14 13 4 2
11 15 10 9 1 0 0 9 1 9 13 2
19 11 9 1 9 11 11 11 9 13 4 1 1 9 1 9 1 0 13 2
27 15 11 7 11 11 1 9 13 4 13 16 0 9 1 1 14 10 9 1 9 1 9 11 14 13 4 2
31 11 11 1 11 11 0 9 1 12 9 0 13 13 4 16 11 12 11 9 13 7 15 15 9 2 9 2 0 13 4 2
11 15 1 9 1 11 1 9 13 9 13 2
25 15 9 1 11 1 15 9 13 4 13 16 11 12 0 9 13 2 15 9 11 11 1 0 13 2
9 15 11 11 15 9 14 13 4 2
15 11 1 10 9 1 9 1 11 11 1 15 9 1 13 2
13 9 13 1 1 1 11 11 1 9 1 13 4 2
17 11 1 0 13 16 11 11 7 0 9 1 1 11 9 0 13 2
11 9 11 1 15 9 1 15 9 13 4 2
14 9 9 11 15 1 0 13 2 15 15 9 14 13 2
22 15 0 9 1 9 1 13 16 0 9 1 1 14 11 9 1 15 13 1 9 13 2
7 15 9 1 15 9 13 2
30 11 1 0 9 1 9 0 13 4 4 7 15 0 7 0 9 1 1 0 9 3 9 9 13 1 9 13 4 4 2
21 11 2 11 7 11 1 0 7 3 0 9 1 13 1 1 9 9 13 4 4 2
20 9 1 10 9 0 9 1 9 13 15 1 9 7 9 1 9 13 4 4 2
28 11 2 11 2 1 9 13 9 1 13 4 16 11 1 9 1 3 0 9 1 9 1 10 9 14 13 4 2
40 11 1 15 9 1 11 1 12 0 9 13 10 12 9 1 9 13 4 15 10 9 1 9 13 4 7 15 0 12 9 1 11 2 9 7 9 13 4 4 2
25 10 9 1 11 11 1 9 1 15 13 1 9 13 4 16 15 9 7 0 9 1 0 9 13 2
24 9 1 11 1 15 9 13 4 2 9 1 9 2 2 11 11 2 1 9 1 9 13 4 2
44 3 0 3 11 2 11 2 1 15 9 1 11 1 2 9 1 9 2 13 4 13 4 16 15 9 7 0 9 1 9 13 15 1 7 15 9 1 0 13 1 9 13 4 2
27 11 11 1 9 1 0 3 11 11 1 11 11 11 1 11 1 11 11 11 1 9 1 10 9 13 4 2
13 15 10 12 9 1 1 12 1 15 15 9 13 2
35 12 0 9 1 11 9 9 12 9 1 11 11 11 11 13 7 11 1 9 1 11 9 1 12 9 1 1 15 0 9 1 9 13 4 2
28 9 1 13 16 9 9 11 11 11 1 9 1 11 9 13 1 13 0 9 1 0 9 1 1 10 9 13 2
16 9 1 15 1 1 11 7 11 9 11 11 1 0 13 4 2
18 0 9 11 9 2 11 11 7 11 1 11 11 11 1 14 9 13 2
32 11 1 12 0 9 1 13 1 3 11 1 11 1 9 9 1 13 16 15 10 9 1 9 1 1 9 13 1 9 1 13 2
18 7 16 15 9 0 14 13 4 2 16 15 9 1 9 13 4 4 2
22 11 1 13 16 11 1 0 9 1 11 1 9 1 9 1 9 13 1 9 13 4 2
17 15 13 16 9 1 13 1 1 11 1 9 7 9 0 13 4 2
8 15 15 10 9 1 0 13 2
21 15 13 16 15 0 13 4 16 0 9 1 0 9 11 1 9 1 13 0 13 2
19 9 11 11 1 0 9 1 11 11 1 11 11 1 15 9 0 13 4 2
41 9 1 11 1 0 9 1 10 9 1 0 13 1 9 13 4 2 15 9 1 1 13 4 11 11 11 11 1 9 0 9 1 13 1 9 1 13 4 4 4 2
26 11 11 1 1 15 9 1 13 4 12 9 1 13 4 7 12 9 1 0 13 1 9 13 4 4 2
23 10 9 1 9 0 9 1 13 1 1 15 3 0 9 7 15 9 1 9 0 13 4 2
18 15 9 1 11 1 9 1 1 9 11 11 1 15 9 0 13 4 2
17 15 1 0 9 1 11 11 1 11 1 9 1 0 13 4 4 2
39 9 1 13 4 16 0 9 1 9 9 1 9 7 0 9 1 9 7 9 1 9 13 1 1 13 4 4 2 7 11 1 9 1 10 15 14 14 13 2
23 11 1 13 13 16 11 10 9 1 9 1 13 4 15 1 15 9 1 9 0 13 4 2
36 0 13 16 11 0 9 1 9 1 9 1 13 1 1 11 1 9 13 1 1 13 4 4 16 11 11 0 13 1 9 1 9 13 4 4 2
34 3 11 1 15 1 11 1 11 9 1 1 0 9 1 13 1 9 1 1 9 13 4 7 15 0 9 1 0 13 1 9 13 4 2
17 0 11 9 1 1 11 11 13 0 9 1 12 9 13 13 4 2
31 0 9 1 9 1 14 11 0 9 1 13 11 11 1 9 13 4 7 11 1 9 1 0 13 1 9 1 13 4 4 2
31 15 11 1 1 3 10 9 13 0 13 2 15 11 1 9 9 1 9 1 13 1 1 11 1 9 13 1 1 13 4 2
48 11 9 11 11 1 1 2 0 9 11 7 9 0 2 0 9 13 13 4 4 16 11 0 9 9 1 9 1 11 1 9 13 7 11 1 9 13 4 16 15 15 1 15 0 9 14 13 2
17 11 1 14 15 9 15 13 16 15 10 9 9 14 13 4 4 2
25 11 10 9 1 14 9 1 9 1 13 16 11 13 11 9 9 1 1 15 9 14 13 4 4 2
25 11 1 1 2 11 7 11 1 9 9 1 9 1 13 1 0 13 7 15 11 1 9 1 14 13
15 11 1 13 13 16 15 10 9 1 15 0 9 14 13 2
17 11 1 9 13 16 13 9 1 13 1 9 1 9 13 4 4 2
13 11 2 11 11 1 11 1 12 0 9 13 4 2
12 9 1 0 9 1 3 9 7 9 13 4 2
16 3 1 9 1 11 9 1 10 9 13 4 8 3 13 4 2
38 11 9 14 12 12 9 11 2 11 11 2 11 2 15 11 9 1 10 14 3 13 4 16 3 1 0 0 9 1 9 1 9 1 1 9 13 13 2
25 9 1 9 13 4 9 1 13 1 9 13 2 7 9 9 9 14 13 1 1 1 9 14 13 2
13 15 1 9 1 3 2 3 14 13 9 13 4 2
17 9 13 9 1 9 2 9 1 9 13 11 9 1 1 9 13 2
23 9 1 0 9 1 13 16 15 9 11 1 10 3 13 4 15 1 10 9 13 4 4 2
28 9 1 9 7 0 9 1 9 1 13 16 10 9 1 9 9 1 13 4 1 1 1 9 0 13 4 4 2
10 9 9 13 1 3 9 13 4 4 2
14 9 1 3 2 3 9 1 11 9 1 13 4 4 2
13 15 14 12 2 12 9 1 9 9 13 4 4 2
20 9 1 9 2 3 13 13 4 7 9 13 1 3 14 15 3 0 13 4 2
25 9 1 13 13 16 10 9 13 1 9 9 14 13 4 4 7 14 9 2 9 1 14 9 13 2
31 11 11 11 1 11 9 1 0 11 1 9 9 13 1 9 1 11 1 0 9 9 11 11 1 0 13 1 9 13 4 2
30 9 1 9 13 16 10 9 1 11 11 11 2 11 2 3 11 1 9 9 1 13 9 1 9 1 0 13 1 13 2
21 9 1 9 11 11 1 10 9 1 9 1 9 13 4 9 13 1 9 13 4 2
51 11 9 11 11 1 9 9 1 9 1 0 9 1 1 1 13 16 11 1 1 11 1 1 9 13 1 1 10 9 0 13 7 15 12 9 1 11 9 1 9 0 13 1 1 14 3 14 9 0 13 2
23 11 13 4 16 9 1 9 9 1 1 15 15 9 14 13 7 15 9 9 14 13 4 2
5 10 9 15 13 2
8 11 11 11 11 1 9 13 2
9 9 14 10 9 1 9 9 13 2
19 15 10 9 1 9 13 0 13 16 15 9 1 9 1 10 9 13 4 2
16 16 15 13 16 10 9 1 11 14 15 9 1 13 14 4 2
14 16 15 10 9 1 9 14 13 16 10 0 9 13 2
16 7 10 9 0 13 4 16 11 11 1 15 13 1 15 13 2
17 11 1 9 13 16 15 15 9 1 9 13 4 1 0 9 13 2
36 15 13 16 9 1 15 15 14 13 16 15 9 1 0 13 1 9 15 9 13 7 11 1 9 11 1 9 1 15 11 11 1 13 4 4 2
15 11 1 13 16 11 1 10 9 1 0 9 13 13 4 2
11 11 9 9 9 1 9 1 1 9 13 2
19 0 9 9 7 11 9 11 1 0 12 0 9 1 9 13 1 13 4 2
26 11 11 0 10 9 1 9 13 16 15 9 1 0 9 9 1 11 9 1 13 1 9 13 4 4 2
17 12 0 11 11 1 11 1 9 9 11 1 11 0 13 4 4 2
25 11 11 11 0 11 11 11 11 11 1 9 13 1 14 3 11 9 1 15 15 9 1 13 4 2
30 9 9 9 2 9 2 11 11 1 11 1 13 16 11 9 1 9 1 11 9 1 10 0 9 1 9 1 13 4 2
26 11 9 1 13 4 16 11 1 0 9 9 1 0 9 1 13 1 9 1 9 1 0 13 4 4 2
25 16 2 11 1 15 1 1 0 9 13 1 3 15 0 13 4 16 11 1 1 10 9 13 4 2
11 10 9 1 12 7 12 9 13 4 4 2
9 15 1 9 11 1 9 13 4 2
28 10 3 11 9 11 1 1 1 10 10 9 13 1 1 11 9 1 0 9 1 9 13 1 9 13 4 4 2
20 11 1 9 9 1 9 9 1 13 4 4 7 15 15 0 14 13 4 4 2
14 9 9 1 9 0 10 9 1 15 9 13 4 4 2
18 9 9 1 13 16 9 9 0 10 9 1 11 1 9 13 4 4 2
30 9 1 13 4 4 16 15 9 15 9 3 9 11 11 7 9 11 11 13 2 9 1 15 9 9 9 1 0 13 2
30 11 1 12 9 1 13 16 10 10 9 13 1 1 9 9 1 12 9 11 0 11 11 11 11 1 9 13 4 4 2
18 7 9 1 0 15 11 11 7 11 11 0 9 15 1 14 13 4 2
45 3 11 0 10 0 9 1 0 13 1 3 11 1 9 9 9 9 11 11 11 1 11 1 12 9 9 1 13 16 11 1 11 1 9 1 9 1 9 9 13 1 9 13 4 2
9 15 1 15 9 13 4 4 4 2
13 3 1 15 11 0 10 9 1 14 9 13 4 2
21 16 2 9 1 10 9 13 4 4 16 15 1 15 9 9 7 0 9 14 13 2
21 15 1 15 11 0 13 1 9 13 4 2 15 11 11 15 1 0 9 13 4 2
16 9 1 0 9 1 0 9 1 12 9 1 15 9 13 4 2
24 9 7 9 1 10 9 1 10 9 2 15 13 7 15 14 13 2 1 0 9 13 4 4 2
13 9 1 14 0 9 1 9 9 13 4 4 4 2
23 0 9 7 9 2 9 1 9 14 13 2 15 1 9 14 13 2 1 10 9 13 4 2
36 0 9 1 0 9 1 9 2 9 7 9 9 1 9 1 9 0 14 13 7 9 1 9 0 13 4 4 16 9 15 0 9 14 13 4 2
16 9 1 1 10 9 14 0 9 1 15 9 1 14 9 13 2
31 12 9 1 9 1 9 11 11 1 13 13 16 9 10 9 13 15 10 9 1 10 9 13 16 15 9 9 13 9 13 2
7 15 9 1 13 4 4 2
17 0 9 9 11 11 1 13 13 16 9 1 1 9 9 0 13 2
10 7 15 0 9 1 9 13 4 4 2
12 9 1 15 9 1 9 9 9 13 4 4 2
18 7 15 0 9 2 9 7 9 15 15 13 4 15 15 9 13 4 2
27 16 11 11 11 1 9 9 11 11 1 13 16 0 9 2 9 1 10 9 1 9 9 1 13 4 4 2
21 15 15 15 14 9 1 9 14 13 7 15 14 9 14 13 1 9 13 4 4 2
18 9 1 1 14 9 1 1 9 7 9 0 9 1 9 13 4 4 2
32 9 1 13 4 4 4 16 15 1 10 9 0 13 1 15 15 1 13 4 2 7 3 9 13 7 9 1 9 13 4 14 2
31 11 11 1 0 9 3 14 0 13 15 9 13 1 9 1 13 11 11 11 11 11 11 0 9 11 1 9 13 4 4 2
51 15 0 9 7 0 11 11 11 11 11 11 11 1 11 1 0 9 13 14 12 0 9 1 13 1 3 11 11 1 9 15 9 1 0 9 1 1 1 15 1 9 7 0 0 9 1 9 13 1 13 2
24 11 11 11 11 1 0 9 13 1 0 9 9 1 0 9 1 0 13 1 9 13 4 4 2
24 7 11 11 1 0 9 13 1 9 1 15 0 9 1 9 15 13 2 15 15 0 14 13 2
15 15 1 1 9 9 13 1 1 11 11 11 13 4 4 2
30 15 9 1 0 9 1 0 13 1 13 11 11 1 0 9 15 11 11 1 0 9 13 1 9 1 9 1 13 4 2
31 11 11 1 11 11 11 11 13 1 14 3 14 11 11 1 9 11 11 1 9 1 9 1 12 9 1 15 9 13 4 2
44 11 11 1 10 9 1 10 9 13 4 16 15 15 9 2 11 11 14 11 11 1 9 13 4 2 1 0 9 3 13 7 10 9 1 3 14 9 13 1 9 14 13 4 2
25 16 15 3 1 13 4 4 16 9 1 9 3 2 3 15 13 15 11 1 9 1 0 13 4 2
22 10 9 1 9 13 1 9 1 11 11 11 2 11 11 1 11 9 1 13 4 4 2
18 10 3 15 11 1 9 11 11 1 1 14 9 2 9 13 4 4 2
38 16 9 9 1 0 9 1 13 16 11 11 1 9 0 9 1 9 1 1 2 9 0 9 1 9 1 9 11 11 1 1 0 9 2 9 13 4 2
18 15 11 11 11 11 1 9 11 11 11 7 0 9 1 14 13 14 2
11 9 1 9 1 1 14 9 2 9 13 2
17 15 10 9 1 9 7 9 1 9 9 1 1 14 9 13 4 2
18 0 11 11 11 11 1 9 1 11 11 11 1 9 1 13 4 4 2
23 3 11 1 0 9 11 11 1 11 7 11 11 1 9 1 9 13 4 1 9 13 4 2
31 3 11 1 9 11 11 1 13 16 11 1 11 9 1 1 11 11 1 11 9 1 13 1 9 13 3 0 9 13 4 2
31 15 11 1 10 9 1 9 13 4 13 16 15 9 1 9 12 0 9 1 1 13 4 15 15 9 12 1 11 1 13 2
8 15 11 15 9 13 4 4 2
27 15 13 16 11 7 11 9 14 0 9 1 13 4 4 16 10 9 1 14 11 1 14 1 13 4 4 2
19 10 15 9 15 13 16 11 1 1 10 0 0 9 13 15 14 3 13 4
29 11 1 10 9 11 1 11 1 13 10 9 1 13 4 15 11 1 9 1 1 11 1 9 1 0 13 4 4 2
27 11 1 10 9 1 14 0 9 13 16 11 1 10 9 11 11 1 11 1 9 1 1 0 13 4 4 2
7 3 10 9 1 11 15 13
26 11 1 9 1 2 9 15 13 16 11 7 11 9 14 0 13 4 7 9 9 1 9 14 13 13 2
24 15 0 15 13 16 15 9 1 9 13 4 7 9 1 1 15 10 9 13 4 15 9 13 2
12 15 9 1 9 11 1 9 1 9 13 13 4
18 11 7 11 1 15 11 1 9 9 1 9 1 14 13 4 13 4 2
6 2 15 15 9 13 2
8 15 9 9 1 13 4 4 2
8 9 1 9 9 14 13 4 2
7 15 15 9 15 13 14 4
11 15 11 1 13 1 9 1 13 4 4 2
22 15 13 16 15 3 0 13 16 11 9 1 11 9 9 13 7 15 11 11 13 4 2
24 15 13 16 11 1 15 9 7 11 11 9 1 13 4 15 15 0 9 1 11 1 9 13 2
26 15 13 16 15 0 9 1 9 12 0 9 1 14 1 13 4 15 15 0 9 1 0 9 1 13 2
22 15 13 16 15 1 14 9 9 1 0 14 13 7 15 11 1 14 1 13 4 4 2
29 11 11 11 9 11 11 11 1 9 1 9 9 1 9 13 1 13 11 1 9 13 1 12 10 9 13 4 4 2
12 11 1 11 1 10 9 1 0 9 13 4 2
27 9 1 13 13 16 9 9 1 0 9 7 9 1 10 9 1 9 13 1 15 0 7 0 9 14 13 2
21 9 1 0 0 9 13 4 11 1 13 4 16 15 0 9 1 15 9 14 13 2
28 11 9 1 9 1 13 1 9 13 4 11 1 13 4 16 0 0 9 1 3 1 9 14 14 13 4 4 2
9 15 9 1 1 9 1 9 13 2
16 11 1 13 13 16 9 1 0 9 7 9 1 0 9 13 2
13 10 9 7 9 1 10 9 1 0 9 13 4 2
17 15 10 9 0 13 4 16 9 1 0 9 1 15 9 14 13 2
15 15 13 16 9 1 0 9 13 1 9 0 9 0 13 2
17 9 9 2 9 1 9 1 9 9 1 15 9 0 13 4 4 2
24 11 1 9 1 11 11 11 2 11 2 9 1 1 9 10 9 9 1 0 9 13 4 4 2
14 11 0 9 1 9 15 14 9 9 13 9 13 4 2
10 16 15 9 9 9 14 0 13 4 2
15 15 13 16 0 9 1 9 1 9 1 15 9 14 13 2
27 11 1 9 13 4 9 9 1 13 16 9 9 7 9 9 1 13 0 9 15 9 13 1 0 13 4 2
21 9 1 9 1 1 9 7 15 1 0 9 1 1 0 9 14 13 4 4 4 2
18 15 9 1 13 9 13 7 15 1 9 13 1 0 9 0 13 4 2
18 11 11 11 9 1 0 9 13 1 1 12 0 9 13 4 4 4 2
15 0 0 10 9 1 15 13 1 1 9 9 0 13 4 2
11 15 1 9 9 15 0 9 1 0 13 2
17 9 13 1 9 1 9 1 1 9 1 9 9 14 0 13 4 2
24 9 1 9 1 0 9 1 0 9 7 9 9 1 11 1 15 13 9 1 15 0 13 4 2
11 9 1 11 11 1 10 0 9 0 13 2
24 11 11 1 9 1 9 1 9 1 1 11 1 13 4 9 1 9 1 9 13 1 13 4 2
21 9 1 1 9 9 11 11 11 1 13 16 11 11 1 0 9 9 1 9 13 2
25 15 13 16 9 1 15 0 9 1 10 0 13 7 0 9 1 9 2 9 13 1 13 4 4 2
27 15 13 16 13 9 0 9 1 9 13 2 7 15 15 14 13 16 10 9 10 9 1 9 1 13 4 2
30 11 11 1 9 1 13 16 9 1 13 1 1 11 1 0 9 1 0 7 0 9 1 9 1 9 1 9 13 4 2
14 11 10 9 1 13 1 1 9 1 10 0 9 13 2
18 10 9 1 11 11 11 2 11 7 11 9 1 9 14 13 4 4 2
15 16 15 1 1 1 0 9 1 0 9 9 13 4 4 2
18 9 1 0 0 9 9 1 9 11 1 1 14 0 13 1 9 13 2
18 10 9 1 1 14 9 1 10 9 12 2 12 12 9 13 4 4 2
13 11 1 13 16 9 10 9 1 9 1 13 4 2
16 15 14 0 13 16 9 12 2 12 11 11 9 1 9 13 2
10 11 10 9 1 1 12 12 9 13 2
10 9 1 9 1 0 9 14 13 4 2
24 9 9 1 12 9 1 9 1 13 16 11 1 9 1 1 9 1 9 9 12 0 9 13 2
25 15 11 1 9 13 14 13 16 10 0 9 1 9 1 13 16 10 9 9 1 9 1 14 13 2
13 16 2 9 10 9 1 13 1 9 1 9 13 2
35 9 1 11 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 11 2 11 2 11 11 2 11 2 11 7 11 1 9 0 13 2
12 10 9 1 9 1 11 11 9 13 4 4 2
5 15 0 9 13 2
17 15 1 11 1 9 1 13 9 1 9 1 14 9 9 13 4 2
21 11 11 9 1 1 14 11 1 12 9 7 12 9 9 1 1 9 0 13 4 2
18 11 11 1 12 9 1 1 9 0 9 1 1 3 0 9 1 13 2
26 11 11 1 11 9 9 1 0 9 1 12 9 13 4 7 11 9 9 1 12 9 9 1 9 13 2
6 9 11 11 1 13 2
7 0 9 9 1 13 4 2
20 16 11 1 9 0 9 1 9 13 7 9 13 14 9 1 9 0 13 4 2
14 11 11 1 1 9 1 12 2 12 9 1 9 13 2
22 9 1 9 9 9 11 11 11 11 1 14 12 9 1 10 9 13 1 9 13 4 2
27 9 1 12 9 1 13 12 12 1 10 9 9 1 9 12 12 9 1 9 12 12 9 1 9 13 4 2
19 16 9 1 9 1 9 9 1 9 13 4 2 7 15 0 9 14 13 2
19 9 1 1 11 1 11 1 12 0 2 0 9 1 12 9 0 13 4 2
20 9 1 11 9 1 9 9 13 4 9 9 1 9 1 3 9 9 13 4 2
6 15 15 0 14 13 2
8 0 9 1 1 9 13 4 2
25 12 0 9 1 11 1 9 1 7 11 1 9 1 9 1 0 9 7 9 9 1 9 13 4 2
25 15 11 1 11 11 11 7 11 1 11 11 0 13 4 2 15 11 1 9 1 0 13 4 4 2
15 16 2 11 11 1 9 1 13 9 1 12 9 13 4 2
27 11 11 11 11 1 9 13 1 0 13 11 9 9 1 9 14 12 12 9 0 9 1 12 9 13 4 2
8 12 9 1 0 13 4 4 2
22 12 9 1 9 9 1 12 9 1 9 1 9 13 1 9 14 11 11 1 13 4 2
10 10 9 9 1 0 13 4 4 4 2
14 15 9 1 9 9 9 1 0 9 13 1 3 13 2
32 9 1 9 1 12 9 7 9 1 10 12 9 1 1 13 9 1 0 9 1 1 14 12 2 12 9 9 9 1 3 13 2
21 11 2 11 1 9 1 12 9 1 1 13 9 1 15 0 16 15 0 9 13 2
14 11 1 0 9 1 1 14 12 9 9 9 13 13 2
17 15 1 9 1 11 11 11 11 9 1 13 1 9 13 4 4 2
9 11 9 9 1 12 9 9 13 2
18 16 11 7 11 9 9 1 12 2 12 9 9 13 1 9 13 4 2
16 11 1 11 9 9 1 1 13 9 1 14 12 9 9 13 2
15 11 1 11 9 9 1 9 9 12 9 13 1 9 13 2
23 9 1 3 10 12 9 9 11 1 12 7 11 1 12 9 9 1 1 13 9 1 13 2
26 11 1 12 9 9 1 1 13 9 1 9 1 9 14 13 7 14 12 9 9 14 9 1 3 13 2
21 11 1 9 9 1 9 7 12 9 1 0 9 1 1 0 9 0 9 0 13 2
20 9 1 9 1 1 9 1 12 9 9 1 13 9 0 9 1 0 13 4 2
38 0 9 1 11 11 1 12 2 12 9 2 11 1 12 9 2 11 1 12 9 2 11 1 12 2 12 9 7 11 1 12 9 9 13 1 9 13 2
23 11 1 0 9 11 11 1 11 11 1 11 9 1 9 3 13 4 1 15 9 14 13 2
16 9 14 15 13 16 9 9 11 11 11 1 9 1 0 13 2
9 11 1 9 1 14 9 0 13 2
22 15 9 9 1 9 11 11 1 13 4 9 1 15 9 0 13 1 9 1 14 13 2
17 11 9 11 11 11 1 9 13 4 1 9 1 9 13 4 4 2
41 7 9 1 0 9 11 11 1 0 9 1 9 13 4 1 9 1 14 15 0 13 4 16 9 1 11 11 1 3 9 1 9 13 4 1 9 14 13 4 4 2
26 11 1 12 9 1 12 9 1 11 1 9 1 9 13 4 1 3 15 11 9 1 9 13 4 4 2
25 9 1 9 1 13 13 16 10 9 14 0 13 4 4 16 11 9 1 15 9 1 9 13 4 2
22 3 9 7 0 9 1 11 15 9 13 1 0 13 4 16 15 11 1 0 11 13 2
17 15 1 14 11 1 11 1 11 9 1 14 0 9 13 4 4 2
21 9 9 1 13 13 16 16 11 11 11 13 16 3 14 11 1 0 9 13 4 2
18 11 1 0 9 15 13 16 15 9 7 9 1 1 0 9 13 4 2
27 15 0 9 1 9 9 14 13 4 7 9 2 9 1 1 13 4 1 9 1 9 1 0 9 13 4 2
13 11 9 1 9 1 14 15 15 9 13 4 4 2
33 7 11 11 1 9 1 9 1 9 1 11 1 9 1 9 13 1 9 15 9 1 13 4 2 15 1 9 1 9 1 9 13 2
18 9 9 1 1 10 15 9 14 13 4 16 10 9 1 9 13 4 2
16 15 15 0 13 4 16 3 15 9 9 1 15 9 14 13 2
28 15 2 15 11 9 15 3 13 1 9 13 4 4 16 9 1 10 9 0 13 4 1 3 3 15 9 13 2
21 9 11 1 11 9 0 9 1 9 13 0 9 13 4 1 9 9 1 13 4 2
9 9 0 9 1 12 9 1 13 2
11 9 1 9 0 13 9 9 13 4 4 2
10 15 1 15 1 9 14 13 4 4 2
20 9 1 9 9 1 13 7 15 11 1 14 9 13 1 3 9 1 13 4 2
34 9 1 0 9 1 9 1 13 4 9 1 1 15 9 11 2 0 9 2 11 2 11 11 1 9 1 0 15 9 1 13 4 4 2
16 15 12 9 15 13 15 1 10 3 0 12 9 1 13 4 2
8 15 9 1 15 1 9 13 2
18 9 13 1 15 9 1 9 14 13 2 15 3 1 15 9 13 4 2
13 9 1 1 9 9 1 1 9 1 9 1 13 2
12 9 1 12 9 1 1 9 0 13 4 4 2
8 9 1 0 9 13 4 4 2
26 11 1 11 11 11 9 15 9 1 9 1 9 1 13 4 0 9 7 9 1 1 0 13 13 4 2
21 11 11 11 11 11 1 13 4 16 9 1 10 12 9 1 12 9 8 13 4 2
10 15 9 1 14 15 9 1 9 13 2
11 0 9 1 12 9 14 9 13 4 4 2
13 9 1 9 1 1 11 11 11 1 9 13 4 2
25 9 11 1 13 16 11 1 9 1 10 9 1 10 9 1 9 13 16 11 1 15 14 13 4 2
13 15 1 15 9 1 9 9 1 9 1 9 13 2
21 10 12 9 1 13 1 10 9 11 11 11 2 11 11 11 2 1 9 1 13 2
10 10 9 1 9 1 0 9 13 4 2
15 11 11 1 15 1 1 9 9 1 10 9 1 9 13 2
16 10 9 15 0 13 4 4 2 16 15 15 0 13 4 4 2
26 9 11 1 15 9 1 13 4 16 9 1 15 9 1 9 1 1 10 12 9 1 9 9 13 4 2
15 9 9 1 9 1 10 9 10 14 10 9 13 4 4 2
17 0 2 0 9 1 9 13 1 14 9 1 9 0 13 4 4 2
30 11 11 11 1 11 11 1 9 9 11 11 11 1 9 11 1 9 1 9 0 13 4 13 16 15 14 0 9 13 2
13 9 1 15 9 1 1 1 9 14 13 14 4 2
10 15 9 1 9 1 13 4 9 13 2
13 9 1 10 14 9 1 9 1 9 13 4 4 2
17 11 1 9 1 14 12 9 1 9 12 9 1 0 14 13 4 2
19 7 11 1 12 9 1 9 13 9 1 15 9 1 9 9 13 4 4 2
14 9 1 1 0 9 13 1 15 9 14 13 14 4 2
31 11 11 11 1 9 9 11 11 1 13 13 16 10 9 1 9 0 9 14 9 11 1 13 4 2 7 0 14 13 4 2
22 9 9 14 0 9 1 13 4 2 7 11 1 9 1 10 9 14 0 13 14 14 2
27 15 13 10 9 14 0 13 16 9 1 10 9 1 1 9 13 4 4 4 2 15 15 9 14 13 4 2
9 7 9 1 14 10 9 13 4 2
43 11 11 11 1 9 9 11 11 11 1 13 13 16 15 12 11 11 11 1 9 1 3 2 3 9 14 13 4 4 2 15 9 1 3 2 3 9 13 1 10 9 13 2
16 9 9 0 9 11 1 0 9 9 2 11 2 1 9 13 2
19 10 9 1 9 9 1 9 0 9 1 13 4 15 15 9 10 13 4 2
30 11 11 1 9 11 11 1 11 1 13 16 12 0 0 9 1 11 11 11 11 11 2 11 2 1 9 0 13 4 2
13 9 9 10 9 1 11 11 1 13 1 13 4 2
15 15 13 16 9 9 1 13 1 9 9 13 4 4 4 2
13 15 0 13 1 9 12 0 9 1 13 4 4 2
10 15 13 16 15 0 9 13 4 4 2
21 12 9 1 1 10 9 10 0 9 9 9 1 0 11 1 0 13 1 0 13 2
26 15 13 16 10 9 1 0 13 4 1 3 11 10 9 1 9 1 0 13 4 15 1 0 9 13 2
14 3 11 7 11 10 12 9 13 15 1 10 9 13 2
33 11 0 9 1 9 13 1 2 11 11 11 11 2 11 2 9 13 15 12 9 1 0 9 7 11 11 11 2 11 2 13 4 2
39 9 11 1 0 9 9 1 0 9 11 11 11 11 11 1 9 1 11 11 11 11 11 1 9 1 1 11 1 11 1 0 0 9 1 0 13 4 4 2
20 11 1 0 9 12 9 13 7 15 0 7 9 9 1 13 4 1 0 13 2
35 9 2 9 9 1 9 1 9 1 9 13 4 11 1 13 16 9 1 9 1 13 1 1 11 11 11 11 0 9 1 9 13 4 4 2
15 15 13 16 9 1 9 1 1 10 0 9 14 13 4 2
34 15 1 9 1 9 1 13 1 1 10 9 1 0 13 4 7 15 1 15 0 9 1 9 13 4 15 1 15 15 9 13 4 4 2
26 11 11 13 1 10 9 1 11 11 1 11 1 9 1 0 9 1 9 1 9 1 13 3 9 13 2
21 15 12 9 1 11 1 9 13 16 11 11 1 9 7 15 1 12 1 9 13 2
12 16 10 9 1 15 15 9 1 9 14 13 2
21 11 1 10 9 11 1 11 11 1 13 4 11 11 11 11 11 13 4 4 4 2
18 15 0 9 13 4 9 1 13 11 1 13 16 9 1 10 9 13 2
20 15 1 0 11 9 9 9 1 13 12 9 1 9 14 13 9 14 13 4 2
40 10 9 1 9 1 9 9 2 0 9 2 11 11 1 0 9 1 9 13 4 11 1 13 16 11 11 1 12 11 9 1 13 1 3 15 9 1 13 4 2
53 11 11 7 0 9 1 9 9 1 0 9 1 0 9 1 9 1 9 13 4 11 11 11 1 13 16 15 1 1 0 9 1 9 9 1 9 7 9 1 9 1 1 0 11 11 11 1 0 13 15 9 13 2
22 15 13 16 13 4 0 2 0 9 1 11 11 7 11 11 1 0 9 13 0 13 2
33 11 11 1 11 11 11 11 11 11 1 0 13 9 1 9 13 4 11 11 1 9 9 13 11 11 1 0 13 4 1 9 13 2
24 9 9 1 1 11 9 1 0 9 13 1 12 9 1 9 1 0 13 4 1 9 13 4 2
15 11 1 9 9 1 0 13 1 9 1 9 0 13 4 2
14 12 12 9 1 1 14 12 12 9 1 9 13 4 2
18 9 1 13 16 11 11 1 9 9 13 11 11 1 0 13 4 4 2
29 9 1 9 1 10 9 9 13 4 16 16 0 9 1 1 15 9 7 9 13 4 16 15 14 0 13 4 4 2
10 9 1 11 11 11 1 9 0 13 2
17 11 9 11 1 0 9 1 1 15 9 1 11 1 3 9 13 2
10 13 1 1 12 9 9 14 0 13 2
14 11 11 1 9 11 1 0 9 9 1 0 13 4 2
10 15 9 9 0 0 9 1 13 4 2
16 15 1 11 1 0 9 9 1 3 11 11 1 13 4 4 2
15 10 3 15 13 15 9 0 13 4 7 9 9 13 4 2
18 15 9 1 3 7 3 0 9 1 9 13 7 9 1 14 9 13 2
14 9 1 11 1 11 11 11 11 11 1 14 14 13 2
20 15 1 11 1 0 9 11 14 13 2 7 15 10 9 1 3 3 13 4 2
14 11 9 1 9 12 9 1 0 9 1 0 9 13 2
17 11 9 11 11 1 15 9 1 0 9 13 4 15 0 9 13 2
13 9 1 13 16 3 10 0 9 11 11 1 13 2
30 9 7 9 9 1 9 13 1 1 15 9 9 1 14 13 15 9 1 9 13 4 2 15 12 9 1 9 13 4 2
15 7 12 0 9 9 9 9 1 1 13 9 1 13 4 2
23 0 9 1 1 1 15 9 14 13 4 4 16 15 9 1 7 9 1 9 1 13 4 2
15 13 9 1 12 0 9 13 4 7 10 9 1 9 13 2
15 15 9 1 3 7 3 0 9 1 9 1 14 9 13 2
33 11 11 1 11 1 9 9 13 4 1 3 15 1 13 9 1 0 2 0 13 1 1 9 1 10 9 9 9 1 9 13 4 2
21 9 1 13 1 1 0 12 9 1 9 1 9 13 7 15 1 9 9 13 4 2
32 11 1 0 9 1 1 15 9 11 11 2 11 11 7 11 11 1 11 11 13 1 10 9 1 12 9 9 9 1 13 4 2
19 9 13 13 11 1 9 11 11 1 0 9 9 1 9 1 13 4 4 2
20 15 1 11 11 1 13 4 14 12 9 0 9 9 1 9 1 3 9 13 2
18 10 9 1 9 13 4 7 10 9 9 1 10 9 1 9 13 4 2
15 9 9 1 12 0 9 7 12 9 1 9 13 4 4 2
18 11 9 11 11 1 9 1 12 9 13 1 3 11 1 9 13 4 2
29 12 0 9 1 11 1 12 12 9 1 0 9 7 12 2 12 12 1 12 9 1 9 1 0 13 1 9 13 2
33 9 13 1 3 14 11 1 9 1 14 9 1 9 2 9 13 7 9 1 1 0 13 1 3 9 9 11 11 11 1 9 13 2
34 10 9 1 11 1 14 9 1 1 9 13 4 9 9 1 15 9 14 13 2 7 15 9 11 1 11 11 11 1 9 3 0 13 2
23 11 7 11 1 9 11 11 1 15 9 1 3 9 1 1 9 13 11 0 9 13 4 2
10 11 11 1 13 16 15 3 0 13 2
13 11 1 13 16 15 0 9 1 1 0 9 13 2
17 15 13 16 15 9 1 14 11 1 9 1 9 13 4 4 4 2
34 15 1 11 1 9 9 9 9 11 11 11 1 9 13 4 1 9 13 14 9 1 1 9 1 14 13 9 1 9 1 9 13 4 2
19 9 1 9 1 0 13 1 1 0 9 13 4 7 0 9 14 13 4 2
38 11 11 1 11 1 13 1 1 12 9 9 13 1 9 13 4 12 0 9 1 9 1 9 1 9 7 9 9 1 0 9 1 1 9 1 9 13 2
9 10 9 11 9 1 0 14 13 2
23 7 15 1 11 9 1 12 0 9 1 9 13 1 9 1 9 9 1 1 0 13 4 2
15 9 1 10 9 1 11 1 12 9 1 9 13 4 4 2
31 11 1 9 1 0 9 0 13 1 1 11 11 11 1 9 1 3 0 9 11 1 9 10 9 1 1 0 13 4 4 2
23 11 0 9 9 1 9 12 12 9 1 1 12 12 9 1 9 9 0 13 4 4 4 2
24 15 1 14 15 9 1 9 10 13 4 15 11 11 11 11 11 1 1 1 9 13 4 4 2
27 15 1 0 13 4 9 9 1 1 14 12 12 9 15 9 1 9 1 11 11 11 1 9 13 4 4 2
22 11 1 9 0 13 4 1 9 13 14 11 1 9 12 12 9 9 1 13 4 4 2
21 9 1 1 0 9 7 9 13 4 11 1 1 11 1 14 12 9 13 4 4 2
11 10 9 13 14 9 1 9 3 9 13 2
16 11 1 9 12 9 1 9 1 9 12 12 9 13 4 4 2
21 0 9 1 1 10 9 15 1 10 9 12 12 1 9 1 13 4 1 9 13 2
24 9 9 1 9 11 11 1 1 9 1 9 1 10 9 15 10 9 1 0 13 1 9 13 2
23 0 13 16 0 11 1 14 9 10 9 1 0 13 4 1 3 9 3 9 13 4 4 2
34 0 9 1 11 1 9 2 9 9 9 1 1 13 1 9 9 1 9 1 1 9 11 11 1 0 9 1 3 13 1 9 13 4 2
14 10 9 1 11 11 1 9 11 11 9 13 4 4 2
33 10 9 11 1 9 7 0 9 11 11 1 9 13 4 1 1 10 9 0 13 4 4 2 15 1 9 9 13 0 13 4 4 2
30 11 15 9 1 11 1 11 1 13 0 9 9 1 9 1 11 7 11 11 1 9 1 1 1 9 0 13 13 4 2
15 11 1 15 9 9 1 10 9 1 13 1 9 13 4 2
23 3 11 9 1 1 9 13 4 7 13 4 4 16 15 11 11 1 9 9 1 9 13 2
29 13 4 4 4 16 10 3 15 15 0 9 1 9 1 11 2 11 11 1 9 9 1 12 9 1 14 9 13 2
26 11 1 11 9 11 11 1 9 1 13 16 16 11 11 1 9 9 1 9 13 16 15 3 9 13 2
33 9 1 10 9 1 0 9 13 16 15 11 11 1 15 13 16 9 9 1 15 10 9 13 2 15 3 10 0 9 13 4 4 2
20 15 13 16 9 9 9 1 9 1 1 11 11 1 1 9 1 9 13 4 2
14 16 2 11 9 10 9 1 15 15 14 13 4 4 2
13 9 9 1 11 11 1 9 13 1 9 13 4 2
21 11 1 12 9 1 13 16 0 13 16 10 9 1 15 11 1 3 9 14 13 2
12 7 9 9 15 10 9 1 9 13 14 4 2
19 11 11 1 11 1 9 9 1 11 9 13 1 9 1 9 0 13 4 2
25 15 1 14 11 11 1 9 9 11 11 1 9 1 9 0 13 1 1 12 12 9 9 14 13 2
18 9 9 11 11 11 7 9 11 11 11 1 9 1 9 0 13 4 2
21 10 9 1 11 1 11 11 11 0 11 11 11 1 11 9 13 1 9 13 4 2
14 9 1 9 13 16 11 11 1 12 9 1 9 13 2
18 15 0 9 9 1 15 9 1 0 13 1 0 9 0 13 4 4 2
15 11 1 11 9 1 9 1 1 1 11 1 9 13 4 2
34 11 11 11 11 1 1 1 0 0 0 9 11 11 1 13 16 10 9 0 7 0 0 9 1 13 4 2 15 11 1 9 1 13 2
22 15 13 16 9 9 1 1 9 1 0 9 1 14 13 7 13 1 9 0 13 4 2
33 15 1 11 11 1 9 1 11 11 1 11 1 9 0 13 4 7 0 9 1 9 13 1 3 11 11 1 15 9 0 13 4 2
37 11 11 1 11 11 11 11 11 1 12 0 9 1 0 13 1 9 1 9 13 4 4 2 15 1 0 9 1 9 9 0 13 1 9 13 4 2
24 11 11 11 1 9 1 11 1 13 9 1 9 1 12 12 9 1 10 9 1 9 13 4 2
25 13 4 4 16 0 9 1 9 13 1 1 12 12 9 1 9 1 9 1 9 14 13 4 4 2
14 7 11 1 12 12 1 9 1 0 13 4 4 4 2
22 9 1 1 9 1 11 11 1 11 1 1 12 0 9 1 9 1 9 13 4 4 2
13 0 9 9 1 9 1 9 2 9 14 13 4 2
9 10 9 1 3 13 4 4 4 2
20 9 7 9 9 1 9 13 1 1 15 9 1 0 3 9 1 0 13 4 2
17 15 1 9 9 9 1 9 1 9 2 11 2 1 14 9 13 2
30 15 11 11 11 2 11 7 11 1 9 1 9 1 13 4 11 2 11 9 1 9 13 7 9 9 9 1 9 13 2
21 2 11 11 11 11 11 2 1 1 11 11 1 0 9 1 14 0 13 4 4 2
21 15 1 11 2 11 2 11 2 11 7 11 11 1 9 1 14 0 13 4 4 2
51 16 9 1 11 9 1 13 4 15 0 9 14 13 7 0 9 1 1 2 11 11 11 11 2 1 1 10 0 9 1 10 9 1 9 13 4 15 11 11 7 11 11 1 9 1 14 9 13 4 4 2
17 13 4 4 16 11 11 1 9 1 11 10 0 9 13 4 4 2
25 11 1 9 1 9 9 1 9 9 1 9 1 13 4 9 1 13 4 11 11 11 1 9 13 2
25 9 1 13 16 11 11 1 10 9 1 14 2 0 9 2 9 1 9 1 9 1 9 13 4 2
15 11 11 1 1 9 1 0 9 1 15 9 14 13 4 2
20 9 1 11 11 11 11 2 11 11 11 11 7 11 11 11 11 14 0 13 2
26 9 9 1 11 2 11 1 9 1 11 2 11 9 1 12 9 1 1 9 13 1 9 1 9 13 2
18 11 2 11 1 12 9 0 9 1 1 12 9 1 9 1 9 13 2
11 11 1 10 9 1 11 9 13 4 4 2
16 11 7 11 1 1 11 1 0 9 1 0 9 1 9 13 2
17 12 9 1 1 9 2 9 7 9 1 12 9 1 9 13 4 2
22 9 1 9 13 4 1 3 11 1 11 11 11 7 11 1 11 11 11 11 0 13 2
19 15 1 12 9 1 0 9 1 0 2 0 7 0 9 1 9 9 13 2
23 11 1 11 11 11 11 7 0 11 11 11 1 9 1 1 0 9 1 13 1 9 13 2
13 10 12 9 1 1 11 1 11 11 1 9 13 2
10 11 1 15 11 9 1 0 13 4 2
18 0 13 16 12 9 1 1 11 1 15 11 1 15 0 11 9 13 2
22 11 1 9 1 13 16 9 1 1 15 11 1 0 9 1 1 9 13 1 9 13 2
15 11 1 14 11 11 1 11 1 0 9 1 9 13 4 2
15 10 9 1 11 11 7 15 9 1 0 9 14 0 13 2
17 12 9 1 9 1 1 0 9 1 11 1 9 9 9 13 4 2
21 11 1 1 15 9 11 2 11 1 0 9 7 9 1 12 9 11 13 4 4 2
18 10 9 1 11 1 11 11 11 11 11 7 11 11 11 11 0 13 2
12 11 1 11 11 2 11 11 11 1 9 13 2
26 9 1 9 11 11 11 2 11 2 2 11 7 11 1 12 0 9 1 0 9 1 13 4 4 4 2
18 10 9 1 11 7 11 1 14 12 9 1 9 9 9 13 4 4 2
22 9 1 11 9 15 9 1 9 13 1 3 11 9 1 9 1 9 0 13 4 4 2
25 15 9 1 9 9 1 9 13 7 9 1 9 8 13 1 9 13 4 9 1 13 4 1 13 2
10 0 13 4 16 9 1 9 13 4 2
26 9 1 9 1 0 9 9 1 13 7 9 13 14 12 9 1 9 9 1 0 9 1 13 13 4 2
32 9 1 10 9 9 1 0 15 9 1 1 1 9 13 1 9 13 4 4 7 9 1 9 1 1 9 9 1 13 4 4 2
27 9 1 0 9 11 11 1 0 9 13 2 15 9 9 1 9 1 14 0 14 13 2 15 15 13 9 2
18 11 9 1 12 9 1 13 16 10 9 0 9 1 9 13 4 4 2
25 11 1 13 16 10 9 9 9 13 4 4 7 3 9 7 9 1 9 1 9 1 9 13 4 2
34 12 0 9 11 1 13 16 2 11 0 2 9 1 3 12 9 1 9 1 13 4 7 3 10 9 1 9 13 9 1 13 1 13 2
27 12 9 9 1 9 13 13 4 4 9 1 1 0 9 8 13 4 4 4 2 15 14 13 14 4 4 2
9 0 13 14 9 1 9 13 4 2
15 9 9 1 0 9 1 1 13 7 9 1 0 13 4 2
28 11 1 1 2 15 1 9 1 0 13 9 1 0 11 1 1 1 9 13 7 15 9 1 13 9 13 4 2
13 9 0 2 0 7 0 0 9 14 13 4 4 2
21 11 1 10 9 1 1 9 13 16 15 9 1 13 16 15 9 1 9 13 4 2
18 16 15 13 13 2 16 15 15 13 4 16 15 9 1 15 13 4 2
22 3 14 15 15 9 1 1 13 2 16 13 16 0 9 13 10 9 9 13 4 4 2
13 10 9 1 15 15 9 1 1 14 13 1 13 2
20 9 9 7 9 1 1 9 9 9 1 13 1 11 15 9 13 3 13 4 2
6 7 2 15 9 13 2
31 11 1 9 1 9 13 4 11 11 11 11 11 2 11 2 1 9 9 1 12 9 1 11 1 9 9 1 9 13 4 2
23 10 9 1 0 9 1 11 11 11 11 11 1 11 9 1 9 1 9 13 4 4 4 2
21 11 1 13 4 16 9 1 9 1 9 1 9 9 1 1 9 13 4 4 4 2
25 11 1 1 10 12 9 11 1 11 1 11 11 9 1 0 9 9 1 9 1 9 13 4 4 2
16 15 9 9 0 13 1 1 11 1 11 1 12 10 9 13 2
17 15 0 9 1 12 9 9 9 13 1 1 0 0 9 9 13 2
29 11 1 0 9 11 1 13 13 16 10 9 1 10 9 15 1 0 9 1 9 13 4 4 15 10 9 1 13 2
32 11 1 9 1 1 12 9 0 9 1 9 1 0 9 2 7 14 12 9 2 12 9 9 9 7 12 9 9 9 13 4 2
10 15 1 15 12 9 1 9 9 13 2
36 16 0 9 15 9 13 4 15 10 9 14 12 9 13 4 7 0 9 1 12 9 9 1 13 4 2 7 15 1 9 9 12 9 1 13 2
21 10 9 1 10 0 9 9 12 9 14 9 7 11 9 9 12 9 14 9 13 2
17 15 10 9 13 15 11 15 9 9 9 1 9 1 13 4 4 2
18 10 9 1 15 9 2 9 13 1 1 9 1 9 2 9 14 13 2
12 10 9 12 0 7 0 0 9 1 1 13 2
18 11 1 0 9 13 14 15 15 0 9 1 10 9 1 13 4 4 2
36 11 11 11 11 1 0 9 1 13 1 0 0 9 11 11 1 15 1 11 9 11 11 11 1 0 13 4 15 9 1 13 1 9 13 4 2
30 11 1 11 1 11 1 9 13 4 15 1 13 9 12 9 1 0 13 7 9 1 9 1 1 0 13 1 13 4 2
12 9 1 13 16 11 3 0 7 0 9 13 2
19 9 1 10 9 1 15 15 0 9 13 1 9 1 1 1 13 4 4 2
23 0 13 16 11 1 11 1 9 1 13 15 9 11 11 1 9 9 1 9 13 4 4 2
48 9 1 13 4 1 12 9 1 11 1 11 1 15 9 1 13 16 11 1 9 2 11 11 2 1 11 1 15 1 0 9 1 9 1 9 13 7 9 1 9 1 0 13 1 9 13 4 2
11 11 1 13 16 15 15 1 0 9 13 2
26 11 1 13 16 15 9 11 11 1 11 1 13 4 0 12 9 1 0 9 1 9 13 1 13 4 2
10 15 15 9 1 9 1 9 13 4 2
17 11 1 13 16 15 15 9 1 9 1 0 9 13 4 4 4 2
11 15 10 9 1 0 9 1 13 4 4 2
14 11 15 1 11 1 9 9 13 4 1 3 0 13 2
22 15 13 4 16 15 14 9 1 15 0 9 7 9 1 9 1 1 14 13 4 4 2
18 15 0 9 1 0 13 7 15 11 1 9 9 13 4 3 0 13 2
28 15 9 11 11 1 9 1 9 13 4 1 9 0 13 4 15 10 0 9 1 0 7 0 2 0 9 13 2
22 11 11 1 11 11 11 11 11 11 11 1 14 13 15 9 0 13 1 9 13 4 2
17 11 1 13 16 15 9 1 10 0 2 0 9 1 3 14 13 2
45 11 1 13 16 15 9 1 9 1 15 14 9 1 15 9 14 13 2 7 15 15 13 4 4 4 16 11 1 0 0 9 1 0 9 1 9 13 1 1 15 13 4 4 4 2
30 11 1 13 16 9 13 1 3 15 9 14 13 4 16 9 9 9 1 9 9 1 1 10 9 1 9 13 4 4 2
10 11 11 1 14 9 1 9 13 4 2
14 11 9 11 11 1 9 1 11 1 9 13 4 4 2
13 15 1 15 1 1 9 0 13 15 11 13 4 2
22 9 9 1 13 16 11 11 11 1 9 9 1 9 13 1 11 11 1 9 13 4 2
10 15 1 15 0 9 1 9 13 4 2
8 15 9 9 11 11 1 13 2
27 9 1 1 13 1 9 0 13 4 11 9 11 11 1 15 0 9 1 11 11 1 9 1 9 14 13 2
19 7 15 9 14 13 7 15 9 1 15 9 13 4 9 1 9 13 4 2
14 10 9 1 13 9 1 11 11 1 1 3 9 13 2
14 11 9 13 1 14 3 3 15 9 1 1 13 4 2
10 15 15 0 9 1 0 14 14 13 2
22 7 15 0 9 10 3 15 9 1 9 1 9 1 9 1 9 1 9 13 13 4 2
21 3 14 11 9 1 13 13 4 15 0 9 1 2 11 0 13 2 1 9 13 2
11 15 1 11 11 11 1 1 9 13 4 2
26 11 1 11 11 11 2 11 2 1 9 11 11 1 13 13 16 11 11 11 1 9 9 13 4 4 2
26 11 1 13 16 15 11 1 9 2 11 2 11 2 11 7 0 9 1 1 13 4 9 0 13 4 2
20 11 1 13 16 16 11 9 9 1 9 13 4 4 16 15 9 0 13 4 2
23 15 1 9 1 9 2 11 2 11 2 11 7 9 1 1 9 13 4 9 0 13 4 2
19 11 11 2 11 11 11 11 11 2 1 9 13 10 9 11 13 4 4 2
20 11 1 13 16 11 1 9 1 9 1 9 0 13 1 1 15 11 13 4 2
12 11 1 10 9 15 9 13 1 9 13 4 2
18 11 1 13 16 15 9 11 7 11 11 1 9 1 15 9 14 13 2
23 15 13 16 11 9 1 1 13 4 9 1 12 9 13 7 15 15 14 0 9 13 4 2
15 15 13 16 15 9 1 1 0 13 4 9 3 13 4 2
23 15 1 14 15 12 9 1 9 1 11 7 11 1 11 11 3 14 13 1 9 13 4 2
30 15 13 16 15 0 9 1 15 9 1 13 1 1 12 0 9 13 1 9 13 1 10 9 1 9 13 4 4 4 2
31 15 13 16 15 13 4 16 11 7 11 1 1 0 9 0 13 7 12 9 1 1 10 9 1 9 9 1 1 13 4 2
17 15 13 16 9 9 1 0 9 1 0 9 1 13 4 4 4 2
38 9 9 13 1 1 9 1 9 9 1 9 1 0 9 1 9 13 1 9 1 11 1 10 9 0 9 13 4 15 0 9 1 9 1 9 13 4 2
19 11 2 11 1 1 9 11 11 11 11 1 0 9 1 9 13 4 4 2
34 10 3 13 9 15 0 9 1 9 13 1 1 9 9 1 9 13 4 2 9 9 9 11 11 11 9 9 9 1 9 13 4 4 2
15 11 1 10 9 1 1 0 9 1 11 1 9 13 4 2
33 15 9 1 12 9 1 15 1 13 4 15 15 15 1 15 14 9 13 1 9 13 4 13 16 9 9 9 1 9 1 9 13 2
41 9 1 11 1 9 13 1 11 9 11 1 0 9 1 9 1 1 9 1 9 1 0 9 13 4 7 11 1 11 1 9 1 9 13 1 1 9 13 4 4 2
58 16 11 13 9 15 13 9 14 13 4 4 16 14 9 1 9 1 15 1 0 14 13 4 4 7 11 1 0 9 1 9 1 13 11 1 10 9 1 10 9 13 16 11 9 1 15 11 9 13 1 9 13 1 14 9 13 4 2
13 15 9 1 9 1 11 1 9 3 14 13 4 2
42 9 9 1 0 11 11 1 9 2 9 11 11 1 9 11 11 1 1 11 1 9 13 1 9 10 9 3 13 15 11 9 1 9 1 14 12 9 1 10 9 13 2
16 15 9 13 4 16 11 1 12 12 9 9 1 1 13 4 2
31 16 11 1 0 9 9 1 1 10 0 9 1 9 13 4 2 7 15 11 9 9 1 9 1 11 1 9 3 14 13 2
26 11 9 11 11 1 1 2 11 11 1 9 1 9 13 4 4 7 9 13 15 14 9 1 9 13 2
12 11 9 1 11 0 9 1 3 13 4 4 2
15 3 0 11 9 9 1 11 1 9 1 0 9 13 4 2
11 2 15 11 1 0 9 13 0 14 13 2
20 15 9 1 1 1 9 13 1 9 13 7 15 11 1 9 1 9 13 4 4
20 13 9 14 15 15 14 13 4 16 9 1 9 1 14 9 13 0 14 13 2
11 9 1 9 7 9 9 1 13 0 13 2
30 11 11 1 14 15 9 1 9 1 9 1 9 13 9 13 1 11 1 11 1 9 1 14 10 9 3 13 4 4 2
21 11 1 13 13 16 15 9 1 9 3 13 4 7 15 11 1 13 0 14 13 2
20 2 11 9 0 9 1 9 13 7 11 9 1 15 9 1 9 1 9 14 13
18 9 9 1 11 1 11 9 9 1 1 9 9 1 9 0 13 4 2
19 15 1 9 9 1 2 11 11 11 11 11 11 2 0 9 13 4 4 2
18 9 9 1 10 9 1 12 9 9 13 4 15 9 9 14 13 4 2
23 0 9 11 1 13 11 9 9 1 1 9 15 9 1 1 0 9 1 9 13 4 4 2
19 0 13 16 11 11 1 11 9 1 0 9 1 9 0 13 4 4 4 2
31 10 9 1 9 2 9 9 2 9 9 7 11 11 2 9 9 7 15 9 9 9 1 1 0 9 1 0 13 4 4 2
23 9 9 1 11 11 1 11 1 10 12 9 9 1 9 9 13 1 9 9 1 13 4 2
22 7 15 7 9 1 14 12 9 0 13 4 4 2 10 9 1 0 13 3 0 13 2
32 11 11 9 1 11 11 11 11 11 1 9 1 1 12 9 1 13 0 9 1 0 0 9 11 1 9 13 1 9 13 4 2
19 9 9 11 11 1 13 16 15 1 11 1 9 1 9 14 13 4 4 2
22 0 13 16 11 1 9 11 9 1 1 13 10 9 1 12 9 1 9 13 4 4 2
15 10 9 11 9 1 9 9 9 9 1 9 1 13 4 2
9 10 0 0 9 9 1 13 4 2
12 9 1 1 15 7 12 9 1 9 13 4 2
15 9 1 10 9 1 9 13 4 2 7 15 9 0 13 2
12 9 15 1 10 9 1 9 14 13 4 4 2
19 11 1 1 10 9 1 9 1 12 9 13 4 15 11 11 13 4 4 2
16 15 10 9 13 4 16 10 9 0 9 1 13 4 4 4 2
28 11 1 11 11 1 0 9 1 11 11 11 11 11 11 9 11 11 2 11 11 7 12 0 9 1 0 13 2
19 11 11 11 2 11 2 1 9 1 9 13 9 11 1 15 9 13 4 2
26 9 1 1 13 4 0 9 1 9 11 2 9 11 11 11 2 9 11 11 7 9 11 11 0 13 2
24 9 1 9 1 9 1 13 4 13 4 10 9 9 0 7 0 12 9 1 9 1 0 13 2
30 11 1 9 9 1 9 9 1 9 1 0 9 13 1 11 1 9 13 4 1 3 9 15 9 13 4 1 9 13 2
24 11 1 10 9 1 11 1 9 1 9 1 9 13 2 15 9 1 9 1 0 9 13 4 2
30 9 13 16 11 2 11 11 1 10 9 1 9 7 9 1 9 1 12 1 12 9 14 9 1 9 13 4 4 4 2
24 9 9 1 9 2 9 1 9 9 1 9 13 1 13 9 11 11 11 11 3 10 0 13 2
16 9 1 10 12 9 1 9 9 1 9 13 1 9 13 4 2
17 16 15 15 13 1 9 13 16 9 1 9 1 10 9 13 4 2
26 15 1 11 1 11 11 11 11 1 1 11 11 11 1 10 9 1 9 13 7 0 9 1 9 13 2
17 10 9 1 9 9 11 11 11 7 9 9 11 11 14 0 13 2
22 11 11 1 13 9 1 1 11 11 1 9 13 16 9 9 1 9 9 10 13 4 2
21 7 2 11 11 9 1 1 9 9 1 9 9 1 9 1 13 10 0 14 13 2
15 0 9 9 14 0 9 1 9 9 13 1 13 4 4 2
33 16 9 2 9 1 9 14 13 4 7 0 9 9 14 13 16 9 9 1 9 1 12 1 12 9 14 9 1 1 9 13 4 2
18 11 9 9 1 0 9 2 9 1 9 9 1 15 3 0 14 13 2
12 15 11 11 1 1 3 10 9 13 4 4 2
24 9 1 9 1 12 9 7 9 9 7 9 1 12 9 1 9 1 9 2 9 13 4 4 2
16 0 9 1 1 1 11 11 0 9 1 14 9 13 4 4 2
16 9 1 9 9 1 9 1 9 1 9 2 9 13 4 4 2
17 9 13 4 4 4 15 9 14 9 1 9 1 0 9 13 4 2
38 9 9 9 1 9 1 14 9 13 4 4 4 16 0 9 1 9 1 9 1 13 4 9 2 9 1 1 11 1 9 1 9 13 1 9 14 13 2
21 10 9 0 9 1 0 9 1 9 12 2 12 9 1 9 2 3 13 4 4 2
10 0 12 9 1 1 15 0 9 13 2
35 0 12 9 1 1 0 9 1 0 9 1 9 1 14 12 9 14 9 1 9 1 1 0 9 1 9 9 1 9 1 9 14 13 4 2
14 15 0 9 9 1 14 12 12 1 9 13 4 4 2
20 9 9 7 9 1 9 1 11 1 15 1 15 9 1 9 14 13 4 4 2
18 15 14 11 2 11 1 9 9 1 12 12 1 9 13 1 9 13 2
26 11 11 11 11 1 11 1 0 9 1 11 9 1 9 1 9 1 9 13 1 9 1 3 13 4 2
17 15 13 16 9 14 15 9 1 13 4 15 0 9 13 4 4 2
29 11 1 9 2 11 2 9 1 9 9 1 11 1 9 1 13 16 9 1 15 9 13 7 15 15 9 13 4 2
20 10 9 11 1 14 15 9 1 12 15 9 13 7 9 1 15 9 13 4 2
21 11 11 1 13 16 9 1 15 0 9 9 1 9 1 9 13 9 13 4 4 2
28 9 1 9 1 1 9 9 9 2 9 7 9 9 1 11 11 11 2 11 2 1 3 13 9 13 4 4 2
12 9 9 2 9 1 1 14 13 4 4 4 2
14 9 1 15 10 9 1 13 1 9 14 0 13 4 2
17 11 1 13 16 11 11 9 1 10 9 1 10 0 9 13 4 2
10 15 9 1 9 14 9 13 4 4 2
10 15 1 0 9 1 9 1 9 13 2
10 3 11 7 11 1 15 0 9 13 2
10 11 7 11 1 1 9 9 0 13 2
28 15 1 14 11 1 9 1 1 1 0 11 2 11 11 1 9 1 9 1 15 3 13 1 9 13 4 4 2
21 0 0 9 11 7 0 9 11 1 9 1 10 9 1 13 1 0 9 13 4 2
24 16 12 9 1 0 9 1 14 10 9 1 12 9 3 13 1 10 2 10 9 13 4 4 2
25 0 9 11 7 10 9 1 3 0 0 9 11 1 9 1 13 10 9 1 13 1 9 13 4 2
15 11 1 13 12 9 1 12 9 1 0 9 1 9 13 2
10 10 9 1 12 0 9 0 13 4 2
16 10 9 15 2 15 9 1 9 1 9 9 13 1 1 13 2
25 11 1 0 9 9 11 11 1 13 13 16 11 12 0 13 9 13 7 11 1 15 9 13 4 2
56 11 1 0 9 11 2 11 1 9 1 1 13 9 1 11 11 11 7 11 1 11 11 11 11 11 1 14 13 16 9 9 1 9 13 7 11 1 13 9 1 12 0 9 1 1 14 10 9 1 9 2 9 1 9 13 2
17 15 1 10 9 1 9 1 10 10 9 1 13 0 13 4 4 2
15 15 9 1 3 0 0 9 13 11 11 1 13 4 4 2
17 16 15 12 9 1 1 9 2 9 1 1 11 11 13 4 4 2
22 11 1 9 11 11 11 1 13 16 15 10 9 1 3 14 11 11 11 1 1 13 2
27 11 11 11 1 11 1 3 13 4 16 11 1 13 1 0 9 9 1 9 0 11 9 1 0 9 13 2
18 15 1 14 9 11 1 0 11 9 1 12 0 9 13 1 9 13 2
18 11 9 1 13 1 1 9 1 11 11 7 11 11 1 11 13 4 2
10 16 0 9 1 9 9 13 4 4 2
14 10 9 11 1 9 1 9 11 11 1 9 1 13 2
32 15 13 16 11 11 9 1 13 4 9 10 9 1 9 13 4 4 7 10 0 9 1 9 1 10 9 1 9 13 4 4 2
12 11 1 11 0 11 9 1 1 0 9 13 2
16 11 1 13 16 10 0 9 1 9 9 1 13 1 0 13 2
9 7 9 15 1 1 13 4 4 2
17 15 13 16 11 11 1 10 0 9 14 11 1 0 13 13 4 2
24 11 9 11 11 7 11 9 11 11 1 11 1 13 1 9 1 11 9 1 9 1 13 4 2
26 15 13 16 10 9 1 15 1 1 9 13 4 4 7 3 10 9 1 9 1 9 13 0 14 13 2
40 9 9 1 13 16 11 1 13 9 1 9 1 10 0 9 1 9 1 9 13 7 15 12 9 0 13 4 4 16 11 9 1 10 9 1 1 0 9 13 2
24 11 1 11 1 9 1 9 1 0 13 1 9 1 15 13 16 15 9 1 9 13 4 4 2
36 11 1 13 16 9 1 1 15 1 1 9 13 4 16 10 9 1 9 13 4 7 16 9 1 1 15 13 4 16 15 9 1 0 13 4 2
9 15 15 1 1 9 13 4 4 2
42 11 1 11 1 9 1 0 13 1 9 1 11 1 13 16 11 1 9 11 1 9 1 9 1 1 13 7 11 1 9 13 1 3 14 15 1 1 15 9 13 4 2
18 11 1 13 2 4 9 13 4 11 7 11 10 3 13 13 4 4 2
29 11 1 9 15 9 13 4 13 16 11 11 11 1 11 9 1 1 12 9 9 11 11 1 11 9 1 9 13 2
27 9 14 0 11 11 11 11 1 13 4 16 0 11 1 9 0 9 1 13 16 15 1 9 13 4 4 2
39 11 1 11 11 11 11 11 1 11 1 9 1 1 11 11 1 9 1 9 0 13 4 13 2 15 11 11 11 11 13 4 4 2 15 15 1 9 13 2
21 11 11 11 1 0 9 1 1 1 12 0 9 1 11 11 1 11 13 4 4 2
24 11 1 11 1 13 16 15 11 9 1 1 11 11 11 1 1 11 1 0 9 1 9 13 2
14 11 1 13 16 15 0 11 11 1 11 0 13 4 2
16 15 1 15 11 1 13 7 15 9 9 1 9 14 0 13 2
31 11 1 0 9 9 1 9 1 11 11 1 9 1 9 13 4 13 16 11 9 1 9 1 1 15 0 7 0 9 13 2
22 7 14 15 1 12 9 1 0 9 13 7 15 11 11 9 1 1 9 13 4 4 2
31 11 1 13 16 11 13 4 16 11 0 9 1 3 13 7 10 9 13 4 15 9 1 0 9 1 1 1 9 13 4 2
12 15 13 2 15 9 13 4 16 15 0 13 2
10 15 0 9 15 1 10 9 13 4 2
17 12 9 1 15 0 13 4 16 15 15 0 9 1 9 14 13 2
34 15 13 1 16 15 10 10 9 13 4 16 11 0 9 1 1 0 13 2 11 1 13 16 15 1 9 13 1 1 0 9 14 13 2
12 16 15 15 1 15 13 16 15 3 9 13 2
7 15 10 9 14 13 13 2
25 11 1 9 13 16 11 1 11 7 11 1 1 0 9 13 4 4 7 15 1 9 13 4 4 2
20 15 13 16 0 9 15 13 16 10 9 9 7 9 1 1 14 13 4 4 2
27 15 13 16 10 9 11 1 9 9 9 11 11 11 7 11 1 9 9 9 11 11 1 1 13 4 4 2
29 11 1 13 16 16 9 11 7 11 1 0 13 7 9 15 0 13 4 16 9 1 15 14 9 0 14 13 4 2
22 15 13 16 15 0 9 13 16 0 11 11 11 9 1 11 13 1 9 13 4 4 2
31 11 1 11 9 11 11 1 11 9 1 9 1 9 1 11 11 11 11 11 11 1 9 13 1 11 1 9 13 4 4 2
22 11 11 1 0 9 1 11 1 13 16 11 7 11 1 0 9 1 0 9 13 4 2
39 11 1 9 11 11 11 1 11 11 1 15 13 16 11 11 11 1 10 9 1 9 13 4 15 13 4 4 16 11 1 11 1 0 9 1 11 9 13 2
16 15 13 16 11 7 11 1 15 0 9 1 0 9 13 4 2
23 11 1 11 1 10 9 1 10 0 9 13 1 9 13 15 10 9 1 0 9 13 4 2
23 15 9 13 16 11 9 1 9 11 1 9 1 11 1 9 1 0 9 1 10 0 13 2
29 11 1 13 16 15 9 13 4 16 11 9 1 9 1 9 9 1 10 13 1 1 11 9 1 9 13 4 4 2
24 11 11 11 1 11 9 1 9 1 1 0 9 1 9 1 9 1 0 9 1 0 13 4 2
21 15 13 16 12 9 10 9 1 9 1 9 13 4 4 15 12 9 1 0 13 2
33 11 11 11 1 11 1 11 11 1 11 11 9 1 11 9 1 11 11 11 11 11 1 9 1 1 9 1 9 1 10 9 13 2
35 10 9 1 0 9 11 11 11 7 11 11 11 2 11 11 1 11 11 11 11 2 11 11 11 11 11 7 9 1 9 7 9 0 13 2
23 11 11 11 1 13 16 11 9 1 9 1 1 15 0 9 1 9 1 15 9 14 13 2
12 12 9 1 1 0 9 1 10 9 13 4 2
28 3 1 12 9 1 0 13 4 11 11 1 13 16 13 1 9 1 11 11 11 11 9 1 10 9 13 4 2
21 9 1 1 9 1 13 1 1 3 1 15 11 11 11 1 0 13 4 4 4 2
20 11 1 13 16 11 9 1 11 11 11 1 0 9 1 10 9 13 4 4 2
24 15 13 16 0 9 1 0 13 1 1 9 9 9 1 0 13 15 9 1 9 1 0 13 2
27 11 1 13 16 9 9 11 1 9 1 9 1 0 13 1 1 11 11 11 11 11 9 13 13 4 4 2
22 0 9 1 1 11 11 11 11 11 1 3 9 1 3 0 12 12 9 1 13 4 2
16 10 9 1 1 9 1 10 9 14 9 12 9 9 13 4 2
9 0 9 1 12 9 9 13 4 2
21 11 11 10 9 1 1 9 1 0 9 9 0 13 1 1 9 7 9 0 13 2
28 9 9 2 9 9 2 9 9 2 9 9 7 9 1 0 9 1 13 1 9 1 9 9 1 1 13 4 2
28 10 9 1 1 11 11 1 12 9 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 1 13 4 2
31 2 11 11 11 11 11 2 9 1 1 11 11 13 9 1 13 1 11 11 1 0 11 11 11 13 1 9 13 4 4 2
41 9 0 13 4 15 13 16 11 1 0 9 1 13 1 1 3 0 9 1 9 1 9 2 13 4 9 7 0 0 0 9 1 0 13 14 10 9 13 4 4 2
18 11 1 9 1 9 11 11 1 9 13 9 14 13 1 9 13 4 2
31 0 9 11 11 1 9 1 9 11 1 1 15 9 2 11 11 11 11 11 2 1 10 3 0 9 13 1 9 13 4 2
7 15 0 9 1 9 13 2
25 9 1 0 9 11 7 11 1 1 13 4 4 7 15 11 11 1 9 1 0 9 13 4 4 2
38 11 1 9 13 1 9 1 1 9 1 10 9 1 0 9 1 1 9 13 4 13 4 16 15 9 1 9 7 10 9 1 0 9 1 1 9 13 2
16 7 9 1 0 9 1 1 15 10 9 1 9 13 4 4 2
33 11 1 0 12 9 1 13 4 16 0 9 1 9 2 9 9 2 13 9 7 0 9 1 11 11 1 9 1 15 9 13 4 2
26 15 13 13 16 15 14 9 15 10 9 1 1 0 13 7 9 15 14 9 1 15 0 13 13 4 2
17 15 13 4 16 9 1 0 9 1 1 1 9 9 13 4 4 2
11 9 1 15 9 1 0 13 4 4 4 2
44 11 1 9 1 9 1 0 9 2 11 1 0 9 1 9 13 4 9 9 1 9 2 7 11 1 9 9 1 9 13 4 9 1 9 1 9 9 1 10 9 1 9 13 2
32 15 1 2 11 11 11 11 11 2 1 11 7 11 1 11 11 11 1 13 9 1 1 1 0 9 9 1 9 13 4 4 2
24 11 1 11 1 15 0 9 2 11 11 11 11 11 2 1 1 11 11 1 0 13 4 4 2
32 7 10 9 15 15 9 1 3 14 9 13 1 1 13 16 10 9 0 7 0 9 1 0 13 7 15 9 9 1 13 4 2
17 15 13 16 9 1 1 11 1 9 15 9 1 9 14 13 4 2
23 9 1 9 9 1 0 9 1 13 1 1 9 9 11 11 1 11 1 0 9 13 4 2
9 9 1 9 9 11 1 9 13 2
12 10 9 9 9 1 0 13 1 10 9 13 2
20 9 9 9 1 0 9 9 13 1 3 10 9 0 9 13 1 9 13 4 2
17 9 10 9 1 9 1 9 0 9 1 13 1 1 9 13 4 2
32 7 10 9 9 7 15 9 1 0 9 1 9 1 13 4 9 9 1 1 9 1 9 2 9 7 9 10 13 1 9 13 2
21 15 11 13 4 16 10 9 1 9 1 0 9 1 13 1 9 1 9 13 4 2
13 3 9 1 0 9 1 9 14 15 9 1 13 2
18 9 9 10 9 1 9 1 9 1 9 14 13 1 9 13 4 4 2
22 15 1 1 15 10 9 1 9 7 10 9 1 0 9 1 9 13 9 13 4 4 2
8 14 11 1 9 10 0 13 2
13 15 9 1 15 10 9 1 9 9 1 13 4 2
8 9 9 1 14 9 13 4 2
11 7 9 1 10 9 9 14 0 13 4 2
19 10 0 9 1 13 4 9 9 11 11 11 1 10 9 1 9 1 13 2
23 16 15 1 15 11 9 11 11 1 1 11 7 11 1 9 1 0 2 0 13 4 4 2
35 0 11 11 11 11 1 9 1 1 11 11 11 1 11 11 1 0 11 11 11 11 1 9 13 4 1 9 1 0 9 0 13 4 4 2
10 11 1 15 1 0 9 0 13 4 2
24 9 1 13 4 16 11 1 9 1 0 9 1 0 9 1 9 14 13 1 9 1 13 4 2
27 9 1 3 1 9 13 4 11 11 11 1 14 11 1 9 1 9 13 4 11 1 9 1 3 13 4 2
30 11 1 11 1 0 9 13 4 11 1 10 9 1 1 9 13 4 16 15 9 1 13 14 14 9 1 9 13 4 2
14 11 1 11 9 11 1 11 1 12 9 1 9 13 2
15 11 1 9 9 11 11 1 10 9 1 9 1 9 13 2
29 11 1 13 16 11 1 11 1 13 16 0 9 1 0 11 2 11 11 11 1 11 1 9 13 1 15 9 13 2
30 11 1 13 16 11 1 0 9 1 0 9 1 13 9 1 9 1 12 0 9 1 9 13 4 2 15 0 9 13 2
25 11 9 1 9 1 14 1 11 1 10 9 1 11 1 9 1 13 1 12 0 9 13 4 4 2
32 11 9 11 11 11 1 13 16 15 1 0 9 1 15 0 9 13 4 16 15 14 9 9 1 0 0 9 1 14 13 4 2
18 7 9 11 1 11 1 1 11 1 9 13 10 9 1 13 4 4 2
23 15 13 16 11 11 13 4 10 9 9 13 2 7 15 15 14 0 0 9 1 14 13 2
17 15 13 16 11 1 9 1 9 9 1 9 1 9 0 13 4 2
11 15 13 9 0 9 1 9 14 0 13 2
35 11 1 9 1 9 0 13 4 11 9 11 11 11 1 13 16 15 1 9 1 7 15 1 15 13 2 15 11 1 13 1 10 9 13 2
5 15 15 9 13 2
8 15 1 0 9 15 14 13 2
18 7 2 11 11 1 9 1 9 13 1 9 1 1 15 9 14 13 2
25 3 10 9 15 11 11 1 12 9 1 1 13 9 1 0 15 9 1 15 15 9 14 13 4 2
15 9 1 13 13 16 15 9 15 11 11 14 13 4 4 2
38 9 9 11 11 1 15 1 1 9 13 4 13 16 13 4 4 11 11 1 15 11 1 10 9 1 9 13 4 7 11 11 1 9 9 1 13 4 2
19 16 2 10 9 1 1 11 1 13 16 11 3 0 9 1 9 13 4 2
19 10 9 13 4 1 16 15 11 1 0 9 1 10 9 1 9 13 4 2
11 15 13 13 16 9 15 1 13 14 4 2
16 11 1 13 16 11 1 16 15 13 4 16 15 0 14 13 2
17 11 11 11 11 1 14 11 1 9 1 0 9 0 9 13 4 2
17 11 9 11 11 1 13 16 11 1 9 13 15 0 9 14 13 2
17 9 1 1 15 9 15 1 12 10 9 1 1 0 13 4 4 2
19 9 1 12 0 9 1 9 13 10 9 1 9 1 13 1 9 13 4 2
25 15 1 9 9 9 7 0 9 13 9 1 15 13 1 9 13 4 4 16 15 14 15 9 13 2
16 11 1 11 0 9 1 9 1 10 9 15 0 13 4 4 2
12 11 1 14 10 9 0 9 1 9 1 13 2
17 15 12 9 1 12 9 1 9 13 7 9 12 9 13 13 4 2
14 0 9 1 1 9 1 9 15 9 0 13 4 4 2
11 9 14 9 1 10 9 1 13 4 4 2
20 9 1 9 1 9 13 1 1 9 14 9 13 9 9 13 1 13 4 4 2
14 9 1 13 1 1 9 1 14 9 9 0 13 4 2
12 10 9 1 12 9 1 9 1 13 4 4 2
12 15 9 1 9 1 14 12 9 0 13 4 2
12 10 9 1 11 1 9 1 9 13 4 4 2
19 9 1 9 13 16 10 9 15 13 4 7 15 9 9 1 15 0 13 2
13 11 9 12 9 10 9 1 9 14 13 4 4 2
17 7 3 1 9 1 9 7 0 9 1 1 1 9 1 13 4 2
23 11 1 12 0 9 9 1 9 13 16 9 1 0 9 0 9 1 3 0 13 4 4 2
17 9 1 0 13 1 1 1 12 9 1 9 1 9 13 14 4 2
39 9 1 11 11 1 9 1 11 1 11 11 1 9 1 1 13 4 9 1 9 9 1 10 9 1 3 0 13 4 1 1 1 11 1 9 9 13 4 2
12 9 1 13 12 9 1 9 1 3 9 13 2
12 10 3 12 9 1 9 13 9 13 4 4 2
10 9 7 9 1 9 9 0 13 4 2
19 9 1 0 13 1 12 9 1 12 9 7 9 1 9 14 0 13 4 2
25 9 1 12 9 1 10 9 1 9 2 9 7 9 2 9 1 1 14 15 9 1 9 13 4 2
14 9 1 9 1 13 4 9 1 9 13 4 4 4 2
13 0 9 1 1 9 9 1 9 1 0 13 4 2
15 9 1 11 2 11 11 1 9 1 1 9 14 13 4 2
18 9 1 9 9 1 9 2 9 13 13 4 12 9 1 9 13 4 2
6 15 9 13 4 4 2
22 9 1 11 11 1 9 1 11 1 9 11 11 11 1 1 1 11 11 13 4 4 2
22 9 1 9 9 1 9 1 9 9 1 13 15 0 13 1 1 9 1 9 1 13 2
18 9 1 9 0 14 13 15 9 9 1 9 1 3 9 0 13 4 2
8 15 11 11 9 14 13 4 2
23 10 9 1 9 1 9 1 11 1 9 14 12 12 9 11 11 1 1 9 9 13 4 2
9 3 11 11 1 14 9 13 4 2
15 12 9 9 1 9 7 0 9 1 3 9 2 9 13 2
13 9 9 1 13 1 3 14 15 9 13 4 4 2
9 9 1 15 13 9 13 4 4 2
11 15 9 13 14 9 1 9 13 4 4 2
18 16 15 1 14 9 2 9 2 9 2 9 7 9 1 9 13 4 2
13 9 1 11 9 0 12 0 9 1 9 13 4 2
16 9 1 9 9 7 11 0 10 9 1 9 1 9 13 4 2
15 9 2 9 7 9 1 14 12 12 1 10 1 9 13 2
9 12 9 9 1 14 13 4 4 2
22 9 9 1 9 13 1 1 9 9 13 4 2 7 15 9 1 9 1 14 13 4 2
18 9 1 9 11 11 1 10 9 9 7 9 1 9 14 0 13 4 2
12 9 1 9 13 1 3 9 1 9 0 13 2
41 9 1 11 2 11 11 3 14 11 9 1 13 9 1 14 3 15 1 9 13 2 16 9 13 9 13 1 9 14 13 4 2 15 9 1 9 1 0 13 4 2
20 3 9 1 9 9 1 9 2 9 13 13 4 12 9 11 1 9 13 4 2
5 15 9 13 4 2
16 11 1 9 11 11 1 9 10 13 1 9 14 13 4 4 2
23 3 9 1 9 0 13 7 15 15 1 9 1 0 9 7 9 13 1 9 13 4 4 2
21 10 9 1 9 1 13 1 1 9 1 0 9 1 1 11 11 1 9 13 4 2
15 13 4 4 4 16 11 1 10 9 1 9 13 4 4 2
15 11 1 13 4 16 15 1 13 4 9 0 7 0 13 2
30 11 9 1 11 0 11 9 1 12 0 9 11 1 9 7 12 0 9 1 1 9 7 9 9 13 1 9 13 4 2
35 11 9 1 9 0 13 1 11 1 13 4 16 10 9 11 11 1 9 1 9 1 9 7 0 2 9 9 2 1 0 9 0 13 4 2
13 10 9 11 1 13 7 15 9 1 9 9 13 2
14 9 1 9 1 9 1 14 9 10 9 1 13 4 2
19 9 1 1 11 11 9 13 9 13 4 7 15 15 12 9 1 13 4 2
28 11 1 15 9 1 13 4 16 9 1 9 1 14 15 9 1 9 2 9 2 1 3 13 9 1 13 4 2
16 10 9 9 7 15 9 2 1 1 9 15 9 13 13 4 2
27 15 13 16 9 1 9 1 1 1 15 15 9 14 13 7 15 15 14 9 14 13 16 3 9 15 13 2
56 11 1 10 9 1 15 9 14 13 16 11 9 11 11 1 15 0 9 11 1 9 2 11 2 1 13 4 2 7 15 10 9 14 13 4 4 4 16 11 11 11 9 1 9 1 13 14 10 9 1 3 13 13 13 4 2
22 7 10 9 1 11 1 9 1 9 1 13 4 4 7 11 1 9 13 4 4 4 2
37 11 9 11 11 1 9 10 9 1 9 13 4 16 11 0 9 1 1 14 11 11 1 13 1 9 13 4 2 15 15 9 1 1 13 4 4 2
17 15 0 9 1 1 9 1 9 0 13 1 9 14 0 13 4 2
15 15 13 16 9 1 1 9 1 9 1 15 9 14 13 2
41 11 1 13 16 11 1 15 9 11 11 1 13 4 9 13 4 4 4 2 9 1 11 11 0 9 1 13 1 9 1 1 14 12 9 1 1 11 1 13 4 2
16 12 9 1 15 11 1 10 9 13 15 14 13 4 4 4 2
11 9 1 10 9 1 15 9 9 14 13 2
17 11 1 10 9 1 13 11 11 1 9 1 9 13 1 9 13 2
31 11 11 11 11 11 1 11 11 1 13 9 1 1 1 9 1 13 16 16 15 1 9 13 4 16 15 15 9 13 4 2
28 12 9 1 9 1 9 1 11 9 1 13 16 15 11 9 11 11 14 13 4 4 16 15 10 0 9 13 2
11 15 15 10 9 1 9 13 4 4 4 2
30 9 1 0 7 9 1 0 13 1 1 9 9 11 11 1 12 9 13 4 2 15 15 0 9 1 0 13 4 4 2
19 9 1 1 9 9 1 1 9 1 1 0 12 9 1 14 9 1 13 2
21 15 9 1 9 1 14 11 1 11 9 1 1 13 4 12 9 1 9 13 4 2
44 11 1 9 1 1 9 1 13 16 15 15 0 13 1 1 9 13 4 4 16 9 13 1 10 9 9 1 0 13 7 15 9 1 9 13 4 15 15 9 1 1 0 13 2
27 10 9 1 11 1 9 11 11 11 1 9 13 16 9 1 10 9 1 3 0 9 9 1 1 13 4 2
20 15 1 9 1 13 16 15 10 9 1 15 1 0 9 1 9 2 9 13 2
47 9 1 9 0 13 1 1 1 9 1 9 1 0 9 13 4 11 1 13 16 9 1 9 1 9 13 1 1 15 0 9 1 10 11 9 1 10 9 1 9 13 16 10 9 0 13 2
14 15 9 1 13 16 15 15 9 1 0 9 13 4 2
18 9 1 11 1 9 1 9 1 9 1 3 13 4 1 9 13 4 2
11 15 1 11 11 9 9 1 1 13 4 2
23 11 1 11 1 9 1 12 9 1 13 0 9 1 10 14 10 12 9 1 9 13 4 2
12 9 1 14 12 9 1 0 13 1 9 13 2
16 12 9 9 11 1 12 9 1 11 1 11 11 1 0 13 2
23 9 9 11 11 1 9 1 12 9 1 9 13 7 12 9 1 0 13 1 9 13 4 2
28 11 9 1 9 9 11 11 11 11 1 13 16 12 9 1 11 1 11 11 11 7 9 1 13 4 4 4 2
19 11 2 11 7 11 1 0 9 1 14 14 12 9 1 9 13 4 4 2
14 9 1 13 1 9 1 12 9 7 12 9 0 13 2
17 11 1 13 16 12 9 1 9 11 11 1 0 13 4 4 4 2
15 9 1 13 1 1 11 1 9 1 12 9 14 0 13 2
27 11 2 11 11 2 11 11 1 13 16 15 13 4 16 9 1 9 1 1 9 1 9 13 1 9 13 2
20 9 1 9 7 11 11 1 9 11 1 13 16 3 15 0 9 1 9 13 2
12 15 1 13 10 9 1 3 1 9 13 4 2
20 9 1 1 0 9 1 9 13 1 1 13 1 9 9 1 9 0 13 4 2
23 9 1 0 0 11 11 1 13 16 9 1 9 1 9 13 4 7 9 9 1 13 4 2
19 11 1 9 1 0 11 1 9 1 9 1 11 1 9 1 9 13 4 2
25 11 1 11 11 11 7 11 1 11 11 11 1 1 13 9 1 11 1 9 1 9 1 9 13 2
34 0 9 9 1 1 9 9 11 11 1 12 9 1 1 12 9 1 10 9 1 13 9 1 11 1 9 1 9 1 9 1 9 13 2
17 15 13 16 11 1 10 9 1 9 13 1 11 1 9 13 4 2
25 11 1 12 9 1 9 1 1 12 0 9 1 9 13 15 11 11 1 9 1 11 1 13 13 2
10 16 15 11 9 1 15 9 14 13 2
59 11 1 11 1 9 1 15 12 9 13 4 15 11 11 11 1 11 1 12 9 1 13 9 9 1 1 11 1 13 4 9 1 9 1 0 13 4 13 4 16 9 0 9 0 13 7 15 10 9 1 15 9 1 9 14 13 4 4 2
16 9 11 11 11 1 15 9 1 9 1 9 1 0 13 4 2
22 11 1 10 9 1 13 1 9 9 1 9 1 11 1 9 9 1 9 13 4 4 2
41 9 1 12 9 1 11 1 9 1 9 13 4 11 1 3 11 9 1 9 9 1 1 13 1 9 13 4 2 3 15 9 1 0 9 1 1 14 9 13 4 2
36 11 2 11 2 1 9 1 11 1 13 4 11 1 9 1 11 1 3 13 1 9 13 4 13 4 16 11 2 11 9 1 10 0 9 13 2
16 16 10 9 9 9 1 11 1 9 13 1 1 13 4 4 2
15 12 9 13 9 1 0 9 0 9 9 1 9 13 4 2
49 11 9 1 9 1 1 9 13 1 9 0 13 1 3 11 1 9 9 9 1 10 0 13 2 11 1 11 11 11 13 7 0 9 7 9 1 9 1 11 9 1 13 1 9 13 1 13 4 2
25 10 9 11 1 9 1 14 12 9 1 11 1 0 13 1 11 9 1 9 1 9 0 13 4 2
23 11 1 0 9 9 1 1 10 9 1 3 13 9 1 3 10 0 13 1 9 0 13 2
21 11 11 9 1 9 1 13 4 11 1 11 0 9 1 3 13 1 9 13 4 2
10 11 1 9 11 11 11 1 1 13 2
52 11 1 9 1 0 13 1 9 1 1 9 1 1 11 9 11 11 1 13 16 15 11 9 1 3 14 0 9 1 9 1 13 4 2 7 0 9 1 13 4 9 1 1 11 9 1 1 15 9 13 4 2
14 9 10 9 1 9 13 16 9 1 3 9 13 4 2
26 11 1 9 13 16 11 9 1 3 9 1 0 9 7 9 1 9 13 7 11 0 9 1 0 13 2
76 0 11 11 11 11 1 9 1 0 10 9 1 11 1 1 11 1 11 11 2 11 11 2 11 11 7 11 11 11 2 11 11 1 11 11 2 11 11 7 11 11 2 11 11 11 1 11 11 11 2 11 11 11 1 11 11 11 2 11 11 1 11 11 7 11 11 11 11 1 11 11 11 1 9 13 2
20 11 1 0 9 1 0 9 1 9 1 11 9 1 13 1 9 13 4 4 2
45 11 1 11 1 1 9 0 13 1 9 1 9 1 13 4 9 1 9 13 4 13 4 16 11 11 1 9 1 11 7 11 11 1 13 4 9 9 1 0 9 1 3 0 13 2
52 12 9 1 9 13 4 0 11 11 11 11 1 13 16 11 1 15 13 16 2 10 9 13 4 2 7 11 11 1 10 9 16 9 11 1 9 1 9 13 2 9 1 9 1 0 9 1 9 14 13 4 2
19 9 1 14 12 12 9 15 13 15 0 13 1 0 9 14 13 4 4 2
22 3 14 12 12 9 15 13 15 10 13 1 1 1 0 9 1 9 1 13 4 4 2
31 15 13 9 1 13 1 13 4 4 16 9 1 13 1 10 9 1 1 12 9 1 9 1 9 2 9 14 0 9 13 2
18 9 9 1 9 13 16 10 9 1 13 1 1 0 9 9 13 4 2
10 16 0 13 1 9 0 13 4 4 2
35 11 11 11 1 9 9 11 11 11 1 1 9 1 12 9 9 0 9 9 2 12 9 0 9 9 7 14 12 9 0 9 9 1 13 2
19 7 0 9 1 12 9 9 1 14 12 12 9 15 13 15 3 0 13 2
10 15 1 0 0 9 14 0 14 13 2
33 11 11 11 11 2 11 2 11 1 0 9 9 11 11 1 13 16 9 7 10 9 12 9 1 13 1 0 9 0 13 4 4 2
13 9 1 9 1 1 15 0 9 14 13 4 4 2
22 9 11 1 9 13 16 9 11 11 11 1 1 10 9 1 12 9 1 9 0 13 2
15 7 0 9 1 0 13 1 1 9 9 13 1 9 13 2
15 10 9 1 11 1 9 14 1 12 9 1 0 13 4 2
11 7 15 15 10 10 9 9 13 4 4 2
25 0 9 1 1 9 1 1 11 9 1 0 9 1 1 13 9 9 1 13 9 1 0 13 4 2
20 15 9 1 3 13 9 1 9 1 9 0 9 1 13 1 9 13 4 4 2
21 16 9 1 9 7 9 1 9 9 1 9 1 14 13 16 9 10 9 1 13 2
24 0 11 11 1 11 1 0 9 1 0 9 1 1 9 1 9 1 12 9 1 9 13 4 2
16 9 1 1 9 1 9 1 13 4 9 1 9 9 13 4 2
23 9 9 14 10 9 13 4 4 16 9 0 13 7 11 1 11 1 1 12 9 9 13 2
20 7 2 9 1 13 9 1 9 1 9 7 9 9 1 9 1 9 13 4 2
22 9 1 9 1 1 9 10 9 0 13 4 16 15 3 13 1 9 14 0 13 4 2
20 11 0 9 9 1 9 1 13 13 16 9 1 9 9 1 1 13 4 4 2
10 15 9 1 3 13 1 9 13 4 2
10 0 12 9 1 9 3 13 4 4 2
20 11 11 1 9 1 1 9 1 9 7 9 1 9 9 1 9 1 0 13 2
24 9 9 1 9 1 9 1 1 14 13 7 9 1 9 13 1 3 14 15 0 14 13 4 2
12 15 3 9 1 1 9 1 9 13 4 4 2
24 15 9 1 9 1 9 14 13 7 2 9 1 9 7 9 1 9 10 13 1 9 14 13 2
15 16 2 0 9 1 15 9 1 13 7 9 14 10 13 2
23 11 1 9 11 1 14 12 9 1 11 9 1 0 9 1 11 1 9 9 1 13 4 2
11 9 9 11 11 11 1 10 9 13 4 2
13 11 1 13 16 9 1 10 9 9 1 0 13 2
21 9 1 11 7 11 11 9 9 1 1 9 12 9 14 12 9 9 9 13 4 2
16 14 12 9 1 9 9 0 13 1 3 9 0 13 4 4 2
12 10 9 1 9 9 3 14 9 13 4 4 2
15 9 15 12 9 1 0 9 13 9 1 9 13 4 4 2
23 10 3 0 9 1 9 1 9 13 4 9 1 10 9 9 1 9 14 13 4 4 4 2
28 0 11 7 11 9 1 11 9 1 1 0 9 10 9 9 1 0 13 1 9 1 9 1 9 13 4 4 2
17 11 3 0 9 1 1 12 13 2 15 1 9 1 0 9 13 2
12 9 9 1 15 1 12 9 9 13 4 4 2
13 10 9 1 11 11 11 11 1 14 9 0 13 2
29 11 1 0 12 9 1 13 16 15 14 9 0 9 15 9 1 9 13 4 4 7 15 3 10 0 9 1 13 2
14 9 1 13 1 3 12 9 11 1 9 13 4 4 2
33 11 1 9 9 11 11 11 1 13 16 11 7 11 1 9 1 13 4 9 1 13 1 9 1 9 1 1 15 10 9 13 4 2
9 10 9 9 1 9 13 4 4 2
26 15 0 9 1 9 9 13 1 13 11 1 12 0 9 11 11 7 11 11 9 9 1 0 9 13 2
27 9 1 9 7 0 9 1 1 0 9 1 9 13 4 12 9 1 11 2 11 1 0 9 1 0 13 2
10 15 1 0 9 10 9 1 0 13 2
17 11 11 1 13 16 11 11 11 1 0 9 1 15 9 14 13 2
11 10 9 15 10 9 1 9 13 4 4 2
25 9 1 9 1 1 0 9 1 11 11 1 13 16 10 9 1 11 1 11 11 1 3 13 4 2
14 9 1 0 13 1 3 12 9 1 11 1 9 13 2
15 10 3 11 11 9 9 1 12 9 1 9 1 13 4 2
51 11 11 1 13 16 10 9 1 9 1 9 1 11 11 7 11 11 11 1 10 9 1 0 9 1 0 9 1 13 9 7 9 1 13 4 4 4 2 15 1 11 1 12 9 0 7 0 13 4 4 2
19 9 7 0 9 1 9 1 1 15 9 13 4 12 9 0 13 4 4 2
19 11 1 9 13 10 9 1 11 11 3 11 1 13 1 1 9 0 13 2
12 15 10 9 1 11 1 11 11 1 9 13 2
12 15 1 2 11 1 0 9 1 9 13 4 2
28 11 1 11 1 11 9 1 11 1 0 9 1 9 13 1 9 15 9 1 0 13 4 2 15 9 13 4 2
17 0 9 9 11 1 10 9 1 11 1 9 1 13 1 9 13 2
33 11 1 9 13 1 3 14 15 9 9 0 9 11 1 9 1 9 13 0 9 1 13 15 11 1 9 1 9 1 9 14 13 2
16 11 1 11 9 1 12 9 1 11 1 1 0 13 4 4 2
26 15 9 11 1 15 13 7 9 1 9 1 0 13 9 1 13 4 15 11 1 3 9 1 13 4 2
20 11 1 11 11 11 1 11 11 1 13 2 9 1 15 9 1 0 9 13 2
21 3 1 9 1 0 9 1 9 1 10 9 1 13 4 15 9 1 13 4 4 2
24 9 1 13 13 16 11 1 9 1 9 1 9 1 9 1 9 1 1 1 13 1 9 13 2
24 11 1 12 9 9 1 13 1 3 11 2 11 0 11 1 9 11 1 0 9 3 13 4 2
25 9 9 1 13 9 1 9 1 9 1 12 9 1 1 9 1 3 13 9 1 9 1 13 4 2
23 9 1 13 16 10 9 11 1 9 12 9 14 9 1 9 1 9 1 9 1 9 13 2
19 15 15 9 1 13 4 4 15 12 9 1 9 1 9 1 0 9 13 2
31 10 9 1 9 11 1 11 11 11 1 13 4 7 15 1 12 12 12 12 9 2 14 12 12 9 2 1 9 13 4 2
27 11 1 1 10 9 1 11 1 0 9 7 9 1 9 1 0 9 1 1 1 9 1 0 9 13 4 2
26 15 1 11 1 9 1 1 9 9 9 13 13 4 11 1 11 11 11 9 9 1 0 13 4 4 2
23 0 13 16 11 1 0 11 1 12 12 9 1 9 0 13 7 9 1 12 9 9 13 2
22 9 1 9 1 0 3 9 13 4 11 1 11 9 9 1 9 13 14 9 13 4 2
21 10 9 3 9 9 1 0 9 1 9 13 4 4 2 3 15 9 1 14 13 2
41 9 9 1 9 1 0 9 1 1 9 9 1 15 0 9 13 1 9 0 9 1 9 2 0 11 9 1 0 9 14 13 7 15 0 9 13 13 4 4 4 2
33 10 9 1 15 14 0 13 4 4 16 11 1 1 9 1 9 13 1 0 9 1 1 11 1 15 3 10 9 14 13 4 4 2
19 10 9 1 14 13 9 9 1 11 1 9 0 2 14 2 9 13 4 2
16 0 9 1 11 7 11 1 15 0 9 1 0 9 13 4 2
23 10 12 9 1 14 12 0 9 1 11 1 1 11 7 11 1 9 1 9 13 4 4 2
22 11 1 9 9 1 10 13 12 9 9 13 7 10 9 1 14 15 3 0 9 13 2
17 14 11 7 11 1 9 13 16 11 1 12 1 12 9 9 13 2
11 11 7 11 1 1 12 9 9 13 4 2
23 9 9 1 11 1 0 9 1 0 9 1 9 13 4 15 15 9 1 0 9 0 13 2
36 9 1 15 14 0 13 4 4 16 11 11 1 1 11 1 15 14 15 9 9 13 11 7 0 0 9 13 1 9 1 9 1 9 14 13 2
11 14 0 9 9 13 1 1 10 14 13 2
10 10 9 9 13 14 3 13 4 4 2
23 9 1 1 10 9 13 16 11 1 9 1 9 13 1 1 15 9 1 0 14 13 4 2
22 11 1 0 14 13 1 0 9 0 11 9 1 0 9 14 13 14 13 4 4 4 2
29 9 1 1 0 9 1 1 11 1 11 1 11 11 1 9 1 11 2 11 11 2 11 2 9 1 9 13 4 2
14 11 1 12 9 1 12 2 12 9 1 9 13 4 2
18 9 1 0 13 4 12 9 1 12 9 9 1 10 12 9 9 13 2
7 10 9 11 11 1 13 2
10 11 11 1 0 9 1 9 13 4 2
24 0 9 1 11 1 11 11 11 11 1 0 9 1 1 12 9 1 9 7 9 1 9 13 2
27 9 1 11 1 0 13 1 9 13 11 11 11 2 11 11 2 11 11 11 2 11 11 11 7 11 11 2
48 11 11 2 11 2 1 10 9 1 9 13 4 4 15 13 11 11 11 11 2 11 11 11 2 0 11 7 11 2 11 2 1 9 11 11 11 1 9 11 11 11 2 11 11 7 11 11 2
14 15 1 1 11 11 1 13 10 9 9 1 9 13 2
7 11 1 9 13 4 4 2
18 11 1 0 9 9 1 9 1 9 1 13 12 9 1 10 9 13 2
20 10 9 1 12 9 1 0 9 1 1 9 1 1 10 9 0 13 4 4 2
26 15 1 11 1 11 13 1 9 1 9 1 11 11 1 11 1 9 1 0 13 1 9 1 9 13 2
27 9 9 1 9 1 1 1 13 4 1 11 1 13 16 10 9 1 11 9 11 11 1 9 9 13 4 2
11 11 11 1 0 9 1 9 13 4 4 2
17 11 11 1 13 16 9 1 13 12 9 1 1 9 13 4 4 2
10 9 1 9 1 9 11 1 13 4 2
18 11 1 10 9 1 9 13 16 3 14 9 1 0 9 14 13 4 2
18 11 11 1 13 16 9 1 11 11 11 2 11 2 1 1 13 4 2
9 11 1 1 12 9 0 13 4 2
35 11 9 11 1 11 1 1 13 4 11 2 11 2 11 1 12 0 9 1 9 1 0 13 4 9 9 1 0 9 0 13 1 13 4 2
22 9 9 15 14 13 4 4 16 9 1 13 4 9 1 1 1 9 14 13 4 4 2
27 9 9 9 1 9 9 11 11 11 1 9 1 13 16 13 4 9 9 1 9 1 9 14 13 4 4 2
18 9 9 1 13 4 4 16 13 4 9 11 1 15 9 1 9 13 2
11 11 1 13 16 9 1 9 15 0 13 2
41 11 1 9 1 10 9 15 9 9 1 9 13 4 4 2 1 9 13 15 9 1 9 11 1 1 1 13 4 4 7 15 11 1 11 11 1 9 13 4 4 2
23 9 14 13 1 9 1 12 9 1 13 16 9 9 1 0 9 1 9 13 4 4 4 2
11 15 9 1 1 1 0 9 13 4 4 2
13 9 9 1 9 1 1 15 11 11 13 4 4 2
19 9 1 13 16 11 9 1 0 9 1 9 1 9 14 10 0 13 4 2
14 15 10 9 0 13 1 1 1 14 9 0 13 4 2
38 0 9 9 1 9 9 1 1 9 9 13 4 0 0 11 11 11 1 13 4 16 11 11 1 9 9 9 13 1 13 1 0 9 0 13 4 4 2
13 9 1 9 1 9 13 4 14 15 10 9 13 2
21 15 13 16 11 2 11 7 11 13 11 1 9 9 9 9 13 1 13 4 4 2
16 11 1 13 16 11 9 9 1 1 0 9 0 13 4 4 2
22 11 0 9 13 7 15 11 1 9 9 13 1 13 1 15 9 1 9 13 4 4 2
15 15 13 16 9 9 9 9 9 1 1 3 0 9 13 2
16 15 13 16 15 10 9 13 16 9 9 9 1 9 13 4 2
31 3 1 15 9 1 9 13 4 13 16 15 11 1 15 1 9 13 4 16 15 11 11 11 11 1 11 1 1 9 13 2
15 15 13 16 11 2 11 9 9 1 0 13 4 4 4 2
12 11 11 1 1 15 9 1 0 9 13 4 2
15 15 11 1 9 1 0 0 9 1 0 7 0 9 13 2
13 11 1 13 16 11 1 11 1 0 9 13 4 2
23 15 9 13 4 13 16 11 1 15 9 1 9 0 13 15 9 1 9 1 0 9 13 2
18 11 1 0 9 1 13 9 1 1 11 15 13 0 9 13 4 4 2
21 15 15 13 4 16 11 1 10 9 1 9 9 1 1 0 9 1 9 14 13 2
15 11 1 11 1 9 1 9 1 9 1 15 0 9 13 2
33 0 9 1 3 0 9 9 13 4 11 1 11 1 10 9 1 14 0 13 15 15 11 1 9 9 1 9 13 1 9 13 4 2
25 11 11 11 2 11 2 1 0 9 11 11 1 0 9 1 9 13 9 1 13 1 9 13 4 2
12 9 1 11 9 1 0 11 9 1 13 4 2
38 15 11 1 9 1 1 9 1 9 1 9 9 9 1 9 1 13 16 11 9 1 11 9 1 13 4 9 2 9 13 4 15 11 11 1 13 4 2
19 15 1 1 11 9 1 1 9 11 1 9 1 13 1 9 13 4 4 2
22 9 1 13 16 0 9 13 1 3 9 1 11 1 9 2 1 9 9 13 4 4 2
16 15 9 1 1 0 9 13 1 1 1 15 9 13 13 4 2
13 15 15 14 13 4 16 11 0 9 1 13 4 2
22 15 9 1 13 4 11 9 9 11 11 1 3 15 9 11 1 11 11 11 1 13 2
20 11 1 11 1 9 0 13 1 1 9 9 9 1 0 9 13 1 9 13 2
26 9 11 1 12 9 0 9 9 1 9 1 0 13 1 1 9 10 9 9 1 9 1 0 9 13 2
20 9 9 11 11 11 1 13 16 9 9 9 1 9 1 15 9 14 13 4 2
25 15 13 16 9 0 9 9 1 0 9 13 1 3 14 9 1 9 1 0 0 9 1 3 13 2
40 11 1 13 16 9 9 1 15 9 14 13 15 1 15 0 9 1 0 9 13 1 3 14 9 9 1 1 0 9 1 9 2 9 2 1 3 9 1 13 2
20 15 13 16 9 1 9 1 0 9 0 13 1 1 9 1 9 0 13 4 2
33 15 1 9 9 1 9 1 9 1 9 1 3 13 2 0 9 1 9 1 9 13 7 0 9 1 9 0 13 1 9 13 4 2
29 15 13 16 9 11 1 9 1 0 13 12 0 9 13 2 16 12 12 9 1 15 14 9 1 0 9 14 13 2
23 11 11 2 11 2 11 2 11 2 11 7 11 11 1 12 9 0 9 1 9 14 13 2
20 11 1 13 16 9 1 9 1 0 9 1 9 1 9 13 4 1 9 13 2
31 15 1 0 9 1 0 13 1 1 11 1 12 9 9 1 1 14 0 9 1 9 7 9 1 9 1 9 13 4 4 2
11 15 9 1 9 13 1 9 1 9 13 2
14 11 11 1 1 12 9 9 15 1 9 13 4 4 2
15 15 1 12 9 0 9 9 1 0 9 1 0 13 4 2
13 10 9 1 1 12 9 9 1 0 14 13 4 2
26 11 1 0 9 11 11 1 11 1 9 1 1 1 14 11 7 11 1 0 9 13 1 9 13 4 2
24 15 15 9 1 1 12 9 1 13 4 16 9 10 9 1 0 9 1 9 14 13 4 4 2
14 11 9 1 13 0 9 1 10 9 1 9 13 4 2
12 0 9 1 10 9 1 9 1 9 13 4 2
16 9 1 11 1 15 11 9 1 10 9 13 4 13 4 4 2
14 16 2 15 15 11 1 15 10 9 1 9 13 4 2
37 11 1 1 2 9 1 11 11 9 1 9 1 11 1 0 9 9 1 9 1 14 13 4 1 1 1 11 1 9 1 9 13 4 13 4 4 2
13 11 1 13 4 16 15 3 1 10 9 1 13 2
31 9 1 11 1 15 13 4 13 4 4 4 2 9 13 4 4 7 15 9 1 10 9 11 11 1 10 1 13 4 4 2
9 10 9 15 11 1 14 13 4 2
18 9 1 11 1 13 4 2 13 1 9 1 9 0 9 1 0 13 2
18 11 1 13 13 16 10 9 11 1 9 1 1 1 8 13 4 4 2
23 15 13 4 16 2 11 11 2 1 9 11 11 11 1 11 1 0 9 1 9 1 13 2
16 11 15 9 9 1 9 1 11 1 9 1 9 13 4 4 2
21 9 1 11 9 13 4 4 16 0 9 1 1 0 9 1 13 4 3 0 13 2
16 16 2 9 1 15 15 14 13 4 16 11 10 9 14 13 2
20 11 1 13 4 2 10 9 11 11 1 15 15 11 9 1 8 13 4 4 2
17 15 9 11 1 1 11 11 9 9 1 9 11 11 13 4 4 2
10 15 14 11 1 10 9 0 13 4 2
38 10 9 1 11 0 9 1 9 0 13 4 4 2 15 0 11 2 11 11 11 1 13 4 16 9 1 0 13 1 11 1 0 9 13 4 4 4 2
21 11 9 1 0 9 1 9 1 1 11 1 13 2 9 0 9 13 3 0 13 2
23 11 1 1 11 1 13 2 10 9 15 9 14 13 7 15 9 1 10 9 13 3 13 2
20 11 1 13 4 2 10 9 1 9 15 11 11 11 7 11 9 1 13 4 2
19 15 9 1 9 1 1 1 9 13 1 11 1 9 1 14 9 13 4 2
22 11 1 10 9 1 11 11 1 11 9 1 0 9 7 11 1 8 13 4 13 4 2
27 15 12 9 1 11 7 15 0 9 11 11 1 9 1 11 11 11 1 11 1 1 1 9 13 4 4 2
14 15 1 11 11 10 9 1 9 1 9 13 4 4 2
27 9 1 11 1 9 11 11 1 15 13 13 4 4 2 15 1 0 10 9 1 15 9 14 13 4 4 2
37 11 1 13 4 2 9 1 9 2 9 13 4 9 1 9 2 9 1 9 7 0 13 4 9 1 9 1 1 1 15 15 9 14 13 4 4 2
12 0 9 15 9 13 4 16 10 9 0 13 2
13 10 9 1 12 9 9 1 1 0 13 4 4 2
17 11 1 1 2 15 15 9 1 1 12 9 1 10 9 0 13 2
32 11 1 12 9 1 0 9 9 9 11 11 7 12 0 9 1 9 13 1 9 1 11 11 1 1 1 9 9 1 13 4 2
13 9 1 10 9 1 9 9 1 14 0 13 4 2
12 11 1 9 1 9 1 9 1 0 13 4 2
30 0 13 16 11 11 1 9 1 1 0 9 1 9 7 9 1 0 0 9 1 0 13 1 3 11 9 1 13 4 2
22 9 1 1 9 9 1 9 9 1 9 1 9 7 10 0 9 1 9 9 13 4 2
14 15 1 9 1 9 9 1 15 9 1 13 4 4 2
16 9 1 12 9 1 13 0 9 1 1 11 1 0 13 4 2
19 10 9 1 1 0 9 13 7 9 1 0 13 1 9 0 13 4 4 2
20 9 1 10 9 1 0 9 11 11 2 11 2 9 1 9 1 9 13 4 2
35 12 9 9 1 11 1 15 9 13 4 16 15 9 1 9 1 0 13 7 10 0 9 1 1 0 9 1 1 9 15 9 13 4 4 2
21 9 9 1 13 13 16 9 1 9 1 0 13 1 1 1 15 1 0 9 13 2
18 12 9 3 11 11 11 2 11 2 1 1 12 1 9 0 0 13 2
25 11 9 1 9 11 11 1 13 7 11 2 11 1 9 1 9 0 13 1 9 9 1 13 4 2
19 11 2 11 1 11 11 1 9 13 1 1 9 9 1 9 14 13 4 2
9 7 9 1 15 9 1 13 4 2
22 11 2 11 1 11 11 1 11 11 11 13 1 1 9 1 9 13 1 9 13 4 2
47 11 11 1 9 11 11 11 1 11 11 11 11 1 1 11 11 1 13 4 9 1 9 9 9 1 13 1 9 1 9 13 4 1 3 10 9 1 9 1 11 1 0 9 1 9 13 2
13 16 9 1 13 13 16 15 0 9 1 9 13 2
22 11 1 9 11 11 1 13 13 16 9 1 9 1 9 13 1 9 13 4 4 4 2
10 9 9 1 1 11 1 10 9 13 2
20 15 1 9 9 7 9 1 9 1 15 15 1 9 2 9 13 9 13 4 2
8 9 1 9 1 9 13 4 2
16 9 1 9 11 11 1 9 0 13 1 9 13 7 0 13 2
24 11 11 11 11 1 15 9 1 13 16 9 1 9 13 1 15 14 9 1 9 1 13 4 2
10 15 13 16 0 9 1 9 13 4 2
38 9 1 12 0 0 0 0 7 0 9 1 9 1 11 11 1 11 1 9 9 1 9 0 13 7 15 9 1 9 1 9 1 15 9 0 13 4 2
60 9 9 11 11 11 2 9 11 11 11 2 9 11 11 11 2 9 11 11 2 9 11 11 11 2 9 11 11 7 9 11 11 11 1 12 0 9 1 0 9 1 1 1 12 9 1 9 1 9 1 9 13 1 9 1 15 9 0 13 2
40 9 9 1 1 12 11 11 11 11 11 11 11 1 9 1 9 9 1 1 0 9 1 3 14 9 9 13 4 1 1 11 11 11 11 13 1 9 13 4 2
27 9 1 13 16 0 2 0 9 0 13 1 1 1 9 9 1 12 12 1 10 9 15 14 0 13 4 2
40 7 0 0 0 7 0 9 1 13 13 16 9 9 1 9 9 1 14 0 13 4 4 4 7 9 9 1 13 13 16 9 1 9 9 1 0 13 4 4 2
30 11 11 11 1 0 9 9 11 11 1 11 11 11 2 11 2 1 15 9 1 9 1 3 14 9 1 9 13 4 2
17 15 13 13 16 11 11 1 0 9 9 1 1 15 9 13 4 2
32 0 13 16 9 7 0 9 1 9 14 13 1 9 1 15 0 13 4 1 0 11 11 1 1 9 1 0 13 4 4 4 2
31 11 1 13 13 16 9 9 1 9 1 9 9 1 9 1 1 11 11 1 11 11 1 13 4 9 9 1 9 14 13 2
18 11 1 9 11 11 11 1 9 11 11 1 9 13 15 12 9 13 2
23 11 1 15 11 11 11 7 11 11 1 1 1 13 4 9 1 9 13 1 9 13 4 2
16 0 13 16 11 1 15 0 9 1 9 9 1 9 13 4 2
22 9 9 1 15 12 9 1 0 13 4 1 3 11 11 1 9 1 0 13 4 4 2
46 9 9 11 1 15 9 11 11 1 9 1 11 15 13 16 15 9 1 0 9 13 4 2 7 9 2 9 11 11 15 9 11 1 1 11 11 11 13 1 1 0 13 4 4 4 2
22 11 1 9 2 9 11 1 9 1 1 11 1 1 9 13 1 9 11 1 14 13 2
29 11 1 9 11 0 13 7 9 1 15 9 1 9 1 1 9 2 9 1 11 9 1 11 11 11 0 13 4 2
7 11 10 9 1 0 13 2
18 7 9 1 9 1 9 1 15 10 9 15 1 9 1 9 13 4 2
12 9 14 1 9 11 11 1 15 0 13 4 2
15 11 1 9 1 11 11 11 13 1 1 0 13 4 4 2
21 11 11 1 10 9 1 0 15 9 1 12 9 1 11 11 11 1 9 13 4 2
22 0 9 1 13 4 10 9 1 12 0 9 13 2 15 9 1 0 9 13 4 4 2
12 10 9 1 3 11 1 9 1 13 4 4 2
25 11 11 11 1 9 12 9 0 13 7 3 10 9 1 9 1 9 1 15 3 14 0 13 4 2
13 11 11 1 10 9 1 9 1 10 9 13 4 2
20 15 10 9 1 15 11 11 11 0 13 2 15 0 9 1 9 13 4 4 2
15 16 2 0 9 1 9 2 9 1 9 0 13 4 4 2
29 15 15 9 1 9 11 11 11 1 13 4 11 13 1 0 13 4 4 2 15 14 15 1 3 15 9 14 13 2
41 0 11 1 11 11 0 11 1 9 9 1 9 13 1 9 1 9 1 1 9 1 0 9 9 11 11 11 11 1 9 1 12 0 9 1 9 1 9 13 4 2
15 9 1 15 9 13 1 1 12 9 1 9 13 4 4 2
25 11 1 1 11 11 1 0 9 0 9 9 11 11 11 11 7 11 11 1 9 9 1 9 13 2
22 11 11 11 11 11 1 1 9 9 1 9 7 15 1 13 4 9 9 1 9 13 2
21 15 1 9 9 1 0 9 7 9 9 1 9 1 10 0 13 1 9 14 13 2
28 0 13 16 11 11 0 11 1 11 9 1 0 11 11 1 11 11 0 12 9 1 13 1 9 13 4 4 2
9 10 9 9 1 12 9 0 13 2
28 9 7 9 9 1 1 15 1 12 9 1 13 4 4 4 2 7 12 9 1 13 4 1 9 13 4 4 2
9 15 1 12 9 0 13 4 4 2
23 11 1 11 11 11 0 11 9 11 9 1 13 0 9 1 13 12 9 1 13 4 4 2
47 11 9 1 9 1 12 11 9 1 12 9 1 11 11 11 11 11 1 13 11 11 1 13 11 9 1 13 9 1 1 15 3 0 13 7 0 9 1 9 9 9 13 1 9 13 4 2
37 0 9 11 11 11 1 9 1 11 1 13 13 10 9 1 11 11 11 2 11 11 11 2 11 11 11 7 11 11 1 11 0 11 9 0 13 2
42 3 1 12 9 9 1 10 9 1 9 13 16 9 9 1 9 11 11 11 11 1 12 0 9 11 11 11 1 9 13 7 15 11 1 9 1 9 1 3 9 13 2
23 15 13 16 9 9 1 9 13 4 7 11 1 13 1 3 9 13 4 7 9 13 4 2
25 15 11 11 1 9 13 16 11 11 1 13 9 1 0 13 0 9 1 0 7 0 9 13 4 2
38 11 1 9 1 11 1 9 1 0 9 13 4 10 9 1 13 16 11 1 10 0 9 1 0 9 1 3 13 4 16 12 9 1 9 13 4 4 2
23 15 11 11 9 11 11 11 1 10 9 1 11 1 1 15 9 1 9 13 1 9 13 2
45 11 9 1 11 1 9 1 9 13 4 13 16 10 9 15 11 11 1 0 13 7 15 1 15 9 13 1 1 15 1 9 13 4 12 9 1 1 0 9 1 13 9 13 4 2
23 11 11 1 11 7 11 11 2 11 2 1 3 11 11 11 2 11 2 1 9 13 4 2
29 9 15 11 1 9 9 11 11 1 1 9 1 1 9 1 9 13 4 11 11 11 11 11 11 1 10 9 13 2
23 10 9 1 1 1 15 13 16 9 1 13 1 10 9 1 1 11 1 9 13 4 4 2
29 11 1 13 16 9 1 1 11 1 9 1 3 9 13 4 4 7 15 3 13 1 10 9 1 9 13 4 4 2
31 10 9 1 11 1 11 1 0 9 1 15 9 1 9 1 13 1 1 13 4 4 0 2 0 9 9 1 14 9 13 2
19 15 13 16 11 1 9 1 9 1 9 13 4 16 0 9 15 13 4 2
20 0 13 16 15 1 11 1 0 9 9 7 9 1 9 1 1 13 4 4 2
23 15 1 11 1 0 9 2 9 9 7 9 1 9 1 11 1 9 13 1 9 14 13 2
25 9 1 1 11 1 11 1 9 1 11 1 9 13 7 9 1 13 0 9 9 1 9 1 13 2
31 10 9 1 12 9 1 11 11 11 2 11 2 9 1 0 9 9 1 11 11 1 9 1 0 13 4 1 9 0 13 2
16 9 1 11 11 11 1 11 11 11 1 1 1 0 13 4 2
15 15 9 9 1 0 0 9 1 3 13 1 9 13 4 2
14 11 11 11 1 9 1 1 9 1 10 9 13 4 2
37 11 11 11 1 9 9 11 1 9 9 1 12 9 1 9 1 13 16 11 11 11 1 1 1 9 0 9 7 9 1 0 9 1 9 13 4 2
34 15 13 16 9 1 9 9 1 1 1 9 13 4 9 11 11 11 1 0 9 1 9 1 0 9 1 9 13 1 9 13 4 4 2
32 11 11 1 11 11 11 2 11 2 1 1 0 13 4 4 7 0 9 1 13 15 9 9 1 0 9 13 1 9 13 4 2
9 15 9 11 11 1 13 4 4 2
24 10 9 1 11 11 1 11 11 11 2 11 2 1 9 1 1 12 9 9 0 13 4 4 2
16 11 11 1 9 1 1 11 1 9 1 10 9 13 4 4 2
20 0 9 1 11 11 2 11 2 1 9 9 1 10 9 1 9 13 4 4 2
23 11 11 11 11 10 9 1 9 1 9 13 4 4 7 10 9 1 15 0 13 4 4 2
24 15 15 1 9 13 1 1 9 1 9 11 11 1 9 1 9 1 12 9 9 13 4 4 2
15 15 9 7 0 9 1 9 1 14 0 13 4 4 4 2
11 9 1 11 11 11 1 15 9 13 4 2
17 9 12 9 1 1 9 1 9 7 9 1 9 2 9 0 13 2
17 0 0 9 1 1 14 11 11 7 11 11 13 9 1 0 13 2
22 9 1 1 11 11 11 1 1 9 13 4 9 1 9 1 13 9 0 13 4 4 2
33 9 1 13 13 16 9 1 9 14 0 13 7 9 1 14 9 14 13 7 15 9 1 0 13 4 2 15 9 1 9 14 13 2
59 10 9 13 16 0 9 11 11 1 9 1 13 11 11 11 2 11 2 1 9 1 11 11 11 1 9 1 9 0 13 4 4 7 11 11 1 15 1 9 13 4 16 10 9 9 14 13 4 4 7 15 9 14 0 14 13 4 4 2
12 15 15 3 14 9 1 0 13 1 13 4 2
11 9 1 12 3 0 9 13 11 11 11 2
70 10 9 1 0 9 9 1 9 1 1 13 4 4 7 13 4 4 16 11 11 11 11 11 11 1 0 9 1 9 1 0 14 13 4 4 10 9 15 11 9 7 11 11 1 12 2 12 0 9 1 10 9 1 0 9 0 13 1 1 11 11 11 1 9 13 1 9 13 4 2
18 10 12 9 1 9 13 1 3 15 9 1 1 14 9 9 0 13 2
14 11 9 11 11 1 11 1 9 13 4 9 13 4 2
31 7 0 11 11 11 11 1 11 9 11 11 1 13 4 13 13 4 16 11 1 1 9 9 15 10 9 1 13 13 4 2
22 11 1 9 1 9 1 9 13 1 1 11 1 0 11 11 11 11 1 9 1 13 2
23 11 1 15 9 1 10 15 13 4 15 11 1 13 1 3 11 1 9 1 9 14 13 2
28 11 9 1 14 9 2 9 1 11 13 7 11 11 1 1 1 15 9 14 13 1 11 1 0 9 13 4 2
12 9 13 11 9 15 11 13 15 11 15 13 2
17 7 15 15 1 13 1 3 10 9 1 15 13 1 9 14 13 2
32 9 9 1 1 11 11 1 1 15 0 13 4 16 11 1 1 9 9 1 11 1 9 1 9 3 11 1 9 1 13 4 2
26 11 1 9 1 11 9 1 9 1 9 13 0 13 4 16 11 9 1 9 15 11 0 13 4 4 2
24 9 1 13 4 4 16 11 9 1 11 1 11 1 1 15 0 9 1 13 4 1 9 13 2
15 9 9 1 1 11 1 15 10 9 1 9 13 4 4 2
54 11 11 1 13 1 0 13 4 0 11 11 7 9 1 9 11 11 1 11 1 13 16 11 9 14 11 2 11 11 11 1 0 13 1 9 1 13 7 9 1 11 9 1 10 9 1 3 13 1 9 1 9 13 2
27 11 2 11 1 9 9 11 1 0 13 4 4 4 7 9 10 9 1 0 9 1 9 14 13 4 4 2
14 11 1 10 9 1 0 13 1 1 9 0 13 4 2
13 11 11 1 15 1 1 0 7 0 9 13 4 2
41 11 1 13 16 9 10 9 1 11 11 11 11 11 11 1 0 9 13 1 9 1 0 13 15 14 11 2 11 1 1 9 11 1 0 9 9 1 9 13 4 2
23 9 1 13 4 4 16 11 1 9 0 13 7 11 9 1 15 0 9 1 9 14 13 2
23 11 1 13 16 10 9 11 9 1 11 9 1 14 9 11 13 1 9 13 15 0 13 2
27 11 1 11 1 11 1 0 9 7 0 9 1 9 1 0 13 4 13 2 11 9 1 9 0 13 4 2
11 15 11 1 0 9 13 1 14 9 13 2
32 9 9 1 11 11 1 12 9 1 11 11 11 1 9 13 4 0 9 1 9 1 9 1 12 9 1 9 1 9 13 4 2
11 10 9 9 2 9 1 0 9 1 13 2
32 9 1 13 16 9 16 0 12 9 1 9 1 9 1 0 13 16 15 9 15 14 13 16 15 15 9 1 0 14 13 4 2
16 15 0 9 1 13 4 1 0 9 1 13 13 0 14 13 2
32 11 1 15 9 1 9 1 11 11 11 1 10 9 0 13 4 2 15 15 9 11 1 13 4 1 3 9 1 9 13 4 2
20 10 9 1 0 13 4 4 16 9 1 10 9 13 4 1 1 1 13 4 2
37 15 1 9 9 9 1 11 11 11 1 15 9 1 9 1 9 13 4 16 15 11 9 1 9 7 9 1 13 9 1 1 9 9 1 9 13 2
12 9 1 15 1 9 9 9 1 9 13 4 2
15 9 1 10 9 0 13 4 9 1 9 1 0 9 13 2
23 9 1 11 2 11 7 11 1 0 9 1 0 9 9 13 1 9 13 0 9 13 4 2
18 11 11 11 1 9 1 9 15 13 9 1 9 1 10 9 13 4 2
21 0 13 16 10 9 1 10 9 11 1 13 4 4 4 7 11 1 3 13 4 2
27 11 1 1 15 9 13 4 4 7 0 9 1 0 9 1 9 1 1 9 1 15 9 0 13 4 4 2
17 11 11 11 11 1 15 10 9 9 1 1 13 1 9 13 4 2
48 15 10 9 13 1 10 9 7 15 1 9 7 9 9 1 1 0 9 1 1 10 0 9 1 1 10 9 1 1 0 13 4 10 14 9 15 9 10 9 9 2 9 2 1 1 1 13 2
9 16 10 9 0 13 10 9 13 2
21 9 1 13 13 16 15 13 4 1 10 9 0 7 0 9 1 10 0 13 4 2
27 15 15 0 9 1 0 13 7 0 0 9 1 1 15 13 7 9 1 1 15 0 13 1 10 9 13 2
11 15 1 0 0 9 1 0 14 13 4 2
22 9 1 1 15 9 1 9 12 9 1 1 13 7 15 9 11 2 11 1 0 13 2
17 0 9 15 9 13 7 3 3 1 12 9 1 1 15 9 13 2
40 11 11 11 11 2 11 11 11 11 11 2 1 9 11 11 11 1 13 4 16 9 11 11 11 2 11 2 1 0 14 13 2 7 9 1 3 0 13 4 2
14 11 1 9 11 2 11 1 9 1 0 13 4 4 2
28 11 1 11 11 11 11 11 11 1 0 12 9 1 11 1 13 16 2 11 1 0 13 4 1 15 9 14 13
17 11 1 13 16 11 1 9 1 1 9 1 0 9 13 4 4 2
23 15 3 13 16 11 11 1 9 1 0 13 4 16 0 9 1 1 1 9 13 4 4 2
8 9 10 0 9 1 9 13 2
37 9 1 9 1 13 16 11 11 11 2 11 2 1 0 13 4 1 11 11 1 10 9 1 10 0 9 1 1 1 9 13 1 9 13 4 4 2
21 15 13 16 0 10 9 1 10 9 9 1 1 1 0 9 1 9 13 4 4 2
14 0 0 9 1 9 1 1 15 3 14 12 9 13 2
17 11 1 13 16 9 14 1 0 9 1 1 0 9 9 10 13 2
10 15 11 1 14 15 14 13 4 4 2
35 15 13 16 10 9 11 11 1 1 9 9 14 12 12 12 12 9 13 2 7 0 9 10 9 1 1 10 9 12 12 12 12 9 13 2
22 11 11 1 11 1 9 7 9 7 0 0 9 9 1 9 13 4 12 9 1 13 2
31 9 1 0 13 4 16 15 15 14 0 9 0 0 9 7 9 1 9 9 9 2 9 2 13 1 1 0 14 13 4 2
32 9 11 11 11 7 9 11 11 11 1 9 1 9 1 13 16 10 15 14 9 9 1 13 1 9 15 15 9 1 14 13 2
30 9 1 0 13 16 11 2 11 1 1 0 9 1 9 1 1 0 9 13 1 1 15 9 1 0 14 13 4 4 2
17 0 13 16 9 1 11 1 15 10 9 1 9 13 1 9 13 2
37 11 1 12 9 9 1 9 1 0 12 9 9 1 9 13 4 4 16 11 11 11 11 11 11 11 1 9 9 13 1 9 9 1 0 13 4 2
24 10 9 1 9 13 4 4 16 11 11 1 0 0 9 1 9 0 13 1 9 13 4 4 2
18 9 1 9 1 9 11 11 1 9 9 1 9 0 13 1 13 4 2
23 11 11 11 11 11 11 11 1 13 16 15 15 1 0 9 9 1 12 0 9 0 13 2
23 11 1 9 1 9 1 11 1 13 16 11 1 11 9 9 1 9 1 9 13 4 4 2
21 15 11 9 1 9 9 1 9 1 9 1 0 0 9 1 9 1 9 14 13 2
36 9 1 0 9 1 9 1 9 13 4 15 13 13 16 11 9 14 15 9 9 7 9 13 1 9 1 9 1 9 1 14 9 13 4 4 2
28 11 1 11 11 11 1 13 13 16 3 0 9 1 12 13 1 1 11 1 0 9 0 14 13 4 4 4 2
13 15 13 16 11 9 1 9 1 9 13 4 4 2
29 9 9 7 9 9 1 9 1 3 2 3 9 13 1 0 11 11 1 11 11 1 9 1 9 13 1 9 13 2
17 15 9 9 7 11 11 9 9 9 1 0 9 13 1 9 13 2
23 11 1 11 11 1 9 13 16 11 9 1 9 1 1 9 7 9 1 1 1 9 13 2
11 11 1 11 11 1 9 13 1 9 13 2
23 11 1 11 11 11 1 13 16 9 9 1 9 13 14 15 0 9 1 1 13 4 4 2
12 15 9 9 1 9 1 9 14 0 13 4 2
13 15 11 11 1 1 0 0 9 1 9 14 13 2
21 11 1 11 11 1 0 9 9 1 9 1 13 1 1 1 0 9 1 9 13 2
19 11 1 11 11 1 9 1 9 1 9 14 13 1 1 9 1 9 13 2
22 11 1 11 11 1 11 11 11 1 9 0 14 13 1 1 0 11 9 1 9 13 2
18 11 1 11 11 1 12 9 1 9 1 12 9 9 13 1 9 13 2
10 9 9 9 1 11 1 9 0 13 2
24 11 1 13 9 1 1 11 1 12 9 1 9 0 13 2 7 11 1 9 1 12 9 13 2
22 3 11 11 1 11 2 11 9 1 0 9 13 4 12 9 1 1 12 1 9 13 2
22 9 9 1 11 9 1 9 13 1 1 11 11 1 10 12 9 1 14 9 13 4 2
10 9 9 1 1 11 1 9 13 4 2
16 11 1 11 1 11 11 7 11 11 9 1 15 9 3 13 2
17 11 2 11 1 11 11 11 11 1 11 9 1 9 0 13 4 2
11 15 12 9 1 9 1 9 1 9 13 2
24 11 1 13 9 1 1 11 1 11 1 11 11 11 1 11 1 11 11 1 12 11 1 13 2
18 11 1 11 1 11 11 1 11 1 11 11 1 12 9 1 0 13 2
11 3 11 1 11 9 1 9 3 13 4 2
27 11 11 11 11 1 9 1 0 13 9 1 11 1 11 11 11 1 11 1 11 11 1 12 9 1 13 2
18 11 1 11 1 11 11 1 11 1 11 11 1 12 9 1 0 13 2
39 11 9 1 10 9 1 0 11 11 11 15 9 13 1 0 13 2 7 9 1 11 9 1 11 1 11 11 1 11 1 9 11 11 1 12 9 1 13 2
20 11 1 11 1 11 11 1 11 1 9 11 11 11 1 12 9 1 0 13 2
17 11 1 11 1 11 11 1 11 1 11 11 1 12 9 1 13 2
22 11 1 11 1 11 11 1 11 1 11 11 11 1 0 9 1 12 9 1 0 13 2
20 10 9 11 1 11 1 11 1 11 1 11 11 1 12 9 1 9 1 13 2
19 11 1 11 1 11 11 1 11 1 11 11 11 1 12 9 1 0 13 2
21 3 11 11 1 11 1 11 11 1 11 1 11 11 14 11 1 12 9 1 13 2
9 11 1 10 9 11 1 13 4 2
17 11 11 11 1 0 9 11 11 11 1 0 9 1 9 13 4 2
29 11 2 11 1 11 11 9 1 11 11 11 11 1 15 0 9 11 9 11 11 11 1 12 9 1 9 1 13 2
19 11 11 1 11 1 12 9 1 11 9 1 11 11 9 1 9 0 13 2
29 11 1 11 11 9 1 9 1 11 1 11 11 2 11 2 1 15 0 9 11 1 11 11 1 12 9 1 13 2
19 11 11 1 0 11 1 9 13 4 11 1 11 11 9 1 9 0 13 2
9 7 11 9 11 1 9 1 13 2
22 11 11 1 11 9 11 11 11 11 1 13 2 7 11 9 1 11 1 9 3 13 2
21 11 11 1 0 11 11 1 11 1 11 2 11 7 11 9 1 15 9 0 13 2
19 11 1 11 1 9 1 9 13 4 11 1 11 11 9 1 9 0 13 2
24 11 1 0 9 11 1 12 9 1 9 0 13 2 7 11 11 11 1 15 12 9 13 4 2
32 11 11 11 1 3 3 9 13 7 9 1 9 1 9 1 12 9 9 1 9 13 11 11 1 12 9 3 9 13 4 4 2
33 11 1 11 1 12 9 3 9 13 1 3 9 1 15 11 11 1 9 1 13 1 9 13 4 2 16 11 9 15 15 14 13 2
14 9 9 11 11 1 9 1 9 1 1 11 13 4 2
5 15 11 13 13 4
22 15 1 9 1 11 9 1 9 1 11 1 0 13 4 4 9 1 1 1 9 13 2
6 11 11 1 0 13 2
24 9 1 1 14 11 1 12 9 9 1 1 9 13 4 13 16 9 3 15 1 13 4 4 2
21 2 15 1 9 1 9 1 13 16 11 0 9 7 9 1 1 9 13 4 4 2
24 15 9 1 9 13 16 15 11 1 9 1 9 0 13 7 9 1 9 0 13 1 9 13 2
16 11 9 1 14 12 9 13 7 10 9 15 9 13 13 4 2
34 9 1 11 9 1 15 14 13 16 15 11 1 1 9 1 0 14 13 7 15 9 1 9 2 9 0 13 1 9 1 9 13 4 2
32 9 1 9 1 15 14 13 16 15 10 9 13 16 11 1 1 10 9 1 1 9 14 13 4 2 15 9 9 13 4 4 2
26 11 11 11 1 9 13 4 11 11 1 11 11 1 0 9 9 1 1 0 9 13 1 9 13 4 2
18 0 13 16 11 11 11 11 9 1 12 9 1 10 1 9 0 13 2
18 11 11 1 9 1 15 1 0 9 1 9 1 13 11 9 1 13 2
34 11 9 1 9 1 11 1 9 1 9 9 1 9 1 2 0 0 9 2 7 2 9 2 1 0 0 9 1 9 9 13 13 4 2
29 9 1 9 1 11 9 11 11 1 13 16 9 1 9 9 9 1 1 9 0 13 15 15 9 1 13 13 4 2
29 10 9 11 1 9 9 1 9 1 0 9 13 1 11 1 10 9 13 4 7 15 12 9 1 9 0 13 4 2
19 11 1 1 0 9 1 1 11 1 0 9 1 11 1 9 13 4 4 2
34 11 11 1 9 9 9 11 11 11 1 11 9 9 7 9 11 11 1 11 0 11 9 1 9 1 9 1 9 1 1 9 9 13 2
26 11 1 11 1 11 1 11 1 0 9 9 11 1 9 9 11 1 1 13 1 9 1 1 9 13 2
28 12 9 1 1 14 12 9 1 9 1 1 11 9 7 11 9 9 1 12 9 1 1 9 9 1 9 13 2
17 11 13 1 3 11 7 11 1 9 1 13 16 15 9 0 13 2
23 15 13 16 10 0 7 0 2 0 9 1 13 4 11 7 11 1 1 0 9 13 4 2
11 12 9 1 1 15 9 1 9 14 13 2
25 11 1 0 11 11 11 7 11 11 11 11 11 11 2 11 11 1 0 13 1 9 1 14 13 2
16 16 9 9 0 13 4 1 1 1 15 9 13 4 4 4 2
20 15 1 11 1 11 9 9 0 13 1 1 0 9 13 1 9 13 4 4 2
25 9 1 11 11 11 11 11 1 13 16 15 15 1 9 9 0 13 1 1 10 15 9 14 13 2
19 15 13 16 15 10 13 4 4 2 15 15 1 0 9 1 9 13 4 2
20 7 12 9 1 9 13 1 3 11 7 11 1 9 7 9 1 9 13 4 2
24 15 13 16 9 0 13 1 1 11 11 1 13 4 9 1 13 4 9 9 14 13 4 4 2
17 15 1 0 13 4 1 11 1 9 14 11 11 1 0 13 4 2
16 15 13 16 11 2 11 11 9 1 1 9 1 9 14 13 2
15 11 1 11 7 11 1 13 4 16 11 15 0 13 4 2
18 15 0 9 1 0 13 1 1 0 9 1 1 1 9 1 9 13 2
18 9 9 9 1 11 9 1 9 0 9 1 11 11 1 9 13 4 2
19 11 9 1 15 9 1 12 9 1 1 9 9 13 1 9 13 4 4 2
34 9 9 9 1 9 2 11 2 1 15 9 1 13 16 11 9 2 0 2 9 2 11 1 0 13 1 14 12 12 9 0 13 4 2
22 2 11 2 1 9 13 4 11 11 11 1 13 16 9 1 9 1 11 1 9 13 2
21 0 13 16 11 9 1 9 0 13 1 3 14 10 9 11 11 1 0 13 4 2
40 11 9 1 11 1 11 11 1 11 11 11 1 11 9 1 0 9 1 9 1 11 11 11 11 2 11 2 1 9 11 11 1 12 0 9 9 1 9 13 2
17 11 1 11 1 9 1 10 9 1 13 9 1 13 1 9 13 2
25 15 13 16 9 1 13 4 4 9 1 0 13 1 1 0 9 1 9 1 9 1 9 13 4 2
18 7 11 1 0 9 1 1 15 0 9 1 14 0 13 1 9 13 2
18 7 11 1 9 1 13 0 11 11 1 9 1 9 15 0 14 13 2
16 3 2 11 1 0 9 1 15 15 1 15 9 13 0 13 2
36 11 11 1 11 1 9 1 11 1 0 9 1 11 9 11 11 7 9 11 11 11 1 11 9 1 13 11 11 11 1 12 9 0 9 13 2
17 11 1 11 1 0 9 1 13 16 11 1 9 9 1 13 4 2
18 15 9 1 0 7 15 14 0 13 1 9 1 0 13 1 9 13 2
26 9 1 11 1 1 11 11 11 11 2 0 9 9 11 11 11 7 9 9 11 11 11 1 9 13 2
23 9 1 11 9 1 11 1 9 11 11 7 11 1 9 9 11 11 11 11 14 0 13 2
35 11 1 9 9 11 11 1 9 1 1 9 1 13 16 11 10 9 9 1 10 9 7 9 1 9 13 4 15 9 1 9 3 13 4 2
21 7 11 1 9 1 13 16 9 0 15 13 15 15 0 9 1 14 0 13 4 2
14 15 9 1 9 1 9 9 1 1 9 2 9 13 2
21 11 9 1 11 11 1 11 1 1 0 9 11 11 1 11 11 1 9 13 4 2
8 10 9 15 11 11 1 13 2
10 16 15 15 0 9 14 13 4 4 2
26 11 11 1 0 9 1 9 11 11 11 11 1 11 1 11 11 11 1 9 13 1 0 9 13 4 2
11 15 13 13 16 10 9 1 15 9 14 2
30 7 11 11 11 1 9 1 11 11 1 0 9 1 11 11 11 1 9 13 1 9 13 1 1 9 11 1 13 4 2
27 11 9 1 9 9 13 11 11 1 9 1 11 11 1 11 11 1 9 1 9 13 1 9 13 4 4 2
28 0 13 16 15 1 9 1 10 9 13 1 9 1 11 11 1 11 11 1 0 9 1 9 0 13 4 4 2
35 9 11 11 7 9 11 11 11 1 9 1 13 16 16 11 11 0 9 9 1 1 9 13 4 16 10 9 9 9 1 9 13 4 4 2
35 9 1 0 13 16 9 1 9 1 9 14 13 1 9 1 10 9 14 13 4 4 16 9 9 1 9 2 9 2 1 9 13 4 4 2
23 0 13 16 11 11 1 9 14 13 1 3 11 1 11 11 1 11 11 1 9 13 4 2
33 9 1 0 9 1 10 9 13 1 9 1 9 1 11 11 1 11 7 15 0 9 11 11 1 0 9 1 9 0 13 4 4 2
15 9 1 10 9 1 9 1 1 12 9 1 9 13 4 2
15 16 9 1 11 1 9 11 11 1 0 9 13 4 4 2
19 11 15 12 9 1 9 1 12 0 9 1 15 9 1 9 13 4 4 2
28 15 1 9 1 0 9 1 10 9 0 13 1 9 13 7 15 1 11 11 11 1 1 9 0 13 4 4 2
33 11 9 1 11 11 11 1 1 1 0 9 1 1 11 1 1 12 12 1 9 13 15 15 9 1 0 9 1 12 9 10 13 2
18 9 1 13 0 2 0 9 1 12 9 1 12 9 1 9 13 4 2
31 0 9 1 1 2 11 9 1 11 9 1 11 9 1 11 1 9 9 9 1 1 13 9 1 12 0 9 13 4 4 2
21 13 4 9 1 1 1 12 9 2 9 9 2 12 9 7 12 9 0 13 4 2
32 3 12 0 9 1 11 9 1 14 11 9 1 9 1 0 0 9 1 9 11 11 11 14 11 1 9 13 4 9 13 4 2
17 11 11 11 1 0 9 1 9 1 13 4 12 9 1 13 4 2
24 15 1 14 11 9 1 0 9 1 0 9 9 9 9 1 9 1 9 13 4 9 13 4 2
18 11 11 11 1 15 9 13 4 2 15 15 15 9 1 13 4 4 2
17 11 11 1 9 9 1 9 1 9 9 1 9 1 9 13 4 2
23 11 11 11 11 1 1 9 9 1 1 14 0 9 1 9 1 9 1 9 13 4 4 2
26 9 9 9 1 1 0 9 0 13 16 9 1 9 1 1 10 9 1 9 1 9 0 13 4 4 2
16 9 1 10 9 1 11 11 11 11 1 9 1 9 13 4 2
31 10 9 1 13 1 3 9 1 9 15 13 16 11 11 11 11 1 9 1 9 9 1 1 14 12 0 9 0 13 4 2
13 15 1 14 9 9 1 10 9 1 9 13 4 2
26 3 0 9 1 9 1 13 9 7 0 9 1 10 9 1 9 13 1 1 9 1 10 9 13 4 2
20 9 1 1 9 1 10 9 13 15 1 10 9 1 0 9 14 13 4 4 2
28 10 9 1 9 1 1 11 11 11 11 1 9 1 14 0 9 0 13 4 7 9 1 9 14 9 13 4 2
14 3 9 1 9 9 1 13 15 13 1 9 13 4 2
14 15 1 11 11 11 1 1 14 9 1 0 13 4 2
14 16 0 9 1 15 14 9 1 1 0 9 0 13 2
22 3 9 1 0 12 9 1 1 10 9 1 1 12 12 9 1 9 1 9 13 4 2
9 10 9 1 12 9 9 0 13 2
31 11 11 1 13 13 16 10 9 1 13 4 1 9 1 9 9 1 10 9 13 7 0 9 13 1 10 9 10 0 13 2
16 10 9 1 0 9 9 1 9 9 13 12 12 9 13 4 2
26 15 1 14 15 0 7 0 9 1 12 12 9 1 9 13 7 9 1 0 9 14 12 12 9 13 2
12 10 0 0 9 1 10 9 1 1 13 4 2
22 12 0 9 1 11 1 11 9 11 11 1 0 9 1 9 11 11 1 0 13 4 2
30 0 13 16 10 9 1 11 1 11 11 11 11 1 11 1 9 13 4 11 11 1 15 1 0 13 1 9 13 4 2
34 15 13 4 4 16 11 11 11 1 1 15 0 9 0 9 1 0 13 1 1 11 11 11 11 1 1 15 15 14 9 13 4 4 2
35 10 9 1 9 1 9 11 11 11 7 11 11 1 11 1 9 11 1 11 1 9 1 1 13 16 15 1 9 1 10 9 13 4 4 2
7 15 9 1 9 13 4 2
25 9 9 11 1 11 1 12 9 1 11 1 1 12 9 9 1 13 9 11 9 10 0 13 4 2
26 9 1 13 13 16 10 9 1 9 13 1 0 9 7 0 9 9 1 10 14 10 12 9 10 13 2
23 11 11 11 2 11 2 1 12 0 9 1 13 16 9 15 14 0 9 9 13 4 4 2
9 9 9 1 11 1 9 13 4 2
7 10 9 11 1 14 13 2
20 11 1 9 11 11 11 1 13 16 9 1 9 13 1 15 10 9 10 13 2
24 15 0 9 1 13 4 9 13 4 4 7 10 14 10 12 9 1 9 1 9 13 4 4 2
10 3 10 9 1 9 13 9 13 4 2
8 15 1 15 9 13 4 4 2
11 9 1 9 1 0 9 13 4 4 4 2
14 10 9 1 9 13 1 1 11 1 12 9 13 4 2
17 12 0 9 11 0 11 11 11 11 11 11 11 1 13 4 4 2
15 10 9 1 10 9 1 9 1 9 13 1 0 9 13 2
20 10 0 9 9 7 9 9 1 9 13 1 9 1 13 1 1 13 4 4 2
16 12 9 11 1 14 9 1 13 4 7 15 9 1 9 13 2
24 11 1 9 11 11 1 13 16 12 0 9 1 9 13 1 1 13 4 4 9 1 9 13 2
17 15 13 16 15 12 9 9 13 1 1 11 11 11 1 9 13 2
20 15 1 3 1 12 9 1 10 0 9 1 9 1 9 1 9 13 4 4 2
9 10 9 1 12 9 9 13 4 2
11 3 9 1 9 1 14 9 13 4 4 2
9 15 9 1 9 10 13 4 4 2
16 0 9 1 9 1 9 7 9 1 9 1 14 9 13 4 2
20 2 11 2 1 9 2 11 11 2 1 15 11 11 1 9 1 8 13 4 2
34 11 1 9 2 11 11 11 11 11 2 1 11 1 9 13 4 16 10 9 2 11 2 9 1 13 4 15 12 0 9 1 9 13 2
18 10 9 1 9 11 11 11 1 11 11 11 1 12 9 0 13 4 2
20 11 1 9 13 4 16 2 11 11 2 15 9 9 2 11 2 1 0 13 2
14 2 11 2 1 11 11 9 11 11 1 9 13 4 2
39 11 11 1 2 11 2 1 10 9 1 9 1 9 13 1 9 13 4 9 1 10 0 9 9 1 15 9 7 9 11 1 7 15 1 0 13 1 13 2
28 9 13 9 1 9 13 1 9 9 1 9 13 4 9 1 0 9 1 11 1 0 9 1 9 9 13 4 2
18 10 9 9 1 9 12 9 1 1 12 9 9 9 1 1 0 13 2
26 11 1 11 11 11 1 9 1 10 0 9 1 11 11 9 1 0 9 1 1 10 9 1 9 13 2
25 9 11 11 11 1 11 11 7 11 1 11 11 11 11 7 11 1 11 11 9 1 1 0 13 2
9 0 0 9 1 14 3 13 4 2
8 9 1 11 1 14 9 13 2
17 9 1 11 11 9 12 12 9 1 9 9 1 15 9 13 4 2
19 10 9 1 11 11 11 11 1 11 11 1 12 9 1 14 13 4 4 2
16 11 9 1 9 13 9 1 9 0 9 1 0 9 1 13 2
19 9 1 1 11 11 9 1 9 1 13 1 0 9 1 9 13 4 4 2
26 11 11 1 11 1 11 11 9 1 9 1 9 9 11 11 1 9 9 1 9 11 11 1 13 4 2
56 15 1 2 11 9 1 11 11 11 2 11 2 1 9 1 13 16 15 10 9 1 9 13 1 9 13 16 15 11 1 9 1 9 1 13 4 9 11 1 9 9 1 1 9 1 9 13 13 4 9 1 9 1 9 13 2
25 0 9 11 11 11 1 0 0 9 11 11 1 9 1 11 1 9 9 11 1 13 1 9 13 2
53 11 1 9 13 4 1 9 13 4 11 1 15 9 1 13 16 9 1 1 11 1 9 13 4 16 11 11 9 1 0 0 9 11 11 9 9 1 1 9 13 1 1 15 9 9 11 11 1 9 13 4 4 2
28 11 11 9 1 12 0 9 2 0 9 2 1 9 9 1 0 9 1 13 1 9 1 9 9 13 4 4 2
33 9 11 1 3 12 10 9 1 9 9 1 9 13 4 4 4 7 11 1 10 12 0 9 1 0 9 1 9 9 13 4 4 2
9 15 1 12 12 9 1 9 13 2
12 15 9 11 7 11 1 9 1 1 13 4 2
20 9 9 9 9 1 9 0 13 4 4 7 11 11 1 15 0 13 4 4 2
47 11 11 11 11 11 11 1 0 9 1 9 1 13 16 10 9 9 1 0 9 1 15 14 13 4 4 4 16 15 3 13 0 9 1 9 9 1 9 13 15 0 9 1 13 14 4 2
15 11 1 13 16 10 3 9 3 13 1 9 14 13 4 2
30 16 11 1 14 0 7 0 9 9 1 1 14 12 9 1 9 13 2 7 9 1 0 15 14 9 1 15 14 13 2
19 11 1 13 16 10 0 9 1 9 13 4 2 15 15 1 9 14 13 2
17 15 11 1 9 13 4 13 16 9 13 1 1 15 9 14 13 2
30 9 9 1 9 1 0 9 1 9 13 1 10 9 13 2 16 0 9 1 9 1 0 9 1 9 12 9 14 13 2
22 0 12 9 1 9 7 9 1 13 4 1 9 1 12 9 1 9 13 1 9 13 2
18 11 1 0 13 16 9 15 11 11 7 11 11 1 13 3 0 13 2
13 9 9 9 1 9 11 11 1 0 13 4 4 2
10 11 11 1 9 1 9 13 4 4 2
19 0 12 9 1 9 1 9 13 4 4 15 10 9 1 0 9 13 4 2
36 11 1 13 16 0 12 9 1 11 11 1 9 1 9 1 15 9 14 13 4 4 2 16 10 12 0 9 1 9 1 13 9 13 4 4 2
29 0 9 1 14 9 13 1 14 9 13 4 4 2 7 10 9 10 9 1 1 1 0 13 16 15 9 13 4 2
24 11 11 11 1 13 16 11 9 1 9 1 9 9 7 11 1 11 9 1 9 13 4 4 2
19 11 1 9 11 11 1 13 16 9 9 1 11 11 9 1 3 13 4 2
29 7 15 0 9 1 0 13 4 4 16 9 1 1 1 13 9 9 1 9 1 9 9 13 1 9 13 4 4 2
12 15 1 9 1 1 9 1 9 0 13 4 2
25 14 12 9 1 9 1 13 11 11 11 11 1 9 11 11 11 1 11 9 1 0 13 4 4 2
12 11 1 11 9 11 11 9 1 0 13 4 2
18 15 11 1 11 1 1 11 11 1 9 1 14 9 14 9 13 4 2
12 15 12 12 12 9 1 10 1 9 13 4 2
44 9 1 1 11 1 10 9 1 10 9 1 12 9 13 2 7 3 14 2 11 11 2 1 9 9 2 9 0 13 4 7 12 9 1 12 9 1 9 1 10 9 14 13 2
21 11 1 0 9 14 10 14 9 1 1 9 1 9 13 1 9 1 9 1 13 2
23 11 11 11 1 11 2 11 2 11 7 11 9 1 14 12 9 9 1 9 13 4 4 2
14 11 1 15 1 9 1 9 13 1 0 9 0 13 2
17 15 1 11 1 9 1 9 11 9 1 11 9 1 13 4 4 2
25 9 1 1 11 11 9 9 1 9 9 11 11 1 9 13 4 16 11 11 11 1 13 1 13 2
14 0 9 1 9 1 12 0 9 9 1 9 13 4 2
15 9 9 1 11 9 11 11 9 1 9 1 0 13 4 2
38 11 11 9 9 9 11 11 1 1 2 11 11 11 1 9 1 9 13 4 16 11 1 15 12 0 9 13 7 12 12 12 9 9 14 13 4 4 2
23 15 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 7 11 11 9 0 13 2
22 9 1 1 11 11 11 9 1 3 10 9 1 9 10 2 0 13 1 9 13 4 2
14 10 9 1 15 9 1 14 12 12 9 1 9 13 2
20 9 11 11 1 1 9 1 9 1 1 10 9 15 13 3 0 13 4 4 2
22 11 10 9 9 1 9 13 11 7 9 2 3 1 9 1 9 1 9 13 4 4 2
15 15 14 15 12 14 9 10 2 10 9 1 13 4 4 2
21 0 9 9 1 14 1 9 11 11 1 0 13 1 0 9 1 0 9 13 4 2
35 9 11 1 11 1 1 9 9 1 9 13 1 11 15 1 3 12 9 13 4 4 7 15 0 9 13 2 15 15 9 9 14 13 4 2
14 15 0 9 1 9 1 9 11 11 1 13 4 4 2
26 11 1 1 15 3 0 9 13 16 15 10 9 1 9 1 9 13 4 4 15 15 9 13 4 4 2
33 11 1 3 13 1 3 14 11 11 1 9 1 9 11 11 7 11 1 0 9 11 11 1 12 9 1 9 1 0 13 4 4 2
14 11 11 1 14 15 0 9 1 13 1 9 1 13 2
34 9 1 9 9 11 11 1 9 1 9 1 13 16 9 1 11 1 9 13 1 3 13 4 16 15 9 1 13 1 1 12 9 13 2
11 3 9 1 1 15 3 0 13 4 4 2
26 15 15 1 9 1 13 2 15 1 1 15 9 1 9 1 9 1 13 1 3 14 15 13 4 4 2
12 10 9 15 14 9 7 0 9 13 4 4 2
26 15 9 13 4 9 1 13 4 16 0 12 9 1 15 0 13 4 7 15 1 15 0 9 13 4 2
25 16 2 3 9 1 9 13 1 9 11 1 1 9 0 13 16 15 15 0 9 1 13 4 4 2
31 11 9 1 1 15 15 0 9 1 14 12 9 1 8 13 4 2 7 0 13 1 1 15 0 9 9 1 14 13 4 2
19 0 13 16 11 1 9 0 13 1 1 11 9 9 1 14 14 13 4 2
12 10 9 9 1 13 4 16 15 0 9 13 2
18 7 11 1 9 9 13 16 15 11 1 11 11 1 0 13 4 4 2
21 15 1 1 11 1 13 16 9 1 12 9 11 1 15 9 0 13 1 9 13 2
18 15 0 9 1 1 9 2 9 7 9 1 9 14 0 13 4 4 2
8 15 1 15 10 9 14 13 2
17 15 0 9 1 13 4 9 14 13 4 7 15 15 9 14 13 2
11 15 1 12 12 9 15 9 13 4 4 2
13 9 1 1 11 15 1 10 0 0 13 4 4 2
29 0 13 16 0 9 9 1 1 14 11 9 1 9 13 4 4 7 9 1 15 13 1 9 1 9 13 4 4 2
16 7 0 9 1 9 1 15 13 1 1 0 9 13 4 4 2
19 11 0 9 1 0 14 13 4 7 11 13 1 3 15 3 0 13 4 2
21 11 11 1 11 11 11 11 1 13 16 11 11 11 1 0 9 13 4 0 13 2
11 15 13 16 15 13 1 9 13 4 4 2
15 11 1 13 16 10 9 9 1 1 12 9 1 9 13 2
12 11 11 11 11 11 11 11 1 9 14 13 2
21 11 1 13 16 11 11 11 11 1 9 1 0 9 1 9 13 4 0 9 13 2
9 7 10 9 15 9 13 4 4 2
17 9 9 11 11 11 1 9 1 13 9 1 0 9 0 13 4 2
33 9 9 1 15 12 9 1 13 16 10 9 9 1 9 1 15 9 1 13 1 1 9 1 9 9 1 0 13 1 9 13 4 2
16 15 10 9 14 13 2 15 9 1 15 9 2 9 14 13 2
41 9 11 1 11 9 2 11 11 11 11 11 2 9 1 11 11 11 11 11 11 1 13 2 2 10 9 13 4 4 15 14 9 1 15 9 1 9 14 13 4 2
14 16 15 14 13 4 2 16 13 15 9 1 9 15 13
11 9 1 11 11 11 11 11 14 0 13 2
42 7 15 13 9 1 2 10 0 9 14 0 9 1 9 1 13 1 9 13 4 4 2 7 10 9 9 13 1 1 10 9 0 13 16 15 1 3 9 13 4 4 2
36 10 9 15 9 1 9 9 1 15 9 2 9 14 13 2 10 9 1 9 13 13 4 7 13 4 16 15 9 13 1 1 3 0 9 13 2
15 9 9 11 1 13 16 9 1 15 13 9 1 13 4 2
15 15 9 1 9 13 16 15 9 7 9 14 15 9 13 2
19 15 13 16 10 10 14 9 9 1 0 9 13 4 1 9 1 14 13 2
26 9 1 9 1 9 7 0 9 1 1 11 1 11 11 1 12 9 1 12 9 9 1 1 9 13 2
27 0 9 1 0 12 9 11 11 2 11 7 11 1 0 9 1 9 1 1 12 9 1 9 1 9 13 2
22 11 1 11 11 1 12 9 9 2 11 1 12 7 11 1 12 9 1 1 9 13 2
12 15 1 12 9 9 1 9 11 1 13 4 2
9 10 9 1 9 1 0 9 13 2
42 0 9 1 9 1 10 0 9 1 9 1 9 13 4 2 15 9 1 11 11 11 11 2 11 2 2 11 11 11 11 11 2 11 2 7 9 11 11 0 0 13 2
12 11 11 1 9 1 11 1 9 13 4 4 2
17 3 0 9 1 9 9 1 13 4 9 1 0 9 13 4 4 2
37 0 9 1 1 14 11 11 1 14 11 7 11 1 12 9 13 4 4 2 7 11 7 11 1 3 12 7 12 9 1 0 9 0 13 4 4 2
21 10 9 1 11 11 1 10 12 9 0 13 4 2 15 1 11 1 12 9 13 2
8 11 11 1 12 9 13 4 2
9 12 9 1 11 9 13 4 4 2
23 11 1 12 9 13 4 7 12 9 11 11 11 1 1 7 12 9 11 1 1 13 4 2
13 9 1 0 7 9 9 0 9 1 13 0 13 2
21 15 13 13 16 9 9 1 0 9 1 1 9 1 9 9 1 0 9 14 13 2
21 11 11 1 9 1 1 2 0 9 1 9 9 1 9 1 9 9 1 13 4 2
8 10 12 9 9 13 4 4 2
11 10 9 1 12 9 9 1 9 13 4 2
42 9 1 9 1 13 4 9 1 9 13 4 16 9 2 9 9 1 9 1 13 0 9 1 1 0 9 1 9 13 4 16 0 9 1 9 9 1 0 13 4 4 2
27 11 11 1 0 9 9 1 9 1 1 9 1 0 9 1 9 9 9 9 11 11 11 1 10 9 13 2
42 11 11 11 1 13 16 10 9 1 9 9 13 4 4 7 10 0 0 9 1 9 2 9 9 9 1 9 2 9 7 9 9 14 9 13 1 9 13 4 4 4 2
50 9 1 9 1 9 1 9 9 13 4 11 11 11 1 13 16 16 11 11 1 9 1 1 9 9 1 9 1 9 12 9 13 14 4 4 16 9 1 9 0 13 1 12 1 12 9 1 9 13 2
15 15 13 16 15 1 9 1 0 9 1 14 9 13 4 2
15 15 13 16 9 1 0 9 13 15 3 14 13 4 4 2
18 15 13 16 0 9 1 9 1 9 13 1 0 9 10 0 13 4 2
26 0 9 1 9 1 9 1 10 9 13 4 7 15 8 0 9 1 1 9 1 9 1 13 4 4 2
29 15 13 16 3 10 14 10 0 9 1 9 11 7 9 2 9 9 9 1 13 15 9 1 0 9 13 4 4 2
12 15 1 0 9 1 9 1 15 9 14 13 2
20 15 13 16 9 1 0 9 1 9 13 1 9 0 9 9 1 1 13 4 2
42 9 1 9 1 1 9 1 9 1 13 1 1 1 15 13 16 15 9 1 9 1 9 1 1 7 9 1 1 9 7 9 1 9 1 1 0 2 0 9 13 4 2
46 15 13 16 10 9 1 9 1 1 9 1 9 9 0 13 4 16 9 1 9 13 4 1 9 7 10 9 1 0 9 1 0 10 0 9 1 3 9 9 1 0 13 4 4 4 2
27 10 9 1 9 13 4 4 16 15 9 9 1 1 10 9 0 13 16 9 1 15 3 9 0 13 4 2
32 15 13 16 10 9 9 1 1 10 9 14 0 13 4 16 10 9 1 9 9 1 13 1 9 1 9 15 1 0 9 13 2
14 10 0 9 1 14 10 9 0 13 1 9 13 4 2
32 11 11 11 11 1 1 1 0 9 1 1 11 11 11 11 14 1 0 9 1 9 9 1 13 4 1 9 13 4 4 4 2
21 9 1 9 13 1 1 1 11 11 2 11 1 1 9 13 1 9 14 13 4 2
10 9 9 1 9 1 15 9 13 4 2
43 9 9 1 9 11 11 11 1 13 16 11 11 11 11 1 0 9 1 1 11 11 11 11 14 1 0 9 1 15 15 14 9 1 15 9 9 1 14 13 4 4 4 2
26 9 0 13 9 1 0 13 4 4 16 15 9 13 1 1 1 11 11 11 1 1 1 9 13 4 2
34 9 1 15 14 13 4 4 16 11 11 11 11 1 0 9 1 9 13 1 1 1 11 11 2 11 1 1 0 9 9 1 13 4 2
56 15 1 11 11 11 1 9 9 1 9 1 1 14 10 0 9 2 9 9 1 9 2 9 9 1 9 2 9 9 2 9 9 2 0 9 7 0 9 1 11 11 11 11 1 0 9 1 9 1 13 1 9 13 4 4 2
11 11 1 9 1 9 13 15 0 9 14 2
26 11 11 1 11 1 10 0 9 1 3 13 4 11 2 11 11 1 1 12 9 9 1 9 0 13 2
15 9 1 1 11 11 1 0 9 11 1 14 9 13 4 2
18 7 11 11 1 9 7 11 1 0 9 11 1 9 3 10 13 4 2
14 15 12 12 9 1 9 1 1 9 0 13 4 4 2
16 11 1 9 11 1 9 1 1 1 12 12 9 10 13 4 2
12 11 11 11 11 11 1 9 1 9 0 13 2
11 9 1 9 7 9 9 1 9 13 4 2
11 11 11 1 13 4 9 0 9 1 13 2
17 16 11 1 9 1 9 1 1 1 15 9 13 1 9 13 4 2
23 9 11 2 11 1 1 11 11 1 1 0 9 1 9 1 9 1 0 9 1 9 13 2
22 15 10 9 14 0 13 2 15 11 11 1 1 9 1 9 9 1 0 13 4 4 2
16 15 0 13 1 1 12 12 9 1 0 9 1 9 13 4 2
17 11 11 11 11 2 11 2 1 12 9 1 10 9 13 4 4 2
12 9 1 1 9 1 9 0 9 1 9 13 2
27 9 9 1 9 1 9 1 9 1 11 11 11 1 13 4 4 16 9 9 1 10 9 1 3 9 13 2
26 9 1 9 1 9 1 15 11 11 11 2 11 2 1 9 1 10 9 1 9 1 9 1 9 13 2
39 9 1 15 9 1 12 9 9 1 0 9 1 9 1 0 13 2 12 9 1 9 1 9 7 12 9 1 9 1 12 9 1 0 13 1 9 14 13 2
16 9 1 11 1 0 10 9 1 10 9 1 0 13 4 4 2
23 15 13 4 4 16 9 1 1 10 9 1 1 10 9 9 9 9 1 1 0 9 13 2
14 15 10 9 1 9 13 1 1 0 9 13 4 4 2
40 9 1 9 1 9 1 15 13 4 14 0 13 4 4 16 11 11 1 11 11 1 1 15 12 12 9 9 1 9 1 9 0 9 1 9 0 13 1 13 2
26 9 1 1 2 9 1 0 0 13 1 15 9 1 9 1 9 9 15 0 9 0 14 13 4 4 2
24 9 1 9 13 4 4 16 11 11 9 13 16 15 9 1 10 9 1 9 1 9 13 4 2
21 11 1 11 11 11 1 11 9 1 9 1 11 1 9 13 1 9 3 13 4 2
19 11 1 13 13 16 10 9 1 9 13 14 10 9 1 9 0 14 13 2
18 3 11 1 11 1 9 2 9 9 9 13 1 15 9 14 13 4 2
36 0 11 11 11 11 1 1 9 1 0 11 11 11 1 13 16 0 11 9 1 9 13 14 11 11 9 1 0 9 1 9 14 13 4 4 2
22 0 11 11 11 1 11 11 1 9 9 1 1 11 1 13 4 4 9 1 9 13 2
15 15 1 12 9 1 0 9 1 0 9 1 9 9 13 2
25 11 1 1 1 0 12 0 9 1 13 4 4 16 11 11 1 1 0 9 1 0 13 13 4 2
39 3 11 1 9 13 16 0 11 11 11 11 1 11 9 1 1 9 2 9 9 1 9 1 9 1 0 9 13 2 7 11 1 11 1 3 0 13 4 2
25 11 1 12 9 1 1 9 9 1 9 1 9 13 1 1 9 2 9 9 9 13 1 9 13 2
25 11 11 7 11 11 1 9 1 9 1 9 2 9 9 9 1 9 1 9 0 9 1 0 13 2
13 11 1 11 1 9 2 9 1 9 1 9 13 2
20 15 11 1 13 16 11 1 9 9 1 13 4 15 9 2 9 0 13 4 2
23 15 0 9 2 9 1 9 9 13 13 1 1 11 1 9 2 9 13 4 1 9 13 2
21 15 11 1 10 9 14 13 16 15 11 1 12 0 0 0 0 9 1 9 13 2
25 9 9 9 1 1 11 1 13 16 15 9 13 4 4 16 11 1 0 9 1 0 13 4 4 2
14 11 1 11 11 1 13 11 1 9 1 3 9 13 2
25 15 13 16 11 1 11 11 1 9 7 9 1 9 13 1 1 15 9 13 4 2 15 0 13 2
41 9 2 9 1 9 1 15 15 9 14 14 13 2 7 0 3 13 16 11 9 2 9 1 9 1 11 1 9 1 13 4 7 10 9 1 9 3 13 4 4 2
16 15 13 16 11 1 0 2 0 9 1 11 0 9 13 4 2
10 15 9 9 1 14 9 13 13 4 2
15 15 0 2 0 9 1 11 1 9 1 14 3 9 13 2
19 15 13 16 11 1 9 1 1 11 1 10 9 13 4 2 15 0 13 2
12 11 1 15 0 9 1 1 0 9 9 13 2
21 11 11 11 1 9 1 1 11 11 11 9 1 13 4 15 9 1 13 4 4 2
36 0 9 1 9 13 4 9 1 0 9 11 11 1 9 1 13 16 15 12 9 1 9 1 1 11 11 1 9 13 1 1 9 9 14 13 2
23 11 11 1 9 1 10 9 1 3 9 13 4 9 1 0 13 1 11 0 0 9 13 2
14 15 1 12 9 1 9 1 10 9 1 9 13 4 2
15 11 1 9 1 13 15 9 1 10 9 1 9 13 4 2
26 9 1 9 11 11 1 9 1 13 16 15 15 1 3 1 9 1 9 13 7 15 0 13 4 4 2
15 3 1 15 9 1 9 13 16 9 1 13 4 4 4 2
28 9 9 1 9 11 11 1 13 1 15 13 16 15 10 9 1 14 13 2 15 9 15 9 9 1 0 13 2
26 0 11 11 11 1 15 0 11 9 3 11 1 11 11 11 1 15 0 9 1 13 4 0 13 4 2
25 11 9 1 11 11 1 11 1 0 9 1 1 11 12 9 1 1 9 13 4 1 13 13 4 2
36 11 1 15 11 9 0 13 4 1 12 0 9 1 0 9 1 1 11 1 12 9 1 9 1 0 9 1 13 4 10 9 0 13 4 4 2
15 11 1 11 9 11 11 1 9 1 12 9 1 13 4 2
21 0 9 1 15 9 13 4 16 12 9 1 9 1 1 9 15 9 1 9 13 2
36 11 1 11 9 0 13 1 15 1 9 10 9 1 13 4 4 16 11 2 11 1 1 13 9 1 13 11 1 11 1 15 0 9 13 4 2
37 0 9 2 11 2 1 9 1 1 11 1 11 1 0 11 9 1 9 13 4 1 1 15 11 1 11 1 10 9 13 4 11 1 13 4 4 2
13 15 1 9 1 11 1 11 9 1 9 10 13 2
17 11 9 11 11 11 11 11 1 9 1 0 13 11 1 11 13 2
35 9 9 9 11 1 11 1 9 9 1 13 11 11 1 9 1 9 1 13 4 7 11 1 10 9 1 11 11 1 9 1 9 13 4 2
25 3 0 0 9 1 9 11 1 9 1 0 13 1 0 9 9 1 9 1 9 13 4 4 4 2
24 15 1 14 0 11 11 11 11 11 11 14 11 11 1 13 4 10 9 1 9 13 4 4 2
15 15 13 13 16 15 10 9 1 9 9 1 13 4 4 2
14 9 10 9 1 9 15 0 9 1 1 13 4 4 2
28 11 1 9 11 11 1 13 16 11 1 11 11 7 11 11 1 1 1 11 11 1 9 1 9 1 13 4 2
11 11 9 1 1 9 1 9 13 4 4 2
9 15 11 11 1 9 1 0 13 2
11 11 11 1 9 1 15 9 13 13 4 2
18 0 13 16 10 0 9 9 1 11 11 1 13 4 9 9 0 13 2
13 10 9 9 9 9 1 9 14 0 13 4 4 2
15 15 13 16 10 9 1 9 1 10 9 1 9 0 13 2
13 15 15 9 1 13 9 13 4 1 9 13 4 2
31 15 13 16 0 10 9 1 10 9 1 9 9 1 9 13 1 9 1 13 9 7 9 1 0 9 1 13 4 4 4 2
15 15 13 16 9 1 0 9 1 9 9 15 1 0 13 2
18 10 9 1 0 13 1 3 0 0 9 1 13 1 9 13 4 4 2
16 10 9 9 7 9 1 9 1 13 1 14 0 9 13 4 2
25 11 1 12 9 1 11 1 13 16 9 1 11 1 0 13 4 10 9 12 2 12 9 0 13 2
27 0 13 16 11 1 1 11 11 2 11 11 11 11 7 11 11 11 14 1 9 1 14 10 9 0 13 2
26 9 1 0 9 1 0 11 11 1 11 11 1 9 13 4 11 11 1 1 9 1 0 9 13 4 2
35 12 9 1 10 9 1 11 9 11 11 2 11 11 11 2 15 9 9 2 11 0 9 1 11 7 0 9 1 0 9 0 13 4 4 2
29 11 9 1 9 1 11 0 0 9 1 1 9 1 0 12 9 1 13 9 1 13 4 9 1 0 9 13 4 2
49 15 1 14 9 9 1 1 1 0 9 7 0 9 1 9 1 13 11 11 11 11 2 11 2 7 11 11 1 1 1 13 4 1 9 1 9 1 1 1 0 9 1 14 9 1 13 4 4 2
31 9 9 9 11 11 11 1 13 16 9 9 1 0 9 1 13 4 0 9 1 12 1 10 9 1 0 13 4 4 4 2
17 15 1 11 0 9 1 0 9 1 12 9 0 13 4 4 4 2
31 9 1 11 11 11 11 11 1 13 16 9 1 9 1 9 13 4 1 9 1 13 4 9 1 0 9 13 4 4 4 2
20 15 1 9 9 2 9 2 9 9 2 9 7 0 9 1 9 9 13 4 2
12 11 9 1 11 9 11 11 1 0 13 4 2
11 15 11 9 11 11 1 9 13 4 4 2
17 11 11 11 11 11 1 13 16 11 11 1 9 1 9 1 13 2
7 15 9 13 4 4 4 2
15 11 1 11 1 11 11 11 11 11 1 9 0 13 4 2
18 15 11 1 0 9 11 11 11 1 11 2 11 2 11 1 13 4 2
25 16 2 11 1 11 11 11 11 1 9 13 1 9 1 1 11 11 9 1 9 1 0 13 4 2
15 15 13 4 1 16 11 9 1 11 1 9 13 4 4 2
14 15 1 15 13 16 15 1 9 13 15 0 14 13 2
10 15 1 1 15 14 13 14 4 4 2
27 9 9 1 9 1 1 11 11 11 11 1 11 1 0 13 16 9 9 1 9 1 9 0 14 13 4 2
28 9 1 11 11 11 11 11 1 1 1 0 9 1 9 1 15 9 1 13 16 15 9 9 0 14 13 4 2
15 10 15 14 9 13 4 4 2 15 0 13 4 4 4 2
18 9 1 9 1 9 1 9 1 1 1 15 13 16 9 0 13 4 2
21 9 9 1 9 1 1 1 11 1 13 16 15 10 10 9 1 15 9 14 13 2
14 15 13 16 3 14 0 9 1 9 1 9 13 4 2
20 15 1 9 9 1 9 1 11 1 13 4 9 1 9 0 13 1 9 13 2
18 9 1 11 9 11 11 1 9 1 9 1 9 0 13 1 9 13 2
37 11 1 9 9 1 0 12 9 13 4 4 2 7 11 9 11 11 9 9 1 9 13 1 1 9 9 1 9 3 13 1 9 1 13 4 4 2
23 9 9 1 9 15 1 14 13 2 15 1 15 15 9 9 1 9 1 9 13 4 4 2
7 10 9 0 9 1 13 2
17 11 1 0 9 13 1 9 1 13 9 1 0 9 0 13 4 2
16 11 11 1 9 13 1 1 9 1 0 9 1 9 13 4 2
27 11 11 15 0 13 13 4 16 15 9 9 1 1 10 15 9 14 13 15 1 15 9 1 9 13 4 2
16 0 11 1 11 9 9 1 9 11 0 9 9 13 4 4 2
31 15 13 16 0 10 9 1 9 9 0 13 1 1 15 15 9 1 9 1 15 9 1 13 4 9 1 13 1 0 13 2
11 9 1 10 9 1 13 1 9 13 4 2
16 11 7 15 9 9 1 13 9 1 13 1 9 13 4 4 2
12 15 9 1 0 9 1 12 9 7 9 13 2
16 15 9 1 15 9 1 13 9 14 1 13 1 13 4 4 2
22 11 1 13 16 9 1 10 3 1 15 9 1 9 7 11 1 9 9 13 4 4 2
21 15 13 16 16 15 1 9 1 13 15 9 9 1 13 4 16 9 15 9 13 2
19 9 14 1 9 1 11 11 11 1 1 1 9 1 9 1 9 13 4 2
17 11 14 9 9 1 9 1 9 13 1 15 9 14 13 4 4 2
33 0 9 9 1 1 11 11 1 3 13 1 0 9 9 11 11 1 11 1 13 16 15 11 11 11 2 11 2 1 13 4 4 2
31 11 1 13 16 11 9 11 11 1 11 13 1 9 13 1 3 10 9 0 13 4 4 2 15 1 1 15 9 13 4 2
35 11 1 15 11 9 1 9 1 13 16 15 0 9 1 11 11 1 11 13 1 9 1 11 13 4 2 7 15 11 13 1 9 13 4 2
10 7 2 15 15 9 1 9 14 13 2
9 9 1 11 1 15 0 9 13 2
28 11 11 1 9 1 1 1 0 9 9 13 1 11 1 13 16 11 1 15 9 1 15 14 10 0 9 13 2
19 15 13 16 15 0 9 1 9 1 13 15 1 15 11 1 0 13 4 2
18 0 12 9 1 9 1 13 11 11 11 11 12 9 3 9 1 13 2
15 11 1 11 1 9 9 9 1 0 9 9 13 4 4 2
21 11 1 1 0 11 11 11 11 1 9 1 1 9 1 9 1 9 13 4 4 2
13 11 1 11 1 0 9 1 12 9 0 13 4 2
34 15 1 9 1 1 11 1 9 9 1 12 9 1 11 11 1 12 9 1 9 1 9 1 9 1 11 11 11 1 0 9 13 4 2
10 10 9 1 10 9 12 12 9 13 2
33 3 1 9 9 1 13 4 16 9 1 11 1 9 1 10 9 0 13 4 10 9 1 3 10 9 1 15 9 1 9 13 4 2
13 15 1 1 9 1 12 12 9 0 9 13 4 2
19 11 1 1 11 11 1 10 9 1 9 0 13 1 15 9 14 13 4 2
38 9 9 1 9 13 4 16 9 1 9 1 9 13 1 3 14 9 14 13 7 9 1 9 1 9 13 4 15 9 1 12 12 9 1 0 9 13 2
43 11 11 1 11 11 11 11 2 11 11 2 9 2 9 9 2 9 2 9 9 2 9 9 2 9 9 9 9 2 9 2 9 9 7 9 9 1 9 1 9 13 4 2
25 11 11 11 1 11 9 11 1 13 4 16 9 9 1 0 9 1 9 1 9 1 9 13 4 2
32 15 13 16 9 1 9 2 9 2 9 2 9 2 9 7 9 1 14 13 1 9 1 10 9 1 9 1 13 4 4 4 2
37 11 11 11 11 2 11 2 1 0 11 11 11 11 11 1 0 9 1 1 1 11 1 13 16 11 1 9 11 1 9 1 13 14 4 4 4 2
21 9 11 1 9 1 11 1 9 13 4 7 15 11 11 11 11 1 9 9 13 2
13 15 13 16 9 1 9 1 9 1 12 9 13 2
28 15 9 9 9 13 2 9 1 9 14 13 2 9 1 9 2 9 2 9 7 0 9 9 1 14 13 4 2
15 7 10 9 1 3 13 1 1 0 9 13 1 9 13 2
14 11 1 13 16 0 10 9 1 9 1 9 13 4 2
36 9 1 9 1 0 9 1 9 1 13 1 3 14 9 2 0 9 1 9 2 9 1 9 7 9 1 9 1 12 2 12 13 4 4 4 2
31 15 13 16 11 11 1 9 1 9 1 9 13 1 1 10 9 1 9 13 4 7 13 1 1 1 15 9 9 1 13 2
14 11 11 9 1 1 13 11 11 1 9 13 4 4 2
16 15 9 15 9 1 0 9 1 1 0 9 1 14 13 4 2
32 11 11 11 2 11 2 0 0 9 1 9 1 9 1 11 1 15 11 11 11 2 11 2 11 1 9 13 1 9 1 13 2
31 11 1 11 11 11 11 1 11 1 15 9 1 13 16 15 11 1 11 11 1 9 13 4 2 15 10 0 9 13 4 2
22 15 13 16 15 15 3 0 9 13 16 15 10 0 13 7 3 9 9 13 1 13 2
28 11 1 13 16 0 9 1 11 1 9 9 13 1 1 1 15 11 11 1 9 1 9 13 1 1 0 13 2
38 11 11 1 0 9 1 9 1 1 11 7 11 11 11 2 11 2 1 3 9 13 7 0 11 1 11 1 15 12 9 1 9 9 0 13 4 4 2
20 15 13 16 11 1 10 9 1 1 11 1 9 9 7 9 1 1 9 13 2
27 9 11 1 13 1 9 9 1 0 9 1 9 1 9 1 13 4 1 9 11 11 1 0 9 1 13 2
27 11 11 11 11 1 11 11 1 0 9 9 1 1 1 9 1 9 13 1 3 9 13 15 1 13 4 2
22 10 9 10 9 1 13 4 2 15 11 1 0 9 9 13 1 0 3 9 13 4 2
19 15 1 15 9 9 13 1 3 14 9 7 9 1 9 13 4 4 4 2
34 3 10 0 9 1 1 9 1 9 9 11 1 9 13 4 2 16 16 9 9 1 11 11 11 1 2 11 11 2 1 9 1 13 2
34 15 1 1 13 4 1 11 1 13 16 3 10 9 11 1 13 4 4 7 11 1 11 1 1 0 9 13 1 1 15 13 4 4 2
11 15 13 16 9 11 1 9 13 13 4 2
23 9 1 0 9 1 1 14 15 0 13 16 15 9 13 16 9 9 1 15 9 15 13 2
9 15 15 0 9 1 0 9 13 2
26 3 9 1 10 9 1 12 9 14 0 13 16 0 12 9 1 15 9 1 15 9 1 9 14 13 2
14 10 9 1 9 11 11 1 9 1 14 9 13 4 2
29 9 1 10 9 1 1 9 1 15 14 13 1 9 13 4 16 15 9 1 13 4 14 11 1 9 13 4 4 2
35 9 1 11 11 1 0 9 13 3 10 9 13 1 0 9 13 7 11 11 1 12 9 9 0 13 1 1 9 1 9 7 9 13 4 2
21 9 1 14 1 9 1 9 11 11 1 11 1 0 9 1 9 1 9 13 4 2
17 15 13 16 11 1 9 1 9 1 9 13 2 15 10 9 13 2
12 11 1 9 1 9 1 10 9 10 0 13 2
24 15 1 9 1 0 9 11 1 11 1 9 9 1 11 11 1 13 4 11 1 9 13 4 2
17 7 11 1 11 1 9 1 1 14 11 1 9 1 13 4 4 2
17 15 1 11 1 1 0 9 1 11 1 0 9 1 9 13 4 2
28 15 9 1 11 1 11 1 9 9 1 12 2 12 1 13 1 1 9 9 1 9 12 2 12 1 13 4 2
27 11 1 9 1 1 11 1 15 9 1 11 11 1 1 12 9 9 1 9 12 2 12 1 0 13 4 2
14 0 9 1 14 9 15 9 1 9 9 13 4 13 2
22 0 9 1 12 9 9 9 11 11 1 0 0 9 1 9 9 1 9 13 13 4 2
25 10 9 1 1 11 7 11 1 0 0 9 1 9 1 9 3 13 1 1 3 9 1 9 13 2
19 15 9 13 1 1 9 2 0 9 7 0 0 9 3 0 13 4 4 2
51 11 11 11 11 11 11 2 11 2 9 9 9 1 11 11 1 12 0 9 1 13 4 13 16 15 15 13 16 0 9 7 0 9 1 13 1 9 1 1 0 9 9 13 1 9 1 9 13 4 4 2
14 9 1 10 9 0 9 1 9 1 1 9 13 4 2
26 2 11 11 11 2 7 0 9 1 9 1 15 1 1 0 9 9 0 0 11 11 1 0 13 4 2
11 15 1 0 9 1 9 7 0 9 13 2
27 0 9 1 11 9 1 1 11 11 1 13 0 0 9 1 0 9 1 12 12 9 1 9 0 13 4 2
14 15 10 9 12 9 11 1 0 9 9 1 13 4 2
12 0 12 12 9 3 9 9 1 13 4 4 2
18 7 11 11 11 1 0 9 9 1 1 12 12 9 9 13 4 4 2
15 11 1 9 9 1 0 9 13 1 9 14 13 4 4 2
23 0 11 9 11 11 11 1 12 9 3 9 1 0 9 1 1 9 1 9 13 4 4 2
25 15 13 4 16 9 9 11 11 1 1 9 1 13 4 9 1 1 11 9 1 1 13 4 4 2
20 15 13 16 11 1 0 11 11 11 1 15 9 1 9 13 1 1 13 4 2
22 11 1 13 16 11 2 11 7 11 1 0 11 9 9 9 1 15 9 1 0 13 2
17 15 13 16 9 0 13 4 4 16 9 9 1 1 3 9 13 2
24 15 1 9 13 14 11 1 13 16 15 11 1 1 13 1 9 1 1 9 14 13 4 4 2
15 10 9 0 9 1 13 9 9 1 9 1 0 13 4 2
33 15 13 4 1 16 15 15 9 1 13 2 15 13 16 15 15 0 9 1 1 1 9 13 1 1 11 9 1 13 4 4 4 2
16 11 1 13 16 11 7 11 1 9 1 9 0 13 4 4 2
19 11 11 2 11 11 2 11 11 7 11 11 1 9 1 9 13 4 4 2
22 11 11 1 11 2 11 2 11 2 11 11 7 12 0 9 1 9 11 1 13 4 2
10 10 9 1 9 9 9 13 4 4 2
20 11 1 13 16 11 11 1 11 11 1 9 1 9 13 1 9 13 4 4 2
18 11 1 13 16 11 1 1 13 1 9 9 1 9 1 13 4 4 2
16 15 13 16 15 15 0 9 9 1 0 13 1 9 13 4 2
9 9 1 9 13 15 10 0 13 2
26 0 9 1 9 1 11 11 1 9 9 1 9 13 4 0 9 1 9 13 1 1 11 13 4 4 2
17 0 13 16 11 1 14 12 9 1 11 1 9 1 9 13 4 2
23 15 13 4 16 9 15 9 1 13 4 4 7 15 9 9 9 1 1 13 4 4 4 2
19 11 11 11 1 0 12 2 0 9 9 1 13 9 1 9 10 0 13 2
20 15 9 13 16 11 11 11 1 9 2 9 1 0 9 1 1 0 9 13 2
9 11 11 1 9 1 9 1 13 2
9 11 11 1 11 1 9 11 13 2
11 15 1 15 11 1 11 1 11 9 13 2
18 11 1 11 11 1 0 11 2 11 11 11 1 0 9 13 0 13 2
14 10 0 9 9 1 0 13 1 0 9 13 4 4 2
31 11 1 13 1 0 0 9 11 11 11 1 9 11 11 1 11 1 9 13 4 13 16 11 1 9 1 13 9 0 13 2
15 9 1 9 13 16 11 9 1 9 9 1 0 9 13 2
26 15 10 14 9 13 16 11 11 2 11 1 1 9 1 14 9 1 9 1 9 1 9 13 4 4 2
30 15 13 16 16 11 0 0 11 11 11 11 1 9 7 15 9 1 9 13 4 16 15 11 1 9 1 0 9 13 2
18 15 11 9 1 1 11 0 11 11 1 9 9 1 0 13 4 4 2
9 3 10 9 11 11 1 9 13 2
12 15 11 1 9 15 0 7 0 9 13 4 2
14 10 9 11 1 11 1 0 9 1 9 13 4 4 2
18 0 9 9 1 10 9 1 11 11 1 0 13 1 9 13 4 4 2
17 12 9 1 13 16 11 1 10 0 9 1 9 13 4 4 4 2
22 15 13 16 16 11 9 1 9 1 1 0 9 1 9 13 4 16 15 9 0 13 2
34 11 1 0 0 9 11 11 1 9 11 11 1 13 16 11 1 10 9 14 13 4 4 4 16 15 9 1 9 9 1 0 9 13 2
7 9 0 9 13 4 4 2
24 10 9 1 10 9 13 16 15 9 1 1 9 7 0 9 1 9 1 9 13 1 14 13 2
15 14 10 9 1 9 13 1 9 15 1 9 13 4 4 2
5 10 9 14 13 2
43 15 1 13 16 15 0 9 1 9 9 1 13 9 1 1 13 2 15 9 1 1 13 4 2 16 9 1 9 13 16 9 1 9 9 1 13 9 1 9 10 13 4 2
13 13 14 15 14 3 15 12 9 0 13 4 4 2
32 9 9 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 7 11 11 1 11 1 9 0 13 4 2
15 7 11 11 2 11 11 7 11 11 3 13 4 4 4 2
20 9 1 11 11 15 9 7 11 11 11 1 0 9 1 9 1 1 0 13 2
20 10 9 1 11 11 11 1 13 16 10 10 9 1 9 1 1 0 9 13 2
8 15 9 1 9 1 9 13 2
12 9 1 1 11 11 1 9 1 9 13 4 2
19 15 11 1 13 16 9 1 13 4 15 9 1 9 13 1 9 13 4 2
11 7 10 9 1 1 15 0 14 13 4 2
13 15 2 11 15 10 9 1 0 13 1 9 13 2
12 11 11 1 14 9 1 13 1 0 9 13 2
9 7 15 9 1 9 13 4 4 2
14 11 11 1 9 1 15 11 11 1 9 1 13 4 2
19 15 13 13 16 9 9 1 9 9 1 13 9 1 1 3 15 1 13 2
21 11 11 1 15 9 1 9 13 4 11 1 9 1 12 9 9 13 1 9 13 2
22 15 13 13 16 12 9 9 1 0 13 0 9 1 9 10 9 1 9 13 4 4 2
35 9 11 11 1 13 16 9 1 9 9 1 13 10 9 1 0 14 13 16 15 15 15 9 13 4 4 2 15 15 0 13 15 9 13 2
10 11 7 11 11 1 14 15 9 13 2
25 11 11 1 11 11 1 11 9 11 11 11 1 9 1 13 11 9 1 11 1 0 13 4 4 2
19 11 1 9 13 16 9 9 1 15 11 1 9 1 1 9 0 14 13 2
34 9 1 13 16 11 9 11 1 0 9 1 14 1 11 1 9 13 1 9 13 16 9 0 9 1 11 9 1 10 9 9 13 4 2
34 13 4 4 16 11 9 11 11 1 14 11 11 11 11 11 1 9 13 15 11 7 0 11 9 1 9 1 13 15 9 1 0 13 2
14 11 0 9 3 11 11 1 0 2 9 1 0 13 2
20 15 1 11 1 15 2 11 11 2 9 0 13 1 9 9 9 1 13 4 2
25 9 1 13 16 9 1 1 12 0 9 9 1 1 12 0 9 9 10 9 11 1 1 13 4 2
12 15 12 9 9 7 12 9 9 14 13 4 2
14 11 1 10 15 9 9 13 1 9 1 9 13 4 2
21 15 9 13 16 15 9 9 7 11 1 13 1 9 1 9 0 9 1 13 4 2
15 16 15 1 11 1 10 9 1 9 9 1 0 13 4 2
32 11 11 1 1 10 9 1 12 0 9 1 9 13 1 0 9 1 13 4 9 1 1 1 9 1 1 9 2 9 0 13 2
9 10 9 11 1 9 1 13 4 2
47 11 11 11 11 11 1 9 1 1 13 16 0 9 1 1 0 9 1 0 9 1 11 11 1 1 10 9 0 13 1 3 11 11 1 9 13 4 7 15 15 1 1 10 9 13 4 2
17 15 13 16 0 9 1 15 1 1 9 11 11 1 1 13 4 2
31 0 9 1 10 9 1 9 1 10 14 10 12 9 1 9 13 1 0 11 11 11 11 11 11 1 9 1 0 13 4 2
12 10 9 1 9 9 1 1 13 15 9 13 2
16 11 11 11 11 11 11 1 10 9 1 9 1 3 0 13 2
18 0 9 0 13 0 9 1 10 9 9 1 10 9 1 0 13 4 2
29 11 9 11 11 1 13 16 11 9 1 10 9 1 0 13 9 1 15 9 9 1 12 0 9 1 0 13 4 2
43 9 1 10 9 13 4 4 2 15 12 9 1 1 15 0 9 1 0 13 2 0 9 12 9 0 13 7 9 1 15 1 0 9 1 9 0 13 14 1 9 0 13 2
17 11 1 9 0 13 1 3 15 9 1 9 13 4 1 9 13 2
16 9 1 9 9 9 1 10 9 13 1 14 9 13 4 4 2
27 9 0 13 4 11 11 11 1 13 16 0 9 1 9 1 12 12 9 1 10 9 1 0 13 4 4 2
18 15 13 16 12 9 1 1 9 1 10 12 9 1 9 0 13 4 2
25 9 1 10 9 14 13 4 4 16 16 15 9 1 9 14 13 4 4 16 15 9 9 13 4 2
21 11 9 11 11 1 11 11 11 1 9 1 1 9 7 11 9 1 3 9 13 2
15 0 9 1 13 1 9 1 1 15 9 1 14 9 13 2
17 11 1 15 0 9 13 4 13 16 15 0 9 1 0 9 13 2
12 11 11 1 9 1 0 9 1 1 13 4 2
14 15 13 16 9 1 9 1 10 9 12 0 9 13 2
23 15 9 1 0 14 9 13 2 2 9 15 11 1 9 1 3 0 9 1 0 13 4 4
12 9 1 1 15 10 9 11 9 1 9 13 2
36 15 13 16 10 9 1 0 9 9 11 1 0 9 1 9 1 13 7 3 0 9 11 1 11 1 11 11 1 9 1 14 15 1 9 13 2
16 9 11 11 7 9 11 11 1 9 14 15 9 1 9 13 2
17 15 13 16 11 1 11 14 0 9 1 1 11 11 11 11 13 2
10 3 11 1 11 11 11 11 11 13 2
9 15 10 9 1 13 1 9 13 2
25 11 11 1 9 1 9 1 10 9 13 4 2 7 9 1 9 1 9 10 0 14 13 4 4 2
17 11 1 9 1 9 1 13 4 9 1 10 9 9 1 0 13 2
10 3 2 3 9 13 9 13 4 4 2
18 9 1 1 1 10 14 9 13 14 15 9 1 15 13 4 4 4 2
17 3 15 13 13 4 7 15 1 9 2 9 1 9 9 13 4 2
19 12 9 1 1 9 1 9 9 1 1 1 9 1 12 2 12 9 13 2
6 16 15 11 14 13 2
12 9 1 1 14 15 10 9 1 10 13 4 2
16 11 1 11 11 9 1 13 4 9 11 1 9 1 13 4 2
51 11 9 1 9 1 9 9 1 0 11 11 2 11 2 1 9 7 0 11 11 11 11 1 9 11 11 11 1 9 1 1 9 13 4 9 1 12 1 10 9 1 1 9 1 0 13 1 9 13 4 2
14 0 0 9 11 1 11 1 9 13 1 9 13 4 2
28 9 1 11 1 9 1 12 9 1 9 1 11 11 11 11 1 1 9 1 0 9 1 9 1 9 0 13 2
11 9 9 11 1 11 11 11 1 9 13 2
28 11 1 11 1 11 9 1 9 14 13 1 9 13 4 9 1 9 0 13 1 1 11 11 1 1 9 13 2
11 16 11 1 15 1 1 15 9 14 13 2
39 11 1 1 9 13 1 1 11 11 11 11 11 2 11 11 1 9 11 11 2 11 11 11 11 11 7 0 11 2 11 2 9 11 11 11 11 14 13 2
15 15 1 11 11 1 9 1 0 9 13 9 1 9 13 2
17 3 11 1 9 2 9 1 9 1 0 9 1 14 9 13 4 2
27 11 11 11 1 11 11 11 11 7 11 11 11 11 1 1 9 13 9 1 0 9 1 9 2 9 13 2
23 11 2 11 2 9 11 11 1 13 13 4 4 16 11 11 11 14 15 9 1 9 13 2
14 15 1 15 14 9 1 1 1 13 1 0 14 13 2
10 11 1 9 15 15 1 13 4 4 2
17 9 9 11 11 1 9 13 4 16 11 9 1 15 9 14 13 2
23 9 1 13 13 16 11 1 9 1 11 15 9 13 1 3 9 7 9 9 1 9 13 2
28 9 1 1 12 9 1 11 2 11 2 1 0 9 7 11 9 1 0 9 13 2 15 11 1 9 13 4 2
32 15 1 11 11 1 9 9 11 11 7 9 9 1 9 11 11 11 1 1 11 13 7 11 1 1 9 13 1 9 0 13 2
16 11 1 13 16 11 1 15 9 1 9 13 1 9 13 4 2
19 15 1 11 1 11 1 0 9 11 11 11 7 0 11 9 1 9 13 2
25 11 1 9 1 9 9 1 9 1 1 11 2 11 2 1 0 9 1 9 1 0 9 13 4 2
27 15 13 16 3 12 9 1 1 11 2 11 2 9 1 9 13 7 15 1 12 9 1 1 11 9 13 2
20 15 13 16 9 9 1 9 1 11 2 11 2 1 12 9 1 9 13 4 2
30 15 13 16 11 2 11 2 1 11 1 15 9 9 1 9 13 4 7 15 11 13 2 7 11 1 11 11 11 13 2
21 3 11 11 11 7 11 11 11 1 9 1 11 1 13 9 1 0 9 13 4 2
22 11 1 13 16 15 11 2 11 2 9 9 1 9 13 7 9 1 15 9 14 13 2
28 16 11 1 9 13 16 11 1 15 9 1 1 0 9 13 4 2 15 11 2 11 2 0 9 1 9 13 2
30 11 11 1 9 1 9 9 9 1 11 9 1 11 1 11 7 11 11 1 12 0 9 9 1 1 11 0 13 4 2
37 9 9 1 0 9 9 11 1 0 9 9 1 0 9 11 11 1 11 11 1 9 1 0 9 1 13 4 1 9 13 1 3 11 0 13 4 2
15 9 1 9 1 1 11 11 11 11 1 0 13 4 4 2
18 9 1 1 9 1 9 13 4 16 11 1 0 9 9 15 9 13 2
33 15 1 9 1 11 11 11 1 9 13 4 16 11 1 0 9 1 9 1 13 1 9 1 0 9 9 1 1 11 0 13 4 2
39 10 9 1 11 1 11 1 9 1 9 0 13 4 2 7 9 1 9 1 1 9 1 13 1 3 9 9 9 1 0 9 9 1 1 11 0 13 4 2
14 9 9 1 11 1 11 11 1 1 9 0 13 4 2
27 11 1 13 4 4 16 11 11 9 11 11 7 11 11 11 11 1 11 11 1 0 9 1 9 1 13 2
29 9 1 1 11 10 0 13 7 15 0 9 13 4 4 16 10 9 1 11 1 0 9 1 9 1 13 4 4 2
23 11 1 0 9 1 9 1 13 4 1 9 9 9 1 9 1 11 11 1 14 13 4 2
33 9 9 9 11 11 1 9 1 1 1 9 1 9 13 4 16 11 1 14 9 1 1 13 4 4 7 15 9 1 14 13 4 2
38 10 9 9 9 9 1 9 1 13 11 1 9 1 1 3 10 9 1 13 4 2 10 9 1 9 9 9 1 14 11 1 11 11 1 13 4 4 2
30 9 1 10 9 1 12 9 1 14 11 1 0 9 1 13 4 1 9 0 13 4 7 9 9 1 11 0 13 4 2
30 9 1 13 16 11 1 9 9 1 14 11 11 11 1 11 11 11 7 9 9 1 0 9 11 11 1 9 13 4 2
13 15 0 13 4 16 11 11 11 1 9 1 13 2
26 9 1 1 11 0 13 1 3 11 1 9 1 1 13 4 12 12 1 9 14 0 13 13 4 4 2
28 9 1 0 12 12 1 9 1 9 1 11 1 13 4 16 15 12 9 1 0 9 1 9 1 13 4 4 2
28 11 9 11 11 7 15 9 11 11 1 9 1 9 1 11 11 1 9 11 11 9 1 0 9 13 4 4 2
39 9 9 1 15 3 0 7 0 9 1 11 1 9 11 11 11 1 13 13 16 16 10 9 9 1 13 4 7 9 9 13 4 16 15 15 9 14 13 2
35 11 1 11 11 11 11 11 11 1 9 1 15 13 11 1 15 13 4 16 15 15 11 1 15 9 13 1 0 13 15 15 3 13 4 2
10 3 13 2 2 15 14 9 13 4 2
23 11 9 1 9 11 1 13 16 15 1 1 15 14 9 15 9 7 11 1 14 13 4 2
13 9 1 9 1 9 13 13 11 9 1 13 4 2
22 15 13 2 2 15 14 15 9 13 4 2 7 15 9 1 9 1 0 14 9 13 2
12 9 2 9 7 0 9 9 1 9 13 4 4
29 9 1 11 1 10 9 1 9 13 16 9 1 0 9 9 13 14 14 0 9 2 9 7 9 0 13 13 4 2
23 9 1 9 1 1 0 13 1 9 1 9 9 1 13 14 2 16 11 1 13 4 4 2
8 10 9 9 9 1 14 13 2
38 9 2 9 12 9 9 13 9 1 9 9 1 9 14 13 4 4 2 7 3 15 0 9 1 9 13 1 0 13 4 2 15 13 1 14 9 13 2
47 11 1 13 16 15 11 0 15 12 9 1 9 1 9 1 1 15 9 13 4 15 15 10 9 10 0 13 4 16 9 13 4 9 9 1 9 13 1 1 9 13 1 10 9 13 4 2
16 11 11 1 11 1 13 0 9 1 9 0 2 0 13 4 2
16 0 9 1 1 9 2 9 9 7 0 9 1 0 9 13 2
28 11 7 3 1 9 1 13 0 9 1 1 9 9 7 9 10 9 9 1 13 4 4 2 15 9 0 13 2
29 11 11 1 9 1 1 0 2 0 9 1 12 9 1 9 13 4 7 11 1 12 9 1 13 4 1 9 13 2
12 10 3 12 9 1 10 9 0 14 13 4 2
24 15 1 11 11 1 9 11 9 1 9 0 9 1 1 9 1 0 9 1 12 9 13 4 2
17 9 1 12 9 1 10 9 0 13 4 15 9 1 9 0 13 2
19 11 1 0 9 11 9 12 9 9 13 2 15 9 1 12 9 10 13 2
11 9 9 1 9 9 13 4 13 4 4 2
16 9 9 1 13 13 16 10 9 0 12 9 0 13 4 4 2
30 11 1 11 9 11 11 11 1 13 13 16 9 1 1 9 10 0 13 4 4 7 14 10 9 9 1 13 4 4 2
19 11 2 11 7 11 11 1 11 13 1 10 9 10 9 1 13 4 4 2
26 11 2 11 9 1 13 1 14 10 9 9 15 0 9 1 12 9 1 1 12 9 1 9 1 13 2
14 11 9 9 1 10 0 7 0 9 0 14 13 4 2
18 9 9 1 13 0 9 1 1 12 9 1 10 13 0 13 4 4 2
20 9 1 9 1 13 1 1 12 9 1 9 9 1 9 9 13 4 4 4 2
19 11 11 1 9 1 13 4 16 9 1 1 15 12 9 1 9 13 4 2
22 11 11 11 11 11 1 0 12 9 1 13 16 14 10 9 9 9 1 13 4 4 2
24 11 13 1 12 9 1 0 13 4 4 2 7 11 1 11 13 4 12 9 1 11 13 4 2
14 9 1 14 9 0 13 1 9 9 14 13 4 4 2
17 0 9 9 11 11 7 11 11 1 14 0 9 1 9 13 4 2
19 9 1 9 1 1 0 9 1 9 1 1 1 9 9 1 13 4 4 2
42 11 11 11 2 11 2 11 11 11 2 11 2 11 11 2 11 2 11 11 11 2 11 11 2 11 2 11 11 14 12 9 1 1 12 9 1 9 1 13 4 4 2
30 11 11 1 11 9 1 1 11 1 9 1 0 9 13 1 1 11 9 1 1 9 1 9 1 13 12 9 0 13 2
17 9 14 12 9 1 9 14 13 1 1 9 9 13 14 13 4 2
13 10 3 9 14 12 12 9 12 9 15 13 4 2
9 10 9 15 0 9 0 13 4 2
25 0 9 15 9 1 9 1 1 13 14 13 16 11 11 9 1 12 0 9 9 1 13 4 4 2
11 9 9 1 1 12 9 1 14 13 4 2
11 10 9 0 9 14 0 9 1 13 4 2
10 15 0 9 1 9 14 0 13 4 2
13 9 1 9 1 13 9 1 0 9 1 9 13 2
12 11 9 11 7 9 9 11 1 9 0 13 2
10 9 0 9 9 1 9 13 4 4 2
28 11 9 9 13 14 10 9 7 9 13 16 9 1 11 1 1 1 13 4 7 13 4 10 9 0 13 4 2
10 15 13 9 1 14 9 13 4 4 2
21 15 13 13 10 9 1 15 12 9 1 1 9 7 9 1 9 13 11 13 4 2
27 0 9 1 13 4 11 1 13 16 11 1 9 12 1 11 1 9 1 13 4 4 16 9 0 14 13 2
21 15 13 4 16 9 7 11 15 9 13 7 15 9 1 15 11 13 1 9 13 2
26 11 1 12 9 1 9 1 11 13 12 9 1 15 1 9 7 9 13 1 10 9 13 4 4 4 2
59 0 9 1 13 4 11 1 11 1 13 16 11 1 9 1 11 1 1 10 0 9 13 4 4 7 15 15 13 14 4 4 7 15 11 1 9 13 7 14 11 1 10 3 1 13 1 9 13 4 15 15 10 9 1 0 14 13 4 2
44 11 1 13 16 15 9 1 0 9 13 4 4 2 7 3 14 15 9 1 15 9 13 16 15 11 13 4 4 15 15 9 11 9 1 1 13 1 0 9 14 13 4 4 2
28 11 1 13 16 11 13 1 9 13 15 9 1 9 1 14 9 13 4 7 9 1 15 13 1 9 13 4 2
40 9 1 9 11 1 0 9 1 13 16 11 1 9 1 9 1 11 1 9 1 15 14 0 14 13 4 4 15 15 13 16 15 9 1 14 15 14 13 4 2
43 16 2 2 11 11 11 11 11 11 2 1 9 1 1 10 9 11 11 11 11 11 1 9 1 0 13 4 4 15 2 11 2 0 11 1 12 0 9 1 0 13 4 2
16 10 9 1 9 9 11 11 7 15 9 11 11 1 13 4 2
13 0 9 1 10 9 14 12 12 0 9 1 13 2
38 9 1 13 9 1 1 1 9 1 9 1 9 1 9 1 0 13 4 9 1 13 4 16 0 9 1 0 13 1 1 9 1 9 1 0 9 13 2
23 15 1 14 9 1 13 16 0 9 1 1 1 9 1 9 1 14 9 0 13 4 4 2
14 16 11 9 1 1 1 15 9 1 3 9 13 4 2
27 11 9 1 3 9 12 9 14 9 1 9 1 13 4 4 3 10 9 9 12 9 14 9 13 4 4 2
22 0 13 16 9 11 2 11 1 9 1 9 0 9 1 14 12 12 9 10 13 4 2
21 11 1 13 16 9 1 0 9 1 0 13 1 1 9 9 1 15 9 14 13 2
13 16 0 9 1 9 13 1 9 13 4 4 4 2
9 7 15 1 12 9 9 13 4 2
16 10 3 11 1 12 12 9 9 9 1 1 9 0 13 4 2
24 11 1 13 16 9 1 0 12 9 1 13 0 9 1 1 1 9 1 9 1 0 9 13 2
23 15 13 16 10 9 1 9 1 9 12 12 9 1 0 9 1 13 12 12 9 13 4 2
26 15 13 16 9 9 1 1 13 4 9 1 1 0 9 1 15 9 1 9 13 1 15 9 14 13 2
15 9 1 13 0 9 1 9 1 11 11 1 9 0 13 2
14 11 11 1 10 3 9 9 1 0 0 9 0 13 2
15 15 9 11 2 11 1 1 12 9 1 9 13 4 4 2
15 9 1 1 0 9 1 12 12 9 9 9 1 9 13 2
32 11 1 0 9 1 12 0 9 9 1 12 0 9 9 1 9 1 15 1 9 13 7 12 12 9 9 13 1 9 13 4 2
17 0 9 11 1 11 1 11 1 15 9 11 1 9 1 9 13 2
25 9 1 9 9 1 9 7 12 0 9 1 1 11 0 13 9 1 1 12 9 11 13 4 4 2
12 9 1 15 1 15 1 9 14 13 4 4 2
35 9 1 0 9 1 9 13 4 16 11 1 12 9 9 1 12 0 9 11 1 11 11 1 15 9 13 0 13 4 7 3 15 9 13 2
33 9 1 9 0 13 11 13 11 11 11 11 11 11 1 13 16 9 1 1 9 1 9 1 12 12 9 9 13 1 14 9 13 2
14 15 1 1 11 0 0 9 1 9 13 4 4 4 2
14 15 15 9 11 11 7 11 9 1 12 9 1 13 2
15 10 9 1 15 12 0 9 9 1 13 4 1 9 13 2
33 9 9 13 1 15 9 1 9 7 9 11 1 15 12 9 13 4 7 13 16 10 9 15 9 7 11 9 11 1 1 0 13 2
18 0 9 11 1 12 9 13 15 15 0 9 1 0 9 13 9 13 2
14 9 1 0 13 4 1 3 11 1 15 1 9 13 2
12 0 9 9 15 9 11 13 1 0 13 4 2
40 0 13 16 11 1 12 0 9 1 1 9 1 9 1 0 14 9 11 11 11 1 11 1 12 9 9 9 1 9 11 11 11 1 12 9 1 9 13 4 2
23 11 11 11 11 11 1 9 1 11 1 13 9 1 0 9 15 9 1 14 13 4 4 2
17 11 1 11 9 1 13 4 10 9 1 10 9 0 13 4 4 2
10 10 9 1 10 9 1 9 14 13 2
25 7 9 1 1 1 11 1 9 9 11 11 1 13 16 9 1 9 13 4 1 15 9 14 13 2
18 15 13 13 16 15 14 0 13 16 9 1 15 9 14 13 4 4 2
21 11 1 9 13 4 16 11 1 11 11 7 11 1 9 1 15 9 1 9 13 2
15 11 11 11 1 10 9 1 0 9 1 9 13 4 4 2
22 11 1 9 9 11 11 1 9 1 9 13 4 13 16 11 11 11 1 9 0 13 2
19 10 9 1 10 9 1 9 14 13 16 11 1 9 1 9 15 13 4 2
15 15 13 16 14 15 0 9 1 9 1 9 14 13 4 2
14 0 9 1 10 9 1 9 10 9 1 14 13 4 2
18 0 13 16 15 1 10 9 9 1 1 1 12 0 9 13 4 4 2
22 10 9 1 13 4 4 16 11 11 1 11 9 1 11 1 9 1 9 14 13 4 2
13 15 11 11 9 9 1 9 1 13 9 13 4 2
12 7 16 9 14 13 16 9 1 9 13 15 2
15 11 1 13 4 16 11 11 11 1 9 1 9 13 4 2
18 9 9 1 0 9 1 9 1 11 9 1 0 9 1 9 13 4 2
10 9 1 0 9 1 1 13 4 4 2
14 11 9 1 14 15 13 4 4 16 0 9 0 13 2
13 15 11 9 1 9 1 9 1 9 13 4 4 2
30 11 11 1 0 9 9 1 11 1 0 0 9 11 11 11 2 11 2 11 11 11 11 9 1 11 11 1 0 13 2
19 11 1 10 9 1 0 9 1 9 1 11 1 0 13 1 9 13 4 2
11 11 1 9 11 11 1 11 1 0 13 2
14 11 11 11 15 9 1 11 11 1 0 9 9 13 2
19 15 1 1 11 1 13 16 15 11 1 12 9 1 15 9 1 0 13 2
10 3 10 9 9 11 11 1 13 4 2
20 7 0 9 1 9 1 9 1 13 9 1 1 15 12 9 1 1 13 4 2
13 3 1 9 1 1 11 1 12 9 13 4 4 2
25 7 3 1 11 11 11 1 10 9 1 9 13 4 16 11 1 12 9 1 9 1 0 13 4 2
14 15 13 16 15 1 1 12 9 1 1 9 13 4 2
27 11 9 1 9 1 13 16 11 1 3 9 2 9 2 9 7 9 7 9 1 0 9 1 9 13 4 2
11 7 15 9 1 9 1 13 4 4 4 2
23 10 9 9 1 11 1 12 10 0 9 11 7 9 1 14 0 9 11 11 14 0 13 2
20 0 9 9 1 9 0 13 1 1 13 4 4 9 1 13 9 13 4 4 2
29 9 1 0 9 1 9 1 9 1 1 13 1 9 1 11 1 0 9 13 4 9 1 15 9 1 9 13 4 2
38 9 1 11 11 11 1 14 15 9 1 0 13 4 4 2 7 11 1 9 1 1 15 0 9 9 11 2 11 2 1 10 9 1 12 9 14 13 2
12 9 11 1 9 1 0 13 4 1 9 13 2
54 11 9 11 11 1 9 1 11 9 1 11 1 13 9 1 13 4 16 0 9 10 9 1 0 13 4 7 15 0 9 13 16 0 9 1 15 1 13 1 9 1 9 1 13 4 4 16 9 1 15 15 9 13 2
18 7 11 1 0 9 9 11 2 11 2 1 10 9 1 13 9 13 2
13 11 11 1 13 13 16 15 9 1 9 1 13 2
9 0 9 1 9 1 9 13 4 2
15 16 9 1 9 1 9 13 4 16 15 9 1 1 13 2
34 11 9 1 1 11 0 9 1 9 11 11 11 1 9 13 16 9 1 1 10 9 9 3 13 2 15 11 2 11 2 14 0 13 2
34 11 1 0 9 15 13 16 10 0 9 1 0 0 9 1 1 14 9 1 9 13 4 2 7 0 9 1 15 1 0 9 14 13 2
21 9 1 9 13 4 16 9 1 9 1 0 13 4 1 11 10 9 1 9 13 2
13 11 1 13 13 16 15 9 1 9 0 14 13 2
23 0 9 1 13 4 4 10 9 15 13 15 9 10 9 1 13 15 0 0 9 1 13 2
41 10 3 11 11 1 11 11 1 9 1 9 1 13 16 15 9 1 9 1 10 9 13 4 2 15 9 13 4 4 7 9 1 9 1 9 13 1 9 13 4 2
22 9 1 9 1 9 13 1 1 11 11 11 11 1 9 1 9 13 1 9 13 4 2
15 15 1 10 9 7 9 1 9 1 9 1 9 13 4 2
21 11 11 11 11 11 13 4 16 9 1 10 9 1 9 1 1 0 13 4 4 2
15 16 9 15 15 9 13 4 16 9 15 10 0 9 13 2
21 15 9 1 0 9 1 1 13 4 7 0 9 1 0 9 0 13 1 0 13 2
27 11 1 1 11 11 13 1 1 15 11 11 11 1 9 1 14 9 1 9 13 1 1 0 13 4 4 2
22 9 1 13 13 11 1 1 12 9 13 1 1 10 9 1 15 0 9 14 14 13 2
28 11 1 9 1 9 1 9 14 0 13 4 4 2 7 15 10 9 1 9 1 1 9 1 9 14 13 4 2
19 9 1 9 14 9 13 1 1 9 1 9 14 0 9 1 0 14 13 2
14 9 1 9 10 9 1 9 1 14 13 4 4 4 2
16 15 9 14 9 7 9 1 14 12 9 1 0 13 4 4 2
12 9 1 9 13 9 1 9 0 13 4 4 2
34 0 9 1 9 1 3 13 1 3 11 1 15 9 1 13 9 1 13 1 1 11 11 7 11 11 11 2 11 2 1 9 13 4 2
31 11 1 11 1 0 13 9 1 9 7 0 9 1 1 14 0 9 1 13 1 1 0 9 1 9 1 9 1 9 13 2
24 11 0 11 11 11 1 9 1 10 12 0 9 1 11 1 1 1 9 13 1 9 13 4 2
18 9 1 1 10 9 1 9 13 4 4 4 16 10 9 1 9 13 2
9 10 9 1 9 9 0 13 4 2
40 9 1 10 9 1 14 9 13 4 16 11 11 1 11 11 11 2 11 2 1 11 1 9 1 11 1 9 0 9 1 1 12 12 9 13 1 9 13 4 2
23 10 9 1 9 9 9 7 9 1 9 1 13 4 16 9 1 3 9 9 13 4 4 2
21 10 9 11 11 1 9 1 0 9 1 9 9 1 0 13 1 9 13 4 4 2
43 0 13 16 11 11 9 11 11 1 11 1 13 4 16 15 11 1 0 13 4 16 11 11 1 13 9 9 1 13 9 1 13 1 1 15 10 9 1 9 1 9 13 2
13 9 1 1 11 1 12 12 1 10 9 13 4 2
12 11 1 11 11 1 9 1 9 13 4 4 2
19 11 11 1 13 4 16 11 9 1 1 13 4 1 9 9 13 4 4 2
24 9 1 13 16 11 11 11 2 11 2 1 11 1 9 9 1 9 1 1 0 9 13 4 2
15 11 9 1 1 9 13 11 1 14 9 13 1 0 13 2
15 11 11 0 9 1 0 11 9 9 9 1 9 1 13 2
11 15 1 11 11 1 12 9 11 1 13 2
26 15 1 11 1 12 0 9 0 9 11 2 11 7 11 1 12 2 12 9 9 1 9 13 4 4 2
11 11 11 11 11 1 1 9 13 4 4 2
16 9 1 9 13 16 9 0 9 1 9 13 1 9 14 13 2
31 0 11 11 11 11 1 0 11 9 1 13 4 11 11 7 11 1 10 9 1 9 13 4 15 9 7 9 9 13 4 2
25 9 1 9 13 16 11 1 9 1 1 9 1 9 0 13 1 1 9 9 1 9 13 4 4 2
23 0 13 16 9 11 1 0 0 11 11 11 11 13 4 15 11 1 9 1 9 13 4 2
23 12 0 9 1 13 13 16 11 1 9 1 1 10 9 1 9 13 1 1 0 9 13 2
16 9 1 9 1 0 9 13 1 1 0 9 13 4 4 4 2
30 11 11 11 1 11 1 11 11 1 9 13 1 10 9 1 0 11 1 11 9 1 12 9 1 9 13 4 4 4 2
12 9 1 15 1 0 9 1 13 14 4 4 2
38 10 9 1 9 1 11 1 9 1 1 10 9 1 9 13 2 15 1 11 1 9 11 9 1 1 0 13 7 11 11 1 9 13 1 9 13 4 2
24 12 10 9 1 13 16 9 11 1 9 1 1 9 1 13 1 15 0 9 9 13 4 4 2
25 15 11 2 11 1 15 14 9 1 9 1 9 13 11 1 9 1 9 13 1 9 13 4 4 2
13 11 2 11 1 9 9 1 9 13 4 4 4 2
12 10 10 9 1 9 1 9 13 4 4 4 2
23 11 9 11 11 1 11 1 11 1 9 7 11 11 2 11 2 9 11 11 1 9 13 2
22 12 9 1 11 1 0 9 1 11 1 9 13 1 1 0 9 1 9 2 9 13 2
25 11 1 1 12 9 1 9 1 1 9 1 9 1 13 16 15 11 1 9 1 9 2 9 13 2
20 0 9 1 10 9 13 11 2 11 1 9 13 1 1 9 9 1 9 13 2
12 11 9 9 10 9 11 2 11 1 13 4 2
18 10 9 1 11 1 9 1 13 4 9 1 1 0 13 4 4 4 2
18 15 9 1 11 1 13 4 16 11 11 1 11 15 9 13 4 4 2
15 15 1 11 1 11 1 10 9 1 15 9 13 4 4 2
19 16 2 11 11 1 0 11 1 13 16 9 1 15 1 15 9 14 13 2
11 11 0 9 13 7 15 15 9 13 4 2
14 15 13 16 11 9 1 10 9 1 9 7 9 13 2
20 16 11 2 11 2 9 11 11 3 1 9 1 9 1 1 9 13 4 4 2
30 9 1 11 1 9 13 1 1 11 2 11 2 11 2 9 9 1 1 1 15 13 16 15 9 9 0 9 0 13 2
13 10 9 10 9 1 9 0 13 1 9 1 13 2
33 9 14 1 0 9 1 13 4 0 9 1 9 1 13 1 1 11 11 11 11 1 9 9 1 0 11 11 1 11 1 9 13 2
8 15 9 11 9 11 11 13 2
33 11 11 11 11 9 11 11 1 9 1 13 10 9 9 1 9 1 0 9 1 9 1 13 1 1 0 9 1 9 2 9 13 2
14 9 11 1 11 11 11 1 3 13 1 0 14 13 2
12 12 9 13 14 4 16 0 15 13 4 4 2
21 15 11 11 1 11 11 11 11 11 1 13 12 9 1 9 1 9 13 4 4 2
22 11 1 11 1 13 4 9 1 12 0 9 1 0 9 1 0 13 1 9 13 4 2
20 11 1 9 1 0 13 4 11 1 11 9 1 0 13 4 1 9 13 4 2
27 10 3 11 11 1 11 1 9 1 11 1 9 1 0 13 4 13 4 16 9 1 3 13 4 4 4 2
39 11 1 11 11 1 11 1 13 9 1 9 9 9 2 11 11 11 2 11 11 11 11 1 11 11 1 9 9 9 1 9 1 0 13 1 9 13 4 2
13 11 11 11 2 11 1 9 1 1 9 1 13 2
27 11 1 11 11 11 1 12 10 0 9 11 11 1 14 11 11 1 11 9 1 0 13 1 9 13 4 2
17 9 1 15 1 9 13 14 0 9 1 9 1 9 13 4 4 2
24 11 1 13 4 16 11 1 0 9 1 0 9 11 1 9 9 1 0 9 1 13 4 4 2
12 11 11 1 10 9 9 1 12 9 1 13 2
29 11 11 11 11 11 1 11 1 11 9 1 11 11 1 0 2 0 9 1 0 7 0 9 13 1 9 13 4 2
21 15 13 16 11 9 1 13 1 9 9 9 1 1 9 9 1 9 1 0 13 2
15 11 1 9 1 15 0 13 4 4 16 15 0 14 13 2
18 11 2 11 2 1 14 11 1 11 9 1 13 4 1 9 13 4 2
24 11 1 9 1 9 13 4 13 4 16 15 11 1 9 13 4 2 7 15 15 9 14 13 2
28 15 13 16 15 11 1 9 1 15 9 14 13 2 16 15 1 12 9 1 1 9 9 1 9 13 4 4 2
13 15 13 16 9 1 10 9 1 0 9 13 4 2
38 10 3 9 9 1 9 0 13 13 4 16 11 1 11 11 1 11 11 11 1 0 13 4 4 4 7 15 11 11 1 0 13 1 15 9 14 13 2
20 11 11 11 11 15 9 9 9 2 11 2 1 13 1 9 1 13 4 4 2
15 11 11 1 10 12 11 1 9 1 9 1 9 13 4 2
17 9 1 9 11 1 9 1 13 9 1 13 9 1 3 13 4 2
23 15 11 11 1 13 13 16 9 1 9 13 1 10 9 1 15 1 15 9 14 13 4 2
17 9 1 1 11 11 1 10 9 11 11 1 9 1 12 9 13 2
15 15 9 1 9 7 15 10 9 9 13 1 9 13 4 2
20 9 1 1 15 10 9 1 0 9 1 9 1 9 1 13 4 1 9 13 2
37 9 1 12 9 1 1 10 9 1 9 1 15 13 1 14 9 13 15 0 9 11 2 11 1 1 1 13 4 9 1 15 9 1 9 13 4 2
22 11 11 11 11 1 1 11 1 11 2 11 1 9 13 1 9 14 13 15 9 13 2
19 11 11 1 13 16 11 11 11 1 9 1 9 9 13 1 9 14 13 2
9 15 13 16 9 9 1 9 13 2
6 15 15 1 14 13 2
9 15 9 13 1 9 14 14 13 2
27 12 9 9 9 1 9 1 1 11 11 11 1 9 11 11 11 1 9 1 9 1 9 1 9 13 4 2
9 11 1 15 13 4 15 0 13 2
12 3 14 9 12 9 13 15 9 13 13 4 2
23 11 11 1 0 7 0 9 1 9 1 9 1 1 11 11 9 9 1 1 0 14 13 2
15 11 11 11 1 13 13 16 9 1 9 1 10 9 13 2
20 10 9 1 9 13 15 0 13 1 1 11 0 9 14 13 1 1 0 13 2
19 7 9 1 1 11 11 1 1 1 15 1 1 15 9 0 14 13 4 2
19 9 1 1 2 11 11 1 9 1 13 1 0 9 1 9 12 12 13 2
10 15 11 1 13 12 12 1 13 4 2
12 15 1 11 11 10 9 1 13 0 14 13 2
34 11 11 1 1 2 0 9 9 1 11 2 11 2 11 9 9 1 1 10 0 9 1 9 1 1 0 9 13 1 9 13 4 4 2
14 9 1 0 9 1 9 1 13 4 14 10 9 13 2
15 7 11 11 1 15 1 15 1 1 15 9 14 13 4 2
20 11 11 11 11 11 11 1 1 2 9 1 9 1 0 9 11 11 1 13 2
25 7 11 11 11 1 9 2 9 13 15 9 9 1 9 1 1 0 9 0 13 1 1 0 13 2
15 9 1 0 7 0 9 1 9 1 3 9 13 4 4 2
10 0 9 10 9 1 13 10 0 13 2
22 15 13 13 16 11 11 16 15 10 9 1 9 13 16 15 10 9 13 4 4 4 2
19 9 11 1 9 9 9 1 12 9 12 12 0 9 1 9 13 13 4 2
16 3 11 1 9 1 0 9 1 9 1 13 9 1 9 13 2
13 9 9 1 9 1 1 1 15 9 14 13 4 2
15 11 9 9 1 9 11 1 9 1 9 0 13 4 4 2
18 9 1 9 1 1 0 9 13 4 2 7 9 1 15 9 13 4 2
50 13 4 4 16 11 9 9 0 11 11 11 1 0 9 1 13 1 12 0 11 9 11 0 9 1 12 9 1 1 9 1 1 13 15 3 1 0 12 9 11 1 13 15 9 1 13 0 13 4 2
22 9 1 9 10 9 13 15 0 9 1 9 1 13 16 12 9 11 1 13 13 4 2
9 9 1 9 1 13 9 13 4 2
17 9 9 1 9 1 9 9 1 9 11 7 9 1 9 1 13 2
21 11 1 9 1 9 9 1 9 1 1 13 4 7 9 9 9 1 13 9 13 2
13 9 11 1 15 1 1 9 7 9 1 9 13 2
28 15 1 9 11 1 9 1 1 13 4 7 10 9 15 9 1 11 9 9 13 7 9 1 9 1 0 13 2
17 9 1 9 13 14 9 1 9 13 9 1 9 9 9 13 4 2
18 10 9 1 11 9 9 1 9 11 1 9 1 9 0 13 4 4 2
18 9 1 9 13 16 9 10 9 1 9 0 13 1 9 13 4 4 2
15 3 11 9 9 9 9 11 1 9 1 12 9 9 13 2
7 9 1 9 1 9 13 2
19 0 9 1 9 1 9 1 1 1 11 1 13 16 15 9 1 9 13 2
10 9 12 10 9 1 9 1 13 4 2
24 11 1 11 1 11 7 11 9 1 9 13 4 13 16 15 10 9 1 9 1 9 14 13 2
23 3 9 9 9 11 11 1 14 9 7 0 9 1 9 7 9 1 0 13 1 9 13 2
30 11 11 11 1 12 0 9 1 9 1 9 1 11 1 12 9 0 13 0 9 1 9 1 9 1 0 9 13 4 2
13 11 1 13 16 15 9 1 12 10 9 13 4 2
26 9 1 15 14 13 4 16 9 9 9 7 11 9 9 1 1 0 7 0 9 1 0 13 4 4 2
11 15 1 11 1 9 9 9 1 9 13 2
30 10 9 1 11 1 9 9 9 11 11 1 10 9 7 9 14 1 0 9 1 9 7 9 1 0 13 1 9 13 2
25 9 9 9 2 9 9 1 0 9 1 1 11 11 11 11 11 1 9 9 1 1 0 13 4 2
7 9 1 12 9 0 13 2
17 9 9 1 1 9 2 11 2 11 2 1 11 1 9 13 4 2
14 9 1 9 1 9 9 1 9 13 1 9 13 4 2
17 11 11 1 0 9 1 0 9 9 1 11 11 1 9 13 4 2
19 0 11 1 9 1 9 1 1 9 1 9 14 13 4 7 3 9 13 2
13 9 1 9 1 1 9 1 9 12 9 0 13 2
37 15 1 14 15 9 1 9 14 13 15 9 1 9 1 11 1 12 9 1 0 13 4 4 7 15 1 9 1 13 0 9 1 9 1 3 13 2
21 9 1 0 9 9 1 3 11 1 0 11 11 11 11 11 11 1 9 13 4 2
26 15 1 9 9 13 14 0 9 1 9 1 11 11 11 11 11 1 9 1 13 4 7 9 13 4 2
34 15 11 1 9 11 11 1 12 9 13 4 11 11 1 9 1 9 13 2 15 9 1 13 16 15 1 9 1 9 14 13 4 4 2
10 15 13 16 9 1 0 14 13 4 2
21 15 1 9 1 9 1 0 9 9 13 7 15 0 13 1 9 13 9 13 4 2
28 10 3 9 9 1 11 11 1 0 9 9 11 2 11 1 9 9 11 11 7 0 9 11 11 14 13 4 2
33 3 12 9 1 9 11 11 11 1 13 1 3 14 15 9 14 13 15 9 1 9 1 9 12 9 12 9 1 1 0 13 4 2
31 9 9 11 11 14 12 9 9 1 13 9 1 1 14 13 2 7 9 13 0 9 9 2 9 0 13 1 0 14 13 2
21 15 1 14 0 9 1 14 13 1 3 9 1 9 12 9 1 1 0 13 4 2
18 14 12 9 12 9 3 14 9 1 9 9 13 14 9 9 13 4 2
30 15 1 9 1 13 16 9 0 14 13 7 11 1 14 0 13 9 1 13 1 9 13 2 7 0 9 9 13 4 2
37 15 1 9 11 11 1 0 9 1 0 13 1 9 13 7 9 1 15 9 13 4 11 1 12 9 1 9 1 0 9 1 0 13 1 9 13 2
20 15 1 14 15 0 9 1 9 0 13 15 9 1 0 9 1 13 3 13 2
29 9 11 1 1 11 1 12 9 1 9 9 0 9 1 13 4 1 15 0 12 9 1 12 9 1 9 13 4 2
8 12 9 12 14 9 1 13 2
9 10 9 1 12 9 0 13 4 2
16 9 1 12 1 9 0 13 1 15 11 11 8 13 4 4 2
13 0 9 1 11 1 0 9 1 9 13 4 4 2
18 9 1 9 13 14 11 1 9 9 7 11 9 9 9 1 13 4 2
17 9 1 12 9 1 9 1 9 9 1 1 9 0 13 4 4 2
33 0 9 1 1 11 9 9 11 1 12 14 9 1 12 9 9 1 9 11 1 9 1 9 1 0 9 1 9 13 13 4 4 2
26 9 9 11 1 10 3 13 4 16 3 1 13 4 12 9 1 13 1 9 1 9 9 9 13 4 2
12 15 1 9 1 9 0 9 1 9 13 4 2
25 9 10 0 13 16 12 9 1 9 1 14 9 13 4 2 7 9 1 0 0 9 0 13 4 2
9 15 11 7 11 9 2 9 13 2
33 10 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 7 11 0 13 4 2
30 10 9 1 9 1 0 9 13 2 15 9 1 11 2 11 2 11 7 11 1 9 0 13 11 2 11 8 13 4 2
10 9 1 9 13 9 9 1 13 4 2
32 9 1 9 1 9 1 1 9 1 13 13 2 7 9 1 9 13 1 9 13 4 7 9 1 9 13 4 0 9 13 4 2
12 9 1 9 1 13 16 15 3 9 13 4 2
20 15 1 15 15 1 0 14 13 4 7 15 15 1 1 9 14 13 13 4 2
19 9 1 9 1 9 1 9 1 9 1 1 1 13 9 1 13 4 4 2
17 10 9 1 9 13 9 1 9 1 9 0 9 1 13 4 4 2
16 3 14 10 9 9 11 1 13 3 10 9 1 9 13 4 2
9 9 9 11 0 11 13 4 4 2
17 11 11 11 2 11 2 1 11 1 0 0 9 1 9 13 4 2
43 11 1 13 13 16 3 9 1 10 0 9 1 14 9 9 1 9 13 4 4 7 0 9 9 1 9 2 9 13 4 4 4 3 11 12 9 1 1 1 3 13 4 2
23 9 1 1 11 1 1 9 1 10 9 1 0 9 1 9 7 15 9 1 9 13 4 2
21 15 1 2 9 10 9 1 0 9 1 0 13 1 0 9 1 14 10 9 13 2
18 10 9 9 1 0 9 1 0 9 1 9 13 1 9 13 4 4 2
31 0 11 11 11 1 9 9 1 11 11 2 11 11 11 11 11 1 2 11 11 11 11 11 2 1 1 1 13 4 4 2
15 9 1 10 9 1 11 11 1 12 9 1 9 13 4 2
24 10 9 1 11 9 11 11 2 11 9 11 11 7 11 2 11 11 11 11 11 11 0 13 2
23 11 1 11 11 11 11 11 1 9 1 1 15 13 12 0 9 1 12 9 1 0 13 2
11 10 9 1 9 1 3 9 13 4 4 2
13 10 9 1 9 11 1 12 0 9 1 13 4 2
27 0 9 1 9 1 1 1 11 13 1 3 11 1 11 1 11 11 0 9 1 13 12 9 1 0 13 2
22 11 9 9 1 9 11 11 1 13 16 10 9 1 9 12 1 12 9 1 1 13 2
15 11 1 13 16 9 0 9 1 13 0 9 1 13 4 2
26 9 1 3 9 13 1 1 1 1 15 13 16 15 10 9 13 15 9 1 9 1 0 9 13 4 2
10 9 9 1 9 1 9 13 4 4 2
12 15 1 9 1 9 1 9 13 1 9 13 2
15 11 11 11 2 11 2 1 11 1 11 1 0 9 13 2
38 10 9 1 12 9 1 11 15 1 13 11 1 11 1 11 9 1 9 13 4 4 2 15 0 13 4 16 11 1 1 15 0 2 0 9 14 13 2
12 15 2 11 1 9 13 1 9 14 14 13 2
12 10 9 15 1 15 10 12 9 13 4 4 2
24 11 15 15 12 9 1 1 2 11 11 2 1 12 7 12 9 1 9 1 9 13 4 4 2
16 11 1 9 13 16 9 1 9 12 2 12 9 1 13 4 2
32 16 11 11 1 9 9 1 13 12 9 1 9 1 1 0 9 1 9 0 13 1 3 0 9 1 9 14 13 4 4 4 2
13 15 9 15 9 1 13 7 15 9 1 3 13 2
37 15 13 16 11 1 15 9 1 9 1 9 13 4 2 7 15 15 9 1 9 0 13 4 4 15 15 9 1 0 13 4 7 15 9 9 13 2
13 15 12 9 1 9 13 2 15 1 12 0 13 2
16 11 1 9 1 9 1 11 1 9 13 1 9 0 13 4 2
21 11 1 11 1 12 9 7 12 9 1 15 9 1 13 15 9 9 12 13 4 2
16 7 2 12 9 1 11 1 1 15 1 0 9 0 13 4 2
20 11 1 15 9 9 13 4 7 0 9 13 1 15 9 1 13 4 1 13 2
16 3 1 11 7 11 1 9 13 16 9 1 9 3 13 4 2
16 7 15 9 14 13 1 1 15 9 1 1 1 13 4 4 2
47 11 1 11 11 11 11 2 11 11 11 11 7 11 11 11 7 0 11 9 11 11 1 10 0 9 1 9 13 1 1 11 1 9 11 1 9 7 11 11 11 11 11 1 9 13 4 2
36 9 9 1 13 13 9 1 1 11 11 11 1 0 9 11 11 1 9 15 0 9 1 13 16 15 11 1 15 9 1 15 9 0 13 4 2
29 15 13 16 15 11 11 11 1 9 9 9 1 13 4 9 1 12 9 1 11 1 15 9 1 9 0 13 4 2
17 0 13 16 11 9 9 9 1 15 3 1 9 1 13 4 4 2
28 11 1 9 1 13 16 15 15 9 11 1 1 11 11 11 1 9 13 15 9 1 12 12 9 0 13 4 2
25 15 15 14 9 13 16 15 15 12 9 1 11 11 11 1 10 9 1 12 12 9 0 13 4 2
29 7 11 1 11 1 9 11 0 11 11 1 9 1 13 4 4 9 1 1 1 15 14 9 1 9 1 9 13 2
32 9 9 1 11 1 9 1 13 4 16 11 1 9 1 12 12 9 0 13 4 4 7 15 1 14 15 9 1 13 4 4 2
29 15 1 9 1 9 1 15 14 13 4 16 11 1 9 11 1 11 11 1 9 1 12 12 9 0 13 4 4 2
26 9 9 1 11 1 10 12 12 9 1 1 1 14 9 13 15 11 1 1 9 9 9 13 4 4 2
14 10 9 1 9 1 12 9 1 1 9 13 4 4 2
14 10 9 11 7 15 9 1 11 1 9 1 13 4 2
40 9 1 12 0 9 1 0 9 1 9 1 3 9 13 1 3 11 11 9 9 11 11 1 9 2 9 9 1 9 1 13 14 9 9 1 3 9 13 4 2
18 15 13 16 10 0 9 9 2 9 7 9 1 9 1 13 4 4 2
23 11 11 1 1 13 9 1 15 13 16 9 9 1 9 9 1 9 1 10 14 9 13 2
30 9 11 1 0 11 2 11 2 11 1 13 4 9 1 0 9 1 9 1 12 0 9 1 9 1 9 13 4 4 2
41 11 11 7 11 1 0 9 1 1 13 4 9 1 9 1 0 13 4 11 11 11 1 9 1 0 9 1 1 9 1 0 9 1 0 13 1 9 13 4 4 2
27 9 1 13 4 4 16 9 1 9 1 13 9 1 15 9 1 1 0 2 0 9 14 13 4 4 4 2
28 12 9 1 10 9 1 9 11 1 13 4 16 15 10 10 9 13 15 9 1 9 1 1 9 0 13 4 2
24 10 9 14 10 9 9 1 0 9 14 13 4 4 2 16 11 1 9 1 9 13 4 4 2
20 14 12 9 1 13 4 9 1 13 4 16 3 0 9 9 9 1 9 13 2
9 9 1 14 9 10 14 0 13 2
13 11 9 1 12 9 1 14 12 9 13 4 4 2
12 15 9 13 4 4 2 15 14 10 9 13 2
9 9 1 0 9 1 0 9 13 2
11 12 9 1 9 1 9 3 0 13 4 2
33 13 1 10 9 1 14 15 1 13 16 9 9 7 9 1 9 9 1 9 1 13 1 1 13 9 1 13 9 0 13 4 4 2
23 15 1 9 9 15 9 7 9 1 1 9 1 0 9 1 1 13 1 0 13 4 4 2
16 10 9 14 9 1 9 14 15 0 9 1 15 13 4 4 2
20 15 1 0 9 0 9 1 9 13 4 9 2 9 1 9 1 13 4 4 2
21 9 1 13 4 4 16 9 9 1 9 1 1 9 1 9 1 14 9 13 4 2
25 9 1 15 9 1 13 4 2 15 10 14 9 1 13 13 16 9 13 1 15 10 9 13 4 2
32 10 9 11 1 1 1 9 13 1 0 13 4 4 4 2 7 10 9 1 11 1 9 1 13 1 9 0 13 4 4 4 2
25 11 1 13 16 10 9 1 14 9 7 9 1 0 9 13 4 4 2 16 9 1 13 4 4 2
17 15 1 9 9 1 9 9 1 9 1 10 9 7 9 13 4 2
20 9 1 9 11 1 9 1 0 13 1 1 9 9 1 9 9 13 4 4 2
12 9 13 1 1 1 12 9 0 13 4 4 2
13 11 1 9 1 9 1 15 9 1 0 13 4 2
14 9 1 11 1 9 1 1 9 13 9 13 4 4 2
33 0 9 11 1 13 9 1 13 0 9 9 11 11 1 9 9 1 9 1 9 7 9 9 1 9 13 13 9 9 1 0 13 2
22 9 1 9 1 0 7 0 9 1 1 9 13 3 9 1 1 13 1 0 9 13 2
21 9 9 1 9 13 1 9 1 9 1 13 16 9 9 1 1 14 9 0 13 2
14 9 1 13 16 9 1 9 1 9 1 0 9 13 2
15 11 1 9 1 1 9 1 9 1 1 12 9 0 13 2
24 11 1 0 9 9 7 9 9 11 11 1 9 1 9 1 9 13 1 1 1 9 13 4 2
13 9 1 10 3 14 9 1 12 9 1 14 13 2
7 9 13 15 13 4 4 2
18 11 11 1 11 11 11 1 13 4 16 9 1 0 9 11 1 13 2
21 11 11 1 11 11 11 11 1 9 13 1 3 9 1 9 1 1 10 9 13 2
23 11 1 13 16 11 15 9 9 13 7 12 0 9 13 1 1 15 9 1 9 13 4 2
26 15 13 16 9 1 10 9 13 4 15 9 1 0 9 1 9 1 9 1 13 3 1 0 13 4 2
25 11 1 9 1 11 11 11 11 11 1 11 1 11 11 11 11 1 9 13 1 9 13 4 4 2
29 11 11 1 13 4 16 15 9 9 9 1 13 4 4 15 1 15 0 9 1 9 13 1 9 14 14 13 4 2
21 11 1 1 16 11 1 9 13 4 16 9 1 12 12 9 9 0 0 13 4 2
37 11 11 1 11 1 11 1 11 9 1 9 13 1 9 1 11 11 11 2 11 2 7 11 11 11 11 1 15 9 12 9 1 13 1 9 13 2
35 11 1 9 1 13 1 1 1 11 1 1 9 0 13 4 1 13 11 9 1 3 9 1 9 1 9 13 1 9 1 10 9 0 13 2
20 9 1 13 16 12 9 1 11 11 9 9 7 11 11 11 15 9 0 13 2
15 7 9 1 9 14 13 2 15 9 1 9 1 9 13 2
28 0 9 1 9 1 1 0 9 1 9 0 13 1 11 0 9 11 11 9 1 9 2 9 11 1 13 4 2
36 11 1 10 9 1 12 9 1 9 1 11 1 9 1 1 9 13 7 9 1 0 0 9 1 9 13 1 1 12 0 9 0 13 4 4 2
29 9 1 1 11 1 11 11 1 11 1 13 4 11 11 1 1 13 4 9 1 9 1 10 10 9 13 4 4 2
26 10 9 1 11 11 11 11 2 11 2 1 9 1 9 14 1 13 4 9 1 12 9 13 4 4 2
12 15 1 12 9 1 11 1 0 13 4 4 2
11 11 1 11 11 11 1 11 1 9 13 2
27 11 7 11 1 9 1 1 9 1 0 0 9 11 0 9 1 10 9 1 0 13 1 0 9 13 4 2
20 11 14 9 1 1 9 2 9 7 0 0 9 1 9 1 1 9 13 4 2
34 15 9 9 1 9 13 4 7 9 1 9 0 13 4 7 15 1 11 1 9 1 9 13 1 11 1 0 9 1 1 9 13 4 2
25 11 9 1 1 9 1 9 13 1 3 11 11 0 13 4 4 2 15 15 9 13 4 4 4 2
19 10 9 1 9 1 0 9 11 1 11 1 11 1 0 13 4 4 4 2
23 11 1 9 11 7 9 11 11 1 14 10 9 1 0 13 1 9 1 0 13 4 4 2
13 11 7 11 9 1 13 4 9 1 14 13 4 2
26 11 1 2 9 9 9 2 11 11 11 11 11 2 11 2 1 12 9 1 13 0 9 1 9 13 2
27 15 9 1 1 11 2 11 2 11 2 11 7 0 9 9 1 0 9 1 9 13 1 1 9 13 4 2
17 11 7 11 1 1 11 11 7 11 11 1 14 10 9 13 4 2
18 9 1 1 11 0 9 1 9 11 1 11 7 0 9 1 13 4 2
24 11 1 10 9 1 3 9 13 4 4 7 15 15 7 9 1 0 9 1 13 4 4 4 2
14 9 1 9 9 0 11 11 1 9 13 1 9 13 2
27 9 1 13 16 0 9 1 11 1 0 9 1 9 13 1 9 9 10 9 9 1 9 13 1 9 13 2
20 15 9 11 1 11 11 1 11 11 11 1 11 1 9 1 13 13 4 4 2
21 9 1 9 13 16 0 9 11 11 1 12 9 1 9 1 0 13 1 9 13 2
43 9 1 9 1 9 11 1 11 1 11 1 0 9 13 4 13 16 15 1 10 9 1 0 9 13 16 9 0 9 1 0 13 9 2 11 13 2 9 13 13 4 4 2
25 15 13 16 9 1 9 1 9 1 9 1 10 9 1 13 4 4 16 10 9 1 9 13 4 2
13 11 1 13 16 10 9 1 9 11 1 13 4 2
13 0 13 16 11 11 11 11 11 1 9 14 13 2
16 11 1 13 16 11 11 11 1 10 15 14 9 1 9 13 2
14 11 1 11 1 11 11 11 1 13 1 9 13 4 2
31 9 9 11 11 1 13 13 16 11 1 9 1 9 7 12 9 9 1 9 1 9 1 11 0 9 1 9 13 4 4 2
17 11 1 15 9 1 9 1 11 1 11 9 1 9 14 13 4 2
14 11 9 1 13 16 11 14 13 16 11 1 13 4 2
12 15 10 9 1 9 1 0 9 13 13 4 2
27 11 11 1 11 1 11 11 1 1 11 1 11 11 11 1 9 9 13 1 9 1 9 1 3 9 13 2
28 11 11 1 9 11 11 11 1 13 16 11 1 0 9 1 9 1 13 4 1 1 9 9 13 1 9 13 2
20 9 9 11 11 1 14 11 1 9 1 15 13 9 13 16 10 9 0 13 2
22 15 13 16 11 1 11 11 1 9 13 1 1 14 13 15 10 9 1 9 13 4 2
44 9 11 11 11 2 11 11 11 2 11 11 11 2 11 11 7 11 11 1 12 0 9 1 1 11 1 13 16 11 1 0 9 1 9 13 1 9 13 9 1 9 13 4 2
40 0 9 1 11 11 2 11 2 7 11 9 1 9 1 9 13 4 15 13 16 11 1 0 9 13 9 1 9 2 9 7 9 1 9 1 13 1 9 13 2
22 11 11 2 11 2 7 11 9 1 9 9 13 1 11 11 1 9 1 0 13 4 2
49 11 1 9 1 1 13 16 11 11 1 3 2 3 10 9 13 4 16 0 9 1 13 4 0 9 1 0 9 1 9 1 9 13 1 1 15 0 9 1 9 1 12 10 9 13 1 9 13 2
22 15 13 16 11 11 15 0 9 7 9 1 9 9 1 9 13 1 13 14 13 4 2
37 15 13 16 11 11 1 15 9 1 11 11 1 0 9 1 13 4 16 9 1 9 1 9 1 1 0 9 1 0 9 1 9 13 4 4 4 2
21 11 11 1 11 1 13 15 0 9 1 11 1 13 16 9 10 0 13 4 4 2
46 11 1 13 16 11 1 13 4 9 1 9 1 1 11 11 1 11 11 1 3 9 1 9 13 7 9 1 0 9 1 13 4 15 9 11 11 11 11 11 11 1 13 1 9 13 2
44 9 9 13 1 11 11 1 9 1 9 1 1 1 9 1 13 4 1 15 13 16 15 0 9 1 13 15 9 15 9 13 4 15 15 13 4 4 16 15 10 9 13 4 2
28 9 11 1 11 1 12 9 1 15 9 1 9 13 9 13 4 7 3 1 15 1 14 9 13 9 13 4 2
15 9 1 9 13 9 9 1 9 1 9 9 13 4 4 2
11 9 1 12 0 9 14 0 13 4 4 2
14 9 1 9 1 1 11 1 0 9 1 13 4 4 2
10 15 1 15 15 1 14 9 13 4 2
10 15 9 1 9 1 14 9 13 4 2
17 11 1 1 13 9 1 9 1 1 1 9 1 9 1 0 13 2
12 9 1 15 1 1 11 9 9 1 9 13 2
22 9 9 1 9 1 13 12 9 1 9 13 4 9 1 1 11 1 0 9 1 13 2
33 9 1 1 11 1 11 9 11 11 11 9 1 9 9 1 9 13 1 9 11 1 9 13 4 7 9 14 15 9 13 4 4 2
17 15 9 13 1 11 1 9 1 11 1 9 11 1 13 4 4 2
15 7 11 12 9 3 11 11 1 1 9 1 13 4 4 2
38 9 1 9 1 15 1 1 11 1 9 9 7 9 9 1 9 13 0 9 1 1 9 13 1 9 13 4 2 7 9 1 9 1 9 13 4 4 2
13 9 2 9 9 13 1 3 0 11 13 4 4 2
11 9 1 9 1 10 9 1 0 13 4 2
31 10 9 1 13 9 1 9 14 13 4 7 9 1 10 9 1 0 9 13 4 9 1 0 13 1 9 0 13 4 4 2
22 15 1 9 1 9 1 11 1 11 1 0 9 11 1 15 9 1 15 13 4 4 2
12 11 0 12 9 1 10 9 1 13 4 4 2
16 11 1 11 1 13 4 1 11 11 15 13 1 9 13 4 2
27 13 4 4 4 16 11 11 1 12 9 1 14 11 1 13 1 9 13 4 2 7 9 14 13 4 4 2
14 11 11 1 13 16 11 15 1 15 9 13 4 4 2
25 10 9 1 1 1 15 11 1 9 13 9 13 4 7 3 1 15 1 9 13 4 9 13 4 2
26 11 9 11 11 1 9 0 13 1 1 9 1 0 9 11 11 1 9 1 11 1 9 13 4 4 2
22 9 1 9 11 11 1 13 16 9 1 12 9 1 9 11 1 9 13 4 4 4 2
20 11 1 13 16 15 9 0 13 1 1 11 1 12 9 1 9 13 4 4 2
31 15 13 16 16 11 0 9 1 1 9 2 13 9 1 9 14 13 4 16 15 9 1 0 13 1 9 13 4 4 4 2
15 15 13 11 1 1 11 1 9 13 9 1 9 13 4 2
12 15 10 9 1 9 1 9 1 9 13 4 2
17 15 1 11 1 9 1 9 1 11 1 9 1 0 13 4 4 2
32 11 1 9 1 11 1 9 1 11 11 2 11 1 10 9 0 14 13 7 15 0 9 13 4 9 13 1 9 13 4 4 2
8 11 11 11 1 0 11 13 2
13 15 11 1 9 13 1 9 0 9 1 0 13 2
9 15 11 1 9 1 9 13 4 2
16 9 1 10 9 1 11 11 11 1 9 11 1 9 13 4 2
20 0 9 1 9 9 1 9 1 13 11 11 1 11 9 13 0 14 14 13 2
12 11 1 11 1 9 1 12 9 1 9 13 2
23 12 9 1 13 9 1 15 1 9 14 13 1 0 9 1 1 11 9 0 13 4 4 2
16 15 1 12 9 1 13 9 1 9 11 1 0 13 4 4 2
15 10 12 9 1 11 11 1 11 1 10 12 9 13 4 2
15 15 11 2 11 1 12 9 7 11 1 12 9 0 13 2
12 10 9 15 0 9 1 12 9 10 13 4 2
11 0 9 1 1 12 9 1 9 13 4 2
11 7 0 9 1 11 1 12 9 13 4 2
10 11 1 0 9 1 12 9 13 4 2
10 11 15 0 9 1 13 1 0 13 2
8 11 1 14 12 9 13 4 2
18 11 1 10 9 10 12 9 13 4 7 0 9 1 12 9 13 4 2
22 11 1 9 11 1 3 14 15 12 9 1 9 13 4 15 0 9 1 14 13 4 2
15 10 9 1 10 9 11 2 11 9 11 11 1 13 4 2
15 15 12 9 1 11 1 1 11 9 1 1 1 0 13 2
16 0 9 13 1 3 11 1 13 16 0 9 15 0 9 13 2
24 13 4 4 16 11 1 15 9 9 1 9 13 4 7 11 11 1 11 9 1 9 13 4 2
22 11 9 7 11 11 11 11 11 1 9 9 13 4 11 1 10 0 9 1 9 13 2
17 15 11 1 9 1 9 1 0 9 1 0 9 1 9 13 4 2
15 11 1 13 9 1 11 3 0 9 1 1 1 13 4 2
20 11 1 9 13 7 15 12 9 9 13 1 9 1 11 1 0 13 4 4 2
9 15 9 11 9 1 1 1 13 2
19 9 9 1 1 11 1 9 1 15 2 15 1 9 1 9 9 13 4 2
13 11 1 13 13 16 11 1 1 0 9 13 4 2
18 16 11 14 11 2 11 2 11 11 1 13 16 9 9 10 0 13 2
12 15 11 1 15 11 1 9 1 9 13 4 2
12 16 11 7 0 9 1 15 9 13 4 4 2
24 11 1 13 16 15 0 11 1 9 1 16 11 2 11 1 9 13 4 16 9 10 0 13 2
37 11 1 9 7 0 11 11 11 16 11 1 9 13 4 4 7 11 1 12 9 9 13 1 11 11 11 11 1 9 11 11 10 9 0 13 4 2
10 15 11 2 11 1 11 11 1 13 2
58 10 9 11 11 9 1 13 11 11 2 11 2 2 11 11 2 11 2 2 11 11 11 2 11 2 2 11 11 2 11 2 2 11 11 11 2 11 2 2 11 11 2 11 2 7 9 11 11 11 2 11 11 2 0 13 4 4 2
49 0 9 1 13 1 1 9 11 9 11 11 11 2 11 2 2 11 9 7 11 1 9 11 11 11 2 11 2 2 11 1 0 9 11 11 2 11 2 7 9 11 9 11 11 2 11 2 13 2
16 9 1 1 1 9 9 1 9 3 0 0 13 4 4 4 2
23 9 9 15 15 0 13 4 4 16 9 1 0 9 13 1 1 0 9 13 3 0 13 2
22 9 1 13 13 16 0 9 14 13 1 1 1 9 1 0 9 14 13 4 4 4 2
12 0 9 1 1 14 12 12 9 1 9 13 2
23 11 11 11 11 11 11 11 11 11 11 14 0 9 9 1 3 9 13 1 9 1 13 2
24 9 9 1 9 1 1 9 1 9 13 1 1 11 11 1 11 9 11 11 1 9 13 4 2
17 11 1 15 0 9 0 13 9 9 1 9 13 1 1 13 4 2
18 7 2 9 3 14 9 9 1 12 12 12 9 0 13 1 9 13 2
20 15 9 13 16 9 9 9 9 1 9 1 9 1 3 14 15 9 13 4 2
24 11 11 11 1 13 4 1 11 11 11 1 9 9 9 1 1 1 9 1 9 13 4 4 2
13 11 1 13 16 9 0 9 1 9 1 13 4 2
16 11 11 11 1 0 9 1 13 0 13 1 9 0 13 4 2
13 10 9 12 12 9 9 9 0 13 4 4 4 2
24 9 1 9 13 16 0 9 1 9 1 12 12 9 9 9 0 13 1 9 0 13 4 4 2
15 9 0 13 1 12 9 14 9 1 9 13 1 9 13 2
24 15 1 9 1 0 0 2 0 9 1 9 0 13 1 9 0 13 1 9 13 4 4 4 2
17 9 0 9 1 1 9 1 9 0 13 1 14 9 13 4 4 2
21 11 11 3 9 1 9 13 1 9 9 1 10 0 9 1 9 13 4 4 4 2
11 10 9 1 15 9 1 9 14 13 4 2
21 15 1 11 11 10 9 1 9 1 2 11 11 11 11 2 0 13 4 4 4 2
17 9 9 1 9 1 13 4 11 11 10 9 9 13 4 4 4 2
17 11 11 1 9 2 11 11 11 11 2 1 10 9 13 4 4 2
26 9 1 1 15 9 1 14 12 9 9 1 9 13 2 7 14 12 9 9 9 1 9 13 4 4 2
27 15 1 9 1 13 0 3 10 9 1 9 13 4 4 4 2 15 9 1 1 3 9 1 9 13 4 2
18 10 2 11 11 11 11 2 1 1 0 0 9 1 9 9 13 4 2
21 10 9 1 10 9 1 9 13 4 16 15 9 1 9 1 10 14 10 9 13 2
21 9 1 9 1 10 9 1 13 4 16 15 13 0 9 1 10 14 10 9 13 2
9 10 9 1 10 14 10 9 13 2
27 11 11 11 11 1 9 11 11 1 1 10 9 1 9 1 10 14 10 12 1 12 9 9 13 4 4 2
18 15 13 16 10 9 11 1 2 11 11 11 11 2 0 13 4 4 2
31 10 9 1 0 9 1 10 9 9 1 10 0 0 9 1 13 4 2 15 10 14 10 12 9 9 1 9 13 4 4 2
21 10 9 1 10 9 0 9 1 0 13 2 16 9 1 9 1 9 0 13 4 2
15 15 1 10 0 2 0 9 1 1 15 0 13 4 4 2
28 9 1 9 1 15 1 9 14 1 10 9 1 15 9 1 9 9 1 9 13 15 9 1 3 10 13 4 2
13 15 15 9 14 12 12 9 1 9 13 4 4 2
11 15 12 10 9 13 15 15 1 13 4 2
16 9 9 1 9 13 1 1 15 10 9 1 10 9 14 13 2
19 11 11 2 11 11 2 11 11 7 11 11 1 9 10 9 15 1 13 2
12 9 9 11 1 9 11 14 3 11 1 13 2
32 0 9 1 9 9 11 11 11 13 4 16 11 2 11 2 11 7 11 14 10 9 1 1 14 0 9 1 9 13 13 4 2
7 11 1 15 14 14 13 2
8 11 1 14 15 14 13 4 2
21 13 0 13 16 0 9 1 9 1 1 9 1 1 13 1 9 14 13 4 4 2
9 16 15 0 9 1 13 4 4 2
16 11 1 9 11 3 0 13 7 15 1 0 15 9 1 13 2
21 9 11 9 9 1 11 13 4 4 7 10 9 9 9 1 9 13 1 13 4 2
11 11 1 9 9 1 1 1 15 13 4 2
17 15 9 1 10 9 15 9 1 9 1 14 13 1 1 8 13 2
22 3 14 10 9 15 10 9 15 12 9 1 0 0 11 1 13 1 14 13 4 4 2
9 11 1 1 11 1 14 9 13 2
10 15 15 15 3 13 1 13 4 4 2
13 11 1 15 15 1 1 11 1 13 11 11 13 2
13 15 13 1 9 9 1 13 9 9 1 13 4 2
10 7 0 13 1 1 15 10 9 13 2
12 3 11 1 1 15 0 9 13 14 0 13 2
11 9 1 11 15 1 1 9 13 4 4 2
13 11 7 11 1 14 11 1 9 1 13 13 4 2
20 11 1 9 11 11 11 11 1 1 14 15 9 11 1 1 11 13 4 4 2
10 0 11 9 1 0 9 13 4 4 2
16 11 1 14 15 9 1 1 0 9 1 0 9 13 4 4 2
14 7 9 1 0 9 11 1 9 1 9 10 14 13 2
31 11 1 9 1 12 9 1 1 13 4 4 7 11 0 9 1 15 1 13 4 14 3 14 10 9 1 9 13 9 13 2
19 9 9 11 1 9 11 14 3 9 11 7 9 11 1 1 11 1 13 2
28 9 1 9 11 1 11 1 1 12 11 11 13 4 7 15 15 15 1 9 1 1 0 9 9 1 14 13 2
32 9 1 9 1 9 11 0 12 9 9 1 11 9 9 13 4 1 12 9 1 9 13 4 7 12 0 9 1 0 13 4 2
20 15 1 1 11 2 9 9 2 11 11 1 13 16 9 9 14 12 9 13 2
8 10 9 9 9 1 1 13 2
13 9 1 9 0 13 1 1 9 3 14 13 4 2
22 12 9 1 9 1 0 13 4 4 4 7 9 1 11 11 11 1 9 13 4 4 2
18 11 11 1 11 11 11 1 13 16 9 0 9 1 13 4 4 4 2
16 0 9 1 13 4 9 1 9 9 1 1 3 1 0 13 2
11 9 13 1 9 1 9 14 13 4 4 2
11 10 9 1 1 9 1 9 13 4 4 2
14 9 1 9 1 1 11 11 11 1 0 13 4 4 2
11 9 1 12 9 7 12 9 14 0 13 2
19 9 1 13 16 10 9 1 9 13 0 9 9 9 9 1 13 4 4 2
16 11 11 1 9 1 9 1 9 1 15 9 3 13 4 4 2
13 9 1 15 0 13 1 9 1 9 13 4 4 2
22 9 1 12 0 9 1 1 0 9 9 1 11 1 9 9 1 15 0 9 14 13 2
15 11 1 11 11 1 1 11 11 1 13 9 9 1 13 2
20 9 9 11 11 11 1 15 9 9 1 9 13 14 11 11 1 9 13 4 2
15 15 9 1 15 0 9 13 7 15 9 9 1 13 4 2
20 11 9 1 14 9 13 1 9 14 13 7 9 14 13 1 9 1 13 4 2
14 11 1 11 11 1 9 13 7 9 1 9 0 13 2
21 7 9 15 0 13 4 15 9 11 1 11 1 9 1 0 9 1 9 9 13 2
12 9 10 9 1 9 13 1 1 0 13 4 2
12 11 11 1 11 1 1 13 11 9 0 13 2
18 11 11 9 13 4 2 7 15 9 3 3 9 1 9 13 4 4 2
18 0 13 1 3 1 0 9 11 1 11 11 1 1 1 15 13 4 2
12 9 1 10 9 1 9 1 9 13 4 4 2
9 15 15 9 9 14 0 13 4 2
58 0 13 16 11 9 1 9 1 9 0 13 1 11 11 1 11 9 1 9 13 4 4 7 15 9 1 11 9 1 1 15 11 11 11 7 11 11 1 1 15 9 1 13 1 1 13 4 15 15 11 1 9 1 9 13 4 4 2
34 0 12 9 1 11 7 11 1 0 11 9 1 13 4 0 9 1 1 11 11 11 1 0 9 1 9 9 15 9 1 13 4 4 2
29 14 12 9 1 1 10 9 11 1 9 9 1 10 9 14 12 9 9 13 1 1 9 9 1 9 13 4 4 2
15 11 1 0 9 1 1 15 13 4 9 1 9 13 4 2
14 11 1 13 4 9 1 14 15 9 1 3 9 13 2
42 3 2 10 0 9 1 10 9 9 9 1 1 14 9 9 1 3 1 1 11 11 11 11 11 11 2 11 1 1 1 0 0 9 1 9 13 1 0 9 13 4 2
15 10 9 9 9 1 13 1 1 3 9 1 13 4 4 2
11 15 9 1 11 11 11 0 13 4 4 2
13 15 1 11 1 0 0 9 1 9 13 4 4 2
31 15 13 16 3 1 1 10 9 1 1 10 9 14 11 11 11 1 0 9 13 1 1 9 9 1 9 13 4 4 4 2
15 15 0 9 1 9 13 10 9 9 1 9 13 13 4 2
23 9 1 9 9 1 1 10 9 1 0 9 9 1 13 10 9 1 1 15 0 9 13 2
10 10 9 15 0 9 1 1 1 13 2
27 15 13 16 11 11 11 11 1 0 9 1 1 9 0 0 9 1 15 9 13 1 9 14 13 4 4 2
14 9 1 10 9 0 9 1 0 9 1 9 13 4 2
29 15 3 0 9 1 15 9 13 1 9 13 2 3 9 1 0 9 1 13 0 9 1 15 13 1 14 9 13 2
31 15 13 16 10 9 9 1 9 13 1 1 11 1 0 9 1 1 14 12 9 9 11 11 11 1 9 1 9 13 4 2
21 11 11 9 11 11 1 13 16 0 9 14 15 10 9 1 0 9 1 13 4 2
14 9 7 0 9 1 15 1 9 1 0 9 13 4 2
14 11 11 1 13 16 9 1 0 9 1 9 13 4 2
21 15 13 16 11 11 11 11 11 11 2 11 10 9 12 9 1 9 13 4 4 2
33 9 1 9 9 1 1 0 9 1 14 9 13 4 2 15 0 9 7 9 9 1 9 13 4 7 9 9 1 14 0 9 13 2
29 11 11 11 11 11 11 1 9 9 11 11 11 1 13 16 10 9 9 1 11 7 11 11 1 0 9 13 4 2
15 10 9 11 11 11 1 9 9 1 1 13 4 4 4 2
23 15 13 16 11 11 1 11 11 1 9 1 1 1 12 9 1 9 9 13 4 4 4 2
18 11 1 11 11 11 1 11 11 11 13 1 9 9 1 13 4 4 2
19 16 9 1 9 13 4 4 16 10 9 11 9 1 0 13 4 4 4 2
28 15 13 16 14 12 9 1 1 11 9 1 13 9 1 1 9 9 1 1 0 9 1 9 14 13 4 4 2
17 11 9 11 11 1 13 0 9 1 0 9 1 9 13 4 4 2
18 0 9 1 1 13 10 0 9 1 15 3 9 9 1 9 13 4 2
21 11 0 9 9 1 0 10 9 1 9 9 13 15 3 0 13 1 9 13 4 2
27 11 11 11 11 11 11 1 11 1 13 9 1 9 1 0 9 13 4 15 3 0 13 1 9 13 4 2
24 11 11 11 1 10 9 1 0 13 4 11 1 0 9 9 1 1 15 9 11 1 13 4 2
24 11 9 11 11 1 14 11 1 9 11 1 13 9 1 13 4 16 15 10 9 1 0 13 2
19 15 11 1 9 13 4 16 9 1 10 9 1 15 15 9 1 1 13 2
13 15 11 1 3 0 13 4 1 9 0 13 4 2
14 0 11 11 11 11 1 10 9 1 0 9 13 4 2
10 11 1 11 1 10 0 13 4 4 2
15 11 1 9 13 1 9 13 14 11 9 1 9 13 4 2
17 9 1 0 10 9 1 9 9 13 15 3 0 13 1 9 13 2
20 11 9 1 15 9 1 3 0 13 1 1 11 11 1 9 9 13 4 4 2
17 15 9 3 1 13 11 13 11 1 11 11 13 11 1 9 13 2
7 15 9 1 12 9 13 2
19 15 13 16 9 1 9 11 1 9 1 9 1 1 0 9 13 4 4 2
15 11 9 11 11 1 11 1 3 0 13 1 9 13 4 2
20 11 1 12 0 9 13 4 15 13 4 16 9 1 15 1 9 1 9 13 2
29 16 15 13 4 16 9 1 9 9 0 13 7 11 1 0 9 1 13 1 1 13 4 4 2 16 15 0 13 2
12 9 15 0 7 0 9 1 9 13 4 4 2
16 9 1 15 9 13 1 0 9 1 9 1 15 0 9 13 2
9 9 2 9 2 1 13 4 4 2
8 15 9 2 9 2 13 4 2
37 11 1 11 11 11 1 9 1 9 1 13 12 9 1 11 11 11 11 1 9 11 1 15 10 9 0 13 15 9 1 10 0 9 3 13 4 2
29 9 1 1 10 9 9 1 9 1 9 1 10 7 0 0 13 4 1 10 9 1 9 10 9 1 13 4 4 2
26 15 13 16 15 13 0 9 13 16 0 9 1 14 9 9 1 1 9 1 9 13 4 13 4 4 2
19 9 11 1 9 11 1 0 9 9 1 0 9 1 14 0 9 13 4 2
22 9 1 13 4 4 16 14 12 1 12 9 1 14 9 1 15 0 9 13 4 4 2
24 15 9 0 10 9 1 3 14 13 4 4 4 2 15 1 1 3 0 9 13 14 14 4 2
25 15 13 16 0 0 9 9 1 13 10 9 1 9 9 1 0 13 1 1 14 13 4 4 4 2
28 9 0 13 1 10 9 1 10 9 1 0 13 4 4 7 15 9 9 9 1 0 0 9 1 13 4 4 2
13 15 9 1 9 1 0 9 10 0 13 4 4 2
11 9 1 9 13 12 0 9 13 4 4 2
24 15 9 0 9 0 13 4 4 7 0 9 1 9 1 12 9 14 15 1 13 14 4 4 2
51 11 11 11 1 9 1 0 12 9 1 9 13 4 9 11 1 13 16 9 1 0 9 14 13 1 1 14 11 1 9 1 12 9 1 1 11 11 11 11 1 0 9 1 9 3 13 14 4 4 4 2
21 7 0 13 4 1 9 1 9 1 14 9 1 9 1 9 10 9 9 13 4 2
66 15 9 1 0 9 1 9 1 13 4 1 13 4 1 9 1 1 9 7 9 1 9 1 1 1 0 9 1 9 1 0 9 1 14 0 13 7 15 3 13 1 1 9 9 1 1 14 9 1 15 9 7 9 1 13 1 9 1 0 13 4 1 9 14 13 2
21 9 9 1 9 1 11 11 11 7 9 11 1 9 1 9 1 1 3 9 13 2
36 9 1 9 1 11 1 1 9 13 1 9 13 4 11 2 11 1 1 13 9 9 1 9 1 9 1 9 13 2 15 11 1 0 9 13 2
28 11 1 13 13 16 11 1 15 14 9 1 1 9 14 13 4 7 9 9 9 2 9 1 9 1 0 13 2
41 9 1 9 1 1 10 9 1 13 4 0 11 11 7 11 9 11 11 1 13 16 10 9 13 4 4 16 11 1 15 9 9 1 9 13 4 10 9 13 4 2
17 15 13 13 16 15 11 1 10 9 15 9 1 1 13 4 4 2
58 15 0 11 1 13 9 1 1 9 11 11 1 10 9 1 14 9 13 15 13 4 4 16 11 11 11 11 1 9 1 9 1 11 1 3 2 3 9 1 13 4 4 16 15 7 14 11 1 3 13 7 14 0 9 1 0 13 2
38 11 1 13 16 0 9 10 9 1 0 9 14 13 4 7 9 9 1 9 1 0 9 1 1 9 1 9 9 1 0 9 1 1 14 13 4 4 2
31 15 14 1 11 1 11 11 0 13 4 7 15 11 1 9 13 4 13 16 15 9 9 1 10 9 1 0 13 4 4 2
14 15 9 13 16 9 1 11 1 1 9 13 4 4 2
10 15 1 9 9 1 9 0 13 4 2
36 9 1 1 1 11 11 11 11 11 11 1 13 16 11 15 1 1 9 1 13 4 4 16 10 9 0 9 7 0 9 2 9 1 0 13 2
13 15 1 9 9 1 14 15 9 14 13 4 4 2
20 15 13 16 9 16 15 1 9 13 13 4 2 16 9 9 1 1 0 13 2
19 11 11 1 13 16 0 9 15 14 9 1 15 9 0 13 1 0 13 2
17 7 15 9 15 14 13 16 15 15 9 1 9 0 13 4 4 2
19 11 1 16 15 0 13 16 15 15 3 15 9 1 1 1 13 4 4 2
40 11 1 9 1 11 9 1 10 14 9 13 16 10 9 1 10 9 9 1 14 13 4 4 2 15 0 9 9 1 0 0 9 1 1 0 9 13 4 4 2
15 11 9 1 11 1 9 9 11 11 1 0 0 9 13 2
8 10 9 12 0 9 1 13 2
25 11 9 11 11 11 1 10 9 1 11 1 9 11 11 11 7 0 9 11 11 1 9 1 13 2
13 9 1 9 1 11 11 1 13 1 9 13 4 2
10 11 10 9 11 1 11 11 1 13 2
19 11 1 13 16 9 13 1 1 15 11 1 9 11 11 11 1 13 4 2
38 9 1 9 13 4 9 9 11 11 11 1 10 9 1 9 0 13 4 16 11 15 14 11 9 1 13 7 15 1 11 9 1 9 0 13 4 4 2
42 16 11 1 9 11 1 0 9 1 9 13 2 7 11 1 15 13 4 15 9 1 13 4 16 16 10 9 0 9 1 9 13 4 4 16 15 9 0 13 4 4 2
43 0 9 11 11 1 9 13 16 11 1 11 9 9 1 11 1 9 1 9 13 4 4 7 15 1 0 9 0 14 13 4 4 15 1 15 9 1 9 13 0 14 13 2
32 11 1 11 1 9 11 1 10 9 1 0 13 4 15 13 4 4 16 11 1 10 9 1 13 4 1 1 15 9 13 4 2
21 16 2 9 9 1 9 1 13 4 16 0 9 1 1 11 0 9 13 4 4 2
40 0 9 11 11 11 1 0 9 13 1 3 15 11 1 9 1 13 1 9 13 4 7 13 16 9 10 9 1 7 11 1 9 1 9 1 11 1 9 13 2
17 9 1 9 13 4 1 1 11 1 11 1 9 1 0 13 4 2
21 0 13 16 9 9 9 1 11 1 9 1 11 1 0 9 1 9 0 13 4 2
44 13 4 4 16 11 1 12 11 9 1 1 11 9 9 1 15 9 9 13 4 7 3 1 15 0 9 1 9 9 9 1 1 0 13 4 15 10 9 1 11 9 13 4 2
27 11 11 11 11 1 13 16 9 1 0 9 1 9 13 1 1 9 9 1 9 13 1 9 3 9 13 2
33 15 9 1 11 11 1 11 11 1 9 1 0 9 1 9 7 9 13 9 1 1 9 1 13 4 9 1 9 1 10 9 13 2
28 11 1 13 16 11 11 1 0 13 4 0 11 11 1 9 1 9 9 0 13 1 9 1 15 9 14 13 2
29 10 9 1 9 1 10 9 13 4 2 15 1 16 10 9 13 4 7 9 9 9 1 15 1 0 9 13 4 2
15 15 13 16 9 1 9 1 9 13 1 9 9 1 13 2
8 10 9 1 15 9 14 13 2
13 10 9 1 12 2 12 9 1 1 0 13 4 2
11 0 9 1 14 9 9 7 9 13 4 2
29 9 9 1 10 9 13 1 1 9 9 9 1 14 9 13 4 2 15 1 14 9 13 1 9 13 4 4 4 2
15 9 1 11 1 0 9 0 13 1 1 14 9 0 13 2
37 15 9 1 10 9 1 0 13 4 16 16 9 15 1 9 13 4 16 15 0 13 4 4 7 16 15 0 9 9 13 4 16 15 9 13 4 2
22 15 13 16 9 7 9 1 9 1 9 1 10 9 13 4 9 1 1 0 14 13 2
28 15 1 9 1 9 13 4 11 11 1 13 16 9 1 13 9 9 1 0 9 1 1 0 9 13 4 4 2
11 15 9 11 11 1 9 1 3 9 13 2
43 11 11 1 11 1 13 4 16 11 1 9 11 2 11 1 9 1 1 0 13 4 1 12 12 1 9 1 9 1 13 9 1 9 1 9 14 13 4 1 9 15 13 2
19 9 1 10 9 1 9 13 1 1 11 1 11 11 1 1 9 13 4 2
21 9 11 11 7 9 11 11 1 9 1 10 9 12 9 9 1 9 13 4 13 2
28 9 1 13 4 4 16 9 11 1 9 9 1 15 1 1 9 1 9 13 4 4 2 7 15 14 13 4 2
19 9 1 9 1 9 13 16 9 1 9 1 11 11 1 9 1 9 13 2
22 9 9 1 11 1 11 11 11 11 2 11 2 1 9 3 13 4 1 9 13 4 2
32 9 1 13 4 16 0 9 9 1 1 11 11 11 1 9 1 9 1 9 1 1 11 11 11 11 11 11 1 9 3 13 2
16 16 11 1 9 9 1 1 1 9 9 1 9 1 9 13 2
47 11 1 0 9 7 11 1 11 1 9 11 11 2 11 11 1 9 11 11 11 7 11 1 9 11 11 11 1 13 16 9 9 7 0 9 1 9 1 1 11 1 9 3 13 4 4 2
32 11 11 11 1 9 1 9 13 4 16 15 0 9 9 13 4 4 9 9 1 1 0 9 1 1 0 9 9 1 9 13 2
33 11 9 11 11 11 1 11 1 15 13 16 15 9 9 9 1 9 1 13 0 11 1 9 1 9 13 1 0 9 1 1 13 2
20 15 13 16 9 1 15 7 0 10 9 1 1 11 11 11 1 9 13 4 2
20 0 13 16 10 9 9 1 9 1 13 1 3 9 9 1 1 13 4 4 2
17 11 1 13 16 0 11 9 1 9 1 9 10 9 1 13 4 2
10 15 13 4 9 1 9 3 0 13 2
27 11 9 11 11 1 13 16 0 11 11 11 1 9 1 1 11 11 9 1 9 1 0 9 13 4 4 2
20 15 13 16 11 1 15 0 9 11 1 9 13 4 15 15 9 13 4 4 2
31 11 1 11 11 11 11 1 9 9 1 1 11 1 13 16 15 9 9 1 0 9 1 1 0 9 1 1 1 13 4 2
22 15 1 12 9 1 11 1 12 12 9 1 9 1 11 11 1 9 13 4 4 4 2
15 11 9 1 10 0 9 9 11 2 11 1 0 13 4 2
12 15 1 12 12 9 1 9 13 1 9 13 2
40 11 1 15 12 0 9 1 9 1 15 13 16 11 11 11 7 11 11 1 9 1 1 9 1 0 9 1 9 13 7 15 1 11 1 11 9 1 9 13 2
20 15 13 16 9 1 11 1 9 13 9 1 9 13 1 1 13 4 4 4 2
21 9 1 9 1 9 0 13 1 11 1 9 13 1 9 1 9 13 4 4 4 2
20 11 1 13 16 9 1 0 9 1 0 9 0 13 1 9 9 13 4 4 2
21 15 13 16 9 1 9 1 1 0 11 11 9 1 14 0 9 0 13 4 4 2
24 9 1 0 9 2 0 9 7 0 9 1 0 9 1 1 11 11 9 1 14 9 0 13 2
33 0 11 9 11 11 11 7 9 9 11 11 1 11 11 1 9 1 1 9 1 9 13 1 1 11 1 11 11 11 1 9 13 2
18 11 9 1 11 11 11 9 1 11 11 11 13 9 1 14 9 13 2
26 9 1 0 9 11 11 11 2 11 11 7 0 9 1 1 11 1 9 1 9 2 9 7 9 13 2
11 11 10 9 1 1 12 9 1 1 13 2
16 12 9 1 0 0 9 1 13 9 1 10 9 13 4 4 2
21 10 9 1 0 9 7 9 9 1 0 9 1 13 0 9 1 11 1 9 13 2
18 11 7 0 9 1 9 13 1 1 14 12 9 9 9 1 0 13 2
24 11 9 1 11 11 11 13 9 1 9 13 2 15 9 1 11 1 9 1 9 1 9 13 2
14 15 1 1 10 9 9 1 9 14 13 4 4 4 2
23 11 1 11 7 11 9 1 13 9 9 1 1 9 9 9 7 9 1 10 9 13 4 2
18 7 11 2 11 7 11 1 10 9 9 9 13 14 13 4 4 4 2
23 11 9 1 9 1 13 16 11 1 10 9 9 1 10 9 1 9 0 13 4 4 4 2
28 11 9 0 2 11 2 9 1 11 1 0 9 1 14 11 11 7 11 11 0 9 2 11 2 13 4 4 2
18 9 1 0 0 9 1 14 10 9 1 13 4 4 1 9 13 4 2
11 11 11 1 9 1 9 13 4 4 4 2
15 11 1 10 9 9 13 9 1 10 9 13 4 4 4 2
19 11 11 9 1 15 12 9 1 1 10 9 1 9 1 9 13 4 4 2
13 11 1 9 1 10 9 1 10 9 13 4 4 2
19 11 11 1 11 2 11 7 11 1 1 10 9 1 9 13 4 4 4 2
13 11 1 0 9 7 9 11 1 14 10 9 13 2
17 11 1 11 1 10 9 1 15 15 9 15 10 9 13 4 4 2
26 11 11 1 11 9 1 12 0 9 1 13 1 12 9 1 9 13 4 2 7 12 9 0 13 4 2
18 11 9 1 11 1 9 9 13 10 9 1 9 1 9 13 4 4 2
12 10 9 12 9 1 14 10 0 13 4 4 2
26 11 11 1 13 9 1 1 2 11 2 0 10 9 1 9 1 15 1 12 9 1 13 4 4 4 2
18 12 0 9 1 1 12 1 0 9 1 1 9 1 9 13 4 4 2
21 9 1 13 11 11 11 1 11 1 0 9 1 9 1 9 1 9 13 4 4 2
48 9 1 9 1 11 1 13 16 15 11 2 11 11 11 11 11 11 2 1 9 1 9 1 0 9 13 1 1 13 4 2 15 14 10 9 1 1 0 9 7 9 1 1 9 13 4 4 2
10 10 9 1 10 9 1 12 9 13 2
25 11 11 1 12 0 9 1 13 16 9 13 1 3 14 9 1 0 9 1 1 1 9 13 4 2
8 11 9 1 13 9 14 13 2
20 15 9 1 13 1 1 9 1 9 13 7 9 1 9 13 1 9 13 4 2
41 9 1 0 9 7 9 1 9 1 13 4 9 1 0 9 13 4 11 11 1 3 10 0 12 9 1 13 4 16 15 10 9 1 13 1 1 15 13 4 4 2
58 9 9 2 11 11 2 1 1 1 0 9 1 9 13 4 9 11 11 11 2 9 11 11 7 9 11 11 11 1 9 1 10 9 1 13 4 16 15 11 11 11 7 11 11 11 1 9 7 9 1 9 1 0 9 1 9 13 2
38 11 11 7 11 11 1 9 1 1 11 11 2 11 2 11 11 2 11 2 11 2 11 7 11 1 9 7 9 1 9 1 9 3 10 13 4 4 2
24 9 1 10 9 1 0 9 1 13 4 16 15 12 9 1 1 10 9 1 0 9 0 13 2
50 11 11 11 9 11 11 11 1 11 1 13 16 0 0 9 1 1 1 0 9 13 1 1 9 1 0 9 1 11 11 11 0 13 1 11 9 1 9 1 15 13 9 1 9 1 9 13 4 4 2
42 11 11 11 1 9 11 11 11 1 15 11 1 9 1 9 1 13 16 9 1 9 1 1 1 9 13 1 15 14 9 1 1 11 11 11 11 1 15 9 13 4 2
45 3 11 9 1 15 0 9 1 0 9 1 0 13 4 9 13 16 11 1 1 1 0 9 1 0 9 13 1 1 3 15 0 9 1 1 1 0 9 1 9 0 14 13 4 2
48 15 13 16 15 10 9 1 9 13 13 4 2 7 9 1 9 1 11 7 11 9 1 9 1 9 13 4 4 7 9 1 13 4 4 16 9 9 1 13 15 14 0 9 14 13 4 4 2
30 0 11 11 11 11 1 9 1 0 10 9 1 9 14 1 11 1 11 11 11 1 9 1 9 1 9 0 13 4 2
32 9 1 0 9 1 0 9 0 11 11 11 11 1 9 13 1 3 12 9 1 9 11 1 0 9 1 1 0 13 4 4 2
24 15 1 9 1 11 1 0 9 11 11 11 7 11 11 1 0 11 11 11 1 9 13 4 2
33 11 9 1 0 9 1 0 9 1 9 9 9 1 0 9 3 0 9 13 4 4 3 9 9 1 9 1 9 13 2 8 4 2
17 9 1 9 10 15 1 9 11 1 0 11 11 11 1 13 4 2
14 15 9 1 9 1 9 9 13 1 3 14 13 4 2
19 9 1 15 11 7 9 1 10 9 1 9 1 9 13 1 9 13 4 2
11 7 11 1 15 1 14 15 9 14 13 2
25 11 9 1 0 9 13 4 11 11 11 1 11 11 11 11 1 13 0 10 9 9 1 0 13 2
13 15 1 14 11 11 11 14 9 1 0 14 13 2
17 11 1 9 11 11 1 9 1 9 1 0 9 1 9 13 4 2
15 0 9 1 9 13 1 14 3 11 11 9 1 13 4 2
28 15 1 9 1 0 11 11 7 0 9 11 11 11 11 1 1 12 0 9 1 9 1 9 1 9 0 13 2
23 9 9 11 11 1 11 1 9 1 9 13 4 15 0 9 2 9 7 9 1 9 13 2
61 0 9 11 11 11 11 1 12 0 9 2 9 11 11 2 11 11 11 11 2 11 11 11 2 11 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 11 11 2 11 11 11 2 11 11 11 1 9 1 14 9 13 4 2
9 9 1 14 11 1 9 13 4 2
39 9 11 11 11 1 11 1 1 9 1 0 9 7 0 9 11 11 2 11 11 11 2 11 11 2 9 11 11 11 7 11 11 11 1 9 1 9 13 2
60 12 9 1 11 2 11 7 11 1 13 0 9 2 11 1 1 11 1 13 9 2 11 11 1 9 9 7 11 1 9 1 0 9 1 10 10 9 1 13 4 7 0 13 9 1 1 9 0 13 4 9 9 7 0 9 1 9 13 4 2
16 0 9 1 9 0 13 1 1 12 9 1 9 14 13 4 2
15 15 1 12 9 1 9 0 9 1 1 0 13 4 4 2
19 15 11 11 11 11 1 9 13 4 4 2 15 15 9 0 13 4 4 2
11 9 9 15 11 11 13 4 1 9 13 2
8 15 9 9 11 15 1 13 2
18 11 9 11 11 1 9 9 9 13 11 1 9 1 1 1 9 13 2
17 11 1 1 15 0 9 11 11 7 9 1 0 9 14 0 13 2
26 11 11 11 1 11 9 9 1 0 9 1 1 9 1 9 13 4 15 15 12 9 0 13 4 4 2
9 15 1 15 9 2 9 1 13 2
10 15 1 11 1 9 9 14 13 4 2
33 0 13 16 10 9 1 9 1 11 1 10 0 9 1 11 1 11 1 9 1 1 1 0 9 1 0 13 4 1 9 13 4 2
16 11 1 9 11 12 11 9 1 9 1 9 1 9 1 13 2
42 11 7 11 1 9 9 1 9 1 9 13 4 9 9 1 9 1 11 11 11 1 15 1 9 13 7 9 9 9 1 1 1 13 4 0 9 1 9 13 1 13 2
27 11 9 11 11 1 9 1 9 1 11 1 13 4 13 16 9 1 10 9 15 9 1 11 1 9 13 2
26 9 9 1 13 16 11 11 11 11 2 11 2 3 9 13 4 4 7 15 0 9 12 12 9 13 2
29 15 13 16 10 9 1 11 11 11 1 0 9 1 9 1 9 13 4 4 15 1 1 0 9 9 0 13 4 2
20 9 1 11 1 11 9 1 1 1 0 9 1 9 9 13 1 9 13 4 2
24 15 13 16 0 0 9 1 0 0 9 1 9 1 13 3 13 4 9 9 1 0 9 13 2
11 15 9 9 1 9 1 9 13 4 4 2
15 16 10 0 9 1 11 1 9 1 1 9 13 4 4 2
32 9 1 13 16 11 1 9 9 1 3 3 13 4 4 4 7 12 0 9 9 1 0 9 1 13 1 9 13 4 4 4 2
27 11 1 11 11 11 1 11 2 11 9 1 11 9 9 1 11 9 1 1 9 9 1 9 1 13 4 2
15 10 9 1 1 10 9 1 9 9 10 9 1 0 13 2
18 0 12 9 1 0 9 9 1 9 1 9 1 9 1 9 13 4 2
25 9 9 1 9 1 13 16 9 1 0 11 2 0 2 1 9 1 9 13 9 9 1 13 4 2
28 10 9 1 1 11 11 2 11 7 11 11 2 11 11 11 1 10 9 1 12 9 1 11 9 1 13 4 2
12 3 1 9 9 1 9 1 3 0 13 4 2
16 9 9 1 0 13 1 1 9 9 1 9 13 4 4 4 2
20 9 1 0 9 1 13 1 1 9 2 3 1 9 1 9 13 4 4 4 2
23 3 11 11 11 1 11 2 11 9 1 0 9 1 11 1 11 9 1 9 13 4 4 2
24 11 1 0 9 1 0 9 1 1 11 1 9 1 11 2 0 9 1 1 9 9 0 13 2
17 10 9 1 15 1 12 1 10 11 2 0 9 13 4 4 4 2
35 11 11 11 11 11 2 11 2 1 12 9 11 11 1 13 16 11 9 1 13 4 4 9 1 11 1 12 1 10 9 13 4 4 4 2
17 0 13 16 11 1 11 1 0 9 1 15 9 0 13 4 4 2
22 11 1 9 1 13 16 0 9 1 11 1 9 1 9 7 9 9 13 4 4 4 2
29 11 1 9 13 16 11 1 0 9 1 12 1 10 0 9 13 4 4 4 2 7 11 11 1 15 9 13 4 2
10 15 14 12 9 1 1 9 0 13 2
27 0 13 16 11 9 1 9 1 0 9 1 0 9 11 1 11 2 0 9 1 1 9 9 9 13 4 2
11 10 9 1 11 1 12 12 9 0 13 2
18 11 1 15 9 13 16 10 9 1 11 1 12 9 0 13 4 4 2
10 0 9 11 9 1 1 13 4 4 2
21 11 1 9 13 16 11 1 9 11 11 11 1 10 0 9 10 9 1 0 13 2
24 16 11 1 15 14 13 13 16 15 0 9 11 1 1 14 15 9 9 9 13 13 4 4 2
14 0 13 16 11 1 9 11 11 2 11 1 13 4 2
9 11 1 11 1 12 9 0 13 2
22 11 1 1 11 1 0 9 1 12 0 0 9 1 9 11 1 0 9 1 0 13 2
11 10 10 9 1 9 11 1 13 4 4 2
22 11 1 11 13 4 1 9 1 11 11 11 9 11 11 12 9 14 0 14 13 4 2
26 11 9 9 3 2 3 14 13 9 9 1 15 13 16 11 1 11 1 0 13 1 15 9 14 13 2
13 16 11 9 1 11 1 0 9 13 1 9 13 2
32 9 1 9 15 13 16 9 9 1 11 11 1 11 11 11 1 9 1 15 15 0 9 1 0 13 16 11 1 11 0 13 2
18 7 9 1 15 9 1 13 10 0 9 1 0 9 0 14 13 4 2
35 11 1 11 9 9 1 9 1 11 1 13 4 16 11 9 1 11 1 14 0 13 4 16 9 1 0 7 0 9 9 1 0 9 13 2
15 7 15 13 16 12 9 1 0 13 1 15 9 14 13 2
13 0 3 10 9 10 9 1 10 9 13 4 4 2
16 7 10 0 9 15 13 2 15 9 13 1 15 9 13 4 2
11 15 1 15 11 1 9 13 4 4 4 2
23 11 1 13 16 9 11 9 1 9 13 7 15 0 13 1 1 0 2 0 9 13 4 2
12 15 0 9 0 0 13 15 0 0 13 4 2
18 15 1 0 10 9 1 1 12 0 9 0 9 9 1 9 13 4 2
21 15 11 11 2 11 2 11 2 11 7 0 0 9 9 1 9 1 0 13 4 2
14 15 13 4 1 16 0 9 1 11 1 10 9 13 2
18 15 9 1 13 16 15 9 14 14 13 15 9 1 1 1 15 13 2
24 11 1 11 1 11 1 11 0 13 1 9 1 1 9 9 13 4 7 15 0 9 13 4 2
11 7 9 1 13 16 15 15 9 14 13 2
20 12 9 1 9 1 11 11 1 13 16 9 11 1 9 13 1 1 0 13 2
19 15 1 11 2 11 7 11 9 1 11 11 11 1 9 13 4 4 4 2
16 15 11 1 9 1 0 9 1 9 13 7 15 9 13 4 2
17 11 11 11 2 11 2 1 11 11 1 0 9 1 9 13 4 2
21 9 9 11 11 1 13 16 11 9 1 11 1 9 13 1 15 15 9 14 13 2
7 16 15 14 13 14 4 2
31 11 1 9 9 1 9 13 1 13 4 9 1 9 1 11 11 11 11 2 11 2 1 11 11 1 9 1 9 13 4 2
25 9 1 13 13 16 11 11 1 15 1 1 3 11 9 1 9 13 9 1 1 15 9 13 4 2
20 11 1 9 1 9 13 1 1 11 1 9 1 11 13 1 14 9 13 4 2
13 15 1 1 9 1 11 1 9 1 14 13 4 2
17 11 1 9 11 11 11 1 11 1 11 11 11 11 1 9 13 2
11 9 1 1 15 11 11 1 12 9 13 2
52 9 1 9 1 11 1 9 9 1 9 13 1 9 1 1 11 9 1 13 1 9 9 1 9 1 9 7 11 1 0 9 1 9 14 13 1 9 1 1 11 1 9 1 9 13 1 14 9 13 4 4 2
21 11 11 1 9 1 1 9 11 11 1 13 16 11 11 1 9 1 15 9 13 2
24 11 11 1 13 16 15 11 11 1 9 13 4 16 9 11 1 1 9 1 1 15 9 13 2
17 15 13 16 15 1 1 11 1 11 1 11 1 9 1 13 4 2
11 7 15 1 15 1 15 9 14 13 4 2
14 11 9 1 0 9 1 0 9 9 1 9 14 13 2
24 15 13 13 16 11 9 1 0 12 9 9 1 9 1 1 11 11 1 11 1 9 13 4 2
29 11 11 11 11 11 11 1 9 1 13 9 1 0 9 7 9 1 0 7 0 9 13 1 9 1 9 13 4 2
22 15 9 7 9 1 0 12 9 1 11 11 11 11 2 11 2 1 0 13 4 4 2
14 9 11 1 2 11 11 2 1 9 1 0 13 4 2
15 11 1 13 13 16 9 1 13 9 1 9 3 13 4 2
13 3 1 9 1 0 7 0 14 9 13 4 4 2
9 9 1 11 1 9 1 13 4 2
28 11 9 11 11 11 1 13 13 16 10 9 7 9 1 9 1 1 0 7 0 9 1 0 9 3 13 4 2
30 11 11 11 1 9 1 13 4 9 1 10 9 1 9 13 4 16 9 9 7 9 1 15 1 9 1 1 9 13 2
30 11 1 0 9 11 11 1 9 1 1 9 1 1 1 9 1 0 9 1 0 9 13 9 1 12 9 0 13 4 2
24 9 1 1 11 1 9 1 0 9 9 1 9 10 9 1 13 7 15 0 9 1 9 13 2
17 9 1 9 1 0 9 1 9 13 7 15 12 9 0 13 4 2
28 11 1 9 11 1 11 11 9 11 11 1 9 1 1 9 1 9 1 9 13 1 1 9 9 1 9 13 2
11 9 9 1 15 14 12 9 0 13 4 2
14 11 1 14 11 9 1 9 1 12 9 0 13 4 2
27 9 1 1 12 9 1 9 1 0 9 10 9 1 9 13 7 9 13 9 1 15 2 15 13 4 4 2
18 9 1 1 9 1 0 9 2 9 7 0 9 1 9 1 9 13 2
26 11 1 9 1 0 9 1 9 1 0 9 13 7 12 2 12 9 1 13 0 9 1 9 14 13 2
27 9 1 12 9 1 12 0 0 9 1 9 1 1 9 1 1 11 11 1 9 1 1 1 9 13 4 2
9 11 11 9 1 9 1 9 13 2
9 9 9 1 11 1 15 9 13 2
21 9 1 1 0 9 1 12 9 1 13 9 1 0 9 1 11 1 1 9 13 2
16 10 9 1 11 1 15 9 1 12 9 1 0 13 4 4 2
31 10 9 1 12 0 9 11 11 7 11 11 1 9 1 9 13 4 13 16 15 10 9 13 15 15 1 11 11 13 4 2
23 0 9 1 9 1 15 9 1 13 4 16 9 13 1 9 1 15 9 11 11 13 4 2
15 11 1 12 0 0 9 1 11 1 9 1 9 13 4 2
19 9 1 11 1 9 1 9 7 9 0 13 0 9 1 1 13 4 4 2
21 11 11 11 1 13 4 16 9 14 0 9 1 9 9 1 9 14 13 4 4 2
40 9 11 11 11 7 11 11 1 11 11 11 11 11 1 9 1 9 9 11 11 11 11 1 9 1 9 13 1 11 11 11 1 9 0 13 4 10 9 13 2
14 9 1 9 1 11 1 12 12 9 13 1 9 13 2
23 9 1 9 1 11 11 11 11 1 15 10 9 1 0 9 13 1 9 1 9 13 4 2
26 7 11 11 2 11 1 9 1 1 1 11 0 11 11 11 1 13 4 12 9 1 9 1 9 13 2
57 7 11 1 12 9 7 12 9 1 12 9 9 1 9 0 9 1 0 9 1 1 13 2 15 9 1 1 9 1 1 1 14 13 4 4 7 9 1 9 1 1 1 9 1 9 9 14 13 4 1 15 1 9 13 4 4 2
38 11 9 9 1 9 1 11 11 7 11 1 9 7 9 1 9 13 1 9 1 0 13 4 11 1 13 4 16 0 9 15 14 9 1 1 0 13 2
18 11 9 1 11 1 11 11 11 1 0 9 1 9 1 9 13 4 2
20 11 1 9 1 0 0 9 1 11 1 9 11 11 1 10 9 1 9 13 2
20 9 1 9 13 16 10 9 1 12 1 12 12 9 9 1 9 1 9 13 2
18 10 9 1 9 1 9 13 1 3 9 1 12 9 9 13 4 4 2
25 11 1 13 16 9 9 7 9 13 1 9 1 0 12 1 12 9 1 12 12 9 10 9 13 2
17 13 4 9 9 1 9 11 2 11 2 11 2 11 13 4 4 2
12 11 9 1 11 1 14 9 1 9 13 4 2
14 11 1 13 9 1 9 1 9 1 12 9 9 13 2
21 15 1 14 9 1 11 11 1 11 11 1 0 9 1 9 1 0 9 13 4 2
12 10 9 1 12 12 9 9 9 1 9 13 2
27 11 1 13 4 4 9 9 1 0 9 1 11 1 12 9 12 9 1 1 12 1 15 15 1 9 13 2
23 11 11 1 0 10 0 9 1 1 9 9 1 1 0 9 1 0 9 14 13 4 4 2
12 11 1 0 9 1 9 11 11 1 13 4 2
20 0 9 1 1 12 9 1 1 13 1 9 1 12 9 15 9 13 4 4 2
25 7 11 1 11 1 1 14 11 9 13 4 7 12 9 1 15 11 9 1 9 13 4 4 4 2
12 11 1 11 9 1 11 11 9 13 4 4 2
17 10 12 9 1 11 1 0 9 1 14 9 1 9 13 4 4 2
16 0 9 1 13 13 16 10 9 1 9 1 11 1 9 13 2
7 16 15 11 0 9 13 2
35 0 9 1 9 1 11 12 1 1 12 9 1 9 13 4 4 7 15 12 9 11 2 12 9 11 7 12 9 11 9 1 1 13 4 2
29 11 1 11 7 11 11 1 0 9 11 11 11 1 9 1 1 0 11 1 1 13 1 9 13 1 9 13 4 2
17 15 1 14 9 1 9 1 10 9 1 9 13 1 9 13 4 2
37 11 11 11 1 9 11 11 11 1 15 12 9 9 1 13 16 11 1 9 9 13 7 9 1 9 9 13 4 1 1 9 1 0 9 14 13 2
38 11 1 13 16 15 10 9 1 9 13 16 10 9 1 9 13 4 16 9 1 10 9 1 9 14 13 2 16 11 11 11 11 1 12 9 14 13 2
23 15 1 14 15 9 1 1 1 13 4 9 1 10 9 1 0 9 0 13 1 9 13 2
17 15 13 16 11 1 9 1 11 1 0 7 0 9 0 13 4 2
48 11 1 9 1 0 7 9 9 13 4 11 1 11 1 0 0 9 11 11 1 11 1 12 9 9 1 13 16 11 1 9 1 14 1 11 1 1 1 9 13 15 9 1 13 4 4 4 2
39 11 9 9 1 9 1 0 9 1 1 11 9 1 9 11 11 11 11 1 9 1 1 1 15 11 7 11 1 9 1 0 9 1 0 13 1 9 13 2
23 15 13 16 11 9 1 11 9 1 9 1 0 13 4 2 15 9 1 9 1 9 13 2
27 11 1 13 16 15 9 1 9 7 11 1 9 1 1 1 11 11 1 11 1 11 9 1 1 9 13 2
11 15 13 16 9 1 15 1 13 4 4 2
31 10 9 1 11 1 13 16 0 9 13 1 11 11 9 1 9 1 15 9 1 9 13 1 9 1 15 9 14 13 4 2
40 11 11 9 9 11 11 1 9 1 1 11 11 1 9 1 1 9 13 1 9 1 15 13 16 11 1 15 1 10 9 1 11 9 1 15 9 14 13 4 2
27 11 1 11 9 1 11 2 11 11 9 1 11 9 9 9 1 12 9 1 12 9 1 9 13 4 4 2
10 9 1 12 9 7 12 9 0 13 2
24 11 1 9 9 11 11 1 13 16 10 9 1 9 13 4 1 9 1 14 12 9 13 4 2
26 15 1 9 2 9 2 11 1 13 4 16 10 9 1 12 9 7 12 9 1 12 9 13 4 4 2
17 11 1 0 9 1 9 1 1 1 13 16 9 1 9 12 13 2
8 15 9 7 9 13 4 4 2
15 9 1 9 1 13 12 9 1 9 13 4 9 13 4 2
16 3 13 4 4 16 10 9 1 9 9 13 4 13 4 4 2
12 15 0 9 9 13 7 0 0 9 13 13 2
17 9 1 9 7 9 1 9 1 1 1 15 9 14 13 4 4 2
15 3 14 9 9 1 9 1 10 9 1 9 13 4 4 2
43 11 11 1 16 11 1 9 1 0 11 11 11 1 12 9 9 1 13 1 9 13 4 2 7 11 7 11 1 9 1 11 11 1 9 1 1 0 9 0 13 4 4 2
35 11 11 11 11 11 11 9 11 11 1 13 16 11 11 11 11 11 1 0 9 1 1 11 2 11 1 10 0 9 1 0 9 13 4 2
20 15 1 11 7 11 1 9 1 12 0 9 1 0 9 9 13 4 4 4 2
26 11 11 11 1 9 1 11 11 11 1 9 1 11 1 9 7 9 1 13 4 4 9 1 9 13 2
26 15 13 16 11 7 11 1 9 1 9 0 13 4 4 7 10 9 11 1 13 1 9 13 4 4 2
26 11 9 16 15 0 9 0 9 1 0 7 0 13 4 4 2 15 11 1 9 1 13 13 4 4 2
20 12 9 11 2 11 2 11 11 2 11 2 11 7 11 1 10 9 0 13 2
17 10 9 1 11 1 13 1 0 9 11 1 1 1 13 4 4 2
22 15 1 0 11 11 11 1 1 0 9 1 9 1 0 9 9 9 13 4 4 4 2
54 9 1 1 0 9 1 12 0 9 11 2 11 2 11 2 11 11 2 11 2 11 2 11 7 11 11 1 14 10 9 1 9 9 13 4 16 11 2 11 1 9 1 9 1 13 9 1 9 9 0 13 4 4 2
25 11 1 13 16 11 11 11 11 11 1 0 9 1 1 9 1 9 1 12 12 9 0 13 4 2
6 0 9 11 1 13 2
15 11 11 1 9 1 9 1 0 9 1 9 13 4 4 2
11 9 1 10 9 1 0 9 3 13 4 2
19 15 13 16 9 11 9 1 0 9 1 9 9 0 13 1 0 9 13 2
29 11 11 1 11 1 1 13 1 11 11 11 11 1 9 1 9 11 9 1 1 9 1 9 1 13 1 13 4 2
19 15 9 9 1 0 13 4 7 3 13 4 4 2 7 9 3 13 4 2
11 9 1 9 2 9 1 15 9 14 13 2
14 9 1 0 9 1 10 9 1 9 13 4 4 4 2
10 15 9 1 9 13 1 9 13 4 2
31 11 11 1 14 11 13 11 1 13 1 11 11 11 11 11 11 1 15 0 9 1 12 9 9 1 9 12 9 0 13 2
12 11 1 13 1 3 15 0 9 11 9 13 2
9 11 1 13 9 3 11 13 4 2
18 9 1 0 11 9 9 1 9 12 13 4 12 9 1 9 13 4 2
11 14 12 12 9 9 11 9 1 1 13 2
19 10 3 9 1 9 1 13 1 9 13 4 7 9 13 4 3 13 4 2
15 9 1 9 14 12 9 1 1 14 9 1 13 4 4 2
16 16 10 9 1 14 10 9 1 9 9 9 1 13 4 4 2
11 15 1 15 9 1 9 0 13 4 4 2
14 3 1 11 9 1 14 12 9 1 9 1 13 4 2
11 11 9 1 10 9 14 12 12 9 13 2
9 15 1 15 9 1 9 13 4 2
16 9 1 15 1 9 12 13 4 12 9 1 0 13 4 4 2
14 11 1 3 0 9 1 11 0 11 11 14 13 4 2
16 9 1 0 9 1 11 7 11 9 1 0 9 1 9 13 2
15 10 3 0 9 1 12 9 9 1 1 14 0 13 4 2
33 9 9 11 11 1 13 16 9 1 10 9 1 9 14 14 0 13 2 7 10 0 9 1 10 9 1 0 9 1 13 4 4 2
12 15 0 9 1 10 9 1 9 13 4 4 2
10 9 1 9 0 9 9 1 13 4 2
38 11 2 11 1 0 9 11 11 11 11 1 11 1 0 2 0 13 16 0 11 11 11 1 9 1 1 15 9 1 9 1 15 9 14 14 0 13 2
12 11 0 11 11 11 1 9 13 9 13 4 2
18 11 1 13 16 15 9 1 0 11 2 11 2 11 14 0 9 13 2
20 15 10 9 1 15 9 1 9 14 14 13 15 9 1 9 1 9 13 4 2
12 9 1 15 13 1 15 15 0 13 4 4 2
31 10 9 1 11 9 1 9 13 4 2 15 10 9 1 15 9 14 13 7 15 0 9 1 9 13 1 9 13 4 4 2
38 15 13 16 9 11 1 11 11 9 1 9 1 9 1 1 15 9 13 7 15 1 11 11 1 9 1 0 13 9 1 9 7 15 9 1 1 13 2
19 15 13 16 11 1 0 9 1 15 9 10 9 1 0 13 1 0 13 2
38 11 1 12 9 1 13 1 11 1 11 11 11 1 9 1 1 11 1 13 16 10 9 1 11 1 12 9 1 13 9 1 9 1 9 13 4 4 2
22 15 10 9 14 9 1 1 13 2 7 10 9 1 9 1 1 14 15 3 13 4 2
19 12 9 1 9 1 15 13 16 11 11 1 11 11 11 1 9 13 4 2
20 9 1 10 0 9 13 4 15 0 9 1 13 4 4 16 15 15 13 4 2
19 0 9 1 11 2 11 9 1 0 9 1 0 9 1 9 13 4 4 2
22 15 13 16 11 11 11 1 10 9 1 9 13 4 16 15 11 1 15 9 13 4 2
19 11 1 10 9 1 9 13 4 16 11 0 9 1 3 0 9 13 4 2
37 16 2 0 9 1 1 1 11 1 10 9 1 11 1 10 9 1 9 13 2 15 1 15 9 1 0 9 1 9 13 1 0 9 13 4 4 2
32 11 1 9 1 9 1 0 9 0 11 9 1 12 9 1 9 13 4 4 7 0 9 1 0 9 1 9 14 13 4 4 2
25 9 1 0 13 4 9 9 1 9 1 13 4 1 1 11 1 11 1 9 9 1 9 13 4 2
23 11 11 11 11 11 1 11 11 11 11 2 11 2 1 9 1 10 9 9 1 9 13 2
27 11 11 11 11 1 11 11 11 2 11 2 1 9 1 1 10 9 1 9 1 1 11 11 1 13 4 2
32 10 9 1 1 9 9 13 1 9 1 13 10 9 13 4 4 4 2 15 11 2 11 7 11 1 13 9 13 4 4 4 2
22 9 1 1 2 11 1 9 1 9 13 11 11 11 1 1 11 1 0 13 4 4 2
15 15 10 9 9 1 13 9 1 15 0 13 4 4 4 2
30 13 4 16 11 9 1 11 11 11 1 9 1 11 1 9 13 4 11 11 11 11 1 0 12 9 1 9 13 4 2
25 15 1 9 14 1 9 1 11 11 11 11 1 11 1 11 11 11 13 4 1 9 13 4 4 2
23 9 1 13 13 16 11 1 10 9 9 1 13 1 1 9 13 1 9 9 13 4 4 2
29 11 11 11 11 1 9 1 13 13 16 10 9 1 11 11 11 1 9 1 9 1 9 10 9 1 13 13 4 2
22 15 9 1 11 1 0 12 9 1 9 13 4 2 15 11 2 11 7 11 0 13 2
26 9 1 14 12 9 1 1 11 11 11 1 9 1 11 1 10 9 9 1 13 1 9 13 4 4 2
36 15 13 16 15 3 10 9 9 1 13 1 1 10 9 13 2 7 11 1 1 1 11 11 11 1 13 4 1 1 9 0 13 4 4 4 2
30 11 11 11 11 11 11 2 11 2 1 12 9 0 13 4 2 15 9 9 9 11 11 11 11 1 9 9 1 13 2
9 3 1 9 11 11 11 14 13 2
6 15 9 10 15 13 2
17 11 11 1 10 9 1 9 1 13 9 1 9 1 9 9 13 2
15 15 13 16 15 9 9 13 4 4 4 15 9 0 13 2
14 3 11 1 11 2 11 2 11 11 1 9 0 13 2
12 9 9 13 16 10 9 1 15 15 14 13 2
9 11 11 1 9 1 1 9 13 2
5 9 15 14 13 2
15 0 9 1 9 13 15 9 13 10 9 1 0 13 4 2
5 9 1 15 13 2
13 11 11 11 1 10 9 1 14 9 1 9 13 2
10 11 7 11 1 9 15 15 1 13 2
11 9 1 1 1 9 1 10 9 13 4 2
14 15 11 1 13 9 1 9 13 1 9 14 13 4 2
24 11 11 1 11 11 1 12 9 1 12 9 1 12 9 13 7 9 15 12 9 9 13 4 2
14 10 9 1 9 1 10 9 9 1 9 1 9 13 2
7 12 9 1 10 13 4 2
10 9 1 9 13 1 1 15 9 13 2
19 11 11 1 11 11 1 13 11 1 9 1 11 9 1 9 13 4 4 2
13 11 13 16 3 9 0 13 4 4 7 14 13 2
8 9 1 15 9 15 14 13 2
10 11 1 14 9 1 11 11 13 4 2
8 9 1 15 9 15 14 13 2
13 10 9 1 14 0 9 1 9 1 9 13 4 2
4 15 9 1 13
12 11 1 12 9 9 9 2 11 11 2 13 2
10 16 3 9 1 9 1 15 13 4 2
9 9 9 1 9 3 12 9 13 2
7 9 1 15 9 1 13 2
18 11 1 11 2 11 11 1 13 1 1 9 1 15 9 1 9 13 2
20 15 15 0 14 13 16 10 9 1 12 9 1 9 1 0 9 13 4 4 2
33 15 13 1 16 0 9 1 10 9 1 15 3 14 15 1 13 1 9 13 4 2 15 15 11 11 1 11 1 9 1 0 13 2
8 11 9 1 13 2 3 13 2
10 15 15 9 13 16 9 1 15 13 2
7 9 1 15 13 2 9 2
16 11 11 2 11 11 7 11 9 11 11 1 1 10 9 13 2
13 10 9 1 9 1 1 9 13 4 9 9 13 2
10 3 9 9 9 1 9 13 4 4 2
23 9 1 0 7 0 9 1 9 15 9 7 9 1 9 1 1 9 1 0 13 4 4 2
20 9 1 9 1 13 4 9 1 10 9 1 9 13 1 9 1 9 13 4 2
17 15 13 13 16 0 3 15 0 9 1 0 9 1 9 13 4 2
24 11 9 1 0 9 2 11 1 1 0 9 9 1 9 7 15 9 9 14 9 13 4 4 2
20 16 10 9 1 9 10 9 14 13 16 10 0 9 1 9 14 13 4 4 2
21 11 9 1 9 1 13 4 4 16 9 1 9 1 9 1 9 0 9 1 13 2
13 0 9 9 9 1 1 10 12 9 0 13 4 2
25 11 9 1 9 1 13 13 16 15 14 13 16 9 1 9 0 13 1 9 1 0 13 4 4 2
6 9 10 14 0 13 2
37 11 11 11 11 11 11 11 1 9 9 11 11 1 13 13 16 15 9 1 9 9 1 13 4 4 2 15 9 1 1 0 9 1 9 13 4 2
15 15 13 16 10 9 1 9 1 9 13 4 1 9 13 2
26 11 11 11 11 1 9 9 1 9 11 11 1 13 13 16 0 9 0 7 0 9 1 13 4 4 2
28 15 13 16 0 9 2 15 9 1 9 1 1 1 13 4 4 2 1 0 9 1 9 1 0 13 4 4 2
26 15 13 16 9 1 0 9 1 9 1 9 7 15 1 13 4 9 1 9 14 9 1 13 4 4 2
8 0 9 13 4 13 4 4 2
21 0 9 11 11 11 1 13 13 16 0 9 1 9 1 9 13 4 1 9 13 2
29 15 13 16 9 1 9 1 0 9 1 0 9 1 9 1 9 0 13 1 9 13 2 7 9 1 15 14 13 2
16 9 1 9 1 0 0 9 11 11 1 9 10 13 4 4 2
12 11 15 9 1 9 9 2 12 13 4 4 2
21 11 1 11 11 9 1 3 0 9 13 2 7 11 1 11 11 0 9 1 13 2
27 11 11 1 9 1 12 9 1 9 0 13 4 2 15 11 12 12 9 1 9 1 1 0 9 1 13 2
17 9 1 0 9 11 7 11 11 1 9 12 12 9 13 4 4 2
16 3 9 9 11 11 12 12 1 9 1 1 0 9 1 13 2
22 9 1 0 9 1 13 4 11 1 0 9 11 11 12 12 9 1 9 1 9 13 2
14 11 11 12 12 9 1 9 1 1 0 9 1 13 2
16 10 0 9 1 12 9 3 0 9 1 9 0 13 4 4 2
13 11 11 1 11 1 3 0 9 0 13 4 4 2
22 11 9 11 7 11 1 12 12 9 1 9 1 1 11 1 9 1 0 9 13 4 2
22 11 11 11 1 9 11 11 12 12 9 1 9 1 1 11 1 1 0 9 1 13 2
38 0 9 9 11 11 12 12 9 1 9 1 1 11 1 9 1 0 9 1 13 2 7 11 1 9 11 11 1 10 9 1 12 9 1 13 4 4 2
116 11 1 9 1 9 1 0 0 9 1 11 11 2 9 9 2 12 12 9 2 2 11 11 2 9 2 12 12 9 2 2 11 9 2 9 9 2 12 12 9 2 2 11 11 2 9 2 12 12 9 2 2 11 11 2 9 9 2 12 12 9 2 2 11 11 2 9 9 2 12 12 9 2 2 11 7 11 11 2 9 2 12 12 9 2 2 9 11 7 9 2 12 12 9 2 2 11 11 11 2 12 12 9 2 7 9 11 11 2 12 12 9 2 0 13 2
18 0 9 15 13 16 0 9 10 9 1 12 9 1 14 13 4 4 2
24 15 13 11 9 1 11 11 2 15 12 12 9 1 9 1 1 10 9 1 0 9 1 13 2
26 0 9 14 12 0 9 1 9 13 4 16 11 1 9 9 1 9 1 12 9 1 12 12 9 13 2
15 12 0 11 9 1 0 9 13 4 1 3 1 0 13 2
17 9 9 1 9 1 9 1 9 1 0 9 1 9 3 9 13 2
21 9 1 9 9 9 1 9 1 12 9 14 9 1 9 1 9 0 13 4 4 2
19 10 9 11 9 1 9 9 9 1 9 1 15 9 1 9 14 13 4 2
15 0 9 1 11 1 13 9 1 10 0 0 9 13 4 2
42 15 11 11 11 11 11 11 1 9 1 9 2 11 2 1 3 13 7 11 1 11 11 9 9 1 9 13 4 0 0 9 1 9 1 12 9 13 1 9 0 13 2
16 11 1 9 11 1 13 10 9 1 12 9 1 9 13 4 2
29 7 9 1 15 14 13 16 9 1 0 9 1 13 9 1 1 15 13 4 16 9 1 9 1 14 9 13 4 2
23 9 9 9 1 9 11 11 11 1 13 16 10 9 15 2 9 9 2 9 1 14 13 2
42 0 9 1 0 0 9 1 9 1 1 11 11 11 11 1 9 1 0 13 4 13 16 9 1 9 9 1 9 1 12 9 1 0 9 1 0 13 1 9 13 4 2
23 7 15 0 13 4 16 15 1 9 9 1 9 1 1 1 13 4 10 9 3 13 4 2
31 15 13 4 1 16 9 9 1 9 1 12 9 1 0 9 1 0 15 13 4 2 11 1 15 14 13 1 9 13 4 2
30 0 13 16 9 9 9 1 9 1 12 9 1 0 9 1 13 1 9 11 1 9 9 1 9 1 1 13 4 4 2
29 11 11 11 1 9 1 9 1 12 9 14 9 7 9 1 9 1 12 9 14 9 1 9 1 9 13 4 4 2
40 0 9 1 0 9 1 9 1 9 13 1 11 11 1 9 1 9 1 12 9 14 9 1 9 1 9 13 7 9 1 9 1 15 9 1 9 14 13 4 2
16 9 9 9 1 9 1 14 15 9 1 9 14 13 4 4 2
24 3 9 1 11 11 11 11 11 11 1 9 1 9 2 11 2 1 3 13 1 9 13 4 2
41 9 1 9 1 1 11 11 11 11 11 11 11 1 13 16 15 9 1 9 1 9 1 1 9 7 0 9 14 9 9 1 1 9 9 13 1 9 13 4 4 2
8 7 15 0 9 0 14 13 2
23 9 1 11 9 9 1 9 13 4 0 0 9 1 9 1 12 9 13 1 9 13 4 2
23 9 1 11 11 11 1 9 9 1 9 11 11 11 1 1 13 1 9 1 9 13 4 2
33 15 1 9 1 11 11 11 1 0 9 13 7 10 9 1 9 1 9 1 1 9 1 9 13 1 12 9 1 0 9 13 4 2
21 11 11 1 11 1 9 7 9 1 9 11 11 1 9 12 9 1 1 13 4 2
14 9 1 10 9 11 1 9 1 0 9 1 13 4 2
17 9 1 11 1 9 9 1 9 0 13 4 1 9 13 4 4 2
18 0 13 16 11 1 11 1 11 1 11 11 11 1 9 13 4 4 2
20 11 1 9 7 10 0 9 1 11 1 9 1 9 0 13 1 9 13 4 2
12 11 1 10 9 1 11 11 1 9 13 4 2
47 9 1 9 11 11 7 11 11 11 1 0 9 11 11 11 1 9 1 13 16 9 11 11 7 9 11 11 1 0 9 1 9 1 0 9 1 1 11 9 12 9 1 9 0 13 4 2
14 11 1 9 1 9 1 9 13 1 1 9 13 4 2
17 15 9 1 13 4 11 11 1 9 12 9 1 1 13 4 4 2
20 10 9 1 11 1 9 11 11 7 11 11 1 11 11 1 9 0 13 4 2
24 9 1 11 11 1 11 1 11 1 9 9 1 9 1 0 13 1 9 1 9 13 4 4 2
17 9 1 13 4 16 11 1 14 9 1 9 1 9 1 13 4 2
10 15 9 1 0 9 1 9 14 13 2
19 15 1 14 9 9 1 9 1 0 13 1 0 9 1 9 14 13 4 2
25 15 1 9 1 9 1 1 1 11 1 9 1 9 1 0 12 9 1 0 14 13 4 4 4 2
25 15 1 2 11 11 1 11 11 1 11 1 9 1 9 13 1 11 11 1 9 1 0 13 4 2
34 0 13 16 11 11 11 2 11 1 11 1 11 9 1 12 9 1 9 12 1 0 9 11 11 1 9 1 1 15 9 13 4 4 2
12 11 1 11 11 1 10 9 1 9 13 4 2
24 10 9 1 13 4 11 11 1 11 1 9 1 9 1 0 9 1 13 4 1 9 13 4 2
20 11 9 11 11 1 0 9 13 1 9 11 11 1 9 9 1 9 13 4 2
31 9 14 13 9 1 1 9 1 15 9 0 13 4 4 7 11 9 1 1 1 15 9 1 9 1 0 15 14 13 4 2
25 7 2 15 0 13 16 11 9 11 11 1 9 11 1 12 9 1 9 9 1 13 4 4 4 2
8 3 11 11 15 11 1 13 2
23 11 1 11 11 1 9 1 9 1 13 4 2 9 2 1 9 14 13 1 9 13 4 2
21 11 1 13 16 11 9 9 1 1 9 1 0 9 1 15 9 1 9 13 4 2
10 11 1 13 16 15 9 1 9 13 2
14 7 11 9 11 11 1 15 11 1 0 9 9 13 2
16 3 11 11 1 0 9 11 1 15 14 13 1 9 13 4 2
19 11 1 0 9 11 11 1 9 9 1 11 1 9 0 13 1 9 13 2
24 15 13 4 1 16 11 11 1 9 1 10 9 13 4 2 11 1 13 16 15 9 11 13 2
14 3 11 11 1 9 1 0 9 14 0 13 4 4 2
16 11 1 1 9 2 9 13 1 11 11 10 9 11 1 13 2
18 15 11 1 0 9 11 11 1 9 1 11 1 0 9 1 0 13 2
7 15 15 15 1 9 14 13
24 11 11 1 9 1 0 13 1 9 11 7 11 1 0 9 1 1 9 9 1 13 4 4 2
23 10 9 1 9 9 11 11 2 11 11 7 11 11 1 1 11 11 7 11 11 0 13 2
27 11 11 1 0 11 11 11 1 11 11 1 9 1 1 0 9 1 9 1 11 9 11 1 9 13 4 2
28 11 1 11 11 2 11 11 2 11 11 7 11 11 11 1 0 9 1 9 1 1 9 1 9 13 4 4 2
17 15 14 1 11 1 11 1 9 9 9 1 13 0 13 4 4 2
23 9 9 1 13 13 16 11 1 9 1 9 0 9 9 1 9 9 1 1 1 13 4 2
16 11 11 1 9 9 1 11 1 9 1 9 1 9 13 4 2
40 9 9 1 11 11 1 9 0 13 4 1 9 1 1 0 11 11 1 9 11 11 11 1 13 16 11 1 1 11 1 9 1 12 0 9 1 0 9 13 2
13 11 11 1 0 9 14 11 1 9 13 4 4 2
12 7 11 9 11 11 11 1 15 9 13 4 2
24 12 9 1 9 1 11 1 13 4 16 11 11 1 11 1 9 9 1 15 14 13 4 4 2
26 0 9 1 9 1 9 1 9 1 10 9 7 10 9 1 13 1 1 9 1 14 9 0 13 4 2
16 15 1 11 11 11 11 1 9 1 9 1 9 13 4 4 2
20 11 11 1 9 9 13 1 12 9 1 9 1 9 9 1 9 0 13 4 2
14 10 9 1 9 1 10 9 1 9 1 0 13 4 2
24 11 11 11 11 1 9 1 9 9 1 9 1 9 1 9 1 1 11 1 9 1 9 13 2
9 9 1 9 1 0 9 13 4 2
29 0 9 1 1 11 2 11 2 11 7 11 1 10 10 9 1 9 13 4 2 15 11 9 1 13 1 13 4 2
13 9 1 9 9 1 13 1 9 11 11 1 13 2
10 9 13 16 10 9 1 9 11 13 2
24 15 1 10 10 9 1 14 9 13 4 2 15 1 9 1 9 1 9 1 0 13 4 4 2
16 15 11 11 2 11 2 11 2 11 2 11 7 11 0 13 2
28 11 1 9 1 9 9 1 9 1 9 10 9 3 13 4 15 11 9 11 11 11 1 0 9 13 4 4 2
17 10 9 1 9 13 16 9 9 1 1 15 9 14 13 4 4 2
27 9 1 13 13 16 11 9 1 13 9 1 15 15 9 14 13 4 16 10 9 1 9 0 2 0 13 2
28 11 1 11 1 12 9 7 9 9 13 1 9 13 2 16 11 1 11 1 11 9 1 9 13 1 9 13 2
9 9 1 0 9 15 0 14 13 2
27 11 11 1 10 9 2 9 1 9 0 13 2 15 9 1 9 9 1 9 1 11 11 1 11 13 4 2
23 15 11 1 9 14 1 9 13 7 11 11 1 11 1 13 1 11 1 9 1 0 13 2
26 9 9 11 11 13 4 16 10 14 9 15 14 13 16 0 11 11 1 10 9 1 14 9 0 13 2
16 15 13 1 9 9 1 9 1 9 1 9 1 13 4 4 2
28 11 1 0 9 1 9 13 1 0 11 2 11 9 11 11 11 1 0 9 9 11 1 14 9 1 9 13 2
23 0 9 9 1 13 4 16 11 1 11 1 11 2 11 1 9 9 13 1 9 13 4 2
16 9 1 1 12 0 11 1 9 2 9 11 1 13 4 4 2
15 0 9 1 15 2 11 11 2 1 9 13 4 4 4 2
17 13 4 4 4 16 11 1 13 0 9 1 1 15 1 9 13 2
21 10 9 1 14 15 1 9 0 13 4 16 11 1 11 1 0 13 4 4 4 2
48 11 1 2 11 11 2 1 11 1 1 1 13 16 11 11 1 11 1 13 9 1 1 11 1 14 9 13 2 7 0 0 0 9 9 1 9 1 11 1 0 13 1 9 1 9 13 4 2
13 9 1 1 11 11 1 12 0 9 1 9 13 2
16 11 9 1 1 11 0 9 11 1 9 1 9 1 13 4 2
10 15 15 11 11 1 1 11 13 4 2
10 11 11 2 0 9 2 1 9 13 2
12 15 15 11 11 11 1 0 9 13 4 4 2
32 9 9 9 1 9 13 4 16 10 9 11 11 1 13 4 2 15 11 1 11 1 11 1 1 9 9 13 1 9 13 4 2
11 9 1 1 12 9 9 9 13 4 4 2
15 10 9 11 1 12 9 1 9 11 11 1 9 1 13 2
12 11 1 10 9 3 14 0 0 13 4 4 2
31 10 9 1 0 9 1 13 13 16 11 11 11 13 1 11 1 15 13 10 9 13 16 11 1 1 9 1 9 14 13 2
7 9 1 14 9 14 13 2
9 15 1 9 1 9 13 4 4 2
29 9 1 9 13 12 9 11 7 11 15 1 13 4 2 7 9 1 9 1 9 1 12 9 1 1 15 13 4 2
8 7 10 9 1 13 14 4 2
15 11 11 11 1 11 1 11 2 11 1 9 1 9 13 2
23 11 1 13 16 9 1 9 1 9 11 2 11 1 9 7 9 1 9 13 4 4 4 2
24 9 1 9 11 1 1 1 9 0 13 1 14 9 1 12 0 9 15 9 13 1 0 13 2
16 10 9 9 11 11 7 11 11 1 1 13 9 1 0 13 2
26 11 1 9 13 4 9 9 1 11 1 9 1 13 4 0 9 1 1 12 9 1 9 14 13 4 2
24 11 1 9 13 1 0 9 1 9 1 9 13 7 0 9 1 9 1 9 0 9 1 13 2
17 15 13 13 16 9 1 0 9 1 9 9 9 1 13 4 4 2
21 11 1 11 2 11 1 9 1 9 1 9 1 9 1 9 13 1 9 13 4 2
22 15 1 11 1 11 11 11 1 0 0 9 13 10 9 1 9 1 13 1 13 4 2
27 9 1 9 13 1 12 0 9 1 2 11 11 2 1 13 16 11 7 11 11 1 9 14 12 1 13 2
12 11 11 1 9 11 11 1 9 1 9 13 2
23 7 11 13 4 16 9 11 11 7 11 11 1 1 13 9 1 0 9 1 0 13 4 2
25 15 1 9 2 9 9 7 9 11 11 1 1 13 7 0 0 9 9 1 9 1 13 4 4 2
19 16 2 11 11 7 11 11 1 11 7 11 11 1 9 1 9 13 4 2
35 11 11 1 9 9 13 1 3 14 11 11 11 1 9 13 15 0 13 4 4 16 11 7 11 1 1 9 1 9 11 2 11 14 13 2
20 9 1 9 1 13 13 16 15 9 1 0 9 1 9 1 14 0 14 13 2
35 11 11 1 0 9 1 13 10 9 9 1 9 10 9 13 1 3 0 13 4 16 15 9 1 14 14 9 1 9 9 13 4 4 4 2
23 16 2 11 1 9 13 16 9 1 0 9 1 13 11 11 14 10 9 1 0 13 4 2
21 9 1 11 2 11 1 1 11 7 11 1 9 13 1 0 9 1 14 9 13 2
33 11 11 1 9 13 4 11 11 11 1 13 16 15 11 1 9 1 0 9 1 9 0 13 1 0 13 16 10 9 0 13 4 2
22 15 0 11 1 9 1 10 9 1 9 13 1 9 13 4 9 1 9 1 9 13 2
18 15 11 11 1 9 1 2 10 15 1 13 1 9 12 1 14 13 2
24 11 1 9 1 1 1 11 7 11 1 9 1 9 11 1 13 1 9 1 0 13 4 4 2
32 10 9 11 1 13 4 15 13 1 9 11 1 13 1 9 1 0 13 4 4 7 15 9 1 9 13 15 9 1 9 13 4
20 16 2 9 1 9 1 0 0 9 1 0 9 1 9 14 0 13 4 4 2
12 0 9 11 9 1 11 1 13 1 9 13 2
24 11 11 1 11 11 1 9 1 9 13 4 13 4 16 11 9 0 9 1 9 1 13 4 2
8 15 15 9 14 13 4 4 2
26 9 11 11 7 9 11 11 11 1 15 9 1 13 16 9 1 0 9 0 13 1 9 14 14 13 2
33 16 9 1 0 13 4 16 11 11 11 11 2 11 2 1 13 4 16 9 9 1 9 10 9 1 0 9 1 1 1 13 4 2
32 9 1 11 1 9 1 9 1 13 16 10 9 1 9 1 9 7 9 1 0 0 10 9 9 1 1 15 1 14 13 4 2
17 15 14 0 13 4 16 11 9 9 2 9 9 1 0 9 13 2
41 11 2 11 9 1 15 0 9 1 0 13 4 11 12 0 9 9 1 9 1 1 11 1 1 9 7 9 9 1 0 9 13 1 9 2 11 2 1 9 13 2
21 11 1 13 13 16 15 1 12 9 1 1 9 1 9 1 3 13 1 9 13 2
30 0 9 11 1 11 2 11 9 1 9 1 9 0 13 1 3 0 9 12 9 10 0 9 1 9 13 1 0 13 2
76 9 1 1 11 1 1 1 9 1 14 13 4 7 15 1 10 9 1 9 1 0 13 4 1 9 13 15 11 7 11 1 11 11 3 14 13 2 11 7 11 0 9 1 9 1 9 13 4 12 13 2 11 1 11 1 1 9 9 9 13 7 12 9 1 9 1 9 9 1 1 11 9 14 0 13 2
23 9 1 11 9 1 0 13 4 1 1 1 11 1 9 1 13 9 9 11 1 13 4 2
19 11 1 9 13 1 3 12 9 1 1 0 0 0 9 13 4 4 4 2
44 11 11 11 1 9 1 9 9 1 0 9 1 1 11 1 10 0 9 1 9 1 1 9 1 0 13 1 9 1 1 11 11 1 9 13 4 4 9 1 0 9 13 4 2
10 9 1 11 1 9 9 9 11 13 2
20 10 9 1 0 9 9 11 11 7 11 11 1 0 0 9 11 1 9 13 2
25 11 11 1 9 11 11 1 13 16 9 1 0 9 1 9 15 1 9 9 11 11 13 4 4 2
22 11 9 1 11 11 1 11 11 9 1 9 11 11 11 1 0 13 4 1 9 13 2
29 9 1 13 13 16 15 1 12 9 1 1 9 9 1 13 9 1 9 1 12 9 9 1 9 1 0 9 13 2
35 12 9 1 1 9 9 13 1 9 0 11 9 1 11 1 13 11 11 1 1 0 11 11 7 11 1 0 9 11 11 11 1 13 4 2
32 11 1 11 1 9 11 11 11 1 12 9 1 0 9 1 13 16 11 1 11 9 1 9 1 13 10 9 1 10 9 13 2
19 12 9 9 11 1 12 9 1 11 11 1 13 4 9 1 14 9 13 2
27 11 11 11 11 11 1 13 4 16 9 1 1 13 4 9 1 13 1 1 0 0 9 1 9 13 4 2
13 9 1 9 1 1 9 1 9 1 9 13 4 2
17 9 1 9 1 13 1 1 3 14 11 1 9 1 9 13 4 2
21 11 1 0 9 1 1 9 9 1 15 9 9 9 13 1 0 9 13 4 4 2
17 15 13 16 11 1 11 1 1 1 0 13 1 9 13 4 4 2
17 15 1 9 9 13 1 11 2 11 7 11 11 0 13 4 4 2
13 11 11 1 11 1 1 9 9 13 1 9 13 2
14 11 1 9 1 9 9 13 1 14 9 13 4 4 2
31 9 9 1 9 1 9 1 0 13 4 11 1 13 16 9 2 9 9 1 13 0 0 9 0 9 9 1 9 14 13 2
16 15 13 16 9 9 9 1 9 1 0 9 1 13 4 4 2
10 15 3 14 15 9 9 1 13 4 2
11 10 9 9 1 0 9 1 0 13 4 2
58 3 1 9 1 9 1 11 1 13 16 9 1 0 9 9 9 13 2 0 9 9 1 9 9 13 7 9 1 9 2 9 7 9 1 9 1 1 0 7 0 9 9 9 1 1 9 1 9 7 9 7 9 1 9 1 9 13 2
20 11 11 11 1 9 1 15 13 16 15 1 12 9 1 9 1 9 13 4 2
11 10 9 1 11 9 1 9 1 0 13 2
16 11 2 11 9 9 1 9 1 11 11 1 9 13 4 4 2
15 12 9 1 10 9 1 9 1 9 13 1 9 13 4 2
29 15 13 16 9 7 9 1 1 13 9 1 13 1 9 1 11 1 11 7 11 11 1 12 0 9 13 4 4 2
22 11 11 1 13 16 11 11 1 0 9 1 0 13 1 10 9 9 9 1 13 4 2
21 11 7 11 9 9 1 1 11 2 11 9 1 12 9 11 9 9 1 13 4 2
17 9 1 9 1 13 16 9 9 9 12 9 11 1 0 13 4 2
11 7 11 13 1 3 14 10 9 13 4 2
10 9 1 9 1 9 13 4 4 4 2
26 11 0 9 1 9 1 10 9 9 13 4 11 1 0 9 7 15 9 1 9 13 4 9 13 4 2
33 11 1 9 11 11 11 7 15 9 11 11 1 1 0 13 4 0 12 0 9 1 9 1 11 1 9 1 14 0 13 4 4 2
31 16 15 14 0 9 1 10 0 9 1 9 14 13 4 2 7 9 1 9 13 16 15 11 2 11 2 11 1 9 13 2
41 11 1 9 9 11 11 7 15 9 11 1 9 11 1 9 11 9 1 14 12 9 1 11 1 1 13 11 9 1 0 9 1 12 9 1 1 13 9 1 13 2
10 10 9 11 7 11 9 1 1 13 2
17 9 1 9 0 9 1 9 12 9 1 1 13 7 9 1 13 2
20 9 1 0 9 1 9 12 9 1 1 12 9 1 9 0 13 1 9 13 2
14 12 9 1 9 1 0 9 1 1 9 1 9 13 2
10 15 9 15 9 1 9 13 13 4 2
12 12 9 1 9 2 9 9 1 13 4 4 2
10 15 1 15 9 1 9 13 4 4 2
11 9 1 1 1 9 14 9 1 1 13 2
11 9 1 0 0 9 1 15 9 13 4 2
8 9 1 15 9 13 9 13 2
27 9 1 13 9 1 9 1 9 13 4 16 9 1 11 7 15 9 11 1 11 1 9 9 14 9 13 2
37 15 1 10 9 9 1 9 11 7 15 9 11 0 12 9 1 1 13 2 15 9 1 11 1 9 11 9 1 1 1 0 9 1 0 13 4 2
18 11 7 11 1 9 1 9 11 1 0 12 0 9 11 11 1 13 2
14 15 1 9 9 11 7 12 0 9 11 11 14 13 2
11 9 1 10 9 1 9 1 0 13 4 2
18 9 1 9 7 15 9 1 0 13 1 1 12 12 1 9 13 4 2
22 11 1 9 1 11 11 7 11 1 13 4 2 7 9 7 15 9 1 0 14 13 2
11 9 1 14 12 9 1 15 9 14 13 2
10 16 2 11 1 9 9 1 9 13 2
42 9 2 9 7 9 9 1 0 9 1 9 13 12 9 1 9 1 1 0 9 1 9 1 1 0 9 9 13 2 7 9 9 13 14 15 9 15 9 14 13 4 2
36 11 2 11 2 9 11 11 1 1 9 0 13 4 7 9 9 1 9 11 11 11 1 9 1 9 9 9 11 1 15 0 9 1 9 13 2
28 11 1 9 1 12 9 1 11 9 11 11 1 12 9 1 9 13 1 9 13 4 15 1 9 0 13 4 2
27 9 1 0 11 11 11 1 1 2 9 0 9 1 11 11 11 1 9 1 0 9 1 9 13 4 4 2
21 15 13 9 9 1 0 9 11 1 11 1 11 11 1 1 11 1 9 13 4 2
45 9 9 1 1 1 11 11 11 1 9 1 9 0 13 1 9 13 1 3 11 9 11 11 11 1 11 1 13 16 15 11 1 9 9 1 1 0 9 1 15 14 9 14 13 2
38 11 11 1 9 1 9 1 1 9 1 1 1 0 9 1 9 9 1 9 13 1 3 15 1 14 11 11 1 11 1 13 1 9 14 0 13 4 2
16 11 1 13 16 15 9 1 15 9 1 9 1 14 13 13 2
27 9 1 11 11 0 13 1 3 11 1 1 1 11 1 9 1 9 13 1 9 13 4 9 0 13 4 2
22 0 9 1 0 9 1 1 11 11 9 1 1 9 1 9 1 0 9 13 4 4 2
32 10 9 1 11 1 11 11 11 11 11 11 11 9 11 11 11 7 9 1 0 9 7 9 9 1 9 1 9 1 9 13 2
59 11 9 1 0 9 11 11 11 1 15 9 1 13 16 9 1 0 9 1 9 1 9 13 9 1 9 13 1 0 9 7 9 14 1 11 1 0 9 1 9 0 13 1 3 0 9 1 0 13 1 1 9 1 0 9 13 4 4 2
33 11 1 13 16 9 13 9 1 13 4 0 9 1 1 1 9 10 0 13 4 4 7 10 9 0 0 9 0 13 4 4 4 2
24 10 9 1 11 11 1 14 0 13 4 4 4 7 9 2 9 1 9 9 13 4 4 4 2
32 11 1 13 16 15 14 0 9 1 13 1 1 0 9 9 9 1 1 12 9 12 9 9 9 1 0 9 9 1 9 13 2
20 15 1 9 1 11 11 7 11 11 1 1 11 1 0 9 1 11 13 4 2
31 10 9 1 11 1 12 0 9 1 12 9 1 1 11 2 9 9 7 0 0 9 1 0 9 1 1 12 9 0 13 2
7 15 12 9 11 1 13 2
26 15 1 11 11 2 11 11 2 11 11 11 11 2 11 2 9 7 11 11 1 9 1 9 13 4 2
11 3 2 11 1 15 1 0 14 13 4 2
23 15 15 1 12 12 9 0 13 4 7 12 12 9 1 0 2 0 9 1 9 13 4 2
20 0 9 7 9 13 1 9 1 0 10 9 9 1 15 14 9 13 4 4 2
15 11 1 12 9 2 0 9 9 7 0 9 14 13 4 2
25 11 1 9 9 1 12 9 9 7 15 9 9 13 1 11 1 11 11 11 1 14 9 13 4 2
8 15 9 13 0 9 13 4 2
37 10 9 1 11 1 9 9 1 9 9 9 11 11 11 2 9 9 9 11 11 11 7 11 11 7 9 11 11 1 9 7 9 1 14 9 13 2
24 10 9 1 1 0 13 4 9 1 11 11 11 1 9 11 11 11 1 14 0 13 4 4 2
23 10 9 11 1 11 11 11 1 12 9 7 9 1 9 13 9 1 0 9 0 13 4 2
23 11 1 9 9 9 11 11 1 9 2 9 1 9 13 4 7 15 1 9 0 13 4 2
16 9 13 16 15 0 9 1 9 1 12 9 1 9 8 13 2
29 11 1 11 1 11 11 11 11 11 1 0 9 11 1 1 12 9 0 13 7 15 9 7 9 1 9 13 4 2
11 15 1 12 12 9 1 9 1 9 13 2
24 11 9 11 11 1 1 2 9 1 9 10 9 1 13 4 2 15 0 9 1 9 13 4 2
18 11 1 11 1 9 1 9 9 11 11 11 1 1 9 0 13 4 2
19 11 10 0 9 1 1 13 9 1 12 12 9 1 9 13 1 9 13 2
16 15 10 9 1 9 1 9 1 12 12 9 1 9 13 4 2
27 11 1 11 11 11 11 11 11 1 11 9 1 9 11 11 1 1 9 1 10 9 1 9 0 13 4 2
21 11 1 9 9 1 9 1 0 10 9 1 1 12 12 9 1 9 13 4 4 2
18 11 1 11 11 1 9 9 1 1 14 9 1 9 0 13 4 4 2
14 9 1 1 15 1 12 12 9 1 9 13 4 4 2
26 11 1 9 1 0 9 9 1 9 1 11 1 9 9 11 11 11 1 1 14 9 0 13 4 4 2
45 11 9 1 13 16 11 1 10 9 1 11 11 11 2 9 2 9 9 2 11 11 2 11 2 11 11 11 2 11 11 11 11 2 11 11 11 11 7 0 9 1 9 13 4 2
16 10 9 1 9 11 1 14 12 9 1 14 0 13 4 4 2
24 9 11 1 11 7 11 9 1 9 1 11 9 1 9 1 9 1 1 9 0 13 4 4 2
21 9 1 11 9 1 9 3 10 13 1 1 10 9 1 9 1 9 1 9 13 2
10 10 9 1 15 9 1 9 13 4 2
27 9 1 1 11 9 1 9 1 9 1 9 1 9 2 9 1 1 10 9 1 9 2 9 14 0 13 2
16 10 9 1 13 0 11 11 1 11 1 11 9 1 9 13 2
31 0 13 16 9 11 9 9 11 11 1 15 9 11 11 1 9 11 1 9 11 9 11 9 11 11 1 1 0 13 4 2
13 11 1 9 11 13 2 7 11 1 9 11 13 2
39 15 1 14 12 9 1 11 9 1 9 1 10 9 1 9 13 4 2 7 3 1 9 1 10 9 1 9 1 10 9 1 1 1 9 14 13 4 4 2
15 9 1 14 1 0 9 1 11 9 1 9 13 4 4 2
27 10 9 1 9 13 1 1 9 1 12 12 9 0 9 7 12 12 9 0 9 1 9 0 13 4 4 2
41 16 10 9 1 9 14 13 4 2 7 9 1 9 1 9 1 9 1 9 13 7 9 1 15 14 9 11 9 1 9 1 15 9 1 15 9 14 13 4 4 2
12 9 1 11 0 0 15 14 9 14 13 4 2
51 7 9 13 4 1 9 1 0 9 13 1 11 11 7 11 11 1 13 16 15 1 15 1 9 14 13 4 4 7 16 11 11 11 1 13 1 9 13 4 4 16 9 1 9 1 0 13 4 4 4 2
22 7 12 9 9 13 1 3 9 1 13 4 11 9 1 9 1 9 14 13 4 4 2
24 11 9 1 9 1 13 13 16 15 15 15 9 14 13 15 13 1 13 1 15 9 14 13 2
12 16 15 9 1 15 14 9 14 13 4 4 2
24 10 13 0 9 1 1 15 1 9 0 11 11 1 11 1 11 9 1 9 1 13 4 4 2
14 10 9 1 1 14 11 9 1 0 9 10 9 13 2
16 3 9 1 11 9 1 9 13 1 9 13 1 13 4 4 2
23 7 11 9 1 9 11 1 13 13 16 15 9 1 9 1 9 0 13 1 1 9 13 2
22 7 9 11 1 11 9 1 9 13 1 9 13 7 14 13 10 9 15 15 13 4 2
39 3 10 9 1 9 1 11 9 1 11 11 1 13 13 16 16 11 9 1 13 4 4 9 1 0 13 4 4 16 15 14 9 2 9 1 9 14 13 2
33 15 13 16 16 11 9 1 9 9 9 1 15 13 4 16 15 10 9 1 15 9 14 13 2 16 9 15 9 0 13 4 4 2
35 9 1 1 1 9 9 11 11 1 13 13 16 9 1 9 1 9 9 9 9 1 13 4 4 4 7 9 1 1 14 15 9 13 4 2
18 11 1 1 15 11 1 9 14 11 11 9 1 1 0 13 4 4 2
14 9 1 9 1 9 1 9 14 13 1 9 13 4 2
17 11 1 10 9 1 9 13 1 1 9 9 11 1 9 13 4 2
27 11 1 0 13 4 11 1 12 0 9 1 9 9 1 9 0 13 1 9 1 0 9 0 13 4 4 2
14 11 1 14 11 9 1 1 11 1 9 0 13 4 2
20 11 9 11 11 1 10 9 1 9 1 9 1 9 14 13 1 9 13 4 2
31 11 1 9 11 11 1 13 13 16 10 9 1 9 1 0 13 9 9 13 10 9 7 9 1 9 1 15 9 14 13 2
20 15 13 13 16 11 11 1 15 9 13 9 9 13 1 9 15 13 4 4 2
27 15 13 16 11 1 9 13 16 9 1 9 1 9 14 13 1 9 9 1 1 11 11 1 0 9 13 2
16 9 1 1 9 13 16 11 11 0 9 1 9 13 4 4 2
30 11 7 11 1 1 14 15 11 7 11 1 14 9 1 9 13 7 9 1 9 1 0 13 1 9 13 4 4 4 2
20 11 1 11 9 1 11 11 1 1 9 1 9 1 0 9 1 9 13 4 2
11 9 1 12 9 7 12 9 0 13 4 2
14 9 1 12 9 14 13 4 7 12 9 0 13 4 2
32 0 9 1 1 12 9 1 10 9 1 13 4 1 9 13 14 9 11 11 11 1 9 1 0 9 1 11 1 1 9 13 2
36 3 14 9 0 9 1 1 13 3 1 0 9 13 4 2 15 9 1 14 9 11 7 12 9 1 9 13 4 2 7 12 9 0 13 4 2
11 9 1 9 1 13 16 9 9 0 13 2
11 9 13 16 9 1 12 14 12 9 13 2
21 12 0 9 1 9 1 11 9 1 11 1 0 9 0 11 1 9 1 9 13 2
12 9 9 1 0 9 13 2 7 9 13 4 2
12 10 9 1 9 9 1 12 9 1 13 4 2
17 15 1 1 12 9 9 9 2 12 10 9 7 9 0 13 4 2
16 12 0 9 1 9 1 9 9 1 9 1 9 1 9 13 2
11 15 15 1 14 0 13 1 9 14 13 2
9 9 1 9 13 9 0 13 4 2
51 9 1 0 9 13 1 15 7 14 12 9 13 4 4 4 2 0 9 1 11 1 11 9 1 9 13 16 15 9 1 0 9 0 9 1 3 13 7 0 9 1 0 13 0 13 16 15 9 13 4 2
41 11 2 11 7 11 11 1 9 1 9 13 16 0 9 1 9 1 0 9 1 9 1 9 13 4 4 4 7 9 0 9 1 15 9 0 13 1 13 4 4 2
24 11 1 9 11 11 11 1 13 16 11 11 1 0 9 1 9 1 0 9 0 13 4 4 2
31 15 16 0 9 1 14 0 9 1 0 13 1 9 13 4 16 9 9 1 1 15 1 13 1 1 0 15 9 14 13 2
42 11 1 0 9 11 11 1 13 16 9 9 1 9 1 13 4 11 11 1 9 16 0 9 1 14 0 9 1 0 13 1 9 13 4 16 15 0 9 0 13 4 2
21 11 1 13 16 11 11 11 11 11 1 15 11 1 9 0 9 1 13 4 4 2
35 11 11 11 1 9 11 11 11 1 13 16 9 9 1 9 13 16 11 9 9 2 0 9 2 9 7 9 1 1 9 1 10 9 13 2
29 11 11 1 9 11 11 1 13 16 9 11 11 11 2 11 2 1 12 9 9 7 12 9 9 1 1 0 13 2
16 11 9 11 11 11 2 11 2 1 14 10 9 13 4 4 2
15 9 9 11 1 9 1 1 11 1 9 13 0 14 13 2
38 16 15 10 9 1 9 13 13 7 14 0 11 1 0 0 0 9 1 13 13 7 0 11 1 9 9 1 13 13 16 15 15 1 0 9 14 13 2
11 3 0 9 1 1 14 15 0 0 13 2
22 11 1 0 11 11 11 0 9 1 9 1 9 1 9 13 1 1 0 13 4 4 2
22 11 1 9 13 16 0 11 1 9 11 11 1 0 0 9 1 9 1 0 13 4 2
16 0 10 9 1 15 0 9 1 9 0 9 1 13 4 4 2
18 3 11 1 11 1 9 1 11 1 9 1 9 1 9 13 4 4 2
31 11 1 0 9 1 0 0 9 11 11 1 9 1 1 1 9 1 9 1 9 1 10 9 1 13 1 9 13 4 4 2
16 0 9 9 9 1 9 1 9 1 1 0 9 1 0 13 2
11 11 1 12 9 1 0 13 4 4 4 2
25 3 0 9 1 12 9 9 0 13 10 9 13 4 16 11 9 1 9 1 9 1 0 14 13 2
14 0 10 9 1 12 9 1 9 1 0 13 4 4 2
23 3 12 0 9 1 9 1 13 13 16 0 9 15 9 1 9 1 9 0 13 4 4 2
20 11 1 14 15 12 9 7 15 0 9 1 9 1 1 9 1 9 13 4 2
20 11 1 1 1 13 4 4 16 9 1 0 9 1 1 1 9 13 4 4 2
15 0 9 1 10 14 10 12 0 9 1 0 13 4 4 2
11 15 1 12 1 10 9 13 4 4 4 2
33 16 15 12 0 9 13 7 15 9 1 9 7 9 1 15 9 9 13 4 16 3 9 9 1 13 1 1 3 9 1 9 13 2
12 13 4 4 9 3 15 9 1 9 13 4 2
12 9 1 9 9 1 10 9 1 9 0 13 2
17 9 15 13 16 9 1 9 13 1 1 9 9 13 4 4 4 2
48 9 13 4 16 9 1 0 13 1 0 9 0 9 1 9 14 13 2 0 9 1 9 1 9 7 0 0 9 14 13 1 3 14 9 1 0 9 13 1 14 3 9 1 9 13 14 13 2
31 16 9 1 9 1 9 13 4 0 9 1 9 9 9 1 9 13 4 4 2 15 9 1 9 1 3 9 13 4 4 2
31 11 11 11 1 13 4 4 0 9 9 1 0 9 9 11 11 13 4 16 9 1 9 14 12 2 12 0 9 13 4 2
29 12 9 9 14 9 1 14 9 13 13 4 4 4 7 10 9 1 9 1 9 1 9 13 1 9 13 4 4 2
19 11 13 4 16 15 9 15 9 1 9 14 13 15 9 3 9 1 13 2
42 11 11 11 11 11 1 11 1 13 16 0 11 11 11 1 13 9 1 0 12 9 1 13 10 0 0 9 1 9 1 13 1 1 9 1 12 12 9 1 9 13 2
28 11 1 13 16 0 12 9 1 11 1 13 0 9 1 13 9 1 9 13 1 1 3 0 9 1 9 13 2
16 0 9 1 13 9 1 9 1 1 12 12 9 1 9 13 2
20 7 0 0 9 1 13 9 1 9 1 1 14 12 12 12 9 1 9 13 2
38 11 1 11 11 11 2 11 2 7 11 1 0 9 2 11 11 11 11 11 2 1 13 16 0 0 9 10 9 1 0 9 1 9 13 1 0 13 2
18 15 13 16 9 9 15 9 1 9 13 7 11 11 15 15 9 13 2
27 11 1 0 9 11 11 1 9 14 1 0 9 1 9 1 9 1 1 11 11 1 9 1 3 9 13 2
34 9 1 11 11 1 1 11 1 0 9 1 11 1 11 9 1 9 1 9 13 4 9 1 1 0 9 9 1 1 9 1 9 13 2
32 11 1 13 16 11 1 11 1 11 1 1 1 12 9 1 9 0 13 1 9 1 1 1 0 9 1 1 0 9 13 4 2
20 15 13 16 9 1 9 1 15 0 13 4 4 16 9 1 9 1 9 13 2
26 9 1 9 1 1 9 10 9 13 13 4 16 15 14 9 1 9 1 9 1 9 1 13 4 4 2
13 15 13 16 15 9 1 15 13 1 9 14 13 2
9 15 0 9 1 9 13 13 4 2
19 0 9 1 9 1 9 13 2 7 0 9 1 1 15 9 1 14 13 2
28 15 13 16 16 9 12 9 1 9 1 9 9 1 9 13 1 0 13 4 16 15 9 9 1 9 9 13 2
24 11 1 13 16 9 1 13 12 9 0 13 4 4 2 7 15 9 13 1 14 13 4 4 2
14 0 9 1 1 15 9 1 10 12 9 1 9 13 2
32 11 11 7 15 9 1 9 1 9 13 4 15 13 16 15 14 0 9 13 4 4 7 9 1 9 9 1 9 13 4 4 2
14 15 13 16 9 0 11 9 1 9 1 13 4 4 2
21 11 1 0 9 11 11 2 0 9 11 11 7 11 11 1 14 9 1 0 13 2
38 11 11 11 1 11 1 13 16 11 11 11 1 0 0 9 1 9 1 1 9 9 1 9 9 0 13 1 11 1 1 1 9 14 13 4 4 4 2
37 11 11 1 0 9 1 9 9 1 1 11 11 1 0 9 9 1 1 1 9 13 1 3 11 1 9 1 13 16 15 1 1 15 9 14 13 2
30 15 1 11 1 11 1 11 1 0 13 1 12 9 11 2 11 7 11 11 11 1 9 9 0 13 1 9 13 4 2
43 9 9 11 11 11 1 11 1 11 11 1 9 13 16 15 11 1 13 11 11 11 2 11 2 1 9 1 11 1 12 12 9 1 9 1 9 13 1 0 0 13 4 2
35 15 0 2 0 9 1 11 1 13 16 15 11 1 0 9 13 4 4 15 11 11 11 11 1 13 4 11 11 11 1 9 13 4 4 2
19 11 11 11 11 11 1 11 1 9 9 11 1 9 13 1 14 9 13 2
25 9 1 1 1 0 9 9 1 11 1 13 16 9 1 11 1 9 1 14 12 9 1 9 13 2
22 15 9 13 16 11 1 9 9 1 9 0 13 1 9 13 2 15 13 4 4 4 2
23 15 9 1 15 15 9 14 13 4 2 7 11 0 9 1 0 13 1 9 14 13 4 2
27 15 13 7 14 9 0 9 1 0 9 0 13 7 15 1 9 1 11 1 14 9 1 9 9 13 4 2
44 11 1 9 13 16 11 11 1 9 13 16 11 15 9 9 1 9 1 9 13 1 12 12 9 0 13 4 2 7 11 1 9 1 14 1 14 10 9 1 0 9 13 4 2
21 15 13 16 16 9 13 14 4 16 11 7 0 9 7 15 9 1 14 9 13 2
13 15 9 1 12 12 9 1 15 9 14 13 4 2
37 11 1 13 16 11 9 1 1 11 1 11 1 0 9 9 1 9 13 14 0 14 13 2 7 15 9 1 1 12 9 11 11 11 13 13 4 2
23 10 9 11 11 11 1 9 13 4 15 9 1 9 1 9 1 9 15 13 4 4 4 2
14 15 11 11 1 11 11 1 9 1 14 0 9 13 2
21 9 1 11 11 1 13 16 11 1 9 1 9 1 1 9 1 9 1 9 13 2
15 15 9 11 1 9 9 11 1 0 11 11 1 13 4 2
27 15 13 16 11 1 11 11 1 13 1 9 1 1 9 9 10 9 1 11 1 12 0 9 14 0 13 2
34 11 11 11 1 9 11 11 1 11 1 0 2 0 9 9 7 11 11 9 1 1 11 9 1 9 13 11 9 1 9 13 4 4 2
17 11 1 10 9 1 11 1 0 9 13 1 9 13 4 4 4 2
18 3 11 11 1 0 9 9 11 11 1 11 1 0 9 13 13 4 2
17 7 11 1 10 9 1 11 1 10 9 1 9 1 13 4 4 2
18 11 1 11 1 9 2 9 9 1 11 9 11 11 9 13 4 4 2
14 10 9 0 9 11 11 1 9 1 1 0 13 4 2
20 7 11 1 9 13 4 1 9 1 11 11 11 11 11 1 9 13 4 4 2
13 11 1 10 12 9 1 11 9 13 1 0 13 2
35 16 11 13 4 16 10 12 9 1 11 1 9 13 1 1 1 11 0 9 9 7 11 9 11 11 1 11 11 9 1 1 15 9 13 2
8 3 11 1 11 9 0 13 2
16 11 7 11 1 10 9 1 11 1 0 9 1 11 13 4 2
29 15 11 1 11 1 9 13 2 15 11 1 11 1 13 11 11 1 9 13 4 4 7 11 9 1 9 13 4 2
12 7 11 11 1 9 13 1 9 1 14 13 2
18 15 11 1 11 9 1 9 13 11 1 0 9 13 1 9 13 4 2
30 16 16 11 11 1 11 1 9 14 13 4 16 11 10 9 1 0 9 1 1 13 4 7 15 0 9 11 1 13 2
27 16 11 1 0 9 7 9 11 11 11 1 13 13 16 15 11 1 9 7 9 1 1 9 13 4 4 2
16 15 1 1 11 1 11 1 11 11 7 11 1 9 13 4 2
26 15 15 9 1 9 13 4 4 15 15 15 0 9 1 14 9 13 4 7 15 9 9 1 9 13 2
25 11 11 1 9 1 0 9 1 0 9 7 9 9 11 11 11 1 0 11 11 11 0 13 4 2
20 0 9 9 7 11 7 11 1 11 1 9 13 4 11 11 11 1 9 13 2
13 11 11 11 1 9 1 11 10 0 13 4 4 2
23 3 9 9 1 1 11 1 9 2 9 7 9 9 1 0 9 0 13 1 9 13 4 2
10 11 11 1 0 9 9 1 13 4 2
9 15 11 1 11 1 0 9 13 2
17 15 1 15 11 2 11 7 11 1 14 11 1 9 13 4 4 2
17 15 11 2 11 2 11 7 11 1 9 1 1 1 9 13 4 2
13 11 1 11 1 9 1 15 9 9 0 13 4 2
10 15 9 9 1 11 1 0 0 13 2
17 0 9 1 15 11 11 11 11 1 9 9 1 9 1 9 13 2
23 11 9 11 11 11 11 11 11 2 11 2 1 9 1 1 0 9 1 9 13 4 4 2
15 15 1 11 9 9 1 9 1 0 9 13 4 13 4 2
30 9 1 1 9 1 9 1 13 9 1 9 9 9 1 0 9 13 1 9 1 9 9 1 0 13 1 13 9 13 2
19 15 1 14 9 1 9 1 9 1 9 9 13 1 14 11 10 0 13 2
24 16 0 9 1 9 1 15 10 9 14 13 7 15 1 10 9 1 0 13 4 1 9 13 2
37 11 9 1 11 11 11 2 11 11 2 11 7 11 11 1 11 9 1 0 13 4 1 1 11 15 9 1 0 0 13 1 10 9 13 14 13 2
28 9 1 1 2 9 0 9 1 9 1 10 9 13 13 4 7 15 10 0 9 13 1 9 14 13 4 4 2
34 9 1 0 9 1 11 1 0 9 11 1 9 9 13 1 9 13 1 1 11 1 9 13 4 16 15 15 10 9 14 13 4 4 2
30 0 13 16 3 11 1 12 9 1 9 11 1 0 13 1 9 13 4 4 2 7 15 15 11 1 14 0 13 4 2
12 9 1 14 12 11 9 10 9 1 9 13 2
31 9 1 11 2 11 2 11 2 11 7 11 1 0 9 9 1 9 1 9 7 9 1 0 13 1 9 1 9 13 4 2
23 9 1 1 2 0 9 11 7 11 1 11 1 0 9 7 0 9 13 1 14 9 13 2
39 11 9 11 11 1 0 0 7 11 1 11 2 11 11 11 11 1 12 9 3 11 13 1 9 1 9 1 9 3 14 3 13 1 9 0 13 4 4 2
40 11 11 9 1 9 9 1 9 1 9 1 9 15 9 13 4 1 0 13 9 9 11 13 11 1 11 1 13 0 9 1 1 15 9 13 9 13 4 4 2
52 16 0 9 1 9 1 13 4 15 10 9 9 1 9 13 4 4 2 7 0 9 1 13 13 16 11 1 9 0 9 11 11 11 2 9 9 11 11 7 11 9 1 9 9 11 11 1 13 15 9 13 2
31 11 1 9 1 1 9 13 4 13 16 15 1 11 11 11 1 9 9 7 15 11 11 11 1 9 14 3 0 9 13 2
35 9 1 1 2 11 1 0 9 1 13 16 15 14 11 11 1 9 1 13 4 9 9 1 9 9 1 1 14 9 1 9 0 13 4 2
32 9 13 4 16 11 15 11 9 1 1 9 9 11 11 1 13 1 9 1 13 16 9 1 9 11 11 1 9 13 4 4 2
11 15 10 10 0 9 1 14 13 4 4 2
34 11 9 1 15 14 9 13 16 11 0 9 1 9 13 11 1 0 9 1 13 1 0 9 1 15 9 1 3 1 9 13 4 4 2
22 9 9 1 10 9 0 9 1 13 12 9 13 7 15 9 13 12 1 13 4 4 2
34 15 10 9 1 13 4 11 1 15 1 9 9 13 4 4 16 9 1 9 1 0 13 1 9 1 15 9 1 0 14 13 4 4 2
25 11 1 9 1 9 1 1 11 9 1 9 7 11 1 13 9 1 9 1 0 9 13 4 4 2
23 7 11 9 11 1 9 1 13 9 1 13 9 1 0 9 1 1 1 0 13 4 4 2
25 0 3 11 9 9 9 1 0 9 1 1 11 1 9 1 13 0 9 1 13 14 4 4 4 2
51 16 10 9 1 0 9 1 15 1 9 11 11 11 1 15 0 9 14 13 4 2 7 13 4 4 16 11 11 7 11 1 13 9 1 10 0 13 7 9 13 14 15 15 9 13 1 14 9 1 13 2
27 9 1 12 0 9 1 13 16 9 9 1 11 1 11 1 9 1 12 0 9 11 1 0 9 14 13 2
18 9 9 9 1 13 12 9 1 1 13 4 9 1 14 10 0 13 2
18 11 1 9 13 14 11 11 1 9 3 14 13 1 9 14 13 4 2
35 9 11 1 9 11 11 1 2 9 9 2 1 0 13 1 9 13 4 0 9 1 9 1 13 4 16 11 1 15 0 9 14 13 4 2
16 3 15 9 1 9 13 7 15 15 0 9 0 13 4 4 2
22 10 3 9 1 13 4 16 11 11 11 11 1 11 1 13 4 16 3 13 15 4 2
22 0 9 1 9 9 9 9 11 11 1 9 1 13 16 15 15 11 1 9 13 4 2
22 11 1 15 13 16 11 1 9 1 9 1 9 13 1 15 9 1 9 13 4 4 2
13 15 9 1 0 13 4 15 9 0 13 4 4 2
21 11 1 13 16 11 1 9 0 9 13 1 14 13 2 15 14 9 1 13 4 2
21 15 13 16 10 9 1 0 9 1 14 13 4 4 7 9 15 0 13 4 4 2
42 0 13 16 12 9 9 1 11 11 1 11 1 9 9 1 1 9 1 1 9 1 0 13 4 0 9 11 11 1 9 1 1 3 1 9 0 13 4 13 4 4 2
11 11 1 9 11 1 1 9 13 4 4 2
26 16 10 9 11 1 9 1 1 0 13 4 2 3 11 11 1 9 1 15 15 9 9 14 13 4 2
29 11 1 9 1 9 1 0 13 1 12 0 9 9 1 9 9 1 15 9 2 12 9 9 9 2 1 13 4 2
9 0 9 1 14 10 9 13 4 2
34 11 9 11 11 1 9 7 11 11 11 1 9 9 1 9 1 1 11 1 13 0 9 9 1 9 9 1 9 1 9 14 13 4 2
14 9 9 1 9 9 1 1 11 9 1 9 13 4 2
27 9 9 1 9 1 0 2 0 9 1 13 4 16 12 9 0 11 9 1 1 9 9 13 0 14 13 2
23 11 1 3 13 4 13 4 16 11 1 1 1 9 1 9 9 1 13 1 9 14 13 2
12 3 11 1 13 16 9 15 14 13 4 4 2
25 0 3 11 7 11 11 1 13 13 16 11 11 11 1 9 1 13 1 15 9 2 9 14 13 2
28 11 1 9 11 11 11 1 13 2 15 13 13 16 11 9 9 14 13 16 15 11 1 15 0 9 14 13 2
23 9 1 12 9 1 13 4 9 9 1 9 1 11 1 13 16 10 15 9 1 9 13 2
21 11 1 0 9 9 11 11 11 1 13 16 11 1 10 14 9 13 4 4 4 2
12 11 10 9 7 9 1 15 14 13 4 4 2
17 7 15 10 9 1 12 9 1 13 1 9 9 1 9 13 4 2
19 11 1 9 11 11 7 11 11 1 11 11 1 14 9 9 1 9 13 2
21 11 1 13 16 0 11 2 11 2 11 7 11 9 1 11 1 15 9 14 13 2
29 11 1 0 9 11 11 1 13 11 10 9 0 9 13 4 16 9 9 1 15 0 9 13 1 15 9 14 13 2
15 15 1 14 11 9 1 11 1 9 15 0 14 13 4 2
24 11 11 1 11 7 11 1 9 13 7 15 1 15 14 9 11 1 9 13 1 0 14 13 2
13 7 11 11 2 11 7 11 1 11 1 9 13 2
21 15 13 16 14 11 1 11 1 9 1 12 9 13 15 15 0 9 13 4 4 2
22 0 11 1 13 4 11 1 12 10 9 1 9 1 13 1 11 1 0 9 13 4 2
41 9 11 11 7 9 11 11 1 1 9 1 11 11 11 11 2 11 2 1 0 9 11 11 1 0 9 13 4 11 7 9 1 0 9 11 11 1 3 9 13 2
21 11 1 11 2 11 9 1 0 9 13 4 13 16 15 3 9 9 1 9 13 2
26 15 13 16 11 1 0 9 2 9 1 9 1 8 13 1 1 0 7 0 9 1 11 14 0 13 2
31 9 1 9 13 1 9 1 15 0 9 1 9 9 11 11 7 11 9 1 9 1 9 13 11 11 1 14 3 9 13 2
22 11 1 13 1 9 1 9 9 1 9 1 1 11 1 10 9 0 13 4 4 4 2
7 11 14 9 1 9 13 2
19 10 9 1 9 7 9 1 15 9 13 1 1 3 2 3 13 4 4 2
16 3 11 1 11 1 13 4 9 1 9 13 1 9 13 4 2
41 11 1 0 9 1 13 11 1 11 0 13 1 3 9 9 1 9 1 15 1 1 13 4 9 1 9 1 3 0 13 16 15 10 9 1 15 9 14 13 13 2
33 11 1 11 11 11 2 11 7 11 9 9 1 11 1 9 1 9 0 13 11 11 1 11 11 1 13 4 9 1 9 13 4 2
40 9 1 9 9 0 13 4 12 0 9 9 11 11 11 7 11 11 11 1 13 1 9 13 1 3 14 11 1 9 11 11 1 1 13 1 9 13 4 4 2
7 9 1 11 1 9 13 2
45 9 1 15 9 1 12 9 1 13 4 14 9 11 11 11 1 11 9 13 1 9 13 4 4 2 7 9 13 4 16 9 1 12 0 9 1 13 4 9 1 14 0 13 4 2
16 12 0 9 1 14 12 9 1 9 13 1 1 0 13 4 2
45 11 1 11 11 11 11 1 11 1 0 9 9 1 11 1 9 13 4 13 16 11 1 9 1 3 9 13 1 9 13 7 15 14 9 15 13 16 15 11 1 0 9 0 13 2
20 11 15 0 9 13 4 4 16 15 15 14 13 2 15 15 15 13 14 4 2
25 16 2 11 1 0 9 9 1 9 1 9 7 9 1 14 9 13 1 9 13 1 9 13 4 2
21 0 13 16 11 11 11 1 11 9 1 1 11 7 11 1 1 9 3 13 4 2
42 11 1 9 13 4 13 16 11 1 9 13 1 1 1 11 1 13 9 1 9 9 9 9 13 1 3 15 14 13 2 9 1 9 13 1 3 14 10 9 15 13 2
35 11 1 13 16 15 9 1 1 13 4 4 16 16 11 10 9 1 9 14 13 4 16 15 9 1 1 13 9 1 9 9 1 14 13 2
26 15 13 16 9 9 11 11 11 1 10 9 1 9 13 4 16 0 9 2 9 11 1 1 15 13 2
9 11 11 1 11 1 3 9 13 2
24 11 7 11 9 1 1 9 1 9 1 13 4 9 1 11 1 9 1 9 1 1 13 4 2
34 11 9 11 11 11 2 11 11 7 11 11 11 11 1 11 9 1 1 9 13 13 4 7 12 9 11 9 11 11 1 13 14 4 2
13 10 11 9 1 11 1 9 13 4 14 13 4 2
32 11 1 10 9 11 9 1 1 13 4 7 9 1 9 1 1 13 13 9 11 11 1 15 9 1 1 13 1 9 13 4 2
29 9 1 1 9 11 11 1 11 11 11 1 1 13 4 13 4 2 7 15 11 1 1 13 1 3 13 4 4 2
22 11 11 11 11 11 11 11 11 7 11 9 11 11 1 11 1 9 13 4 13 4 2
27 11 1 9 1 9 1 1 13 4 1 3 9 1 13 16 11 9 1 0 9 1 1 0 13 4 4 2
24 11 9 9 1 9 11 11 7 11 9 11 1 9 1 15 9 1 9 13 1 9 13 4 2
22 11 11 11 1 13 16 11 9 1 15 9 1 9 13 1 9 15 0 13 4 4 2
24 9 1 13 16 0 9 1 1 1 9 13 1 1 15 11 1 9 9 1 9 1 9 13 2
27 11 1 15 9 1 9 9 13 15 11 9 11 11 11 1 9 1 9 9 1 9 1 9 13 4 4 2
15 11 9 3 3 1 13 4 2 15 10 9 13 13 4 2
18 15 1 11 1 13 16 15 15 9 0 13 4 15 1 9 9 13 2
10 15 1 12 9 1 9 9 13 4 2
20 11 1 11 11 1 11 9 1 9 0 9 11 11 1 9 9 0 13 4 2
29 10 9 1 9 9 1 0 12 9 11 1 9 11 11 7 9 1 9 11 11 1 9 9 14 9 13 4 4 2
17 11 1 11 11 1 0 11 11 1 11 11 1 0 13 4 4 2
17 11 9 1 0 9 11 11 9 1 3 13 15 9 1 13 4 2
23 15 13 16 15 9 7 9 1 1 10 10 14 9 13 2 15 9 1 9 1 13 4 2
15 15 9 1 13 16 15 11 1 1 1 15 9 14 13 2
24 15 1 9 9 1 0 9 11 11 1 13 9 13 0 9 13 4 11 9 1 3 9 13 2
33 9 9 1 9 9 0 14 13 4 2 15 1 9 1 0 9 13 7 11 1 9 9 13 1 9 1 13 4 15 9 13 4 2
17 15 9 1 9 1 3 1 9 1 1 11 1 9 13 4 4 2
18 10 9 1 0 9 11 11 1 11 9 1 9 11 1 9 13 4 2
14 15 1 11 9 1 11 7 9 11 9 13 4 4 2
20 15 1 11 9 1 9 11 1 9 1 9 1 15 9 1 9 13 4 4 2
24 11 1 9 1 9 13 4 1 3 15 11 11 11 1 9 1 9 1 13 1 9 13 4 2
9 15 11 11 1 9 1 0 13 2
20 15 11 9 1 9 13 4 13 16 11 9 1 11 9 1 9 14 14 13 2
23 11 9 9 1 9 13 4 4 7 9 1 10 9 1 14 9 3 13 15 9 13 4 2
24 11 1 11 9 1 11 1 0 12 0 9 1 0 9 11 11 1 11 9 1 0 13 4 2
16 10 9 1 11 11 11 1 9 1 1 14 0 13 4 4 2
37 9 1 15 0 9 1 13 16 10 9 1 9 7 11 1 9 9 1 9 1 9 13 1 11 11 11 2 11 2 1 9 9 9 1 13 4 2
15 9 1 9 0 13 1 1 9 1 10 14 9 14 13 2
15 15 1 9 1 9 9 11 2 11 2 11 7 11 13 2
33 9 1 1 9 1 0 9 1 9 13 16 0 9 1 9 0 9 1 13 4 4 7 15 11 11 1 11 9 1 13 4 4 2
30 11 7 11 11 1 10 12 9 1 0 13 4 4 7 11 9 1 0 0 9 1 1 15 1 1 0 13 4 4 2
20 15 1 9 9 1 9 1 9 1 15 9 13 7 15 15 9 13 4 4 2
43 15 12 9 1 9 1 2 0 9 2 13 1 7 11 1 9 1 9 13 1 11 11 11 7 11 11 11 11 1 11 11 11 1 12 0 9 9 13 1 9 13 4 2
14 10 9 1 9 2 9 7 9 9 1 14 9 13 2
25 15 9 13 16 9 0 13 1 1 15 10 11 1 12 9 1 1 9 9 9 1 9 1 13 2
37 11 11 11 11 11 1 11 1 13 16 2 11 1 9 1 9 1 13 4 9 14 10 9 1 12 9 9 13 15 3 11 2 11 1 9 13 2
16 10 9 1 11 1 0 9 9 2 9 2 9 7 9 14 13
24 9 1 3 13 16 2 11 1 9 0 9 1 1 10 13 7 0 9 1 15 0 9 13 2
17 15 15 12 0 9 9 13 1 1 10 9 1 9 1 9 13 4
27 11 1 13 4 16 11 11 11 1 9 1 13 1 3 14 15 9 9 13 1 9 9 1 9 13 4 2
20 9 1 9 7 11 1 9 1 1 3 13 9 1 11 1 9 13 4 4 2
27 9 1 13 1 3 3 15 11 11 14 13 4 4 16 15 1 9 7 11 1 9 1 1 9 0 13 2
14 15 11 11 9 9 1 11 1 0 9 13 4 4 2
31 11 11 11 1 9 1 10 9 1 13 1 1 9 0 13 1 1 0 9 1 0 9 7 9 9 11 11 1 15 13 2
31 11 11 1 9 15 14 13 4 16 9 15 0 2 0 9 1 9 13 1 3 14 11 1 9 1 1 9 13 4 4 2
19 0 9 1 15 1 9 0 0 9 1 15 9 13 1 9 13 4 4 2
15 7 9 1 0 9 1 11 1 9 1 9 13 4 4 2
22 11 11 11 11 11 13 4 16 0 9 1 15 1 9 1 9 13 1 9 13 4 2
20 9 15 13 16 0 9 15 1 12 9 1 12 9 1 15 9 13 4 4 2
16 11 11 1 9 1 9 2 9 13 9 13 1 9 13 4 2
16 15 1 10 9 1 10 9 11 11 1 11 1 9 13 4 2
25 9 1 11 11 11 1 9 1 0 9 1 0 9 7 9 9 1 13 12 9 9 13 4 4 2
28 10 9 9 1 0 13 1 1 11 11 11 1 9 1 0 9 1 11 1 0 9 1 9 1 9 13 4 2
19 10 9 1 11 1 9 1 0 9 1 13 9 1 9 14 0 13 4 2
20 11 1 11 11 11 1 9 9 11 11 1 9 13 1 9 1 0 13 4 2
33 11 1 9 11 11 1 13 16 11 1 0 11 11 11 1 9 9 11 11 1 9 13 1 9 1 11 1 11 1 0 13 4 2
25 11 1 15 1 12 9 1 0 13 1 1 11 1 12 9 1 12 12 9 13 1 9 13 4 2
20 11 11 11 11 11 11 1 11 9 1 1 9 1 0 9 13 4 4 4 2
27 11 11 11 1 15 11 9 1 1 11 1 11 11 11 11 7 11 1 11 11 1 9 9 1 0 13 2
25 11 1 9 9 11 11 11 1 11 1 13 16 11 1 9 1 9 1 9 15 9 14 13 13 2
19 9 1 9 9 11 11 11 7 9 9 11 11 11 11 1 9 11 13 2
20 15 15 9 1 9 13 1 3 14 9 9 1 13 4 4 9 1 9 13 2
25 11 11 11 15 11 13 7 9 1 9 13 1 3 9 9 1 9 9 1 9 9 13 1 13 2
14 11 1 11 11 11 11 1 11 11 1 9 9 13 2
12 15 14 11 1 9 1 1 9 9 1 13 2
26 11 11 1 0 11 11 7 15 0 9 9 1 1 9 1 9 1 9 10 0 9 1 13 4 4 2
17 16 15 0 13 4 16 15 9 1 1 13 1 13 14 4 4 2
19 10 9 11 1 15 9 1 12 9 11 11 7 11 11 1 9 1 13 2
17 12 9 11 11 1 0 9 1 9 13 1 3 0 13 4 4 2
37 15 13 16 9 1 11 11 9 1 9 1 1 0 9 13 4 2 7 10 9 1 9 1 9 0 13 7 15 9 1 9 1 15 9 14 13 2
16 15 0 13 14 10 9 1 9 0 13 4 15 0 13 4 2
29 11 11 11 11 11 11 11 1 13 16 9 11 2 11 1 11 9 1 1 13 9 9 1 9 1 9 13 4 2
18 15 0 13 4 9 7 9 9 1 12 9 1 0 13 4 4 4 2
27 11 1 13 16 9 1 9 1 10 0 9 1 9 1 1 13 4 9 1 11 11 1 15 0 9 13 2
42 15 9 13 16 0 11 11 1 9 1 0 0 9 0 13 1 1 15 9 7 9 1 0 9 13 4 7 10 9 1 9 2 9 7 9 9 13 1 9 13 4 2
19 9 1 9 2 9 2 9 2 9 7 9 1 15 9 1 0 13 4 2
20 0 11 11 11 11 1 0 11 9 1 12 9 1 1 9 9 1 9 13 2
14 9 1 1 9 9 1 9 1 10 9 1 9 13 2
17 11 11 1 11 0 11 11 11 11 11 11 1 9 1 9 13 2
17 11 7 11 1 9 1 0 9 1 1 10 9 1 0 13 4 2
16 0 9 9 9 1 1 0 9 9 1 9 9 0 13 4 2
24 11 1 9 1 0 0 9 9 11 11 1 11 1 11 11 1 9 13 1 0 9 13 4 2
34 11 11 11 11 2 11 2 1 9 11 11 1 13 16 11 1 9 1 12 9 1 9 9 7 9 9 1 1 9 1 0 9 13 2
26 15 13 16 9 9 2 11 11 11 11 2 9 1 1 9 9 9 7 9 9 9 1 9 13 4 2
20 0 9 11 1 11 11 11 7 0 9 9 1 1 12 9 1 9 13 4 2
21 14 12 0 9 1 11 1 12 9 9 7 9 9 1 1 9 1 9 13 4 2
31 11 1 11 9 1 1 11 9 1 13 9 1 13 4 9 1 9 1 1 0 9 1 9 1 9 13 1 9 13 4 2
14 16 9 1 15 1 1 9 1 15 9 14 13 4 2
11 10 9 11 9 1 1 11 9 1 13 2
29 11 1 0 9 11 1 13 13 16 16 9 1 0 9 1 13 4 9 1 0 9 1 1 1 15 9 14 13 2
11 15 13 13 16 10 9 1 9 0 13 2
23 11 1 9 9 11 11 11 1 13 13 16 15 9 1 9 1 1 1 15 9 14 13 2
13 15 3 10 9 1 9 13 1 9 13 4 4 2
24 10 9 1 11 1 9 9 11 11 11 1 13 16 15 15 1 9 1 12 9 13 4 4 2
15 10 9 1 13 9 1 9 1 14 15 15 13 4 4 2
17 11 11 11 1 0 9 1 9 9 1 9 1 9 13 4 4 2
12 15 13 16 15 10 9 1 9 1 13 4 2
27 11 1 0 0 9 1 9 9 11 11 1 13 13 16 9 1 9 1 9 13 10 9 7 9 13 4 2
13 15 13 16 15 0 9 1 15 9 13 4 4 2
24 11 1 13 16 15 11 1 15 1 1 9 0 13 10 9 1 3 14 9 13 1 9 13 2
13 9 9 1 1 13 9 0 9 2 9 13 4 2
52 3 9 14 11 11 1 9 1 9 9 1 9 1 13 4 2 3 9 1 9 1 9 1 13 0 9 2 11 1 11 0 13 1 11 1 9 7 11 11 11 11 14 1 13 11 11 9 1 9 1 13 2
30 10 9 1 1 10 9 9 9 7 9 1 9 14 13 7 0 9 1 15 9 15 13 16 15 9 1 1 9 13 2
15 9 1 9 1 14 11 11 1 9 1 9 0 13 4 2
18 9 1 0 9 1 15 13 0 9 1 9 9 1 0 13 4 4 2
19 15 1 9 1 3 2 3 14 9 1 11 11 1 12 12 9 13 4 2
34 10 9 1 13 9 13 16 0 9 9 1 11 11 1 9 13 1 9 13 4 7 9 1 9 1 15 1 1 9 9 14 13 4 2
13 11 11 9 11 11 15 9 1 13 9 1 13 2
16 15 9 14 0 2 0 13 7 0 15 0 9 14 13 4 2
35 3 15 14 9 1 9 1 9 13 1 9 13 7 9 1 0 9 1 1 3 9 10 9 14 13 4 7 0 9 1 1 15 0 13 2
24 3 1 15 11 9 1 11 13 1 9 13 4 15 11 11 11 1 9 1 1 9 13 4 2
10 0 14 9 9 15 9 1 13 4 2
26 9 1 9 1 9 1 9 1 9 1 14 11 11 11 11 1 9 1 1 10 9 9 14 13 4 2
13 15 0 11 11 1 15 1 9 13 1 9 13 2
23 11 9 1 9 1 9 1 1 15 9 1 0 13 1 14 0 13 7 0 14 13 4 2
9 15 9 9 1 1 13 4 4 2
20 9 1 1 1 11 2 9 9 7 9 1 13 9 2 9 1 9 13 4 2
29 9 9 9 1 13 14 11 1 15 1 13 16 15 9 9 13 7 9 1 9 13 1 15 10 15 9 14 13 2
30 10 9 15 9 9 11 1 0 9 1 0 13 7 9 9 11 1 1 0 9 13 1 1 14 11 0 9 1 13 2
21 11 11 1 0 9 1 1 11 9 1 0 13 1 9 14 10 9 13 14 4 2
17 11 1 9 9 1 13 14 11 11 1 0 9 1 9 13 4 2
31 11 11 11 1 12 9 1 9 1 0 9 13 7 9 1 0 9 1 9 13 1 14 9 9 1 9 1 0 9 13 2
25 11 11 1 11 1 11 11 9 1 9 9 1 9 1 9 1 9 1 9 1 0 9 13 4 2
12 9 1 0 9 9 0 13 1 9 13 4 2
9 11 11 1 13 2 15 0 13 2
23 0 13 16 11 9 1 9 1 9 1 1 9 9 0 13 1 3 9 13 4 4 4 2
15 7 3 1 10 9 1 9 1 9 1 9 0 13 4 2
11 9 1 9 1 9 1 9 1 9 13 2
40 0 9 1 9 1 9 1 9 13 4 7 3 1 11 11 11 1 15 9 1 0 9 9 14 0 14 13 2 7 9 1 1 0 9 0 13 1 9 13 2
30 11 11 1 9 1 9 1 9 1 13 4 12 0 9 1 13 4 16 0 9 1 9 1 3 9 14 13 4 4 2
9 9 1 9 13 4 3 0 13 2
14 15 9 13 4 4 16 9 1 9 1 9 13 4 2
56 9 11 11 11 7 9 11 11 11 1 9 1 11 11 1 9 1 9 13 1 11 11 11 11 7 9 1 9 9 13 4 9 1 9 1 0 13 4 7 9 11 11 1 9 1 0 13 4 13 16 15 0 9 13 4 2
20 9 1 15 0 9 1 13 16 9 1 15 1 9 1 9 13 0 9 13 2
25 9 1 13 16 3 14 9 1 9 1 9 14 0 13 4 4 15 1 9 1 9 1 9 13 2
25 15 9 1 13 0 9 1 15 0 14 13 16 9 1 14 15 9 1 9 13 1 9 13 4 2
9 9 1 9 1 13 4 0 13 2
29 11 11 1 13 9 13 1 0 0 9 1 1 9 13 1 9 13 1 11 11 1 0 9 1 9 13 4 4 2
31 9 1 9 1 9 1 1 0 9 1 9 13 4 11 11 2 11 9 7 9 9 2 11 11 2 1 9 0 13 4 2
8 9 9 1 14 9 13 4 2
32 9 1 9 13 4 4 16 9 1 0 9 2 9 9 7 0 9 1 1 9 13 4 1 9 0 9 1 0 13 4 4 2
45 9 9 11 11 11 2 9 11 11 11 7 9 11 11 11 1 9 1 11 1 11 11 11 7 11 11 11 7 9 1 12 9 1 9 13 4 11 11 1 9 1 9 13 4 2
22 11 11 10 0 9 1 9 14 1 0 9 9 7 9 1 9 1 13 4 9 13 2
69 11 11 1 11 11 2 11 1 9 7 11 11 11 1 0 9 1 9 1 1 0 9 1 9 9 1 9 7 9 1 0 0 0 9 1 9 13 4 11 11 11 11 2 11 11 11 2 11 2 11 11 11 2 11 11 11 7 11 11 1 15 0 9 1 9 13 4 4 2
23 11 11 1 13 4 9 13 1 9 1 0 9 1 1 9 13 1 15 9 0 13 4 2
28 10 9 1 11 11 11 2 11 11 11 7 11 11 11 1 1 9 13 2 15 9 9 1 0 13 4 4 2
22 11 11 1 13 4 16 0 9 1 9 1 3 13 1 1 9 1 0 9 13 4 2
63 9 1 12 9 1 10 9 1 0 9 1 13 15 9 1 9 13 1 12 9 1 9 13 4 13 4 16 12 9 1 10 9 1 0 9 1 9 0 14 13 2 16 15 15 15 9 1 13 4 7 10 9 1 9 1 3 9 9 14 13 4 4 2
31 9 1 1 2 9 1 10 9 1 0 14 13 4 4 16 15 9 12 9 1 10 9 1 13 7 15 12 9 1 13 2
35 11 11 1 9 1 9 0 13 7 12 9 1 0 13 1 9 13 4 13 4 16 10 9 1 9 1 9 1 1 0 9 0 14 13 2
23 9 1 9 1 9 9 1 0 13 15 15 9 1 1 13 1 9 13 1 9 13 4 2
7 15 1 12 9 0 13 2
37 0 9 0 13 9 1 0 9 9 13 1 9 1 0 11 11 1 11 0 9 1 13 1 9 1 11 1 9 13 1 1 11 1 9 13 4 2
12 9 1 11 11 1 13 9 1 9 13 4 2
24 11 11 1 2 11 11 2 1 13 16 15 11 11 1 1 15 9 13 1 9 13 4 4 2
21 9 1 9 1 9 14 13 4 11 1 13 16 15 11 1 1 9 9 14 13 2
14 11 1 9 13 4 13 16 9 11 1 10 0 13 2
14 15 1 15 11 9 11 11 1 13 9 14 13 4 2
14 9 1 13 16 15 0 9 1 14 9 1 9 13 2
30 11 1 13 16 15 11 2 11 2 11 2 11 11 2 11 7 11 1 13 1 10 9 1 15 9 1 9 0 13 2
16 15 13 16 11 11 1 9 1 9 7 9 9 12 13 4 2
30 9 1 9 13 16 11 11 1 1 14 12 9 1 1 14 15 12 9 1 15 9 1 9 9 1 9 0 13 4 2
17 9 1 1 15 15 9 1 9 1 9 13 10 9 1 9 13 2
17 9 9 9 1 9 13 4 11 1 13 16 15 9 9 9 13 2
12 15 9 1 9 9 9 1 9 9 13 4 2
22 9 9 1 13 13 16 11 1 9 9 11 11 15 0 9 1 9 13 13 4 4 2
9 9 1 10 9 1 9 14 13 2
12 11 11 11 7 11 11 1 9 13 4 4 2
11 10 9 10 9 1 13 4 1 9 13 2
21 3 10 9 1 9 1 0 9 11 11 11 1 9 1 9 1 9 1 13 4 2
19 9 11 1 13 4 16 15 11 1 9 13 1 9 9 1 9 1 13 2
31 7 9 9 1 13 13 16 9 1 13 11 1 9 9 11 11 1 15 9 13 11 11 11 1 10 9 1 9 13 4 2
15 15 1 11 11 1 14 15 10 9 1 0 13 4 4 2
12 0 13 16 10 3 9 11 11 1 1 13 2
16 9 9 1 13 13 16 9 1 11 11 1 9 1 9 13 2
14 10 9 1 0 9 11 11 1 9 1 13 4 4 2
14 11 11 1 9 1 9 1 9 1 9 13 4 4 2
36 9 1 10 9 1 9 13 4 4 16 11 11 1 9 1 9 1 13 4 4 4 2 7 9 9 1 13 13 16 15 15 9 1 13 4 2
19 7 0 0 13 16 11 1 10 9 1 11 11 11 11 1 0 9 13 2
24 11 1 3 0 9 2 9 9 7 9 2 9 9 1 9 11 11 1 11 1 9 13 4 2
6 15 12 9 1 13 2
33 11 0 11 1 11 11 9 9 1 1 2 15 9 11 1 12 9 0 13 13 4 16 11 1 15 11 0 9 1 0 9 13 2
17 15 9 1 11 1 11 11 11 1 10 9 1 9 0 13 4 2
22 11 1 0 9 1 13 4 4 16 0 9 15 9 7 9 11 7 11 15 1 13 2
29 16 9 1 10 9 1 9 14 13 4 4 16 14 12 12 9 9 1 9 1 9 11 1 9 10 9 1 13 2
20 0 13 16 9 11 1 11 1 11 13 1 3 11 1 9 1 9 13 4 2
14 11 11 11 1 15 9 9 1 15 12 0 9 13 2
13 9 9 13 1 1 15 0 9 1 9 13 4 2
23 15 9 9 11 11 1 13 16 11 11 2 11 1 0 11 15 9 1 3 0 9 13 2
9 10 9 1 9 2 11 2 13 2
26 10 14 0 9 1 0 14 13 10 9 13 15 10 0 9 1 9 9 1 15 14 0 13 4 4 2
31 10 3 0 9 1 14 10 9 1 9 7 9 15 9 1 0 9 1 14 15 0 9 13 4 1 9 0 13 4 4 2
19 11 11 11 1 13 9 1 14 0 9 1 0 10 9 0 13 4 4 2
82 16 15 11 9 1 13 10 9 1 9 7 9 9 1 13 13 16 0 2 0 9 1 9 1 0 9 9 15 1 9 1 13 4 2 15 1 9 1 9 1 15 9 1 9 1 9 13 4 7 15 10 9 1 10 0 13 16 3 0 9 1 0 10 9 1 9 7 9 1 9 1 15 14 0 9 15 9 14 13 4 4 2
68 11 1 11 9 1 11 1 9 9 1 9 13 4 10 14 9 1 9 9 1 13 4 11 11 11 11 1 9 11 11 9 13 4 16 9 1 9 1 9 1 9 1 15 9 1 9 9 1 13 4 7 9 10 9 3 13 4 4 15 15 1 9 14 8 13 4 4 2
11 9 13 4 14 0 9 0 2 11 2 2
19 10 9 2 11 2 14 12 9 1 12 9 9 0 13 1 9 13 4 2
23 15 1 1 11 13 4 16 15 14 12 9 1 9 7 9 13 9 1 9 13 4 4 2
30 11 11 11 1 9 11 1 1 10 9 1 9 1 10 0 9 14 0 13 2 15 15 15 10 9 1 9 13 4 2
20 15 15 9 1 1 9 14 9 1 1 0 13 4 7 9 14 13 4 4 2
18 11 11 13 4 16 9 1 1 9 9 1 9 1 10 0 13 4 2
23 15 1 9 13 12 9 2 9 2 1 9 2 15 11 1 11 1 9 1 13 4 4 2
26 0 9 1 9 1 13 10 9 1 9 13 1 3 2 9 14 10 10 9 0 13 1 14 9 13 2
35 0 9 1 0 9 13 1 10 9 1 0 9 13 16 3 9 9 1 10 14 0 9 13 4 7 15 9 3 9 1 15 9 13 4 2
25 15 1 10 9 1 9 1 9 13 16 15 9 1 1 12 1 1 12 9 1 1 0 13 4 2
10 15 10 9 1 14 0 9 13 4 2
32 11 1 1 11 1 9 1 12 9 1 12 10 9 13 15 15 9 1 12 9 13 4 7 15 13 4 16 15 12 9 13 2
14 10 9 11 1 1 11 1 10 0 9 1 9 13 2
9 11 11 11 1 11 1 9 13 2
10 15 0 9 7 9 1 0 9 13 2
21 11 1 13 16 0 9 1 9 11 1 9 1 9 7 9 1 0 9 13 4 2
16 11 7 0 9 1 0 0 9 1 15 0 9 13 4 4 2
10 15 13 16 15 1 1 0 9 13 2
14 15 1 11 1 9 1 9 13 1 15 9 14 13 2
11 15 11 1 10 0 9 1 9 13 4 2
33 11 1 11 1 1 11 11 13 1 1 10 9 1 9 13 4 4 7 11 10 9 1 13 4 1 9 1 15 9 13 4 4 2
33 15 2 9 10 9 1 9 13 4 7 9 10 9 1 13 4 2 9 1 0 12 9 1 10 0 9 1 9 13 1 9 13 2
38 15 13 16 11 11 2 11 11 2 11 11 2 11 7 11 11 1 0 9 1 0 9 7 9 1 0 9 1 9 1 9 1 13 1 9 13 4 2
25 15 13 16 10 9 1 11 2 11 9 1 0 9 1 11 11 1 9 1 9 2 9 13 4 2
31 15 9 1 15 15 13 1 9 13 4 16 11 7 11 1 9 1 10 9 1 9 13 7 11 2 11 9 15 1 13 2
31 15 13 16 10 0 9 1 10 9 13 4 16 11 1 11 11 13 1 1 14 12 9 14 9 1 9 1 9 13 4 2
10 11 0 3 9 1 1 11 13 4 2
17 9 0 13 1 3 15 10 9 1 3 0 9 1 0 13 4 2
35 11 1 12 0 7 0 9 1 11 1 11 11 1 12 9 1 9 13 1 9 10 9 0 13 4 2 15 9 1 15 9 14 13 4 2
28 9 9 1 14 13 1 0 11 1 15 11 13 1 9 0 13 4 4 2 16 9 7 9 13 15 0 13 2
29 12 9 1 9 14 12 0 11 3 0 9 11 9 1 13 4 2 15 9 13 1 1 0 9 1 13 4 4 2
19 11 11 9 1 9 13 15 11 1 0 7 9 1 0 0 9 13 4 2
32 11 9 1 15 9 13 4 11 1 13 16 15 0 9 1 1 13 9 1 9 0 13 1 9 13 2 7 15 9 14 13 2
20 11 1 10 9 1 1 11 11 11 1 9 11 11 1 9 9 1 0 13 2
14 11 1 13 16 16 0 9 1 11 1 10 9 13 2
8 7 9 1 1 15 0 13 2
29 0 13 16 9 1 0 7 0 9 1 9 1 1 13 4 0 9 1 1 15 11 11 1 10 9 9 13 4 2
28 9 2 9 7 9 9 1 9 14 9 13 4 2 7 11 1 9 1 9 9 1 9 10 13 4 4 4 2
15 0 11 9 1 10 9 12 9 1 1 12 9 1 13 2
26 9 13 1 9 1 13 1 10 9 9 1 9 3 0 13 2 15 9 1 9 7 9 14 0 13 2
36 3 2 15 1 9 13 1 9 9 13 4 4 7 3 14 15 11 11 1 0 9 1 0 9 1 13 1 3 0 9 1 0 13 4 4 2
30 0 13 16 0 11 11 11 11 1 0 9 11 1 15 9 13 4 16 9 9 1 0 9 1 9 9 0 13 4 2
16 10 9 1 9 13 16 9 9 1 9 1 9 10 13 4 2
23 15 1 15 0 13 4 16 9 1 13 9 13 1 9 1 14 9 1 9 9 13 4 2
19 15 9 13 1 9 1 12 9 1 9 13 4 9 15 9 9 13 4 2
19 11 11 1 9 13 16 9 9 1 14 9 9 1 1 1 9 13 4 2
27 0 9 1 15 9 15 13 16 12 1 1 12 9 1 9 9 13 7 15 1 9 7 9 14 0 13 2
24 10 9 1 0 13 1 3 10 0 9 9 1 10 9 1 9 3 13 1 9 13 4 4 2
20 9 1 9 15 13 4 4 16 11 11 2 11 11 1 10 9 1 13 4 2
24 7 11 11 1 10 9 1 9 13 7 9 9 1 9 10 13 1 9 1 9 9 13 4 2
28 9 1 13 13 16 15 9 9 1 13 4 16 11 1 9 9 0 13 1 9 10 0 9 1 13 4 4 2
24 11 1 9 1 1 10 9 1 9 1 9 9 13 4 4 7 9 14 0 13 4 4 4 2
13 9 1 12 9 1 9 13 9 9 9 0 13 2
12 9 9 1 9 1 9 7 9 14 0 13 2
18 11 1 9 9 9 9 11 11 11 1 13 13 16 10 9 0 13 2
12 11 11 1 9 13 1 9 9 13 4 4 2
20 0 9 1 10 9 9 1 13 4 7 9 12 9 1 9 9 0 13 4 2
25 11 11 11 1 11 1 11 11 2 11 11 1 9 13 4 1 0 9 1 9 1 13 4 4 2
34 0 11 11 11 1 9 1 1 11 1 9 1 9 13 4 16 11 1 1 0 9 9 1 9 1 9 9 1 0 14 13 4 4 2
13 15 15 14 0 13 16 10 14 9 9 9 13 2
20 11 11 11 1 11 1 1 0 9 9 1 11 1 9 1 9 1 9 13 2
19 15 13 16 10 9 11 1 9 9 1 9 1 13 4 13 4 4 4 2
22 15 13 16 9 7 0 9 9 1 15 2 15 1 0 13 1 9 1 9 0 13 2
22 15 15 14 0 13 4 16 0 9 1 1 13 1 9 1 1 10 9 9 13 4 2
14 15 15 10 15 1 1 1 10 9 13 0 14 13 2
33 11 1 13 16 9 7 0 9 1 0 2 0 13 1 9 9 9 1 1 13 2 15 0 0 9 9 9 1 9 13 4 4 2
40 9 1 2 9 2 1 9 13 4 15 11 1 9 13 16 11 11 1 13 9 1 1 15 2 10 9 2 13 4 2 15 15 1 0 14 13 4 4 4 2
15 11 9 1 1 0 9 1 9 14 10 9 1 12 13 2
46 11 1 0 9 0 9 9 1 9 0 13 4 13 16 0 9 1 15 10 0 9 9 1 0 9 1 1 1 13 4 15 11 9 1 13 4 15 15 0 9 9 1 12 9 13 2
41 15 13 16 15 14 10 9 9 1 9 1 13 2 15 9 15 0 9 1 9 13 14 7 9 9 9 9 1 0 13 14 9 9 9 1 1 1 13 4 4 2
50 0 13 16 11 1 10 9 10 9 1 13 4 2 15 11 11 1 11 1 12 0 11 9 9 13 4 4 7 10 9 1 0 11 11 11 11 11 7 0 11 11 11 11 1 1 9 13 4 4 2
15 0 9 9 1 9 1 9 15 11 11 1 13 4 4 2
21 11 11 11 11 11 11 1 9 1 10 9 1 13 11 11 11 1 9 13 4 2
25 11 10 9 1 15 9 1 9 1 0 9 1 15 9 14 13 1 9 13 1 9 13 4 4 2
21 7 15 1 14 11 11 11 1 10 9 1 13 9 1 9 1 9 0 13 4 2
24 9 1 9 1 1 11 11 1 0 9 9 1 9 1 9 1 11 1 1 9 1 9 13 2
18 10 9 13 11 11 11 1 11 1 14 10 9 1 0 13 4 4 2
13 7 11 10 9 1 0 9 1 9 13 4 4 2
12 1 11 11 2 10 9 1 10 9 0 13 2
16 11 11 11 11 11 11 11 1 9 1 15 15 9 14 13 2
30 11 11 1 9 1 1 1 13 9 1 9 1 15 13 16 15 9 9 1 0 13 13 4 2 15 15 14 13 4 2
8 7 15 10 15 9 14 13 2
22 9 1 1 1 13 4 9 1 9 15 15 13 4 13 4 16 9 1 15 14 13 2
30 11 1 11 1 11 11 1 10 9 1 15 13 4 9 13 4 16 10 9 1 0 9 1 0 9 1 0 9 13 2
13 9 1 9 1 1 13 9 1 11 10 0 13 2
12 16 2 15 0 9 9 1 9 1 13 4 2
24 9 1 0 9 1 9 13 9 15 0 13 4 16 11 1 15 9 1 14 15 9 14 13 2
19 15 2 11 1 0 9 1 0 9 1 9 1 9 13 1 9 13 4 2
15 7 11 11 11 11 11 1 15 9 1 10 9 13 4 2
26 11 1 13 13 1 3 0 9 9 1 9 1 9 2 9 7 0 9 1 14 13 1 9 13 4 2
34 11 9 7 11 1 9 11 1 11 1 11 11 11 7 11 2 11 11 1 9 1 1 15 9 1 13 16 15 9 0 13 4 4 2
18 15 15 0 9 1 9 13 16 15 9 1 9 13 7 3 9 13 2
14 11 1 13 16 11 1 11 9 1 9 13 4 4 2
15 13 4 4 16 11 1 9 13 1 15 0 13 4 4 2
6 15 9 13 4 4 2
33 11 7 15 9 1 1 11 1 9 1 13 13 4 4 9 1 1 1 15 13 16 10 9 3 10 9 1 9 1 1 13 4 2
14 15 13 16 11 11 1 12 9 1 9 13 4 4 2
17 15 0 12 9 1 10 0 13 4 4 4 7 15 9 3 13 2
20 11 1 11 11 1 9 13 4 11 1 13 16 15 11 1 0 9 13 4 2
11 15 15 14 15 13 15 1 9 14 13 2
21 10 9 1 11 1 11 1 0 9 1 13 1 15 9 11 1 9 1 0 13 2
16 10 9 1 11 11 1 9 11 11 11 1 14 0 13 4 2
26 9 9 11 1 1 12 9 1 13 9 1 13 4 1 1 12 9 13 4 7 12 9 0 13 4 2
19 12 9 1 9 0 13 4 4 2 15 11 11 11 1 9 13 4 4 2
24 9 1 1 9 15 13 2 15 9 9 1 9 13 4 7 9 12 9 0 9 1 13 4 2
8 9 1 10 12 9 0 13 2
18 10 9 11 1 11 1 13 4 4 7 11 1 15 9 13 4 4 2
24 12 9 1 11 1 0 9 1 9 13 4 4 7 9 1 0 9 1 1 9 13 4 4 2
8 9 1 1 9 0 13 4 2
34 0 12 9 1 11 1 0 9 12 1 12 2 12 9 1 13 1 1 0 0 11 9 1 9 1 9 1 9 13 9 13 4 4 2
29 0 9 1 1 9 14 10 9 1 13 16 15 15 9 0 9 1 13 4 7 15 15 1 13 1 9 13 4 2
14 15 1 11 1 9 0 9 11 11 1 13 4 4 2
20 9 1 9 1 11 1 13 1 9 11 1 9 1 1 9 1 14 13 4 2
21 9 10 0 0 9 1 13 1 9 1 15 1 13 4 11 1 0 13 13 4 2
33 0 12 9 1 11 1 0 9 12 1 12 2 12 9 1 13 1 1 11 1 9 1 9 1 9 1 9 13 9 13 4 4 2
15 7 10 9 10 0 14 13 16 15 1 3 13 4 4 2
45 10 9 1 13 4 9 1 9 13 4 4 16 9 1 1 14 9 1 9 0 9 1 13 4 7 11 1 1 12 9 3 15 15 1 3 13 7 9 9 13 1 9 13 4 2
31 11 11 1 9 13 1 12 0 11 11 1 13 16 11 11 1 13 9 1 1 11 11 1 11 0 9 1 13 4 4 2
14 10 9 15 1 9 12 1 12 9 1 13 4 4 2
16 15 1 11 1 3 10 9 11 11 11 1 9 13 4 4 2
15 10 9 15 1 9 12 1 12 9 1 9 13 4 4 2
21 15 13 16 12 9 11 1 9 8 10 13 4 4 16 15 1 9 14 13 4 2
26 15 13 9 1 9 13 4 13 16 10 9 11 11 11 11 13 7 3 15 11 7 11 1 9 13 2
24 11 13 1 16 3 10 9 11 1 15 1 13 4 16 3 15 0 11 9 11 11 14 13 2
29 9 1 13 1 3 15 9 1 9 1 11 13 1 3 14 15 11 9 1 1 15 1 13 1 1 13 4 4 2
14 12 9 14 15 11 1 9 1 9 14 0 13 4 2
23 9 1 15 9 13 14 9 1 15 1 14 10 9 11 1 0 9 1 13 1 9 13 2
19 7 3 12 9 3 11 11 1 9 11 1 9 9 13 1 1 13 4 2
25 0 9 1 9 1 11 1 11 1 0 9 1 9 13 1 3 11 1 0 9 1 9 13 4 2
24 0 9 1 9 1 13 4 9 1 0 9 1 12 9 1 0 9 1 9 13 1 9 13 2
29 11 1 0 11 11 11 11 1 0 9 1 1 12 9 1 11 1 0 11 11 11 1 9 9 0 0 9 13 2
15 9 9 1 14 12 9 1 11 11 1 1 0 13 4 2
19 3 2 11 7 11 1 0 9 9 1 11 1 9 13 1 9 13 4 2
40 0 9 1 9 9 1 11 1 11 1 0 9 1 9 0 13 1 3 11 1 0 9 1 9 1 12 9 1 15 9 1 11 13 9 7 9 1 9 13 2
16 10 9 1 11 1 15 9 1 13 16 15 12 0 9 13 2
14 15 13 13 16 15 9 9 1 9 13 1 0 13 2
29 9 1 0 9 1 9 13 4 15 0 9 1 11 7 9 1 1 9 13 4 9 1 0 14 13 1 9 13 2
8 15 13 16 9 15 1 13 2
16 11 1 13 16 15 12 9 3 0 9 1 9 13 4 4 2
23 10 9 1 11 1 13 16 15 15 13 15 15 0 13 16 15 9 13 1 1 0 13 2
15 15 13 16 15 11 1 9 1 13 0 13 4 9 13 2
24 0 9 1 0 12 9 1 0 10 9 1 11 11 7 11 11 11 2 11 1 1 13 4 2
15 11 2 11 1 13 16 15 9 9 1 9 13 13 4 2
31 0 9 1 9 9 1 9 9 1 9 11 11 1 11 1 11 13 1 9 13 4 13 16 11 12 9 9 13 4 4 2
16 11 1 11 11 11 11 1 0 9 1 1 11 1 9 13 2
32 11 1 11 1 9 9 9 2 9 1 0 13 1 3 11 1 9 13 7 15 0 9 1 14 15 9 13 15 0 13 4 2
9 11 0 9 11 1 11 1 13 2
33 3 2 11 1 11 11 11 11 1 10 9 1 9 13 4 13 16 15 9 11 1 0 9 1 10 0 9 13 1 1 0 13 2
41 11 11 11 2 11 2 9 9 1 9 1 13 1 9 1 0 9 1 1 11 11 11 11 11 9 12 9 3 10 9 9 1 9 7 9 1 9 13 4 4 2
15 15 9 1 9 1 15 11 11 1 15 9 1 0 13 2
51 11 11 1 11 1 9 7 9 1 1 9 13 4 9 1 1 0 11 11 11 11 11 11 11 1 10 9 1 0 13 4 4 1 9 13 15 1 10 9 9 1 9 13 12 12 9 13 4 4 4 2
17 15 1 1 11 11 11 1 0 9 1 9 14 13 4 4 4 2
19 9 1 1 15 9 9 1 1 1 15 0 9 11 11 11 1 13 4 2
27 3 14 13 4 4 4 16 9 9 1 9 7 9 1 1 9 1 1 10 9 0 9 1 0 13 4 2
14 0 9 9 13 0 9 0 13 1 9 13 4 4 2
25 9 1 14 2 6 15 9 1 9 2 2 9 1 13 15 14 9 1 9 1 9 13 4 4 2
30 12 9 1 1 10 9 1 9 11 2 11 11 1 0 9 2 0 9 1 9 7 9 1 9 1 1 9 13 4 2
48 7 9 9 11 1 1 1 9 14 13 1 10 9 1 13 1 11 1 0 9 7 9 0 11 1 9 11 11 1 11 11 1 12 9 0 13 10 9 9 1 15 0 9 2 9 13 4 2
45 9 9 0 13 9 1 2 11 11 11 2 9 1 10 9 1 13 9 1 9 1 9 7 15 9 1 3 11 11 1 9 1 0 13 1 1 14 9 0 13 1 9 13 4 2
25 11 11 1 9 9 9 11 11 11 7 9 11 11 11 1 9 9 1 0 9 11 11 1 13 2
27 3 11 1 11 2 11 9 1 1 0 9 7 9 1 3 9 9 1 12 9 0 13 1 9 13 4 2
33 10 9 1 1 9 1 9 11 11 1 9 11 1 10 0 9 2 6 15 9 1 9 2 10 9 1 13 4 9 2 13 4 2
16 11 11 1 14 15 0 13 4 7 9 13 4 11 11 1 2
10 15 1 10 9 1 15 9 14 13 2
12 10 9 1 9 1 9 11 11 1 13 4 2
58 9 1 15 14 13 4 16 9 11 2 9 9 11 11 7 9 11 11 1 1 15 9 13 4 16 10 9 1 9 7 9 1 10 9 13 1 9 9 1 0 13 9 2 9 7 0 9 1 3 11 11 1 9 1 0 13 4 2
23 14 12 9 9 13 1 9 1 15 10 9 1 0 9 1 12 9 9 13 0 13 4 2
47 16 15 1 15 0 9 14 13 7 9 1 0 13 9 1 10 9 0 13 16 2 10 9 1 9 1 9 1 13 1 9 1 10 9 9 1 0 13 9 1 9 7 9 1 1 9 13
35 9 2 9 1 9 13 4 16 15 1 9 9 11 11 1 11 0 11 11 11 1 14 10 9 1 13 4 7 11 11 1 9 13 4 2
15 7 15 1 0 9 7 9 1 3 1 9 14 0 13 2
25 9 9 1 11 11 7 11 11 1 9 1 9 1 1 1 9 0 13 1 9 1 9 13 4 2
44 11 9 1 11 11 1 9 1 1 11 1 0 9 1 9 13 4 1 9 1 1 9 1 9 11 11 1 13 16 15 1 1 14 10 9 9 9 1 9 0 13 4 4 2
28 9 1 9 1 11 1 13 16 9 9 1 3 14 13 4 1 9 15 1 9 1 9 1 9 13 4 4 2
28 15 13 16 11 9 7 11 11 9 1 15 9 1 1 14 15 1 7 15 9 1 9 0 13 4 4 4 2
24 11 1 9 7 11 11 11 1 9 9 11 1 11 1 11 11 1 0 9 1 9 13 4 2
9 15 11 11 1 15 9 13 4 2
14 10 9 1 9 1 11 1 9 1 14 9 13 4 2
20 11 11 1 13 16 10 9 1 11 2 11 7 11 11 11 1 9 13 4 2
23 15 13 16 15 10 9 1 0 9 1 9 13 1 1 11 7 11 9 1 9 13 4 2
19 11 1 13 16 15 9 13 16 12 9 9 1 9 13 1 15 9 13 2
20 10 9 1 9 1 9 13 1 1 15 9 11 11 11 1 12 9 11 13 2
13 10 9 1 15 9 1 12 2 12 0 9 13 2
18 11 1 13 16 15 9 1 9 1 11 9 1 15 0 9 14 13 2
28 11 1 11 1 11 13 11 1 9 9 11 11 1 9 13 7 9 1 9 7 9 1 3 13 1 9 13 2
22 9 1 1 13 12 9 1 9 1 15 1 7 15 9 1 13 9 1 14 9 13 2
33 11 7 11 9 9 1 9 1 0 0 9 1 9 12 9 1 13 12 13 1 9 1 9 2 11 2 1 11 1 9 13 4 2
40 11 11 11 11 1 9 1 11 1 11 7 11 9 9 1 9 7 9 1 1 0 9 1 0 0 9 9 1 12 9 9 1 9 1 14 0 9 13 4 2
26 11 11 11 11 1 10 14 10 12 9 9 12 9 1 1 9 1 0 11 11 11 1 0 13 4 2
8 7 0 9 9 1 14 13 2
24 11 1 11 11 11 11 11 11 2 11 11 11 11 11 11 7 11 11 11 11 11 0 13 2
34 11 1 11 1 9 1 1 13 1 11 11 11 11 2 11 2 1 11 1 11 2 11 2 11 2 11 2 1 9 1 9 13 4 2
11 15 11 7 11 1 11 11 1 13 4 2
60 11 11 11 11 7 11 11 11 11 1 9 1 11 1 15 13 16 9 9 11 11 1 9 1 11 1 12 9 1 0 9 1 9 11 11 11 11 11 2 11 2 7 9 9 2 9 7 9 2 1 13 0 9 1 9 1 1 0 13 2
25 11 1 13 16 10 9 1 14 12 12 9 12 9 1 12 9 14 9 1 9 1 9 13 4 2
7 10 9 1 9 0 13 2
30 11 1 13 16 10 9 1 1 9 1 12 14 9 1 13 4 7 15 9 1 13 7 13 1 14 15 9 14 13 2
12 15 13 16 0 9 1 1 15 10 0 13 2
16 0 9 7 9 13 1 9 1 9 1 14 15 10 0 13 2
26 15 13 16 15 1 11 1 9 1 12 12 10 9 13 15 0 9 1 12 12 12 9 14 9 13 2
15 15 13 16 15 11 11 11 11 1 9 1 9 13 4 2
15 10 9 9 7 9 9 9 1 9 1 14 3 0 13 2
19 0 9 1 13 16 11 1 11 1 11 1 15 12 9 14 0 13 4 2
14 15 1 11 1 11 11 1 0 9 14 13 4 4 2
32 11 1 9 9 11 11 1 9 13 16 11 1 11 11 11 0 13 4 1 10 9 1 0 13 4 4 9 1 9 13 4 2
22 11 11 1 12 12 1 10 9 7 0 9 1 9 9 9 1 9 1 13 4 4 2
20 9 1 9 1 9 1 0 10 9 1 9 12 12 9 0 9 13 4 4 2
14 10 9 1 9 1 14 9 13 14 15 9 1 13 2
15 0 9 1 9 13 1 11 11 11 7 11 0 3 13 2
21 9 1 13 9 13 1 10 0 9 7 9 1 0 9 14 9 13 1 1 13 2
11 9 1 10 9 1 9 14 0 14 13 2
14 7 2 15 0 9 0 9 7 9 1 13 4 4 2
19 9 1 12 12 1 10 0 9 10 9 9 1 9 1 9 13 4 4 2
14 10 9 1 9 13 4 4 15 9 1 9 0 13 2
18 0 9 1 9 13 1 10 9 0 0 9 1 3 14 13 4 4 2
11 0 9 1 9 13 1 11 0 3 13 2
14 11 1 9 13 4 9 1 9 12 12 1 10 13 2
6 15 1 10 9 13 2
9 15 1 10 9 7 9 9 13 2
27 9 9 1 14 9 1 1 3 1 1 9 1 9 1 9 9 1 9 1 0 9 9 1 9 1 13 2
14 10 9 1 9 1 12 1 1 12 1 9 0 13 2
10 9 9 1 9 14 3 0 14 13 2
11 10 9 1 13 15 14 9 1 9 13 2
19 16 9 9 1 9 1 9 13 1 9 13 1 15 9 14 0 13 4 2
34 9 9 1 1 3 1 10 9 1 9 1 0 10 9 9 13 2 9 13 1 1 9 9 1 10 9 13 1 1 10 9 13 4 2
18 9 9 1 9 1 10 0 9 1 9 1 12 2 8 9 0 13 2
26 0 9 15 13 16 9 1 9 2 9 1 9 1 13 1 0 11 9 1 9 1 14 10 9 13 2
18 16 15 1 10 9 1 9 1 0 9 9 1 15 9 1 13 4 2
31 2 11 11 2 1 13 4 9 1 9 1 0 14 10 9 0 9 14 15 13 15 9 1 0 9 9 14 13 4 4 2
9 3 0 9 9 7 9 1 13 2
13 15 1 9 1 9 9 1 9 1 13 4 4 2
32 9 1 1 10 9 14 3 13 16 9 9 7 9 9 1 12 0 9 9 13 1 3 14 0 9 1 9 1 13 4 4 2
22 0 9 15 13 16 10 9 10 0 7 0 0 9 1 9 1 14 9 13 4 4 2
16 12 11 9 1 9 1 9 1 11 1 12 9 13 4 4 2
35 9 7 11 11 1 0 9 1 1 3 11 11 11 1 11 11 1 11 1 11 2 11 1 1 11 1 12 9 9 13 1 9 13 4 2
32 9 9 3 9 9 13 1 9 13 4 4 2 3 11 11 1 15 13 1 9 1 9 1 1 9 13 1 9 13 4 4 2
23 0 9 1 9 1 11 11 11 1 11 11 2 11 2 1 10 9 9 1 9 1 13 2
27 11 11 11 11 11 1 13 4 16 15 13 1 9 1 11 1 11 11 11 2 11 2 1 0 13 4 2
27 11 11 11 11 2 11 2 1 9 1 15 0 9 13 2 15 15 11 11 11 1 9 13 4 4 4 2
35 15 1 11 9 1 9 1 11 2 11 1 1 11 1 12 9 9 9 1 1 12 9 11 11 9 13 1 1 11 1 9 13 4 4 2
29 15 1 11 11 1 15 13 4 12 9 9 1 9 1 0 13 4 4 16 15 12 12 9 0 13 1 0 13 2
31 9 1 11 11 1 10 9 13 16 10 9 1 9 13 4 1 0 9 9 9 1 14 9 1 9 13 1 9 13 4 2
16 0 12 9 9 9 1 0 9 1 1 1 0 13 4 4 2
40 11 1 9 1 1 12 9 15 14 13 4 3 13 16 9 11 2 11 1 1 10 9 1 1 0 0 9 1 9 1 9 1 13 4 12 9 13 4 4 2
10 15 13 1 9 1 9 14 13 4 2
14 10 9 1 9 14 13 4 7 15 9 13 4 4 2
39 9 1 10 9 13 4 16 9 11 2 11 1 1 11 1 0 9 1 9 1 9 12 12 13 7 12 9 1 9 13 1 11 1 12 12 1 9 13 2
17 7 2 0 9 1 9 1 9 13 1 1 0 9 12 12 13 2
14 10 9 12 9 9 1 9 10 13 12 12 13 4 2
23 11 1 0 9 9 1 10 9 1 0 13 1 3 10 9 1 12 12 9 10 13 4 2
20 11 1 9 15 11 1 9 9 13 15 9 9 1 9 10 0 9 1 13 2
38 11 1 9 11 11 11 1 9 1 9 1 13 16 3 14 15 9 12 9 9 9 1 13 2 7 15 14 9 1 12 9 1 10 9 9 14 13 2
11 15 10 9 13 16 11 9 9 14 13 2
24 11 11 1 11 1 0 9 1 11 1 3 0 9 9 11 1 9 9 1 1 9 13 4 2
19 9 7 11 1 9 1 9 1 1 11 11 1 0 11 11 1 13 4 2
23 11 11 11 1 9 1 13 4 16 11 9 1 10 9 1 11 1 9 13 4 4 4 2
31 11 11 1 12 9 1 1 15 1 9 9 9 11 11 11 1 9 13 7 15 3 11 1 9 11 11 1 13 4 4 2
18 9 1 13 16 15 1 11 1 0 9 11 11 1 13 4 4 4 2
14 11 1 9 13 16 15 11 9 1 9 13 4 4 2
15 7 15 13 2 15 15 1 13 4 9 1 0 14 13 2
13 11 1 0 13 16 15 9 10 0 7 0 13 2
20 15 13 2 15 15 1 11 1 9 11 1 9 2 9 1 1 13 4 4 2
12 15 9 13 16 11 3 14 15 9 13 4 2
55 0 13 16 12 9 1 14 11 1 11 11 11 1 13 11 11 1 1 9 9 13 1 9 0 13 4 2 7 11 1 15 1 10 9 14 13 4 4 16 9 1 11 1 9 7 9 1 0 9 1 14 9 13 4 2
38 11 1 11 11 11 1 11 11 1 11 1 9 9 1 1 13 4 9 1 9 13 4 13 16 15 9 1 0 9 1 0 9 1 9 13 4 4 2
35 0 13 16 12 9 1 14 11 11 1 11 1 12 0 9 9 11 11 11 11 11 2 11 2 1 3 9 9 1 9 1 9 13 4 2
33 11 1 11 9 1 11 9 1 0 9 1 0 9 1 9 1 13 1 9 1 12 9 3 9 1 9 11 9 1 1 13 4 2
40 10 9 1 9 1 13 4 11 1 3 9 9 1 9 13 2 3 11 11 11 1 11 1 11 7 11 9 1 15 1 1 12 9 1 1 9 9 13 4 2
18 11 1 12 0 9 7 11 1 9 1 14 0 9 1 9 13 4 2
7 9 1 11 1 9 13 2
21 15 13 16 9 1 1 12 9 9 1 9 13 15 1 12 1 15 13 4 4 2
19 15 13 16 9 9 1 9 1 10 9 0 13 16 15 15 9 14 13 2
12 15 9 1 1 9 1 10 9 9 13 4 2
12 12 9 1 1 12 1 9 13 4 4 4 2
9 15 12 1 0 9 1 13 4 2
12 9 11 1 12 9 1 13 9 1 13 4 2
9 15 1 9 1 15 9 14 13 2
25 3 11 1 0 11 1 13 4 16 11 1 0 9 1 9 1 15 0 9 15 9 14 13 4 2
22 11 9 11 11 1 13 16 11 11 11 1 15 1 1 9 9 1 9 9 13 4 2
23 11 1 9 9 11 11 1 13 16 11 11 11 9 1 1 9 0 13 9 13 4 4 2
32 11 1 11 11 11 11 1 9 13 16 11 1 11 11 11 2 11 2 9 1 15 9 1 13 1 1 9 1 11 9 13 2
19 15 1 11 1 12 9 7 11 9 1 9 1 9 0 9 1 9 13 2
23 10 9 1 15 9 13 10 9 11 11 1 11 1 13 1 9 1 1 14 3 13 4 2
23 3 11 11 1 9 11 11 11 1 9 1 11 9 1 9 11 11 11 1 9 0 13 2
40 9 1 9 13 4 16 11 9 1 9 0 9 1 13 9 10 9 1 13 2 15 9 11 1 11 1 1 9 1 1 11 9 1 13 9 1 9 13 4 2
21 10 9 1 12 0 9 2 11 11 11 11 11 2 9 1 11 1 0 13 4 2
29 10 9 1 0 9 1 9 13 4 4 16 9 1 9 1 3 8 13 11 9 1 1 11 1 11 11 13 4 2
21 8 13 1 9 9 9 1 9 1 1 13 7 15 9 1 9 7 9 13 4 2
39 9 1 9 13 4 4 16 9 1 9 1 1 9 14 13 4 2 15 10 9 1 9 13 16 9 1 9 13 1 3 15 0 9 1 9 14 13 4 2
23 9 1 9 1 9 1 1 1 9 13 4 4 4 7 3 15 0 9 1 13 4 4 2
47 9 1 9 13 4 4 16 11 11 2 11 1 11 11 1 9 1 0 9 1 0 11 1 12 9 1 13 1 9 13 4 4 2 7 0 9 1 10 14 10 12 9 1 9 13 4 2
33 11 1 11 11 11 1 11 1 11 11 11 11 1 9 13 11 7 11 1 9 1 0 9 1 12 0 9 9 13 1 9 13 2
39 11 1 1 10 9 1 9 1 1 11 1 9 1 13 16 0 9 1 9 1 9 1 13 4 15 11 7 11 1 1 14 9 1 0 9 9 13 4 2
29 11 1 13 16 10 9 1 0 9 0 7 0 9 1 0 13 4 4 7 15 0 9 1 9 0 13 4 4 2
6 15 10 9 13 4 2
12 15 13 16 11 1 15 9 1 9 13 4 2
36 11 1 1 9 1 9 9 13 4 11 1 13 16 15 11 1 12 9 0 0 9 1 9 1 1 12 12 9 1 0 9 1 9 13 4 2
21 15 13 16 10 9 11 11 11 1 9 1 13 4 16 0 9 1 9 13 4 2
25 11 1 13 16 15 11 1 1 0 9 13 4 7 11 11 1 15 9 1 10 9 1 13 4 2
18 11 11 1 9 1 0 9 1 9 1 9 1 14 9 13 4 4 2
34 16 10 9 1 11 1 9 1 9 9 1 13 4 11 2 11 2 11 1 12 9 1 1 1 15 9 1 9 13 1 9 13 4 2
34 11 1 11 9 1 11 9 1 0 9 1 13 4 1 9 1 1 11 1 11 11 11 11 1 15 9 1 9 13 1 9 13 4 2
43 11 1 13 16 15 14 10 9 13 4 16 11 11 1 0 9 1 10 9 1 9 13 1 1 9 13 13 4 7 15 15 1 10 9 1 15 9 9 0 14 13 4 2
38 15 13 4 1 16 15 11 1 9 13 1 9 1 9 13 4 4 11 1 13 16 15 10 9 1 9 14 13 4 4 16 15 12 0 9 1 13 2
22 11 1 11 13 1 9 1 1 1 13 4 1 15 13 16 15 1 15 9 14 13 2
26 9 1 9 11 1 0 9 1 12 14 9 1 12 9 1 9 13 7 9 1 13 9 13 4 4 2
24 9 1 12 9 9 1 9 13 1 0 13 4 2 15 0 9 1 11 1 0 13 4 4 2
13 9 1 12 9 7 12 9 1 12 9 0 13 2
11 9 1 1 1 10 9 14 13 4 4 2
11 9 1 9 1 12 0 9 0 13 4 2
13 9 1 9 1 11 1 11 9 0 9 0 13 2
17 9 1 9 1 13 1 13 9 1 10 9 1 0 9 0 13 2
11 11 9 1 9 1 9 0 13 4 4 2
12 9 1 9 1 9 1 1 11 13 4 4 2
26 0 9 1 1 11 1 11 1 11 9 14 12 7 12 9 1 1 12 9 1 0 0 12 9 13 2
10 15 9 1 9 1 14 9 13 4 2
9 9 1 15 1 14 9 13 4 2
12 9 1 11 1 9 1 13 9 13 13 4 2
4 11 0 13 2
22 9 1 11 1 0 13 7 14 3 13 3 13 2 10 9 1 13 9 13 4 4 2
15 9 1 13 13 16 15 9 9 9 13 1 3 14 13 2
14 9 1 11 1 9 1 9 13 9 1 3 13 4 2
11 15 15 9 13 4 7 15 9 13 4 2
17 3 9 1 11 1 9 1 12 9 13 7 9 1 14 9 13 2
18 11 15 1 9 1 13 4 9 1 9 1 13 12 9 1 13 4 2
7 9 15 13 13 13 4 2
29 9 1 9 1 10 9 1 15 9 13 15 3 1 9 1 9 1 13 4 9 1 9 1 9 13 13 9 13 2
15 9 1 9 13 0 3 11 1 9 11 9 1 1 13 2
15 11 1 9 1 13 7 15 9 1 0 13 0 13 4 2
19 3 15 9 1 13 9 1 1 0 13 2 15 11 0 9 1 13 4 2
20 11 1 9 1 13 16 11 14 15 13 14 15 9 1 13 4 7 13 4 2
13 9 1 14 1 14 0 9 1 9 0 13 4 2
14 15 1 9 1 11 1 9 1 14 11 1 9 13 2
14 9 1 1 11 9 9 14 12 9 1 9 1 13 2
22 9 1 9 9 7 9 9 9 9 1 14 13 4 2 15 1 9 1 9 13 4 2
21 10 9 1 13 9 1 0 9 9 13 4 4 7 15 9 13 1 0 14 13 2
11 9 15 13 2 15 9 14 13 4 4 2
14 9 10 9 1 0 9 1 9 13 9 13 4 4 2
26 3 9 1 9 1 9 1 13 1 13 11 9 14 12 9 9 1 9 1 14 10 9 1 9 13 2
11 9 9 1 9 1 1 9 1 9 13 2
23 11 2 11 11 11 11 1 11 1 11 9 11 11 1 9 1 11 1 0 9 13 4 2
22 9 1 13 13 16 11 1 10 9 1 9 1 9 1 9 1 9 0 13 4 4 2
30 11 11 1 12 9 1 9 1 13 4 16 9 1 9 16 9 9 1 1 13 4 16 2 11 1 9 3 0 13 4
28 11 9 11 11 1 11 1 9 1 9 1 13 16 9 11 11 1 10 9 1 9 1 9 1 9 13 4 2
15 11 1 10 9 10 9 13 4 15 9 9 1 0 13 2
14 3 2 15 9 1 9 1 9 1 1 1 13 4 2
17 3 2 10 9 1 9 13 9 1 9 13 1 9 13 4 4 2
11 11 11 1 10 9 1 0 9 13 4 2
23 11 1 13 16 11 1 1 10 9 1 9 1 1 14 11 1 0 9 1 9 13 4 2
10 15 9 1 0 9 0 13 4 4 2
18 11 9 1 13 16 15 11 1 11 1 10 9 1 9 13 1 13 2
24 11 1 9 13 4 16 11 1 3 9 14 13 2 15 1 1 9 1 0 9 13 4 4 2
12 0 9 1 0 9 1 13 15 0 14 13 2
14 16 0 9 1 10 10 9 1 11 11 1 9 13 2
36 9 9 15 12 12 7 15 10 1 9 1 9 15 13 4 15 13 7 13 1 9 14 11 11 1 0 9 1 0 13 4 9 1 13 13 2
13 15 9 1 9 9 1 9 1 0 9 13 4 2
26 10 9 1 9 1 10 9 1 9 13 1 9 9 9 1 13 4 7 15 10 9 13 4 4 4 2
18 15 9 13 4 7 10 9 1 9 9 11 11 1 9 9 1 13 2
17 11 1 9 9 11 11 1 0 13 4 9 9 1 1 9 13 2
24 11 11 1 3 1 10 9 13 4 4 16 12 12 7 15 10 1 9 13 1 9 13 4 2
11 14 12 9 1 10 9 0 13 4 4 2
18 15 1 9 1 9 2 9 1 11 11 1 9 0 14 13 4 4 2
20 11 11 1 12 9 3 0 9 1 9 2 9 1 9 13 9 13 4 4 2
26 9 9 9 11 11 11 1 13 16 9 14 1 11 11 1 1 1 9 9 1 9 0 13 4 4 2
29 15 15 13 4 4 16 12 12 7 15 10 9 1 9 1 9 15 13 4 15 9 7 13 1 0 9 13 13 2
18 10 9 1 9 9 1 1 9 7 9 2 9 1 0 9 13 4 2
12 10 9 9 9 11 11 1 9 9 1 13 2
29 9 9 11 11 1 13 13 16 15 1 11 11 1 14 9 13 1 9 13 4 7 15 15 9 13 4 4 4 2
9 15 3 9 1 0 13 4 4 2
9 9 9 9 1 13 1 9 13 2
10 14 10 9 1 13 9 14 13 4 2
15 10 9 1 11 1 10 9 9 9 1 0 13 4 4 2
6 10 9 0 13 4 2
36 15 13 16 15 1 11 11 1 11 11 1 12 12 7 15 10 1 9 1 2 15 9 13 4 15 9 11 11 1 0 9 9 1 13 4 2
7 10 9 13 4 4 4 2
13 15 11 1 0 12 9 1 9 10 13 0 13 2
23 9 9 13 1 0 9 1 9 11 1 0 11 11 7 11 1 1 0 9 8 13 4 2
17 7 11 1 9 1 0 9 7 11 12 9 12 9 14 9 13 2
25 9 1 12 9 1 13 4 4 16 0 7 0 9 1 11 1 11 1 9 13 1 12 9 13 2
30 15 1 9 1 12 10 0 9 13 4 15 1 12 7 15 10 1 0 9 1 9 1 12 9 1 0 9 9 13 2
28 11 11 11 1 9 1 13 4 10 9 1 12 9 1 0 9 9 9 1 9 1 12 9 1 1 0 13 2
21 15 1 10 9 1 1 11 1 11 1 10 0 0 0 9 12 9 14 9 13 2
11 15 1 0 12 9 9 9 1 1 13 2
35 11 11 11 1 1 1 0 9 1 9 1 15 11 11 11 14 14 13 7 15 11 1 1 11 11 1 1 1 9 1 9 3 13 4 2
36 11 1 11 11 1 10 9 13 1 9 13 4 16 16 9 1 0 9 1 9 0 13 4 16 11 1 9 1 0 9 1 1 3 13 4 2
19 11 1 11 1 1 12 12 12 9 1 10 1 0 9 1 9 13 4 2
21 15 1 11 1 0 9 1 0 9 1 1 14 0 9 13 1 9 13 4 4 2
25 11 11 11 11 11 7 11 11 11 11 11 11 11 11 1 1 9 1 9 1 9 13 4 4 2
12 9 1 9 9 1 11 1 0 9 13 4 2
23 15 13 4 16 9 9 0 7 0 9 3 13 1 1 9 1 9 1 9 13 4 4 2
26 9 11 2 11 1 9 1 0 9 1 1 1 9 1 9 1 12 9 1 9 1 9 13 4 4 2
23 15 1 9 1 9 1 0 13 1 1 11 11 1 12 12 9 0 9 1 9 13 4 2
19 15 9 1 11 11 1 9 0 13 1 11 1 9 1 14 9 13 4 2
21 15 13 16 10 9 9 9 1 3 0 9 13 7 15 15 0 9 13 4 4 2
18 11 11 1 11 11 11 1 14 9 1 9 1 0 9 13 4 4 2
31 10 9 1 9 1 9 13 4 16 0 9 1 9 13 4 7 15 9 1 0 9 1 13 1 1 9 9 13 0 13 2
31 15 13 16 16 9 1 10 3 0 9 1 3 9 13 1 1 0 9 14 13 16 9 1 9 1 9 0 13 4 4 2
25 11 1 9 9 1 0 9 1 9 13 4 13 16 9 9 7 0 9 1 1 0 9 0 13 2
14 15 13 16 0 9 9 1 0 13 15 9 13 4 2
31 9 0 13 1 0 9 1 14 0 13 4 7 9 1 9 1 0 9 1 0 9 1 9 1 13 1 1 0 13 4 2
13 15 9 13 1 9 1 9 1 14 0 9 13 2
24 15 9 9 1 0 13 1 1 9 1 12 9 9 9 1 1 1 0 13 1 14 9 13 2
18 11 11 1 9 13 16 9 1 9 1 9 1 9 1 9 13 4 2
22 11 9 1 9 1 0 9 0 13 4 11 2 11 2 11 1 9 1 9 13 4 2
17 10 9 1 1 11 1 12 9 13 4 7 12 0 13 4 4 2
21 10 9 1 11 11 11 1 11 7 0 9 1 10 0 9 1 9 1 9 13 2
29 12 0 9 9 1 13 16 11 11 1 11 1 10 12 9 9 9 1 13 4 4 15 9 14 10 9 1 13 2
35 11 2 11 1 9 9 11 11 1 9 1 13 16 10 9 1 11 1 11 11 7 11 2 11 7 11 1 0 9 1 9 1 9 13 2
14 15 1 15 9 1 10 9 7 0 9 9 14 13 2
30 11 9 1 0 9 9 1 9 13 4 16 10 9 1 9 11 1 11 11 1 9 1 13 4 12 9 1 14 13 2
20 11 11 1 13 16 11 1 13 4 9 11 2 9 1 14 15 13 4 4 2
17 15 13 16 10 9 0 13 1 1 15 9 1 9 13 4 4 2
22 11 11 1 13 16 10 9 1 0 12 9 1 1 11 1 0 9 1 13 4 4 2
11 10 9 10 0 9 1 9 1 0 13 2
18 10 9 1 11 9 11 11 11 1 9 9 11 11 1 9 13 4 2
12 15 1 15 10 9 7 0 9 1 0 13 2
14 11 1 13 16 11 9 1 12 9 0 13 4 4 2
21 15 1 11 9 11 9 1 9 1 9 9 1 9 1 1 12 0 9 13 4 2
10 10 9 1 12 9 14 0 13 4 2
17 9 1 9 13 1 13 4 7 15 9 1 9 13 9 13 4 2
18 9 1 0 9 1 12 9 13 4 7 0 9 1 9 13 13 4 2
14 13 4 9 1 9 11 11 1 1 1 13 4 4 2
17 9 1 12 9 9 9 2 12 9 9 7 9 0 13 4 4 2
38 11 0 9 1 9 1 9 1 9 1 15 1 15 9 3 14 13 4 7 10 9 1 13 12 0 9 1 9 12 2 12 9 1 13 1 9 13 2
19 10 9 9 1 9 7 9 9 1 14 10 9 1 0 13 4 4 4 2
15 9 7 9 9 1 9 13 1 3 15 1 9 13 4 2
22 11 9 11 11 2 9 11 11 7 11 11 1 0 9 11 11 10 9 1 9 13 2
31 9 0 12 2 12 9 1 14 9 7 9 1 9 1 13 10 9 13 1 13 4 4 15 1 9 1 9 13 4 4 2
32 10 9 1 0 9 1 14 15 1 9 14 0 13 0 13 4 4 2 16 10 9 0 9 1 9 1 9 13 4 4 4 2
15 9 1 9 9 1 13 4 9 1 1 0 13 4 4 2
15 10 9 1 11 1 0 9 1 14 9 1 9 13 4 2
13 10 9 1 15 15 9 1 13 10 0 13 4 2
27 9 9 1 10 9 1 9 1 11 1 9 13 4 2 10 9 1 14 13 4 1 9 13 4 4 4 2
8 10 9 1 14 0 9 13 2
35 11 1 9 13 15 14 12 9 1 9 13 16 16 9 1 12 2 12 9 9 9 1 11 3 13 4 16 0 3 11 1 13 4 4 2
14 9 3 15 14 11 1 13 4 1 9 1 14 13 2
23 11 1 13 4 9 1 1 15 1 9 13 1 1 9 9 1 14 9 13 4 4 4 2
20 10 9 1 9 9 1 0 9 13 0 13 4 1 9 14 13 4 4 4 2
45 10 9 1 14 11 3 14 11 9 11 11 1 9 1 13 7 10 9 1 9 13 16 10 9 1 1 15 15 0 9 1 1 14 13 4 4 2 15 3 9 13 4 4 4 2
13 9 1 3 0 9 1 11 1 0 9 13 4 2
22 11 1 0 0 9 9 9 1 3 0 9 0 9 11 1 3 0 9 13 4 4 2
15 11 9 2 11 2 1 9 13 1 10 9 1 9 13 2
9 11 14 11 1 10 3 14 13 2
18 12 1 12 1 9 1 11 1 10 9 12 9 0 13 0 9 13 2
12 16 9 1 9 1 11 1 10 9 13 4 2
8 9 11 1 10 9 12 13 2
23 10 9 1 11 1 3 13 1 9 14 11 2 11 2 11 2 11 2 11 7 11 13 2
24 10 9 1 11 1 0 9 1 9 7 15 0 9 1 13 4 9 1 9 9 13 4 4 2
14 11 1 9 1 1 9 1 12 12 9 1 9 13 2
14 0 11 1 9 1 12 12 9 9 1 9 13 4 2
11 7 0 9 1 9 1 8 13 4 4 2
9 11 10 9 1 3 10 0 13 2
13 15 3 10 9 12 13 4 7 9 9 13 12 2
29 11 1 15 9 0 13 4 11 1 9 9 2 0 0 2 11 11 11 1 13 16 0 9 1 9 3 10 13 2
16 7 11 2 11 7 11 1 0 9 1 1 15 9 10 13 2
13 11 1 12 9 1 1 3 10 0 9 13 4 2
19 7 11 1 15 10 14 0 9 13 12 9 1 1 12 9 0 13 4 2
21 9 1 1 9 1 9 1 0 9 11 1 0 9 0 13 12 9 0 13 4 2
11 7 15 12 9 1 1 0 9 1 13 2
26 2 11 11 2 1 9 13 1 3 9 9 11 11 15 3 14 15 0 9 1 0 13 1 0 13 2
19 7 14 15 9 1 1 9 13 2 0 9 2 1 9 14 14 0 13 2
14 10 9 1 9 1 9 9 1 1 9 3 0 13 2
14 15 1 11 1 12 9 1 9 1 13 1 9 13 2
33 15 1 14 9 1 0 9 9 1 15 13 1 0 9 13 4 4 16 2 11 11 2 1 13 9 1 0 2 0 0 13 4 2
19 11 1 9 9 9 11 11 1 13 2 2 15 12 0 9 1 9 13 2
16 10 9 3 0 13 4 4 7 10 9 15 1 0 14 13 4
39 16 2 0 9 9 11 1 13 16 15 11 1 13 1 1 1 0 9 1 15 9 13 1 9 1 14 13 16 0 10 9 1 15 11 1 14 13 4 2
15 11 1 13 2 2 15 11 13 4 7 15 15 9 13 4
19 7 15 13 16 10 9 1 9 8 13 4 1 3 11 1 9 0 13 2
25 9 11 1 13 2 2 15 13 4 4 16 15 9 1 1 0 9 1 10 9 1 13 4 4 2
31 11 1 10 9 1 9 13 1 0 13 1 9 1 11 1 13 2 2 11 1 14 9 13 15 1 15 1 9 13 0 13
28 0 9 1 3 0 13 1 9 1 1 1 9 1 9 9 1 13 2 2 10 9 0 11 1 9 1 13 2
16 9 9 3 0 13 4 16 9 1 9 7 9 1 9 13 4
35 0 9 1 10 0 13 1 9 13 4 11 1 13 2 2 9 1 9 2 9 1 9 1 9 13 4 7 11 1 10 9 14 13 4 4
32 11 11 1 9 7 0 9 1 9 1 1 12 9 9 1 9 1 9 1 11 11 11 1 11 11 1 1 1 13 4 4 2
22 9 13 1 9 1 9 1 9 13 1 9 1 11 1 9 1 15 9 14 13 4 2
36 9 11 11 11 2 9 11 11 2 9 11 11 2 9 11 11 11 7 9 11 11 11 1 0 9 1 9 1 11 11 1 1 1 13 4 2
64 0 9 11 11 2 11 2 11 2 11 11 1 9 11 11 2 11 1 0 9 11 11 7 11 1 11 11 11 1 13 16 15 9 1 1 15 9 13 16 9 1 12 9 0 9 0 2 0 7 0 9 1 13 4 4 7 0 9 1 15 9 0 13 2
37 11 1 13 16 2 16 15 0 9 1 0 9 1 15 9 1 9 13 4 4 16 3 0 9 2 9 2 1 15 9 1 10 9 15 14 13 4
38 15 15 14 13 16 9 1 9 1 14 0 9 1 13 1 1 14 9 13 1 9 14 13 2 16 15 14 14 15 0 9 1 12 3 0 9 13 2
40 11 1 13 16 9 13 1 1 9 1 9 9 1 9 1 1 9 13 4 9 1 0 13 7 9 1 0 9 1 1 0 11 11 11 1 9 0 14 13 2
33 16 2 9 9 1 1 1 9 1 0 13 9 11 11 11 11 1 13 16 2 9 9 9 2 1 9 1 1 0 13 4 4 2
16 10 9 1 9 1 9 1 9 1 9 13 1 9 13 4 2
23 11 7 11 11 11 1 0 9 11 11 11 1 9 13 4 16 9 9 1 1 9 13 2
19 15 13 16 9 1 10 9 1 0 7 0 9 1 0 9 1 9 13 2
20 12 9 9 1 9 9 11 11 1 9 1 11 1 1 1 9 13 4 4 2
19 12 9 7 9 1 9 1 9 1 9 1 9 1 9 1 10 9 13 2
17 11 1 0 9 1 9 1 11 1 14 9 1 9 1 9 13 2
14 16 11 1 15 1 9 13 15 11 1 14 0 13 2
20 15 1 9 1 11 1 11 1 1 1 0 14 13 1 9 1 9 13 4 2
37 11 1 15 1 13 4 9 7 9 1 13 1 9 13 1 9 1 0 13 4 13 4 16 15 9 1 9 0 13 1 1 9 13 1 9 13 2
26 7 9 1 9 13 16 11 1 15 9 1 13 7 15 9 13 1 9 13 12 9 15 0 9 13 2
41 9 9 13 1 3 11 2 11 1 0 9 1 15 0 9 1 11 1 11 11 11 11 1 13 16 11 1 10 9 1 0 13 1 1 0 9 1 9 13 4 2
17 15 11 2 11 9 1 9 1 9 1 9 1 14 0 9 13 2
13 15 13 16 9 9 1 9 1 15 9 14 13 2
42 11 11 11 11 1 9 1 9 1 9 13 4 13 16 11 1 9 9 13 1 1 10 9 3 14 13 16 15 15 9 1 9 1 1 1 15 0 9 1 9 13 2
24 11 2 11 7 11 2 11 9 13 4 1 9 1 15 13 16 9 1 9 1 9 14 13 2
24 9 9 1 9 1 1 1 13 4 1 15 11 11 1 13 1 0 9 1 9 13 1 13 2
26 15 1 15 9 1 9 1 0 13 4 13 16 11 1 9 9 1 11 1 0 9 1 9 13 4 2
22 11 11 2 11 1 9 1 9 2 9 7 9 1 10 9 1 9 1 1 0 13 2
25 15 9 1 9 9 13 4 15 13 16 9 9 1 0 9 1 13 1 1 10 0 9 13 4 2
13 15 13 16 9 9 1 9 1 9 0 13 4 2
16 11 11 1 9 1 0 0 9 1 1 2 0 9 2 13 2
29 9 9 11 11 11 7 0 0 9 1 15 9 9 1 9 7 9 13 1 1 13 4 9 1 1 1 9 13 2
20 0 9 1 9 1 11 11 11 11 11 11 1 9 9 1 9 13 4 4 2
19 10 9 1 0 9 11 1 11 2 11 11 1 13 1 9 1 13 4 2
19 11 1 9 1 10 9 1 11 11 2 11 2 9 11 11 14 0 13 2
12 9 1 11 1 0 9 1 0 9 0 13 2
33 15 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 11 2 11 11 2 11 11 7 11 11 0 13 2
22 7 10 0 9 1 9 13 16 16 9 14 13 4 16 9 1 15 0 9 13 4 2
22 11 9 11 11 1 13 13 16 0 9 1 9 1 9 1 13 1 9 0 13 4 2
16 15 13 13 16 15 10 9 1 15 0 9 14 13 4 4 2
11 11 1 9 1 15 1 0 9 13 4 2
14 0 9 1 9 1 3 0 9 11 11 11 1 13 2
23 9 1 10 9 1 14 9 13 7 9 9 1 11 7 11 1 1 13 9 1 9 13 2
28 9 1 0 13 16 9 9 1 13 4 1 9 1 9 9 1 13 2 7 15 1 15 9 1 9 14 13 2
20 11 9 11 11 1 11 1 11 11 11 1 13 4 1 9 1 0 9 13 2
12 15 13 13 16 11 1 13 4 9 0 13 2
15 15 13 16 9 1 9 1 13 4 1 9 0 13 4 2
10 0 9 11 1 8 13 2 13 4 2
25 11 2 11 11 11 11 11 11 1 13 9 1 1 11 7 11 9 1 0 9 3 0 13 4 2
17 9 11 1 0 9 1 9 0 13 3 2 3 9 1 13 4 2
13 9 15 13 4 16 9 1 9 12 1 13 4 2
22 3 1 3 2 3 12 12 9 9 1 9 13 9 9 7 0 9 1 9 13 4 2
11 0 11 1 12 9 1 3 9 13 4 2
28 11 11 1 9 1 9 13 13 9 9 1 11 11 11 11 1 3 9 1 9 13 9 1 0 9 13 4 2
10 9 0 9 13 4 15 12 9 13 2
22 9 12 9 1 9 12 9 1 14 9 14 13 16 11 11 1 9 13 9 13 4 2
32 15 9 13 16 9 14 12 9 11 2 11 11 11 11 11 11 1 11 9 1 9 9 1 9 13 1 10 9 0 13 4 2
11 10 9 1 12 9 9 3 1 0 13 2
23 11 2 11 1 1 14 12 9 9 1 11 2 11 7 11 2 11 9 14 8 13 4 2
8 15 9 9 0 9 13 4 2
23 10 9 9 13 2 10 9 9 1 14 12 9 9 13 4 4 15 3 12 1 13 4 2
22 9 9 13 4 16 9 1 14 12 12 9 14 9 13 4 15 14 12 1 9 13 2
22 9 1 3 12 9 1 9 13 1 9 1 9 12 9 1 13 4 15 12 13 4 2
11 11 11 0 9 1 9 2 9 13 4 2
21 11 1 11 11 7 11 9 9 1 13 0 9 1 9 1 0 9 13 4 4 2
15 11 7 11 1 0 9 1 9 1 9 1 9 0 13 2
10 9 9 9 12 12 9 1 0 13 2
28 9 1 13 4 9 12 12 9 1 9 1 12 12 9 1 9 1 9 1 1 9 1 9 0 13 4 4 2
51 9 1 11 1 12 9 1 12 7 11 1 12 9 1 12 9 9 1 0 14 13 4 4 7 0 9 1 1 11 1 12 9 9 1 12 9 7 12 9 9 1 12 9 9 1 3 13 0 14 13 2
19 15 1 1 0 12 2 12 9 1 9 1 9 9 3 13 1 9 13 2
35 11 11 11 2 11 2 1 11 1 11 11 1 0 9 9 11 11 11 1 0 9 1 9 1 9 13 1 1 12 9 1 9 13 4 2
13 11 1 15 9 1 11 11 11 1 9 13 4 2
12 15 1 1 9 9 1 15 9 13 4 4 2
13 9 9 1 9 1 9 13 1 1 9 13 4 2
14 15 1 11 1 9 1 0 9 11 11 0 13 4 2
12 9 9 1 11 1 0 9 1 9 13 4 2
14 15 15 9 11 11 1 11 11 11 1 9 13 4 2
20 9 9 1 11 1 1 0 9 0 13 1 1 15 3 12 9 9 13 4 2
38 7 9 9 1 0 9 9 1 0 14 13 1 15 9 1 11 1 1 0 12 9 1 11 1 0 9 0 13 1 9 1 0 13 1 9 13 4 2
37 11 1 9 1 13 13 15 11 11 1 3 12 9 0 13 1 0 0 9 1 9 14 13 2 15 10 9 10 9 10 0 15 13 4 4 4 2
35 11 1 11 11 1 0 9 1 1 12 9 9 9 13 4 7 11 11 1 11 1 9 0 13 1 9 14 13 1 9 0 13 4 4 2
60 11 1 1 1 9 1 0 9 1 11 11 11 1 9 11 1 11 1 1 9 14 13 1 9 1 9 13 4 7 9 13 4 16 11 11 1 1 9 13 1 9 9 1 13 1 14 13 1 1 1 11 11 11 1 15 9 13 4 4 2
28 11 11 2 11 2 1 13 4 16 11 1 10 9 1 9 13 1 1 12 9 1 9 1 15 9 14 13 2
13 9 1 13 13 16 12 9 1 1 0 9 13 2
35 11 11 2 11 2 0 9 1 9 11 11 1 11 1 13 16 15 1 0 13 9 1 10 9 14 13 16 15 11 1 0 13 4 4 2
51 11 11 0 0 0 9 9 1 9 9 2 9 9 7 0 9 1 0 9 1 9 1 1 9 9 7 9 1 0 9 1 9 1 13 12 9 1 1 0 13 9 1 9 1 9 1 9 13 4 4 2
16 0 9 1 9 1 15 13 16 11 15 1 9 13 13 4 2
13 7 9 1 9 1 13 10 9 1 1 9 13 2
23 11 1 9 13 16 10 12 9 1 11 7 11 11 2 11 2 1 9 0 2 0 13 2
21 15 13 16 11 11 2 11 2 11 1 11 1 9 1 11 9 1 12 9 13 2
54 15 9 1 11 11 1 10 9 1 15 9 13 13 15 15 13 4 16 11 9 1 9 1 14 11 1 9 0 13 15 11 1 13 16 11 1 9 13 16 9 1 9 7 9 1 1 10 9 1 9 13 4 4 2
30 11 1 11 1 11 11 11 1 9 1 9 1 13 4 12 9 1 9 1 11 1 13 16 15 11 1 0 9 13 2
24 11 1 0 9 11 11 1 11 1 11 1 0 9 11 11 11 7 11 11 11 1 9 13 2
17 9 1 1 15 13 16 15 11 7 11 1 9 13 15 13 4 2
21 11 1 15 0 9 7 11 1 0 9 11 11 1 9 1 1 9 13 4 4 2
16 11 1 11 11 11 1 0 9 15 11 7 11 1 9 13 2
18 0 0 9 0 13 1 3 11 0 9 1 0 9 9 13 4 4 2
19 15 13 16 11 7 11 1 9 1 0 9 1 9 1 15 9 14 13 2
21 15 13 16 12 0 9 13 7 15 1 9 0 13 1 1 15 15 9 13 4 2
18 9 1 1 11 1 1 15 9 1 9 1 9 13 1 15 9 13 2
42 15 13 4 1 16 15 15 11 1 9 11 9 11 11 11 1 11 9 1 13 9 1 0 9 1 9 13 1 15 9 13 4 2 15 15 9 13 1 9 13 4 2
15 15 9 1 15 10 9 1 9 1 14 13 1 1 13 2
34 11 11 1 9 11 11 1 11 1 13 16 16 11 9 11 11 1 9 1 9 1 13 4 9 9 13 16 15 3 9 14 13 4 2
30 9 14 1 11 11 11 1 13 0 9 1 1 11 1 9 1 9 7 11 11 11 1 9 9 1 9 13 4 4 2
41 15 11 11 11 1 0 9 1 0 13 4 11 1 13 16 11 1 15 14 10 9 1 9 13 4 1 9 13 4 2 15 1 11 11 11 1 13 1 9 13 2
12 15 13 16 11 15 9 1 9 13 4 4 2
18 15 13 16 9 1 9 1 0 0 13 4 1 9 1 15 9 13 2
36 15 13 16 11 1 9 13 4 2 16 15 9 1 11 11 1 9 1 0 9 11 11 1 11 11 11 1 13 1 13 0 9 0 13 4 2
29 15 1 1 0 9 1 9 13 4 11 11 1 9 11 11 1 9 1 13 16 15 11 1 9 14 13 4 4 2
15 15 13 16 15 14 11 1 1 9 11 11 1 13 4 2
17 11 1 11 1 11 9 11 11 12 9 3 9 1 13 4 4 2
18 12 0 9 1 0 9 1 15 1 0 2 0 9 0 13 4 4 2
24 9 9 11 11 1 11 1 13 16 9 1 11 9 1 1 0 9 9 1 12 9 13 4 2
7 15 3 14 9 13 4 2
30 0 9 1 1 9 1 1 9 1 9 9 1 9 2 11 9 9 7 0 9 1 0 9 9 1 13 4 4 4 2
46 11 9 1 12 9 11 11 7 11 11 1 9 9 1 10 9 13 4 1 1 9 1 1 0 14 13 1 9 9 9 9 11 11 11 1 11 1 9 11 1 1 9 0 13 4 2
11 0 9 1 9 1 12 0 9 0 13 2
23 11 2 11 1 3 0 9 1 9 11 11 11 1 11 1 11 9 1 0 13 4 4 2
30 11 1 0 9 10 9 1 9 1 11 7 11 1 0 9 1 9 9 13 1 9 1 12 12 9 1 9 0 13 2
17 11 2 11 9 1 13 4 1 9 0 11 11 11 1 13 4 2
31 11 11 1 1 1 12 0 9 1 0 9 1 1 10 0 9 1 0 11 1 12 9 1 9 1 1 0 13 4 4 2
24 10 9 1 9 1 0 9 7 15 9 1 0 9 1 1 12 0 0 9 14 13 4 4 2
12 10 9 1 1 12 9 1 0 13 4 4 2
37 11 11 1 13 4 9 1 9 14 13 7 2 11 11 11 2 0 9 1 12 9 1 1 1 13 4 16 15 0 15 14 0 11 11 11 13 2
19 11 11 1 11 7 11 1 0 9 1 13 4 9 9 9 1 0 13 2
9 10 9 1 10 9 13 4 4 2
33 0 11 11 11 11 1 13 4 9 1 9 11 1 1 1 13 4 7 13 4 16 15 0 9 1 1 9 1 12 0 9 13 2
23 11 1 13 16 15 9 13 15 9 13 4 16 11 1 15 9 10 10 9 1 13 4 2
15 15 13 16 11 1 0 9 9 1 1 14 11 13 4 2
29 11 0 9 9 11 1 3 0 9 1 1 13 7 0 9 1 15 9 1 12 12 9 1 9 0 13 4 4 2
23 11 11 11 1 13 4 11 11 11 1 1 11 1 13 4 1 0 0 11 11 9 13 2
28 11 1 9 12 9 1 10 10 13 7 15 2 9 2 7 2 11 11 11 2 1 9 1 14 13 4 4 2
37 11 11 1 9 1 11 13 4 10 12 9 11 9 10 9 3 2 3 13 4 15 9 13 9 1 1 13 4 7 15 9 9 9 1 13 4 2
29 11 9 1 10 9 1 1 9 1 15 0 13 4 4 7 15 13 1 10 9 1 11 1 13 1 1 13 4 2
18 9 1 1 9 1 12 9 1 0 13 1 3 11 1 13 4 4 2
17 10 9 11 1 9 12 9 10 9 13 15 0 9 13 4 4 2
10 11 11 2 11 9 11 1 13 4 2
20 11 1 15 10 9 1 0 13 4 7 15 9 2 9 2 14 13 4 4 2
38 11 11 11 11 11 11 1 11 1 13 16 0 9 1 13 4 4 16 0 9 1 9 9 1 13 1 13 1 1 9 1 0 9 1 9 14 13 2
18 15 13 16 9 1 9 13 16 9 0 13 1 3 9 9 13 4 2
18 15 13 7 9 9 1 9 9 9 1 10 9 1 9 1 13 4 2
33 16 2 9 1 3 9 1 13 4 7 15 12 0 9 11 11 2 11 1 9 12 13 12 9 1 11 1 1 0 13 4 4 2
11 11 11 1 9 11 11 1 10 9 13 2
22 7 9 1 9 9 1 12 9 1 1 14 15 1 13 9 1 0 13 4 4 4 2
16 12 14 9 11 11 1 9 1 12 9 9 1 9 13 4 2
25 10 9 1 0 12 9 1 3 9 1 8 13 2 3 0 9 1 13 9 14 0 13 4 4 2
13 9 1 1 11 11 1 9 13 1 9 14 13 2
10 10 9 9 9 1 1 14 13 4 2
25 11 1 0 9 1 10 9 9 13 4 2 15 9 1 0 13 4 12 9 9 1 0 13 4 2
21 15 14 1 0 9 1 9 1 13 13 1 12 9 1 11 11 13 1 0 13 2
16 0 9 1 9 13 4 16 10 9 1 0 9 13 4 4 2
36 0 9 9 11 1 1 12 0 9 1 9 1 9 1 1 11 11 11 7 0 11 11 11 2 11 2 1 9 11 11 9 1 0 14 13 2
19 0 9 9 11 11 11 11 11 1 10 9 1 1 9 1 8 13 4 2
38 0 11 11 11 1 11 1 13 16 11 1 11 11 2 11 2 1 0 9 7 9 1 0 13 1 3 1 11 1 9 1 0 0 9 13 4 4 2
26 15 13 16 15 11 10 9 1 9 1 1 15 15 9 9 15 13 15 10 9 15 0 9 1 13 2
49 11 1 9 13 4 11 1 11 1 10 9 1 9 1 9 13 1 1 11 1 13 1 9 9 7 14 11 1 1 11 11 1 9 1 0 9 13 1 1 10 9 2 9 13 1 9 13 4 2
22 11 11 11 1 1 11 1 13 1 9 9 1 10 9 0 9 2 9 13 4 4 2
25 11 1 1 13 1 11 11 1 9 1 9 1 13 4 9 9 1 9 1 0 13 1 9 13 2
39 11 1 12 9 9 1 10 0 9 1 0 13 1 12 9 1 11 11 0 11 11 1 11 11 1 13 16 15 9 13 4 16 11 10 9 1 9 13 2
33 15 14 10 0 9 15 11 1 9 1 13 15 13 4 16 0 9 1 9 15 13 7 9 7 0 9 1 9 0 9 15 13 2
21 11 15 9 1 0 9 13 1 1 3 14 11 1 0 9 7 9 13 4 4 2
22 3 14 0 11 11 1 12 9 10 9 1 9 1 9 1 11 1 9 13 4 4 2
29 9 9 9 1 12 0 9 1 15 9 0 13 1 9 1 13 16 11 11 9 1 12 9 11 0 13 4 4 2
17 11 1 11 11 0 11 11 11 1 10 0 9 1 9 13 4 2
20 9 1 13 16 0 7 0 9 1 9 1 9 1 9 13 3 0 13 4 2
20 0 13 16 11 9 13 1 1 11 11 11 1 0 9 1 9 13 4 4 2
18 0 9 1 9 10 9 1 9 1 14 9 1 0 9 1 9 13 2
17 12 9 0 11 2 11 11 1 0 9 1 9 14 13 4 4 2
15 15 1 9 1 1 0 9 1 9 13 0 13 4 4 2
15 9 1 0 9 15 13 16 9 0 9 13 0 14 13 2
21 9 1 13 16 11 7 11 1 0 9 1 10 0 9 1 0 13 4 4 4 2
32 9 1 15 14 13 16 11 11 9 1 10 0 9 1 9 13 13 4 2 15 1 13 9 1 9 11 1 9 13 4 4 2
10 10 0 9 1 0 13 4 4 4 2
16 9 1 0 9 1 1 9 1 9 9 1 13 4 4 4 2
14 9 1 9 9 1 1 15 9 14 13 4 4 4 2
21 11 11 11 1 13 4 16 0 9 1 9 1 10 9 11 1 9 13 4 4 2
21 15 11 1 9 1 11 1 0 9 9 1 3 2 3 9 13 1 9 13 4 2
28 11 1 0 9 1 3 3 13 4 13 16 15 10 14 0 13 7 9 1 1 15 13 1 10 9 13 4 2
17 15 1 9 9 1 11 1 9 1 11 12 9 9 1 9 13 2
42 11 11 11 1 11 1 11 11 11 11 1 9 1 11 9 11 11 1 13 4 12 9 1 13 16 11 1 9 11 1 0 9 9 1 9 1 0 9 13 4 4 2
16 15 9 1 0 9 1 9 1 11 1 9 1 9 13 4 2
25 10 9 1 11 11 11 11 2 11 11 11 11 11 7 11 11 11 1 10 0 9 1 9 13 2
11 0 9 1 9 14 10 9 1 0 13 2
20 15 9 11 11 2 11 11 2 9 9 11 11 7 9 11 11 14 0 13 2
34 11 1 11 1 1 11 11 11 11 2 11 2 1 9 1 1 15 9 1 13 16 0 9 1 12 9 1 1 9 1 0 9 13 2
28 15 13 16 15 9 14 0 9 2 9 7 9 9 1 13 9 1 11 1 9 1 1 9 1 1 0 13 2
8 11 11 11 1 0 13 4 2
15 11 1 11 1 12 9 1 9 1 9 1 9 9 13 2
17 15 9 13 16 10 9 1 12 9 1 9 1 10 9 0 13 2
23 11 11 1 0 9 1 1 11 1 9 1 0 13 1 11 1 9 1 14 3 9 13 2
28 11 11 11 11 1 11 11 2 11 2 1 9 1 9 13 4 13 4 16 9 1 15 10 0 7 0 13 2
38 7 12 0 9 1 15 9 1 9 13 16 15 11 11 2 11 2 7 11 11 1 1 9 1 9 1 9 13 15 9 1 9 13 0 13 4 4 2
11 11 10 9 1 0 9 13 1 0 13 2
42 11 1 11 11 11 11 1 11 1 9 1 0 9 1 11 1 13 16 11 2 11 1 0 9 2 9 7 0 9 1 9 7 9 1 10 9 7 0 9 0 13 2
31 15 9 13 16 11 11 1 9 1 9 1 0 9 13 15 15 0 9 1 9 1 1 1 10 0 7 0 13 4 4 2
37 15 11 1 10 9 1 1 9 13 16 15 0 9 1 3 10 9 1 0 13 7 9 13 4 4 16 11 1 11 11 11 11 1 0 9 13 2
31 12 0 9 1 11 1 11 1 9 1 0 13 4 13 16 11 11 7 11 11 1 9 0 0 9 1 1 13 4 4 2
17 15 12 9 1 1 9 9 1 0 9 1 9 13 1 14 13 2
29 15 13 16 9 9 9 1 11 11 1 9 11 2 11 11 2 9 9 7 9 1 1 1 0 9 13 4 4 2
31 9 9 1 1 13 1 9 1 0 2 0 7 0 9 13 1 1 9 13 1 9 1 10 9 1 15 9 13 4 4 2
26 11 11 11 11 11 1 10 9 1 9 13 1 3 10 9 1 10 9 1 15 9 7 9 13 4 2
30 9 1 1 1 13 4 4 0 9 1 9 1 1 13 4 9 9 1 10 9 1 9 10 9 1 15 9 13 4 2
37 9 1 10 9 1 10 9 1 9 13 16 9 1 0 13 1 3 15 0 9 1 9 1 1 9 1 1 9 9 9 1 14 9 0 13 4 2
34 9 1 13 0 9 1 9 1 13 16 9 2 3 7 9 1 9 1 13 1 9 1 1 9 9 1 13 0 9 1 0 14 13 2
10 15 1 10 9 1 9 14 13 4 2
19 9 1 10 9 1 11 11 9 9 1 1 1 14 13 4 1 9 13 2
17 10 9 1 12 9 1 1 9 1 0 9 1 9 9 13 4 2
40 9 1 0 13 4 11 11 11 11 11 11 11 1 13 16 10 9 9 1 1 10 0 9 1 1 9 13 15 15 9 2 9 7 0 7 0 0 9 13 2
14 10 9 1 9 7 9 9 1 0 13 1 9 13 2
15 11 1 11 1 11 2 11 11 11 1 15 9 13 4 2
14 11 1 13 16 11 1 12 9 1 13 0 13 4 2
47 3 2 0 9 7 11 11 11 1 15 9 1 13 2 9 9 9 9 7 0 9 11 11 1 15 9 9 1 9 1 9 1 9 1 13 16 11 1 9 1 1 11 1 0 13 4 2
15 0 9 1 10 9 1 13 15 9 15 14 13 4 4 2
15 16 0 11 11 11 1 11 1 9 1 0 9 13 4 2
29 9 9 1 12 0 9 1 11 2 9 9 11 11 7 11 11 7 11 11 1 9 9 1 0 9 1 9 13 2
22 11 1 0 13 16 15 9 1 9 11 1 0 13 2 15 12 9 9 13 13 4 2
18 15 13 16 15 14 0 9 1 1 9 9 1 9 1 9 13 4 2
41 11 1 0 9 1 1 1 9 1 1 11 1 9 1 9 13 4 11 1 9 11 1 9 13 13 16 0 9 1 9 13 4 16 11 12 0 9 14 13 4 2
24 15 13 16 15 1 1 11 1 14 12 9 13 4 2 7 15 0 11 1 9 13 0 13 2
22 11 1 13 16 11 1 15 9 1 0 13 4 16 16 11 1 15 9 1 13 4 2
23 15 13 16 10 9 13 16 15 9 9 1 0 7 0 9 1 10 9 1 9 13 4 2
33 15 13 9 11 11 2 11 2 1 9 2 10 9 9 1 9 1 0 13 1 3 14 11 7 0 9 1 3 13 4 4 4 2
17 15 11 2 11 7 11 11 1 10 9 9 1 1 1 0 13 2
13 15 12 0 9 1 9 14 1 9 13 4 4 2
37 0 0 0 9 2 11 11 2 1 15 0 12 9 0 13 4 13 4 16 11 11 1 9 7 11 1 9 11 11 14 10 9 1 0 9 13 2
15 10 9 1 9 13 2 0 9 15 12 9 13 4 4 2
26 10 9 1 15 11 1 11 1 9 1 9 13 4 15 15 10 9 1 2 0 2 13 0 13 4 2
13 15 9 1 13 16 10 9 1 9 9 14 13 2
22 9 1 1 11 11 1 9 13 1 9 1 2 11 11 11 11 2 9 1 9 13 2
15 16 0 9 1 9 14 1 12 12 9 1 9 13 4 2
31 9 1 10 9 1 0 13 4 4 16 11 11 1 12 9 1 1 12 1 15 0 13 4 15 0 9 1 9 13 4 2
29 9 1 9 1 11 1 0 11 11 2 9 1 1 9 13 1 0 9 11 7 11 11 11 11 1 9 0 13 2
32 12 0 9 9 2 11 11 2 1 10 9 1 15 9 1 13 4 16 0 9 1 1 9 7 9 1 9 14 0 9 13 2
15 16 9 9 1 13 4 10 9 1 9 13 15 0 13 2
24 9 1 1 1 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 9 13 13 4 2
10 7 11 1 11 12 9 13 4 4 2
17 15 10 9 1 0 9 1 9 1 1 1 0 13 4 4 4 2
25 11 11 9 11 2 11 2 11 2 7 11 2 11 2 11 2 1 0 9 1 9 9 1 13 2
16 11 9 11 11 1 13 16 15 0 9 13 0 13 0 13 2
37 11 11 16 11 7 0 7 0 11 11 1 9 1 13 13 4 2 16 0 0 9 1 14 10 12 9 1 12 9 1 13 1 9 9 13 4 2
25 16 2 11 11 7 11 1 13 1 9 1 12 0 7 0 2 0 9 1 9 1 13 4 4 2
31 9 1 0 9 1 1 10 9 1 13 4 11 11 1 13 16 10 9 0 11 11 7 11 1 9 1 1 3 0 13 2
17 13 9 7 9 1 0 9 1 1 1 15 1 9 13 4 4 2
22 15 1 11 2 11 2 11 7 11 1 9 1 13 1 12 9 1 9 13 4 4 2
28 11 11 1 13 16 9 1 12 9 9 9 1 1 1 11 11 1 12 2 12 9 1 1 0 13 4 4 2
20 9 0 13 1 0 11 11 7 11 1 0 9 1 9 14 0 13 4 4 2
9 11 11 1 15 1 9 13 4 2
12 11 1 11 1 0 9 1 1 0 9 13 2
28 15 1 11 2 11 11 2 11 2 11 2 11 2 11 7 11 1 12 9 1 14 12 9 1 9 13 4 2
22 15 12 12 1 9 0 13 7 0 9 1 0 12 12 1 9 1 9 1 9 13 2
32 9 9 1 12 0 9 1 1 9 1 10 9 13 2 9 1 9 2 9 13 7 9 7 0 9 13 1 12 9 0 13 2
11 15 9 9 9 1 12 9 14 0 13 2
26 15 9 9 13 4 15 11 2 11 2 11 2 11 7 11 11 11 9 1 0 9 1 9 0 13 2
10 11 1 12 9 11 1 9 1 13 2
7 15 11 9 14 0 13 2
47 9 13 9 9 1 9 13 1 9 1 13 11 1 0 9 9 11 11 11 1 11 0 9 2 11 1 11 1 11 9 11 11 11 1 9 7 11 11 1 12 9 1 9 1 9 13 2
26 11 1 9 1 11 1 12 12 1 9 1 1 11 11 1 12 12 1 9 1 12 9 1 9 13 2
17 9 1 0 9 1 9 9 1 12 9 1 9 1 9 13 4 2
32 11 1 11 1 12 9 7 11 11 1 12 9 1 9 9 1 9 1 9 1 9 1 1 11 11 1 12 9 9 13 4 2
16 11 1 9 1 1 12 9 9 0 13 1 9 1 9 13 2
13 11 9 11 11 1 0 9 1 9 9 1 13 2
14 9 1 1 9 1 9 9 7 9 1 14 9 13 2
19 7 9 1 1 9 2 9 1 0 9 7 9 1 9 0 14 13 4 2
21 11 1 13 4 16 11 1 0 9 9 11 11 1 9 13 1 15 9 14 13 2
16 9 1 13 13 16 11 7 11 1 9 15 0 9 14 13 2
10 9 9 1 13 10 9 13 4 4 2
12 3 2 11 1 1 9 1 0 9 14 13 2
17 11 1 9 1 9 13 9 1 9 0 13 1 14 9 13 4 2
21 9 1 13 13 16 15 15 0 9 13 7 15 14 13 4 16 9 1 15 13 2
24 11 9 11 11 11 1 13 16 11 11 1 9 13 1 9 9 1 15 9 1 9 14 13 2
11 16 2 11 1 1 15 9 10 0 13 2
27 9 1 9 13 9 1 9 0 13 1 9 13 4 15 13 16 11 1 10 9 1 15 9 0 14 13 2
33 1 11 2 15 0 9 13 7 10 9 7 9 1 9 13 1 1 0 9 1 9 13 4 1 9 1 9 1 9 13 4 4 2
13 15 13 13 16 15 10 9 1 14 13 4 4 2
39 11 9 11 11 11 14 11 1 9 1 3 1 0 13 4 7 11 11 1 9 11 11 11 1 11 1 14 9 1 3 3 13 1 1 0 13 4 4 2
24 11 1 11 1 11 1 9 13 15 1 11 11 9 1 11 1 3 13 1 0 13 4 4 2
32 11 9 1 11 1 1 11 11 11 1 9 1 9 13 4 11 1 1 11 11 1 11 1 1 9 1 9 0 13 4 4 2
17 11 9 1 11 7 15 9 1 1 9 2 9 0 13 4 4 2
28 11 7 11 1 9 1 9 13 4 11 1 15 0 13 1 14 9 13 16 11 1 9 9 1 1 0 13 2
23 11 1 11 9 1 15 9 13 16 11 1 9 1 1 0 11 9 1 13 9 13 4 2
10 7 11 1 9 15 0 14 13 4 2
26 11 11 1 15 11 1 1 14 11 1 13 9 9 13 4 4 15 11 1 1 9 0 13 4 4 2
31 9 1 1 11 11 1 11 9 11 1 11 1 9 15 9 13 9 13 7 11 1 11 1 3 0 13 1 9 13 4 2
16 11 1 13 9 11 9 11 11 1 14 9 13 13 4 4 2
26 11 11 14 9 11 1 1 13 9 0 13 13 4 4 2 7 15 15 9 1 9 13 11 13 4 2
16 15 15 0 9 11 1 11 1 13 13 1 9 1 9 13 2
34 11 7 11 1 10 9 9 1 3 13 1 11 1 1 15 14 9 13 4 4 16 11 1 0 9 9 0 9 1 9 1 1 13 2
27 11 11 3 1 9 9 1 9 1 13 7 15 10 9 11 1 1 13 9 13 9 1 9 13 4 4 2
17 9 1 0 9 0 9 1 9 1 15 9 2 9 14 13 13 2
17 15 9 13 4 16 10 14 10 0 9 13 1 1 15 9 13 2
7 15 9 9 1 9 13 2
21 9 2 9 1 1 9 13 1 9 0 9 1 9 1 1 10 9 9 13 4 2
19 11 11 11 1 1 2 9 1 0 9 9 12 12 11 9 9 13 4 2
26 3 2 0 9 1 13 7 0 9 9 0 13 1 1 11 11 11 1 9 1 15 0 9 13 4 2
30 9 1 9 11 11 1 13 13 16 0 9 1 13 1 11 13 1 0 9 1 9 1 12 9 1 9 1 9 13 2
36 11 14 14 3 2 3 13 16 11 11 1 9 1 1 15 1 11 9 1 9 1 1 1 9 14 13 7 11 9 11 11 11 15 0 13 2
10 15 1 2 11 9 1 9 15 13 2
4 15 0 13 2
18 0 9 1 15 9 15 9 7 11 1 0 11 11 11 1 1 13 2
25 11 1 11 11 1 13 1 0 9 1 9 1 1 11 1 12 9 1 9 14 0 13 4 4 2
33 11 1 11 1 15 12 9 9 1 15 0 2 0 9 1 13 16 10 15 13 4 16 11 1 1 1 11 9 1 9 15 13 2
7 15 1 15 9 13 15 2
31 15 13 16 11 9 11 2 11 7 11 11 11 1 11 11 11 2 11 2 1 9 13 7 15 1 9 1 9 13 4 2
16 12 9 1 15 13 16 9 7 0 9 9 1 0 9 13 2
15 0 9 1 9 1 15 9 1 9 0 9 0 13 4 2
19 11 1 13 16 12 2 12 9 9 1 15 1 9 9 2 14 13 4 2
23 11 11 7 14 15 1 9 0 13 7 0 9 1 9 1 15 9 13 1 9 9 13 2
38 11 9 11 11 1 10 9 1 16 15 0 9 1 0 9 1 9 13 1 0 14 13 2 11 1 13 16 15 11 1 10 9 1 15 9 0 13 2
17 15 0 9 1 9 13 1 1 9 1 9 13 4 1 9 13 2
22 11 1 11 1 10 12 9 1 9 1 9 13 4 2 15 12 9 7 12 9 13 2
10 7 11 11 1 11 1 0 9 13 2
29 15 1 1 13 4 1 11 1 13 16 11 11 1 11 1 15 9 14 13 7 15 10 9 1 0 13 13 4 2
36 16 0 9 1 15 9 13 16 11 9 1 11 11 2 11 2 9 11 11 1 9 0 13 1 9 1 1 10 9 11 1 1 13 4 4 2
28 11 11 11 1 0 9 1 9 1 12 10 9 7 9 3 14 0 13 1 9 1 9 1 0 13 4 4 2
17 15 13 16 11 11 11 11 1 10 9 13 1 9 13 4 4 2
30 11 1 13 16 12 9 1 1 10 0 9 1 0 9 1 1 0 13 16 11 15 9 1 9 1 9 1 0 13 2
19 15 9 13 16 11 1 0 9 9 0 13 1 9 1 10 0 14 13 2
11 11 11 11 1 15 0 9 1 3 13 2
37 15 3 13 2 15 9 1 9 1 9 13 1 1 9 14 13 4 7 10 9 1 1 12 9 1 9 9 1 3 13 1 1 0 9 13 4 2
11 15 1 9 13 1 0 9 1 9 13 2
20 11 1 9 13 16 12 9 1 9 1 1 9 13 10 15 13 4 4 4 2
19 11 1 15 14 13 16 11 0 9 1 13 0 15 9 1 3 0 13 2
37 15 13 2 16 9 1 13 9 1 1 15 9 13 4 7 11 1 9 7 0 9 1 9 13 4 2 16 15 9 1 0 9 14 13 4 4 2
32 11 1 13 16 11 9 1 9 0 12 9 1 14 13 4 4 2 7 15 9 1 1 15 9 9 0 13 2 0 2 13 2
21 14 12 9 13 9 2 9 1 15 13 16 12 9 1 9 9 3 13 4 4 2
17 9 10 0 9 13 16 2 0 9 2 1 9 13 4 4 4 2
26 15 10 9 1 9 1 1 0 13 2 15 1 14 15 11 11 11 11 1 2 0 9 2 13 4 2
30 11 1 13 16 11 1 1 15 0 7 3 0 0 2 9 15 13 4 16 0 9 1 0 9 1 9 1 13 4 2
19 0 9 1 9 1 11 1 9 1 0 9 11 11 1 0 9 13 4 2
12 15 15 9 1 9 7 9 1 9 14 13 2
21 2 0 11 2 11 9 11 11 7 0 11 11 11 11 1 9 1 13 4 4 2
20 9 1 15 1 13 4 9 1 0 9 1 9 1 9 13 1 9 14 13 2
20 16 15 11 1 14 0 9 1 1 11 1 2 11 2 11 11 2 0 13 2
29 1 9 2 2 10 9 1 0 13 1 1 15 10 9 13 4 7 15 15 0 9 1 9 1 13 1 1 0 13
35 9 1 15 9 7 9 1 1 1 9 0 13 4 13 16 2 0 9 2 7 0 2 0 9 1 1 13 10 9 1 13 1 9 13 2
27 15 11 7 11 1 0 13 4 15 10 9 1 0 2 0 9 1 13 7 9 1 9 13 1 9 13 2
29 11 11 1 1 9 1 1 0 9 1 13 15 9 1 13 4 11 1 13 16 12 9 1 1 9 1 9 13 2
20 11 7 11 1 9 13 4 9 1 11 11 1 13 9 1 13 1 9 13 2
13 11 1 13 16 15 15 9 1 1 9 14 13 2
26 9 1 9 9 2 9 2 0 9 7 0 9 1 9 9 1 9 13 4 2 15 15 9 13 4 2
23 15 13 16 15 9 1 9 0 13 1 1 11 1 9 0 13 1 3 10 9 13 4 2
45 2 11 2 11 11 2 1 1 0 9 13 1 9 1 9 13 4 11 1 13 16 15 0 2 0 9 13 2 15 15 7 9 9 11 11 11 11 1 11 1 9 13 4 4 2
14 10 9 1 0 9 13 1 1 12 9 14 13 4 2
25 1 11 2 7 11 1 15 0 9 1 2 12 9 1 1 9 2 13 4 9 0 13 4 4 2
32 15 13 4 1 16 15 15 1 11 1 9 11 1 13 13 4 2 9 1 13 16 15 9 1 10 9 11 1 13 13 4 2
22 11 1 13 16 9 1 9 13 1 9 9 1 0 9 1 1 1 10 9 13 4 2
28 9 1 1 9 9 1 9 14 13 1 11 9 11 11 1 9 1 11 1 13 2 2 15 15 13 4 4 2
12 15 10 9 1 3 13 13 1 0 9 13 2
15 15 15 9 1 9 2 15 9 7 0 9 1 9 14 13
32 15 13 4 1 16 15 15 1 11 1 9 11 1 13 13 4 2 11 1 13 16 15 9 1 10 9 11 1 13 14 13 4
29 0 9 1 9 1 9 1 11 1 9 13 1 1 11 15 0 9 1 1 14 11 1 0 9 1 9 13 4 2
24 3 11 1 11 11 11 1 9 13 4 1 9 13 2 15 11 1 3 0 9 9 13 4 2
19 11 11 11 1 13 11 11 1 11 11 1 9 13 1 9 1 13 4 2
17 11 1 13 11 7 11 11 1 0 13 1 1 11 13 4 4 2
23 11 1 1 11 1 0 9 1 11 1 9 1 9 14 13 4 4 0 9 1 13 4 2
20 11 1 10 9 1 9 13 4 15 0 9 1 1 9 1 9 14 13 4 2
21 0 9 1 9 1 0 9 1 14 9 1 9 1 3 2 3 0 13 4 4 2
37 11 9 11 11 1 13 16 11 1 9 1 9 13 1 0 13 4 7 10 9 11 1 0 13 4 16 9 1 13 9 1 15 15 9 14 13 2
31 11 1 13 16 11 7 11 1 11 1 15 9 1 9 13 4 7 15 9 1 10 10 0 9 13 15 1 0 9 13 2
10 11 1 10 9 1 9 14 13 4 2
44 11 1 10 9 1 0 9 13 16 9 9 1 14 9 7 3 11 1 1 1 0 9 1 9 3 3 14 13 4 7 15 13 1 1 11 1 14 0 9 1 9 13 4 2
19 0 9 1 14 11 11 2 11 11 11 7 11 11 1 9 13 4 4 2
16 7 15 11 1 11 11 11 1 1 11 1 9 1 13 4 2
15 11 9 1 11 1 10 9 1 11 1 14 9 13 4 2
28 11 1 13 16 11 1 9 0 13 2 16 15 9 14 1 11 11 11 1 11 1 9 13 9 9 13 4 2
11 10 9 1 1 14 15 11 13 4 4 2
19 11 1 11 11 11 1 1 13 9 1 9 9 1 10 9 1 13 4 2
19 11 1 0 9 3 9 1 9 13 11 9 1 9 13 1 13 4 4 2
13 7 9 10 9 11 1 13 1 9 14 13 13 2
31 16 2 9 11 11 11 1 1 11 1 13 1 9 1 1 11 1 0 9 9 1 9 1 1 1 11 9 1 0 13 2
18 15 0 9 13 15 9 9 0 9 1 0 9 1 9 13 4 4 2
28 9 9 1 9 1 1 11 13 0 11 9 11 11 2 11 11 7 11 11 1 15 1 9 13 9 0 13 2
18 10 10 9 1 13 13 16 15 9 1 9 1 9 9 1 1 13 2
24 13 4 4 4 16 11 1 0 9 1 9 1 1 11 1 9 9 1 9 1 9 13 4 2
23 7 9 9 1 9 11 1 11 11 1 13 4 9 1 0 9 1 9 1 1 14 13 2
9 15 1 14 9 1 9 14 13 2
18 9 10 9 1 0 9 1 9 9 1 13 1 14 9 13 4 4 2
16 11 11 11 1 11 1 0 11 11 11 11 1 9 13 4 2
16 9 1 1 11 1 11 1 15 1 3 13 13 1 9 13 2
14 11 1 10 9 1 9 1 10 9 13 4 4 4 2
14 16 11 10 9 1 11 1 9 1 0 13 4 4 2
10 15 1 9 14 3 9 13 4 4 2
32 9 1 9 15 13 16 11 1 15 1 10 9 11 11 1 10 15 9 14 13 15 9 1 9 1 15 3 7 15 0 13 2
28 9 1 9 13 16 15 9 0 9 7 11 1 1 9 2 9 13 4 16 9 1 15 9 1 9 14 13 2
20 11 11 11 11 1 9 1 11 9 14 12 12 11 9 15 9 1 13 4 2
18 15 1 11 9 9 11 1 9 7 9 1 1 11 1 9 13 4 2
14 9 1 1 11 11 11 9 11 0 11 9 13 4 2
11 15 9 1 10 9 15 9 1 0 13 2
22 10 9 1 11 1 9 1 0 13 4 13 16 15 0 9 13 9 9 1 13 4 2
22 11 1 9 1 15 9 13 4 9 13 16 15 1 15 9 1 9 14 13 4 4 2
22 15 13 16 11 1 9 1 9 7 9 1 1 13 9 1 12 0 9 9 13 4 2
15 0 13 16 11 1 9 7 9 1 0 9 13 4 4 2
11 15 12 9 7 10 9 0 13 4 4 2
8 15 1 9 10 13 4 4 2
19 9 9 11 11 1 9 1 11 1 11 1 9 1 11 11 1 9 13 2
14 11 11 1 9 1 1 10 9 1 0 9 13 4 2
28 11 9 9 9 9 1 9 1 1 11 11 11 11 11 11 11 1 9 7 9 1 1 11 1 9 13 4 2
38 10 9 1 11 11 7 9 9 9 9 1 9 7 0 9 11 11 1 9 1 9 1 9 1 12 9 1 1 14 9 9 1 9 1 14 9 13 2
19 9 13 1 3 11 9 11 11 15 14 9 1 9 1 0 13 13 4 2
25 15 14 12 9 9 11 0 11 11 11 11 11 11 1 9 1 9 1 0 9 9 1 1 13 2
17 15 9 1 13 1 3 14 15 14 12 12 9 0 13 4 4 2
11 11 1 9 1 10 9 9 9 1 13 2
12 10 0 9 0 9 0 13 1 9 1 13 2
11 15 1 9 7 9 9 9 1 13 4 2
20 11 1 9 9 7 9 1 9 1 9 1 9 1 0 9 13 1 9 13 2
45 11 1 9 1 9 13 2 0 9 13 7 0 9 1 9 13 1 13 13 4 9 1 1 1 13 4 12 9 1 9 1 13 16 0 9 1 15 0 13 4 15 0 13 4 2
21 9 1 0 13 1 3 11 1 11 9 1 9 1 9 1 1 1 12 9 13 2
33 10 9 1 9 1 9 7 0 9 9 11 11 2 0 9 1 9 11 11 7 9 9 7 11 9 1 9 11 11 14 0 13 2
26 9 1 1 9 1 12 0 9 9 1 9 1 9 13 1 10 9 1 11 1 9 1 13 4 4 2
11 0 9 9 1 12 9 14 13 4 4 2
22 9 1 1 9 12 9 1 15 9 9 1 1 14 13 7 0 9 1 15 9 13 2
14 9 1 13 1 3 15 12 9 0 9 13 4 4 2
10 0 9 9 1 1 9 14 13 4 2
18 9 1 1 9 1 9 1 15 1 10 9 13 4 15 0 13 4 2
39 9 7 9 1 1 15 13 14 9 13 4 16 16 9 0 9 13 2 0 9 13 7 0 13 7 0 9 13 15 14 12 9 1 15 9 1 9 13 2
16 9 1 1 9 1 0 9 9 0 13 7 15 9 14 13 2
16 11 11 11 1 13 4 12 9 1 0 13 1 9 13 4 2
7 15 0 14 13 4 4 2
7 9 9 1 9 3 13 2
33 11 11 11 2 11 2 1 9 9 1 9 9 7 9 1 1 9 14 13 4 1 1 11 1 15 1 15 9 14 13 4 4 2
30 9 11 2 11 1 1 11 9 9 1 15 0 9 14 13 4 1 1 3 10 9 1 9 13 1 13 4 4 4 2
15 15 11 11 11 2 11 2 1 9 11 11 1 3 13 2
17 3 10 12 9 1 1 12 9 9 9 1 9 11 1 13 4 2
15 7 11 11 1 15 1 10 9 1 9 0 14 13 4 2
38 15 1 11 2 11 1 1 14 9 1 9 1 12 1 9 1 9 1 9 0 13 4 4 7 11 2 11 1 1 9 9 1 0 14 13 4 4 2
25 11 1 9 1 1 9 1 9 1 11 11 11 11 11 1 13 16 9 9 1 13 0 9 13 2
14 7 9 14 13 4 1 1 15 9 14 13 4 4 2
22 3 14 9 13 1 3 10 9 3 13 15 13 4 9 9 0 13 1 9 3 13 2
12 15 11 1 9 11 11 1 3 13 4 4 2
28 3 2 9 9 1 15 1 1 15 14 0 13 1 9 13 4 16 9 11 9 9 1 15 9 13 4 4 2
21 11 1 9 7 9 9 1 0 9 9 1 1 12 9 9 9 1 9 13 4 2
15 16 15 1 9 9 13 11 11 1 9 1 0 13 4 2
17 16 9 1 1 9 12 1 12 1 9 9 9 1 13 4 4 2
15 15 1 0 0 9 1 9 0 9 1 13 4 4 4 2
31 11 11 11 7 11 11 11 3 12 9 9 9 1 9 13 4 4 3 10 9 13 4 16 12 1 9 9 0 13 4 2
21 11 1 0 11 11 11 1 9 11 11 1 1 9 12 9 9 9 13 4 4 2
39 9 9 1 13 16 0 9 1 9 1 11 11 1 0 9 13 1 3 9 13 4 4 1 1 0 12 9 1 9 9 1 1 14 9 0 14 13 4 2
22 9 11 2 11 1 1 12 1 9 1 9 9 9 1 9 1 0 13 4 4 4 2
14 7 9 11 2 11 1 1 1 15 15 0 14 13 2
25 0 9 1 10 0 9 1 12 9 9 9 2 15 12 9 9 0 13 2 13 1 9 13 4 2
19 7 11 11 1 1 1 9 14 13 1 1 15 9 0 14 13 4 4 2
30 10 9 1 14 9 1 9 13 4 4 16 14 12 12 9 1 9 1 9 11 2 11 1 1 10 9 9 0 13 2
16 16 9 1 15 15 9 1 9 13 1 9 1 9 13 4 2
37 3 14 12 12 10 9 1 10 9 1 9 13 4 4 4 15 7 14 0 13 4 7 14 15 1 15 9 1 1 11 9 1 9 13 4 4 2
38 11 11 11 11 1 0 9 1 9 1 10 13 1 1 12 12 9 1 11 2 11 9 9 1 11 1 0 9 1 9 1 13 4 1 9 13 4 2
28 11 11 1 9 1 13 16 0 9 1 9 1 9 1 1 11 1 1 9 11 1 11 1 9 1 1 13 2
20 11 1 13 1 12 9 0 9 9 1 1 11 11 11 1 3 14 9 13 2
22 9 9 11 11 1 3 9 1 11 1 11 1 1 15 9 1 13 1 9 13 4 2
21 7 2 11 1 10 9 1 10 9 13 1 1 9 1 0 9 1 9 13 4 2
25 9 1 13 16 12 9 0 9 1 1 9 1 9 9 11 1 9 13 1 9 0 13 4 4 2
23 11 1 9 13 1 3 1 9 1 9 11 11 11 11 11 2 11 2 1 3 14 13 2
36 11 9 1 9 1 1 9 1 9 1 11 1 13 4 1 9 9 1 9 9 1 9 0 13 1 1 11 1 0 9 1 11 1 9 13 2
27 9 9 1 0 9 1 9 1 9 2 9 2 9 7 9 0 13 1 1 12 0 9 0 13 4 4 2
15 11 11 11 11 11 9 1 9 1 10 9 13 4 4 2
30 9 10 9 0 13 13 4 15 14 0 0 9 1 9 1 15 9 2 9 7 15 9 1 15 9 1 9 14 13 2
13 0 13 16 11 11 1 11 11 11 13 4 4 2
19 9 1 1 9 1 9 0 13 1 9 1 12 9 1 9 1 9 13 2
14 11 2 9 2 9 1 9 1 9 1 9 13 4 2
20 10 9 0 9 1 9 2 9 1 9 7 9 2 9 1 9 1 9 13 2
11 9 1 9 1 15 9 1 9 14 13 2
10 10 9 1 9 1 1 0 9 13 2
18 9 1 9 1 1 15 14 9 12 9 9 1 1 9 13 4 4 2
32 9 1 1 11 11 11 11 11 1 9 1 0 9 7 9 1 0 9 1 9 1 1 10 9 1 9 13 1 9 13 4 2
22 11 11 1 9 1 9 13 1 3 14 0 9 1 1 0 9 9 1 9 13 4 2
16 9 1 15 9 9 1 12 9 1 9 1 9 13 4 4 2
17 9 1 9 13 1 1 0 9 15 2 9 9 2 13 4 4 2
12 10 9 1 15 0 9 14 0 13 4 4 2
42 11 11 11 11 11 1 0 11 9 11 11 1 9 1 13 9 1 2 9 9 2 1 1 0 13 1 3 11 11 11 14 2 9 9 2 1 9 1 13 4 4 2
36 11 11 1 3 0 9 15 13 16 15 15 10 9 9 14 13 4 4 4 2 15 9 1 1 0 11 1 9 1 1 1 0 13 4 4 2
18 15 9 13 16 2 9 9 2 1 9 1 9 1 9 1 9 13 2
22 9 1 1 9 1 1 1 14 9 9 1 1 13 1 9 1 0 13 4 4 4 2
14 7 9 13 16 0 13 1 9 14 14 13 4 4 2
18 2 9 9 2 1 1 10 0 0 9 1 9 1 9 14 13 4 2
24 7 10 9 1 15 14 15 9 1 1 13 4 1 1 1 9 9 0 13 1 13 4 4 2
20 11 11 1 13 9 14 0 9 1 2 9 9 2 13 1 9 1 14 13 2
16 15 13 13 16 9 1 15 0 9 1 15 9 14 13 4 2
13 7 0 0 9 15 14 15 9 1 13 4 4 2
15 9 9 1 10 0 9 14 9 9 1 9 1 0 13 2
23 7 15 1 15 10 9 14 13 2 15 0 11 1 1 1 9 1 1 0 13 4 4 2
28 16 2 11 11 1 13 10 9 1 11 11 7 11 1 9 1 9 13 4 1 11 11 1 10 9 13 4 2
11 7 11 11 11 15 1 14 0 14 13 2
24 11 11 1 0 9 1 13 13 16 11 11 1 9 13 1 1 2 9 9 2 3 0 13 2
19 0 9 1 9 1 9 1 1 2 9 9 2 1 9 3 0 13 4 2
26 15 9 1 9 1 1 9 13 7 9 1 9 1 9 13 1 1 11 11 11 9 9 13 13 4 2
21 1 15 2 9 1 1 9 9 12 7 0 9 1 13 10 9 14 13 4 4 2
14 9 9 1 1 9 9 9 13 1 1 14 0 13 2
19 11 11 11 0 9 1 9 9 9 1 10 0 9 3 0 13 4 4 2
18 15 9 1 10 9 14 13 2 15 1 9 9 1 9 13 4 4 2
13 9 1 0 13 1 0 9 1 9 13 4 4 2
24 10 9 1 9 9 1 9 1 11 11 1 11 1 9 9 9 9 13 1 9 0 13 4 2
20 9 9 1 1 9 1 9 9 9 1 9 1 9 1 0 13 0 9 13 2
18 9 9 1 15 9 1 0 9 13 1 3 9 9 9 1 13 4 2
22 9 9 1 13 9 1 1 0 12 2 12 9 1 9 1 9 1 10 9 0 13 2
22 15 9 1 1 0 9 1 9 1 1 9 13 15 13 1 15 15 9 1 14 13 2
19 9 1 9 1 15 9 0 9 1 14 13 15 15 9 2 9 13 4 2
11 15 1 9 1 10 9 1 9 13 4 2
8 15 1 9 1 9 9 13 2
31 9 1 1 9 9 1 9 1 9 1 13 1 9 13 2 7 15 1 0 13 9 1 1 1 15 9 14 13 4 4 2
17 10 0 9 1 1 9 1 9 1 9 1 0 13 1 13 4 2
17 0 9 9 1 1 14 10 9 0 9 1 0 13 4 4 4 2
34 15 1 0 9 11 9 1 14 11 1 11 9 1 12 0 9 1 9 13 4 4 2 15 9 9 9 1 10 0 9 0 13 4 2
27 9 1 9 1 11 1 13 4 16 11 1 9 9 15 0 9 1 9 9 1 9 1 9 13 9 13 2
11 10 9 0 13 2 15 14 0 13 4 2
24 11 11 11 1 0 9 11 11 1 0 9 1 9 1 11 1 9 1 0 9 13 4 4 2
12 9 1 13 13 16 9 1 9 13 4 4 2
34 9 9 2 9 2 11 11 1 15 13 16 11 1 9 9 1 9 1 1 11 11 1 9 7 9 1 13 4 9 1 9 14 13 2
24 15 15 13 4 16 9 9 1 1 11 1 9 13 7 13 1 9 1 1 15 13 4 4 2
17 11 1 13 16 11 1 11 11 11 11 1 9 12 9 1 13 2
15 10 9 1 13 4 4 16 9 1 0 9 13 4 4 2
17 15 9 1 9 14 13 7 9 14 9 2 3 13 9 13 4 2
12 15 13 16 9 1 9 3 14 13 9 13 2
46 15 13 4 1 16 15 11 11 1 0 9 13 4 4 4 2 11 1 13 16 9 1 10 9 1 1 13 4 9 1 9 15 9 1 3 0 13 4 15 15 9 3 0 13 4 2
20 15 13 16 10 9 1 0 9 1 1 12 0 9 1 9 14 13 4 4 2
39 0 13 16 0 9 11 1 11 1 11 1 0 9 1 9 1 1 10 9 9 1 9 13 1 1 11 1 9 1 9 1 11 11 1 9 13 4 4 2
26 11 11 11 7 0 11 11 11 11 11 1 11 1 11 1 12 9 1 1 10 0 9 1 9 13 2
27 11 11 1 10 9 1 9 13 4 16 11 1 1 15 14 9 1 11 1 9 1 15 9 14 13 4 2
13 11 11 1 9 1 15 0 7 0 9 13 4 2
33 11 9 1 15 1 13 9 1 9 1 11 1 13 16 15 12 0 9 13 4 15 15 14 9 1 14 9 1 0 14 13 4 2
31 10 9 15 10 9 1 9 1 13 16 15 11 11 11 1 11 1 9 9 13 13 15 15 15 11 9 1 14 9 13 2
42 0 9 11 1 11 1 11 1 11 1 7 11 1 11 1 15 9 1 1 0 12 9 1 1 1 11 1 13 16 15 1 15 15 13 4 2 15 15 1 0 13 2
15 11 1 1 11 2 11 1 9 1 10 15 0 13 4 2
16 0 9 1 12 9 0 13 4 4 7 0 9 13 4 4 2
31 11 1 11 1 12 0 0 9 2 11 11 2 1 13 4 9 1 13 16 11 11 9 1 15 0 7 0 9 13 4 2
12 12 9 1 1 0 9 7 9 13 4 4 2
20 11 2 11 1 1 9 7 9 1 9 0 13 1 1 9 9 0 13 4 2
21 15 3 14 0 13 4 4 16 10 9 9 9 1 9 1 9 13 1 0 13 2
33 10 3 0 9 1 15 13 16 11 2 11 9 9 1 13 1 10 9 3 13 4 4 4 7 0 9 11 11 1 0 13 4 2
18 12 9 1 9 13 4 16 15 3 13 7 9 1 12 0 9 13 2
34 12 9 1 9 1 0 9 1 9 13 4 1 9 13 4 11 1 13 16 10 9 1 9 15 0 11 11 11 1 14 9 13 4 2
55 15 13 4 1 16 15 11 1 9 2 9 13 4 1 0 9 1 11 2 11 11 11 11 1 9 13 4 2 11 1 9 13 16 15 0 9 1 13 4 4 16 10 9 10 9 13 15 12 9 1 10 9 0 13 2
6 15 15 9 13 4 2
14 11 1 11 1 11 1 1 0 9 7 9 14 13 2
16 15 13 11 1 9 1 1 11 15 1 9 9 1 1 13 2
10 11 10 9 1 11 1 1 0 13 2
16 9 1 0 7 0 9 9 1 0 9 9 1 13 4 4 2
38 11 7 11 1 9 1 13 11 11 11 1 13 4 4 7 0 12 9 1 9 1 9 13 1 0 9 1 9 1 13 4 1 9 10 13 4 4 2
33 15 16 11 1 0 9 1 9 13 4 16 14 9 1 9 13 4 4 2 16 9 14 9 1 9 9 1 9 1 13 4 4 2
20 11 9 15 9 9 13 15 0 0 9 1 0 9 1 0 9 1 9 13 2
20 0 9 1 11 9 1 9 1 9 13 7 9 1 3 15 9 1 13 4 2
15 11 9 0 9 11 11 7 11 11 1 3 0 9 13 2
26 7 11 11 11 1 9 1 13 4 7 9 9 9 1 9 9 13 9 9 1 15 9 0 13 4 2
7 15 1 11 14 13 4 2
10 0 11 14 3 13 9 1 13 4 2
16 9 13 16 0 9 1 0 0 9 12 9 1 0 13 4 2
17 12 9 1 9 1 1 11 9 1 0 9 1 13 13 9 13 2
12 9 11 11 7 11 11 1 0 10 9 13 2
12 11 1 15 1 12 9 1 9 13 4 4 2
13 10 13 9 11 1 9 1 1 13 4 4 4 2
17 3 11 1 11 1 11 11 1 9 9 1 9 14 13 4 4 2
13 15 3 13 9 1 15 0 9 9 1 13 4 2
27 11 9 9 10 9 1 12 0 9 14 13 7 15 1 1 14 11 1 9 1 9 1 0 13 4 4 2
16 9 1 9 1 1 11 1 9 1 9 10 0 13 4 4 2
17 9 1 9 1 1 11 1 12 0 9 9 1 0 13 4 4 2
18 9 1 1 15 1 14 9 7 0 9 13 4 1 9 14 13 4 2
14 11 1 0 9 1 1 14 9 1 3 13 4 4 2
36 11 1 1 9 1 13 0 9 1 9 10 9 0 13 4 2 15 11 9 11 11 1 9 1 0 9 1 9 11 11 1 9 0 13 4 2
18 7 2 0 9 1 1 0 9 1 11 11 9 1 1 1 0 13 2
17 9 1 9 1 14 12 0 9 13 2 11 1 9 11 11 1 2
20 0 9 9 1 1 11 1 9 11 11 11 1 9 1 9 1 13 4 4 2
21 11 11 1 11 11 9 2 11 11 9 7 11 11 1 9 1 9 13 4 4 2
15 11 7 14 11 1 1 13 11 11 1 9 13 4 4 2
17 11 1 15 9 1 9 7 9 1 12 2 12 9 0 13 4 2
53 11 11 2 9 9 1 1 11 1 0 13 1 11 11 2 7 0 0 9 11 11 11 7 2 9 9 2 11 11 2 2 11 2 11 11 7 11 11 11 1 0 9 1 0 9 1 1 1 0 13 4 4 2
15 11 11 2 11 11 7 11 11 11 9 1 9 13 4 2
12 11 1 9 11 1 0 9 1 9 0 13 2
16 15 13 16 9 7 9 1 12 0 9 3 14 13 4 4 2
16 11 11 1 9 1 9 13 1 1 9 1 9 13 4 4 2
20 9 1 13 13 16 11 11 1 9 1 0 13 4 11 11 1 0 14 13 2
30 11 1 9 1 11 9 1 9 1 9 2 11 11 1 9 1 0 9 7 11 9 9 1 9 1 9 1 0 13 2
18 15 15 14 0 9 13 11 11 1 11 11 1 11 1 9 14 13 2
13 11 11 1 11 11 11 1 9 14 13 4 4 2
18 11 1 9 1 11 1 0 9 1 14 0 9 1 9 13 4 4 2
21 11 9 1 11 1 11 9 1 13 4 11 11 1 0 9 1 0 13 4 4 2
35 10 9 11 1 11 1 9 1 9 13 11 1 2 9 2 1 1 13 11 1 9 1 9 1 9 13 4 1 9 0 13 4 4 4 2
12 7 15 0 9 1 9 1 9 13 4 4 2
24 11 11 11 7 11 11 11 1 11 11 7 11 11 1 12 0 9 9 1 0 13 4 4 2
10 9 1 11 11 7 11 11 14 13 2
15 11 1 0 11 11 11 1 14 9 1 0 13 4 4 2
24 11 11 1 9 9 1 13 4 11 11 1 0 9 1 0 9 1 1 1 0 13 4 4 2
12 9 1 0 9 11 11 14 9 1 0 13 2
13 15 9 11 11 11 1 9 1 9 13 4 4 2
12 9 1 10 12 9 1 14 12 9 0 13 2
9 9 1 9 1 15 9 14 13 2
21 9 1 12 9 0 13 2 15 1 12 9 0 9 1 1 1 0 13 4 4 2
26 11 11 11 1 13 16 9 1 0 9 2 9 9 9 7 9 9 14 1 3 14 9 13 4 4 2
40 11 11 1 11 9 14 9 1 9 1 9 9 13 1 9 1 9 13 4 4 7 9 9 1 9 1 9 1 13 14 4 7 9 1 11 9 1 13 4 2
35 9 9 1 0 0 9 1 13 13 16 10 9 11 1 0 9 11 1 0 13 4 7 3 11 2 11 7 11 0 9 1 15 9 13 2
16 11 11 1 11 9 14 12 9 9 1 9 1 8 13 4 2
23 0 9 0 9 1 1 13 4 15 11 1 1 11 9 9 9 1 9 1 13 4 4 2
30 9 9 1 0 0 9 1 1 9 14 12 9 11 9 1 0 9 1 9 1 9 13 4 1 9 13 4 4 4 2
16 11 1 0 9 7 0 9 1 1 9 1 9 13 4 4 2
10 15 1 9 1 9 3 0 9 13 2
15 15 1 9 1 3 9 1 9 9 1 9 9 13 4 2
23 11 1 0 9 1 9 1 1 14 10 9 1 9 9 9 1 9 1 9 13 4 4 2
31 9 1 9 1 9 13 1 3 14 9 1 10 9 1 9 13 4 4 16 10 9 1 9 1 15 9 1 9 9 13 2
23 9 9 1 9 1 13 13 16 9 9 1 0 9 7 15 9 3 9 1 14 13 4 2
23 0 3 0 9 1 15 14 9 13 16 9 9 1 9 1 1 0 9 11 1 9 13 2
24 9 1 13 13 16 12 0 0 9 1 9 1 9 13 4 9 13 1 9 14 13 4 4 2
24 15 1 1 9 1 9 9 1 1 11 2 11 2 11 7 11 11 11 1 9 3 13 4 2
23 9 1 15 14 9 13 16 9 7 15 9 2 1 11 11 1 15 10 9 13 4 4 2
12 3 15 1 15 1 0 14 13 4 4 4 2
26 9 1 11 1 9 13 1 3 14 0 11 1 11 1 13 4 0 9 1 9 13 9 13 4 4 2
27 9 9 9 1 14 10 9 1 9 13 1 1 9 13 4 15 0 9 1 0 9 8 13 4 4 4 2
13 11 9 11 11 15 9 9 1 13 0 14 13 2
14 15 10 9 1 14 15 9 9 1 9 13 4 4 2
17 10 9 1 1 15 0 9 1 9 1 13 9 1 10 0 13 2
13 11 11 1 13 16 9 15 9 1 9 13 4 2
20 9 1 9 1 1 15 9 9 1 9 14 13 15 15 10 13 4 4 4 2
7 15 15 15 9 14 13 2
13 11 0 9 1 9 1 1 9 1 0 14 13 2
14 15 13 13 0 9 1 14 9 1 9 13 4 4 2
14 10 9 1 15 15 13 4 15 15 9 14 13 4 2
28 15 13 16 11 9 2 11 11 11 2 9 1 0 13 7 2 11 11 2 2 11 2 0 9 1 9 13 2
24 9 9 10 13 1 1 1 13 4 1 15 13 16 15 15 15 14 9 1 9 14 13 4 2
11 15 9 7 9 1 9 1 13 4 4 2
9 15 15 1 1 15 14 13 4 2
29 0 9 1 9 1 9 1 15 9 1 1 1 13 1 15 13 16 15 11 1 12 9 1 9 1 1 13 4 2
10 15 1 9 9 1 1 1 11 13 2
14 15 0 9 1 13 4 9 1 15 10 9 13 4 2
11 15 9 1 0 9 1 0 9 13 4 2
23 15 0 13 4 16 16 13 0 9 1 3 9 14 13 4 16 0 9 0 13 4 4 2
51 11 1 11 1 11 2 11 11 2 11 1 9 13 4 11 1 13 16 2 9 1 0 9 1 1 1 15 3 0 13 2 16 11 7 9 1 0 0 9 0 9 1 12 2 12 9 13 4 4 2 2
21 15 3 13 16 16 9 1 9 14 13 4 16 9 1 0 9 0 13 4 4 2
16 0 9 1 9 13 1 1 0 9 1 15 3 9 13 4 2
12 9 1 1 15 10 10 14 9 13 4 4 2
20 15 10 9 1 2 0 2 13 7 15 0 9 1 0 9 13 1 9 13 4
18 11 11 1 10 9 1 9 1 15 9 1 0 13 1 9 13 4 2
16 15 1 15 10 9 9 9 1 13 9 1 14 9 13 4 2
11 10 9 1 1 0 9 0 13 4 4 2
31 11 1 10 0 9 1 10 9 1 9 13 4 16 15 9 1 13 9 9 1 0 13 1 9 7 9 1 1 1 13 2
17 15 13 2 2 10 9 1 9 9 3 14 9 14 13 4 4 2
14 10 9 12 1 12 12 12 9 1 9 13 4 4 2
18 0 9 1 9 14 13 4 4 7 9 15 0 9 13 1 0 14 13
29 11 1 13 16 16 9 1 9 13 4 16 11 11 11 1 9 1 9 13 4 7 9 7 9 9 1 13 4 2
28 15 13 16 0 9 1 0 9 13 4 4 4 2 7 0 9 16 10 9 13 4 16 9 0 13 4 4 2
25 9 1 0 9 1 9 13 4 15 13 16 9 9 1 9 0 9 1 9 1 13 4 4 4 2
37 15 13 16 10 9 1 9 1 2 11 11 2 11 11 11 11 11 0 13 4 2 15 1 0 12 9 1 12 12 12 12 12 9 9 13 4 2
34 0 11 11 11 9 1 11 9 11 1 9 9 14 1 13 4 1 9 15 13 2 11 11 1 15 9 1 9 13 9 13 4 4 2
30 11 1 11 9 1 0 11 1 9 11 1 11 1 9 1 9 1 13 16 10 9 11 1 0 0 9 1 13 4 2
21 15 13 4 4 16 11 1 10 9 11 9 1 9 1 9 1 13 14 13 4 2
28 12 9 1 15 15 12 14 9 1 13 2 15 14 15 11 9 7 11 1 9 1 1 1 10 15 13 4 2
15 0 13 16 11 9 1 0 11 9 1 14 11 0 13 2
20 11 1 9 9 11 11 1 9 1 11 9 0 2 0 0 9 1 9 13 2
28 9 1 0 9 7 11 1 11 11 1 9 1 1 9 1 9 13 4 9 10 10 14 0 9 13 4 4 2
16 10 9 1 9 9 11 11 1 13 9 11 11 1 0 13 2
18 15 1 0 0 9 11 11 1 0 10 9 1 10 9 9 13 4 2
7 9 1 9 3 13 4 2
14 10 9 11 1 0 9 1 9 1 0 13 4 4 2
15 16 2 15 9 11 11 1 1 14 15 0 14 9 13 2
11 11 15 0 9 11 1 9 13 4 4 2
22 9 11 1 9 1 15 11 1 9 13 4 15 10 9 9 9 11 11 1 9 13 2
12 9 1 1 9 1 1 9 1 0 9 13 2
17 10 9 1 9 13 4 4 2 15 1 9 9 0 13 4 4 2
15 11 1 0 9 9 7 9 1 3 14 13 4 4 4 2
15 9 1 1 11 1 0 9 9 13 15 0 13 4 4 2
28 9 1 13 16 11 1 10 0 12 9 11 1 15 14 9 1 9 2 9 1 1 3 0 9 1 13 4 2
16 10 3 9 1 15 15 9 1 1 3 11 7 11 13 4 2
30 10 9 15 11 9 1 10 0 9 1 9 13 15 15 10 9 11 13 4 7 15 11 11 1 15 9 1 9 13 2
14 7 11 7 15 9 11 11 2 11 1 11 1 13 2
13 16 2 11 1 15 9 9 1 13 14 4 4 2
19 15 11 11 1 14 11 9 1 1 15 9 7 9 1 1 9 13 4 2
14 10 9 1 11 15 9 7 9 1 1 13 4 4 2
11 3 1 9 1 9 1 1 9 0 13 2
27 10 9 1 9 15 9 1 9 13 15 9 9 9 1 12 9 9 1 13 4 7 0 9 0 13 4 2
7 3 1 15 9 13 4 2
5 9 0 9 13 2
27 11 1 15 9 1 10 0 13 4 4 16 9 1 13 1 9 1 3 1 15 9 13 1 0 14 13 2
13 16 2 11 1 1 15 15 1 9 11 1 13 2
7 15 11 11 1 9 13 2
22 11 2 11 11 13 4 4 2 15 11 1 9 2 9 1 15 1 9 0 13 4 2
33 11 1 0 3 0 9 11 1 9 1 9 13 1 1 0 13 4 0 2 0 11 2 11 9 9 11 1 9 1 13 4 4 2
25 11 1 9 2 9 2 1 3 9 13 1 3 11 1 10 0 9 1 9 13 9 13 4 4 2
12 10 9 11 1 0 9 9 11 1 13 4 2
37 11 1 12 9 1 13 16 11 0 11 1 9 9 9 1 0 9 1 1 11 9 12 9 11 1 9 13 16 15 15 9 1 0 13 4 4 2
34 9 1 13 16 10 9 13 14 9 1 9 9 1 13 9 9 9 1 13 4 7 11 1 10 9 1 1 15 2 15 1 9 13 2
19 11 0 12 9 1 12 12 9 1 9 0 13 11 1 9 1 13 4 2
15 15 15 0 9 1 14 12 9 1 11 1 9 1 13 2
19 11 0 0 0 9 13 15 11 1 0 3 0 9 1 9 1 9 13 2
8 11 1 3 0 9 11 13 2
16 11 1 9 1 9 13 1 3 3 11 9 1 15 1 13 2
17 15 0 12 9 1 9 1 1 11 11 1 10 1 15 14 13 2
23 11 1 3 0 9 1 13 1 1 11 1 10 9 1 1 1 9 1 9 0 13 4 2
13 10 9 11 11 1 12 12 9 1 9 1 13 2
19 12 12 9 1 10 9 1 1 0 7 0 9 9 1 9 0 13 4 2
15 11 0 12 9 1 11 7 15 0 12 9 1 9 13 2
10 11 1 11 1 9 1 13 4 4 2
19 11 11 11 1 9 1 11 1 12 9 1 9 1 9 14 13 4 4 2
21 15 2 11 11 11 11 11 2 1 9 11 11 7 11 11 1 9 14 0 13 2
24 11 1 11 11 11 1 11 1 2 11 1 9 2 1 1 0 9 1 9 1 9 13 4 2
30 15 13 16 10 9 1 15 0 9 1 9 9 13 7 9 14 9 1 9 1 0 15 0 9 1 13 1 13 4 2
11 11 0 11 11 11 1 0 13 4 4 2
13 15 13 16 0 9 1 3 13 1 0 9 13 2
14 10 9 1 1 10 9 1 9 1 13 1 9 13 2
24 15 10 9 1 9 1 9 13 4 13 2 11 1 9 1 1 15 10 9 13 1 9 13 2
16 11 1 9 1 13 13 4 0 9 1 15 1 0 9 13 2
19 12 0 9 1 9 1 9 1 11 12 9 1 9 1 0 13 4 4 2
13 15 1 0 11 11 11 2 11 2 1 9 13 2
16 11 1 10 9 1 13 2 15 0 7 0 13 4 4 4 2
12 9 14 9 1 1 15 9 0 13 4 4 2
23 15 10 0 9 15 9 1 0 9 13 7 9 1 9 9 13 4 14 0 13 4 4 2
17 11 1 13 2 9 9 11 7 11 1 9 1 9 13 4 4 2
20 11 1 11 1 10 9 1 9 9 1 9 1 1 12 12 0 9 0 13 2
74 15 10 9 1 1 9 1 9 13 2 9 1 9 1 0 9 9 2 9 7 9 2 9 7 9 1 9 2 0 9 1 9 13 1 1 9 9 1 9 9 1 9 2 0 7 0 9 1 1 9 2 11 11 11 1 9 2 11 1 9 7 11 1 9 1 1 0 0 9 1 9 0 13 2
31 11 1 1 11 11 1 9 13 4 9 9 1 0 12 9 1 1 0 12 0 9 1 11 11 1 14 0 13 4 4 2
15 15 1 11 11 2 11 11 7 11 11 1 9 13 4 2
15 7 11 1 0 9 11 11 15 9 0 13 1 0 13 2
20 16 9 1 13 9 1 11 1 9 1 9 1 9 13 1 9 13 4 4 2
13 7 15 14 15 0 9 8 0 14 13 4 4 2
18 11 11 1 9 13 4 11 9 1 1 11 1 9 9 1 13 4 2
10 15 1 14 15 13 1 15 9 13 2
15 10 9 1 0 9 11 11 7 9 11 11 14 0 13 2
14 9 1 9 1 1 15 0 9 1 9 14 13 4 2
19 9 9 1 1 1 0 11 11 1 1 11 11 1 3 9 13 4 4 2
12 0 9 9 11 11 3 9 13 1 0 13 2
16 11 1 11 11 1 0 0 9 1 1 1 0 13 4 4 2
27 11 11 1 11 11 11 1 9 1 11 11 11 2 11 2 1 9 13 1 11 1 9 1 9 13 4 2
29 16 15 14 13 16 10 9 1 9 1 12 0 9 0 13 4 4 4 7 15 0 12 14 9 1 13 14 4 2
33 11 11 11 1 0 13 4 1 0 9 1 1 1 9 9 1 11 11 11 11 1 13 16 10 9 1 1 0 9 1 9 13 2
7 9 9 1 9 1 13 2
14 10 9 1 0 13 2 13 0 9 0 13 4 4 2
40 10 9 1 9 1 1 11 11 11 1 9 1 9 0 13 4 15 13 16 10 9 15 0 13 15 9 9 1 9 13 13 4 7 15 9 14 13 4 4 2
23 11 1 11 9 11 11 1 11 1 0 11 11 11 1 9 1 12 0 9 1 9 13 2
21 0 9 1 12 0 9 1 0 13 4 4 2 7 12 9 0 9 1 14 13 2
23 11 9 1 9 1 1 2 9 1 13 4 16 9 1 9 1 15 9 14 13 4 4 2
40 15 13 16 0 12 9 1 11 1 9 9 1 9 9 13 1 11 11 11 11 1 9 1 14 13 4 2 7 11 11 1 9 11 11 11 1 9 1 13 2
23 16 2 9 1 10 0 9 1 0 13 4 4 15 11 1 0 9 11 11 9 14 13 2
27 9 11 1 12 0 9 13 7 11 1 15 11 1 9 13 4 4 10 9 15 11 11 14 13 4 4 2
13 9 1 1 2 10 9 1 9 13 4 4 4 2
11 9 1 0 9 1 9 13 4 4 4 2
10 3 10 9 11 11 11 1 1 13 2
32 11 1 11 11 9 1 9 13 1 1 11 11 11 11 11 11 11 1 11 1 15 14 9 1 9 1 9 1 9 13 4 2
14 11 1 9 1 0 9 13 7 15 1 3 9 13 2
14 10 9 1 11 11 1 9 1 11 0 9 13 4 2
45 11 11 11 11 2 11 2 1 9 9 11 11 1 9 1 9 1 13 16 9 1 9 9 9 1 9 13 1 1 9 1 0 9 1 11 1 9 1 9 13 1 9 13 4 2
37 0 13 16 11 1 11 1 12 0 9 1 13 1 14 3 11 1 12 9 9 1 0 13 4 11 1 9 1 9 9 9 1 3 9 13 4 2
19 15 13 4 16 15 1 9 9 9 0 9 1 1 12 9 13 4 4 2
24 16 2 11 1 13 16 2 11 1 9 1 15 3 10 0 13 16 15 0 9 1 13 4 2
34 0 9 1 13 1 9 10 9 1 0 9 0 13 4 4 16 9 1 1 11 1 13 4 4 9 9 1 9 15 14 13 4 4 4
34 15 3 13 16 2 0 11 11 11 1 9 13 1 9 10 0 9 1 9 13 4 15 9 1 0 13 1 1 0 9 13 4 4 2
20 11 11 1 11 11 11 1 11 11 11 1 11 1 12 0 9 1 0 13 2
13 11 9 11 11 1 11 11 11 11 9 13 4 2
31 11 9 11 11 11 2 0 9 11 11 7 11 1 11 9 9 11 11 11 1 12 9 1 9 1 0 9 9 13 4 2
12 10 9 1 12 9 9 1 14 0 13 4 2
23 9 0 11 11 1 11 1 11 11 1 11 11 1 9 1 0 9 1 9 11 1 13 2
15 15 9 1 11 11 1 9 1 0 9 1 0 9 13 2
21 11 1 12 9 1 9 1 0 9 1 9 1 9 1 0 9 1 3 9 13 2
22 15 13 16 0 9 1 12 9 9 13 9 1 9 1 9 1 0 9 0 13 4 2
13 11 1 10 9 1 9 9 7 9 9 9 13 2
13 0 9 7 9 11 11 1 14 0 9 13 4 2
14 9 0 14 13 1 1 15 9 1 0 14 13 4 2
12 15 1 1 15 9 11 11 1 9 9 13 2
21 0 11 9 11 11 1 11 11 11 2 12 12 9 7 9 9 2 9 13 4 2
17 12 0 9 1 14 0 2 12 12 9 7 9 9 2 13 4 2
31 9 13 1 1 11 9 11 11 2 11 9 11 11 2 11 9 11 11 2 11 9 11 11 7 11 9 11 11 0 13 2
17 15 1 9 1 12 0 11 9 2 9 2 1 14 9 13 4 2
34 15 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 11 2 11 11 7 11 11 11 0 13 2
31 10 9 1 0 9 11 11 2 11 11 2 11 11 7 11 11 1 14 9 13 4 4 2 7 15 9 1 0 14 13 2
24 11 11 11 11 11 2 11 2 1 0 11 7 11 1 9 11 1 9 14 1 9 13 4 2
15 10 9 1 12 12 1 10 9 2 9 9 13 4 4 2
17 7 9 0 9 1 9 11 7 11 2 11 1 1 9 0 13 2
19 11 9 1 13 16 10 9 1 1 12 12 12 12 9 1 9 13 4 2
14 10 9 9 13 1 9 1 12 9 1 9 13 4 2
20 11 9 11 11 1 13 16 10 9 9 1 13 1 9 1 9 13 4 4 2
15 9 1 10 9 0 7 0 9 1 1 0 9 13 4 2
11 10 9 9 9 9 1 14 13 4 4 2
14 9 13 1 1 9 1 10 9 9 1 9 13 4 2
21 15 9 1 9 9 9 13 4 4 2 15 9 1 9 9 1 9 13 4 4 2
22 11 11 1 13 13 16 0 9 1 1 15 10 9 9 7 0 9 1 9 13 4 2
33 0 3 11 11 11 11 11 1 13 16 16 0 9 1 11 11 1 9 1 9 13 1 9 13 4 2 16 11 11 3 9 13 2
27 11 9 2 11 2 11 2 11 2 1 0 9 13 9 1 9 15 9 9 1 9 13 1 1 13 4 2
11 15 1 15 9 9 1 14 0 13 4 2
28 3 2 0 9 13 9 2 11 2 11 2 1 0 13 1 3 0 9 1 1 15 9 9 1 9 13 4 2
17 7 15 15 13 4 9 13 4 16 14 12 9 0 13 4 4 2
31 11 1 9 1 9 13 1 11 11 1 9 1 9 1 0 9 9 7 15 1 9 7 9 13 1 9 1 9 13 4 2
21 10 9 10 9 13 15 0 9 1 0 11 9 1 13 9 1 9 1 9 13 2
11 10 9 0 9 1 1 10 3 0 13 2
14 9 1 13 1 3 15 1 13 9 14 0 13 4 2
5 14 3 15 13 2
17 3 14 0 9 1 9 13 4 4 7 9 1 9 9 13 4 2
13 9 1 1 0 9 1 14 9 9 0 13 4 2
43 10 9 14 1 15 14 9 14 13 16 0 9 1 9 13 14 11 11 11 1 9 1 9 1 9 13 4 7 9 1 15 9 13 9 1 3 0 9 1 9 13 4 2
25 15 1 9 9 1 0 2 0 13 1 1 0 9 1 12 12 9 1 10 9 13 4 4 4 2
22 7 0 9 1 1 9 13 15 9 9 1 10 0 9 1 14 0 9 13 4 4 2
26 9 1 11 1 10 9 1 9 13 16 11 11 11 1 1 11 2 11 11 1 9 0 13 4 4 2
30 11 2 11 2 11 11 11 11 11 11 11 1 9 1 1 9 1 13 16 11 2 11 11 1 9 0 13 4 4 2
18 15 13 16 11 11 11 1 1 15 1 10 12 9 9 13 4 4 2
30 12 9 1 9 1 15 13 16 10 9 1 1 13 4 4 9 1 9 13 1 1 9 1 9 0 9 1 0 13 2
18 0 11 11 11 11 1 9 1 9 11 1 0 9 9 13 4 4 2
21 3 11 7 11 11 1 9 1 14 9 10 15 13 16 9 14 9 14 13 4 2
10 11 11 9 1 14 11 13 4 4 2
26 9 9 7 9 9 9 1 10 9 1 1 0 13 4 4 2 15 11 1 13 4 7 15 15 13 2
13 15 15 13 1 9 11 11 11 1 13 4 4 2
19 7 15 14 9 1 0 11 11 11 1 0 7 0 9 9 1 9 13 2
14 0 9 1 0 12 9 1 9 1 9 13 4 4 2
13 10 9 1 11 11 11 1 3 9 13 4 4 2
18 15 1 15 14 9 1 9 13 7 9 1 1 0 9 13 4 4 2
14 12 9 1 9 1 1 0 9 0 13 4 4 4 2
27 11 9 1 9 1 1 9 13 1 9 1 13 4 16 15 15 9 9 1 9 12 12 9 14 13 4 2
10 15 15 15 9 1 9 14 13 4 2
8 16 9 9 12 9 9 13 2
18 11 1 9 10 9 1 13 13 2 15 0 9 1 1 3 0 13 2
13 11 11 1 0 9 1 1 11 1 11 13 4 2
18 11 11 1 9 1 9 9 1 1 9 9 1 0 9 1 9 13 2
15 15 9 9 2 11 2 9 7 11 11 1 9 0 13 2
23 10 0 9 1 10 9 1 14 9 13 2 15 0 9 1 0 9 1 9 13 4 4 2
12 11 1 14 10 9 7 12 9 13 4 4 2
11 11 10 0 9 1 14 11 1 9 13 2
22 16 2 0 9 1 10 9 7 9 1 9 14 13 2 15 1 15 11 1 9 13 2
19 15 11 1 9 1 9 11 1 13 4 4 15 10 9 12 9 0 13 2
10 15 12 9 1 0 9 14 0 13 2
15 10 9 1 15 1 11 7 11 1 10 9 9 13 4 2
37 11 1 12 0 9 11 11 7 11 11 1 0 9 1 15 15 1 1 9 2 9 1 0 11 11 11 1 11 1 12 9 1 3 3 9 13 2
21 11 9 9 1 13 1 3 11 11 11 1 10 9 1 9 13 1 9 13 4 2
27 11 1 11 11 1 12 9 1 3 3 13 15 15 1 1 9 13 7 9 2 9 1 13 1 9 13 2
22 11 11 11 1 11 1 10 9 1 9 1 13 1 9 1 1 11 1 10 9 13 2
26 0 9 12 0 9 1 9 1 13 4 15 15 1 1 13 4 9 1 9 13 1 9 13 4 4 2
23 0 9 9 11 11 11 1 14 11 1 9 1 11 11 1 11 11 11 11 1 9 13 2
36 11 1 13 13 16 0 9 1 1 11 1 12 0 9 1 15 15 1 1 9 2 9 13 1 1 11 9 1 9 1 0 9 13 4 4 2
24 9 1 9 11 11 1 13 16 10 9 1 9 1 11 1 0 9 1 9 1 13 4 4 2
27 11 11 1 9 1 1 9 1 9 13 4 11 11 1 13 16 15 11 1 11 1 13 9 0 13 4 2
15 7 11 9 1 9 1 1 9 1 9 13 14 13 4 2
26 15 1 11 1 10 9 1 0 13 4 13 16 15 11 1 14 0 13 4 4 11 1 14 13 4 2
32 11 1 11 7 11 11 11 1 9 1 15 1 9 13 7 15 9 1 0 13 7 9 9 1 9 9 13 1 9 13 4 2
16 11 1 13 16 10 10 9 13 4 15 15 0 13 4 4 2
19 0 3 11 1 11 1 9 2 9 7 9 1 9 13 1 9 13 4 2
47 11 11 11 2 11 2 1 9 1 10 9 1 9 13 4 16 15 11 11 11 11 2 11 2 1 0 9 7 9 9 9 1 1 0 12 7 12 9 9 1 9 13 1 9 13 4 2
33 11 9 11 11 1 11 1 13 16 15 11 1 11 1 9 11 11 1 0 9 1 12 7 12 9 9 1 13 1 9 13 4 2
21 0 9 11 11 1 12 9 7 12 9 9 9 9 13 11 9 1 13 4 4 2
23 10 9 1 9 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 1 13 4 2
13 3 11 11 1 9 1 9 1 13 10 0 13 2
12 11 1 9 1 1 11 1 3 9 13 4 2
21 11 9 1 9 13 16 15 9 1 9 1 10 9 1 0 9 13 4 4 4 2
19 15 1 13 4 4 4 16 11 1 11 1 11 11 11 1 14 9 13 2
31 10 9 1 0 9 1 9 13 4 4 4 7 11 9 1 11 1 9 9 9 1 9 1 9 1 0 13 1 9 13 2
12 16 11 1 10 12 9 9 1 9 14 13 2
15 15 13 16 15 9 13 0 14 13 2 7 15 0 13 2
17 11 11 11 1 14 9 1 11 1 9 14 13 1 9 13 4 2
35 11 11 1 3 14 13 2 7 15 9 15 13 16 0 9 10 9 1 9 14 13 13 2 15 1 10 0 9 1 0 9 13 4 4 2
27 15 13 16 15 0 9 1 1 1 9 13 7 0 9 1 1 1 11 1 15 9 1 0 13 4 4 2
15 15 11 1 9 13 1 3 15 0 13 1 9 13 4 2
20 15 0 9 13 16 15 10 9 1 9 13 13 4 7 15 9 0 14 13 2
11 11 1 11 1 1 3 15 9 14 13 2
26 7 11 1 11 1 13 11 11 11 2 11 2 1 9 1 15 0 9 1 1 1 9 13 4 4 2
20 11 1 13 16 15 3 14 11 11 7 11 11 11 9 11 11 1 9 13 2
17 11 7 11 1 9 14 1 11 1 9 9 9 1 9 13 4 2
20 15 9 13 13 16 11 1 0 9 0 13 7 15 9 1 15 9 14 13 2
23 11 9 1 9 1 9 13 1 3 11 11 1 9 1 1 11 1 12 10 0 9 13 2
31 11 11 1 1 1 9 0 9 1 13 4 16 9 1 9 1 11 11 1 9 9 1 9 1 13 1 9 13 4 4 2
20 11 11 1 12 9 9 9 1 9 1 1 0 9 1 11 11 14 9 13 2
43 0 3 9 10 9 1 13 4 4 16 11 11 1 9 7 9 9 11 11 1 0 9 9 1 12 12 9 1 9 1 1 1 11 11 1 0 0 9 1 0 13 4 2
28 9 13 4 4 16 11 11 1 9 1 11 11 1 15 1 9 13 1 3 0 9 1 14 9 13 4 4 2
25 9 1 13 16 11 11 1 11 11 1 12 9 1 11 11 7 11 11 1 9 1 0 13 4 2
20 15 0 9 1 11 1 12 9 1 9 9 1 1 1 0 9 13 4 4 2
33 0 13 16 10 9 13 16 11 11 1 12 12 9 1 11 11 11 1 1 11 11 1 11 1 9 1 13 14 9 13 4 4 2
13 13 4 16 12 9 1 9 14 10 9 1 13 2
32 9 13 4 16 11 11 1 0 13 1 3 11 11 2 11 1 11 1 11 11 1 1 12 12 9 1 9 9 0 13 4 2
16 10 9 1 11 11 1 9 7 9 9 11 11 14 0 13 2
22 9 1 1 10 9 1 14 1 11 1 11 7 12 9 1 1 3 14 9 13 4 2
25 15 11 7 11 11 11 11 11 1 11 1 11 11 1 12 12 9 9 2 9 1 9 13 4 2
21 0 9 1 9 1 13 9 1 0 9 1 12 11 9 10 9 1 13 4 4 2
10 10 9 11 1 12 9 1 13 4 2
33 0 9 11 2 11 15 1 0 9 1 9 2 9 1 13 4 4 7 15 9 9 1 0 10 9 2 9 9 1 13 4 4 2
9 10 9 0 10 9 1 0 13 2
18 15 10 0 9 9 1 9 1 10 9 9 1 0 13 1 0 13 2
35 0 9 13 1 1 11 2 11 13 4 1 10 9 15 1 15 9 1 0 14 13 2 15 1 14 15 15 9 2 9 9 14 13 4 2
22 9 1 9 13 1 1 9 1 9 10 9 1 13 4 4 16 15 1 9 14 13 2
49 15 9 1 10 9 1 0 13 1 13 1 3 0 9 13 16 15 15 1 15 9 2 9 9 14 13 2 15 1 14 15 0 9 1 15 9 14 13 16 15 15 13 4 7 9 1 15 13 2
23 9 1 11 11 1 1 11 1 11 11 11 11 11 1 0 11 11 1 9 14 13 4 2
27 11 11 11 11 11 11 1 1 1 9 9 13 4 1 9 1 9 1 15 14 9 0 14 13 4 4 2
31 16 9 1 0 11 2 15 9 11 11 7 0 9 1 11 1 0 11 11 2 11 11 7 9 9 1 14 9 13 4 2
15 11 11 1 15 0 9 1 9 1 9 0 13 4 4 2
22 15 10 0 9 1 1 2 9 11 1 9 1 10 0 9 1 14 0 13 4 4 2
14 15 12 0 9 13 11 11 11 11 11 11 11 11 2
6 15 3 0 9 13 2
14 15 1 11 1 0 0 11 11 14 9 1 0 13 2
14 0 0 9 1 9 1 9 1 9 0 13 4 4 2
22 11 1 11 11 1 9 1 1 11 11 9 1 12 9 1 1 0 13 4 4 4 2
8 16 15 9 9 13 4 4 2
27 10 9 11 9 1 0 9 1 9 13 1 11 7 11 11 11 2 11 2 1 9 1 0 9 1 13 2
33 9 1 0 13 13 11 11 1 9 9 11 11 11 1 9 1 9 1 13 16 9 1 9 11 7 11 1 9 9 1 13 4 2
17 15 15 12 9 1 1 0 9 9 1 9 13 1 9 13 4 2
23 16 15 13 16 9 1 9 1 9 1 11 9 1 0 9 1 1 1 15 9 14 13 2
13 10 9 1 11 7 11 1 12 9 1 9 13 2
23 11 1 11 11 1 13 16 9 1 0 9 12 9 1 1 0 9 9 1 0 13 4 2
20 11 1 11 11 1 13 16 9 1 11 9 1 9 1 13 15 9 14 13 2
28 11 1 13 16 11 1 0 13 1 10 0 9 13 15 11 2 11 2 11 7 0 9 1 9 1 9 13 2
23 0 9 1 1 0 9 11 1 9 9 1 0 0 9 1 9 1 9 9 1 9 13 2
22 9 1 11 11 11 1 9 11 11 1 11 1 9 1 1 10 9 1 9 13 4 2
38 15 13 4 16 15 9 13 16 3 0 9 1 10 9 1 9 0 13 4 2 16 9 1 13 11 0 9 1 0 13 7 9 0 9 1 9 13 2
30 11 1 13 4 16 0 9 1 0 9 1 0 9 14 13 2 16 15 1 10 9 1 9 1 14 9 13 4 4 2
18 9 9 1 3 0 9 13 4 4 1 9 1 13 1 0 13 4 2
25 15 13 16 3 10 9 0 9 1 0 9 1 13 4 2 16 9 9 1 9 1 15 0 13 2
22 11 1 13 16 9 1 0 9 1 9 1 0 9 1 0 9 1 13 15 9 13 2
23 15 10 9 1 9 13 2 15 10 9 1 9 1 9 1 3 0 9 1 0 13 4 2
28 15 13 16 10 9 1 13 13 16 10 9 1 9 1 0 9 7 15 0 9 1 9 1 9 13 4 4 2
27 15 1 9 9 7 9 1 7 9 1 1 15 9 0 0 9 13 4 15 15 0 9 1 9 13 4 2
47 15 13 16 11 1 9 1 9 1 0 9 1 0 10 9 13 4 1 0 9 1 9 1 9 13 4 2 7 0 10 9 1 9 1 9 1 0 13 1 1 9 13 9 13 4 4 2
27 11 15 11 9 1 1 9 7 9 1 9 2 0 9 1 9 2 0 0 9 7 0 0 9 1 13 2
38 11 9 11 7 12 0 9 1 1 11 9 0 13 1 11 11 1 9 1 9 1 9 13 4 0 9 1 11 1 15 9 11 11 1 13 4 4 2
29 0 9 11 1 9 1 9 13 16 15 1 9 9 1 9 1 9 14 13 2 7 15 9 1 9 0 13 4 2
28 15 1 11 11 1 11 9 11 11 1 9 9 1 1 1 0 9 1 9 13 1 9 1 9 0 13 4 2
40 7 11 1 9 1 9 1 1 9 9 1 9 11 11 7 11 11 11 1 11 1 11 11 1 1 9 0 13 11 1 9 1 0 9 1 9 1 9 13 2
8 11 10 9 9 9 1 13 2
14 0 9 1 15 9 1 11 11 11 11 1 9 13 2
34 9 1 13 13 16 9 1 9 7 0 7 0 9 1 13 0 9 1 1 9 1 0 11 1 9 1 1 1 14 13 4 4 4 2
43 11 1 11 11 11 1 11 1 11 9 1 9 0 9 1 0 9 1 3 0 13 1 9 13 4 7 9 1 14 9 1 9 9 1 0 9 1 0 13 1 13 4 2
43 11 1 9 11 11 11 1 0 9 1 9 1 9 9 9 13 1 9 13 4 7 11 1 11 9 1 9 9 1 13 4 9 1 0 9 1 12 9 13 1 9 13 2
16 11 9 1 11 9 1 9 13 4 1 12 9 13 4 4 2
33 11 11 9 1 11 1 11 7 11 1 9 1 1 9 1 9 1 1 1 12 9 1 15 9 1 9 1 9 13 1 9 13 2
28 11 9 1 11 1 12 9 1 13 9 1 9 1 11 2 11 9 1 0 9 9 1 12 9 0 13 4 2
9 9 9 1 11 1 10 9 13 2
40 9 1 1 0 9 1 9 1 0 11 11 1 9 7 0 9 9 1 9 1 11 2 11 9 1 12 9 1 13 9 1 13 1 1 0 9 1 13 4 2
18 11 11 1 9 9 1 1 13 7 9 9 1 9 9 1 1 13 2
21 10 3 15 13 9 1 9 13 1 12 9 0 13 4 15 3 1 9 13 4 2
33 9 1 9 1 9 1 10 9 13 4 16 15 10 0 9 1 15 0 13 7 9 1 15 9 1 9 15 14 9 1 0 13 2
27 15 1 14 9 1 10 9 1 0 14 9 13 4 7 12 9 1 0 9 1 9 1 9 13 4 4 2
10 10 11 1 9 1 9 1 9 13 2
13 10 12 9 11 1 12 2 12 14 10 0 13 2
31 9 9 1 15 11 11 1 1 9 1 9 1 1 11 11 0 9 1 9 13 1 9 1 12 0 9 1 9 13 4 2
22 0 9 9 9 11 1 1 0 12 9 1 1 9 9 1 10 9 1 9 13 4 2
21 10 9 1 9 1 11 1 1 15 0 9 1 0 13 1 9 0 13 4 4 2
48 11 11 11 11 1 9 11 11 1 1 15 1 11 1 15 0 9 1 9 1 9 3 14 13 2 7 10 0 9 1 9 13 4 4 16 9 1 11 1 1 15 0 9 0 13 4 4 2
9 13 4 12 0 9 11 1 13 2
43 0 9 9 11 1 9 1 0 12 9 9 1 9 9 1 13 4 16 0 9 1 9 11 2 11 2 1 1 13 7 9 15 11 1 1 1 12 2 12 14 10 13 2
21 16 10 0 9 0 10 9 1 1 15 11 1 1 13 4 0 9 1 0 13 2
15 0 10 9 1 12 1 10 9 1 9 13 4 4 4 2
11 13 4 4 4 16 15 9 1 9 13 2
15 15 15 1 11 1 1 9 1 9 14 13 4 4 4 2
27 7 11 11 1 0 9 1 9 9 1 13 9 13 4 4 4 16 15 1 15 11 1 1 9 0 13 2
42 16 9 11 1 1 9 1 9 13 1 11 1 1 9 1 15 0 9 1 9 13 4 4 16 15 0 9 1 9 1 9 13 1 3 15 1 9 1 9 13 4 2
25 16 9 13 4 16 3 15 9 1 1 0 9 7 9 10 9 1 0 13 15 9 0 13 4 2
31 11 11 1 9 9 9 11 11 1 1 15 1 11 11 9 1 12 1 9 13 1 12 0 9 1 9 13 4 4 4 2
20 9 1 9 13 16 9 1 1 13 1 10 9 1 9 1 9 12 9 13 2
17 16 11 1 1 9 1 9 1 1 15 0 13 1 9 14 13 2
19 11 11 1 1 15 11 11 11 1 11 1 14 0 9 9 0 13 4 2
18 11 11 11 11 11 11 1 11 1 11 11 1 0 9 1 9 13 2
15 15 9 1 9 9 13 1 11 11 1 9 1 9 13 2
28 11 1 11 1 1 0 9 1 11 11 13 1 9 11 1 9 7 9 9 9 1 1 13 4 0 13 4 2
28 11 1 0 9 1 9 1 9 1 11 1 1 11 2 11 1 11 11 11 11 7 10 0 0 9 0 13 2
20 9 1 11 1 12 0 0 9 1 11 9 1 11 9 1 9 1 13 4 2
14 10 9 1 0 9 0 0 9 13 1 0 13 4 2
13 11 1 11 1 13 16 11 0 0 9 1 13 2
16 11 1 0 9 1 10 9 1 0 13 1 9 13 4 4 2
14 10 9 1 9 1 9 1 1 0 9 13 0 13 2
30 11 1 13 16 11 1 9 1 0 0 9 1 11 11 1 0 12 9 1 0 9 1 9 2 9 13 4 4 4 2
43 15 13 16 11 9 1 9 0 9 1 14 13 4 4 7 10 9 13 16 11 9 1 3 1 9 13 4 9 9 1 9 1 0 0 9 1 13 1 1 9 13 4 2
39 11 11 1 10 0 9 9 1 1 1 0 0 9 1 0 9 13 4 11 1 13 16 9 7 9 1 9 1 3 14 10 9 1 12 0 9 13 4 2
37 11 1 9 9 1 1 1 15 13 16 11 7 11 12 0 0 9 13 7 15 15 0 13 15 9 13 16 0 9 1 9 1 0 9 13 14 2
25 15 13 16 0 9 12 9 1 9 13 4 4 16 0 9 1 10 9 0 13 1 13 4 4 2
17 15 9 10 9 1 10 0 9 13 7 10 0 9 1 9 13 2
23 15 13 16 15 10 9 1 0 13 4 16 11 1 11 11 1 9 3 0 0 9 13 2
21 11 9 11 11 7 11 11 11 11 1 11 9 11 1 11 11 11 1 9 13 2
21 12 9 1 11 1 0 9 9 1 0 7 0 9 1 9 1 9 2 9 13 2
15 11 11 1 11 11 11 1 1 10 9 9 2 9 13 2
13 10 3 12 9 1 0 9 1 9 2 9 13 2
14 11 1 11 12 9 1 0 9 1 11 1 15 13 2
9 11 9 15 11 11 11 1 13 2
14 15 11 1 11 1 1 0 9 9 1 1 1 13 2
15 12 9 1 0 2 0 7 0 9 1 9 2 9 13 2
14 11 1 1 9 9 9 9 1 1 1 14 9 13 2
12 11 9 11 11 14 11 1 0 11 1 13 2
20 9 9 1 9 1 1 11 11 1 11 9 1 9 9 1 9 1 9 13 2
14 9 1 0 9 9 1 9 1 9 13 1 1 13 2
18 11 11 1 0 9 1 13 4 16 14 12 9 0 9 9 1 13 2
12 15 1 0 9 11 11 1 11 9 1 13 2
12 11 1 12 9 1 9 1 9 13 4 4 2
17 10 9 9 14 1 13 9 9 9 1 9 1 0 13 4 4 2
21 9 1 13 4 4 16 9 1 0 9 1 1 10 9 9 1 13 1 0 13 2
23 9 1 9 1 13 9 13 4 4 10 9 1 15 0 13 4 4 9 13 4 4 4 2
16 9 1 13 1 3 15 11 11 1 0 9 11 1 13 4 2
8 15 10 0 9 13 4 4 2
14 9 7 9 9 1 15 1 1 0 13 4 4 4 2
24 11 9 9 1 9 1 1 14 11 1 0 0 9 1 3 13 1 0 9 9 13 4 4 2
27 11 1 11 11 11 1 0 13 4 4 16 15 0 9 1 9 1 0 9 1 1 1 0 9 13 4 2
14 11 1 13 11 1 14 11 1 9 0 13 4 4 2
34 11 1 13 13 16 16 0 9 1 0 9 11 11 11 1 9 1 9 13 1 9 14 13 16 15 0 9 1 0 13 4 4 4 2
25 11 1 11 1 3 13 1 10 9 1 1 11 0 11 1 9 1 15 9 13 1 0 14 13 2
15 7 2 11 1 0 9 9 15 10 9 1 0 14 13 2
15 15 9 13 16 10 9 1 9 9 9 1 1 13 4 2
22 15 1 2 9 3 1 1 11 14 11 1 1 15 9 13 1 1 14 0 14 13 2
26 9 9 7 11 1 9 11 11 0 13 4 4 16 11 1 11 7 11 1 1 12 1 9 13 4 2
19 9 1 12 0 9 1 1 2 11 1 11 11 1 1 9 13 4 4 2
35 11 9 11 11 11 1 9 1 14 9 1 1 1 9 13 4 7 0 9 11 1 13 1 10 9 9 1 12 9 1 1 13 4 4 2
25 9 1 1 11 1 11 1 1 9 13 1 9 1 0 9 1 15 9 13 1 14 9 13 4 2
13 11 1 15 1 15 1 1 15 9 14 13 4 2
18 11 1 0 9 1 9 14 13 1 1 9 11 1 0 13 4 4 2
21 9 9 11 11 9 1 11 1 9 1 3 13 1 10 9 0 9 13 4 4 2
31 0 11 1 9 1 13 16 11 11 1 0 9 9 1 13 4 2 16 9 1 9 1 11 11 1 13 1 9 13 4 2
27 11 1 11 11 11 1 13 16 9 9 1 14 13 14 15 9 1 9 7 9 9 13 1 1 3 13 2
12 9 9 1 9 13 0 13 9 1 13 4 2
18 0 0 9 1 9 1 11 1 15 9 1 0 13 4 10 9 13 2
29 11 1 11 11 11 11 11 1 9 9 1 9 9 1 11 11 1 13 16 9 9 1 13 4 9 13 4 4 2
19 11 1 13 16 15 15 9 1 14 9 1 9 7 9 9 13 4 4 2
14 7 10 9 1 13 13 16 9 1 15 9 14 13 2
20 15 13 16 15 10 9 1 9 13 4 15 9 1 1 1 15 9 14 13 2
15 11 1 13 16 11 11 10 0 9 1 9 13 4 4 2
15 11 1 13 16 11 9 1 13 9 1 15 9 14 13 2
23 15 0 13 16 15 1 9 1 9 13 15 1 11 9 7 9 1 10 9 13 4 4 2
58 0 9 1 0 0 9 2 11 2 1 0 9 1 9 1 9 13 1 1 11 1 9 1 9 1 9 13 4 1 1 11 11 11 11 1 11 1 13 16 9 1 9 1 11 11 1 9 1 0 13 1 10 9 13 4 4 4 2
30 11 1 13 16 11 1 0 9 0 13 7 10 9 9 1 13 4 0 9 1 0 13 1 9 1 13 4 4 4 2
37 15 9 1 13 0 9 9 1 0 13 4 11 1 9 13 16 0 0 9 1 0 13 1 9 0 13 7 15 1 0 9 1 9 13 4 4 2
24 11 11 1 10 9 1 14 9 13 16 9 9 7 9 1 1 0 9 1 9 7 9 13 2
43 11 11 1 9 1 13 4 16 15 1 12 0 0 9 1 9 1 0 13 3 14 0 13 2 16 9 11 2 11 1 9 2 9 1 0 9 1 9 1 1 13 4 2
18 15 1 9 1 9 9 1 13 4 1 1 15 13 3 14 0 13 2
21 11 11 1 9 9 1 13 16 11 1 9 11 11 11 2 11 2 1 13 4 2
25 15 1 14 15 13 16 11 0 9 1 0 0 13 1 1 0 9 9 1 0 13 1 0 13 2
37 11 11 1 10 9 9 1 13 0 9 1 11 1 9 1 9 1 9 13 1 1 11 1 9 1 9 13 1 9 13 1 12 9 1 13 4 2
40 0 0 9 1 11 11 1 9 13 1 0 9 11 11 11 2 11 2 1 9 1 0 11 11 1 10 9 1 9 9 7 9 1 9 13 1 9 13 4 2
33 11 11 11 1 1 11 9 1 13 12 0 9 1 9 1 13 16 11 11 9 1 1 0 9 9 0 13 1 9 13 4 4 2
16 0 12 9 1 1 9 1 9 1 0 9 9 13 4 4 2
29 9 1 13 16 16 15 9 13 16 13 16 11 11 7 0 15 0 9 1 1 13 4 9 9 1 0 14 13 2
10 15 10 9 13 15 1 15 9 13 2
10 0 13 16 9 1 9 11 13 4 2
9 10 9 11 11 11 1 9 13 2
16 0 0 9 1 0 9 9 7 11 1 9 3 0 0 13 2
24 3 11 0 0 9 1 0 9 2 9 13 4 2 3 9 9 1 9 1 9 13 4 4 2
18 9 1 13 4 16 11 1 11 1 13 1 9 1 0 9 13 4 2
10 10 9 1 0 10 9 1 9 13 2
18 16 0 9 1 10 9 1 1 1 0 9 13 1 9 13 4 4 2
41 11 1 11 1 9 2 9 7 9 2 9 0 9 13 1 9 1 9 0 13 4 9 1 13 16 11 11 0 9 1 13 9 1 14 9 2 9 13 4 4 2
17 11 1 11 2 11 7 11 1 3 0 9 13 1 9 13 4 2
12 0 9 1 10 9 1 9 13 4 4 4 2
24 11 11 10 15 14 9 1 0 9 1 0 0 9 1 9 7 9 2 9 1 0 9 13 2
17 11 1 11 1 12 9 9 9 1 10 14 10 12 9 13 4 2
15 9 11 1 9 1 11 11 1 12 0 9 1 13 4 2
10 9 1 1 15 15 9 13 4 4 2
26 11 11 2 11 11 11 1 9 11 11 11 11 1 11 11 1 12 9 1 11 1 9 13 4 4 2
13 9 1 1 2 15 10 9 1 9 13 4 4 2
15 16 9 1 15 1 13 12 0 9 1 0 13 4 4 2
39 0 9 1 9 11 1 0 0 9 1 9 13 4 11 11 1 11 11 1 9 11 11 1 13 16 15 0 14 13 16 13 1 9 1 0 9 13 4 2
37 0 9 1 1 2 11 1 11 11 1 13 0 9 11 11 11 11 1 0 9 13 7 9 9 9 7 0 9 1 9 1 15 14 9 13 4 2
35 11 11 11 11 2 11 2 1 0 9 1 15 9 1 10 9 0 13 1 1 9 1 11 11 11 2 11 2 1 9 1 9 13 4 2
31 11 1 9 11 11 11 1 11 1 13 16 9 9 1 9 1 9 1 9 1 12 14 9 1 10 9 1 9 13 4 2
41 11 1 11 11 11 11 11 11 1 11 1 13 16 10 9 1 9 9 13 4 15 1 9 1 9 2 9 2 9 2 9 7 9 0 9 1 9 13 4 4 2
18 15 13 16 11 1 11 1 0 9 1 10 9 1 0 9 13 4 2
13 10 9 1 9 11 1 11 11 11 11 1 13 2
27 11 1 11 1 13 16 16 15 9 9 7 0 9 0 13 4 16 11 10 9 1 9 13 1 0 13 2
43 0 9 11 7 11 0 9 1 0 9 1 15 13 16 15 9 1 9 1 0 9 0 13 7 15 0 13 1 0 9 13 4 4 16 15 0 9 9 14 13 4 4 2
33 9 9 1 9 1 13 9 9 11 11 11 1 11 9 1 2 11 11 2 1 1 13 1 3 15 15 11 1 11 9 1 13 2
40 9 9 1 13 1 12 0 9 7 12 9 13 1 3 16 15 11 1 15 9 9 1 9 1 9 13 4 9 1 9 11 11 1 9 13 1 9 13 4 2
31 11 1 15 11 11 11 1 13 16 15 11 11 1 1 11 1 11 9 1 12 0 9 2 9 13 11 11 1 9 13 2
37 11 1 1 13 15 9 14 0 13 1 9 1 9 13 4 11 1 13 16 10 9 15 0 9 1 1 15 9 1 0 13 1 9 13 4 4 2
21 15 10 9 13 15 15 1 10 9 1 9 1 9 7 0 9 1 13 13 4 2
34 15 13 16 11 1 9 9 1 9 1 1 13 7 9 0 13 1 13 9 1 1 0 12 9 1 15 12 0 9 9 1 13 4 2
27 16 11 1 13 13 16 12 0 9 9 7 12 9 13 1 3 15 15 15 9 9 1 0 13 13 4 2
16 15 11 11 1 15 9 1 9 3 14 9 13 1 9 13 2
23 11 9 1 9 13 15 9 2 9 1 9 13 1 3 15 11 1 11 1 9 13 4 2
34 11 11 1 9 1 13 10 9 1 11 9 2 3 9 9 11 11 11 7 11 11 1 0 9 1 0 13 1 9 9 13 4 4 2
21 12 1 12 12 1 9 1 10 9 1 9 1 12 9 1 9 0 13 4 4 2
9 10 9 1 12 0 9 13 4 2
14 11 1 13 16 15 15 0 2 0 9 14 13 13 2
20 15 9 1 13 14 0 9 1 12 9 9 9 1 0 2 0 9 13 4 2
31 12 9 9 9 13 4 9 1 9 2 9 1 9 2 9 9 2 9 9 2 9 9 7 0 9 14 1 9 13 4 2
22 11 11 1 13 4 12 9 1 11 11 1 12 0 9 7 12 0 9 9 14 13 2
19 13 4 9 1 10 9 11 1 1 11 1 9 9 9 1 9 14 13 2
10 10 9 1 12 9 1 9 13 4 2
18 3 2 11 9 11 1 11 1 0 11 9 1 12 9 0 13 4 2
31 9 9 1 1 11 9 11 9 1 11 1 1 11 7 0 9 1 0 9 1 9 1 9 11 9 11 11 1 13 4 2
9 15 11 11 9 1 9 9 13 2
5 15 0 9 13 2
27 7 11 9 1 11 1 11 2 11 9 1 1 9 1 1 0 11 9 11 11 11 14 11 1 13 4 2
8 15 11 9 1 13 1 13 2
27 3 2 11 9 1 11 1 11 9 1 11 2 11 7 11 1 1 9 1 9 1 9 1 0 9 13 2
12 10 3 12 11 7 12 9 1 9 13 4 2
30 10 9 1 9 11 1 9 11 11 7 9 9 9 9 1 9 11 11 7 11 2 11 1 11 1 1 1 13 4 2
29 11 11 1 11 1 9 9 1 9 1 13 4 9 1 11 9 11 11 1 2 9 1 9 1 9 2 9 13 2
19 15 13 16 11 1 11 9 1 9 0 0 11 9 1 1 0 14 13 2
11 15 15 9 1 0 9 1 13 4 4 2
22 9 1 14 3 3 15 9 13 16 15 14 10 9 15 9 13 1 2 9 2 13 2
23 15 15 9 9 9 11 11 11 1 10 9 1 9 1 9 13 1 9 1 1 0 13 2
53 11 1 11 11 11 1 9 1 9 1 11 11 1 13 16 11 1 9 9 1 12 12 9 1 9 13 4 9 1 12 9 13 1 1 13 7 15 0 13 4 16 9 0 9 9 1 9 1 1 0 14 13 2
15 15 11 1 9 1 0 11 1 9 1 3 0 9 13 2
14 15 13 16 9 1 10 9 13 4 15 3 10 13 2
12 9 1 13 16 15 0 9 1 9 14 13 2
18 11 9 1 1 11 11 11 9 11 11 11 7 11 11 11 14 13 2
10 11 11 1 0 3 9 1 9 13 2
7 15 15 9 9 13 4 2
26 9 9 1 9 1 9 1 0 9 13 4 9 9 1 11 1 9 13 9 1 12 9 1 13 4 2
13 10 9 1 9 9 1 12 9 14 0 13 4 2
21 15 1 11 9 1 9 1 9 1 9 9 13 9 1 12 9 1 0 13 4 2
19 9 1 1 11 9 1 11 9 1 9 1 9 1 9 1 0 13 4 2
19 11 9 1 13 4 10 9 1 9 1 9 9 12 9 1 13 4 4 2
10 9 9 10 12 9 0 13 4 4 2
14 10 9 9 9 1 15 1 12 9 13 4 4 4 2
20 11 1 1 11 9 1 11 9 1 11 1 14 9 1 12 9 1 13 4 2
21 9 9 9 1 9 9 1 1 13 10 9 1 9 1 12 9 14 0 13 4 2
11 9 1 13 16 9 9 15 14 0 13 2
25 9 1 1 11 1 11 9 1 9 9 11 11 1 9 11 11 11 14 11 1 9 0 13 4 2
22 7 9 1 11 1 11 9 1 0 9 9 11 11 1 15 9 1 13 9 13 4 2
16 11 9 1 11 1 9 1 12 9 1 9 1 13 13 4 2
20 10 9 11 2 11 11 1 9 9 1 1 0 9 1 9 12 12 9 13 2
11 15 0 12 9 1 9 0 13 4 4 2
26 9 1 1 9 9 1 9 1 13 4 7 9 1 13 1 1 0 9 9 13 7 15 9 14 13 2
32 9 1 0 9 1 1 11 11 11 2 11 2 1 0 9 12 9 1 0 9 0 13 12 9 1 0 9 9 1 0 13 2
11 11 11 12 9 13 12 9 1 0 13 2
19 9 1 1 9 0 13 1 3 1 10 0 9 15 9 1 13 0 13 2
27 7 2 9 0 13 1 0 13 4 4 16 10 14 10 9 9 1 9 1 15 15 0 0 9 14 13 2
21 15 1 9 1 9 1 3 13 1 0 7 0 9 9 1 0 9 13 4 4 2
14 10 9 1 9 9 1 3 9 0 13 4 4 4 2
16 0 7 0 9 1 9 13 4 0 9 1 14 9 13 4 2
14 0 9 1 1 14 10 9 1 9 1 9 13 4 2
33 15 0 9 1 1 11 9 11 11 11 1 11 1 9 9 11 11 11 1 9 13 7 9 1 13 9 1 3 13 1 9 13 2
14 11 1 11 1 0 9 1 13 1 0 9 13 4 2
18 15 9 9 1 9 13 16 15 9 1 10 9 1 9 1 9 13 2
25 0 13 16 11 1 11 1 11 1 13 4 16 0 9 1 11 1 9 0 9 1 15 9 13 2
57 16 2 9 9 1 1 2 13 4 4 16 14 10 9 1 9 1 11 1 11 1 10 9 1 0 13 1 9 13 16 15 15 9 1 2 15 9 7 9 0 14 13 2 13 4 2 7 10 15 14 13 15 10 14 0 13 2
13 2 11 1 11 1 9 1 15 0 9 13 4 2
21 15 12 0 9 1 13 16 2 15 13 4 16 11 1 9 1 11 0 14 13 2
20 15 10 9 1 9 2 9 13 1 1 11 11 1 9 2 3 13 13 4 2
18 9 1 1 9 2 9 1 1 15 10 9 3 1 1 0 13 4 4
27 0 9 1 1 0 9 13 4 11 1 11 1 11 1 12 10 9 1 0 0 9 13 1 9 13 4 2
20 11 1 10 9 1 1 10 9 13 1 11 1 9 1 9 13 12 13 4 2
27 11 11 1 9 11 11 1 13 16 11 11 1 0 9 1 12 10 9 1 0 9 1 9 13 4 4 2
20 10 9 1 11 1 0 7 0 9 1 0 9 11 1 0 0 9 13 4 2
31 0 9 9 13 4 10 9 1 1 11 11 1 1 1 9 7 15 12 9 1 9 9 7 13 1 9 0 13 4 4 2
29 11 1 1 1 11 1 1 9 0 13 1 9 1 1 10 9 11 0 0 9 1 1 1 0 13 4 4 4 2
31 11 9 1 11 9 1 9 1 9 13 4 1 9 1 12 9 1 9 1 15 1 9 9 7 9 9 1 13 4 4 2
27 11 1 9 11 11 11 1 0 9 13 2 7 11 1 9 9 11 11 1 11 9 1 9 13 4 4 2
11 0 12 9 1 0 13 1 9 0 13 2
35 0 13 16 11 1 0 11 1 9 1 9 13 4 1 9 1 1 1 14 10 9 9 1 9 1 9 7 9 1 13 1 9 13 4 2
18 11 1 0 0 9 1 1 11 1 9 11 1 14 13 4 4 4 2
17 15 9 1 11 2 11 2 1 9 11 11 1 11 13 4 4 2
18 11 1 9 11 11 1 11 11 1 9 1 11 1 9 13 4 4 2
26 11 1 13 4 9 11 11 11 2 9 9 11 11 7 9 11 11 1 3 15 9 14 13 4 4 2
18 11 13 4 11 11 1 9 1 11 1 0 9 1 9 15 13 4 2
26 12 10 9 1 1 9 1 11 11 1 9 11 11 11 11 1 11 11 1 9 1 0 9 13 4 2
20 15 13 16 11 11 1 9 13 1 9 1 12 9 1 0 13 4 4 4 2
11 0 12 9 1 0 13 1 9 0 13 2
52 10 3 11 1 9 9 2 0 2 11 11 1 13 16 11 9 1 9 13 7 9 13 1 9 1 0 11 9 11 11 0 11 11 7 11 9 11 0 11 1 0 13 9 9 9 1 9 1 0 13 4 2
13 9 1 15 11 11 1 9 1 9 1 13 4 2
20 15 13 16 9 1 9 1 1 11 11 2 11 1 9 9 0 13 4 4 2
21 15 13 16 11 1 9 9 1 9 9 9 1 1 12 0 9 0 13 4 4 2
18 10 9 9 1 1 11 11 0 11 7 11 1 9 1 13 4 4 2
36 11 1 11 11 1 12 9 1 9 9 13 1 9 9 1 9 1 9 13 4 11 9 11 11 11 1 13 16 15 9 2 9 1 1 0 13
41 11 1 12 0 9 1 9 13 4 11 11 11 11 1 9 1 13 9 1 13 16 15 11 11 1 9 1 12 9 1 9 13 1 9 1 9 1 9 13 4 2
9 11 9 1 1 3 0 13 4 2
35 16 2 11 1 15 14 13 16 0 13 16 9 1 9 1 9 13 1 3 11 11 1 9 13 4 11 1 0 9 1 14 9 13 4 2
17 15 13 16 11 1 1 9 9 2 9 1 9 1 0 13 4 2
23 15 13 16 11 11 1 0 9 1 0 7 0 9 1 9 13 1 1 0 9 0 13 2
17 11 1 13 16 9 1 0 7 0 9 1 1 0 9 13 4 2
44 11 11 7 11 1 9 1 9 1 0 9 1 1 1 0 11 1 10 9 1 9 1 9 13 4 4 3 11 7 11 1 0 9 1 9 13 1 9 0 2 0 13 4 2
17 9 1 9 1 1 1 11 7 11 1 12 9 1 9 13 4 2
35 7 0 9 1 11 1 9 13 4 1 1 9 9 1 12 9 9 10 8 13 4 2 7 9 1 1 1 9 9 1 9 0 13 4 2
24 11 2 11 11 11 1 9 1 13 9 9 1 1 9 9 9 0 9 1 0 13 4 4 2
23 9 9 1 1 11 1 9 1 1 1 9 9 1 12 9 10 12 9 9 8 13 4 2
15 7 0 9 9 13 1 9 1 0 9 1 9 13 4 2
12 9 1 1 9 9 13 12 9 0 13 4 2
26 15 1 0 9 1 15 9 14 13 7 10 9 1 9 1 0 13 4 7 15 9 1 0 13 4 2
18 0 9 1 1 11 1 9 9 1 12 9 10 12 9 8 13 4 2
7 9 1 12 9 9 13 2
22 11 1 12 9 9 8 13 4 16 0 9 9 1 12 9 13 12 9 9 13 4 2
25 11 1 13 9 1 1 9 1 9 9 9 1 11 1 11 11 9 1 12 9 1 9 13 13 2
15 7 11 1 12 0 9 1 9 1 1 1 9 13 4 2
25 11 2 11 1 10 9 1 0 9 1 1 9 1 9 1 9 13 1 9 9 1 13 4 4 2
28 9 1 1 9 1 1 9 1 9 1 0 9 1 9 13 4 4 7 11 1 11 11 11 1 12 9 13 2
31 9 1 1 11 2 11 11 11 1 13 12 1 10 9 1 9 1 9 1 1 1 3 2 3 13 1 9 13 4 4 2
42 11 11 1 9 1 9 1 9 1 14 9 1 13 4 10 0 0 9 1 9 1 1 1 12 0 9 1 11 11 1 12 9 1 9 1 0 9 0 13 1 13 2
30 16 11 1 11 1 9 1 13 16 15 9 1 0 9 1 0 9 9 1 1 11 11 11 13 1 9 13 4 4 2
34 11 11 1 1 1 9 1 9 9 9 11 11 1 9 13 16 0 9 1 0 9 1 1 12 11 11 11 13 15 1 9 9 13 2
6 15 1 9 13 4 2
38 11 11 11 1 9 1 0 9 1 11 11 11 2 11 11 11 11 2 11 11 11 7 11 11 11 1 10 0 9 1 9 13 9 0 13 4 4 2
62 9 9 11 11 11 2 9 11 11 11 2 9 11 11 11 7 9 11 11 11 1 9 1 12 9 9 11 11 11 11 1 9 9 1 9 13 1 1 11 11 1 13 16 12 9 1 0 9 9 1 0 13 7 12 9 1 9 1 9 13 4 2
31 9 9 1 9 13 4 4 16 0 0 9 1 14 13 4 0 9 1 9 1 13 4 16 15 9 9 1 1 0 13 2
39 11 11 1 12 0 9 1 1 9 13 15 9 13 1 12 9 1 11 11 11 0 13 13 4 16 15 0 9 1 1 9 9 1 9 15 14 13 4 2
40 9 9 1 10 9 1 0 14 0 9 13 4 9 9 1 9 13 4 7 11 11 1 11 11 1 9 9 1 9 1 9 9 1 9 1 0 13 4 4 2
25 11 11 1 9 1 9 13 1 11 11 1 0 9 9 1 9 1 0 9 1 9 0 13 4 2
11 9 10 9 11 1 9 9 1 0 13 2
21 11 11 11 1 9 1 9 13 4 16 11 9 15 9 1 9 1 1 0 13 2
15 0 9 1 9 1 1 0 9 1 14 9 0 9 13 2
17 11 1 10 9 1 12 0 9 0 13 4 1 9 14 13 4 2
23 3 2 11 11 11 11 11 11 1 9 1 15 7 9 1 1 9 0 13 1 9 13 2
18 15 13 16 0 9 9 1 15 15 9 1 15 9 1 9 14 13 2
20 9 1 9 7 9 1 9 11 11 11 1 1 1 12 9 1 9 13 4 2
32 9 1 9 13 4 11 11 11 1 13 16 11 9 1 9 1 1 9 1 0 7 0 9 1 0 13 1 9 1 13 4 2
12 15 11 1 14 9 1 0 9 13 4 4 2
23 11 1 13 16 15 9 9 1 9 1 13 4 9 1 3 13 1 1 10 0 9 13 2
16 10 9 1 12 0 9 1 9 13 4 1 9 14 15 13 2
23 11 11 1 13 16 0 9 0 0 9 9 1 3 0 9 1 0 13 1 9 1 13 2
22 0 9 0 7 0 9 1 9 1 0 7 0 9 1 0 9 1 9 1 1 13 2
16 15 9 10 9 1 9 7 9 1 9 1 1 0 13 13 2
32 11 1 11 11 11 11 11 11 1 9 2 9 1 0 9 1 3 13 1 1 15 0 13 4 1 9 1 13 1 9 13 2
11 3 2 11 1 9 13 1 9 14 13 2
36 11 11 1 11 11 11 11 13 1 3 13 4 9 1 9 13 4 11 1 13 16 9 15 9 13 4 4 16 15 9 0 9 1 0 13 2
27 3 2 11 11 1 15 0 11 11 11 1 9 14 14 13 7 15 9 1 9 13 1 15 9 14 13 2
27 15 10 9 1 12 0 0 9 1 9 9 1 9 13 1 9 1 12 9 1 13 4 4 1 9 13 2
21 11 11 1 13 16 15 0 9 9 1 10 9 0 2 0 13 1 9 14 13 2
9 7 11 10 9 1 0 14 13 2
28 9 1 13 1 9 2 9 1 9 1 9 1 9 9 1 0 9 1 9 1 1 0 9 13 1 9 13 2
32 9 9 1 11 1 13 16 9 0 12 2 12 9 1 9 1 11 7 0 2 0 11 1 0 9 1 1 13 1 0 13 2
39 11 11 11 2 11 2 1 9 11 11 11 1 13 16 0 12 9 1 9 0 13 4 4 2 7 15 9 1 9 1 15 0 13 1 9 13 4 4 2
45 15 13 16 10 9 9 0 9 1 0 9 1 3 13 4 4 7 16 15 15 10 9 13 4 16 0 12 2 12 9 1 11 7 0 2 0 11 1 0 9 1 9 13 4 2
28 15 1 14 11 1 13 16 11 2 11 7 11 1 0 12 2 12 9 1 0 0 9 7 9 1 9 13 2
38 11 1 11 9 1 9 11 11 11 1 13 16 11 2 11 2 11 2 0 11 11 7 11 1 10 9 1 13 9 1 0 9 1 9 13 4 4 2
32 11 1 13 16 11 11 11 1 0 2 0 9 1 10 9 1 9 13 4 4 7 15 11 2 11 11 1 13 1 9 13 2
17 10 9 1 10 9 9 1 9 1 9 13 4 10 9 1 13 2
23 11 1 13 16 11 1 0 9 7 0 2 0 11 1 0 9 2 9 2 13 4 4 2
32 15 0 12 9 1 11 11 2 11 7 11 1 0 9 2 11 2 13 4 4 2 15 9 1 0 13 1 9 13 4 4 2
22 0 0 9 15 13 16 11 1 0 9 1 1 13 0 9 11 1 1 13 4 4 2
45 15 13 16 0 2 0 11 1 10 9 11 11 11 1 0 9 1 13 9 1 10 9 1 9 1 9 13 4 2 7 0 12 9 1 10 9 1 10 9 1 9 14 13 4 2
32 16 2 10 9 11 11 11 1 0 2 0 9 1 10 9 1 9 13 4 4 7 15 0 2 0 9 1 13 1 9 13 2
26 15 9 1 0 7 0 11 1 11 2 11 2 11 7 11 1 0 12 9 1 9 13 1 9 13 2
22 15 1 11 1 9 1 9 13 16 15 10 9 1 10 9 1 0 13 1 0 13 2
20 11 1 9 1 11 1 12 2 12 9 9 13 2 15 14 9 1 10 13 2
11 9 1 11 1 15 1 9 14 13 4 2
13 10 9 1 10 9 1 9 1 13 1 9 13 2
19 11 1 11 9 1 11 11 11 1 9 1 9 1 0 9 10 0 13 2
16 15 13 13 16 11 1 9 1 0 0 9 1 9 13 4 2
26 11 9 1 0 9 9 11 11 1 13 13 16 11 1 0 9 1 9 9 1 9 13 4 4 4 2
28 16 2 15 15 9 13 4 16 11 1 9 1 9 9 11 11 1 15 9 1 0 13 1 15 9 14 13 2
21 11 1 16 10 9 15 9 1 0 13 16 2 0 9 11 1 1 0 13 4 2
31 11 11 1 0 9 11 11 11 1 13 13 16 11 1 9 1 1 13 1 0 13 16 9 1 0 9 1 9 0 13 2
9 3 2 11 1 15 9 13 4 2
24 11 1 16 10 9 0 13 15 9 13 4 4 2 16 15 9 1 3 9 1 9 0 13 2
23 15 12 9 14 13 16 11 1 9 1 9 7 10 9 1 0 0 9 1 9 13 4 2
20 11 11 1 9 11 11 1 13 13 16 11 1 9 9 1 9 1 14 13 2
19 9 1 9 1 1 0 13 16 11 9 1 1 1 15 9 1 9 13 2
11 16 2 11 1 1 11 1 9 3 13 2
24 3 2 15 9 13 4 4 16 0 9 1 0 0 9 11 1 9 1 9 13 1 9 13 2
14 16 2 11 1 9 1 13 4 15 9 3 10 13 2
22 0 11 9 1 11 11 11 1 9 1 11 7 11 1 9 1 13 1 9 14 13 2
15 15 9 1 14 9 13 7 12 9 1 1 9 3 13 2
17 11 1 11 1 0 9 11 11 11 7 11 11 1 10 9 13 2
27 11 11 11 1 13 13 16 11 11 1 3 11 11 1 13 1 12 9 1 1 0 9 1 9 0 13 2
19 15 13 2 15 9 13 16 11 7 11 1 1 0 9 1 10 9 13 2
16 10 9 1 11 7 11 9 1 1 9 9 1 3 9 13 2
12 11 1 1 14 15 0 0 9 13 4 4 2
29 15 1 1 11 11 11 1 13 16 11 1 13 13 16 11 1 1 0 9 1 15 9 1 15 9 14 13 4 2
28 11 11 1 13 16 11 1 3 11 13 1 12 9 1 9 1 9 1 9 14 13 7 15 9 1 9 13 2
18 15 13 16 11 11 11 1 11 7 11 1 9 1 10 9 14 13 2
26 11 2 11 11 7 11 1 11 11 11 1 9 1 11 7 11 9 1 14 9 0 13 4 13 4 2
24 11 11 1 13 12 9 1 9 1 9 1 13 7 9 1 9 1 13 1 9 13 4 4 2
10 9 1 15 11 1 9 13 4 4 2
6 15 0 9 1 13 2
18 9 1 13 4 4 16 16 11 11 11 13 16 15 14 13 4 4 2
10 10 9 13 9 1 9 9 14 13 2
16 11 1 9 1 13 13 16 11 11 1 15 15 9 14 13 2
8 11 11 1 9 0 13 4 2
11 11 11 1 15 11 1 9 1 0 13 2
9 9 1 1 11 1 9 13 4 2
22 16 15 9 1 9 14 13 16 15 1 0 9 1 9 1 0 11 11 1 9 13 2
12 11 1 11 11 13 16 9 1 13 4 4 2
16 16 15 9 14 13 16 11 9 9 1 1 11 1 9 13 2
6 15 9 11 11 13 2
15 15 9 1 10 9 15 9 1 9 1 1 13 4 4 2
10 10 9 13 9 1 9 9 13 4 2
12 9 1 15 0 9 1 9 1 9 13 4 2
19 11 1 9 9 11 11 1 13 16 11 11 3 0 9 1 9 13 4 2
16 11 11 1 9 11 11 1 13 16 11 11 9 1 13 4 2
14 9 1 9 9 1 3 10 9 1 1 9 13 4 2
28 11 11 11 1 9 9 1 9 9 11 11 11 1 13 13 16 9 1 9 1 9 9 14 13 4 4 4 2
17 15 13 16 15 14 9 1 11 11 9 1 15 9 14 13 4 2
12 11 11 9 1 3 10 9 1 9 13 4 2
7 15 9 1 9 0 13 2
12 11 11 11 11 1 9 1 1 9 13 4 2
25 11 1 11 11 9 9 1 9 9 11 11 1 13 13 16 11 11 10 0 7 9 1 9 13 2
8 15 3 15 9 1 13 4 2
16 9 9 11 11 1 13 16 11 11 15 1 3 13 13 4 2
14 10 9 13 9 13 1 9 13 14 0 9 13 4 2
11 9 11 9 1 0 9 1 9 1 13 2
20 9 7 9 9 1 14 11 11 9 13 0 9 1 9 13 7 9 9 13 2
9 9 1 1 15 9 8 14 13 2
13 15 1 9 9 1 0 9 9 1 0 13 4 2
13 15 9 1 3 1 9 13 1 9 14 13 4 2
22 10 9 1 9 9 1 9 1 13 11 11 11 11 11 1 9 1 9 1 1 13 2
14 15 13 16 9 1 9 9 3 9 1 13 9 13 2
14 11 1 0 9 9 1 1 11 1 9 1 9 13 2
17 15 15 1 10 12 9 1 9 13 15 9 1 1 9 0 13 2
25 15 13 16 11 9 1 3 10 9 13 15 9 9 7 9 9 1 0 9 1 9 13 4 4 2
15 0 9 9 1 1 11 1 12 12 9 1 9 9 13 2
27 11 1 13 16 11 1 9 1 13 1 9 7 9 1 1 10 9 12 12 9 1 9 8 13 4 4 2
7 15 9 13 4 4 4 2
21 15 13 16 9 1 0 9 13 1 0 9 11 2 11 9 1 13 4 4 4 2
31 15 13 16 10 9 1 9 1 9 1 3 1 9 9 13 2 15 9 9 1 9 1 13 1 3 14 8 14 13 4 2
13 10 9 1 10 9 1 10 9 1 13 4 4 2
24 3 2 11 9 1 9 1 13 4 15 14 11 11 11 9 13 1 11 11 9 13 4 4 2
29 15 9 1 0 9 1 1 1 13 16 11 1 9 1 11 1 11 7 11 1 11 9 1 9 13 0 9 13 2
20 11 1 13 16 9 1 9 9 1 14 0 9 13 1 9 13 4 4 4 2
10 15 9 1 11 11 11 9 13 4 2
20 0 9 1 15 9 1 9 13 4 11 1 11 15 12 9 1 13 4 4 2
21 11 1 9 1 11 1 9 9 1 13 11 1 9 1 15 1 9 13 4 4 2
20 9 1 11 14 14 16 15 9 1 14 9 1 9 1 13 1 9 13 4 2
34 9 1 13 13 16 11 1 11 1 9 1 1 11 11 1 12 12 9 13 1 3 2 9 9 1 9 1 10 13 1 9 13 4 2
16 15 15 15 0 9 1 1 2 9 0 9 1 13 4 4 2
14 11 1 13 9 1 1 9 1 9 0 9 1 13 2
41 15 10 9 1 13 9 1 13 4 9 1 9 1 15 9 1 1 13 4 10 9 1 9 13 1 1 9 14 13 4 15 9 1 9 13 1 9 14 13 4 2
16 7 9 1 11 1 13 16 15 10 15 14 9 14 13 4 2
13 11 1 9 1 0 9 13 1 9 1 0 13 2
29 15 10 9 1 0 9 7 15 1 9 1 13 13 16 11 15 9 1 13 4 4 7 15 1 15 9 9 13 2
27 15 9 1 9 1 13 4 4 16 9 1 11 7 15 12 9 11 11 7 11 11 1 9 14 13 4 2
17 16 15 9 15 1 1 15 9 1 9 13 16 9 2 9 13 2
18 9 1 15 14 13 13 16 11 0 9 1 9 1 1 9 14 13 2
43 10 9 9 1 11 15 9 1 9 1 13 4 4 7 12 0 11 9 1 9 1 9 13 4 13 16 9 1 9 0 13 7 10 9 1 11 11 11 1 9 13 4 2
32 9 1 13 13 16 11 1 11 1 14 9 13 7 16 11 13 16 11 11 1 9 1 9 1 1 14 10 9 13 4 4 2
12 9 1 15 1 0 9 1 14 9 0 13 2
11 15 3 2 3 0 9 13 4 4 4 2
16 9 1 12 0 9 11 1 9 14 9 1 9 1 13 4 2
20 11 1 11 9 12 9 9 1 1 9 1 13 4 9 1 0 9 13 4 2
10 12 9 1 1 3 9 7 9 13 2
16 9 1 9 13 1 9 1 9 9 1 9 13 7 9 13 2
11 9 1 15 1 12 9 1 0 13 4 2
20 0 9 1 9 1 1 11 7 11 9 1 0 9 1 0 13 4 4 4 2
25 0 9 1 12 9 9 13 1 3 14 12 9 1 14 10 9 13 4 7 9 9 0 13 4 2
15 9 1 9 13 1 1 9 1 9 7 0 9 13 4 2
22 9 9 0 11 11 11 11 1 9 13 16 11 1 9 0 9 0 7 9 1 13 2
12 0 9 7 0 9 9 1 9 13 4 4 2
30 11 1 13 16 9 9 1 9 13 1 0 11 11 1 1 11 11 11 11 1 3 12 12 9 1 9 0 13 4 2
28 0 9 1 13 16 11 1 12 9 1 9 13 1 3 13 9 7 9 1 9 1 14 9 13 4 4 4 2
39 11 1 11 2 11 1 11 11 1 9 1 9 1 13 11 9 9 7 9 1 9 13 9 1 9 1 11 1 0 9 9 1 9 2 9 0 13 4 2
23 9 1 9 1 1 11 1 9 9 1 9 1 9 1 13 11 11 1 9 1 9 13 2
30 15 1 0 9 1 0 9 1 9 1 9 13 11 1 0 9 1 9 1 9 13 4 2 15 12 9 0 13 4 2
9 9 1 9 9 13 7 9 13 2
20 0 9 7 9 1 9 1 1 10 9 2 9 9 1 1 0 13 4 4 2
16 9 11 1 11 1 14 10 9 9 0 13 1 9 13 4 2
12 9 11 11 1 14 13 16 9 1 9 13 2
25 0 13 16 11 2 11 1 11 9 11 11 1 9 11 1 9 11 11 1 11 11 1 1 13 2
18 9 1 1 9 7 9 1 9 1 9 13 1 13 9 13 4 4 2
20 9 1 1 0 9 1 9 1 9 13 4 4 7 3 9 7 9 13 4 2
44 9 13 9 1 1 9 9 9 0 13 1 15 9 1 15 1 9 1 9 9 13 4 7 9 14 12 9 9 1 9 1 9 1 9 9 1 9 1 9 1 1 13 4 2
7 12 9 11 9 1 13 2
13 9 1 9 0 9 13 7 9 1 9 13 4 2
29 11 11 1 12 0 9 11 7 11 11 1 12 9 1 9 11 11 9 14 12 12 9 9 1 1 13 4 4 2
11 9 13 1 3 14 10 9 9 14 13 2
24 11 1 15 15 9 13 4 15 9 1 14 12 9 1 9 1 1 13 9 1 15 9 13 2
12 12 9 9 1 9 13 4 7 9 14 13 2
24 15 1 0 9 0 13 4 7 12 9 1 9 1 1 11 11 11 1 1 9 1 13 4 2
19 9 11 11 11 11 1 15 9 1 0 13 1 9 13 15 9 13 4 2
15 9 0 13 4 7 9 1 0 9 1 9 9 13 4 2
11 11 1 13 1 9 13 16 15 13 4 2
13 11 11 11 1 9 1 9 13 9 13 4 4 2
18 15 9 1 9 1 10 9 1 9 1 13 0 9 1 9 13 4 2
16 9 1 9 13 1 1 9 1 9 1 9 1 0 9 13 2
22 11 11 1 11 13 4 11 11 1 0 9 7 9 1 12 9 1 0 9 13 4 2
38 11 11 1 9 7 11 11 11 11 2 11 2 1 13 9 2 9 1 1 9 1 13 13 9 1 12 9 1 9 13 4 7 12 15 0 13 4 2
18 10 9 11 1 9 12 9 11 1 11 9 1 11 9 9 1 13 2
19 11 9 1 9 1 9 1 9 7 9 1 9 13 15 1 9 13 4 2
25 15 1 13 9 1 11 9 1 11 11 11 1 9 1 9 1 11 1 12 9 1 9 13 4 2
19 11 9 1 0 9 11 11 7 11 11 1 11 11 11 8 13 4 4 2
8 3 9 1 15 9 13 4 2
22 3 11 1 9 1 13 16 10 9 1 9 1 13 1 9 1 9 13 1 9 13 2
16 10 9 1 11 9 1 9 9 14 0 9 1 0 13 4 2
24 11 1 9 9 11 11 11 1 13 16 11 2 11 11 11 1 11 9 1 10 9 9 13 2
14 10 9 9 2 9 9 9 1 9 13 4 4 4 2
18 7 13 9 1 14 9 1 10 9 1 0 9 1 9 7 9 13 2
10 10 9 9 1 1 11 13 4 4 2
17 10 9 1 1 9 1 9 9 1 11 1 15 9 1 9 13 2
14 15 1 14 11 1 9 1 12 9 9 1 13 4 2
6 7 9 15 14 13 2
32 15 1 15 1 12 9 1 11 1 9 1 9 9 1 9 0 13 9 1 3 13 4 7 9 1 3 13 1 9 13 4 2
13 7 9 1 9 1 9 7 9 1 0 13 4 2
20 15 10 9 1 14 12 9 9 1 9 13 9 1 0 9 1 9 13 4 2
18 15 12 1 9 9 1 13 4 7 12 9 1 9 1 9 13 4 2
19 9 9 1 13 16 15 1 9 1 9 1 12 9 1 9 1 13 4 2
18 15 1 12 1 9 13 4 4 7 12 1 0 9 1 0 13 4 2
31 9 1 13 16 0 9 1 1 0 9 1 11 9 1 10 9 1 9 12 9 9 1 15 9 1 1 0 13 4 4 2
20 7 11 1 9 11 7 11 9 1 9 13 9 1 13 1 9 13 4 4 2
36 3 11 1 9 9 9 9 11 11 11 1 13 16 11 11 2 11 2 1 9 1 1 12 9 1 11 11 1 1 9 1 1 13 4 4 2
31 11 1 3 14 9 11 1 11 9 1 12 9 1 13 3 12 2 12 9 7 12 2 12 9 9 1 9 1 13 4 2
9 9 12 9 1 1 9 13 4 2
8 11 9 1 9 1 15 13 2
27 0 9 1 9 1 13 1 3 14 12 9 13 4 7 11 9 1 9 1 9 7 9 13 9 13 4 2
12 9 1 11 9 1 9 1 14 9 13 4 2
17 11 11 11 11 1 12 0 9 1 11 1 11 1 1 0 13 2
30 11 10 9 11 2 11 11 11 1 9 13 11 13 4 4 15 9 1 11 11 1 13 9 1 9 0 13 4 4 2
28 11 11 1 11 11 7 11 1 11 11 11 9 1 1 0 9 2 0 9 7 0 9 1 9 1 9 13 2
14 11 11 1 11 9 1 1 12 0 9 1 9 13 2
14 15 1 12 9 9 9 1 0 9 9 1 13 4 2
17 0 9 0 9 1 9 1 0 12 9 9 1 9 1 13 4 2
10 12 9 1 9 9 1 10 9 13 2
35 10 9 1 0 9 13 4 16 11 9 1 9 1 9 1 9 14 13 7 10 9 0 13 16 11 0 9 1 0 9 0 13 13 4 2
31 9 9 11 11 1 11 1 13 16 10 9 0 9 1 0 9 7 0 9 1 0 9 1 9 1 9 9 13 4 4 2
19 16 10 9 15 10 9 1 14 13 16 15 9 1 9 1 9 13 4 2
14 0 9 9 1 13 13 1 9 11 1 9 1 13 2
18 15 12 9 1 11 1 9 9 9 0 9 1 0 13 1 9 13 2
13 15 1 11 11 1 11 1 11 1 9 13 4 2
26 15 15 11 11 11 1 11 1 9 1 11 11 1 9 1 11 1 0 9 1 9 13 4 4 4 2
23 11 12 9 1 11 1 1 13 2 7 9 1 15 9 1 1 9 1 0 9 13 4 2
22 0 9 11 11 11 9 1 11 11 7 11 9 11 11 1 9 1 9 13 4 4 2
23 9 1 13 16 11 0 9 9 11 7 11 1 0 9 1 10 9 0 13 1 9 13 2
13 11 15 9 1 1 10 9 1 14 13 4 4 2
40 11 1 11 11 9 13 1 9 1 9 14 13 1 1 11 1 11 11 7 11 1 13 4 4 9 1 1 11 11 11 11 1 11 1 11 9 9 13 4 2
26 11 7 11 12 12 9 1 9 1 12 9 0 9 9 1 1 11 1 11 11 9 13 1 0 13 2
13 9 1 9 1 12 9 1 1 0 9 9 13 2
12 11 11 11 1 9 7 9 9 1 9 13 2
17 15 11 1 11 11 11 11 11 7 11 11 11 11 1 9 13 2
24 7 11 1 13 13 16 11 11 11 1 9 1 11 9 1 9 1 9 1 9 13 4 4 2
30 9 1 13 16 11 1 9 13 4 16 15 11 1 9 1 15 13 9 1 13 1 1 11 11 11 13 1 0 13 2
18 9 1 1 15 1 11 13 4 16 11 11 1 1 0 9 14 13 2
13 0 9 1 11 1 0 9 1 9 1 13 4 2
35 11 11 1 14 9 13 4 4 16 15 11 2 11 2 11 1 1 11 2 11 2 11 2 11 2 9 9 1 15 9 9 1 0 13 2
15 11 11 11 11 11 2 11 9 9 1 14 12 9 13 2
17 15 11 10 9 10 0 9 1 9 1 13 9 0 13 4 4 2
15 0 3 11 11 1 10 9 1 9 1 9 13 4 4 2
14 11 11 1 11 2 11 7 11 1 1 0 13 4 2
20 15 10 9 1 9 11 2 11 7 11 1 9 9 1 9 1 9 13 4 2
32 9 1 10 9 1 13 1 0 9 1 1 0 9 1 9 2 9 10 13 1 0 9 1 3 0 9 11 11 11 0 13 2
10 15 11 11 1 0 9 9 0 13 2
22 11 11 1 9 1 1 0 9 1 1 10 9 1 9 1 1 9 1 3 9 13 2
24 11 9 9 1 0 9 13 1 1 9 1 14 13 4 1 12 9 1 0 9 1 9 13 2
32 11 9 7 9 9 1 9 1 9 1 13 1 1 11 9 12 13 12 9 1 10 9 7 9 9 1 9 1 9 13 4 2
20 9 9 1 13 16 10 9 1 9 12 9 1 1 14 9 9 0 13 4 2
17 11 9 9 1 12 12 9 1 9 9 13 9 9 0 13 4 2
20 3 11 1 10 9 1 13 0 9 1 1 1 9 0 2 0 13 4 4 2
17 10 3 11 11 9 1 0 9 1 9 9 11 1 9 13 4 2
14 11 13 11 1 1 13 1 12 9 1 0 13 4 2
21 0 9 9 1 11 7 11 13 11 1 1 13 1 12 9 1 14 0 13 4 2
29 11 1 11 11 9 1 11 9 9 1 12 9 1 9 1 12 9 1 10 9 1 13 13 15 9 9 0 13 2
11 9 1 10 9 1 0 2 0 13 4 2
27 11 11 1 13 16 15 0 9 9 1 9 1 9 1 0 11 11 11 1 9 1 0 13 1 0 13 2
24 15 1 14 11 7 11 11 1 1 1 15 0 13 1 10 15 9 1 9 13 1 0 13 2
50 11 1 11 11 11 1 11 1 15 9 1 13 16 15 9 9 1 1 11 9 1 1 1 9 1 13 9 1 9 13 1 1 11 1 11 11 11 1 0 13 1 1 9 1 0 13 1 0 13 2
37 11 11 11 2 11 2 1 9 1 9 1 1 9 0 13 1 9 9 1 9 1 9 13 4 9 9 1 9 1 0 9 13 1 9 13 4 2
45 3 9 9 1 11 1 12 9 9 1 15 13 4 0 9 13 1 9 13 4 4 16 10 9 1 0 9 1 9 1 9 0 14 13 7 9 1 1 14 9 1 0 13 4 2
44 10 9 1 11 11 11 11 1 9 1 0 13 4 9 11 11 11 7 9 11 11 11 1 9 1 9 9 1 11 11 2 11 11 7 11 11 11 1 9 13 1 9 13 2
17 10 9 1 12 9 1 10 9 1 9 13 9 0 13 4 4 2
23 9 1 15 9 1 10 9 1 12 9 1 1 0 9 1 12 9 13 1 9 13 4 2
28 9 9 9 1 10 9 1 0 14 13 16 9 1 1 9 0 13 1 1 12 9 0 9 1 0 14 13 2
42 9 1 13 16 15 10 9 1 9 13 16 9 1 9 13 1 3 9 9 10 9 9 1 10 9 1 9 13 16 10 9 1 9 13 1 15 10 9 0 13 4 2
19 9 1 13 16 9 9 1 9 1 0 10 9 1 9 0 13 4 4 2
17 15 1 11 11 11 1 14 12 9 1 9 13 1 9 13 4 2
33 10 9 1 0 9 9 1 13 16 16 9 9 9 1 15 1 9 13 16 15 11 11 11 1 9 1 9 1 15 9 14 13 2
18 9 9 9 11 11 11 1 13 16 11 1 9 9 1 13 13 4 2
16 9 11 1 13 16 15 10 9 9 1 9 1 9 13 4 2
22 15 13 16 15 11 9 1 11 11 7 0 9 1 1 9 10 0 9 1 13 4 2
17 9 11 1 13 16 9 13 1 1 12 0 9 9 13 4 4 2
20 10 9 9 1 9 9 9 13 1 3 13 4 1 9 1 14 9 13 4 2
11 9 11 1 13 16 9 1 9 0 13 2
27 15 1 1 9 13 4 15 13 16 11 1 11 1 0 9 1 9 1 9 1 12 9 1 0 13 4 2
19 9 11 1 13 16 0 9 10 9 1 1 9 1 12 14 9 13 4 2
18 10 9 1 11 1 9 13 1 1 1 9 11 1 15 9 14 13 2
15 15 13 16 9 9 1 12 9 0 9 1 9 13 4 2
12 10 9 1 3 9 13 1 13 4 4 4 2
26 9 11 1 13 16 9 9 1 11 9 1 11 1 12 9 9 1 9 13 1 9 0 13 4 4 2
39 9 1 9 9 1 13 4 1 1 11 11 1 9 0 13 4 1 1 1 9 11 1 13 16 0 11 11 1 10 9 1 1 1 9 13 4 4 4 2
32 11 11 1 9 9 11 11 1 12 9 1 10 10 9 1 0 9 0 13 4 4 2 15 11 11 11 11 1 0 9 13 2
14 9 1 1 10 9 1 1 9 10 9 11 1 13 2
25 9 13 16 15 9 1 1 11 11 11 1 1 14 9 7 0 11 1 9 1 9 1 9 13 2
9 10 9 11 1 0 9 1 13 2
35 11 1 9 1 10 9 11 11 11 11 11 1 11 2 11 7 0 0 9 1 0 9 1 1 10 9 1 9 1 1 0 13 4 4 2
16 9 1 9 9 1 9 2 9 1 9 1 9 14 13 4 2
22 11 11 0 9 1 11 1 12 1 10 9 7 9 1 13 1 1 9 13 4 4 2
35 15 11 11 2 11 2 11 2 11 9 9 11 11 7 11 11 11 1 0 9 1 9 1 9 1 1 1 13 4 12 0 9 0 13 2
24 0 9 1 1 11 1 0 9 0 11 1 9 1 13 1 1 11 1 9 9 13 4 4 2
29 15 13 4 4 4 16 0 9 1 11 1 9 1 12 9 9 11 11 11 7 11 11 11 1 9 14 0 13 2
15 15 1 0 9 9 11 1 0 9 2 9 13 4 4 2
32 9 9 1 1 12 9 1 9 1 9 13 7 15 11 11 1 11 11 11 1 9 1 1 9 7 9 13 1 9 13 4 2
69 2 11 11 11 2 1 0 9 1 1 9 1 0 9 1 0 11 1 0 9 1 11 11 11 2 9 11 2 11 11 2 11 11 11 2 11 11 11 11 2 11 11 11 11 2 11 11 11 2 11 11 11 11 2 11 11 11 11 2 11 11 7 11 11 11 11 0 13 2
40 11 11 11 1 11 9 1 9 11 11 11 1 11 1 9 13 16 11 11 1 11 1 9 9 1 12 9 1 11 1 0 9 1 9 1 9 13 4 4 2
61 11 11 11 2 11 2 1 9 11 11 11 1 15 9 1 13 16 11 1 11 9 1 9 7 11 11 1 15 11 0 11 11 1 11 11 1 9 7 15 1 14 11 11 11 1 13 9 1 9 9 1 1 9 9 13 1 9 13 4 4 2
23 11 1 13 16 15 1 11 1 12 9 1 12 9 1 9 9 1 9 13 4 4 4 2
18 10 9 9 1 1 15 15 1 9 1 9 13 1 9 13 4 4 2
17 15 13 16 11 11 1 10 9 1 12 9 1 9 1 9 13 2
27 11 1 11 9 1 1 9 1 9 13 1 1 0 9 11 1 9 1 13 12 0 9 1 9 13 4 2
46 15 13 16 15 11 11 1 9 9 9 11 11 11 2 0 9 11 2 11 2 11 7 11 11 11 1 9 11 11 1 9 13 7 15 1 9 1 9 1 13 9 1 0 9 13 2
24 11 1 13 16 15 9 1 9 1 9 13 4 4 7 15 1 1 15 0 9 14 13 4 2
26 15 13 16 9 1 9 1 9 11 1 9 11 11 1 9 2 9 1 13 15 11 1 9 0 13 2
19 15 13 16 15 15 0 13 4 4 16 9 1 15 9 2 9 14 13 2
16 15 13 16 9 1 11 1 9 7 9 2 9 0 13 4 2
27 9 13 4 16 11 1 0 11 1 0 9 11 11 1 11 11 1 2 0 9 2 1 9 13 4 4 2
23 11 1 9 1 0 9 1 0 13 4 16 9 1 10 9 1 9 9 9 13 4 4 2
15 9 1 13 4 16 3 0 9 1 10 9 9 13 4 2
25 15 1 9 1 11 11 11 11 7 11 11 1 11 11 1 10 9 1 9 0 13 1 13 4 2
27 11 11 14 11 11 1 9 13 1 11 11 1 9 1 1 0 9 1 9 9 9 1 9 13 4 4 2
19 11 11 1 9 1 9 1 9 13 4 11 11 1 11 11 13 4 4 2
21 11 9 11 11 1 9 1 9 1 0 11 11 1 11 11 1 1 13 13 4 2
9 10 9 1 9 9 1 9 13 2
31 11 1 13 13 16 11 1 1 0 12 9 15 12 9 1 13 4 4 4 7 9 9 1 9 1 9 13 4 4 4 2
44 9 11 11 11 7 9 11 11 11 1 9 1 11 11 1 11 11 1 9 7 11 11 1 13 4 9 1 15 1 0 9 9 1 13 4 9 13 1 0 9 0 13 4 2
29 11 11 1 9 1 13 16 11 1 11 11 1 0 12 9 9 1 1 12 11 11 1 9 1 9 1 0 13 2
26 10 9 15 9 1 9 1 9 1 9 1 0 13 7 9 1 9 1 1 9 1 1 9 13 4 2
22 11 1 9 11 11 11 1 13 16 15 9 1 14 15 9 1 0 13 4 4 4 2
16 9 15 11 1 1 13 1 9 13 1 3 9 1 9 13 2
13 9 1 15 1 14 9 11 11 1 0 13 4 2
24 11 1 13 16 11 11 1 9 1 1 14 11 1 1 9 9 1 9 1 15 9 14 13 2
20 15 1 9 1 13 16 10 9 1 1 11 1 9 1 14 9 9 1 13 2
27 9 1 13 9 9 1 13 4 1 3 11 1 12 9 9 1 0 11 1 9 9 1 9 9 13 4 2
14 9 9 1 13 16 9 1 0 10 12 9 0 13 2
16 11 1 11 13 4 10 9 1 11 11 11 11 1 13 4 2
8 9 1 9 13 4 4 4 2
24 10 9 11 11 11 1 11 11 11 1 13 1 7 13 4 1 14 12 9 1 14 13 4 2
22 11 9 1 0 9 1 10 12 9 7 9 9 1 12 9 9 2 9 13 4 4 2
23 9 1 11 11 1 13 16 9 0 13 1 1 1 9 13 4 9 1 9 13 4 4 2
25 11 1 15 1 1 13 4 4 16 9 1 9 13 1 12 9 1 1 14 9 1 13 4 4 2
17 15 13 16 1 9 9 9 1 14 1 10 9 1 13 4 4 2
11 15 13 16 10 3 15 14 0 14 13 2
8 9 1 9 13 4 4 4 2
32 11 1 11 11 1 9 1 9 1 1 13 9 1 14 12 10 9 1 9 1 13 1 3 11 11 1 9 9 13 4 4 2
13 10 9 11 11 11 1 9 1 9 1 0 13 2
27 10 9 1 9 14 0 13 2 15 9 13 4 16 11 11 1 14 0 9 7 9 1 1 9 13 4 2
18 16 10 12 9 1 11 11 11 1 13 4 9 1 10 9 14 13 2
14 10 9 1 0 9 1 0 9 1 13 13 4 4 2
14 10 10 9 14 13 2 15 0 9 9 1 0 13 2
12 15 11 1 9 1 0 9 13 4 4 4 2
13 10 12 9 11 1 9 1 12 9 1 13 4 2
26 10 9 1 9 1 13 1 9 1 13 13 16 10 9 1 15 9 11 1 9 1 13 1 13 4 2
14 15 0 14 13 4 16 10 9 1 13 1 15 13 2
21 11 11 1 13 13 16 11 1 9 13 1 3 9 1 9 9 13 4 4 4 2
31 11 1 0 9 1 9 13 4 16 11 11 1 0 9 1 9 1 9 13 1 3 9 13 4 9 1 10 9 13 4 2
21 12 9 1 15 9 1 0 13 13 4 4 7 15 9 1 0 9 1 9 13 2
33 11 11 1 9 11 11 1 15 0 9 1 13 4 16 10 9 1 0 9 7 9 1 1 13 9 1 13 10 9 0 13 4 2
21 10 9 11 11 11 11 1 13 4 4 4 7 9 1 9 0 13 4 4 4 2
31 9 1 13 9 7 9 1 9 1 1 15 11 11 11 11 1 0 9 7 9 1 13 9 1 9 14 9 13 4 4 2
23 9 7 9 9 9 1 12 9 11 11 1 10 0 0 9 1 0 9 9 13 4 4 2
27 10 9 10 9 1 9 13 16 11 11 1 13 0 9 1 10 0 9 1 9 1 10 9 1 9 13 2
18 15 9 10 9 1 13 16 15 10 9 9 1 9 14 14 13 4 2
17 10 9 11 11 1 0 9 0 9 1 9 1 1 1 9 13 2
34 11 11 11 11 9 11 11 1 11 1 9 1 13 16 15 1 9 1 13 9 1 9 1 9 1 9 1 9 1 14 9 13 4 2
20 7 2 15 15 9 14 13 16 15 9 13 4 7 15 15 9 1 9 13 2
24 11 1 13 2 9 1 13 9 13 4 4 16 0 9 1 9 1 9 1 10 9 9 13 2
24 11 1 13 16 9 9 1 12 9 9 1 9 1 9 7 9 1 13 9 1 9 13 4 2
12 11 1 9 1 12 0 9 15 13 4 4 2
26 10 9 9 1 11 11 11 1 9 9 1 9 13 7 11 11 11 11 2 11 2 1 3 9 13 2
31 11 1 13 16 15 9 9 1 9 13 3 11 1 9 9 1 9 13 9 2 9 1 9 1 9 7 9 1 9 13 2
25 15 13 16 15 0 9 13 16 0 9 1 1 11 1 0 9 1 0 9 0 9 0 13 4 2
11 15 1 9 1 9 1 14 9 13 4 2
15 7 2 15 15 14 0 9 0 9 1 9 1 13 13 2
30 15 13 4 16 0 9 1 9 1 9 1 0 9 1 0 9 13 4 7 10 9 1 15 3 9 0 13 0 13 2
19 11 11 11 11 11 9 11 11 14 9 11 11 1 9 1 9 13 4 2
26 15 13 16 16 0 9 9 1 9 1 9 1 13 4 4 16 3 15 9 1 0 9 13 4 4 2
21 15 13 16 15 9 1 13 9 13 1 9 7 9 1 9 9 1 13 4 4 2
13 0 9 1 0 9 9 2 9 13 1 9 13 2
23 11 9 11 11 13 4 16 9 1 9 1 1 9 1 9 1 9 1 0 13 4 4 2
15 16 9 1 9 1 13 1 9 1 0 9 13 4 4 2
45 11 11 11 11 11 11 7 11 11 11 11 11 11 1 9 1 13 7 9 9 11 11 2 11 11 11 7 11 1 11 11 1 9 1 9 13 3 2 3 0 13 4 4 4 2
12 11 13 4 16 9 1 10 9 1 9 13 2
18 10 9 11 11 2 11 2 11 2 11 7 11 1 15 9 14 13 2
21 9 13 4 4 4 11 11 1 11 11 1 11 11 11 1 9 13 4 4 4 2
20 9 1 0 9 1 9 13 1 1 11 11 1 14 9 1 9 13 4 4 2
13 11 11 7 11 9 1 12 13 4 1 9 13 2
17 11 9 1 1 10 12 9 9 9 1 12 14 9 1 1 13 2
24 11 11 1 9 2 9 1 9 1 9 1 13 4 11 11 1 9 1 9 13 4 4 4 2
15 11 11 11 1 9 1 9 1 11 1 0 9 13 4 2
26 11 11 11 11 11 1 9 11 11 1 9 1 1 0 13 9 1 11 1 14 13 4 1 9 13 2
14 11 11 11 11 11 1 9 1 14 9 0 14 13 2
16 0 9 15 2 0 11 2 1 1 9 1 14 13 4 4 2
19 7 9 1 0 9 1 3 13 4 11 11 1 13 1 1 0 14 13 2
23 11 9 1 9 13 16 10 9 9 1 13 11 11 1 13 1 9 1 0 9 14 13 2
16 0 9 1 0 9 1 1 1 9 2 9 13 1 9 13 2
32 15 1 9 15 13 4 4 4 16 9 1 0 9 13 1 9 1 9 1 9 9 1 1 9 1 13 1 1 9 13 4 2
19 16 2 9 1 1 9 1 9 1 9 1 0 9 1 9 13 4 4 2
19 3 2 9 1 9 1 13 1 9 1 9 9 1 0 9 13 4 4 2
19 11 11 11 11 2 11 2 1 9 1 9 11 11 1 13 1 9 13 2
28 15 13 4 4 4 16 11 11 1 11 1 9 7 9 9 1 11 1 13 4 9 1 15 9 13 4 4 2
18 15 1 9 9 13 15 14 9 1 9 0 9 1 9 13 4 4 2
12 10 9 12 9 1 1 12 9 1 0 13 2
32 0 13 16 11 11 1 9 1 11 11 11 2 11 2 1 9 1 11 11 1 9 13 15 0 9 1 9 1 9 13 4 2
21 15 1 11 11 1 10 9 15 2 15 9 1 9 13 1 1 9 13 4 4 2
12 11 11 1 9 11 11 1 9 13 4 4 2
24 12 12 12 9 1 11 11 1 11 9 1 1 9 1 9 11 1 10 14 0 13 4 4 2
28 0 9 1 11 11 1 12 9 9 7 11 1 9 11 11 1 9 13 4 10 9 1 9 9 13 4 4 2
25 11 1 11 1 11 9 1 9 13 1 9 13 7 15 0 9 9 1 9 13 1 9 13 4 2
15 11 0 9 1 9 9 1 9 11 1 11 11 1 13 2
29 10 9 1 11 11 2 11 2 11 7 11 1 10 9 2 15 11 1 9 13 2 1 11 11 9 1 9 13 2
21 15 13 16 10 9 1 9 1 11 0 9 1 0 9 9 0 13 1 9 13 2
31 9 9 1 1 2 10 9 1 0 11 11 11 11 11 11 1 9 1 10 0 9 0 9 1 9 9 1 14 9 13 2
33 11 1 11 11 11 11 1 11 9 1 1 12 9 1 1 9 9 7 9 1 0 9 1 0 9 1 9 13 1 9 13 4 2
27 11 11 1 11 13 1 9 10 9 1 1 13 4 2 7 11 1 11 9 14 10 9 13 1 9 13 2
33 11 1 11 11 11 11 7 11 11 11 11 11 1 1 11 9 12 9 13 9 1 1 12 9 1 1 0 9 1 0 9 13 2
37 11 7 11 11 1 11 1 9 1 1 15 14 0 13 16 9 2 9 2 9 2 9 7 9 9 9 9 9 1 9 1 3 0 9 13 4 2
17 12 9 15 11 2 11 11 11 1 9 1 9 1 0 9 13 2
34 11 11 1 9 11 11 1 1 9 9 1 1 3 0 11 2 11 7 11 2 11 9 9 1 9 1 14 12 9 1 1 9 13 2
17 0 13 16 2 11 11 11 11 2 10 9 1 9 1 9 13 2
25 10 9 1 1 11 2 11 7 11 2 11 1 1 1 9 1 9 9 1 9 9 9 13 4 2
25 11 11 1 11 1 11 11 11 11 2 11 11 11 7 11 11 11 11 11 11 1 14 9 13 2
27 15 0 0 9 1 9 9 1 1 12 9 1 1 13 9 1 9 9 9 9 1 14 9 1 9 13 2
15 15 16 12 9 13 4 9 13 16 10 3 13 4 4 2
37 11 1 9 9 1 11 11 11 11 1 13 1 11 11 11 11 2 11 2 1 9 1 9 1 9 13 1 9 1 11 1 9 1 9 13 4 2
22 0 9 1 14 15 9 0 13 4 11 1 10 9 1 9 13 1 1 9 13 4 2
38 11 1 9 11 11 1 13 13 16 11 9 1 0 9 1 13 10 9 13 4 16 9 1 10 9 7 10 9 1 11 1 1 9 1 9 13 4 2
16 11 11 2 11 2 1 14 9 1 9 1 0 9 13 4 2
28 9 1 9 11 11 11 1 13 16 9 1 9 1 9 1 9 13 4 11 1 9 1 9 14 13 4 4 2
38 0 9 1 14 9 14 1 11 11 11 1 13 13 4 16 9 1 10 9 1 9 1 13 1 1 0 0 9 1 9 9 13 9 1 9 13 4 2
11 7 9 1 9 1 9 1 9 13 4 2
31 9 1 13 13 16 11 15 0 9 9 13 7 0 0 7 9 1 9 1 15 9 1 0 9 1 15 9 1 9 13 2
5 15 10 9 13 2
13 15 13 16 11 11 11 1 9 1 0 14 13 2
12 16 15 15 1 1 9 1 15 14 14 13 2
19 11 1 0 9 13 4 11 1 0 11 11 11 11 11 1 11 11 13 2
17 9 1 1 11 11 11 7 0 9 1 1 15 9 1 9 13 2
14 9 1 1 11 0 9 2 9 1 1 15 13 4 2
21 9 1 1 11 1 9 1 9 1 1 9 11 1 9 13 1 1 11 1 13 2
32 11 11 1 11 11 11 1 13 9 1 9 11 2 11 2 11 1 9 11 11 1 13 9 1 9 11 11 1 0 13 4 2
23 16 2 9 1 0 9 11 11 11 1 13 9 1 12 9 1 0 9 1 0 13 4 2
31 3 1 11 11 1 11 11 7 11 11 1 9 1 9 13 4 0 9 1 9 1 11 7 11 11 1 0 13 4 4 2
34 11 7 11 1 9 1 9 1 1 11 11 1 9 13 4 7 11 9 1 9 1 11 7 11 1 0 13 1 9 1 9 13 4 2
24 14 12 9 1 9 1 9 13 1 3 11 11 1 0 11 11 1 15 9 0 13 4 4 2
52 9 11 11 7 9 11 11 1 9 1 12 9 1 15 9 1 11 1 0 9 13 1 11 1 9 0 13 9 1 0 13 4 13 16 15 15 9 14 13 16 11 9 1 13 0 9 1 9 1 0 13 2
26 9 1 1 10 9 7 9 1 9 1 15 0 13 4 16 9 1 13 9 1 15 0 9 13 4 2
9 9 1 1 11 14 0 9 13 2
33 9 1 13 9 1 9 1 9 1 13 4 9 1 3 13 16 16 11 1 9 14 13 4 16 0 7 0 9 1 9 13 4 2
17 9 1 1 9 1 9 9 1 0 9 1 0 9 1 9 13 2
15 3 15 0 9 1 9 1 10 1 9 14 13 4 4 2
64 9 1 11 11 1 9 0 9 1 9 13 4 9 1 9 13 11 11 11 1 11 2 11 1 1 9 1 1 13 4 9 1 13 1 9 1 12 9 1 0 9 7 12 12 9 9 1 9 13 7 9 14 13 1 12 9 1 0 9 1 9 14 13 2
25 9 1 9 1 0 9 1 15 14 13 16 9 1 9 1 11 7 11 1 0 13 4 4 4 2
29 0 13 16 11 9 1 1 1 0 9 11 11 7 9 1 1 1 0 9 11 11 1 9 1 15 9 13 4 2
20 9 1 13 0 9 1 12 9 1 9 13 4 4 7 12 9 0 13 4 2
10 10 9 1 12 9 14 13 4 4 2
8 9 1 9 9 13 4 4 2
13 12 12 1 10 0 9 9 9 1 9 1 13 2
15 9 9 9 7 9 9 9 9 1 9 14 0 14 13 2
23 9 11 2 11 1 9 1 1 12 9 9 9 7 12 9 9 9 9 1 9 13 4 2
30 0 9 1 9 10 12 0 9 9 1 9 9 1 9 13 1 7 14 9 13 4 4 7 15 9 0 13 4 4 2
30 9 1 13 4 12 9 1 9 13 4 11 11 11 11 1 13 16 9 1 1 15 14 9 1 0 14 13 4 4 2
62 7 9 9 1 12 9 9 9 9 2 11 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 7 11 2 11 2 1 15 13 0 9 1 1 9 13 1 9 13 4 4 2
35 11 1 13 16 0 12 9 1 1 11 11 2 11 11 11 7 11 11 11 11 11 1 13 0 9 1 15 14 9 1 9 14 13 4 2
10 11 11 1 9 1 3 9 13 4 2
15 9 1 0 9 1 0 13 1 10 9 1 0 9 13 2
16 11 11 11 7 11 11 11 11 11 1 9 1 9 13 4 2
25 11 11 1 13 16 9 1 1 0 7 0 9 1 15 14 9 9 1 9 13 0 14 13 4 2
33 11 1 11 11 11 1 15 9 13 4 11 1 0 13 4 16 15 9 9 1 11 1 11 1 9 1 0 13 1 9 1 13 2
34 11 1 11 1 10 9 1 9 13 4 7 11 11 11 11 1 11 1 9 13 4 4 16 11 11 1 14 0 9 15 0 14 13 2
18 11 1 9 11 11 11 11 2 7 9 1 9 11 11 1 9 13 2
9 11 11 11 11 14 11 1 13 2
37 11 11 1 9 1 9 13 16 11 1 9 1 1 11 1 13 16 11 1 16 9 9 1 0 9 0 13 4 16 15 11 1 14 9 13 4 2
18 9 9 1 15 2 0 9 2 1 9 1 1 1 14 13 4 4 2
14 15 13 16 15 14 11 11 1 0 9 14 13 4 2
22 9 1 13 16 11 1 13 16 9 15 9 9 9 1 9 9 1 0 13 1 13 2
28 11 1 9 13 16 9 9 1 0 9 1 11 11 1 0 13 9 1 11 11 1 9 7 9 10 13 4 2
14 15 9 11 1 9 1 1 12 0 9 0 13 4 2
21 11 1 1 11 7 11 11 11 1 11 1 0 9 1 1 1 9 2 9 13 2
29 9 1 13 4 16 11 1 11 1 11 11 1 1 11 1 10 9 1 11 1 11 11 11 1 14 9 13 4 2
15 15 1 1 12 9 1 9 15 1 10 9 13 4 4 2
18 7 12 9 1 1 10 9 9 1 13 4 15 0 13 4 4 4 2
25 11 1 3 0 9 11 11 1 9 1 11 11 11 11 1 12 9 9 13 1 9 13 4 4 2
28 0 9 1 11 11 1 9 9 1 1 1 11 1 0 0 9 1 9 1 1 9 9 9 13 1 0 13 2
11 10 0 9 1 9 9 12 12 9 13 2
14 15 13 16 11 11 11 1 1 11 12 0 9 13 2
12 9 14 9 12 12 9 9 1 9 13 4 2
21 2 11 9 12 9 1 1 9 14 0 13 7 15 0 9 1 13 1 9 13 2
20 16 9 1 15 14 9 10 9 1 13 1 0 13 16 15 1 12 0 9 13
38 11 1 0 2 11 11 11 2 1 13 9 1 1 2 9 9 13 1 1 9 0 13 2 7 9 1 1 11 1 11 1 0 9 1 0 9 13 2
44 9 1 1 2 11 10 9 1 1 9 1 9 13 4 4 16 9 1 10 9 7 9 1 1 9 1 9 13 1 9 1 1 15 9 1 0 9 1 3 9 1 13 4 2
16 0 13 16 10 9 1 9 1 9 1 9 9 1 10 13 2
21 11 1 1 9 1 9 14 10 13 15 1 0 9 9 1 9 1 9 13 4 2
26 15 13 2 2 15 1 9 9 1 9 1 9 1 1 1 15 14 13 4 2 7 15 9 13 4 2
13 15 9 1 9 13 7 0 9 1 14 9 13 2
32 15 14 15 14 13 4 16 9 1 10 9 15 1 13 2 7 12 9 14 3 13 16 9 9 1 0 9 8 13 4 4 2
20 9 1 10 9 1 0 13 1 1 15 1 12 9 1 0 9 9 13 4 2
23 9 1 9 1 9 1 1 14 0 13 4 1 9 1 9 9 14 13 1 9 13 4 2
22 16 2 9 9 13 15 0 13 4 4 16 9 1 9 2 9 14 9 1 0 13 2
34 10 9 1 10 9 0 13 4 9 11 11 1 13 13 16 0 0 9 15 9 1 0 9 7 15 0 13 1 1 1 15 14 13 2
14 15 0 14 13 16 10 9 9 1 1 0 14 13 2
14 11 9 9 1 0 13 7 15 9 1 9 13 4 2
15 15 13 16 10 9 15 0 14 12 9 1 13 4 4 2
13 10 9 1 9 15 15 9 9 1 1 13 4 2
14 15 15 14 15 0 9 13 4 15 15 9 13 4 2
20 11 1 9 13 16 15 14 9 1 1 1 15 9 12 9 1 0 13 4 2
20 15 15 9 1 1 1 9 13 1 3 9 2 9 7 9 1 9 13 4 2
17 15 1 15 0 9 1 9 1 9 7 9 1 1 1 13 4 2
20 9 11 11 15 14 15 1 0 13 4 15 15 0 9 9 1 0 13 4 2
15 15 0 9 13 16 9 9 2 9 1 10 9 13 4 2
18 11 1 13 16 11 15 9 13 7 15 1 15 9 3 0 13 4 2
27 15 1 13 9 1 9 13 11 1 13 4 9 0 13 4 7 10 9 9 1 1 3 9 13 4 4 2
30 12 0 9 11 11 14 15 15 0 9 9 13 4 7 15 0 9 13 4 15 15 0 9 9 1 14 0 13 4 2
30 15 13 4 16 9 15 9 1 10 9 1 15 9 13 4 4 16 3 0 9 1 9 1 15 15 14 9 13 4 2
11 11 14 15 1 1 11 1 9 13 4 2
34 12 0 9 9 1 13 13 16 9 1 9 1 3 0 14 13 4 4 2 7 14 15 9 1 14 15 1 9 13 14 0 14 13 2
11 9 1 13 14 9 13 4 9 9 1 2
30 9 15 13 16 9 1 12 1 9 9 1 13 4 1 9 15 13 2 9 9 1 2 9 9 1 7 9 9 1 2
28 9 9 1 9 0 0 0 13 2 10 9 1 9 15 14 0 0 13 2 15 15 9 13 9 13 4 4 2
10 3 9 9 1 9 1 1 15 13 2
45 11 11 1 9 11 1 1 9 9 1 10 0 9 1 1 0 0 9 1 0 9 2 9 2 9 7 9 9 1 9 1 9 7 9 7 9 9 1 9 1 9 1 9 13 2
12 9 9 1 9 1 15 0 9 14 13 4 2
15 9 7 9 9 1 9 15 14 9 1 9 13 4 4 2
16 15 9 2 9 7 9 9 1 9 1 9 13 4 4 4 2
50 11 11 11 1 9 11 11 1 1 15 9 10 9 1 13 15 2 9 9 2 1 0 9 13 4 4 4 16 0 9 1 2 15 1 14 9 1 10 9 9 9 7 9 1 9 13 1 13 4 2
11 9 1 1 2 11 1 0 11 1 13 2
11 9 1 15 9 1 0 9 14 13 4 2
25 7 16 11 1 11 1 9 9 1 13 4 0 13 4 16 0 9 1 1 9 13 1 13 4 2
13 9 9 1 9 9 9 11 1 14 0 13 4 2
19 9 9 1 10 9 1 9 1 0 9 13 2 15 9 13 4 4 4 2
24 11 11 11 1 9 9 11 11 13 4 2 2 9 1 9 13 1 9 1 12 9 3 13 2
14 9 1 9 9 1 13 1 9 1 0 9 13 4 2
18 2 9 1 9 13 14 10 9 9 0 0 9 1 9 13 4 4 2
7 9 1 9 1 14 13 2
10 9 1 9 15 13 15 9 0 13 2
10 10 9 9 9 1 11 1 14 13 2
46 9 1 1 2 16 15 9 9 10 9 1 9 9 8 13 4 15 9 9 1 9 10 9 1 13 16 9 1 13 14 9 1 11 0 9 1 10 13 4 7 15 9 13 9 13 2
14 9 0 0 9 1 1 9 1 0 9 3 0 13 2
7 15 0 9 9 1 13 2
13 9 1 10 9 1 9 1 9 0 13 4 4 2
26 15 1 9 9 0 9 13 1 15 9 1 13 4 4 7 15 10 9 0 9 1 0 13 4 4 2
29 9 14 1 15 1 13 9 9 1 12 9 10 13 2 7 9 1 9 13 16 15 12 9 1 10 9 14 13 2
13 7 0 9 1 15 15 0 0 14 13 4 4 2
24 9 9 1 13 16 16 0 9 14 9 13 16 9 1 10 9 1 0 0 13 4 4 4 2
30 10 3 9 14 13 1 1 9 1 3 15 9 13 9 13 4 7 10 9 1 9 12 9 9 1 3 13 4 4 2
32 9 9 1 1 11 1 11 1 12 9 1 9 14 1 10 12 9 9 13 4 7 10 9 1 1 12 9 0 9 13 4 2
10 15 15 1 10 12 9 1 9 13 2
26 0 9 15 12 9 1 9 13 7 13 0 9 9 14 13 1 1 15 12 9 1 10 9 13 4 2
32 11 11 2 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 7 9 1 10 9 1 9 1 10 9 13 4 2
13 15 10 9 1 9 1 0 9 13 1 9 13 2
10 9 1 3 0 9 0 9 1 13 2
9 0 11 1 14 12 9 9 13 2
26 16 15 13 9 0 13 4 4 15 15 3 10 13 4 7 3 14 12 9 9 15 1 13 4 4 2
20 15 1 0 11 11 1 9 3 0 13 15 9 1 12 9 10 9 13 4 2
21 10 9 1 10 12 9 9 0 13 4 4 7 15 1 9 12 9 9 13 4 2
14 0 12 9 1 1 0 11 11 1 9 0 13 4 2
17 15 9 12 9 1 1 12 9 9 13 4 15 12 9 10 13 2
20 0 9 0 11 11 1 9 14 13 7 10 9 1 14 12 9 9 13 4 2
8 16 0 9 12 9 0 13 2
16 7 0 11 11 1 12 9 9 13 16 12 9 9 13 4 2
27 9 1 1 11 11 1 9 1 12 9 1 12 1 1 12 9 9 13 4 15 9 1 12 9 10 13 2
18 11 1 12 1 1 12 9 9 13 4 15 9 1 12 9 10 13 2
13 0 11 1 1 0 11 1 9 14 0 14 13 2
12 0 11 1 9 1 12 9 10 9 13 4 2
11 15 12 1 1 14 12 9 9 13 4 2
24 11 1 12 9 9 13 4 7 10 9 1 12 9 9 13 4 15 9 1 12 9 10 13 2
13 9 1 9 1 9 12 9 1 10 13 4 4 2
11 7 0 9 15 12 9 1 14 13 4 2
16 11 1 9 1 9 1 12 9 9 1 9 0 13 4 4 2
11 11 1 11 1 0 9 12 9 9 13 2
8 11 1 9 12 9 9 13 2
23 9 9 1 9 13 16 0 12 2 12 9 9 15 14 13 16 9 13 1 9 13 4 2
18 11 11 11 11 1 11 1 9 1 9 1 3 15 9 0 13 4 2
9 10 9 10 12 9 9 8 13 2
11 9 12 9 7 9 12 9 8 13 4 2
8 9 1 0 9 11 1 13 2
13 9 9 9 7 9 1 14 0 13 4 4 4 2
9 15 1 9 1 0 9 13 4 2
27 9 9 1 9 11 11 1 11 1 15 13 16 10 9 11 1 9 12 9 1 14 0 13 4 4 4 2
15 11 1 9 1 10 12 12 12 12 12 9 0 13 4 2
17 10 9 1 1 12 12 12 12 12 0 13 7 12 1 9 13 2
16 12 12 12 12 12 9 1 1 12 12 12 9 0 13 4 2
16 9 1 1 2 0 9 1 9 13 1 12 9 9 0 13 2
9 0 9 1 12 9 9 0 13 2
18 0 9 1 9 9 12 13 4 2 7 0 9 1 0 9 12 13 2
46 9 1 13 16 11 11 1 0 9 1 1 0 9 1 9 12 9 1 0 9 1 10 9 13 4 4 7 0 9 1 1 0 9 9 9 1 9 12 9 1 9 9 13 4 4 2
18 0 7 0 0 9 13 1 9 1 0 9 15 15 9 13 4 4 2
19 0 0 9 1 1 13 4 1 11 11 9 1 0 9 15 11 14 13 2
22 10 9 11 1 0 9 1 0 0 0 7 0 9 1 9 1 13 4 13 4 4 2
34 11 11 9 1 9 1 9 13 1 0 9 2 11 11 11 2 2 11 2 1 0 13 4 16 15 11 14 15 9 1 0 9 13 2
15 15 1 14 10 9 1 9 9 14 11 1 14 13 4 2
20 9 1 15 14 9 1 9 13 1 11 11 11 10 9 1 1 9 13 4 2
19 15 9 11 1 13 1 9 1 10 13 2 16 15 9 3 0 13 4 2
33 11 11 11 2 11 2 9 14 1 9 9 1 9 1 9 2 9 13 1 9 11 11 2 11 2 1 0 2 0 0 9 13 2
15 11 1 9 1 9 15 9 9 9 11 11 1 15 13 2
25 15 1 10 9 1 3 11 11 9 1 13 1 0 9 10 13 3 11 1 9 1 9 14 13 2
20 9 9 1 13 13 16 10 9 1 0 0 0 9 1 10 9 13 4 4 2
20 15 9 1 13 7 15 9 1 1 15 9 13 7 9 13 1 14 9 13 2
16 15 1 9 1 1 15 9 1 1 10 9 1 9 13 4 2
36 3 14 11 11 9 15 14 9 7 9 8 13 4 4 2 7 15 9 0 0 9 1 9 13 1 9 7 9 13 1 9 1 1 13 4 2
45 11 9 1 0 0 9 1 9 13 1 11 1 11 1 9 11 11 1 12 9 11 11 2 11 2 2 11 11 11 11 2 11 2 7 11 11 2 11 2 9 1 13 4 4 2
28 11 13 9 11 1 11 13 4 7 15 9 1 13 1 3 12 9 9 15 11 11 11 11 11 1 13 4 2
19 15 15 1 9 13 16 9 7 3 1 10 9 1 15 9 13 4 4 2
14 7 15 11 0 9 1 9 9 0 13 4 4 4 2
16 15 0 9 1 16 13 4 16 11 1 15 9 14 13 4 2
8 15 15 9 1 9 1 13 2
19 10 3 9 1 11 1 12 0 0 9 1 11 13 1 14 9 13 4 2
19 10 9 1 9 1 10 9 13 4 2 15 15 7 15 9 1 13 4 2
18 11 11 1 9 12 9 11 11 1 9 1 0 9 9 1 13 4 2
18 15 1 12 9 1 9 1 15 8 13 4 7 0 9 1 13 4 2
23 9 13 1 11 0 9 1 15 9 11 11 1 13 11 10 9 15 9 1 0 14 13 2
13 15 11 1 14 13 2 7 10 9 0 14 13 2
18 15 0 9 1 10 9 1 0 13 16 11 1 9 13 4 4 4 2
7 0 9 9 1 3 13 2
17 10 9 13 16 11 1 13 1 1 15 9 1 1 14 13 4 2
15 16 9 1 0 9 1 15 1 1 9 13 4 4 4 2
15 15 10 9 9 1 15 9 2 9 2 1 0 9 13 2
35 15 9 1 9 9 13 4 1 1 11 9 1 9 9 11 11 1 13 16 11 1 9 7 9 1 0 9 11 1 9 1 13 4 4 2
6 15 9 13 4 4 2
40 0 13 16 11 1 0 11 11 11 11 1 11 9 1 9 1 0 9 13 11 1 11 11 11 1 13 4 11 11 11 11 11 1 9 13 1 9 13 4 2
25 11 11 1 9 11 11 1 13 16 12 9 1 11 1 9 1 10 9 1 9 2 9 13 4 2
15 11 1 1 9 1 9 0 13 1 9 13 4 4 4 2
12 16 12 9 9 2 9 1 9 13 4 4 2
15 9 1 10 0 9 14 13 1 9 1 11 1 9 13 2
27 9 1 1 11 11 1 12 9 0 9 11 11 11 1 9 1 0 9 1 9 13 11 0 13 4 4 2
20 11 2 11 1 11 11 1 11 9 1 9 1 1 1 11 1 9 13 4 2
20 9 1 1 10 9 1 15 9 13 4 2 10 9 1 10 9 14 9 13 2
31 11 11 1 12 9 1 13 16 0 9 1 9 1 13 1 1 15 10 14 10 9 1 13 9 1 0 13 1 9 13 2
48 11 1 9 1 9 1 9 1 13 4 16 11 1 11 11 1 13 4 1 11 11 11 11 11 1 9 1 11 1 13 9 1 15 9 11 7 15 9 11 11 1 1 11 11 14 0 13 2
15 7 11 11 1 13 4 16 11 10 9 1 0 14 13 2
13 9 9 1 1 9 1 9 1 9 13 4 4 2
19 9 1 0 9 1 13 9 1 11 1 0 2 0 9 1 9 13 4 2
17 11 1 11 1 9 1 9 13 4 9 13 4 9 1 13 4 2
11 15 9 1 9 1 9 1 9 13 4 2
31 10 3 9 9 1 13 9 1 11 9 11 1 11 11 0 9 9 1 3 9 13 7 9 7 9 9 1 1 9 13 2
11 11 9 1 10 9 1 9 1 9 13 2
30 0 13 16 9 9 1 13 9 1 11 1 11 9 1 9 13 4 4 2 7 11 1 12 9 1 9 13 4 4 2
35 9 9 1 0 11 1 11 1 9 1 0 9 1 9 13 1 9 9 1 0 13 1 9 1 9 1 11 1 0 9 1 9 13 4 2
24 0 13 16 11 1 9 1 11 1 9 9 1 13 12 9 1 0 9 1 9 13 4 4 2
44 9 1 10 9 1 11 1 14 12 9 1 1 0 9 9 13 2 9 9 1 1 9 1 0 13 7 9 9 1 9 1 13 1 9 13 1 9 11 9 1 0 13 4 2
29 13 4 4 16 11 1 10 9 1 9 7 9 9 1 9 13 2 15 15 14 12 9 11 13 1 9 13 4 2
18 7 15 9 1 14 13 1 14 12 9 9 1 0 9 9 13 4 2
10 14 12 9 9 1 3 9 13 4 2
11 15 1 9 1 9 1 9 9 13 4 2
18 9 1 14 15 9 9 1 13 7 9 13 9 1 15 1 13 4 2
7 9 1 9 13 4 4 2
12 9 1 11 11 1 12 9 1 9 13 4 2
27 9 1 9 13 1 9 9 11 1 9 11 11 9 2 9 1 1 9 1 13 7 9 13 1 9 13 2
13 15 1 9 7 13 9 1 1 0 9 14 13 2
13 0 9 9 2 9 13 1 9 1 0 13 4 2
17 13 9 1 9 1 13 1 9 13 1 10 9 1 9 13 4 2
8 15 9 1 9 13 9 13 2
47 3 9 2 9 1 9 1 13 0 9 9 1 9 11 11 11 1 9 1 12 9 1 9 1 11 2 11 9 0 11 11 11 11 1 1 9 12 9 1 9 12 9 1 9 13 4 2
24 9 9 1 9 9 11 11 11 9 1 13 7 11 11 1 9 1 0 9 13 1 9 13 2
36 10 3 9 9 1 13 9 1 11 9 12 9 11 1 11 11 0 12 9 9 9 9 1 3 9 13 7 9 7 9 9 1 1 9 13 2
14 9 1 9 1 9 1 9 7 9 1 0 13 4 2
10 9 1 15 9 9 9 9 1 13 2
25 9 1 9 1 13 9 1 9 13 1 9 13 2 7 13 9 1 9 9 1 1 14 9 13 2
20 9 1 13 9 11 11 7 0 9 1 9 2 9 13 9 1 0 13 4 2
16 9 1 10 9 1 12 2 12 9 1 1 9 0 13 4 2
31 11 11 1 11 1 11 11 1 11 11 1 11 11 1 11 9 1 9 1 9 13 1 9 1 9 13 4 9 0 13 2
42 9 9 11 11 11 1 9 1 9 1 1 11 1 11 9 1 9 1 11 1 9 9 1 1 11 1 0 9 9 1 9 1 9 13 1 9 1 15 9 13 4 2
12 9 1 13 16 0 9 1 3 14 9 13 2
27 9 1 11 11 1 9 11 11 11 11 1 12 0 9 9 1 11 1 3 9 13 1 9 0 13 4 2
25 11 1 13 16 9 1 0 13 4 4 4 7 15 1 11 1 9 13 1 9 13 4 4 4 2
19 15 1 11 11 1 9 1 10 9 1 11 1 9 9 9 13 4 4 2
22 11 1 11 9 1 0 9 9 1 0 13 1 3 10 9 1 9 1 9 0 13 2
15 9 1 11 1 11 11 1 0 9 1 13 1 9 13 2
28 11 11 1 11 1 9 13 1 12 9 1 9 1 1 9 1 9 13 7 13 1 9 1 0 13 4 4 2
15 0 9 9 1 11 1 11 1 9 13 1 3 0 13 2
34 11 11 11 2 11 2 1 9 11 11 1 11 1 9 13 16 15 1 12 9 1 11 1 9 1 0 9 1 9 9 1 9 13 2
38 11 1 13 16 11 11 2 11 1 11 11 11 11 1 1 13 9 1 0 13 9 9 11 1 9 1 12 9 1 0 9 1 1 0 13 4 4 2
20 11 1 1 11 1 9 1 9 1 12 1 12 9 1 13 4 1 9 13 2
11 15 9 9 9 9 7 11 9 9 13 2
36 16 11 1 9 0 13 16 11 1 0 9 1 9 1 9 9 3 13 4 4 2 16 15 13 16 10 9 11 7 11 9 1 1 0 13 2
47 15 15 13 4 16 9 9 1 10 9 11 11 1 15 13 4 2 15 15 13 16 11 1 13 9 1 9 9 1 13 9 1 9 11 9 1 8 13 7 11 11 9 11 11 1 13 2
16 11 1 10 9 1 14 1 11 1 14 10 14 9 13 4 2
8 10 0 9 1 9 11 13 2
20 0 9 1 1 10 9 13 10 9 9 1 12 12 1 10 9 0 13 4 2
28 11 1 9 1 13 16 10 9 9 9 13 4 10 9 1 10 9 14 13 0 9 1 9 13 9 1 13 2
14 15 13 16 9 9 0 9 1 0 9 1 14 13 2
8 15 0 9 11 11 9 13 2
22 11 2 11 9 1 13 4 0 9 1 10 9 13 15 0 9 11 11 11 14 13 2
17 11 0 11 11 11 1 9 1 9 1 1 11 1 10 9 13 2
46 11 11 11 11 2 11 2 1 9 11 11 11 11 1 9 1 13 16 15 11 2 11 9 1 13 4 9 1 9 13 7 10 9 1 13 16 9 1 13 4 9 11 11 14 13 2
18 10 9 11 1 11 2 11 9 1 0 9 11 11 1 13 4 4 2
24 9 1 0 9 13 1 9 1 11 11 7 12 9 9 1 11 11 2 11 1 0 13 4 2
10 3 1 15 9 1 0 13 4 4 2
24 9 1 1 9 1 1 11 11 13 13 4 2 7 11 2 11 9 1 15 15 9 14 13 2
16 9 1 9 1 1 11 1 11 11 1 11 11 1 9 13 2
26 11 1 1 1 11 11 1 0 9 9 0 13 11 11 1 9 1 9 1 9 13 1 9 13 4 2
24 12 0 9 1 11 1 11 13 1 9 13 4 4 2 7 9 1 15 1 9 13 4 4 2
30 11 1 11 11 11 7 11 11 11 1 9 9 7 0 9 1 0 13 1 9 13 1 1 11 13 1 9 13 4 2
23 9 1 9 1 13 4 11 1 9 11 13 7 11 11 11 7 11 11 11 1 9 13 2
24 9 9 13 1 3 9 9 1 9 12 0 9 13 7 9 1 3 1 9 1 9 0 13 2
6 15 9 1 13 4 2
14 15 13 16 9 9 1 9 1 15 10 9 13 4 2
17 15 1 14 15 13 16 15 9 1 9 13 1 1 9 0 13 2
11 15 10 9 1 11 11 1 13 4 4 2
26 15 13 16 9 1 10 9 1 10 9 13 16 11 11 11 1 3 3 10 9 1 15 9 13 4 2
36 15 13 16 9 1 1 13 1 1 9 1 11 11 1 9 11 1 9 1 9 13 2 16 10 9 1 0 9 1 9 13 9 1 9 13 2
20 9 7 9 9 1 15 3 13 4 16 15 3 15 9 1 9 13 4 4 2
16 11 11 11 1 1 14 13 4 2 10 15 14 13 4 4 2
26 9 1 0 9 15 9 1 9 9 13 1 1 9 11 1 11 11 1 2 11 11 11 2 1 13 2
17 7 2 15 9 9 1 9 1 3 1 10 9 3 13 4 4 2
12 9 1 9 8 9 1 14 10 9 13 4 2
11 15 9 1 13 9 1 15 9 14 13 2
11 9 1 10 9 9 1 13 9 1 13 2
11 11 1 0 9 1 11 9 13 4 4 2
16 15 12 9 1 9 1 9 1 3 13 13 1 9 14 13 2
15 12 9 1 9 1 9 1 9 9 13 1 0 14 13 2
16 9 1 13 4 15 15 0 9 1 9 1 9 3 13 4 2
23 9 9 2 9 1 9 13 16 9 1 13 1 3 9 15 0 9 1 14 0 13 4 2
30 9 1 10 9 15 9 1 1 9 13 1 1 0 13 4 15 14 13 14 7 9 1 15 11 1 9 14 14 13 2
30 15 9 13 16 10 9 1 9 1 0 9 15 15 9 13 7 9 1 9 1 12 9 1 9 1 13 1 9 13 2
13 10 10 9 1 9 1 9 1 0 13 0 13 2
23 12 9 1 9 1 1 9 2 9 15 9 1 9 9 1 1 9 1 0 13 4 4 2
18 7 15 14 9 9 14 13 4 4 16 9 9 1 15 9 14 13 2
29 9 1 9 9 13 1 9 1 10 9 1 9 13 16 9 1 9 1 11 12 0 0 9 1 1 1 0 13 2
35 15 14 13 4 4 16 9 9 15 9 9 13 4 16 11 11 11 1 15 15 1 10 9 7 9 0 13 4 15 1 3 14 9 13 2
42 9 9 13 1 7 0 9 1 10 9 1 15 9 14 13 16 9 1 12 9 1 10 9 1 13 1 9 13 4 2 10 9 15 15 13 15 1 15 9 0 13 2
19 15 9 10 9 14 13 4 16 9 1 0 9 1 9 1 15 9 13 2
11 7 15 9 1 1 9 1 9 0 13 2
19 10 9 1 9 9 13 1 9 13 4 4 15 1 15 9 15 0 13 2
19 9 1 9 9 1 9 1 0 9 7 0 9 2 9 1 9 15 13 2
14 11 1 0 0 13 1 1 11 11 11 1 9 13 2
18 10 9 10 9 1 11 11 1 0 9 1 9 13 0 13 4 4 2
27 15 1 11 1 9 9 1 11 11 1 0 14 13 4 4 7 11 2 11 7 11 1 9 15 0 13 2
25 11 1 9 1 15 10 14 9 13 7 3 0 9 15 9 7 9 1 13 1 9 1 13 13 2
42 11 1 0 9 13 1 11 2 11 2 11 7 11 1 10 9 1 9 13 1 1 9 9 1 9 1 11 11 1 11 11 1 0 9 13 1 9 10 3 13 4 2
33 11 11 11 11 1 1 13 1 10 9 1 1 11 11 11 11 11 2 11 2 1 9 1 1 1 11 11 1 9 0 13 4 2
38 10 9 1 10 9 9 13 2 15 12 9 11 11 11 1 13 4 9 1 9 1 1 1 9 9 1 13 7 0 12 9 9 9 9 1 0 13 2
36 11 9 1 9 9 7 9 9 1 11 11 1 9 13 4 4 7 0 9 1 1 11 11 7 11 11 1 1 9 1 9 14 13 4 4 2
17 9 1 0 12 9 1 9 9 9 1 1 1 13 4 4 4 2
16 11 2 11 7 11 1 9 9 11 11 1 13 4 4 4 2
22 11 11 1 9 9 11 11 11 11 1 11 11 11 1 10 9 1 9 1 13 4 2
37 15 1 11 11 11 11 11 1 15 9 1 9 11 1 10 9 13 4 7 0 13 4 16 15 1 1 11 11 1 3 9 9 13 4 4 4 2
22 9 11 1 13 13 16 11 9 1 13 1 10 0 9 1 1 9 3 0 14 13 2
12 15 10 9 1 10 9 13 1 9 13 4 2
19 16 9 1 13 9 13 15 9 1 9 13 16 3 13 15 9 13 4 2
14 10 9 9 1 1 0 9 13 1 9 13 4 4 2
14 10 9 13 9 9 1 13 12 9 9 1 13 4 2
12 9 9 1 2 9 2 9 9 1 13 4 2
14 9 9 1 9 13 1 1 1 0 9 0 13 4 2
35 15 1 3 13 14 15 9 15 9 1 0 0 9 1 13 15 9 7 9 1 9 1 1 0 9 9 1 14 15 9 1 13 4 4 2
32 10 9 1 1 9 1 13 4 1 9 1 9 0 13 1 9 15 0 14 13 4 4 2 16 15 9 1 13 4 4 4 2
13 9 9 9 1 2 9 2 9 9 1 13 4 2
22 10 9 1 10 9 7 9 13 4 4 2 16 10 9 15 0 9 1 14 13 4 2
13 16 15 9 1 11 11 13 16 13 13 4 9 2
19 9 1 11 9 1 13 7 13 4 15 9 2 9 7 9 1 0 9 2
25 15 14 10 9 1 9 13 1 9 13 16 9 2 9 13 1 1 3 14 10 9 1 9 13 2
23 10 9 1 15 8 13 8 13 2 10 9 9 9 1 1 9 2 9 9 1 13 4 2
19 15 15 9 13 1 9 2 9 7 9 13 1 9 14 0 13 4 4 2
20 11 11 1 13 16 11 7 0 9 1 0 2 0 9 1 9 0 13 4 2
18 9 1 0 9 1 15 0 9 1 9 2 9 7 9 13 4 4 2
32 11 11 11 11 1 1 1 11 7 0 9 9 1 9 1 1 11 11 2 11 1 11 2 11 11 11 2 1 9 13 4 2
9 15 1 11 11 1 9 0 13 2
40 9 9 9 1 9 1 1 11 11 11 11 11 1 9 0 10 9 11 2 11 2 11 7 11 1 0 11 1 9 1 12 9 0 0 9 1 0 13 4 2
31 11 11 1 0 13 1 11 1 9 2 11 11 2 1 9 1 11 11 1 0 12 9 1 9 9 13 1 13 4 4 2
28 11 11 11 11 1 9 1 11 1 12 0 9 1 1 0 9 11 11 11 11 1 9 1 14 9 13 4 2
9 9 11 11 7 11 1 1 13 2
12 11 9 9 1 1 11 1 0 9 13 4 2
18 15 9 1 14 9 13 4 7 10 0 9 1 9 14 13 4 4 2
10 9 1 1 9 9 1 9 13 4 2
21 11 1 9 1 0 0 9 1 9 13 12 0 11 11 0 9 14 11 13 4 2
19 15 3 11 11 1 1 13 4 7 10 9 1 15 11 1 1 13 4 2
13 11 1 0 9 1 15 9 1 1 0 9 13 2
19 15 1 0 9 1 0 9 13 1 3 15 9 1 13 9 1 1 13 2
11 11 1 9 11 11 14 9 1 1 13 2
16 11 9 1 13 7 10 3 3 11 1 9 15 9 1 13 2
7 15 9 1 0 13 4 2
10 15 1 15 12 0 9 13 4 4 2
10 15 9 1 9 1 0 0 13 4 2
20 11 9 1 0 9 9 11 1 13 16 9 1 9 9 1 1 14 9 13 2
30 11 11 1 9 11 11 1 15 13 16 15 10 9 1 3 0 13 7 15 1 15 14 13 4 1 9 1 14 13 2
16 11 1 0 9 13 9 13 16 9 1 9 9 1 9 13 2
33 15 1 14 11 11 1 15 14 13 16 15 9 9 1 9 1 10 15 9 1 0 13 1 1 0 0 9 13 1 15 14 13 2
26 11 11 1 0 9 1 1 0 0 9 13 1 1 0 0 9 7 15 0 9 1 9 0 13 4 2
36 0 0 9 1 9 1 0 9 1 9 2 0 9 1 9 2 0 9 7 9 1 9 1 9 1 9 13 1 1 0 9 1 0 13 4 2
31 9 1 15 0 2 0 13 4 4 16 11 9 2 9 2 0 9 2 0 9 7 9 1 9 7 9 1 9 13 4 2
32 11 11 1 10 9 1 15 14 0 13 4 16 11 9 1 1 11 11 1 0 0 11 1 13 9 1 9 1 13 4 4 2
31 11 1 1 15 9 13 1 9 1 1 11 11 1 11 2 11 1 0 15 12 12 9 1 0 9 1 0 13 4 4 2
36 9 1 0 0 9 1 11 1 15 9 13 4 13 16 15 1 12 9 7 9 0 13 1 3 2 9 10 9 1 14 9 0 13 4 4 2
28 10 9 1 11 1 2 11 11 2 1 1 1 14 13 4 4 7 15 15 0 0 9 1 13 4 4 4 2
11 9 1 10 9 1 9 1 9 13 4 2
22 11 1 11 1 11 1 13 1 0 9 9 1 1 11 1 9 9 11 13 4 4 2
12 3 0 9 1 14 11 13 9 13 4 4 2
9 9 14 12 12 0 9 11 13 2
12 11 1 9 11 1 9 15 9 13 4 4 2
25 11 13 1 3 11 1 9 3 11 11 11 2 11 2 11 13 7 15 9 9 1 9 13 4 2
13 0 9 1 10 9 11 1 14 11 13 4 4 2
12 12 14 9 11 1 9 11 1 13 4 4 2
12 9 1 10 9 1 0 9 8 13 4 4 2
18 0 9 0 9 1 11 9 9 7 11 11 9 13 11 13 4 4 2
20 10 9 1 0 9 1 11 13 1 1 11 11 1 0 9 13 4 4 4 2
20 11 11 1 11 11 1 0 9 1 13 1 1 0 9 1 14 9 13 4 2
22 11 1 9 1 9 0 13 4 16 10 9 1 13 1 1 14 12 0 9 15 13 2
18 0 9 1 9 1 1 11 2 11 7 11 1 0 9 13 4 4 2
16 15 1 11 1 0 9 14 0 9 1 15 15 13 4 4 2
25 0 13 16 11 1 9 7 9 9 9 1 14 0 9 1 11 11 13 1 1 0 9 13 4 2
19 10 0 9 9 1 13 4 11 7 11 1 0 9 2 9 13 4 4 2
22 0 11 11 11 11 1 11 11 1 11 1 11 1 0 9 0 13 1 9 13 4 2
11 11 11 1 11 1 0 9 13 4 4 2
35 0 13 16 11 1 0 9 1 9 15 0 13 4 4 15 11 1 11 11 1 10 9 1 0 13 11 11 11 1 0 9 0 13 4 2
7 15 11 1 9 11 13 2
13 11 1 13 4 16 11 1 0 9 0 13 4 2
13 15 11 7 15 9 9 1 9 1 0 9 13 2
22 11 1 13 4 16 15 11 1 9 7 9 1 9 1 1 9 1 1 13 9 13 2
16 0 11 11 11 11 1 11 1 9 1 0 9 9 13 4 2
23 15 13 16 11 7 11 11 1 0 9 1 9 13 1 1 11 1 0 9 1 9 13 2
15 15 9 13 16 11 11 1 11 1 0 9 1 0 13 2
25 11 1 0 0 11 11 11 1 11 11 11 1 1 15 9 1 9 7 9 1 0 9 13 4 2
22 11 1 13 16 10 15 14 9 0 9 1 1 15 12 9 0 9 1 9 13 4 2
8 3 9 14 3 1 9 13 2
34 11 1 13 16 15 10 9 1 15 9 14 13 16 15 9 0 13 7 9 9 1 1 1 11 11 7 11 1 1 10 9 13 4 2
32 11 1 10 9 10 9 1 1 13 4 16 15 13 4 16 11 1 11 1 1 0 9 1 1 11 0 9 1 9 13 4 2
21 7 11 1 9 1 10 9 1 9 13 4 16 15 0 9 1 1 9 13 4 2
6 15 15 9 9 13 2
18 15 13 16 9 15 9 1 9 13 15 1 15 9 14 13 4 4 2
33 9 1 1 15 9 12 0 9 13 7 15 9 7 9 1 10 9 1 0 9 1 1 0 0 9 1 1 1 14 13 4 4 2
20 11 1 9 1 1 15 9 11 1 0 9 11 11 1 9 1 1 13 4 2
17 11 1 13 16 15 11 1 1 9 13 15 9 0 14 13 4 2
28 0 11 1 13 16 15 7 11 2 11 1 1 12 0 11 1 1 0 9 9 1 1 9 13 0 0 13 2
35 11 11 11 11 1 0 9 1 0 11 2 11 1 9 1 0 9 1 0 13 1 10 9 14 13 16 0 9 0 9 1 9 13 4 2
25 9 1 13 13 16 0 9 7 9 1 1 14 0 9 1 11 2 11 1 9 1 0 13 4 2
16 9 1 1 0 9 1 1 10 9 1 1 0 9 0 13 2
61 0 13 16 11 1 11 2 11 1 9 1 1 13 9 1 0 9 1 11 2 11 1 1 0 9 0 13 1 9 0 13 4 2 7 11 1 9 11 11 1 13 0 9 1 9 9 1 0 9 0 13 1 9 1 9 1 14 13 4 4 2
21 0 9 1 10 9 1 11 2 11 7 11 1 9 1 9 13 4 0 13 4 2
12 11 1 0 9 1 9 1 0 9 13 4 2
45 12 0 9 1 13 16 0 9 1 14 12 9 1 15 14 11 2 11 1 0 9 1 0 9 1 0 14 13 4 7 15 9 1 1 0 9 1 0 13 4 9 1 14 13 2
29 0 13 16 11 11 11 1 11 2 11 1 9 1 12 2 12 9 0 13 1 1 12 9 1 9 1 9 13 2
20 0 9 1 1 13 4 1 11 2 11 1 9 1 15 9 0 13 4 4 2
20 0 9 1 12 9 13 7 15 9 15 14 9 1 0 13 1 1 0 13 2
23 11 1 11 9 1 11 9 9 9 0 11 9 1 11 1 12 9 1 9 13 4 4 2
14 15 1 3 9 13 1 9 1 9 13 4 4 4 2
15 10 9 1 9 11 11 7 11 11 1 1 1 13 4 2
21 9 1 12 9 1 13 16 10 9 1 10 9 9 13 4 15 15 13 4 4 2
21 9 1 13 16 10 0 9 10 12 9 1 9 1 9 9 1 9 13 4 4 2
11 9 1 9 9 13 1 9 13 4 4 2
13 15 0 13 9 1 10 12 9 1 9 13 4 2
18 10 12 9 12 9 9 1 9 13 1 9 1 9 1 13 4 4 2
15 9 1 13 13 16 15 1 12 0 0 9 1 9 13 2
13 10 9 1 9 1 12 9 1 0 13 4 4 2
8 15 0 9 13 4 4 4 2
13 11 9 1 11 1 0 9 1 9 13 4 4 2
16 15 14 10 9 1 11 7 11 1 10 9 9 13 4 4 2
13 10 15 1 9 1 1 9 1 0 13 4 4 2
23 11 1 1 12 9 1 11 1 11 1 12 7 11 1 12 9 1 9 13 4 4 4 2
10 10 9 12 9 9 1 13 4 4 2
18 9 1 9 1 1 11 7 15 1 1 9 1 9 13 4 4 4 2
31 11 11 11 11 11 11 1 11 1 9 9 1 11 11 11 11 2 11 2 1 9 0 13 1 1 15 0 13 1 13 2
38 9 9 9 9 9 9 1 12 0 9 1 0 13 4 11 1 9 1 10 9 3 9 1 9 7 9 9 0 13 1 1 10 9 13 1 9 13 2
14 10 9 1 15 13 16 15 15 15 9 1 9 13 2
11 15 15 13 4 4 7 15 15 13 4 2
13 10 15 15 9 2 9 7 9 1 0 13 4 2
15 15 13 16 10 9 1 13 1 1 15 0 9 13 4 2
25 15 15 9 1 0 13 7 9 1 3 0 9 1 9 1 15 9 1 1 0 13 1 9 13 2
21 15 1 15 10 9 1 1 12 9 2 9 0 13 4 2 15 0 13 4 4 2
20 11 1 13 16 14 0 9 1 14 9 13 4 4 4 7 9 1 9 13 2
21 15 13 16 15 9 2 9 9 1 9 2 9 7 9 9 1 0 13 4 4 2
30 15 13 16 12 10 9 0 13 4 4 15 10 9 1 9 13 4 16 15 15 0 13 7 10 0 9 13 4 4 2
22 9 7 11 1 3 10 9 1 9 13 4 16 9 1 1 15 10 9 13 4 4 2
36 10 9 1 11 11 11 11 11 11 11 1 13 16 9 0 13 15 15 1 0 14 13 2 16 15 0 13 4 4 16 9 0 9 1 13 2
31 9 1 0 12 9 1 12 12 12 12 9 1 9 1 1 11 11 11 11 11 11 1 11 1 12 9 1 9 13 4 2
48 11 1 9 7 9 1 9 9 1 0 12 0 9 1 9 13 4 15 13 2 9 1 12 12 12 12 9 0 13 7 9 9 1 13 12 9 9 1 1 0 0 9 1 9 1 9 13 2
19 15 13 16 15 9 12 12 12 12 9 1 1 0 9 1 9 13 4 2
28 11 1 13 16 9 9 9 1 9 2 9 9 7 9 9 1 9 1 0 9 1 9 1 9 13 4 4 2
18 11 1 13 16 9 9 1 9 1 0 13 9 1 13 4 4 4 2
34 15 13 16 12 12 12 12 9 1 15 9 1 12 12 9 1 9 0 13 4 4 4 7 12 12 12 12 9 1 9 13 4 4 2
34 15 13 16 9 1 9 1 9 1 9 1 1 0 9 11 11 1 12 12 9 1 9 13 1 3 12 12 9 1 9 13 4 4 2
50 11 1 13 16 0 9 9 1 3 0 13 7 9 9 1 12 2 12 9 1 1 12 12 9 1 9 1 9 13 4 4 7 10 9 0 13 4 1 3 15 9 2 9 1 14 9 1 9 13 2
23 15 13 16 9 9 13 11 9 1 9 9 1 15 9 12 1 13 12 9 13 4 4 2
26 15 13 16 9 9 1 9 13 12 9 7 12 12 12 12 9 9 9 1 0 9 13 4 4 4 2
12 0 9 9 1 15 9 1 12 0 9 13 2
20 15 13 16 0 9 1 9 13 1 1 9 1 9 9 1 9 0 13 4 2
12 9 1 13 9 12 9 3 0 13 4 4 2
31 11 11 11 1 1 1 0 9 1 9 1 13 4 16 11 11 2 11 7 11 1 0 9 1 9 1 9 13 4 4 2
20 10 9 11 11 13 4 4 7 15 1 9 1 9 1 9 14 13 4 4 2
25 11 11 1 11 11 11 1 9 7 11 1 11 1 9 1 2 9 9 2 1 9 1 9 13 2
12 12 0 10 9 1 9 9 9 11 11 13 2
14 11 11 11 1 11 11 11 11 11 1 0 9 13 2
15 0 9 1 11 1 9 11 11 7 9 11 11 11 13 2
24 9 1 13 9 1 13 0 9 9 1 13 9 1 13 11 11 1 10 9 1 9 13 4 2
32 9 1 9 11 11 1 0 13 4 4 7 11 11 1 13 9 1 1 9 1 13 4 16 9 1 9 1 9 13 4 4 2
36 10 9 10 9 1 13 4 4 15 9 14 13 7 9 11 1 1 11 11 2 11 7 11 1 11 11 1 9 1 9 9 1 13 4 4 2
18 10 9 0 9 9 14 13 9 1 9 9 13 4 13 4 9 13 2
9 0 9 1 15 0 13 4 4 2
14 9 11 1 1 9 9 1 0 9 9 1 9 13 2
22 15 13 4 16 11 11 1 15 9 13 1 11 11 11 1 9 1 14 0 9 13 2
22 11 1 10 9 1 11 11 1 9 13 4 4 15 9 11 11 1 9 9 1 13 2
24 11 2 11 7 11 1 0 9 15 3 1 11 11 1 9 0 9 1 13 15 9 14 13 2
31 9 11 1 1 9 1 15 0 13 4 4 16 9 13 15 3 9 1 9 1 13 7 11 11 1 10 9 3 14 13 2
57 11 11 1 9 11 11 13 4 16 15 0 13 16 11 11 11 1 12 0 9 13 7 15 9 1 9 10 9 1 13 4 4 7 9 1 9 13 16 15 9 2 9 2 0 9 7 9 1 1 15 9 14 13 4 4 4 2
29 0 9 11 1 11 1 11 1 12 9 9 1 9 11 11 1 9 1 9 1 9 1 12 9 1 0 13 4 2
19 11 7 11 11 1 11 1 0 13 4 7 11 13 9 1 0 13 4 2
24 15 1 9 10 9 1 0 9 11 11 2 15 9 11 11 7 11 11 1 0 13 4 4 2
13 11 1 9 11 11 1 15 9 1 13 4 4 2
18 9 1 15 11 11 1 11 1 11 11 1 12 9 1 13 4 4 2
28 11 11 11 2 11 2 9 11 11 11 1 9 1 1 0 7 0 9 1 9 1 13 9 1 9 13 4 2
22 11 15 11 9 1 11 1 0 11 11 11 11 1 9 2 9 1 0 13 4 4 2
29 15 11 9 2 9 1 10 2 0 2 0 2 9 1 0 13 1 9 13 2 15 0 9 1 15 14 13 4 2
13 11 9 1 10 9 15 9 1 9 13 14 13 2
27 15 10 9 10 9 13 4 15 11 1 11 1 0 11 2 11 11 11 1 13 4 9 1 0 9 13 2
29 11 9 1 15 9 1 11 1 9 11 11 11 1 9 1 2 0 2 7 2 9 9 2 13 15 0 13 4 2
14 11 1 13 16 11 1 12 12 9 9 13 4 4 2
13 16 2 9 9 15 13 1 3 9 13 4 4 2
16 15 15 13 4 4 4 16 9 1 9 0 9 9 1 13 2
22 11 1 11 11 2 11 1 0 9 1 13 0 9 1 13 0 9 1 9 15 13 2
8 15 15 11 1 15 9 13 2
13 10 9 0 7 9 9 1 0 9 13 4 4 2
21 9 1 0 9 1 10 9 1 11 2 11 2 11 1 9 13 1 9 13 4 2
19 7 0 9 1 9 1 11 1 9 9 11 14 10 9 1 1 0 13 2
25 9 1 10 9 1 14 9 13 16 10 14 9 9 1 15 0 0 9 1 14 13 4 4 4 2
21 11 1 13 0 9 1 1 15 15 13 1 1 0 9 1 9 14 13 4 4 2
30 11 1 9 13 0 9 1 0 9 1 9 9 1 10 9 13 4 4 16 11 2 11 2 11 14 15 1 0 13 2
26 9 9 1 1 12 9 1 1 10 9 13 16 9 9 1 10 0 9 1 9 13 1 9 1 13 2
10 15 15 9 1 0 9 13 4 4 2
20 15 13 4 16 0 10 9 1 11 1 15 9 13 1 9 1 9 13 4 2
40 11 7 11 1 1 13 4 9 9 1 1 15 15 10 9 1 9 1 15 14 13 15 9 1 9 13 4 0 9 13 1 1 0 9 1 9 13 4 4 2
22 11 1 9 1 15 9 1 9 13 4 13 16 9 1 9 9 1 15 9 14 13 2
23 11 1 0 9 9 11 11 11 11 14 10 9 1 11 1 9 13 1 9 14 13 4 2
25 15 13 4 16 11 7 11 9 9 7 9 1 9 0 13 13 4 7 11 1 15 0 9 13 2
12 9 7 9 13 1 15 3 0 9 13 4 2
33 11 1 11 9 1 12 12 9 1 9 1 13 1 9 9 1 13 11 11 11 11 7 15 0 9 11 11 1 1 13 4 4 2
16 9 1 11 1 10 9 1 9 13 1 9 9 1 9 13 2
27 11 1 13 4 16 13 9 1 1 11 11 1 0 9 1 13 4 9 1 9 13 1 9 13 4 4 2
37 11 1 11 9 1 11 1 13 1 0 9 9 1 9 9 1 11 1 9 1 1 9 13 4 1 13 15 1 10 9 1 9 13 1 9 13 2
16 15 13 16 10 9 1 9 0 11 11 11 11 1 13 4 2
13 15 9 9 1 0 9 14 0 14 13 4 4 2
19 11 1 13 16 11 1 9 1 0 13 9 13 1 1 15 13 4 4 2
27 10 9 1 11 1 11 7 11 7 11 7 11 1 1 11 11 1 12 0 9 9 13 1 9 14 13 2
19 15 1 15 11 9 9 1 11 2 11 11 11 1 9 13 0 14 13 2
26 11 1 11 11 1 9 1 9 1 11 11 11 11 2 11 2 1 9 12 0 9 0 13 4 4 2
47 11 1 11 1 9 1 0 15 9 1 13 16 11 1 11 11 7 11 11 9 1 9 0 9 1 9 1 13 4 4 2 7 15 0 9 2 0 9 2 1 9 1 13 4 4 4 2
29 10 9 1 9 2 9 7 0 9 9 1 9 1 9 14 13 4 2 16 16 11 11 1 0 9 1 13 4 2
24 0 11 11 11 11 1 11 1 9 13 4 16 11 11 1 9 1 15 14 0 14 13 4 2
39 15 9 1 12 9 1 0 13 4 10 9 1 13 4 4 16 9 1 13 1 9 7 9 1 1 9 13 7 9 1 0 9 13 1 9 14 13 4 2
24 9 0 13 1 3 11 1 13 16 10 9 1 15 15 14 9 1 9 13 1 1 0 13 2
29 11 1 12 0 9 1 9 9 13 1 1 0 9 1 9 1 9 1 1 3 1 11 9 1 9 13 4 4 2
25 11 1 13 16 9 1 9 1 2 11 11 2 1 1 9 1 9 1 9 9 1 13 4 4 2
59 11 11 1 0 13 9 1 1 11 1 15 9 1 11 9 1 9 2 9 1 1 11 11 11 1 12 12 9 9 13 1 3 9 1 9 14 0 13 1 1 15 9 13 4 2 7 10 9 1 0 9 1 15 9 14 13 4 4 2
27 10 9 0 9 1 9 1 1 11 1 9 1 0 9 0 13 1 1 11 1 15 9 1 0 13 4 2
17 9 1 13 4 4 16 11 9 1 15 1 12 12 9 9 13 2
32 0 9 11 9 1 9 1 13 1 3 0 9 11 11 11 1 9 9 13 1 9 13 4 15 9 1 0 13 4 4 4 2
8 11 11 1 0 13 4 4 2
32 10 9 1 9 1 1 0 9 0 13 1 1 1 11 1 13 4 16 0 9 1 9 1 1 13 4 9 1 9 0 13 2
22 9 1 9 13 1 1 0 9 13 1 1 9 13 7 9 13 1 3 9 13 4 2
46 0 13 16 11 11 1 0 13 4 11 11 1 11 11 1 11 11 1 11 0 12 9 11 11 7 11 11 1 13 1 9 13 4 2 15 11 11 1 11 11 1 9 13 4 4 2
20 11 11 1 9 1 12 9 0 0 13 4 4 7 12 1 9 0 13 4 2
16 10 9 9 1 14 12 9 9 11 11 11 11 11 13 4 2
22 10 9 11 11 1 9 1 14 14 12 9 2 9 9 11 11 11 11 11 13 4 2
18 11 11 1 9 11 11 1 0 13 4 7 12 12 9 0 13 4 2
13 11 11 11 11 1 12 12 9 1 13 4 4 2
56 10 9 11 11 11 1 11 1 15 9 1 13 16 11 11 1 1 9 1 13 4 9 1 1 0 15 9 1 9 14 13 4 4 7 16 13 0 13 16 0 9 1 1 1 15 9 1 1 9 1 1 0 13 4 4 2
43 11 11 1 11 11 1 0 9 1 9 1 0 13 7 10 9 1 9 1 1 1 9 0 13 1 1 9 14 0 13 7 11 2 11 1 15 9 9 13 1 0 13 2
43 11 7 11 1 1 0 9 1 9 13 1 9 1 9 13 4 11 1 11 11 11 1 0 9 1 3 13 1 1 2 0 9 2 7 2 0 2 9 1 9 13 4 2
31 2 11 11 11 2 1 0 12 9 1 11 1 13 4 16 11 7 11 1 9 0 9 1 0 13 1 1 0 14 13 2
29 15 9 13 4 13 4 16 12 9 1 0 9 1 0 9 13 7 0 9 1 1 13 1 1 0 9 13 4 2
45 15 13 4 1 16 12 9 1 9 1 9 7 0 9 1 13 4 1 1 9 7 9 1 9 13 4 2 15 13 16 11 7 11 1 10 0 9 1 15 0 9 1 9 13 2
26 15 13 16 0 9 1 9 1 0 13 1 15 0 9 13 7 9 1 9 1 10 12 0 9 13 2
17 15 13 16 11 7 11 1 0 0 9 1 9 13 1 9 13 2
29 11 1 13 16 15 15 15 1 9 7 0 9 1 9 13 4 7 0 9 1 9 7 9 1 9 1 13 4 2
17 15 15 2 15 1 9 1 9 14 13 1 9 1 9 13 4 2
11 15 15 15 1 9 13 1 9 13 4 2
52 11 1 15 11 11 9 1 0 7 0 9 1 1 9 1 10 0 13 4 11 1 13 16 9 1 9 1 1 0 9 13 1 9 15 1 13 7 0 9 1 13 13 4 2 16 9 9 9 1 13 4 2
17 15 13 16 11 11 1 0 9 1 11 11 1 9 13 4 4 2
14 16 11 12 9 3 13 4 16 11 12 9 3 13 2
46 11 1 13 13 1 11 2 11 11 11 11 1 1 1 15 13 16 0 9 13 1 10 12 0 9 13 4 4 7 0 9 1 15 9 2 9 7 10 0 9 1 9 13 4 4 2
30 11 1 11 1 13 16 15 11 11 11 3 0 13 1 1 11 1 9 0 13 7 15 9 1 13 1 1 0 13 2
36 11 1 11 1 9 11 11 1 15 9 1 13 16 9 1 15 9 1 9 14 13 1 11 11 1 9 1 15 13 4 7 15 9 13 4 2
27 15 13 16 16 11 0 9 13 1 1 15 9 1 9 13 4 2 16 11 1 9 13 1 10 9 13 2
30 11 1 9 9 1 1 12 0 9 0 13 1 9 13 4 13 16 10 9 1 11 11 1 9 1 15 9 14 13 2
13 10 9 3 13 9 13 1 0 9 13 4 4 2
19 0 9 1 13 16 10 9 1 15 11 9 1 0 9 1 9 13 4 2
8 11 1 15 0 9 13 4 2
32 11 1 13 16 12 9 1 1 0 0 9 1 1 11 1 12 9 0 9 1 9 13 1 9 1 10 9 11 13 4 4 2
30 15 9 2 9 7 9 9 11 11 2 11 11 11 11 7 0 7 0 9 7 0 9 9 1 9 11 11 0 13 2
19 15 13 16 15 1 11 2 11 11 11 11 11 11 14 0 9 11 13 2
18 11 1 13 16 11 1 11 11 11 14 10 9 11 1 9 1 13 2
11 15 11 9 1 9 15 0 13 0 13 2
23 15 1 11 11 11 7 11 1 11 2 11 11 1 1 11 1 11 1 9 13 4 4 2
17 0 12 9 1 10 12 9 1 0 0 9 1 9 1 9 13 2
29 11 1 11 9 1 9 13 1 3 13 9 7 9 1 11 9 1 9 2 1 14 12 9 2 9 13 4 4 2
12 11 2 11 11 1 10 0 9 13 4 4 2
26 11 1 0 9 11 11 11 1 11 1 13 16 10 9 1 11 9 12 9 1 1 13 4 4 4 2
15 16 11 11 7 11 1 0 0 9 1 1 9 0 13 2
19 11 1 13 16 11 9 1 9 2 1 14 12 9 2 9 13 4 4 2
16 9 9 9 1 9 1 9 12 9 1 1 13 4 4 4 2
16 15 13 16 9 2 9 1 15 9 1 3 15 9 14 13 2
15 12 12 9 9 1 11 11 2 11 11 0 9 0 13 2
18 0 9 1 13 16 13 9 1 15 1 13 1 9 13 4 4 4 2
19 11 1 1 13 4 10 9 2 9 1 0 9 13 1 13 4 4 4 2
27 3 9 1 1 11 2 11 2 11 2 11 2 11 7 11 9 1 9 2 9 1 14 9 0 13 4 2
13 9 1 9 1 9 7 9 9 1 14 0 13 2
12 10 9 1 9 9 8 13 1 14 9 13 2
28 11 11 11 11 11 11 11 1 11 1 9 1 9 1 1 13 9 1 0 9 1 9 1 9 13 4 4 2
27 9 1 9 1 1 13 0 9 1 3 13 1 1 1 15 0 12 2 12 9 1 14 15 9 13 4 2
21 9 1 12 0 9 1 14 15 0 9 1 9 2 9 1 13 1 9 13 4 2
26 7 3 9 10 9 1 0 9 1 14 10 9 1 13 13 1 9 14 0 13 1 9 13 4 4 2
32 15 13 1 9 1 9 1 1 9 2 9 1 10 9 14 13 7 10 3 14 13 1 9 2 9 14 0 13 4 4 4 2
37 11 11 11 11 1 9 11 11 11 1 11 1 9 1 9 1 13 16 9 1 9 1 1 13 9 1 15 0 9 1 9 13 1 9 13 4 2
20 9 1 10 9 1 9 2 9 13 4 4 7 3 14 15 9 13 4 4 2
15 9 1 9 13 4 16 9 0 7 0 2 0 13 4 2
16 9 10 9 1 9 1 1 9 13 1 9 14 13 4 4 2
18 11 1 13 16 15 14 9 13 1 9 1 9 1 0 9 13 4 2
34 9 1 1 11 1 1 9 9 1 12 9 1 1 13 11 11 11 1 1 11 11 1 11 1 13 1 9 2 9 9 1 9 13 2
8 16 15 9 9 8 13 4 2
16 0 9 1 1 9 9 1 13 4 11 11 1 9 13 4 2
7 11 11 14 9 1 13 2
50 9 1 11 11 1 9 1 0 10 9 1 1 12 0 9 1 9 13 4 9 1 9 11 11 1 13 16 9 1 11 1 10 9 1 9 13 1 9 13 15 15 15 1 0 13 1 9 13 4 2
64 9 10 9 13 2 11 11 2 9 2 2 11 11 2 9 2 9 2 2 11 11 2 11 11 2 11 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 9 9 2 2
40 11 9 1 1 13 9 9 1 1 15 11 0 9 9 11 11 7 15 9 11 11 1 1 11 11 1 11 11 11 1 13 0 9 1 9 9 13 4 4 2
34 0 9 11 1 2 11 11 2 1 9 13 16 15 11 0 0 13 4 11 11 11 1 3 14 9 1 13 1 1 9 13 4 4 2
28 7 0 9 9 11 11 11 11 2 11 2 1 11 11 1 1 0 9 0 13 1 9 1 9 13 4 4 2
10 10 9 15 11 0 11 11 1 13 2
6 11 1 9 11 13 2
33 9 1 3 0 9 9 11 11 7 11 0 9 1 9 9 1 9 13 1 9 1 1 15 14 9 1 10 9 1 13 13 4 2
40 11 11 1 11 7 11 11 1 15 9 1 1 0 9 1 9 13 2 7 11 1 11 11 11 7 11 0 11 11 11 1 1 10 10 9 13 1 9 13 2
31 9 1 13 4 4 16 9 1 9 13 1 1 1 12 9 1 10 9 1 0 9 1 1 9 3 14 13 4 4 4 2
37 11 11 7 15 0 9 11 11 1 9 13 16 11 11 1 11 2 11 11 11 2 1 3 9 1 9 13 1 3 10 9 1 15 9 13 4 2
27 3 11 11 1 13 13 16 9 1 0 9 1 1 0 13 1 1 15 0 9 11 11 1 9 13 4 2
19 11 11 1 12 9 1 13 16 11 11 1 1 3 15 0 9 14 13 2
30 9 1 15 14 13 16 15 11 1 0 13 4 11 11 11 1 0 9 1 1 9 1 13 1 1 9 13 4 4 2
41 11 11 11 11 11 1 11 1 9 1 15 0 9 1 0 13 4 16 2 0 9 9 2 7 2 0 9 2 1 1 11 1 9 13 1 15 9 14 14 13 2
16 15 15 14 13 4 16 11 11 11 11 1 9 13 4 4 2
20 11 11 1 13 16 3 15 9 13 1 1 15 1 11 1 9 14 13 4 2
19 16 15 11 1 9 13 1 9 13 14 4 16 11 15 9 9 1 13 2
42 16 2 9 14 1 0 9 9 11 11 1 11 1 12 9 1 1 13 4 9 1 1 1 15 13 16 2 15 10 9 1 9 13 2 15 13 15 9 1 1 13 2
26 15 13 16 15 11 9 11 11 11 1 9 1 9 13 4 7 15 13 4 16 15 15 1 9 13 2
26 16 2 11 1 13 16 0 10 9 1 13 9 1 1 11 7 11 1 9 1 15 9 14 13 4 2
28 15 13 16 11 11 1 11 9 1 9 2 3 1 9 1 12 9 1 0 9 1 9 9 1 9 13 4 2
51 11 1 0 9 2 9 2 9 1 1 1 11 1 11 11 11 11 1 13 16 16 11 1 11 1 2 9 2 9 2 1 9 13 4 4 2 7 9 9 15 14 15 13 4 7 15 9 1 9 13 2
21 15 13 16 15 9 1 9 13 16 11 11 1 11 1 9 1 9 13 4 4 2
12 15 13 16 2 11 11 1 9 13 4 4 2
22 11 1 11 11 11 10 9 1 1 3 0 9 13 2 7 15 3 0 13 4 4 2
15 11 9 1 13 16 11 1 11 1 9 1 9 13 4 2
30 11 1 9 2 9 1 9 13 4 11 1 13 16 15 9 9 1 0 3 0 9 9 9 1 0 9 9 1 13 2
22 11 1 9 13 16 11 11 1 9 1 1 11 15 15 1 9 1 9 13 4 4 2
21 11 1 0 9 1 9 1 9 0 13 14 0 9 1 11 1 15 1 9 13 2
16 7 15 1 11 1 9 15 1 0 9 1 0 14 13 4 2
57 11 11 1 11 1 13 9 1 10 14 9 13 7 10 9 1 13 1 11 11 1 12 0 9 1 13 4 16 15 15 9 1 9 1 9 1 0 13 4 4 15 11 11 1 9 11 11 1 9 11 11 1 9 1 9 13 2
20 11 1 0 11 11 11 11 11 1 12 12 0 9 1 9 1 9 13 4 2
39 11 1 13 16 15 15 9 14 13 16 12 0 0 9 1 10 0 9 1 9 15 1 13 7 15 15 9 9 11 11 1 9 13 1 10 3 13 4 2
23 2 11 11 11 2 1 13 4 9 1 11 1 13 16 16 15 9 1 14 10 9 13 2
24 7 15 3 14 0 13 2 15 9 13 16 11 1 9 15 9 1 1 9 1 13 4 4 2
7 15 15 15 1 0 13 2
42 10 9 1 1 11 11 1 10 9 1 9 1 9 1 10 9 1 11 11 7 15 9 1 11 1 13 16 15 11 11 1 9 1 9 1 9 13 4 9 1 13 2
30 16 11 7 15 9 1 13 13 16 9 1 10 9 1 9 13 4 4 2 15 11 11 9 1 0 13 9 13 4 2
11 11 1 9 1 13 16 15 0 13 4 2
9 16 15 10 9 1 0 9 13 2
24 16 2 11 1 9 0 13 1 3 11 11 11 7 15 9 1 10 9 1 9 1 1 13 2
30 11 1 13 16 15 9 1 10 9 1 9 13 2 15 13 4 4 16 11 11 1 9 1 11 1 9 0 14 13 2
13 15 1 10 9 1 10 0 9 10 9 1 13 2
27 11 1 10 9 0 11 1 13 4 4 2 10 9 11 1 11 11 11 11 7 11 9 1 9 13 4 2
25 11 1 13 4 4 16 3 11 1 15 9 1 9 1 9 15 9 1 9 13 1 1 13 4 2
14 11 1 13 2 9 9 1 15 15 15 9 14 13 2
30 11 1 9 11 11 1 13 16 10 9 1 9 1 14 9 3 14 13 2 16 11 1 0 0 9 1 9 13 4 2
20 7 15 15 9 1 9 1 9 14 13 4 2 16 15 15 9 14 14 13 2
6 10 13 11 13 4 2
44 16 15 10 9 1 9 13 16 11 2 11 2 1 9 1 1 1 3 14 13 7 11 10 9 1 0 13 16 11 1 11 1 9 8 13 1 1 15 9 1 9 14 13 2
15 15 11 11 11 1 9 1 13 1 15 9 14 14 13 2
34 11 1 13 16 9 1 1 15 1 15 13 14 14 16 9 1 10 9 1 15 1 9 13 1 9 13 7 15 1 9 14 13 4 2
9 10 9 1 15 9 14 14 13 2
15 11 11 11 1 9 9 1 0 9 1 0 9 13 4 2
18 11 11 11 1 9 1 15 2 11 11 11 2 13 1 9 13 4 2
42 10 9 1 11 11 11 1 1 9 2 9 13 9 1 9 14 14 13 7 2 15 10 9 1 11 11 1 1 2 9 12 9 1 9 1 9 1 0 13 4 4 2
23 11 11 11 11 11 1 15 0 9 9 1 0 9 1 1 0 9 13 1 9 13 4 2
23 15 13 13 16 0 9 7 9 1 13 1 9 1 9 1 1 9 1 15 9 14 13 2
21 0 9 9 1 9 1 10 9 9 9 2 11 11 11 2 1 1 14 13 4 2
22 9 1 12 9 0 13 15 9 13 0 9 1 0 9 7 0 9 1 9 13 4 2
8 15 9 1 0 9 13 4 2
16 16 2 9 1 1 15 15 9 1 9 1 9 14 13 4 2
18 11 1 13 13 16 9 9 1 9 1 9 1 14 0 9 13 4 2
15 11 11 11 1 9 1 0 9 1 9 1 9 13 4 2
25 0 7 0 9 1 9 1 1 13 4 1 11 11 11 11 1 0 9 1 15 9 9 13 4 2
22 11 11 1 13 11 1 9 9 7 11 1 11 1 9 13 4 15 0 11 13 4 2
23 11 7 0 11 1 9 9 0 13 1 0 9 11 11 11 1 9 1 0 9 13 4 2
28 15 13 13 11 1 2 15 11 11 7 0 9 9 1 9 9 13 1 11 11 1 9 1 9 13 4 4 2
50 11 1 0 9 9 1 9 1 9 1 13 4 1 13 4 11 9 1 9 1 9 1 13 4 16 11 1 9 9 9 1 9 13 1 1 11 1 12 9 1 14 10 9 1 0 9 1 9 13 2
12 10 3 15 11 2 11 11 7 11 11 13 2
43 9 1 13 13 16 11 7 11 11 11 11 2 11 2 1 9 2 9 1 13 13 16 11 1 11 11 2 11 7 11 2 11 11 7 11 1 0 9 1 14 9 13 2
41 9 1 1 11 1 10 9 1 9 15 1 0 14 13 2 7 0 9 1 13 13 16 11 11 7 11 9 9 1 9 1 13 7 10 0 9 0 11 0 13 2
26 11 1 1 9 1 9 13 4 16 11 1 9 1 11 7 0 11 1 9 13 1 0 9 13 4 2
35 9 1 1 11 1 1 1 9 9 1 10 9 1 0 13 1 9 13 1 1 11 7 11 1 11 1 3 9 13 1 9 14 13 4 2
48 9 1 9 1 9 13 4 13 16 0 9 11 1 11 11 1 12 9 1 1 11 11 11 1 0 11 11 11 1 13 4 16 15 13 13 16 11 1 15 10 0 9 1 9 14 13 4 2
26 11 1 15 1 9 13 4 2 7 15 14 0 9 1 11 1 9 1 9 13 1 9 13 4 4 2
39 11 1 9 9 11 11 11 1 11 1 13 16 11 9 7 0 11 11 11 11 1 11 11 1 9 1 1 13 4 11 9 9 1 9 0 14 13 4 2
29 11 1 15 12 9 9 1 13 16 11 1 9 9 1 13 4 0 9 1 13 4 9 1 9 13 4 4 4 2
13 15 13 16 15 11 1 9 1 0 9 14 13 2
21 11 1 1 10 9 1 9 9 11 11 11 7 9 9 11 11 11 14 0 13 2
31 11 1 11 1 15 9 0 13 1 9 9 1 9 1 0 9 13 4 7 9 1 9 1 9 0 13 1 9 13 4 2
29 0 9 1 13 13 16 11 11 1 0 11 11 1 0 9 1 9 1 0 11 1 9 1 9 1 9 13 4 2
17 0 9 1 10 11 1 1 9 1 9 1 9 1 0 9 13 2
28 11 11 1 9 1 9 1 0 11 1 0 13 1 9 1 9 1 11 11 1 9 11 11 0 9 13 4 2
21 3 11 11 1 14 9 1 15 9 14 13 16 10 11 1 9 1 0 9 13 2
13 15 13 16 9 1 9 1 10 11 10 0 13 2
16 11 1 10 9 13 7 11 1 9 1 9 9 1 13 4 2
22 0 9 1 13 13 16 10 11 1 9 1 0 9 1 9 1 9 1 9 13 4 2
13 0 9 1 10 11 1 1 9 1 0 9 13 2
16 11 1 11 1 1 15 9 1 0 13 1 15 9 14 13 2
19 9 11 1 9 11 11 1 13 16 15 9 1 11 1 0 9 13 4 2
16 15 13 16 11 11 1 9 1 14 12 12 9 1 9 13 2
18 9 9 7 9 1 9 1 13 4 10 9 1 3 2 3 9 13 2
10 15 9 1 0 9 13 1 9 13 2
11 15 9 1 15 9 14 0 13 4 4 2
12 15 9 1 10 9 1 10 10 9 9 13 2
40 9 1 13 13 16 10 11 1 1 9 1 11 1 9 13 1 9 13 9 1 10 9 13 16 15 0 9 1 13 11 7 15 0 9 1 9 14 13 4 2
7 15 9 1 9 13 4 2
33 0 11 11 11 1 11 9 1 1 0 0 0 9 11 11 1 13 4 16 0 7 0 15 2 15 1 0 9 1 9 13 4 2
15 15 15 14 13 16 15 11 1 9 9 13 4 4 4 2
37 3 14 11 11 1 11 11 1 12 0 9 1 9 9 13 2 7 15 11 1 0 0 9 1 1 1 10 0 2 0 7 0 9 14 9 13 2
12 11 11 11 1 11 1 9 1 13 4 4 2
22 15 12 2 0 11 9 1 1 15 0 9 1 9 9 7 0 0 9 1 9 13 2
14 15 11 11 1 2 0 0 9 2 1 14 9 13 2
9 15 15 9 1 9 9 9 13 2
37 12 0 10 0 0 9 1 15 14 13 16 15 11 1 9 1 9 14 13 4 4 16 15 14 0 9 1 9 1 14 11 9 1 9 13 4 2
19 11 11 1 13 16 15 0 9 1 0 7 0 9 13 1 9 1 13 2
13 15 0 13 4 13 4 16 15 9 0 14 13 2
17 15 0 9 1 1 14 0 9 1 9 13 4 1 9 1 13 2
20 15 13 16 11 11 1 0 9 13 10 9 1 9 1 9 0 13 4 4 2
17 11 11 1 11 7 11 1 9 1 13 4 9 1 14 9 13 2
12 15 13 16 11 7 11 0 9 1 9 13 2
15 10 12 9 1 1 9 1 9 1 12 9 1 9 13 2
23 15 15 11 11 1 12 9 9 1 9 13 9 11 11 11 1 9 1 0 9 0 13 2
