14187 11
29 3 15 15 13 1 10 9 0 1 13 10 9 16 15 13 9 1 10 9 7 10 9 16 13 9 1 10 9 2
59 9 1 10 9 1 10 9 7 10 9 0 10 9 0 13 1 12 12 1 10 9 0 2 13 1 10 9 12 16 4 1 13 13 1 12 1 12 12 1 10 9 12 2 7 1 10 9 0 4 1 13 15 1 3 12 1 12 9 2
89 11 2 12 2 11 11 2 10 9 0 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 7 11 11 4 13 13 10 9 16 13 10 0 9 1 10 11 11 1 13 1 10 9 1 10 11 11 11 1 11 2 11 2 3 1 3 1 12 9 1 9 1 10 11 11 1 11 2 8 2 1 10 9 1 10 9 1 9 1 10 9 2 11 11 2
20 10 9 1 9 13 12 9 3 0 1 13 9 0 7 15 16 3 13 9 2
13 13 1 10 10 9 11 7 11 11 10 0 9 2
12 13 10 9 13 1 9 10 9 13 15 0 2
33 7 13 3 0 16 10 9 13 10 9 1 11 11 15 3 15 13 1 11 2 16 13 9 1 10 0 9 7 9 1 10 9 2
23 13 16 13 0 16 10 9 13 9 7 3 15 13 1 10 9 0 1 9 2 2 13 2
19 10 0 9 13 10 9 1 9 2 16 3 13 10 9 1 10 9 0 2
17 13 1 9 1 10 11 11 7 11 11 2 1 11 11 1 11 2
69 10 9 0 1 10 9 1 9 13 10 9 1 9 1 9 7 13 1 10 2 9 1 9 2 16 13 10 9 16 13 1 10 9 7 1 10 9 1 10 9 2 7 10 9 9 2 7 11 11 2 16 13 10 9 1 10 9 16 15 13 1 10 9 1 10 9 1 9 2
30 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 11 11 11 1 10 9 0 1 11 2
29 10 9 1 11 11 2 3 11 11 11 11 11 2 13 10 9 0 0 2 13 1 10 9 1 11 11 2 11 2
18 13 10 13 9 1 13 10 9 2 7 16 13 13 15 3 13 15 2
10 11 11 13 10 0 9 1 10 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
28 11 11 11 13 1 10 9 1 12 9 7 1 10 9 1 11 11 2 1 10 9 1 9 11 2 12 2 2
12 4 13 1 10 9 1 11 1 9 3 13 2
49 4 1 13 1 10 9 10 9 1 11 11 7 13 10 9 1 10 8 3 9 3 3 13 16 3 13 10 9 1 10 9 2 16 15 13 3 10 9 0 16 11 13 1 13 15 1 10 9 2
28 3 13 9 1 13 7 13 1 10 9 1 10 9 1 10 9 13 1 11 1 10 9 0 7 10 9 0 2
4 13 12 9 2
43 10 11 13 10 9 1 10 9 1 10 0 9 7 15 13 1 10 9 16 15 13 11 7 13 3 1 10 9 0 3 13 10 11 12 1 13 0 9 0 1 10 9 2
28 10 9 13 16 10 2 9 2 16 15 4 13 1 13 1 10 9 11 1 10 9 4 13 15 1 10 9 2
21 15 1 10 13 15 1 16 15 4 13 0 2 9 1 11 2 13 1 13 3 2
16 10 9 1 10 12 9 1 11 13 10 0 9 1 10 9 2
27 15 1 10 0 9 1 10 9 13 1 10 9 1 11 1 10 12 9 7 3 10 9 3 13 1 9 2
12 13 9 0 2 0 7 10 9 13 3 0 2
29 1 10 9 1 10 9 11 2 1 9 0 10 9 1 11 2 13 10 9 1 10 11 7 9 1 10 9 11 2
10 11 11 2 9 1 9 0 11 2 2
65 10 9 1 10 0 9 1 10 9 13 13 10 9 0 1 13 10 9 3 3 1 15 2 1 10 11 11 1 10 9 7 10 9 1 11 11 11 11 1 11 2 11 2 13 12 9 1 9 0 1 12 9 13 15 15 3 1 15 1 10 9 0 1 9 2
45 10 9 13 10 9 1 9 7 1 9 1 12 12 12 9 2 15 16 13 4 1 13 10 12 9 1 9 2 3 1 9 1 10 9 1 9 3 0 7 15 13 1 10 9 2
28 1 9 1 11 12 2 13 10 9 7 9 1 10 9 0 1 10 9 11 2 0 1 10 9 1 10 11 2
8 11 1 11 2 10 11 2 2
45 11 13 16 1 9 0 13 12 9 3 9 2 15 2 4 13 16 16 13 1 9 10 11 2 3 2 15 13 10 9 2 16 15 13 15 16 13 1 10 9 0 2 2 13 2
36 1 12 2 10 9 4 13 2 13 1 11 11 1 10 9 1 9 0 1 11 2 16 13 1 12 1 12 9 1 10 9 1 13 1 12 2
66 11 11 2 13 10 12 1 11 1 12 1 11 2 11 13 10 9 2 9 7 9 1 10 9 1 11 11 11 2 3 13 1 10 9 1 13 9 15 13 1 11 10 15 13 0 9 0 1 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2
43 1 9 2 10 9 1 0 9 1 9 13 3 1 10 12 12 9 13 11 2 12 2 2 10 11 2 12 2 7 10 11 11 2 12 2 2 3 1 11 2 12 2 2
65 3 7 2 11 13 10 11 1 10 9 1 11 2 11 15 2 8 2 2 3 13 2 10 9 1 10 9 1 10 9 1 10 11 11 1 11 2 11 11 2 1 10 9 1 10 9 1 9 2 11 11 2 15 15 13 10 9 1 13 1 10 9 1 11 2
44 10 16 10 9 13 10 0 9 0 1 10 9 2 15 13 1 10 9 0 7 1 10 9 1 9 7 9 1 10 0 9 0 2 1 10 15 3 13 10 0 9 1 9 2
31 1 3 2 11 4 13 1 10 10 9 1 9 3 1 13 1 10 9 13 10 9 1 10 11 2 11 11 11 11 2 2
13 10 9 1 9 13 1 12 8 2 5 9 5 2
77 11 11 15 4 13 1 10 9 0 1 10 9 7 1 15 4 13 1 10 9 1 10 9 1 0 9 1 10 9 0 7 9 1 10 15 15 13 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 1 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2 1 13 10 9 2
13 15 15 13 7 3 13 15 16 13 1 3 3 2
20 3 2 7 16 10 9 1 9 13 10 9 1 9 2 13 3 15 1 9 2
14 10 0 9 7 15 13 7 15 13 10 9 1 13 2
27 15 13 1 10 9 2 15 13 10 9 0 1 11 7 3 13 15 1 9 1 16 10 9 13 1 0 2
20 11 11 13 1 9 1 10 11 1 10 9 13 1 10 0 9 0 11 11 2
50 15 1 10 0 9 13 10 9 1 10 11 2 11 11 2 2 12 2 2 10 9 1 11 11 2 12 2 2 7 10 9 0 1 11 11 10 11 2 12 2 7 1 10 9 1 11 2 12 2 2
16 13 15 1 10 9 3 0 13 1 10 11 12 1 10 9 2
22 1 10 9 13 1 10 11 11 11 2 9 1 10 9 1 10 11 1 11 7 11 2
32 11 13 11 1 10 11 13 10 0 9 1 10 9 0 11 2 16 13 10 9 1 10 9 12 2 1 10 9 0 11 11 2
21 1 10 9 15 13 9 1 11 11 2 11 11 2 11 11 2 11 11 7 11 2
23 10 9 0 11 11 4 13 1 10 9 1 10 9 0 0 1 10 9 1 9 7 9 2
16 10 9 1 10 9 0 13 10 9 0 0 7 10 9 0 2
40 1 13 10 9 0 2 0 7 16 10 9 0 15 13 1 13 1 10 9 2 3 4 13 2 9 2 2 16 7 10 9 7 10 9 13 0 1 10 9 2
16 13 10 9 0 7 0 15 13 15 2 7 15 4 13 15 2
11 10 9 13 10 9 1 10 9 1 9 2
42 1 13 9 15 13 9 1 9 0 2 16 10 9 3 4 13 15 1 10 9 0 0 2 7 1 10 9 1 10 9 1 9 0 1 10 9 0 7 10 9 0 2
30 10 9 1 10 9 13 1 3 12 9 16 4 4 13 1 10 9 0 7 3 12 9 16 15 13 1 10 9 0 2
12 11 13 10 9 3 1 11 11 11 11 12 2
14 15 13 10 9 1 10 0 9 1 10 11 1 11 2
32 10 11 11 11 13 10 11 16 10 9 13 3 3 9 15 3 0 1 10 9 0 7 0 9 1 10 9 1 9 7 9 2
33 1 3 0 9 7 1 9 0 2 15 13 16 10 9 13 1 10 9 1 10 9 7 1 10 9 1 10 9 0 1 10 9 2
34 10 11 0 2 11 11 13 13 15 1 10 9 0 1 13 10 9 1 10 9 1 10 9 1 9 1 11 11 1 10 9 16 13 2
26 3 13 9 1 9 7 10 9 0 16 4 13 10 9 1 2 9 16 13 10 9 7 9 0 2 2
27 10 9 1 10 0 11 11 1 11 11 13 10 9 1 10 9 1 9 2 9 2 9 1 9 7 9 2
23 10 9 13 10 9 1 10 9 11 11 15 13 10 9 0 1 10 9 13 1 9 0 2
18 2 16 15 13 1 9 2 15 3 13 10 9 0 2 2 4 13 2
18 11 3 13 11 11 7 10 9 1 10 9 1 9 7 1 0 9 2
22 10 9 13 3 1 10 12 9 1 3 2 16 13 13 1 10 9 16 4 1 13 2
28 10 9 1 10 0 9 16 13 10 9 1 10 9 2 1 12 9 7 0 1 9 2 4 4 13 1 9 2
55 3 3 2 16 13 10 9 1 15 1 10 9 2 1 10 12 9 2 9 8 2 13 16 13 10 0 9 2 1 15 16 15 13 16 1 10 9 1 10 9 13 10 9 0 1 1 10 12 9 5 5 8 1 9 2
28 1 12 2 11 13 11 7 10 9 1 9 0 1 11 2 13 9 1 0 9 1 10 9 1 10 1 9 2
44 1 9 2 11 7 11 2 3 7 10 10 9 2 4 13 9 1 10 0 9 2 7 7 11 15 13 7 13 10 0 9 2 13 15 1 15 1 10 9 1 11 1 15 2
48 9 1 9 1 10 9 1 10 9 13 11 11 7 11 11 2 0 1 10 9 1 10 9 1 10 9 11 11 11 1 10 9 11 11 2 15 3 13 1 10 9 1 10 9 1 9 2 2
69 1 10 9 3 13 11 11 15 13 10 0 9 2 15 9 1 13 1 11 1 10 9 2 11 15 13 9 1 16 10 13 3 7 13 3 13 10 9 2 10 9 1 11 13 1 10 9 7 15 13 1 10 9 16 11 13 8 2 10 15 15 13 7 15 13 1 10 9 2
26 10 9 4 3 13 1 9 1 11 11 10 12 1 11 2 7 3 1 11 10 12 1 11 1 12 2
10 13 10 0 9 1 10 9 0 11 2
16 3 13 9 0 7 3 0 2 1 10 9 1 10 15 13 2
19 13 13 16 10 9 3 13 1 9 1 9 0 2 7 13 1 9 0 2
15 11 15 13 0 1 10 9 15 4 13 1 9 7 9 2
9 10 9 0 13 15 15 11 13 2
54 1 13 1 10 9 1 11 2 10 10 9 16 13 1 10 9 2 13 9 7 13 1 10 2 8 8 2 13 13 10 9 1 13 10 9 1 9 7 9 1 12 9 1 15 1 10 9 1 11 1 11 7 11 2
68 15 4 13 10 9 1 10 10 9 2 13 1 10 9 1 5 16 13 9 1 3 4 1 13 10 9 7 15 1 10 9 13 10 9 7 8 3 4 13 13 15 2 13 1 9 7 3 13 7 3 13 10 9 3 0 16 15 13 1 10 9 2 10 12 1 10 9 8
9 10 9 13 0 7 3 3 0 2
50 11 11 13 10 9 13 1 10 11 11 11 1 11 1 10 11 1 11 11 2 7 13 1 11 11 11 1 10 9 2 11 11 11 1 10 9 2 11 11 11 1 10 9 2 7 11 1 10 9 2
31 11 15 13 1 10 9 1 9 0 1 10 11 2 13 1 11 2 11 7 11 2 1 9 1 3 13 1 9 10 9 2
15 4 13 1 0 9 1 10 9 1 10 9 11 1 12 2
22 13 1 10 9 1 10 9 9 1 9 1 9 1 13 3 16 15 13 1 10 9 2
40 1 3 1 11 11 2 16 13 10 9 3 0 1 10 9 1 9 0 2 10 9 3 0 1 10 9 1 10 9 13 2 11 12 2 12 2 12 7 12 2
29 10 2 11 2 13 10 9 9 16 13 12 0 9 2 15 15 13 16 3 1 10 9 3 13 10 9 1 9 2
11 11 11 1 11 7 11 11 1 11 11 2
9 11 10 11 15 13 12 9 3 2
53 13 1 10 9 1 15 15 13 10 0 9 1 10 9 2 3 7 13 1 9 1 11 11 1 10 11 11 1 10 11 1 11 1 10 11 1 12 7 13 3 1 0 9 0 1 11 11 2 11 7 10 11 2
8 9 1 10 11 11 1 11 2
33 10 9 11 2 13 3 1 10 9 11 11 2 13 0 1 10 9 1 11 2 11 2 10 9 0 1 10 0 9 0 7 0 2
43 10 11 1 11 13 1 10 9 15 1 10 9 0 3 0 1 10 9 1 11 2 16 10 9 0 4 13 15 1 10 9 1 10 9 0 13 1 9 1 10 9 12 2
33 10 9 2 13 1 10 0 9 1 12 9 7 9 1 10 9 0 1 11 2 13 15 16 13 10 0 9 1 9 7 9 0 2
19 3 1 3 12 9 1 10 8 8 2 10 9 4 13 1 10 8 8 2
11 10 9 1 11 15 13 13 1 10 9 2
13 10 9 0 13 1 15 1 10 9 12 1 12 2
31 16 13 1 9 0 2 11 2 11 13 10 9 1 10 9 0 0 1 10 9 7 3 3 2 1 10 9 1 10 9 2
20 10 9 1 10 9 0 13 0 1 9 0 1 9 0 1 9 1 10 9 2
22 10 9 16 10 9 13 0 9 2 13 0 16 15 13 1 11 1 13 1 10 9 2
37 10 9 1 0 9 7 9 15 13 1 9 7 9 1 10 9 2 1 10 12 9 2 9 0 2 2 16 10 9 0 15 13 1 10 9 0 2
50 1 10 9 10 9 1 12 9 0 4 13 13 15 1 10 9 1 10 9 1 16 4 13 1 10 9 12 2 15 0 1 10 9 2 13 10 11 11 10 16 3 9 1 0 9 13 1 10 9 2
34 10 9 0 4 13 3 10 9 0 2 9 1 10 9 4 13 10 9 1 10 9 7 10 9 1 9 15 15 13 10 9 0 2 2
16 1 12 11 4 13 9 1 10 9 2 10 11 11 1 11 2
27 13 1 10 9 2 9 7 9 1 9 0 2 10 9 13 1 10 9 13 3 10 9 1 10 9 0 2
15 13 10 8 1 9 1 0 9 2 7 3 1 9 0 2
24 15 1 10 9 15 13 1 9 1 10 9 3 0 3 2 1 11 2 11 11 2 7 11 2
14 10 9 13 9 1 10 9 0 0 2 9 7 0 2
25 11 13 10 9 0 1 9 7 4 13 1 10 9 1 11 1 9 7 9 15 11 13 1 11 2
28 10 9 0 10 11 4 13 10 0 2 10 11 11 11 11 11 2 1 10 9 1 10 9 7 9 9 11 2
36 7 3 15 13 1 10 9 7 1 9 10 9 1 11 11 2 1 10 9 1 11 2 13 10 11 7 16 15 1 11 11 7 11 10 11 2
28 10 9 0 0 1 10 9 1 9 1 10 9 15 13 1 10 0 9 1 0 9 1 10 16 13 10 9 2
41 4 13 1 12 9 0 1 0 9 2 10 9 0 13 1 9 0 16 13 10 9 7 9 1 10 9 2 1 10 9 0 1 10 9 13 10 9 1 10 9 2
14 13 9 1 10 11 1 11 2 1 10 9 1 9 2
31 9 1 9 13 16 3 13 9 0 7 9 0 15 16 13 1 9 1 10 9 0 0 13 1 11 11 1 11 7 11 2
23 3 2 10 9 13 10 9 7 10 9 13 1 10 9 2 1 10 9 1 10 12 9 2
32 13 1 9 10 9 1 10 9 0 2 4 15 13 15 1 10 9 0 1 10 9 1 10 9 2 2 13 10 9 3 0 2
34 2 11 11 2 13 1 10 12 9 8 10 0 9 1 10 0 9 1 9 2 10 2 11 2 3 13 1 10 9 1 10 0 9 2
24 1 10 9 1 10 9 2 10 9 13 10 9 0 1 2 1 10 15 13 9 7 13 9 2
36 3 1 10 9 2 11 3 13 10 9 1 9 1 11 1 10 9 1 12 2 7 10 9 1 11 12 2 12 2 7 12 4 13 1 12 2
35 1 13 10 9 1 0 9 2 7 1 10 0 9 1 10 9 1 9 2 16 13 0 2 10 9 13 10 9 1 10 0 9 1 9 2
7 3 15 13 10 9 2 2
36 1 9 9 2 9 2 10 9 13 1 10 9 1 11 11 2 13 1 9 1 10 9 1 11 7 11 2 11 7 11 11 7 11 7 11 2
37 10 9 13 13 16 15 13 11 2 13 10 0 9 2 3 4 7 13 3 13 1 10 9 2 3 13 9 1 10 9 1 13 9 1 10 9 2
19 15 13 1 15 1 10 9 16 13 1 10 9 2 16 13 10 9 0 2
25 13 3 9 1 9 0 2 3 9 2 7 13 10 0 9 0 1 12 1 10 11 11 1 11 2
46 1 10 9 13 10 9 1 9 7 9 7 12 9 1 9 1 9 2 3 1 9 0 1 9 2 3 10 9 7 9 1 10 0 8 1 10 0 9 13 1 9 0 13 1 9 2
40 1 10 9 1 0 10 9 1 10 9 4 13 15 1 10 9 1 13 7 13 10 9 1 10 9 0 2 1 10 9 1 10 9 7 10 9 2 9 2 2
21 11 13 10 9 1 11 3 16 0 9 1 10 9 13 10 9 0 7 10 9 2
47 4 13 12 9 2 7 16 3 13 10 9 3 1 10 9 7 1 10 9 2 15 13 0 13 10 9 2 3 10 9 2 9 1 9 2 7 15 13 1 10 9 0 1 9 7 0 2
42 13 10 0 9 1 10 11 11 10 12 1 11 1 10 12 2 1 10 9 1 10 9 1 9 12 1 11 10 11 10 15 13 8 1 9 1 10 2 9 0 2 2
25 10 11 13 10 9 1 16 10 0 9 13 10 0 9 2 1 15 15 10 9 1 2 13 2 2
24 10 9 1 9 13 1 13 10 10 0 9 1 10 9 1 8 8 1 11 1 10 9 12 2
13 1 12 13 1 10 9 11 2 11 1 10 11 2
8 11 15 13 11 1 10 9 2
28 10 9 1 10 11 13 10 9 0 0 12 1 9 1 11 11 11 1 11 2 9 1 10 8 9 1 11 2
14 13 1 9 0 1 16 10 9 15 13 3 1 12 2
38 13 10 9 1 10 9 1 10 9 3 0 1 10 9 0 1 11 1 10 9 11 11 1 10 9 11 11 7 10 9 1 9 1 9 11 11 11 2
37 10 9 11 2 10 9 16 13 1 10 8 7 15 13 0 2 15 4 13 1 10 9 7 4 13 1 10 9 1 10 9 1 10 9 1 9 2
13 3 10 10 9 15 13 3 1 3 1 13 9 2
20 10 9 0 3 13 9 1 10 11 11 7 4 13 3 3 1 10 11 12 2
40 10 9 1 9 7 9 13 10 9 0 7 0 16 15 13 1 12 9 2 1 10 15 15 13 1 13 1 10 9 1 10 9 2 11 7 11 2 12 2 2
18 1 10 9 1 10 9 11 13 1 13 10 11 11 1 10 0 9 2
14 3 2 4 13 3 1 10 11 1 11 2 11 2 2
30 15 13 12 5 1 10 9 1 9 2 15 4 13 12 3 1 10 9 1 8 2 13 2 16 10 9 13 10 8 2
49 3 11 1 12 15 13 1 9 0 2 3 10 9 4 1 13 15 11 1 11 1 12 2 3 11 1 11 1 12 2 7 11 1 11 1 12 1 10 11 1 11 11 1 11 11 13 1 12 2
31 1 13 10 9 0 2 13 1 10 9 3 1 15 1 13 15 1 10 9 1 10 9 1 10 9 7 13 15 12 9 2
7 1 12 13 9 1 11 2
15 10 9 4 13 1 9 2 9 1 9 7 9 1 9 2
57 12 9 3 13 1 10 9 1 10 9 1 11 2 1 10 9 1 10 11 11 11 11 2 8 9 1 10 9 1 10 9 0 2 1 10 9 1 11 1 10 11 11 1 10 12 1 11 1 12 7 10 12 1 11 1 12 2
24 10 9 1 9 1 9 1 9 13 10 9 0 2 13 1 10 9 0 7 10 9 1 11 2
9 3 1 9 16 4 13 9 0 2
11 10 9 1 10 11 11 11 13 10 9 2
64 13 1 9 2 11 11 13 12 9 1 2 11 1 10 11 2 1 10 9 11 11 2 15 1 9 1 12 1 10 9 2 11 1 10 11 2 7 15 1 10 9 0 0 11 11 2 1 10 15 13 10 9 1 11 7 1 10 15 15 13 10 0 9 2
22 10 9 13 9 1 10 9 0 0 0 11 1 8 2 16 15 13 1 10 9 0 2
11 1 9 2 13 10 0 9 1 10 9 2
10 15 13 1 10 0 9 1 10 9 2
48 11 11 11 2 2 11 2 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 10 9 0 0 2 9 1 10 9 0 11 2 0 1 11 11 2 11 11 7 11 11 11 2 2
31 1 10 9 0 13 10 10 9 1 10 9 2 16 1 12 10 11 11 8 13 10 9 1 13 1 12 1 10 9 0 2
37 11 11 1 11 13 10 9 0 1 10 9 1 11 2 0 1 10 9 1 11 1 11 2 1 10 9 1 10 11 11 0 1 10 9 1 11 2
30 1 10 9 15 13 10 9 1 10 9 12 16 13 1 10 9 11 11 13 1 10 11 2 9 1 11 7 11 11 2
31 10 9 13 1 10 9 1 9 15 1 11 11 1 1 11 11 1 13 15 15 4 13 1 10 9 1 9 1 11 11 2
42 1 10 11 1 10 11 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
39 1 10 12 5 9 0 1 9 1 11 10 0 9 11 11 13 10 9 0 1 10 9 11 2 15 13 10 9 0 1 10 0 9 1 10 0 9 11 2
45 3 10 3 0 1 15 13 10 11 2 13 1 10 9 0 1 12 2 10 9 13 0 1 13 12 9 2 1 12 1 0 2 1 10 9 1 10 9 0 1 9 7 9 0 2
18 11 11 13 9 1 11 7 11 2 12 9 16 13 1 10 9 0 2
22 13 10 9 12 2 7 11 7 11 13 1 10 0 9 1 10 9 1 9 2 9 2
16 10 9 13 10 9 3 1 16 10 9 4 13 1 10 9 2
104 10 9 2 11 2 11 11 11 11 11 2 2 13 10 9 1 16 15 2 9 2 3 13 15 9 15 10 9 0 13 1 10 9 7 1 16 15 0 4 4 13 1 9 1 10 9 1 10 9 7 1 9 1 9 0 2 10 9 0 13 0 1 16 10 9 0 1 11 15 13 7 13 1 15 16 13 1 10 9 1 10 9 0 2 2 11 2 9 2 8 9 0 2 2 2 15 15 13 1 11 1 10 9 2
24 13 3 13 1 11 1 10 9 1 12 9 2 1 16 10 9 0 13 16 13 9 1 11 2
19 1 10 9 2 10 9 0 11 13 9 2 9 2 9 2 9 2 9 2
27 1 12 13 10 9 11 11 11 2 11 11 2 15 16 13 1 11 11 2 11 11 13 10 9 1 11 2
16 10 9 13 1 10 9 1 10 11 11 7 13 10 9 0 2
26 15 13 16 1 0 9 15 13 1 10 9 1 11 1 10 11 1 11 11 2 1 3 10 9 9 2
38 13 1 10 9 0 1 11 2 15 13 1 10 12 9 1 9 1 11 1 10 9 7 13 1 10 9 0 1 11 2 11 2 1 10 9 1 11 2
29 10 9 1 10 9 3 13 0 1 10 9 1 10 9 2 3 16 15 13 10 0 9 1 10 9 1 10 9 2
14 1 12 13 1 9 1 10 9 0 10 11 11 11 2
8 10 9 1 10 9 13 0 2
8 13 9 1 9 0 7 0 2
22 1 12 15 13 1 11 7 15 13 1 9 0 1 10 11 11 1 11 2 1 11 2
22 11 13 10 9 7 9 0 2 13 1 10 9 1 11 11 2 1 10 9 1 11 2
34 2 11 2 4 13 1 12 9 1 10 11 11 2 12 9 1 9 1 12 9 2 10 9 0 1 12 2 7 12 9 1 12 2 2
35 3 1 10 9 3 0 2 7 3 0 2 1 10 9 0 2 11 11 15 13 3 1 10 12 1 10 9 12 1 11 2 1 11 11 2
45 10 11 11 11 2 1 9 2 11 11 11 2 13 10 9 0 0 1 12 9 2 12 5 2 1 9 2 1 10 11 11 7 11 11 2 13 1 11 2 11 2 2 11 11 2
31 15 13 12 9 1 1 10 9 0 2 3 1 12 3 9 16 13 1 10 9 7 12 9 1 9 16 13 1 10 9 2
10 11 11 11 11 2 2 13 8 8 2
11 10 9 1 11 15 13 0 1 10 9 2
20 1 9 1 10 12 10 11 11 15 13 1 10 11 11 11 11 2 11 2 2
30 10 11 13 0 1 10 9 1 9 11 2 12 1 10 9 2 7 1 10 9 13 10 9 0 11 2 11 1 9 2
55 15 0 2 15 3 3 2 7 1 10 10 9 13 1 9 2 3 3 2 1 10 9 1 11 2 10 9 1 10 9 1 9 0 2 13 15 1 10 9 1 9 16 10 9 13 0 7 1 10 0 9 1 9 0 2
25 1 12 2 13 1 10 9 1 11 13 1 10 9 0 7 13 1 11 1 10 9 1 10 9 2
55 4 13 1 10 9 1 10 9 13 0 9 2 1 10 9 2 10 9 1 9 13 10 9 3 0 7 13 0 1 10 9 13 10 9 0 16 15 13 15 13 10 9 1 10 9 16 13 13 1 10 9 1 10 9 2
20 10 9 1 12 2 13 9 1 10 9 0 2 13 12 9 3 1 10 11 2
26 11 11 2 8 9 1 10 9 0 2 7 11 1 10 11 2 10 0 9 1 10 9 2 1 15 2
36 1 10 9 2 1 10 9 7 1 10 9 0 1 10 9 1 11 2 15 13 9 10 9 1 9 2 9 0 7 9 16 13 9 1 9 2
44 10 9 13 1 11 13 1 15 1 10 0 9 2 11 7 11 2 11 7 11 2 11 0 2 11 7 11 2 11 2 11 7 11 1 9 0 7 11 7 11 1 9 0 2
32 15 4 4 13 10 9 1 11 9 0 1 13 10 9 7 1 10 3 13 10 9 1 10 9 1 13 10 9 1 10 9 2
24 7 15 9 1 10 9 13 10 9 7 10 9 16 13 2 1 3 13 1 10 0 9 0 2
20 10 9 3 0 7 0 15 13 1 10 9 11 2 16 13 1 10 12 9 2
29 1 10 9 12 13 10 0 9 1 9 10 15 13 10 9 2 3 10 9 11 11 1 13 12 9 1 11 11 2
39 10 9 2 13 2 15 10 9 0 1 10 9 0 13 9 1 9 1 10 9 2 10 9 0 15 13 1 10 9 2 7 10 9 0 13 12 9 0 2
24 11 13 10 9 0 1 10 0 9 1 9 0 2 11 11 2 3 13 1 9 1 9 0 2
23 16 15 13 16 15 1 10 12 9 13 10 9 15 13 3 3 1 4 1 13 10 9 2
14 10 9 4 13 7 13 1 10 10 9 1 9 0 2
18 10 11 11 4 13 1 11 1 11 16 15 13 13 15 1 10 9 2
29 1 9 2 15 1 10 0 9 0 13 10 9 1 10 9 0 1 10 9 1 8 12 1 10 9 1 10 9 2
29 3 2 10 9 1 10 9 1 11 1 13 0 9 4 13 1 11 2 10 9 16 13 10 9 2 1 9 0 2
20 13 10 9 16 13 9 7 10 9 0 1 10 9 7 9 1 10 9 11 2
24 10 9 3 0 2 4 13 1 9 1 10 9 1 10 9 13 1 10 10 9 1 10 9 2
21 10 9 0 0 15 13 1 9 1 10 9 1 11 7 9 1 10 9 1 11 2
23 13 1 10 9 1 11 2 11 12 9 2 11 11 2 11 11 2 11 11 7 11 11 2
17 1 10 9 0 13 10 9 7 10 9 7 13 13 1 12 9 2
25 3 15 13 16 15 13 1 9 2 13 10 9 16 10 9 3 0 7 11 13 10 9 1 11 2
26 10 9 13 10 9 1 10 9 0 2 9 2 1 0 9 1 10 9 2 9 7 0 1 10 9 2
26 13 1 10 0 9 0 7 0 2 1 10 15 15 13 10 9 1 9 7 9 1 10 9 1 11 2
98 10 9 13 10 9 15 13 1 10 9 1 10 9 16 13 10 9 1 11 2 13 10 0 9 15 1 10 9 4 13 1 9 7 1 9 7 3 10 9 1 10 9 15 4 13 2 16 3 9 2 3 10 9 1 0 9 16 15 13 1 10 9 15 13 1 13 10 10 9 1 10 9 1 0 9 7 2 3 1 10 9 1 11 2 10 9 13 1 3 16 3 10 9 4 13 1 3 2
28 1 9 2 15 13 1 10 9 0 13 1 10 9 1 9 1 10 9 0 13 10 0 9 1 9 1 15 2
11 10 0 9 4 3 13 1 9 1 9 2
27 1 10 9 2 13 7 13 10 9 15 13 1 10 9 3 0 1 10 9 0 16 13 10 9 1 9 2
11 10 9 4 13 10 12 1 11 1 12 2
45 10 10 9 3 4 13 1 10 0 11 2 3 7 10 9 13 10 9 1 10 0 9 1 9 1 10 12 9 16 13 10 9 0 1 15 1 10 9 1 11 2 10 9 11 2
65 10 9 0 2 10 12 1 11 1 12 2 15 13 1 11 11 11 2 11 2 9 1 11 11 11 2 11 7 11 11 7 9 1 11 11 11 2 11 2 14 2 0 9 1 10 11 11 2 2 1 10 0 9 13 12 9 2 11 11 2 11 11 7 11 2
64 10 11 1 11 2 11 7 10 11 13 12 1 10 9 13 1 10 9 1 11 2 9 1 10 11 16 4 4 13 1 11 16 13 10 0 0 1 15 1 10 0 9 1 10 9 11 13 1 7 13 3 1 12 9 1 10 0 9 2 10 12 2 12 2
24 10 9 13 1 9 13 1 9 1 9 13 1 10 9 2 7 1 9 7 9 1 10 9 2
26 10 0 9 0 13 9 1 10 11 2 3 13 1 10 9 1 10 11 11 2 13 1 11 11 2 2
9 13 1 10 9 1 11 1 12 2
7 3 0 1 10 9 0 2
56 1 10 9 13 1 10 9 1 10 9 3 13 0 2 1 9 1 7 3 1 10 9 1 2 9 0 2 2 10 9 11 11 2 10 9 9 13 3 1 9 2 10 9 1 10 9 1 11 11 1 10 9 1 9 0 2
75 1 10 0 9 15 0 15 1 9 0 2 12 9 2 1 9 2 12 5 9 2 2 1 10 0 10 9 7 10 1 10 9 3 13 10 9 7 15 13 1 10 11 1 11 1 10 0 9 8 1 10 9 1 9 2 3 3 13 1 13 10 9 2 13 3 0 9 0 1 12 9 7 13 3 2
8 15 13 1 10 11 1 11 2
32 10 9 0 1 10 9 0 2 13 1 10 9 2 15 13 1 10 9 10 12 1 11 1 12 2 1 11 11 2 11 2 2
42 13 3 16 10 12 1 11 1 12 13 10 9 1 9 1 9 2 9 2 9 1 9 7 9 1 9 1 10 0 9 3 15 4 13 10 9 1 10 11 11 11 2
10 10 0 9 13 10 9 1 12 8 2
49 3 13 10 9 13 10 9 1 8 7 9 13 2 1 10 0 9 15 13 10 9 1 16 10 10 10 9 15 4 1 13 10 9 2 7 10 0 9 13 10 9 16 13 1 10 15 16 13 2
21 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 10 9 0 0 2
64 10 9 15 13 10 9 1 13 10 9 0 1 10 9 2 3 7 2 1 10 9 0 2 10 9 13 10 9 1 9 0 1 9 16 15 13 2 16 4 7 13 3 13 10 9 16 13 10 0 9 7 9 10 1 9 7 10 10 9 1 10 9 2 2
21 1 10 9 13 2 1 9 0 13 1 9 0 4 3 13 7 13 1 10 9 2
54 3 1 15 2 13 11 2 10 9 1 11 2 2 3 0 1 9 2 7 11 11 11 2 10 9 9 1 10 9 11 2 3 13 1 11 2 2 15 4 1 13 1 11 1 13 10 9 1 13 2 13 10 9 2
16 1 10 9 10 11 3 13 10 9 1 10 10 9 1 12 2
16 10 9 13 1 13 10 9 0 16 13 10 9 1 10 9 2
11 10 9 1 11 15 13 13 1 10 9 2
35 1 10 9 2 7 1 10 4 13 15 1 10 12 9 0 2 13 10 15 3 1 11 1 10 9 2 10 9 4 13 1 9 1 13 2
73 10 9 16 13 1 9 1 9 1 9 1 10 9 1 10 9 11 11 2 4 13 1 11 11 9 1 10 9 11 11 11 11 9 1 10 9 2 11 1 10 11 7 11 1 11 2 2 3 3 10 9 13 1 10 9 1 10 9 11 11 7 11 2 7 4 13 1 10 11 11 1 11 2
38 15 13 1 10 9 1 11 3 1 10 9 11 11 7 3 1 10 9 0 1 2 10 11 2 2 11 12 1 11 2 13 3 1 10 9 11 11 2
51 1 9 1 10 9 0 2 15 13 10 9 0 1 10 9 1 11 2 10 0 9 0 1 11 2 16 15 13 1 9 1 10 9 0 1 12 9 2 1 16 15 13 10 9 1 10 11 11 11 11 2
21 1 12 4 13 1 10 11 1 9 1 9 2 13 0 7 13 1 12 7 12 2
40 10 12 1 11 1 12 4 13 9 1 10 9 0 1 10 9 1 11 11 1 11 11 1 10 11 7 10 12 1 11 1 12 4 13 1 9 1 10 9 2
21 1 10 9 1 10 15 10 9 13 1 9 7 9 2 10 9 15 13 1 9 2
5 3 3 13 9 2
32 10 9 0 16 2 1 10 13 15 1 10 0 9 0 1 10 9 0 2 4 13 10 9 1 10 9 1 9 1 9 0 2
7 2 3 3 12 9 2 2
22 2 1 15 3 13 10 9 2 7 13 10 9 1 10 9 7 13 15 13 10 9 2
13 10 9 4 13 1 10 9 1 10 9 11 11 2
19 11 11 13 10 0 9 1 10 9 2 10 9 0 1 11 13 11 11 2
7 11 12 1 11 1 12 2
40 3 2 10 9 13 16 2 3 13 9 1 9 3 1 10 9 16 13 13 10 9 2 3 7 13 0 13 1 9 1 0 9 1 9 1 9 1 9 2 2
18 10 9 0 13 1 12 7 12 2 15 0 13 1 12 1 12 2 2
35 1 10 0 9 13 13 15 1 11 11 2 3 15 13 3 1 11 1 11 2 1 10 9 0 13 9 1 10 9 0 1 11 2 11 2
20 11 11 11 13 16 10 9 3 0 13 10 9 1 13 1 15 13 10 9 2
14 13 1 9 13 13 9 1 0 9 2 9 7 9 2
48 10 0 12 1 11 1 12 2 11 11 2 1 11 2 13 10 9 0 1 10 0 9 1 10 9 2 2 1 10 9 1 11 2 13 1 10 9 1 10 9 1 10 9 1 10 8 9 2
19 10 9 1 10 9 1 10 9 13 10 9 3 0 7 15 1 10 9 2
40 3 15 4 13 10 9 2 11 11 2 15 3 4 13 16 10 9 1 10 9 1 10 9 0 15 13 1 10 9 10 0 12 1 11 1 12 5 5 9 2
34 10 9 13 3 1 10 11 11 1 11 1 11 2 11 2 13 1 9 1 10 0 9 1 10 8 1 9 16 4 13 10 0 9 2
16 4 13 10 9 3 7 1 15 1 9 3 0 13 10 9 2
32 1 12 2 10 9 1 11 13 1 10 9 1 9 2 16 11 12 1 11 13 2 13 10 0 9 0 1 10 9 1 11 2
22 1 12 11 15 13 1 9 0 1 11 11 2 3 3 10 9 1 10 9 0 0 2
35 10 12 9 13 3 1 10 0 9 1 10 9 1 10 9 12 10 9 1 12 9 1 10 12 9 2 13 1 10 9 1 9 7 9 2
6 1 9 13 9 0 2
31 10 13 10 9 1 10 9 1 9 1 10 2 9 1 9 2 2 11 11 2 2 1 10 0 8 1 10 11 1 12 2
33 3 1 9 2 10 9 1 10 11 15 4 13 1 9 0 13 1 10 9 2 13 10 9 7 10 9 2 10 11 1 11 11 2
19 10 9 0 15 13 10 9 2 9 2 9 7 10 10 9 1 10 9 2
15 10 9 13 15 13 1 11 16 11 4 4 13 1 11 2
16 16 13 0 1 16 10 9 13 0 4 4 15 1 13 15 2
30 3 7 1 10 9 0 2 10 9 0 1 10 9 13 7 13 1 10 9 0 2 15 16 1 0 13 3 10 9 2
16 1 10 9 10 11 11 9 0 13 11 15 13 10 0 9 2
20 13 3 9 10 9 3 0 2 13 1 10 9 1 10 9 7 10 9 0 2
38 10 12 1 11 1 12 2 10 9 1 10 9 0 1 10 11 1 11 13 1 9 16 12 1 10 9 16 13 15 1 10 9 13 7 12 13 0 2
23 1 15 2 10 11 11 13 12 9 1 7 9 7 9 15 13 1 9 1 10 9 0 2
30 11 4 13 1 0 9 1 9 2 13 10 9 8 2 0 1 11 1 11 11 2 7 13 1 10 9 1 11 12 2
23 15 2 1 10 11 11 7 10 11 11 15 13 1 13 3 15 1 10 9 1 10 9 2
44 10 9 0 2 11 1 11 7 11 1 11 2 11 2 13 1 10 9 1 10 13 15 2 7 11 11 1 11 2 1 10 13 15 1 10 9 1 12 2 13 13 10 9 2
45 10 9 0 0 13 10 9 1 10 9 13 1 10 9 1 10 9 1 11 2 10 9 13 9 1 10 9 1 10 9 1 11 2 3 1 10 9 1 11 7 3 1 10 9 2
16 11 15 13 1 10 0 9 11 2 3 13 1 10 9 0 2
71 10 9 1 11 11 2 11 2 13 10 9 0 2 1 9 0 7 1 9 1 9 13 1 12 1 10 9 1 13 10 9 1 10 9 1 9 1 11 2 13 1 10 9 1 9 0 2 13 1 9 1 9 2 9 7 9 0 2 13 10 9 0 1 10 9 7 9 1 10 9 2
41 10 9 15 13 1 10 9 2 16 3 1 1 9 2 15 4 13 16 13 16 10 9 15 13 3 1 10 9 2 15 1 10 0 9 1 9 1 10 0 9 2
15 10 9 13 10 9 1 10 9 0 1 11 11 1 11 2
14 10 0 9 9 1 10 9 1 10 9 1 1 11 2
33 1 10 9 0 2 11 11 4 13 1 10 9 3 0 2 13 1 10 9 9 1 10 9 11 2 7 0 9 1 10 9 0 2
11 3 15 15 13 10 9 1 11 1 11 2
23 10 9 13 10 0 9 2 13 0 12 9 2 2 11 11 11 11 2 7 2 11 2 2
32 1 11 2 1 9 2 10 10 9 15 13 1 0 9 1 9 1 9 7 9 2 13 10 9 1 10 15 10 9 4 13 2
48 1 10 9 4 13 10 9 1 8 8 2 9 0 7 9 0 2 9 8 1 9 0 7 0 2 16 13 13 1 10 9 1 12 9 13 1 10 3 0 9 7 1 10 9 1 0 9 2
24 11 11 11 2 9 1 10 11 11 13 1 11 2 13 1 11 16 15 13 9 1 10 9 2
11 15 13 2 3 3 2 1 10 9 0 2
58 13 15 15 3 2 10 9 15 4 13 15 3 3 9 1 10 9 1 10 9 7 10 9 2 16 15 13 10 9 16 11 13 1 10 9 1 2 11 2 1 11 11 2 1 10 15 3 15 13 7 3 2 13 10 0 9 2 2
13 10 9 4 1 13 15 10 12 1 11 1 12 2
24 11 1 11 13 10 9 1 10 9 12 7 12 1 10 9 1 11 13 1 10 9 1 11 2
15 13 3 0 1 4 13 1 15 2 9 0 7 3 0 2
55 3 3 2 16 13 9 2 15 13 1 10 9 10 9 1 9 1 10 9 1 9 16 15 4 13 1 10 9 1 11 2 11 2 3 7 1 10 9 3 4 13 10 9 1 3 13 10 11 1 10 9 1 11 12 2
41 1 9 1 11 2 2 11 11 11 11 11 11 11 11 2 13 10 9 0 3 0 1 10 10 9 1 11 11 1 10 0 9 1 11 11 2 10 11 11 12 2
31 3 13 10 9 2 11 11 1 11 7 1 11 2 7 9 1 10 9 2 11 2 10 11 2 11 2 11 7 11 2 2
47 1 13 15 0 10 2 9 11 2 2 11 2 1 9 1 11 11 2 13 10 9 1 10 9 11 11 2 16 13 4 13 9 1 11 2 1 13 9 0 2 9 1 10 16 4 13 2
6 9 7 13 1 8 2
47 11 11 2 13 1 11 1 10 11 1 11 7 1 11 1 11 3 7 10 11 2 13 10 9 0 1 12 2 1 10 9 9 2 13 1 11 2 11 2 1 10 9 13 1 11 11 2
30 1 9 2 16 3 13 0 1 10 12 1 11 2 10 9 16 4 13 9 1 10 0 9 3 13 9 1 10 9 2
20 15 16 13 0 16 2 16 13 3 2 10 9 3 4 3 13 1 10 9 2
18 10 9 1 10 11 11 1 10 9 1 10 9 1 11 13 10 9 2
21 16 3 13 0 13 1 16 11 15 4 13 1 11 2 16 4 13 10 9 2 2
31 16 13 10 9 1 13 1 10 9 2 10 9 13 13 1 10 11 11 2 3 16 10 0 9 13 10 9 1 10 9 2
44 10 9 15 13 1 10 9 1 0 9 0 2 7 13 2 1 10 0 9 1 10 9 2 10 3 0 9 2 1 9 10 9 1 11 13 15 16 15 13 13 10 0 9 2
18 10 0 9 0 13 10 9 1 13 9 0 0 1 10 9 7 9 2
16 10 9 1 9 13 10 9 1 9 1 11 2 1 11 11 2
14 13 0 9 1 9 2 9 2 9 2 0 7 0 2
19 13 10 9 1 12 9 5 2 10 9 15 13 1 10 12 1 12 9 2
10 9 7 9 1 10 9 1 10 9 2
7 13 3 10 9 1 9 2
12 1 10 9 2 15 4 13 9 1 11 11 2
31 1 9 2 16 4 13 1 10 9 1 9 1 10 9 7 9 2 4 13 1 10 9 0 10 9 7 0 9 1 11 2
22 11 13 10 0 9 1 9 0 7 13 1 10 9 1 10 0 9 13 10 9 11 2
17 10 11 1 11 11 1 11 7 10 9 1 11 4 13 10 9 2
22 1 10 0 9 4 4 13 1 13 9 1 9 1 0 9 7 15 4 13 10 9 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 13 1 9 0 7 2 12 5 2 12 5 5 13 9 2
30 10 9 1 10 9 11 2 11 2 13 10 9 16 13 10 9 16 4 13 9 0 2 1 3 10 9 1 10 9 2
28 1 3 1 12 9 13 9 1 10 9 1 10 11 11 1 11 1 10 11 1 11 2 3 7 1 10 9 2
67 7 3 1 10 12 9 9 1 10 9 0 1 10 9 2 4 13 10 9 1 3 9 0 7 1 0 9 2 1 2 10 9 2 2 1 11 11 2 16 13 10 9 1 11 11 7 16 13 10 0 9 1 10 16 13 10 11 11 16 13 10 9 1 10 0 9 2
18 1 12 2 10 9 1 9 13 10 11 1 10 9 1 10 11 0 2
13 10 9 15 13 16 13 10 9 1 9 0 0 2
9 13 3 3 1 10 9 1 11 2
17 11 11 4 13 1 11 11 1 11 7 13 1 11 12 2 12 2
13 10 9 0 1 11 13 10 9 1 12 9 5 2
52 1 10 9 2 10 9 0 1 11 11 2 11 2 11 13 3 7 10 9 0 2 13 0 2 7 13 16 11 2 15 4 1 13 1 10 9 2 1 10 9 2 16 15 4 13 10 9 0 2 13 2 2
20 15 15 13 2 7 11 15 13 16 3 13 10 9 2 7 15 13 1 15 2
15 4 13 10 9 7 13 0 2 15 10 9 7 10 9 2
25 16 3 13 9 0 2 3 13 10 9 0 0 1 10 9 9 1 10 9 1 10 9 0 0 2
51 10 11 11 1 11 13 13 9 0 1 10 0 9 2 1 10 1 10 9 7 0 16 13 15 16 4 13 10 9 1 0 9 7 15 13 10 9 1 12 9 1 9 16 13 15 16 4 13 1 9 2
36 9 2 9 0 7 9 0 13 9 13 1 10 0 9 0 1 13 15 1 10 9 0 16 15 13 1 10 9 12 1 10 9 0 1 11 2
12 13 10 9 0 16 13 1 12 9 1 9 2
21 13 10 0 9 1 13 10 9 2 3 1 16 4 13 1 10 9 9 1 12 2
36 15 13 16 10 9 1 10 9 1 10 9 0 1 13 10 9 13 1 10 0 9 1 10 9 1 9 2 1 15 15 1 10 0 9 0 2
28 10 9 3 4 13 1 10 9 11 1 10 0 9 1 10 9 1 12 2 16 13 1 2 11 2 1 11 2
25 11 13 1 11 16 15 15 13 2 7 15 15 13 16 13 10 9 0 2 7 3 13 15 9 2
32 13 1 10 9 1 11 1 12 2 13 10 9 3 0 1 11 7 10 9 1 13 1 10 9 1 10 9 1 10 11 11 2
29 1 15 2 13 0 13 10 11 1 10 11 2 16 13 3 10 9 1 10 9 1 9 13 1 9 1 10 9 2
19 1 10 9 15 13 1 10 11 1 11 16 13 10 9 0 1 10 9 2
23 1 10 9 1 11 2 13 10 9 1 9 2 9 2 9 7 2 1 0 9 2 9 2
24 10 9 1 10 9 1 10 9 0 15 13 13 1 10 9 10 11 2 1 10 11 1 11 2
19 1 9 2 10 9 15 13 3 16 13 16 10 9 2 11 15 13 0 2
36 11 11 11 11 2 12 1 11 8 1 11 12 2 2 13 10 9 2 9 2 11 2 9 0 2 9 1 9 1 10 9 1 11 1 11 2
27 15 9 3 13 10 9 2 13 10 11 11 11 7 10 9 1 10 0 9 0 1 10 9 1 10 9 2
33 11 11 12 11 11 11 13 10 9 1 9 2 1 9 13 1 10 11 11 12 2 13 1 12 1 10 9 1 9 0 11 11 2
105 1 10 9 1 13 1 9 10 0 9 16 15 4 13 1 10 9 7 9 1 10 0 11 1 10 11 2 11 1 11 2 7 13 9 1 9 1 10 9 1 9 0 2 4 13 15 16 15 13 10 0 9 2 15 4 13 1 16 2 1 3 2 7 3 13 1 10 9 16 13 16 10 9 3 13 9 2 13 15 1 10 9 1 10 15 15 15 4 13 3 9 2 7 16 15 15 4 13 2 3 3 15 13 0 2
45 11 2 11 11 2 2 10 0 9 0 2 13 10 9 3 0 2 13 10 9 1 10 15 13 11 11 2 10 9 1 0 9 1 10 9 0 7 16 13 10 9 0 1 9 2
41 10 9 13 1 12 9 2 2 11 2 1 11 2 2 11 10 11 1 11 2 1 11 11 2 2 11 1 11 2 1 11 7 2 11 1 11 2 1 10 11 2
139 3 13 10 9 2 3 2 10 0 9 0 7 0 1 10 9 0 2 10 9 0 0 7 10 0 9 0 2 16 15 4 13 2 3 3 16 13 10 9 0 1 11 7 10 9 1 10 9 1 10 9 0 1 11 2 7 16 13 12 9 0 1 9 1 10 0 9 1 10 9 1 10 9 2 1 10 13 0 1 12 9 0 1 10 9 1 9 1 10 0 9 1 10 11 11 7 10 9 0 2 1 9 1 16 15 13 10 0 9 1 9 0 1 10 9 0 0 7 2 10 11 11 15 13 0 1 10 0 9 0 1 10 9 1 10 9 0 0 2
15 1 1 11 1 12 2 12 9 1 10 9 13 1 9 2
30 11 10 11 1 10 2 11 11 2 10 9 0 1 11 1 9 1 10 9 2 10 9 1 11 3 4 13 1 11 2
19 3 15 4 13 1 10 9 2 10 9 1 10 9 13 1 8 1 11 2
20 0 2 11 13 1 11 7 1 11 1 10 9 1 9 1 10 9 1 11 2
66 1 10 9 1 10 9 2 10 9 0 1 10 9 0 4 13 1 13 1 14 2 9 1 10 9 1 9 1 10 14 2 9 2 11 2 11 2 2 12 2 9 2 11 11 11 2 11 2 7 11 11 2 11 2 16 13 9 0 1 10 8 2 9 1 9 2
47 1 10 0 9 2 16 13 10 12 1 11 2 11 11 13 10 10 9 1 9 1 13 1 10 9 2 13 10 0 9 1 8 1 10 9 13 1 10 11 11 1 11 1 12 1 11 2
20 10 9 13 10 9 1 9 2 10 9 16 10 15 4 13 7 10 0 9 2
20 15 13 10 9 3 0 2 3 0 1 10 9 7 0 1 10 9 1 9 2
28 10 9 4 13 3 0 2 10 9 13 3 0 7 13 13 15 9 1 10 9 7 15 9 1 10 9 0 2
21 10 9 1 10 9 1 9 1 9 13 1 12 1 10 9 0 1 10 9 0 2
38 1 3 10 9 4 1 13 10 9 0 0 7 10 9 0 1 10 0 11 3 4 1 13 15 1 15 1 10 9 1 9 1 12 2 12 7 12 2
30 10 12 5 1 10 9 1 10 9 1 10 9 1 10 9 13 1 9 0 1 10 9 1 12 9 2 12 9 2 2
113 10 9 1 10 9 1 11 11 13 3 0 1 13 15 1 10 0 9 0 16 13 1 10 11 11 7 1 10 15 13 10 9 11 13 10 0 9 1 10 11 1 11 2 10 9 1 10 9 13 1 10 12 9 1 10 9 1 10 9 1 10 10 9 1 10 9 1 10 12 9 1 10 9 1 10 9 16 15 13 1 10 0 9 1 10 9 16 15 13 1 15 0 9 1 10 9 3 1 10 9 1 10 9 1 11 7 16 3 13 11 1 11 2
30 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 5 12 7 10 9 0 1 9 13 5 12 2
24 10 9 0 2 13 1 10 9 0 2 13 1 10 2 9 2 1 2 9 2 1 10 9 2
38 3 2 10 9 11 4 13 10 9 0 1 10 9 1 10 0 9 1 9 2 11 11 4 13 1 9 1 10 9 1 9 1 10 12 9 1 9 2
16 13 1 9 0 7 13 10 3 0 1 10 9 1 10 11 2
36 3 2 10 9 9 3 13 10 9 7 9 0 0 2 4 13 0 1 10 0 9 0 2 0 0 2 16 15 13 1 10 9 0 2 9 2
90 15 15 13 13 10 0 9 1 10 9 1 11 2 1 10 9 0 0 1 10 12 9 1 10 9 2 10 9 0 2 10 9 1 10 9 2 7 10 9 0 16 15 9 2 7 3 2 7 11 11 2 7 11 1 11 2 1 10 9 1 11 7 11 2 13 2 13 1 11 2 16 10 0 9 15 13 11 2 10 3 0 7 0 1 10 9 1 10 9 2
50 3 2 11 13 16 10 11 3 13 10 9 1 9 1 9 1 9 1 9 1 10 9 1 10 9 0 2 7 1 10 9 2 10 9 1 9 13 3 15 16 13 10 9 1 12 12 9 10 9 2
69 15 13 2 16 1 9 1 10 9 0 1 9 1 9 0 2 1 12 1 11 2 15 12 2 12 2 16 10 9 13 10 9 1 9 0 4 13 3 1 10 9 1 10 9 1 10 9 7 9 1 10 9 1 10 9 1 10 9 2 3 13 1 10 11 1 11 1 11 2
31 1 10 9 0 9 2 13 10 9 1 10 9 2 0 1 10 9 2 10 9 2 10 9 2 7 10 9 1 9 0 2
22 0 13 10 9 16 15 13 10 9 7 3 3 15 2 7 3 10 9 1 10 9 2
36 13 1 10 9 1 9 1 9 0 7 9 2 10 9 13 0 1 10 11 2 1 10 12 9 13 1 11 11 2 3 12 15 13 1 11 2
75 1 10 9 1 9 1 9 0 2 1 9 1 10 12 1 11 1 12 2 10 9 0 1 9 7 9 0 13 1 10 11 16 13 10 9 1 9 2 15 3 3 3 4 13 1 10 9 2 7 16 3 2 13 0 7 1 10 0 9 0 7 0 2 16 13 10 9 13 1 10 8 7 10 9 2
17 13 10 9 16 13 1 9 0 7 0 10 9 0 1 10 9 2
23 4 13 1 10 0 9 2 12 5 2 1 10 9 1 10 11 1 12 1 10 11 11 2
14 9 11 13 10 9 1 10 9 1 10 9 1 11 2
26 10 9 0 11 4 13 13 15 1 10 11 1 11 7 13 3 1 10 11 1 11 1 10 0 9 2
32 13 1 15 16 13 10 9 0 1 10 9 1 11 2 7 3 13 1 3 1 12 9 1 10 11 11 7 1 10 11 11 2
58 3 3 1 10 9 0 2 13 16 10 9 13 3 16 10 11 3 13 9 1 10 9 0 1 7 13 1 10 9 1 10 11 2 1 11 2 10 9 16 13 10 9 13 10 9 2 3 1 10 9 1 10 0 9 1 10 9 2
28 1 10 9 4 13 2 13 7 3 15 13 15 2 1 15 1 10 11 11 2 9 3 13 9 3 9 3 2
10 10 9 4 13 1 10 9 11 11 2
22 11 11 13 10 9 1 9 0 1 10 9 11 2 9 1 10 0 9 0 11 11 2
13 10 9 2 12 2 3 13 9 2 9 7 9 2
22 11 11 13 10 9 1 9 0 16 13 1 10 11 1 10 11 1 10 0 9 0 2
23 10 9 13 1 10 9 1 10 0 9 11 11 2 1 15 15 4 13 10 9 1 9 2
28 3 0 9 2 1 15 1 10 10 9 2 15 13 3 3 7 15 13 10 9 1 10 9 8 3 0 9 2
15 10 9 13 0 2 0 2 0 2 1 8 9 1 9 2
33 1 9 12 9 2 13 3 1 9 2 10 11 2 2 9 1 8 2 9 1 9 2 9 1 9 2 9 2 9 0 7 9 2
14 1 10 9 2 13 13 15 1 10 9 1 10 9 2
28 15 15 13 3 1 15 2 15 13 10 9 1 9 7 3 15 13 12 9 1 9 1 7 13 4 1 13 2
40 10 9 2 1 10 15 15 15 13 10 9 1 11 3 13 15 2 13 13 2 10 2 9 2 2 13 15 1 10 10 9 1 9 0 16 4 13 3 15 2
21 3 10 9 1 9 0 4 13 0 1 9 0 2 7 1 9 1 9 1 9 2
43 13 1 10 9 1 9 2 10 9 1 11 2 1 9 1 10 9 2 1 11 1 12 2 7 10 9 1 11 7 11 11 1 10 11 2 1 11 1 12 2 1 15 2
6 10 9 15 4 13 2
15 1 12 13 1 11 11 7 1 10 9 0 1 11 11 2
8 13 13 1 9 7 3 13 2
28 2 10 9 13 1 10 9 7 13 15 15 16 4 7 13 15 1 9 7 13 10 9 1 10 9 2 13 2
14 15 16 13 1 10 0 9 1 10 11 4 3 13 2
21 10 9 15 13 0 1 10 9 1 10 11 11 2 1 10 9 1 10 9 11 2
8 13 10 12 1 11 1 12 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
12 13 11 11 1 10 11 1 11 12 10 11 2
50 10 9 0 2 10 0 1 10 12 9 16 13 10 9 0 2 13 1 10 9 0 7 10 5 9 1 10 9 2 1 10 9 7 1 10 9 1 10 9 2 3 7 12 1 10 13 0 1 11 2
24 10 9 0 13 1 10 9 7 13 10 9 2 13 16 10 9 15 13 1 9 1 10 9 2
18 1 12 13 10 0 9 1 9 3 0 2 2 10 11 1 11 2 2
12 10 9 1 10 9 13 1 10 9 11 11 2
68 11 4 13 15 3 16 15 13 8 2 1 9 2 10 15 13 10 9 13 10 9 7 13 10 9 0 2 16 15 13 13 3 0 2 7 13 0 13 15 2 15 2 13 16 15 4 13 1 9 7 9 2 13 10 9 7 1 0 9 1 10 9 0 1 10 8 11 2
21 15 13 1 10 9 1 11 2 11 2 3 1 10 9 0 2 2 11 7 11 2
25 10 11 13 10 0 9 1 9 2 3 1 10 9 1 10 9 1 10 9 13 1 10 9 0 2
11 1 15 15 2 3 13 9 1 13 15 2
26 1 9 2 13 10 9 1 10 9 1 11 3 13 9 1 10 9 0 0 2 7 1 10 11 2 2
82 10 9 0 1 10 9 0 2 11 2 1 10 9 1 9 2 2 13 2 7 16 10 9 0 13 1 10 9 1 9 0 15 4 13 1 10 0 9 1 9 2 2 2 10 9 13 1 10 9 0 13 1 10 9 4 13 0 2 7 13 1 0 9 1 10 9 1 10 9 1 9 0 2 16 13 0 1 13 1 10 9 2
19 15 13 1 10 0 9 13 1 9 1 0 9 1 9 13 1 9 0 2
43 1 10 9 1 10 9 0 2 11 13 1 10 10 9 1 10 9 3 10 1 11 2 11 2 11 7 11 2 1 10 15 15 13 11 1 10 9 1 11 1 12 2 2
33 1 12 2 10 9 1 9 8 4 13 1 10 9 1 11 2 1 10 9 1 11 11 2 7 13 10 9 1 11 11 1 11 2
13 1 10 9 2 11 15 13 13 15 1 10 9 2
28 3 13 0 0 1 11 11 1 10 11 1 10 11 16 15 13 10 10 9 1 11 10 11 11 1 10 11 2
32 15 13 1 10 0 9 0 1 10 9 1 9 1 9 16 13 13 1 10 9 16 4 13 9 1 10 9 0 1 10 9 2
14 3 13 0 1 10 9 2 1 0 9 7 9 0 2
18 13 10 9 1 11 11 2 11 7 10 9 1 10 9 11 2 11 2
100 10 12 1 11 4 1 13 1 11 2 1 9 2 10 11 11 1 10 11 2 13 16 10 11 11 13 1 10 12 9 1 13 15 1 3 1 10 9 9 2 10 11 11 13 10 9 1 12 9 7 13 3 12 9 1 9 1 9 2 10 11 11 13 12 9 2 16 13 15 12 9 1 3 1 10 9 0 2 7 10 11 11 13 3 1 12 9 3 1 10 0 9 2 1 10 13 10 12 9 2
20 13 3 1 10 11 1 10 11 1 11 1 12 2 13 10 0 9 1 9 2
26 10 9 1 9 1 10 9 13 1 9 12 7 10 12 5 1 10 9 13 1 10 9 1 9 0 2
31 1 9 2 16 11 13 16 10 9 12 13 1 9 10 11 11 11 2 15 15 13 16 13 16 15 13 1 15 10 9 2
16 10 9 1 9 4 4 13 1 10 9 1 9 0 11 11 2
7 11 13 10 9 1 12 2
36 13 10 9 13 2 9 1 9 2 2 1 9 2 2 11 2 2 3 0 1 10 9 2 2 16 13 1 0 9 1 9 13 1 9 0 2
15 1 10 9 10 9 3 13 1 13 10 10 9 1 9 2
40 1 10 9 0 1 10 9 7 1 10 10 9 1 9 4 13 10 9 2 10 10 9 0 13 10 9 16 13 3 1 9 1 10 9 2 1 9 1 9 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
19 1 10 9 12 7 1 10 9 12 2 10 9 1 10 9 13 11 11 2
44 11 11 13 10 9 1 10 0 9 1 11 2 13 1 10 9 11 11 1 9 1 10 0 9 7 11 1 10 0 1 10 9 1 10 9 2 13 1 9 1 10 9 2 2
20 0 13 3 16 16 4 13 12 7 12 9 1 10 11 3 15 15 13 0 2
23 10 0 9 2 11 11 15 13 1 10 11 2 11 2 9 0 2 11 2 11 7 11 2
38 1 15 15 13 1 9 0 7 0 2 1 10 9 1 9 0 7 10 9 0 2 7 10 9 1 9 0 7 1 10 9 1 9 1 9 1 9 2
51 10 9 13 0 2 7 3 0 7 15 1 10 10 9 1 9 2 0 2 0 2 12 9 1 0 7 12 9 1 9 16 13 0 2 13 15 3 1 12 9 2 3 15 0 1 10 9 0 1 9 2
27 10 9 11 8 1 11 11 7 10 9 0 1 11 13 11 11 1 10 9 1 9 1 10 9 11 11 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
28 11 1 10 9 0 2 9 7 9 2 4 13 1 10 9 2 3 16 3 13 10 9 1 9 1 10 9 2
16 10 9 13 3 0 7 13 0 2 0 2 1 10 9 0 2
41 1 10 9 2 16 13 10 9 1 10 9 0 2 11 13 1 10 9 1 10 9 2 1 13 15 1 9 0 1 10 9 7 13 13 10 9 1 12 13 9 2
28 1 3 13 16 3 13 2 1 10 9 0 2 7 16 15 4 13 10 9 1 9 2 9 2 9 7 9 2
25 3 10 9 13 9 0 1 10 9 3 1 15 2 15 16 13 10 0 7 0 9 1 10 9 2
31 1 9 2 1 9 1 10 11 11 2 11 13 10 9 3 1 10 9 7 13 10 9 1 10 9 11 11 1 10 9 2
25 10 9 1 10 9 9 13 1 9 16 10 9 13 9 1 10 9 2 16 3 15 13 1 15 2
42 11 13 10 9 7 9 0 2 1 10 9 1 11 1 10 11 2 9 1 11 2 1 10 9 1 10 11 2 11 7 9 1 11 2 11 2 11 2 1 2 11 2
41 1 13 15 1 10 9 0 1 10 9 2 10 12 9 13 3 10 9 7 9 1 10 9 2 0 1 10 9 2 16 13 10 9 1 10 9 1 10 0 9 2
20 10 0 9 0 15 4 13 1 13 9 9 1 0 9 1 10 11 2 12 2
30 11 13 3 10 9 0 2 1 15 1 7 4 13 15 1 10 11 11 2 16 15 13 0 9 1 15 1 9 0 2
16 15 13 1 10 9 10 12 1 11 1 12 1 10 0 9 2
11 13 1 11 2 10 12 1 11 1 12 2
37 1 10 11 13 10 9 0 7 1 10 11 11 13 9 3 1 4 13 1 10 9 7 16 13 11 13 0 16 13 9 1 3 1 9 1 3 2
23 3 13 1 9 3 0 1 11 13 9 13 1 11 7 13 15 1 10 11 1 10 11 2
29 1 12 2 10 9 1 11 13 1 10 9 1 11 1 9 1 10 9 7 10 9 1 10 9 0 1 9 0 2
26 10 0 9 13 1 10 9 12 2 7 1 13 1 10 0 9 13 1 12 13 10 9 1 9 0 2
24 3 12 9 3 1 10 9 1 10 9 2 11 13 10 9 10 11 1 10 9 11 1 12 2
43 13 10 9 1 11 11 1 10 9 1 12 9 2 10 12 1 11 1 12 2 1 10 9 1 10 9 11 11 9 1 11 1 12 1 12 2 13 1 9 1 11 11 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
34 10 9 4 13 13 1 9 2 3 16 1 9 1 10 9 1 10 9 11 11 11 2 11 13 0 3 7 16 11 13 10 9 0 2
15 1 9 1 13 10 9 1 9 2 10 9 4 3 13 2
19 10 9 13 1 10 9 1 10 0 11 2 16 13 10 9 1 12 9 2
40 3 13 10 9 1 9 0 1 10 9 2 16 16 4 13 10 9 4 13 15 3 1 10 9 1 7 15 15 13 2 16 13 1 10 10 9 16 15 13 2
29 1 11 1 12 15 15 13 10 9 1 11 2 11 1 10 9 2 1 16 15 13 10 9 12 1 11 1 12 2
21 13 1 12 9 1 10 11 1 10 11 1 11 2 13 10 9 1 10 9 0 2
33 11 13 0 9 7 1 10 9 0 13 3 9 1 4 4 13 1 9 2 3 7 10 9 1 11 11 11 15 4 13 10 9 2
36 10 9 0 2 10 11 11 2 10 11 7 10 9 0 4 13 10 9 3 0 1 9 2 16 15 13 3 1 10 9 0 0 0 1 9 2
50 1 10 0 9 1 10 9 10 9 0 2 13 9 0 2 1 10 9 4 3 13 1 10 9 9 0 2 0 7 9 0 7 2 3 2 1 10 9 1 10 9 7 10 0 11 1 11 1 11 2
27 15 13 16 13 1 10 9 2 7 16 4 13 1 9 16 3 4 13 1 10 0 9 1 10 0 9 2
3 13 0 2
30 1 10 9 4 13 1 10 9 1 11 2 3 11 2 2 7 1 10 9 12 1 10 9 12 15 1 11 1 11 2
61 10 9 10 9 3 0 1 10 9 2 10 9 13 0 1 9 2 13 9 1 10 1 10 11 1 10 9 1 11 2 15 1 10 11 11 7 1 10 11 11 1 10 9 1 10 9 1 11 2 7 10 0 9 0 16 13 10 11 1 11 2
29 3 13 10 9 11 11 11 2 9 0 1 10 9 7 10 9 11 11 2 9 1 9 1 9 1 10 9 0 2
23 10 9 1 10 9 4 13 1 10 9 0 2 3 13 10 9 2 7 2 4 11 13 2
36 13 1 10 11 1 11 10 12 1 11 1 12 7 13 1 10 9 1 13 9 1 10 9 1 9 1 10 12 1 11 16 13 1 11 11 2
7 11 13 10 9 0 0 2
28 10 9 11 13 10 0 9 1 10 9 1 11 2 10 9 1 10 9 11 16 13 9 1 10 9 1 10 11
18 10 9 1 11 4 13 1 11 11 7 13 1 11 11 1 11 11 2
10 11 13 10 9 1 2 9 0 2 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
33 15 13 15 1 10 9 0 3 0 3 1 10 9 7 1 0 9 1 9 2 1 15 15 15 13 1 10 0 1 10 9 0 2
36 10 9 1 9 1 11 2 1 9 2 11 11 11 11 11 11 2 13 10 9 0 1 10 9 1 11 2 3 16 10 9 13 10 9 0 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
44 1 10 11 11 11 2 11 13 1 11 2 11 2 11 2 11 11 2 2 7 1 11 2 11 11 2 1 11 2 10 9 1 10 9 2 2 16 13 1 11 1 10 9 2
43 10 9 15 13 7 13 1 0 9 1 9 10 9 0 11 11 2 8 2 1 10 11 2 11 1 12 5 2 11 2 11 2 2 1 10 9 1 11 2 11 11 2 2
21 10 9 13 3 1 10 9 1 10 9 7 15 13 3 1 15 15 13 11 11 2
8 11 15 13 13 1 10 9 2
25 15 15 10 3 9 13 13 16 10 9 1 10 9 0 13 10 9 0 1 10 9 1 10 9 2
36 10 9 0 7 1 10 15 9 1 10 9 1 10 9 2 15 16 3 13 1 9 15 13 2 10 9 13 0 7 15 13 9 1 10 9 2
16 11 1 11 13 10 9 1 11 1 9 1 9 2 8 2 2
29 1 10 0 9 15 13 10 9 0 1 11 1 12 7 12 1 13 1 10 9 13 1 10 11 11 1 11 0 2
18 16 13 10 0 9 9 2 9 15 13 16 10 9 0 13 3 0 2
59 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 2 3 13 1 2 11 11 2 2 2 11 11 2 7 2 11 11 2 2 13 10 9 0 2 0 9 1 12 9 0 7 10 9 1 0 9 0 1 11 11 7 11 11 2
18 3 15 13 10 9 1 10 2 0 9 2 16 13 13 1 10 9 2
23 13 10 0 9 1 11 2 13 10 9 1 10 15 13 11 7 10 0 9 1 10 9 2
40 10 9 11 4 13 9 7 10 9 13 10 9 16 13 1 11 2 3 13 10 9 3 0 1 10 9 2 15 16 13 13 9 1 10 9 1 12 9 0 2
28 3 4 13 15 1 10 9 7 13 1 10 9 1 10 10 9 0 1 10 11 11 2 11 11 7 10 11 2
19 10 9 0 1 10 9 13 10 11 7 10 11 2 0 1 10 9 11 2
10 13 1 0 9 16 10 9 4 13 2
14 11 1 11 7 11 3 1 9 13 10 9 3 0 2
18 10 9 13 1 9 0 0 2 1 0 9 3 1 12 9 1 0 2
16 13 10 9 0 16 7 15 4 13 2 13 3 0 7 0 2
11 10 9 13 2 3 8 2 7 3 0 2
15 3 11 1 0 9 4 13 1 10 9 1 10 9 0 2
5 15 13 3 3 2
23 1 10 9 13 1 10 12 1 11 1 12 2 11 13 1 12 9 0 13 1 12 9 2
16 1 9 15 13 10 9 1 11 7 1 10 9 10 11 11 2
41 10 9 0 2 16 13 10 9 1 9 2 10 9 2 7 3 0 2 13 10 9 0 1 15 16 4 13 1 10 9 0 2 16 15 13 1 9 1 10 9 2
19 10 9 13 16 15 13 12 9 0 1 4 13 15 16 13 1 10 9 2
94 4 3 7 13 9 1 11 1 10 9 11 11 2 11 1 10 11 11 2 11 1 10 11 11 2 11 1 11 7 15 2 1 11 1 10 12 2 13 13 10 10 9 0 1 10 9 1 10 11 11 7 13 1 10 11 11 11 2 11 2 10 9 7 13 10 9 1 11 11 1 10 11 1 10 0 11 2 10 9 0 15 13 10 9 7 3 13 13 10 9 1 11 11 2
63 10 9 0 13 1 10 9 2 9 1 9 0 1 10 9 2 10 9 0 7 10 9 1 9 1 10 9 2 4 13 16 10 9 13 1 10 9 0 1 10 9 2 3 10 9 0 7 10 9 1 9 9 2 9 7 9 2 4 13 10 0 9 2
22 7 3 1 0 7 0 2 7 1 10 0 9 1 16 10 0 9 3 13 10 9 2
5 10 9 13 11 2
55 3 13 0 1 10 9 1 10 9 2 1 13 15 10 0 9 1 13 7 1 13 10 0 9 1 9 2 7 13 16 3 1 10 0 9 7 9 1 10 9 2 15 13 1 0 7 0 1 13 15 1 10 9 0 2
38 1 9 2 1 9 1 13 10 0 9 2 3 13 1 13 10 9 1 9 1 10 0 9 2 7 1 10 9 11 11 2 10 9 2 13 10 9 2
26 10 9 7 10 9 1 10 9 1 10 9 15 13 1 10 9 7 10 9 1 10 9 1 10 9 2
26 1 10 9 1 10 9 15 13 11 2 10 9 1 11 2 15 15 13 15 15 16 4 13 1 9 2
20 1 12 13 11 11 11 11 2 10 0 9 7 1 12 11 2 10 0 9 2
27 10 9 1 9 14 2 9 0 1 10 9 0 2 16 13 9 2 4 3 13 1 10 9 0 1 11 2
26 10 9 1 9 1 10 9 4 13 1 10 9 1 10 9 0 1 10 9 7 3 2 1 10 9 2
17 1 10 9 0 13 3 15 13 10 9 1 10 9 16 3 0 2
16 1 10 9 15 13 0 9 1 9 1 9 1 9 1 9 2
18 10 9 13 3 15 1 9 1 9 7 10 9 0 16 13 1 9 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
19 3 13 1 10 11 16 13 15 1 10 11 11 1 10 9 1 12 9 2
41 10 9 13 12 9 1 12 1 9 2 9 1 10 9 1 9 1 11 1 10 11 1 10 12 9 0 2 12 8 2 2 3 10 9 1 9 4 1 13 9 2
46 16 10 11 11 13 10 9 1 10 9 5 1 12 2 11 2 3 4 13 1 10 9 1 9 2 13 10 9 1 10 9 2 11 11 11 11 2 2 2 15 13 1 11 2 2 2
19 10 9 1 10 9 15 13 1 10 9 1 10 0 7 0 9 1 11 2
33 13 9 1 0 9 15 13 10 0 9 8 10 9 15 13 10 9 3 0 3 1 10 9 7 9 1 10 9 2 2 13 11 2
27 15 13 2 1 10 9 2 10 0 9 2 10 9 0 3 0 7 3 9 1 10 9 1 10 9 0 2
11 13 1 15 13 3 9 11 11 1 15 2
14 15 4 13 9 1 9 1 11 11 1 11 7 3 2
9 3 3 15 13 1 13 1 11 2
12 12 2 8 2 2 13 1 11 11 1 12 2
16 10 9 1 10 9 11 13 3 0 16 10 9 3 13 0 2
18 1 10 9 4 1 13 10 9 1 10 9 0 10 9 1 10 11 2
10 13 1 9 1 10 9 7 10 9 2
47 1 9 1 12 2 10 9 13 1 12 0 9 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 7 3 11 11 1 10 9 0 2 3 1 11 11 7 13 2 11 12 2 2
40 13 10 11 1 11 11 1 11 1 11 1 10 9 0 1 10 11 1 10 11 2 11 2 11 2 11 2 11 7 11 11 2 13 1 10 9 0 11 11 11
47 10 9 13 10 9 1 10 9 0 2 1 15 15 15 4 13 10 9 1 10 9 16 13 10 9 1 10 11 2 13 10 9 1 10 11 1 10 11 1 10 12 1 11 1 0 9 2
21 13 1 11 7 10 9 1 9 1 12 9 1 15 9 7 10 0 9 1 9 2
12 3 3 2 11 13 10 9 1 10 9 11 2
16 13 10 9 1 11 1 9 2 1 9 15 13 10 9 9 2
32 1 10 9 1 10 9 1 12 2 10 9 0 1 9 1 10 9 13 1 9 12 2 7 10 9 0 1 9 13 9 12 2
8 11 11 11 2 11 2 12 2
14 10 9 0 1 10 9 13 8 2 12 0 9 2 2
24 11 13 9 1 10 9 0 9 12 1 10 11 1 11 16 13 1 10 12 9 1 10 9 2
8 13 10 9 1 9 16 13 2
17 10 9 0 0 2 10 9 0 2 10 9 1 10 9 3 0 2
35 10 9 13 3 0 9 1 9 2 1 10 9 1 9 0 13 1 11 11 1 9 1 10 9 5 7 5 2 1 9 0 1 10 9 2
16 3 13 10 0 9 2 1 9 1 9 7 4 13 1 9 2
16 3 1 10 12 5 1 10 9 13 1 10 9 1 9 0 2
13 10 9 1 9 13 1 12 8 2 2 9 8 2
42 1 13 10 9 1 10 9 0 1 10 9 1 9 1 10 9 0 2 10 9 0 1 9 2 10 9 1 9 1 10 9 7 10 9 1 9 4 4 13 7 13 2
20 1 9 1 11 1 11 3 4 7 13 10 9 1 10 9 1 13 10 9 2
21 1 10 9 1 9 10 9 0 1 10 9 0 11 11 13 10 9 1 10 9 2
21 13 10 9 1 10 9 1 10 9 2 10 9 11 11 7 10 9 11 7 11 2
72 16 10 9 1 13 10 9 1 10 9 1 11 15 4 13 1 10 9 1 11 1 12 2 10 9 13 1 10 0 9 1 11 1 10 3 13 1 10 9 0 2 11 12 4 7 13 1 12 10 0 9 16 13 0 9 1 10 9 1 11 1 11 2 1 3 9 1 10 9 1 11 2
19 7 3 13 1 10 9 12 1 10 0 9 16 15 4 1 13 9 0 2
32 13 1 7 15 13 10 9 7 1 9 1 12 9 16 15 13 2 13 12 9 2 7 10 9 13 1 13 15 1 10 9 2
37 9 1 10 0 9 1 10 9 3 0 1 10 9 7 10 9 3 0 2 11 11 7 11 13 9 0 7 0 16 13 13 10 10 9 1 9 2
7 10 9 13 1 9 0 2
21 13 1 0 1 11 2 7 4 13 3 1 10 0 2 10 9 1 10 11 11 2
39 16 10 9 13 3 12 9 1 15 1 10 11 2 10 9 13 1 12 9 10 9 0 2 13 13 1 10 9 1 11 2 11 1 3 1 10 9 0 2
18 10 12 1 11 2 10 9 11 13 1 12 8 2 12 9 3 2 2
20 13 1 10 11 1 9 0 7 11 1 11 11 10 12 5 1 11 1 12 2
18 1 0 9 10 9 13 10 9 0 7 0 1 10 9 1 10 9 2
30 1 10 9 0 13 10 9 1 10 9 1 10 11 2 11 2 10 0 9 13 13 9 1 11 13 7 13 10 9 2
27 11 2 9 11 1 11 1 11 11 2 13 10 9 1 9 1 10 9 11 1 11 7 10 9 1 11 2
26 13 10 9 0 1 9 7 1 10 4 13 0 9 1 11 2 11 11 2 11 2 11 7 3 11 2
19 10 0 9 13 1 9 0 1 9 1 9 0 7 9 0 1 10 9 2
14 13 3 10 9 2 2 1 15 13 1 10 9 2 2
11 1 9 2 11 13 3 1 9 1 11 2
31 3 15 4 13 10 9 0 2 7 13 9 1 13 9 1 10 9 1 9 2 16 13 10 0 9 1 9 2 9 2 2
20 4 13 1 10 0 9 1 10 11 1 10 11 1 12 1 10 11 11 11 2
28 10 0 9 15 13 1 9 7 0 1 9 0 2 13 1 9 0 2 0 2 9 2 9 7 0 2 0 2
15 3 13 9 1 11 11 2 9 1 10 0 9 16 13 2
23 10 9 4 1 13 1 11 2 3 16 10 0 9 4 13 10 9 3 1 10 9 0 2
47 10 9 12 1 10 11 1 11 1 10 11 11 2 4 13 1 9 10 12 1 11 1 12 2 1 4 13 10 9 1 9 1 9 1 10 9 1 11 16 4 13 9 1 10 11 11 2
23 10 11 11 13 1 10 9 0 10 9 16 13 10 9 1 10 0 9 16 13 1 13 2
19 1 10 9 15 13 10 9 1 10 9 0 13 1 10 9 12 7 12 2
36 10 9 0 13 0 1 10 1 11 2 3 16 3 10 9 0 1 10 9 1 10 9 4 13 10 9 2 1 10 0 9 7 10 9 0 2
22 10 0 9 1 10 9 13 11 11 1 10 9 11 7 11 11 1 10 9 1 9 2
24 10 9 2 1 10 9 2 15 13 3 1 9 16 4 3 13 1 9 1 9 1 10 9 2
12 13 10 9 13 1 12 9 2 9 12 2 2
19 10 9 13 15 0 1 9 1 9 7 9 7 9 1 9 0 2 0 2
15 13 10 9 3 0 1 10 15 16 4 13 1 10 9 2
37 3 15 13 0 1 10 9 0 2 13 1 10 9 1 9 2 13 1 10 9 0 10 12 1 11 1 12 1 10 9 1 10 11 1 10 11 2
16 4 13 10 9 0 7 15 16 13 11 1 10 11 13 0 2
41 1 12 10 12 9 15 13 1 11 2 11 2 13 10 9 1 10 0 9 2 11 2 11 2 1 10 10 9 16 10 0 9 13 10 9 1 10 9 0 11 2
12 11 11 13 10 9 1 9 1 10 9 11 2
29 1 12 13 1 11 1 11 1 10 9 1 11 2 3 13 10 9 1 10 9 0 7 13 10 9 0 1 12 2
13 3 1 13 1 15 4 13 1 10 9 1 11 2
43 11 13 1 12 0 9 0 2 16 1 15 9 1 10 0 9 1 9 16 15 13 1 10 9 0 2 3 13 10 9 7 9 1 10 9 1 3 0 9 1 10 9 2
24 9 0 7 0 4 3 13 10 10 9 0 2 7 16 10 9 3 4 13 9 1 0 9 2
7 13 1 10 9 11 2 2
34 7 16 3 15 15 13 10 9 0 13 1 10 9 2 9 1 10 9 2 13 10 9 1 10 9 1 9 1 4 4 13 10 9 2
23 15 13 10 9 7 11 15 13 15 2 7 3 13 1 9 1 10 13 1 11 1 9 2
28 10 9 1 9 16 15 13 9 1 10 9 1 10 9 1 10 0 9 1 10 9 0 7 10 9 3 0 2
19 10 9 15 13 1 15 1 10 9 0 0 1 10 9 1 10 11 0 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
110 10 9 2 9 2 9 7 9 15 13 3 1 10 9 1 10 9 7 1 15 15 13 10 9 1 9 2 11 2 2 3 1 10 15 13 10 9 1 9 1 9 1 9 2 9 1 9 13 7 9 1 9 0 13 15 1 13 3 1 13 2 10 2 9 2 1 10 9 15 13 16 10 9 13 1 10 0 2 9 1 10 9 2 16 13 1 11 2 1 10 0 11 2 13 10 11 1 10 9 1 11 7 13 1 10 9 1 10 11 2
8 11 15 13 0 1 10 9 2
85 13 1 10 9 0 1 10 9 0 2 16 13 10 11 11 11 2 11 12 1 11 2 11 11 2 11 11 2 3 15 13 10 9 0 10 2 9 2 2 1 10 9 0 2 13 9 10 9 1 10 9 11 11 2 10 9 1 10 9 0 2 10 9 1 10 0 9 2 1 10 9 0 7 10 9 1 10 9 16 13 0 1 10 9 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
30 15 1 10 9 4 13 1 10 9 0 2 1 10 9 11 2 10 11 7 10 11 2 3 7 1 9 1 10 9 2
40 2 11 2 13 3 13 15 1 10 11 11 1 11 7 15 13 15 1 10 9 1 13 10 9 0 2 1 9 2 2 11 2 13 9 10 9 1 10 9 2
21 7 2 15 4 13 2 3 13 1 10 9 0 1 10 9 1 9 1 9 0 2
26 1 10 9 2 10 9 13 10 9 0 7 10 9 0 15 13 1 9 1 10 9 1 9 10 9 2
31 11 2 9 1 10 9 1 10 9 0 8 2 4 13 1 9 12 9 0 1 9 7 9 0 1 9 1 10 0 9 2
27 10 9 1 11 11 1 10 11 13 10 9 0 2 1 11 2 10 9 1 9 1 10 9 1 10 9 2
19 13 10 9 1 9 1 12 2 11 11 1 11 2 1 9 1 11 11 2
48 2 10 9 0 1 9 0 7 0 2 10 9 11 11 2 13 3 1 11 16 11 3 15 4 13 1 10 9 0 2 15 16 15 4 13 13 15 1 10 9 1 9 3 13 1 10 11 2
32 10 9 1 11 3 13 9 0 2 7 10 11 11 3 4 13 15 2 3 7 3 10 11 1 10 11 2 3 3 13 11 2
12 2 8 2 13 10 9 0 1 10 9 0 2
14 10 9 13 10 9 0 1 10 9 3 1 10 9 2
32 1 10 9 15 13 0 1 12 9 1 10 9 1 10 9 0 1 10 11 2 11 1 10 11 2 11 2 11 11 7 11 2
12 4 13 0 9 1 9 7 9 1 9 0 2
39 15 13 0 9 0 2 16 13 10 9 3 0 1 9 7 9 0 2 1 10 15 15 13 1 9 10 9 0 1 11 7 11 2 11 2 11 7 11 2
22 13 9 2 1 12 2 1 10 11 1 9 13 1 9 0 2 11 11 2 11 2 2
17 10 9 0 11 13 10 9 0 1 12 7 10 9 0 1 12 2
24 13 1 12 9 0 1 12 9 0 13 15 2 10 9 1 10 9 4 13 1 9 3 0 2
19 3 1 10 9 10 9 1 9 7 9 0 13 1 10 9 1 10 9 2
30 4 13 16 15 13 1 10 9 1 9 1 10 9 16 4 13 3 2 9 2 9 2 9 2 9 2 9 7 9 2
14 3 13 0 2 0 7 13 0 10 9 1 10 9 2
50 13 10 9 1 12 9 7 13 10 9 9 1 10 9 0 7 9 2 3 1 10 9 1 10 9 7 10 9 0 2 7 1 10 9 2 9 1 10 0 9 1 9 2 9 2 9 7 9 2 2
11 11 15 13 1 13 10 9 1 10 9 2
28 11 2 12 2 7 10 9 0 2 11 2 12 2 2 9 2 3 2 1 13 3 10 9 0 1 10 9 2
21 7 2 16 3 13 2 4 13 9 0 16 13 0 9 1 9 2 2 4 13 2
15 15 13 1 10 9 1 10 9 11 1 15 1 10 11 2
28 13 3 10 9 1 13 9 1 10 9 0 1 10 9 2 10 9 1 9 7 10 9 2 1 13 1 12 2
20 1 10 9 10 0 9 1 11 1 12 9 0 13 1 10 2 11 11 2 2
20 16 10 9 0 15 13 2 15 13 1 10 9 2 2 3 13 0 7 0 2
16 11 11 4 13 3 1 10 9 3 1 10 9 1 11 11 2
25 13 1 12 9 1 9 2 12 9 1 9 0 2 12 9 1 9 1 9 7 12 9 1 9 2
8 1 0 13 12 9 1 9 2
32 3 13 7 13 10 9 1 10 9 2 15 4 13 11 2 1 10 9 1 10 9 2 11 7 10 9 1 10 9 2 11 2
17 13 10 9 0 13 1 10 9 9 9 1 10 9 0 11 11 2
11 10 9 3 4 13 1 10 9 11 11 2
35 10 9 0 1 11 11 2 1 10 0 7 10 9 1 10 9 2 15 13 1 0 9 1 9 2 16 10 9 0 4 13 10 0 9 2
20 11 11 13 0 1 10 9 1 10 9 1 11 11 9 13 9 1 10 9 2
19 4 13 1 9 7 1 13 1 10 9 2 7 1 11 1 12 4 13 2
26 10 0 2 9 2 15 15 13 1 10 9 16 15 13 0 1 9 1 10 9 7 15 13 0 9 2
61 13 10 9 1 10 0 9 1 10 9 2 11 11 2 8 8 8 8 8 8 2 3 7 1 10 9 2 11 11 2 8 8 8 7 1 10 9 1 10 11 11 11 11 2 11 11 11 11 11 2 8 8 8 8 2 8 11 8 8 8 2
19 10 9 1 10 9 4 13 1 11 11 11 7 10 9 1 11 11 11 2
14 13 10 9 1 12 9 2 11 12 2 1 12 9 2
24 3 1 3 11 15 4 13 9 1 16 13 3 3 9 1 13 1 10 9 11 7 1 11 2
20 1 9 1 12 2 10 9 1 9 4 13 1 11 11 1 10 9 11 11 2
8 16 13 1 10 9 13 15 2
14 10 9 13 0 7 3 13 10 9 1 9 3 0 2
30 11 13 10 9 7 9 0 2 1 10 9 1 11 2 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
23 10 11 13 1 10 9 10 9 1 10 9 1 11 16 15 13 1 10 9 1 10 11 2
21 13 10 9 0 0 1 10 9 2 1 9 1 10 9 7 15 0 1 10 9 2
62 7 15 2 10 10 9 13 10 9 11 7 10 9 13 16 15 13 3 2 15 13 1 10 10 9 16 13 7 3 7 13 10 9 2 1 10 9 3 15 15 0 7 10 16 13 0 1 3 10 0 9 5 2 7 1 10 12 9 15 13 0 2
41 15 15 10 10 9 13 1 0 13 16 2 13 1 9 1 9 0 1 10 9 2 10 9 16 15 13 13 10 9 1 10 9 3 7 3 15 7 15 15 13 2
25 11 11 2 11 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 13 10 9 0 2
45 13 1 9 1 13 1 11 11 11 7 13 1 9 1 12 1 11 1 12 1 9 0 2 13 11 11 1 11 2 0 1 10 11 1 10 11 1 11 2 13 9 11 11 11 2
25 10 12 2 15 13 9 1 10 9 1 10 9 0 1 11 10 11 11 2 1 10 9 1 11 2
12 16 13 1 10 9 10 9 13 1 12 5 2
50 3 13 10 9 16 15 13 1 10 9 1 10 9 2 10 9 1 16 10 9 0 15 13 9 1 10 9 13 1 12 9 1 10 9 1 10 9 7 9 7 2 1 9 2 10 9 1 10 9 2
33 10 9 0 1 10 9 13 1 9 0 1 9 7 15 13 1 10 9 16 10 9 1 10 9 1 11 13 3 10 9 1 11 2
27 10 9 15 13 16 13 10 9 1 13 10 9 1 10 9 7 10 9 1 15 16 3 13 10 9 0 2
22 10 0 9 2 3 2 15 13 1 10 9 16 3 1 9 13 10 9 11 1 11 2
30 1 9 2 1 10 11 11 1 11 12 10 9 16 3 13 10 9 4 13 10 12 5 1 10 9 1 9 1 9 2
19 13 10 9 16 13 15 1 10 3 0 7 0 9 1 9 1 10 9 2
22 10 0 9 1 11 1 10 9 0 13 1 10 9 1 11 1 10 12 1 11 12 2
23 1 10 9 1 11 2 1 10 16 13 15 1 9 2 10 9 13 0 9 1 10 9 2
31 1 10 9 0 1 10 9 1 10 9 1 10 9 1 12 2 15 13 15 1 10 9 16 13 10 9 0 1 10 9 2
84 11 3 13 0 10 9 7 9 1 10 9 0 7 1 10 9 16 13 9 1 10 9 0 1 12 2 10 9 0 7 10 9 15 13 0 1 10 9 1 10 9 1 9 2 10 9 13 3 13 1 11 1 10 9 1 11 7 1 10 9 2 7 13 13 1 10 9 0 1 11 10 9 1 10 9 13 7 9 1 10 9 1 12 2
22 2 3 3 15 13 1 10 0 9 7 3 1 10 0 9 2 0 2 0 7 0 2
42 10 1 10 11 13 10 9 1 10 11 1 11 7 10 9 3 0 2 7 10 1 10 11 11 13 3 0 7 1 9 0 2 3 11 13 10 9 3 0 7 0 2
17 11 13 10 0 7 3 4 13 10 9 2 11 3 15 13 0 2
24 10 9 2 16 15 13 1 10 9 1 0 9 2 13 3 10 0 9 16 4 13 10 9 2
31 11 11 12 11 13 3 0 1 10 9 13 1 11 2 7 10 9 13 10 0 9 13 1 10 9 7 1 10 0 9 2
15 10 9 13 3 0 2 16 13 1 11 13 1 13 15 2
19 13 15 0 7 10 9 13 1 2 15 4 13 10 9 13 15 15 2 2
34 3 16 1 11 11 3 4 13 1 10 12 2 11 13 10 9 1 13 10 9 1 11 7 11 2 16 13 1 9 1 10 11 11 2
16 11 4 13 1 2 11 11 11 11 2 10 9 1 9 0 2
20 10 9 4 13 2 1 4 13 1 9 7 13 1 10 9 1 7 15 13 2
27 10 9 1 9 1 15 1 10 9 13 10 9 1 9 0 1 9 3 0 7 0 1 13 0 9 0 2
12 13 10 11 1 10 11 1 10 11 1 11 2
15 10 12 9 13 0 9 0 7 13 9 0 1 0 9 2
12 11 11 2 10 11 2 2 9 0 7 9 2
30 3 1 10 0 9 1 9 2 10 12 1 11 2 10 11 11 13 9 1 9 0 1 9 1 10 9 1 10 11 2
32 10 9 4 13 1 9 2 10 1 3 0 9 0 1 10 11 1 12 2 15 11 13 1 10 9 1 15 1 10 9 0 2
8 2 13 1 10 9 7 3 2
24 11 4 13 1 10 9 0 2 1 15 15 3 13 3 0 16 13 1 10 9 1 10 9 2
12 10 9 1 9 13 1 12 9 2 9 5 2
30 11 13 10 9 1 16 11 13 10 9 1 13 1 11 7 2 3 1 10 9 2 15 13 10 9 1 9 1 9 2
4 2 1 15 2
25 13 3 0 9 2 12 9 2 12 9 1 9 0 7 12 9 1 9 0 2 16 13 12 9 2
21 3 7 2 10 9 1 10 9 12 1 10 9 0 4 13 15 1 10 0 9 2
51 1 9 3 4 13 7 13 10 9 1 10 9 2 15 13 1 10 12 9 9 1 10 9 2 1 13 10 9 1 10 9 1 10 9 1 11 2 13 10 9 2 10 9 11 7 10 9 2 11 11 2
25 10 9 1 10 9 2 3 13 2 13 0 1 12 9 2 13 1 9 7 1 9 13 1 9 2
4 13 9 0 2
14 1 10 9 2 10 9 11 7 11 13 1 10 9 2
29 0 9 16 13 1 11 7 11 3 13 1 16 10 9 2 0 2 13 10 9 7 3 7 16 10 9 13 0 2
31 1 13 10 0 9 0 0 2 4 13 15 10 9 1 10 9 1 10 9 0 2 9 0 1 9 2 1 10 9 0 2
12 1 10 9 2 13 12 9 7 13 12 9 2
22 10 9 13 10 9 10 9 12 2 1 10 9 1 10 9 1 9 1 10 9 0 2
17 10 9 11 7 9 13 0 9 1 10 9 0 13 1 10 9 2
16 11 11 13 10 9 1 9 1 10 9 11 1 10 9 11 2
13 15 13 10 9 1 10 9 1 9 7 10 9 2
33 4 13 7 0 2 1 15 2 1 11 2 11 2 11 2 16 3 13 9 1 10 11 11 11 7 1 10 11 11 11 11 11 2
12 13 16 10 9 4 13 0 1 10 10 9 2
10 15 13 10 9 1 15 13 10 9 2
30 13 1 10 9 1 10 9 11 7 11 7 1 10 9 11 2 3 1 10 0 9 1 11 7 11 11 2 11 2 2
28 10 9 13 13 10 0 9 0 16 13 1 10 9 1 11 2 7 3 13 1 10 11 11 3 1 10 9 2
22 1 10 12 1 11 13 10 9 1 12 9 1 12 9 1 9 2 13 12 9 0 2
8 13 1 9 7 9 1 9 2
16 13 9 0 7 1 10 9 0 13 9 1 9 0 7 9 2
11 10 9 13 0 2 3 1 12 9 2 2
92 10 11 1 10 11 11 13 10 9 15 13 10 9 0 16 13 9 1 11 1 10 9 12 2 1 10 9 1 10 11 2 1 10 9 1 10 9 16 13 10 9 1 10 9 1 10 9 2 10 0 9 1 15 9 7 13 1 10 3 13 9 0 2 16 15 13 1 10 9 0 1 3 13 9 0 1 10 9 2 1 13 15 0 1 10 9 1 9 2 12 2 2
118 10 9 13 16 2 1 10 0 9 2 10 15 13 13 1 16 15 4 13 13 2 13 10 9 16 4 13 1 11 11 12 2 10 9 3 13 2 3 13 9 1 11 11 2 1 15 11 13 3 1 10 9 1 10 9 2 7 1 10 0 9 7 10 9 11 11 2 1 15 13 1 10 9 1 13 15 15 13 2 7 3 1 10 12 1 9 15 13 1 9 1 13 1 9 2 16 13 10 9 1 10 9 1 9 0 1 11 11 2 1 10 0 11 11 2 9 2 2
15 11 13 10 0 9 1 9 1 10 9 1 10 9 0 2
57 1 15 7 10 9 2 10 0 9 11 12 2 12 2 2 13 0 9 1 13 1 15 0 2 10 9 1 11 2 11 2 15 13 1 15 1 10 0 9 1 11 2 16 13 1 10 9 1 10 9 1 11 12 11 1 12 2
46 11 11 2 9 1 10 9 2 15 13 0 1 10 9 2 7 10 9 2 9 15 13 3 7 13 10 9 2 1 10 9 16 13 10 11 2 11 1 10 10 9 7 9 3 13 2
54 13 1 11 12 2 7 13 1 10 9 0 2 16 13 10 9 11 2 10 9 13 1 11 1 9 2 7 13 10 12 1 11 1 12 10 10 9 7 9 2 13 10 9 1 10 11 0 1 11 1 10 11 2 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
49 10 9 1 10 9 1 10 11 11 2 11 11 2 3 4 13 10 9 1 11 2 0 1 10 9 1 10 11 11 1 11 1 10 11 11 2 11 11 11 2 7 10 9 1 11 2 1 15 2
62 1 9 1 10 9 2 10 9 13 2 13 1 9 1 10 10 9 2 1 10 9 7 10 9 13 10 9 2 2 1 0 9 1 10 9 2 1 10 10 9 1 13 10 9 0 3 1 10 9 0 1 10 12 5 9 1 10 11 1 10 11 2
22 10 9 2 3 4 13 16 13 0 9 0 13 1 10 9 7 10 9 1 10 9 2
25 11 13 10 9 3 0 7 10 8 2 9 13 10 9 1 10 15 10 9 13 10 9 1 9 2
14 10 9 13 3 0 2 10 9 3 0 3 7 0 2
21 13 1 11 10 11 2 11 2 2 16 13 9 1 10 0 9 1 11 1 11 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
62 10 9 15 13 16 3 2 15 15 13 1 10 3 10 9 2 2 16 13 10 9 1 10 11 1 9 1 11 2 11 11 11 2 3 7 15 13 10 9 0 1 0 9 1 11 2 12 9 1 11 7 0 9 1 11 2 3 7 10 9 0 2
42 10 9 1 12 9 1 10 9 0 1 11 15 13 3 1 10 9 0 1 11 11 2 1 10 9 1 11 2 1 16 1 10 9 15 4 13 1 9 7 9 0 2
25 16 3 13 10 9 1 16 13 10 9 0 13 1 15 16 15 13 7 13 1 10 9 1 9 2
34 1 12 13 10 9 1 10 9 0 1 9 1 10 9 1 10 11 11 11 15 13 10 9 2 7 1 10 9 0 3 13 10 9 2
55 1 10 9 1 10 0 9 2 10 0 9 2 15 1 9 2 4 13 1 9 1 9 7 9 1 10 9 13 1 10 9 2 1 10 12 9 1 10 9 1 9 2 13 1 9 2 13 1 10 9 11 11 7 11 2
46 13 1 9 10 0 9 1 9 1 9 2 1 10 10 9 9 7 9 2 15 13 16 13 10 9 1 10 16 3 13 15 13 2 16 13 7 3 3 13 9 2 7 15 15 13 2
16 10 9 4 14 2 13 1 12 8 9 1 9 7 9 0 2
7 1 12 13 1 11 11 2
21 10 9 3 1 10 9 13 16 13 10 0 9 7 10 9 13 0 2 3 0 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
30 15 13 3 0 2 13 13 2 1 10 9 2 8 2 2 16 15 13 13 15 10 9 2 3 2 2 7 3 0 2
11 3 13 10 9 1 10 9 0 1 11 2
58 10 9 13 1 10 9 1 16 2 1 9 1 0 9 2 15 13 1 13 1 11 1 9 2 7 11 3 13 7 13 10 9 1 13 1 10 9 2 1 9 13 1 10 9 1 16 10 9 4 13 9 7 13 13 1 10 9 2
13 1 10 12 9 10 9 13 7 3 1 10 9 2
21 10 9 2 7 0 2 4 3 13 1 11 2 10 9 3 15 13 3 0 2 2
23 11 13 2 2 10 9 13 9 16 15 13 1 10 9 7 16 13 3 13 0 7 0 2
20 3 13 1 10 9 1 9 2 3 13 1 9 2 9 0 7 3 1 9 2
39 10 9 13 10 0 9 1 10 9 1 9 1 10 9 2 1 10 9 1 10 9 1 11 11 1 9 1 10 9 1 9 1 11 11 7 10 11 11 2
34 3 13 10 9 13 1 10 9 1 10 11 16 13 9 1 9 0 16 11 11 13 0 2 1 10 9 0 16 3 13 11 11 11 2
20 11 11 13 10 9 1 9 1 10 9 1 10 11 1 10 9 1 10 11 2
35 10 9 1 11 2 1 9 2 11 11 2 11 11 2 2 13 1 12 2 13 15 1 10 12 9 1 10 9 0 1 11 1 10 11 2
52 1 9 1 11 2 1 12 15 13 1 11 2 3 15 13 1 10 9 1 10 9 7 1 10 9 2 7 3 1 10 1 10 9 2 13 10 9 1 10 15 15 13 10 2 0 9 2 7 0 9 2 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
42 1 10 11 1 10 11 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
58 10 9 15 13 10 9 1 13 1 10 9 1 12 9 1 10 0 9 1 0 9 11 11 2 1 9 11 11 12 2 2 12 8 8 2 12 8 1 9 8 8 2 8 7 11 2 12 9 7 9 8 2 8 12 7 9 8 2
14 13 1 9 7 10 9 0 13 10 11 1 10 11 11
13 13 0 1 9 7 13 1 0 9 1 9 0 2
24 4 13 1 13 1 10 0 9 1 15 3 1 12 9 2 7 16 13 1 10 9 2 0 2
15 11 13 10 0 9 1 10 9 1 10 9 11 1 12 2
56 10 9 1 10 9 13 0 9 2 1 10 9 13 10 9 1 10 9 1 16 13 10 9 1 10 9 2 7 1 15 1 9 1 10 9 1 10 9 2 7 10 9 1 4 1 13 10 9 7 10 9 1 10 9 0 2
44 10 9 12 1 11 1 12 2 11 11 13 10 0 9 1 10 13 15 1 10 9 1 9 2 12 9 2 2 11 1 11 11 2 9 13 1 10 9 1 11 1 10 11 2
24 10 9 1 9 13 0 1 0 9 1 9 16 2 1 10 9 2 13 10 9 1 10 9 2
34 13 9 2 1 10 0 9 2 1 2 10 9 1 9 7 9 2 2 10 11 4 13 1 10 9 1 10 0 9 7 9 1 15 2
41 3 1 10 9 0 13 9 1 16 10 11 13 1 10 9 1 13 15 1 10 9 1 10 9 2 15 4 13 10 9 1 10 11 11 7 10 9 3 13 0 2
27 10 9 0 1 10 11 11 13 10 9 1 10 9 1 11 1 12 1 13 1 10 15 1 11 1 12 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
16 3 13 9 1 11 11 0 1 10 0 9 1 11 11 11 2
23 10 9 1 11 4 13 1 10 10 9 1 10 0 9 1 10 9 0 1 10 9 12 2
27 1 10 9 13 1 10 11 11 16 15 13 1 10 9 0 1 11 1 12 1 10 9 1 13 10 9 2
13 2 10 9 13 10 9 1 13 10 9 1 11 2
42 1 12 13 10 9 0 1 10 9 11 11 7 13 3 1 10 9 1 10 9 1 11 11 7 1 10 9 1 10 9 1 12 2 9 1 10 15 4 7 13 15 2
17 10 0 9 0 3 0 1 10 9 0 1 10 9 1 11 11 2
27 10 11 11 1 11 13 10 9 0 0 1 10 9 1 11 2 16 13 1 10 12 9 16 13 10 9 2
12 4 13 3 1 9 1 10 9 0 11 11 2
40 10 0 9 1 10 9 0 7 10 9 1 9 1 10 9 0 4 13 10 11 2 11 2 11 11 11 2 11 7 11 2 12 2 7 11 2 12 2 2 2
32 10 9 4 13 9 1 10 9 1 10 9 2 1 9 1 10 9 13 1 10 11 7 1 10 9 1 10 9 9 1 11 2
64 1 10 0 9 15 13 0 9 2 13 13 2 13 10 9 7 9 1 10 9 1 10 9 2 16 1 9 2 13 10 9 9 1 10 9 1 12 9 2 2 3 7 9 2 15 13 3 10 9 13 10 9 9 3 1 10 9 7 10 15 1 0 2 2
22 10 9 13 10 9 7 9 1 10 9 16 13 13 10 12 9 1 11 10 0 9 2
26 13 15 10 9 16 13 9 0 1 10 9 2 9 2 9 2 9 2 10 9 0 2 10 9 8 2
42 16 4 7 13 1 10 0 9 1 10 9 2 11 2 2 15 3 13 1 9 1 11 2 10 9 2 7 1 10 0 9 1 9 2 11 2 2 10 9 13 9 2
18 13 1 9 7 10 9 0 13 10 11 11 1 10 9 11 11 0 2
34 15 13 1 10 11 1 10 9 0 1 11 11 2 9 2 2 11 11 2 9 2 2 11 11 2 9 2 7 11 11 2 9 2 2
18 1 3 2 10 9 0 4 13 10 9 7 10 9 2 16 13 0 2
22 11 2 8 12 2 3 1 12 2 13 10 0 9 0 1 11 11 1 10 11 11 2
30 13 10 12 1 11 1 12 2 1 10 9 1 10 9 0 7 1 10 9 0 1 11 11 2 1 10 9 11 11 2
53 10 9 0 13 3 1 10 9 1 9 0 16 13 1 10 9 2 9 2 9 7 9 1 9 0 2 9 1 10 9 1 9 8 8 1 9 0 2 7 16 13 1 10 9 11 11 11 1 0 9 1 9 2
29 9 2 9 1 10 9 16 13 9 2 1 9 1 9 2 1 11 2 13 0 9 1 11 13 1 11 10 11 2
17 3 2 10 9 0 4 13 16 3 13 13 10 9 1 10 9 2
26 15 15 13 10 2 9 0 2 1 10 11 2 7 3 0 2 12 9 1 0 7 12 1 9 2 2
14 1 10 9 1 12 2 13 12 9 13 1 10 11 2
63 3 15 13 10 9 0 1 10 11 11 1 10 11 1 10 11 1 10 11 1 10 11 7 11 2 11 2 2 11 11 2 1 10 9 1 10 0 9 1 10 9 1 10 11 11 11 2 1 10 16 4 13 12 9 0 1 10 9 9 1 11 11 2
23 1 9 2 3 15 13 10 9 1 9 7 4 13 1 0 9 1 11 11 7 11 11 2
25 15 4 13 9 1 9 7 4 13 1 13 9 1 10 9 1 10 9 13 9 1 9 1 9 2
49 15 15 13 10 9 1 9 1 9 2 1 10 9 1 10 9 16 15 13 1 10 9 2 3 7 10 9 4 13 1 10 0 9 7 1 15 15 2 10 15 13 10 0 9 15 15 13 15 2
13 10 9 1 11 13 10 9 0 1 11 2 11 2
10 13 1 10 9 10 9 1 10 9 2
20 1 3 13 10 9 1 13 3 1 3 13 1 11 1 10 9 0 3 0 2
20 15 1 10 9 13 1 10 9 13 1 10 0 11 11 7 10 9 11 11 2
31 3 1 13 12 9 3 2 13 15 15 10 9 1 10 9 1 10 11 11 4 13 7 15 13 1 10 11 2 11 11 2
35 10 9 1 11 2 11 11 2 2 13 13 2 10 9 1 10 9 1 11 11 1 11 11 2 4 13 1 9 0 1 10 0 8 9 2
30 13 0 10 9 16 15 13 1 10 9 16 7 3 3 13 1 10 9 2 13 3 10 9 11 13 1 10 9 9 2
29 10 11 11 1 11 11 11 1 12 13 3 10 9 1 9 1 10 9 1 10 9 7 1 15 10 9 1 11 2
11 10 12 1 11 10 9 13 1 10 11 2
18 10 9 11 12 13 10 11 1 11 7 10 11 11 16 13 10 9 2
12 10 9 13 1 11 1 12 1 11 1 12 2
15 13 1 10 9 1 9 1 0 2 0 2 0 7 0 2
35 1 9 2 13 16 16 11 13 3 2 4 4 13 1 10 9 1 9 1 9 2 7 13 13 16 13 3 7 16 10 9 3 15 13 2
26 3 2 13 10 0 9 1 10 9 1 10 9 7 10 9 1 10 9 0 7 1 10 9 1 9 2
62 13 0 2 7 3 0 2 13 3 1 9 1 10 9 1 10 9 1 9 2 9 2 9 1 9 2 9 2 9 1 9 2 9 1 9 7 9 1 9 7 1 9 16 13 1 10 9 1 9 1 9 13 1 9 1 9 13 1 9 1 9 2
41 1 10 9 13 10 0 9 16 13 13 1 10 12 0 9 1 10 9 2 11 11 2 8 2 2 11 2 8 2 2 11 2 8 2 7 11 11 2 12 2 2
7 10 9 3 13 10 9 2
14 13 3 0 2 16 15 13 1 11 10 9 1 9 2
28 10 9 16 13 15 7 3 13 16 13 9 13 16 10 9 13 0 7 15 0 7 15 15 13 15 3 3 2
58 10 9 13 3 0 1 10 12 9 7 3 1 10 0 9 10 9 15 4 13 1 10 9 1 11 2 12 2 2 11 11 2 12 2 7 11 11 2 12 2 2 3 7 1 10 0 10 9 0 13 10 0 7 0 1 10 12 2
19 11 13 10 9 1 0 9 7 9 16 4 13 0 9 1 10 9 0 2
15 10 12 9 0 13 11 2 11 1 11 2 11 7 11 2
38 13 16 10 9 1 10 9 13 1 9 3 7 1 9 7 13 16 10 9 13 10 9 1 15 15 13 2 10 9 1 11 11 2 7 3 10 9 2
13 10 9 13 3 0 7 3 13 13 15 1 9 2
33 1 10 9 15 13 13 10 9 1 10 0 9 2 7 13 3 0 10 9 7 13 16 15 13 15 1 11 2 16 13 10 0 2
22 10 9 13 10 9 1 0 9 1 10 9 2 1 9 1 10 9 3 0 1 9 2
10 3 13 10 9 1 11 1 10 9 2
36 1 10 9 2 10 9 4 13 1 10 9 1 10 9 1 11 1 10 11 2 7 7 10 11 2 13 1 9 9 1 10 11 1 10 11 2
25 11 13 10 9 1 10 0 9 1 3 7 13 1 11 2 1 9 1 10 9 3 1 10 9 2
52 10 9 9 11 1 11 2 1 7 3 0 9 1 9 1 10 9 1 11 2 4 13 0 9 0 7 4 13 10 9 0 9 15 13 13 9 2 13 15 1 10 9 16 3 10 9 0 4 13 10 9 2
8 3 1 10 0 9 1 9 2
56 1 15 2 11 2 16 3 15 13 1 10 0 2 4 13 3 10 10 9 2 3 16 11 2 16 13 10 9 1 9 0 2 15 13 1 9 1 9 2 2 1 15 9 3 13 10 9 3 0 1 10 9 1 9 0 2
18 13 10 9 1 10 9 1 10 9 2 3 2 16 13 1 13 0 2
25 1 13 10 9 2 13 10 9 1 9 7 10 9 1 8 1 10 15 1 10 9 1 9 0 2
36 10 9 13 16 11 11 2 10 9 16 13 1 10 9 1 12 9 1 11 2 4 13 10 9 1 9 15 13 11 7 10 9 1 10 9 2
12 11 11 11 13 1 13 10 8 2 12 11 2
20 13 1 10 9 15 13 10 9 0 16 13 15 0 2 10 9 1 10 9 2
51 10 9 4 13 16 10 2 9 0 2 1 10 9 0 15 4 13 16 13 1 10 0 9 1 10 9 0 1 10 9 2 3 7 10 9 1 9 13 1 9 13 10 9 7 1 10 9 2 4 13 2
19 1 13 1 3 2 15 13 1 10 9 7 13 10 9 1 9 1 9 2
19 3 13 2 10 9 3 13 1 9 1 13 10 9 2 13 10 9 11 2
21 11 13 10 9 1 11 10 12 1 11 1 12 2 13 10 9 0 1 10 9 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
39 10 9 1 9 2 3 13 1 9 1 9 0 2 13 10 9 13 1 10 9 1 9 1 10 12 9 16 13 16 10 9 0 4 13 1 10 9 0 2
18 4 13 1 10 11 11 11 2 10 11 11 11 7 10 11 1 11 2
13 10 9 9 4 13 1 10 9 1 10 10 9 2
27 1 9 1 16 10 9 0 13 0 1 3 1 12 9 2 13 3 0 1 10 0 9 1 9 3 0 2
28 15 13 3 1 9 1 9 2 9 7 15 13 10 9 16 13 10 9 1 0 9 16 15 13 1 9 0 2
17 13 10 9 0 2 1 9 1 0 9 1 10 9 1 10 9 2
34 2 13 9 16 1 10 9 12 3 4 13 15 1 9 2 16 3 15 15 4 1 13 2 2 13 10 9 1 2 15 13 15 2 2
29 12 9 3 1 10 9 1 10 9 2 1 12 13 3 1 10 9 1 11 2 16 3 4 13 1 10 9 11 2
21 13 11 2 11 11 1 10 9 0 2 10 9 11 11 13 9 1 10 11 11 2
20 13 9 1 11 2 10 9 13 13 1 13 10 9 1 10 9 2 12 2 2
18 1 9 1 10 9 13 10 9 16 13 10 9 2 11 1 11 2 2
15 15 13 16 10 9 0 1 11 13 1 10 3 12 9 2
29 9 0 2 0 2 0 7 1 9 0 1 8 9 1 9 0 3 0 7 1 9 0 0 1 8 5 1 9 2
14 11 13 1 10 0 11 1 13 10 9 1 10 9 2
4 11 11 11 2
26 13 16 10 0 9 0 11 11 11 2 2 11 2 2 10 9 0 7 0 2 4 13 1 10 9 2
31 1 12 10 9 1 9 1 9 16 13 10 9 1 9 0 1 9 1 10 9 11 2 11 2 3 4 13 10 9 0 2
24 0 9 2 12 9 1 10 9 1 10 9 1 10 9 16 3 2 15 11 2 13 1 11 2
26 11 15 15 13 1 10 9 2 15 16 13 10 9 1 10 0 9 1 10 11 11 2 11 1 11 2
7 10 9 13 9 0 1 11
10 9 4 13 15 1 10 9 1 11 2
36 11 13 1 9 1 11 7 11 11 13 10 9 0 1 10 9 2 7 13 16 2 10 9 1 15 15 15 10 15 13 13 15 1 0 2 2
21 1 10 9 1 10 11 15 13 10 9 1 0 9 1 10 9 0 1 10 11 2
19 10 9 13 9 9 1 12 9 0 7 10 9 0 7 9 1 10 9 2
18 13 3 1 11 2 3 13 9 1 10 9 2 11 11 11 2 11 2
24 11 11 2 11 11 11 11 2 11 2 11 2 12 1 11 1 12 2 2 13 10 9 0 2
31 10 9 13 1 10 9 0 1 11 7 10 11 2 3 7 13 9 1 9 0 2 1 15 13 1 10 9 1 10 11 2
30 1 10 0 9 16 15 13 1 10 0 9 1 11 2 11 2 16 15 1 15 15 13 1 10 9 0 1 10 9 2
37 1 10 9 1 11 1 10 9 2 11 11 13 1 10 9 1 11 13 10 9 1 10 9 0 1 10 11 7 13 1 10 0 9 1 10 9 2
19 11 7 11 13 10 0 9 1 10 11 7 2 3 2 13 10 0 9 2
11 2 13 10 9 0 1 9 1 9 0 2
21 11 11 13 1 10 9 0 1 10 9 11 2 1 11 11 0 1 10 9 0 2
20 10 11 12 4 13 1 12 2 7 13 1 10 11 12 7 10 11 11 12 2
26 3 2 4 13 1 0 9 1 9 0 16 15 13 1 12 9 0 2 15 1 10 9 1 10 9 2
14 1 12 13 10 11 1 11 1 10 0 9 0 0 2
52 1 9 1 10 9 12 2 10 11 11 1 10 11 1 11 2 3 1 10 9 0 11 11 2 10 11 2 2 13 1 10 9 1 10 0 9 2 13 10 9 0 0 1 10 9 16 15 13 1 10 9 2
27 1 10 9 10 9 0 4 1 13 0 7 10 9 1 10 9 2 1 10 9 7 10 9 2 4 13 2
65 16 10 9 2 11 2 11 2 11 11 2 2 10 9 2 7 11 2 11 11 11 2 2 10 9 2 13 1 10 9 2 13 1 10 12 9 0 2 11 2 11 11 2 2 11 2 11 11 2 7 11 2 11 11 11 2 16 13 1 13 1 10 9 0 2
20 13 10 9 1 12 9 1 15 13 12 9 7 1 3 3 4 13 10 9 2
17 10 9 15 13 3 3 1 10 0 9 1 10 9 0 1 11 2
31 16 10 9 4 13 2 7 15 3 13 1 16 15 13 9 2 1 10 9 7 1 10 9 1 13 2 13 10 9 2 2
69 10 9 11 11 15 13 10 9 1 10 9 16 13 1 10 9 1 10 11 2 11 11 11 2 13 16 13 10 9 1 10 9 15 16 3 13 10 9 1 11 1 10 9 1 10 9 11 16 2 16 15 4 13 9 7 9 1 10 9 2 13 10 9 1 10 9 0 0 2
37 10 9 2 3 7 10 9 15 1 10 9 0 13 13 13 0 1 10 0 9 13 10 9 1 10 9 1 10 9 1 13 0 2 0 7 0 2
49 10 12 1 11 2 10 9 0 1 10 11 11 11 2 13 1 10 12 5 1 10 9 2 13 16 11 4 13 1 10 12 5 1 10 9 2 7 16 11 13 10 12 5 7 11 10 12 5 2
7 15 13 0 9 1 9 2
11 1 10 9 2 10 9 13 10 12 9 2
30 15 1 10 9 1 10 9 1 10 11 4 4 13 1 12 1 11 11 11 1 4 13 1 10 9 13 1 10 9 2
28 11 13 10 9 1 9 9 0 1 12 13 7 13 1 11 11 7 13 1 11 11 2 11 11 7 11 11 2
32 1 10 9 2 10 9 11 13 1 12 10 9 1 10 9 1 10 0 9 0 2 13 1 10 9 1 10 9 1 10 9 2
8 1 9 13 3 0 7 0 2
37 4 13 0 1 10 9 0 1 9 8 2 12 7 13 1 10 9 0 10 12 1 11 1 10 12 1 10 9 1 10 9 1 11 13 12 9 2
20 15 13 1 10 9 0 1 9 2 16 15 13 3 1 10 9 1 10 9 2
16 10 0 9 1 11 15 13 1 12 2 9 1 10 15 13 2
33 1 10 9 11 2 11 7 11 15 13 10 9 1 9 1 10 9 0 2 1 13 15 13 1 9 1 9 2 7 15 13 0 2
28 10 9 4 13 1 11 11 1 2 10 0 9 1 10 9 2 2 16 13 1 10 9 1 11 7 10 9 2
15 15 13 0 1 10 10 9 16 13 1 10 9 1 9 2
25 11 11 11 13 10 0 9 0 1 10 9 1 10 9 12 7 9 1 10 12 2 0 1 9 2
50 1 11 11 15 13 16 13 10 9 1 10 0 11 11 1 11 2 1 15 15 13 16 2 13 1 10 0 9 2 13 10 9 1 10 9 16 15 15 13 1 10 0 9 1 9 1 10 9 0 2
5 11 13 10 9 2
56 9 0 1 10 11 1 11 7 11 11 1 11 2 1 12 2 7 9 0 1 2 10 11 1 11 7 11 1 11 11 2 1 10 11 11 1 10 11 2 1 10 2 11 11 8 11 2 7 1 10 11 11 1 11 11 2
12 3 13 10 9 7 1 10 9 3 15 13 2
18 11 2 3 2 4 13 3 1 11 11 2 11 11 7 11 11 11 2
18 10 9 13 3 3 7 4 13 10 9 7 3 3 13 15 16 13 2
66 1 15 1 10 0 9 1 10 11 2 2 11 2 2 2 3 1 10 9 9 12 2 2 10 9 2 2 13 1 11 13 15 1 2 9 2 2 7 13 15 0 1 16 11 11 2 9 1 10 15 13 11 2 3 13 1 10 9 1 10 11 1 10 11 11 2
19 3 4 2 13 10 9 13 1 15 1 10 9 13 1 10 9 11 2 2
16 10 9 0 13 1 10 9 1 11 1 10 9 1 11 11 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
48 1 13 15 9 1 16 15 13 1 10 9 13 1 10 9 1 13 1 10 9 1 10 13 15 1 9 2 11 13 1 9 2 2 3 15 4 13 1 13 9 2 15 4 13 1 9 2 2
28 1 10 12 10 9 1 9 0 1 10 9 13 1 5 12 2 7 10 9 9 1 10 9 13 1 5 12 2
73 15 13 1 9 1 9 2 9 2 7 9 13 1 9 7 9 7 9 1 4 3 13 1 9 1 9 2 7 3 0 2 13 1 10 9 2 1 10 9 2 2 4 13 9 1 9 1 9 1 12 9 2 1 10 9 4 13 9 2 7 10 9 13 1 9 1 9 2 9 2 9 2 8
32 15 16 4 7 13 1 9 13 16 13 0 9 16 13 3 2 3 13 15 9 13 10 9 7 13 10 8 1 10 9 2 2
32 13 1 9 2 15 13 16 11 13 12 9 1 9 1 9 1 9 0 1 10 9 12 2 9 1 10 12 9 13 1 11 2
17 11 11 4 13 1 11 11 7 10 9 11 11 1 11 7 11 2
20 10 12 1 11 1 12 2 13 9 1 10 9 1 10 9 1 9 1 11 2
30 1 10 9 13 11 11 2 11 2 11 2 10 11 2 11 7 11 1 9 1 9 7 3 16 13 1 10 9 0 2
24 3 2 4 13 1 10 9 1 11 2 9 0 13 1 10 9 13 1 10 9 0 7 0 2
21 3 2 1 0 9 0 2 11 13 10 9 1 11 1 10 12 5 1 10 9 2
13 10 9 0 1 10 11 1 11 11 1 11 2 2
24 1 15 9 1 10 9 10 9 1 11 13 1 10 9 2 1 10 10 9 2 9 7 9 2
39 10 9 1 8 1 10 9 11 11 7 15 1 9 7 9 11 2 15 1 11 2 13 1 10 9 7 9 13 16 13 10 9 2 0 2 1 10 11 2
32 10 12 1 11 1 10 9 12 2 11 4 13 1 9 1 10 9 1 9 2 3 1 11 2 9 2 11 2 11 7 11 2
21 1 10 9 1 10 11 1 10 9 15 13 10 9 13 9 1 9 0 1 11 2
38 11 13 10 9 1 11 2 1 10 7 13 10 0 9 2 1 9 1 10 9 1 9 16 13 9 10 12 1 11 1 12 2 1 10 9 11 12 2
9 10 9 1 10 9 15 4 13 2
44 13 1 9 10 9 1 9 1 10 11 1 13 10 0 9 1 11 2 7 13 9 0 1 10 9 1 10 9 0 1 10 9 2 1 10 13 10 9 11 1 11 7 11 2
24 1 10 0 9 1 10 11 11 13 10 0 9 2 15 13 3 3 1 4 13 1 10 11 2
23 10 0 9 13 3 0 1 10 9 1 10 9 0 2 3 10 9 0 13 0 13 10 9
75 10 9 4 13 1 10 9 1 10 9 11 11 11 7 11 2 11 2 12 9 1 11 2 12 9 1 11 2 12 9 1 11 1 10 11 2 12 9 1 11 2 12 9 1 11 11 2 12 9 1 11 2 12 9 1 11 2 16 13 1 11 1 11 11 1 10 11 7 11 2 1 15 10 9 2
31 10 9 15 13 1 10 9 1 9 7 13 10 9 0 1 10 9 2 10 9 2 10 9 2 10 9 7 10 9 0 2
41 1 10 9 4 13 12 9 1 9 2 12 9 1 9 1 9 2 12 9 1 9 0 2 12 9 1 11 0 2 12 9 1 9 1 9 7 12 9 1 9 2
43 1 10 9 1 10 9 1 10 11 11 2 11 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
49 13 10 9 0 1 10 9 2 13 16 13 10 0 9 2 10 3 9 7 9 2 7 3 15 1 13 12 7 12 9 2 16 13 10 9 7 13 10 9 1 10 9 2 13 10 9 11 11 2
23 10 9 1 10 9 1 9 13 1 10 9 1 10 9 1 10 9 15 13 1 10 11 2
16 1 12 1 9 2 10 9 0 1 10 9 13 10 1 9 2
23 8 8 11 8 8 2 16 13 10 11 12 2 4 13 1 11 11 1 10 9 1 11 2
11 10 9 1 11 15 13 13 1 10 9 2
11 9 0 1 10 11 2 12 2 12 9 2
24 11 11 13 1 10 11 11 1 10 9 1 11 7 10 11 2 1 10 9 1 10 11 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
19 1 10 9 2 10 9 13 12 9 0 1 10 9 0 11 8 11 11 2
17 10 9 13 9 1 9 0 2 9 0 1 10 9 1 10 9 2
44 16 10 9 4 13 10 9 2 11 11 2 10 9 1 9 2 13 13 1 11 16 15 13 1 15 16 13 10 9 1 9 1 10 9 1 11 1 13 15 10 9 0 9 2
31 1 10 9 1 11 2 11 13 1 11 7 1 11 1 10 0 9 1 10 9 1 9 16 4 13 1 11 7 1 11 2
21 7 3 10 9 3 4 4 13 3 1 10 9 0 15 13 3 1 9 1 9 2
26 2 11 2 13 10 9 0 1 10 9 1 13 1 10 9 12 1 10 9 11 11 11 11 1 11 2
17 1 9 2 13 1 9 0 1 10 12 5 1 10 9 1 11 2
33 10 9 15 13 1 12 9 1 9 2 15 1 10 9 1 10 9 2 1 10 1 10 9 7 1 10 9 3 10 9 4 13 2
8 3 2 15 3 13 10 9 2
12 3 13 13 10 9 1 13 10 9 1 11 2
22 10 9 13 9 1 11 11 2 13 1 10 9 1 10 9 0 2 9 1 11 11 2
44 10 0 9 2 10 11 1 11 2 10 11 1 10 11 2 2 10 15 4 13 1 10 12 2 15 13 3 1 12 9 7 13 3 9 1 10 9 1 9 1 10 10 9 2
28 11 11 1 10 13 15 15 13 7 15 13 1 10 9 16 13 1 10 9 1 10 9 13 15 1 10 9 2
29 3 15 13 1 10 9 0 7 13 2 1 10 9 2 10 9 1 11 11 11 11 1 11 1 10 9 1 9 2
33 10 9 1 8 4 13 9 1 13 15 2 4 13 10 9 1 12 1 12 9 7 2 1 15 2 4 13 10 12 9 1 9 2
29 10 9 13 10 11 1 11 16 13 2 13 7 13 9 16 13 9 1 9 1 10 9 7 10 9 1 10 9 2
16 10 11 3 15 13 1 3 1 12 9 1 9 2 3 2 2
39 10 9 0 13 10 9 13 2 15 13 3 1 10 9 7 10 9 0 2 1 10 0 9 1 10 9 2 13 9 2 9 1 9 0 2 9 1 9 2
60 10 9 16 13 10 9 4 13 1 10 9 0 1 10 11 2 11 11 2 7 4 13 9 1 15 2 1 15 2 11 11 11 2 11 11 2 11 11 11 2 11 11 7 10 12 0 9 13 2 11 11 11 2 12 2 7 11 11 11 2
67 1 9 2 16 11 4 13 10 9 1 10 9 1 9 16 11 3 13 2 11 15 13 10 11 1 10 9 2 1 10 9 1 16 16 10 9 13 10 9 1 9 0 2 16 4 13 15 1 10 11 10 12 1 11 2 4 13 10 9 7 3 13 15 1 10 13 2
24 3 10 9 2 16 4 13 15 1 10 9 0 2 13 15 1 10 3 13 1 10 9 0 2
11 11 11 15 13 10 12 1 11 1 12 2
21 11 13 1 13 2 7 16 11 15 13 1 15 7 1 11 2 10 9 13 13 2
37 10 11 13 13 1 10 9 1 10 9 7 16 13 3 13 8 10 9 1 11 7 11 11 2 13 9 2 10 16 3 13 13 10 9 1 11 2
50 10 9 15 13 1 12 9 1 10 9 1 10 9 1 10 11 11 2 10 15 13 10 3 0 1 10 9 2 1 10 9 10 9 11 13 12 9 1 10 11 11 1 10 9 9 1 10 9 11 2
12 10 0 9 13 16 15 13 10 9 9 0 2
26 10 9 1 9 3 13 10 0 13 10 9 16 13 3 13 10 9 16 13 7 10 9 1 9 0 2
24 1 9 1 10 11 11 11 11 4 4 13 1 0 9 2 3 16 13 9 16 13 9 0 2
30 1 11 2 11 13 16 13 3 9 1 13 15 16 15 4 13 1 10 9 2 13 10 9 1 10 9 15 4 13 2
34 10 9 0 0 1 11 11 2 0 2 11 11 11 11 2 13 10 9 13 1 10 9 1 11 11 1 10 9 0 1 11 1 11 2
24 1 16 10 9 3 13 1 9 2 11 13 1 10 9 1 10 9 1 10 9 1 10 9 2
23 3 3 4 13 10 9 1 9 1 0 9 2 9 2 1 10 9 16 13 1 10 9 2
12 13 1 10 11 11 11 1 10 9 0 0 2
22 13 3 10 9 2 13 0 2 13 16 13 15 1 13 10 9 10 9 1 10 9 2
34 10 9 0 15 13 1 10 9 11 11 11 11 2 1 11 2 15 13 16 15 13 1 12 1 10 9 0 7 1 9 1 9 0 2
15 10 9 13 1 10 9 1 15 1 10 9 2 11 11 2
18 11 7 11 13 1 10 9 2 9 1 10 9 2 16 13 10 9 2
29 1 10 9 1 11 11 13 10 12 1 11 1 12 2 10 9 1 11 13 13 10 0 9 1 13 1 10 9 2
46 10 9 1 9 11 13 9 1 10 9 1 11 11 2 7 1 13 9 10 9 13 1 13 7 16 1 9 13 9 1 10 9 1 10 9 2 15 3 15 15 4 13 1 10 9 2
34 1 10 9 1 10 12 2 1 13 1 10 0 9 1 9 0 2 10 9 0 4 4 13 9 1 9 0 0 1 13 1 10 9 2
57 2 10 9 1 16 15 13 16 13 10 9 1 11 2 13 10 9 16 3 15 4 13 2 2 13 1 10 11 11 11 2 1 12 9 2 15 1 10 9 1 10 9 11 10 11 1 11 2 10 9 1 10 9 1 10 9 2
21 15 13 10 9 0 2 1 10 9 1 9 2 15 3 4 13 1 10 11 11 2
59 10 0 9 1 11 1 10 9 1 10 9 1 10 11 15 13 13 0 9 1 13 10 9 0 1 9 3 0 7 0 2 16 13 9 1 13 1 10 0 9 0 1 10 9 1 10 9 10 12 1 11 1 12 2 1 3 12 9 2
55 3 13 0 7 13 1 10 9 2 1 10 16 15 13 10 9 2 7 10 9 0 7 10 9 1 10 9 2 1 10 9 2 13 10 9 1 9 7 1 9 1 3 13 10 9 0 1 10 9 0 1 16 13 2 2
43 3 2 1 10 9 1 0 9 2 3 1 9 11 2 13 10 9 13 1 10 13 1 11 7 13 15 1 10 9 0 2 13 10 9 0 1 10 9 1 10 9 0 2
42 7 2 13 1 10 9 1 9 10 9 11 2 13 10 9 1 2 9 1 11 2 11 2 2 11 2 9 1 10 9 11 11 11 16 13 10 16 3 13 10 9 2
26 1 9 2 13 10 9 2 16 10 9 1 10 9 16 13 0 13 3 0 7 15 13 1 13 15 2
29 11 11 11 2 3 13 1 11 2 13 10 9 0 1 9 1 11 1 9 1 11 2 1 10 9 0 1 11 2
26 1 10 9 2 10 9 13 12 9 2 7 0 2 3 10 9 16 13 12 9 13 1 10 0 9 2
12 10 9 13 0 2 9 1 10 13 7 13 2
25 1 10 9 2 1 12 2 3 1 10 9 16 4 13 3 1 12 2 13 13 10 11 11 11 2
8 13 1 10 11 11 1 11 2
28 10 0 0 9 16 13 1 10 9 3 0 2 3 3 1 10 0 9 2 7 1 10 0 9 1 10 9 2
22 4 13 15 1 9 1 9 7 4 13 3 1 9 1 11 2 9 5 12 8 2 2
32 9 1 10 9 13 1 9 0 2 13 9 1 9 7 9 1 10 9 0 2 13 1 11 1 11 1 10 9 7 11 0 2
20 10 9 0 1 10 9 1 9 13 1 9 0 3 4 13 1 10 9 12 2
12 3 2 13 0 7 13 9 1 10 9 0 2
51 11 11 13 15 1 10 9 3 0 16 4 13 1 10 9 1 9 7 3 13 9 1 10 9 0 2 1 15 15 15 15 13 10 9 0 1 10 9 1 0 9 16 3 4 13 1 10 11 1 11 2
13 3 13 2 1 9 2 1 10 9 7 10 9 2
19 12 2 1 9 1 10 0 9 2 3 13 0 13 10 9 1 9 0 2
9 10 0 9 13 11 11 1 12 2
29 10 11 11 1 11 2 11 2 15 13 1 12 1 10 9 15 10 9 1 10 9 13 1 10 9 9 11 11 2
19 10 9 13 1 10 12 5 7 10 12 5 1 10 9 0 1 10 9 2
40 10 9 2 10 9 2 10 9 0 7 10 2 9 0 2 13 1 15 2 7 13 9 1 15 10 16 3 13 10 11 7 16 3 3 13 1 15 1 9 2
41 10 9 0 1 11 11 4 13 1 9 0 2 10 9 3 1 10 2 9 1 11 2 10 12 1 11 1 12 2 16 13 15 1 10 9 13 1 11 2 11 2
28 10 12 1 11 1 12 10 11 7 10 11 11 1 11 13 10 9 11 1 10 9 1 10 9 1 0 9 2
16 10 9 13 16 10 9 1 10 9 7 1 10 9 13 0 2
15 13 13 10 9 0 4 13 7 13 1 10 9 7 9 2
17 11 13 10 9 1 10 9 13 10 9 1 11 13 1 10 9 2
12 11 13 16 11 4 4 13 16 2 13 2 2
51 12 1 10 12 13 0 1 10 11 11 2 16 13 11 2 9 0 1 10 9 11 2 2 10 11 11 2 9 1 10 9 1 10 9 11 2 7 10 11 11 2 9 1 10 9 1 10 11 11 2 2
67 10 9 13 1 10 0 9 0 10 11 11 2 3 15 13 0 10 11 1 10 9 11 2 11 11 11 2 2 3 15 13 10 9 1 9 1 10 9 1 10 9 0 2 10 11 1 10 11 1 10 11 11 2 13 1 10 11 11 7 10 11 11 1 10 11 11 2
18 10 9 13 10 9 1 10 9 15 13 10 9 1 9 1 10 11 2
7 10 9 15 13 12 9 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
49 1 13 1 10 9 11 15 13 1 11 11 13 10 9 7 10 9 13 3 13 10 9 0 1 13 10 9 3 0 1 10 9 2 16 15 13 10 11 1 10 11 2 13 15 10 11 11 11 2
15 13 10 9 16 13 1 10 9 0 2 9 0 7 0 2
16 11 11 7 11 11 13 9 1 9 7 15 15 13 10 9 2
11 1 12 10 9 4 13 2 3 2 11 2
33 1 12 2 11 13 3 3 1 10 0 9 1 11 11 7 15 13 1 15 1 10 0 9 1 11 11 2 8 2 11 11 2 2
29 3 2 1 10 9 1 10 0 9 1 11 10 9 1 9 1 10 11 3 4 13 10 9 0 1 9 1 11 2
28 1 10 9 2 7 9 1 9 2 13 9 13 1 10 9 1 10 9 2 7 11 11 13 9 1 10 9 2
23 1 10 11 13 10 0 9 1 9 2 13 10 9 2 1 13 10 9 7 13 10 8 2
38 1 9 1 10 9 0 2 10 9 3 4 13 10 9 0 1 10 9 1 10 9 1 11 2 3 13 1 10 9 1 10 0 9 1 10 9 11 2
26 3 1 16 10 11 11 15 13 1 10 11 1 10 11 1 12 2 10 9 4 13 1 10 9 0 2
16 1 10 9 12 2 3 13 1 11 10 9 0 1 10 9 2
26 0 13 10 9 7 9 16 13 1 10 9 16 13 1 10 11 2 13 13 15 7 11 15 15 13 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
20 1 10 11 13 10 9 0 1 10 9 11 2 11 2 7 11 2 11 2 2
20 13 10 9 1 10 12 9 7 1 0 13 9 0 7 13 1 13 9 0 2
12 1 9 12 13 1 10 9 1 12 12 9 2
23 1 10 9 2 3 15 13 10 9 0 1 11 2 13 16 10 9 0 13 0 1 13 2
6 3 13 10 9 0 2
19 11 13 1 12 1 11 2 13 10 9 1 12 9 1 10 9 0 0 2
16 13 9 1 11 1 11 2 1 12 1 12 9 1 10 9 2
19 10 9 16 15 13 13 3 0 7 10 9 16 13 13 3 0 7 0 2
31 10 9 1 10 9 13 1 10 9 7 9 1 10 9 2 3 3 10 9 1 10 0 11 2 11 7 10 9 1 11 2
20 10 9 4 13 10 9 1 10 9 0 11 2 1 0 9 1 10 0 9 2
43 10 9 4 0 1 10 9 16 15 13 1 10 9 1 10 9 16 13 10 11 2 3 7 1 10 9 1 10 11 11 1 11 1 11 7 10 9 0 15 13 10 9 2
11 13 1 15 12 9 1 10 10 9 0 2
11 9 0 1 10 11 11 1 11 1 11 11
23 1 9 10 9 1 10 9 0 13 10 9 1 9 0 1 11 1 13 1 10 9 0 2
10 16 15 15 13 2 15 13 1 15 2
11 2 9 0 7 11 1 9 2 9 0 2
47 10 9 2 1 9 1 10 9 2 13 1 10 2 9 11 2 7 1 10 9 1 10 9 2 16 4 13 1 10 9 16 7 3 15 13 10 12 2 5 7 13 10 9 1 11 11 2
19 11 1 11 13 10 9 1 10 9 1 11 1 10 9 1 10 9 0 2
16 1 10 11 1 11 13 9 1 9 7 0 9 0 3 0 2
13 1 9 2 10 9 0 13 10 9 1 10 9 2
18 13 10 11 2 11 1 10 11 11 1 10 0 9 0 1 10 9 2
19 13 10 9 1 10 0 9 13 1 11 11 3 1 16 11 2 11 13 2
32 10 12 1 11 1 12 2 4 13 16 11 11 15 4 4 1 13 1 10 9 2 13 0 9 0 1 9 1 11 1 12 2
36 4 13 3 1 10 9 11 2 10 9 1 10 9 11 7 11 11 2 13 3 12 9 2 10 9 11 2 10 9 0 7 1 9 10 9 2
18 10 9 13 10 9 0 1 9 12 3 1 10 9 12 1 10 9 2
22 10 9 13 10 9 1 12 1 3 9 16 15 13 1 10 9 15 4 13 7 13 2
18 11 2 1 9 11 1 11 2 13 10 9 0 1 10 9 1 11 2
14 13 9 1 9 7 9 1 10 9 1 10 0 9 2
19 1 0 9 2 15 4 13 10 9 0 2 15 16 4 13 10 9 0 2
11 10 0 9 1 9 15 13 10 9 12 2
18 10 11 1 10 11 13 10 9 0 1 11 11 1 10 11 2 11 2
29 10 9 1 10 11 11 11 13 16 10 9 1 10 9 4 2 13 2 9 0 1 10 9 1 11 2 9 2 2
18 10 9 2 1 10 9 13 1 10 9 1 11 10 9 12 1 11 2
19 10 9 13 1 9 10 3 0 9 1 9 0 1 10 9 1 11 11 2
28 10 9 16 15 13 16 13 1 9 7 9 13 0 2 10 9 13 0 7 10 9 1 10 9 7 15 13 2
50 10 9 4 13 1 13 15 1 10 9 0 2 11 2 11 7 11 2 1 9 1 9 1 9 3 16 1 11 7 1 10 9 1 10 9 3 13 10 9 1 9 16 4 13 15 9 1 10 9 2
38 10 9 11 11 11 13 1 12 10 11 1 11 1 11 7 11 11 11 2 11 2 2 1 10 9 1 13 7 13 10 9 0 7 0 1 11 11 2
31 10 9 1 10 9 15 13 1 11 16 10 9 1 10 9 13 2 15 16 13 10 9 15 10 9 7 9 15 13 0 2
20 15 4 13 1 15 9 1 12 1 10 12 0 9 1 11 1 9 1 9 2
28 10 12 1 11 1 12 2 10 9 1 10 11 4 13 3 1 15 1 10 2 12 9 0 1 10 9 2 2
79 16 15 13 10 9 15 4 13 16 10 9 9 13 1 11 2 7 10 0 12 9 1 10 9 13 15 16 3 15 13 1 11 2 10 0 9 13 1 10 11 1 10 11 1 11 2 11 11 11 2 1 10 9 1 11 2 11 2 1 10 15 2 7 1 11 1 10 9 1 11 2 11 11 11 2 1 10 9 2
28 10 9 15 13 1 9 1 10 9 13 1 10 9 2 3 1 0 9 0 2 0 13 10 9 1 9 11 2
34 1 10 9 13 10 9 0 1 10 9 0 1 10 11 11 2 11 11 2 2 1 10 9 1 10 9 11 7 15 1 10 9 11 2
17 3 1 4 13 2 15 13 7 15 13 1 11 1 11 1 12 2
29 10 11 11 13 10 9 0 13 1 11 2 11 2 11 2 1 10 9 1 10 15 3 15 13 10 11 11 11 2
19 10 9 1 9 13 3 10 9 1 16 10 9 0 8 13 10 0 9 2
23 10 9 0 1 11 11 11 9 1 10 9 0 10 12 11 11 1 10 11 1 10 11 2
48 1 10 9 2 13 9 1 16 11 3 9 1 10 11 11 2 3 1 7 10 11 11 11 13 16 9 13 3 10 9 2 15 15 4 13 16 10 9 13 10 9 1 13 1 10 9 0 2
45 10 9 0 4 13 1 12 9 2 15 1 15 13 1 10 9 0 1 10 9 1 10 11 9 1 11 7 1 10 9 0 1 9 2 3 1 10 9 0 1 10 11 9 0 2
27 1 10 9 2 11 13 1 10 9 10 0 9 2 13 1 10 9 13 10 9 1 10 9 16 13 13 2
9 4 13 1 9 2 15 13 11 2
27 1 10 11 1 10 11 7 10 9 2 10 9 1 10 9 2 8 13 1 10 9 1 10 9 7 9 2
18 13 13 3 10 9 16 13 13 10 9 7 15 13 10 9 1 9 2
27 1 11 7 10 0 9 15 13 13 0 1 10 9 1 11 2 11 13 1 10 9 2 13 1 10 9 2
59 10 9 1 11 11 11 1 10 9 0 4 13 1 10 9 13 16 10 9 11 2 11 4 13 1 9 1 10 9 1 10 16 15 4 13 10 9 1 11 1 9 1 10 9 11 11 2 7 1 10 9 0 1 10 9 1 10 9 2
24 3 3 2 10 12 1 11 1 12 15 13 1 10 9 0 1 11 1 10 9 1 11 11 2
52 10 9 4 13 10 9 1 10 15 2 3 3 1 10 0 9 2 11 13 10 9 1 11 11 2 15 13 1 10 0 9 10 9 1 10 11 11 2 16 13 10 9 0 13 1 10 9 0 2 11 8 2
15 10 0 9 13 15 16 15 13 1 9 1 10 9 8 2
38 1 10 9 13 9 1 10 9 1 10 11 2 11 2 11 7 11 3 10 9 1 10 9 1 10 9 15 13 1 9 1 10 9 1 10 9 0 2
46 16 11 2 3 2 13 13 15 1 10 12 2 4 13 15 1 11 11 3 16 15 13 1 12 9 7 13 10 0 9 2 13 15 0 2 0 7 13 10 9 1 9 7 1 9 2
50 1 9 0 15 13 13 10 0 9 1 9 0 1 10 9 2 3 15 13 9 1 9 0 2 11 11 2 11 11 2 11 11 2 1 9 1 9 9 2 11 11 2 11 11 2 11 11 11 2 2
11 3 13 16 10 9 13 10 0 7 3 2
37 1 0 9 15 13 11 11 11 2 15 1 10 9 3 0 7 0 1 10 9 2 13 10 0 11 1 11 11 7 1 10 0 12 1 10 9 2
22 3 2 11 13 1 13 12 9 1 10 9 1 13 3 1 12 1 10 12 9 0 2
14 4 13 13 10 9 1 9 9 3 1 13 1 9 2
22 1 9 1 10 9 0 1 10 9 2 10 9 13 1 10 9 1 9 1 10 9 2
36 1 15 1 10 9 1 10 0 9 2 16 3 4 13 2 13 10 9 7 10 9 13 1 9 13 1 9 1 9 2 0 1 9 7 9 2
14 11 11 11 13 10 9 0 10 9 9 1 10 9 2
10 1 9 13 16 10 9 0 13 0 2
9 3 4 7 13 16 4 13 9 2
13 1 9 15 13 10 9 1 9 7 15 13 13 2
13 1 15 4 13 10 9 1 10 9 1 10 11 2
23 10 11 1 10 11 13 10 9 1 11 1 10 11 2 16 15 13 1 10 9 1 11 2
29 10 9 1 10 11 1 10 11 1 11 13 10 9 2 13 15 1 15 9 2 1 10 0 9 1 9 11 11 2
45 10 9 1 11 13 10 9 1 9 3 10 9 0 9 1 10 9 0 3 13 13 10 9 0 0 15 16 13 1 10 9 1 9 3 3 0 7 10 9 0 1 10 12 5 2
10 1 12 2 4 13 1 9 1 9 2
24 11 4 1 13 10 9 1 10 9 2 13 1 9 1 11 11 2 11 11 2 11 7 11 2
19 1 10 9 2 10 9 13 1 10 9 1 12 9 0 1 10 9 0 2
26 3 10 12 1 11 1 12 2 13 0 9 1 10 11 11 11 1 11 2 11 4 13 9 1 11 2
30 1 10 11 1 10 11 1 12 10 9 0 1 9 1 10 9 13 1 5 12 7 10 9 0 1 9 13 5 12 2
15 3 2 10 11 13 10 9 1 10 9 1 10 9 11 2
16 3 2 1 12 1 12 13 10 9 3 0 2 15 1 9 2
33 7 15 4 13 10 9 1 10 9 11 16 4 13 2 15 5 13 7 10 9 11 13 3 13 1 10 9 1 10 13 10 9 2
13 10 11 4 13 1 11 2 7 4 13 10 9 2
22 10 9 15 13 1 9 1 9 1 9 9 2 7 13 9 2 9 1 9 7 9 2
16 10 9 2 13 3 1 9 0 2 3 13 9 7 9 0 2
29 10 2 11 11 13 10 9 1 10 9 0 1 10 9 12 3 1 10 9 1 11 1 10 9 0 1 11 11 2
12 11 4 13 10 9 2 11 1 10 11 2 2
48 1 9 2 10 9 1 9 1 10 9 0 4 13 3 7 1 10 9 2 1 10 9 1 10 2 9 2 2 10 15 15 13 1 10 9 1 9 1 10 9 1 9 1 3 1 10 9 2
23 10 0 9 4 13 1 11 11 7 13 1 11 2 11 7 1 10 11 2 13 15 8 2
26 10 9 1 10 9 4 13 1 10 9 2 9 2 9 1 11 11 11 12 10 12 1 11 1 12 2
37 10 11 2 9 1 11 11 11 11 2 11 11 1 11 1 11 2 2 13 10 9 13 13 9 1 10 9 1 9 11 1 10 9 1 12 9 2
19 3 13 13 3 12 9 1 9 1 10 9 16 3 3 4 13 9 0 2
34 3 13 0 1 10 9 1 10 11 15 13 11 2 16 10 9 13 0 10 9 1 9 1 10 9 1 10 9 1 10 11 1 11 2
31 10 0 9 13 10 1 10 9 13 1 11 11 11 7 11 11 2 13 10 12 1 11 1 12 2 1 11 12 1 11 2
21 7 16 10 9 13 10 3 0 2 13 10 1 9 0 2 10 9 3 13 0 2
32 10 9 1 10 9 12 2 13 10 9 1 12 9 1 10 9 1 12 9 5 2 1 10 9 0 1 12 9 1 9 5 2
14 13 10 9 7 13 9 2 15 13 10 9 1 9 2
38 3 1 10 9 0 13 10 0 9 1 9 0 2 1 10 0 9 1 9 2 7 9 1 9 0 13 1 10 9 1 10 9 1 10 9 15 13 2
39 11 13 1 11 11 11 2 9 0 1 9 2 9 2 1 10 9 15 13 11 11 1 11 2 2 3 1 11 11 1 11 2 10 9 1 10 9 11 2
34 1 10 9 0 2 13 10 9 0 0 1 10 9 1 11 2 1 10 9 13 10 9 1 10 9 7 1 10 11 1 10 11 11 2
13 2 10 9 4 13 13 10 12 5 1 9 0 2
39 11 13 10 9 0 7 10 9 2 10 0 9 2 2 9 0 0 2 9 0 1 11 2 13 10 9 0 2 10 9 7 9 9 7 12 9 1 9 2
55 11 11 11 2 11 2 12 1 11 1 12 2 12 1 11 1 12 2 2 1 9 11 7 11 2 13 15 1 10 9 0 3 0 2 3 1 4 13 10 9 0 1 11 2 10 8 8 8 2 9 1 10 9 2 2
20 13 10 9 13 1 10 9 2 11 13 10 9 1 9 2 13 13 1 11 2
21 13 10 9 1 12 9 7 3 15 13 7 10 2 11 2 15 15 13 1 9 2
22 10 0 9 15 13 1 15 9 1 10 12 9 1 9 2 1 10 9 1 0 9 2
12 10 9 16 13 13 0 7 10 9 13 0 2
62 9 1 0 9 0 1 10 9 1 10 11 0 1 10 9 11 11 11 7 1 10 9 1 10 9 0 1 10 9 0 2 11 11 13 1 10 9 1 10 9 0 1 11 11 1 10 9 1 10 9 0 1 10 9 1 11 7 10 9 1 11 2
21 3 9 16 13 10 9 1 0 9 0 16 13 10 9 1 10 11 1 10 12 2
18 10 9 0 0 2 13 10 11 11 11 2 15 13 1 12 1 12 2
6 15 13 16 13 15 2
18 1 12 4 13 1 11 11 2 3 1 13 15 1 11 12 9 3 2
18 16 15 13 1 11 11 2 15 13 1 11 1 13 10 9 1 9 2
20 10 9 4 13 1 10 9 1 11 7 13 1 10 9 1 10 9 13 3 2
27 1 15 1 10 9 2 10 9 1 13 15 1 9 2 10 9 2 9 7 9 1 10 9 13 13 15 2
20 3 13 9 1 10 11 1 9 0 2 15 4 13 1 0 9 1 10 11 2
29 13 10 9 15 13 1 0 9 10 9 1 10 9 1 12 9 0 2 1 10 9 11 11 2 11 2 12 2 2
14 13 16 15 13 16 1 0 9 13 3 1 12 9 2
42 3 13 16 13 10 9 0 2 3 13 16 13 0 1 4 13 15 16 13 1 13 2 2 13 11 2 3 13 1 11 2 16 15 13 10 9 1 10 9 1 9 2
14 1 12 15 13 1 11 16 13 1 10 11 11 12 2
14 10 9 15 15 13 7 15 15 13 16 3 15 13 2
22 4 13 2 10 9 2 1 15 1 10 0 9 1 10 9 0 1 10 11 11 11 2
16 11 13 10 9 0 1 9 1 9 1 10 9 1 10 11 2
24 1 10 9 15 13 10 9 9 2 3 7 9 1 9 7 9 16 13 1 13 9 7 9 2
9 15 13 1 10 9 7 15 13 2
16 11 11 1 11 2 11 2 12 2 11 2 11 2 12 2 2
16 10 9 11 13 15 1 10 12 9 0 1 10 11 1 11 2
22 1 13 15 15 2 15 13 10 11 1 10 9 2 15 16 13 16 15 4 13 0 2
52 10 9 0 4 13 2 3 16 10 9 0 13 1 13 15 1 16 15 16 13 15 13 3 1 10 9 1 9 2 3 3 1 9 1 10 9 1 9 7 9 0 2 7 3 1 10 9 0 7 0 0 2
20 10 9 15 13 10 9 2 10 9 2 9 2 9 1 13 7 10 0 9 2
15 13 13 10 9 1 10 9 2 2 15 13 1 10 9 2
43 16 10 9 0 0 15 13 9 1 10 9 7 10 9 1 10 9 13 3 15 3 2 3 16 1 13 1 12 2 12 2 10 9 13 3 10 9 13 1 10 9 0 2
14 11 13 10 9 7 13 3 10 9 1 9 1 9 2
16 1 10 9 13 1 9 1 9 1 10 9 7 1 10 9 2
17 13 1 12 2 3 13 1 10 11 1 11 11 7 4 13 3 2
38 10 9 1 9 13 1 10 9 1 10 10 9 1 11 3 4 13 1 10 9 1 11 2 15 3 13 10 9 1 9 2 5 2 7 2 5 2 2
17 11 4 7 13 15 1 10 9 10 9 1 10 9 7 13 15 2
20 10 9 0 13 1 9 1 9 0 7 9 0 1 13 2 13 7 13 15 2
14 10 9 15 13 11 11 7 13 1 10 8 11 11 2
23 13 10 9 1 10 9 1 10 0 9 1 11 1 11 7 11 1 11 1 11 7 11 2
4 13 1 11 2
36 1 12 2 11 13 10 2 11 11 11 2 13 1 12 9 1 10 11 11 2 1 9 1 10 9 1 9 1 10 9 2 11 8 11 2 2
17 3 1 10 9 10 9 13 15 0 2 3 7 13 3 15 13 2
17 16 13 15 3 1 10 9 3 15 13 7 4 1 13 1 15 2
16 1 10 15 16 13 10 9 0 1 11 2 3 15 15 13 2
26 1 12 4 13 1 11 2 11 11 2 1 13 10 9 1 10 9 0 13 1 13 10 9 1 11 2
33 10 9 15 12 11 11 11 11 11 11 11 1 10 11 13 1 10 9 2 13 16 2 10 9 13 1 10 9 3 1 11 2 2
13 12 9 3 3 13 10 11 1 12 9 13 11 2
25 1 10 9 1 10 9 2 1 11 11 2 3 15 13 1 9 10 9 1 10 9 13 1 11 2
27 1 10 9 2 3 10 9 1 9 13 1 0 9 2 7 16 10 9 1 9 3 13 2 1 9 2 2
27 9 0 13 10 0 9 1 9 1 9 0 7 0 2 7 10 9 1 11 4 3 13 1 13 10 9 2
12 13 10 9 3 0 7 0 16 13 10 9 2
11 10 0 9 1 4 13 13 10 9 0 2
21 15 13 1 10 9 2 11 2 1 11 2 0 1 10 9 2 11 2 1 11 2
21 13 13 15 1 10 9 1 11 11 2 11 11 7 10 9 1 0 9 3 13 2
32 11 11 11 2 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 13 10 9 7 9 0 1 11 2 11 2 2
36 11 2 11 2 1 2 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 11 2 1 10 9 1 11 7 9 1 11 2
24 1 10 11 11 13 3 0 2 13 15 1 10 9 9 0 10 9 12 1 10 9 1 11 2
24 10 11 2 9 10 9 0 4 13 11 2 13 1 16 11 13 10 9 1 11 13 1 11 2
8 2 15 13 10 0 9 0 2
39 10 9 0 7 8 9 15 13 1 10 9 16 13 10 9 1 9 1 13 10 9 2 13 1 10 9 2 1 7 15 13 10 9 1 10 9 1 9 2
40 11 11 2 11 11 2 1 9 2 2 13 10 0 9 13 1 10 9 1 11 11 7 10 11 7 1 10 9 1 10 9 1 10 11 2 1 10 11 11 2
22 10 11 4 1 13 1 10 11 16 3 4 13 1 10 9 16 13 10 0 9 0 2
15 16 4 3 13 1 10 9 13 3 0 1 10 10 9 2
12 11 3 13 1 9 2 7 13 1 12 9 2
25 15 3 13 10 9 0 1 10 9 2 13 10 9 2 7 3 13 0 16 3 13 1 12 9 2
35 13 1 11 2 1 3 12 9 2 4 13 1 10 9 1 10 11 11 2 1 12 9 1 10 9 2 13 1 10 9 0 1 10 11 2
17 10 9 13 11 2 16 15 13 1 10 9 0 1 10 0 9 2
8 11 15 13 0 1 10 9 2
18 11 2 10 9 1 11 13 1 13 10 9 1 10 11 11 1 11 2
20 1 10 9 1 10 0 9 10 9 15 13 1 9 0 1 10 9 1 11 2
25 3 13 9 13 16 10 11 15 13 1 10 9 1 0 9 2 3 0 7 1 0 9 1 9 2
34 15 13 1 10 0 9 9 1 10 9 16 13 10 11 7 16 15 13 13 1 10 9 1 10 11 11 2 1 11 7 1 10 11 2
26 11 11 13 10 9 2 0 1 10 9 0 1 10 11 2 9 1 11 2 16 13 12 9 1 9 2
17 10 9 1 9 1 10 9 0 1 9 13 1 12 7 12 9 2
20 1 10 15 15 13 10 9 0 13 1 10 9 2 13 1 10 9 7 9 2
27 10 9 13 7 13 2 10 9 15 13 1 10 11 11 11 2 16 13 10 10 9 3 13 1 10 9 2
12 11 11 13 10 9 1 9 1 10 9 11 2
8 13 10 9 1 10 9 12 2
26 3 13 10 9 12 1 11 11 2 10 9 12 1 10 11 11 7 9 11 1 11 7 12 1 11 2
18 15 1 10 9 15 13 2 1 10 9 2 16 13 0 1 13 15 2
17 13 10 9 0 16 13 2 15 13 1 9 13 12 9 1 9 2
15 11 2 12 1 11 1 12 2 12 1 11 1 12 2 2
40 11 11 13 1 12 7 2 1 13 1 10 9 2 11 1 11 13 10 9 1 10 9 16 13 1 10 9 12 9 1 10 9 0 7 1 9 1 10 9 2
33 11 11 1 11 2 9 0 1 9 2 13 1 11 1 13 15 1 10 9 11 11 7 1 10 9 1 10 11 11 2 11 11 2
45 10 9 1 10 9 13 2 0 9 2 8 8 2 12 2 2 11 1 10 9 2 8 8 8 2 12 2 7 9 0 2 8 8 8 8 8 2 12 2 2 15 1 11 11 2
36 11 15 13 1 10 9 1 11 2 7 2 1 9 1 16 11 15 4 13 13 1 9 10 9 2 3 13 0 1 13 1 11 1 10 9 2
29 10 11 11 13 1 10 9 10 9 1 9 1 11 11 16 4 13 10 9 3 3 16 13 13 1 10 9 0 2
12 10 9 4 13 1 10 9 1 9 11 11 2
43 10 9 1 10 9 3 4 13 3 0 2 13 1 9 1 10 0 9 2 13 8 0 9 1 10 9 2 1 12 9 1 9 2 7 10 0 0 9 2 1 12 9 2
45 10 9 0 3 4 13 15 1 13 15 3 2 15 15 13 7 13 16 10 11 0 1 11 11 1 9 1 11 2 9 1 10 11 2 2 15 13 9 0 7 15 13 10 9 2
29 1 0 7 10 9 1 10 9 1 11 11 2 2 11 2 11 11 2 13 10 9 7 10 9 13 1 12 9 2
16 2 11 2 13 10 0 0 1 10 9 1 9 0 0 11 2
23 10 9 2 13 1 10 9 2 10 9 0 11 7 10 9 11 2 16 3 3 13 2 2
18 11 3 13 10 9 2 16 13 0 15 13 16 15 13 1 10 9 2
47 15 13 10 9 1 10 9 7 16 3 13 10 9 3 0 2 13 1 10 9 16 13 1 10 9 1 10 9 2 3 3 0 10 9 2 16 3 13 0 1 10 9 2 7 10 9 2
19 10 9 4 13 1 11 11 7 13 1 11 11 12 2 1 10 9 12 2
30 1 12 15 13 1 10 9 0 1 11 2 11 2 2 16 13 3 1 12 1 10 9 0 2 4 13 9 1 11 2
6 13 12 9 1 9 2
47 1 12 13 10 9 1 9 1 10 9 2 11 11 2 2 11 11 13 10 9 1 10 9 1 10 9 11 11 2 3 16 13 10 0 9 1 10 9 2 2 7 13 10 0 9 0 2
14 1 9 13 10 9 1 9 7 9 0 16 13 0 2
5 9 9 1 11 2
11 13 10 9 16 13 10 12 9 1 15 2
11 11 13 3 10 9 0 1 10 9 0 2
28 3 15 13 10 9 1 11 11 2 10 11 11 2 11 11 11 2 11 11 11 7 10 12 0 1 10 9 2
14 1 10 9 1 12 2 13 12 9 13 1 11 11 2
25 13 10 9 13 1 10 9 1 10 9 1 9 7 10 9 1 10 9 1 10 9 0 13 0 2
30 11 11 11 11 2 13 1 11 1 12 2 13 10 9 1 10 9 7 1 10 9 2 9 1 10 9 12 7 12 2
25 1 9 2 10 9 13 16 15 4 13 10 9 13 1 13 1 10 10 9 2 2 8 8 8 2
17 13 10 9 1 10 10 9 2 16 16 13 12 9 3 13 12 2
5 11 13 12 9 2
25 10 9 13 3 0 2 10 9 2 10 9 1 10 9 2 10 9 0 2 7 15 9 10 9 2
28 11 11 11 2 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 10 9 2 9 7 9 0 0 2
24 11 11 2 1 11 11 13 16 10 9 1 10 9 1 9 15 13 1 10 9 1 9 0 2
37 1 10 9 13 3 9 1 10 9 1 10 11 11 1 11 2 4 13 1 10 9 1 9 1 10 11 11 11 2 9 16 13 1 11 1 12 2
16 1 9 1 15 11 13 10 9 1 10 9 16 13 1 9 2
54 10 0 9 2 13 1 12 7 13 10 11 1 10 11 2 13 10 0 9 1 10 9 0 2 7 13 1 10 9 10 9 1 13 9 1 10 9 0 7 0 16 13 13 10 9 7 13 1 13 10 9 3 0 2
9 10 9 13 9 0 13 1 9 2
17 1 9 13 10 0 9 0 1 9 2 10 11 11 2 9 2 2
14 10 9 1 9 13 15 16 13 2 3 13 3 0 2
62 1 10 12 9 2 10 9 1 11 13 0 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
4 13 1 11 2
32 10 9 1 10 9 0 1 10 9 13 10 11 1 15 11 1 11 2 10 11 1 10 11 1 11 7 10 11 11 1 11 2
28 1 10 11 1 10 11 2 10 9 13 10 9 0 1 2 1 10 15 13 9 7 2 12 5 2 13 9 2
65 16 11 4 13 10 9 0 1 10 9 0 1 12 7 12 7 3 13 10 9 0 1 9 7 9 2 10 12 0 9 1 10 9 11 11 13 1 10 9 1 10 9 1 10 9 1 10 2 9 0 2 16 13 10 0 9 1 1 13 10 9 0 1 11 2
10 10 9 4 4 13 1 10 9 0 2
20 1 9 1 9 1 10 9 15 13 10 9 1 9 1 10 9 1 11 11 2
22 9 2 16 3 15 13 10 9 2 10 9 13 1 10 9 13 9 1 15 3 0 2
13 15 16 13 1 11 1 9 13 15 16 15 13 2
38 10 9 1 9 1 9 1 9 2 13 10 9 9 7 13 0 2 10 9 2 10 9 2 10 9 2 10 9 7 3 10 9 1 10 9 13 0 2
45 13 1 10 9 13 1 10 9 0 2 10 9 1 11 13 10 3 0 1 11 3 1 10 9 7 1 15 15 13 0 1 13 1 9 10 9 0 1 10 9 1 9 1 3 2
26 7 13 10 0 9 15 10 9 13 13 2 7 13 13 1 10 9 16 13 10 9 2 11 11 2 2
27 1 9 1 12 4 13 1 13 1 11 1 9 1 16 4 13 10 9 1 9 1 9 13 1 10 9 2
36 1 10 0 9 10 11 11 1 10 11 7 10 9 2 3 11 1 11 1 10 11 11 11 2 4 1 13 15 1 10 11 11 1 11 11 2
21 3 13 10 9 16 15 13 1 12 9 1 10 9 1 11 7 13 10 9 0 2
23 1 8 2 9 2 4 13 10 11 11 11 11 7 2 9 0 2 10 11 11 10 11 2
21 10 9 1 9 13 11 11 11 1 11 2 9 1 11 1 11 2 11 1 11 2
25 1 11 1 12 2 11 13 10 9 1 13 15 1 12 9 0 13 10 9 1 11 1 10 9 2
16 11 13 1 10 9 1 13 1 10 9 0 10 9 1 11 2
16 10 9 0 13 10 9 0 1 10 9 1 9 1 9 0 2
36 10 9 1 10 9 1 11 15 13 10 12 1 11 1 12 2 16 13 3 16 13 1 11 1 11 11 1 10 0 9 1 10 9 1 11 2
53 11 2 13 1 10 9 16 13 1 11 11 2 7 13 16 11 4 13 10 9 0 2 13 13 1 11 1 13 10 9 2 1 13 15 15 1 11 11 15 15 4 13 13 15 1 13 10 9 1 11 7 15 2
16 13 10 10 9 16 13 16 13 7 13 10 9 1 10 9 2
28 11 11 12 13 1 10 12 1 10 9 1 10 12 1 10 9 2 13 9 1 10 9 11 2 1 9 0 2
6 13 3 0 1 12 2
23 1 9 2 10 9 4 13 10 9 13 15 1 10 9 3 0 2 1 9 7 9 2 2
10 13 10 9 1 10 9 1 10 9 2
19 10 9 1 11 11 13 12 9 1 11 2 12 1 11 7 12 1 11 2
36 1 13 10 9 1 10 9 1 10 9 0 2 0 1 10 11 11 1 11 2 11 7 11 2 11 11 11 2 15 13 1 10 9 1 11 2
18 7 4 1 13 15 9 2 1 12 9 1 9 1 12 8 10 15 2
28 10 9 13 10 9 1 13 9 16 4 13 0 1 10 9 1 8 2 15 16 4 13 10 9 1 10 9 2
27 15 13 10 11 1 0 9 1 10 12 1 10 9 13 1 10 9 1 12 8 1 11 2 11 11 2 2
37 1 12 15 13 2 1 10 9 1 10 9 11 10 11 2 10 9 1 10 9 2 13 10 9 0 1 1 10 9 2 1 10 9 1 10 11 2
33 3 15 4 13 7 10 13 10 9 0 13 1 16 10 9 15 13 1 9 2 7 5 13 9 1 10 9 13 16 13 10 9 2
23 13 13 1 10 9 1 10 9 1 12 2 12 9 2 1 11 2 11 2 11 7 11 2
11 13 9 1 16 13 0 9 1 10 11 2
36 1 10 9 16 13 10 9 2 15 13 10 0 9 1 10 9 2 10 9 1 13 9 1 10 9 0 7 10 9 16 13 1 9 1 9 2
18 13 1 9 1 10 9 1 9 0 2 13 1 10 9 0 1 11 2
17 0 9 0 7 0 4 13 1 11 16 13 9 13 1 10 9 2
18 1 10 9 16 13 1 15 15 1 10 0 9 7 9 1 10 9 2
23 11 11 11 13 10 9 1 9 0 1 9 0 1 13 10 9 0 7 0 1 10 11 2
31 10 9 1 9 0 2 11 11 2 13 10 9 1 9 13 15 1 10 9 11 16 13 10 9 0 1 10 15 1 11 2
20 10 9 16 15 4 13 4 13 0 7 10 9 1 10 9 0 13 3 0 2
22 13 1 10 9 2 7 1 4 13 1 10 9 13 1 10 9 1 9 1 9 0 2
32 1 13 1 10 9 12 2 13 10 9 1 9 1 9 7 9 2 3 1 10 9 1 2 10 11 2 7 2 10 11 2 2
17 1 9 1 10 9 13 1 10 11 11 1 10 9 11 1 11 2
28 10 11 1 10 11 15 13 1 10 9 7 10 9 1 9 1 10 9 1 9 1 10 9 9 1 10 9 2
9 3 13 9 15 0 1 10 9 2
27 11 11 2 3 13 1 9 0 2 13 10 9 1 10 9 11 1 10 9 0 2 13 1 10 9 11 2
17 10 9 0 13 11 11 2 1 9 2 7 11 11 2 1 9 2
59 10 9 1 10 9 1 10 9 0 2 11 11 2 13 16 10 9 4 13 9 0 1 9 7 16 1 15 13 1 2 0 9 16 10 9 7 9 13 10 9 0 3 15 13 10 9 1 8 13 13 9 2 9 2 9 7 9 2 2
32 10 9 3 15 13 10 9 0 13 10 11 11 2 11 7 11 2 16 16 15 13 1 13 10 9 0 2 1 11 7 11 2
49 1 10 12 9 13 16 13 10 9 1 10 9 7 13 2 15 13 16 3 13 0 2 16 15 4 13 10 9 7 16 15 4 13 2 13 10 10 9 7 15 13 1 13 10 9 1 10 9 2
13 3 2 1 0 9 2 10 9 13 9 1 11 2
30 11 2 11 13 9 0 1 10 0 9 1 11 1 9 1 10 9 0 2 1 16 15 13 9 1 10 11 1 11 2
7 13 0 1 10 11 0 2
50 10 9 1 9 13 0 9 3 13 1 3 1 10 9 1 13 2 4 13 10 9 1 9 2 2 1 10 0 9 2 1 10 0 9 2 1 10 9 9 2 9 2 3 4 13 9 1 9 0 2
33 1 9 1 11 15 13 15 1 10 0 9 13 11 2 10 9 1 10 0 9 2 9 2 1 10 11 11 1 3 1 12 5 2
45 1 9 3 1 9 0 2 3 13 1 10 9 1 12 9 2 2 13 10 9 1 9 2 13 9 2 13 9 0 2 13 1 10 9 0 7 4 1 13 1 10 9 10 9 2
23 13 16 4 13 16 15 13 5 12 1 10 9 16 3 13 3 7 13 1 9 10 9 2
16 11 13 10 9 1 9 1 10 9 11 13 1 9 1 12 2
18 1 12 2 11 11 13 10 0 9 13 2 11 1 10 11 11 2 2
58 1 9 2 10 9 16 13 10 0 9 1 9 13 1 12 2 15 16 3 13 10 9 0 2 13 1 9 1 10 0 9 1 10 9 7 1 10 9 2 15 3 4 13 1 9 1 9 7 9 1 10 9 3 0 1 11 11 2
27 10 9 4 13 3 1 10 11 11 10 12 1 11 1 12 1 11 11 11 7 3 3 13 10 0 9 2
31 10 11 0 1 10 9 1 9 1 12 2 16 11 13 1 10 9 4 13 1 10 0 1 9 0 9 1 9 11 11 2
25 10 11 13 10 9 1 9 1 10 11 2 16 1 3 13 4 13 1 10 0 9 2 11 11 2
77 1 10 9 2 11 11 2 1 12 10 9 13 1 9 1 13 15 1 9 7 9 1 16 2 1 10 9 1 9 2 15 13 10 9 1 10 9 0 1 10 15 10 9 4 13 16 13 10 9 7 10 9 2 1 10 9 1 16 16 15 13 1 10 9 2 10 9 1 10 9 0 0 4 4 0 9 2
54 13 0 2 16 16 15 13 16 1 10 9 0 10 9 1 10 9 1 15 1 10 9 13 10 9 1 10 15 2 13 16 10 9 7 10 9 13 1 10 0 9 7 3 13 0 16 10 9 13 9 1 10 15 2
22 10 9 4 13 3 1 11 11 11 2 1 9 1 10 9 11 2 3 1 11 11 2
23 1 9 12 2 4 13 3 1 12 9 7 13 1 13 10 9 1 9 1 9 1 9 2
53 10 9 15 13 1 10 9 0 1 10 9 11 11 2 10 9 1 11 7 9 1 10 9 15 4 1 13 10 9 2 10 9 13 1 10 9 1 10 9 16 13 10 9 0 1 10 9 7 1 10 9 0 2
15 1 12 2 10 9 1 10 11 13 15 1 15 3 0 2
15 3 13 13 10 9 1 10 11 11 11 1 10 11 11 2
20 1 10 9 15 13 10 9 11 11 7 11 11 2 7 13 10 9 0 0 2
32 11 13 16 10 9 13 0 2 15 3 15 4 13 7 16 11 3 15 4 13 1 10 0 1 10 0 9 7 10 0 9 2
21 4 13 1 0 12 9 3 3 2 3 1 4 4 13 1 9 16 13 10 9 2
11 15 13 10 9 0 16 15 13 1 12 2
19 1 10 9 12 2 1 10 11 12 15 15 13 10 2 9 2 3 0 2
50 1 15 16 11 13 10 2 9 2 2 13 16 10 9 13 9 7 13 1 9 0 2 16 13 10 9 1 13 10 0 9 16 15 13 3 1 11 7 11 2 3 7 1 9 2 1 11 7 11 2
46 16 13 10 9 1 9 1 10 9 3 13 10 9 1 9 16 13 2 10 9 13 3 0 7 15 13 2 3 1 10 9 1 10 9 16 3 13 3 9 7 3 15 15 13 13 2
15 9 11 11 10 9 0 13 11 11 11 1 10 11 11 2
11 3 3 10 9 13 3 1 10 9 0 2
20 1 12 13 10 0 9 1 10 9 0 16 13 10 9 1 2 9 0 2 2
9 11 11 13 1 10 9 0 11 2
28 1 10 9 2 11 11 11 2 12 2 13 1 10 9 2 7 4 13 1 11 2 11 1 13 10 0 9 2
12 10 9 1 12 15 13 1 11 2 11 2 2
24 11 7 10 9 1 10 9 15 13 9 1 10 9 7 13 10 0 9 7 11 7 10 9 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
46 1 12 2 1 10 9 0 1 11 2 10 9 13 10 9 1 12 8 12 2 1 10 9 5 12 9 2 1 15 15 10 9 0 1 9 1 10 9 1 3 1 5 12 12 9 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
8 11 11 13 1 11 2 11 2
18 3 13 1 10 9 11 1 12 2 3 13 10 9 16 13 9 0 2
16 10 9 4 13 1 10 9 0 16 15 13 1 9 1 11 2
10 13 1 10 9 0 1 10 11 11 2
24 1 10 9 1 9 1 10 9 15 13 10 9 1 10 11 11 1 10 15 13 10 0 9 2
30 1 10 9 12 2 13 1 10 9 1 9 0 1 9 0 2 11 11 11 2 10 9 1 10 0 9 1 10 9 2
62 2 10 9 13 2 1 10 9 1 9 2 10 9 3 0 1 13 1 9 2 13 2 3 1 13 16 2 1 10 9 2 13 10 9 1 10 8 2 1 10 9 1 11 2 16 13 10 9 1 9 2 0 2 2 13 2 3 0 7 0 2 2
18 11 13 1 13 1 11 16 3 13 15 15 15 13 2 7 11 13 2
20 3 3 13 11 8 2 10 9 16 13 10 0 9 1 11 2 10 8 9 2
22 3 15 13 16 10 9 13 1 10 9 2 13 1 10 9 7 13 9 1 10 9 2
13 13 10 9 7 9 1 0 9 13 1 12 9 2
18 11 13 1 13 16 13 1 10 9 7 4 13 10 0 9 1 3 2
13 11 11 13 10 9 0 13 1 10 9 1 11 2
18 13 1 12 16 10 9 1 10 9 13 13 10 0 9 1 0 9 2
8 10 9 13 15 9 1 15 2
21 9 1 11 3 13 10 9 16 15 13 2 7 4 13 10 9 16 15 4 13 2
22 10 11 1 10 11 11 2 1 9 2 8 8 2 13 15 1 10 12 9 1 11 2
77 11 11 11 3 13 1 11 11 2 12 1 11 1 12 1 11 1 11 2 11 2 2 13 10 9 7 9 0 1 9 0 1 10 9 0 13 9 2 9 0 1 9 2 11 7 0 2 1 10 9 13 9 0 2 3 7 9 1 9 0 3 13 10 9 1 8 1 10 9 1 10 9 1 11 7 11 2
36 2 10 9 0 4 13 1 13 7 13 9 0 1 13 10 9 0 2 0 7 0 2 1 9 1 9 2 13 3 3 10 9 0 11 11 2
27 1 11 8 11 2 11 11 2 4 13 16 3 4 13 10 9 7 1 9 7 1 10 9 1 10 9 2
25 7 7 10 9 0 3 13 2 11 11 2 11 2 11 2 11 2 11 2 11 11 2 7 11 2
43 10 9 0 2 10 8 2 0 2 13 0 9 1 10 9 0 1 9 1 9 2 7 1 10 8 2 0 9 1 9 1 9 2 16 13 10 9 0 1 10 9 0 2
14 10 9 7 10 9 13 10 0 9 1 10 9 0 2
16 10 9 1 11 11 4 13 3 10 9 7 10 9 1 9 2
23 10 9 3 15 13 3 1 10 9 1 0 0 9 2 7 4 13 10 0 9 1 11 2
21 10 9 10 11 4 13 1 9 1 10 9 11 11 1 9 12 1 11 1 12 2
16 11 4 13 16 10 10 9 0 1 9 3 4 13 1 9 2
26 1 10 9 0 0 1 11 2 11 1 11 2 10 9 15 13 1 10 9 7 10 9 1 10 9 2
9 9 0 2 1 9 9 7 9 2
20 11 13 12 9 2 13 10 9 1 11 11 2 7 13 12 5 1 10 9 2
13 10 9 15 13 1 9 10 12 1 11 1 12 2
11 10 9 3 0 1 10 9 0 13 8 2
20 10 9 13 3 9 1 10 12 9 2 7 1 0 9 15 13 10 9 0 2
47 10 9 13 1 10 9 2 13 9 7 9 0 2 10 9 15 13 11 2 11 13 9 1 10 9 0 14 2 0 2 2 13 0 1 9 2 7 13 10 9 1 10 12 9 1 9 2
33 13 10 9 3 15 4 13 16 15 13 11 1 10 9 16 13 1 10 9 1 10 9 7 16 13 16 10 9 0 7 0 13 2
37 1 9 2 16 15 13 13 9 1 10 9 1 9 12 1 11 2 9 1 10 9 0 2 2 10 9 13 10 16 15 4 13 1 13 10 9 2
61 3 2 13 1 10 9 1 10 9 11 2 13 10 0 9 0 1 10 0 9 0 2 4 15 13 1 9 0 1 11 2 1 10 0 9 1 9 1 1 9 2 16 13 0 9 0 2 0 2 7 0 2 0 15 1 12 9 10 9 0 2
20 10 9 11 7 11 1 10 9 0 0 13 1 10 9 1 10 12 1 11 2
13 1 12 9 1 9 2 13 1 10 9 1 9 2
19 15 13 12 2 1 10 12 1 11 1 12 7 10 12 1 11 1 12 2
33 1 10 9 1 9 13 10 11 1 11 2 3 15 4 13 10 9 0 2 7 10 11 1 11 11 11 2 11 11 1 11 2 2
14 10 9 13 13 7 13 1 10 12 9 3 1 12 2
13 10 9 1 9 13 1 12 8 2 5 9 5 2
13 10 9 4 13 1 10 9 12 2 12 7 12 2
17 3 2 10 11 3 3 4 13 7 4 13 10 9 1 10 9 2
38 1 11 1 12 2 10 9 11 12 13 1 10 9 1 12 9 3 2 13 1 10 9 1 10 9 11 12 1 11 7 1 10 9 11 12 1 11 2
3 13 9 2
15 11 11 2 9 1 11 2 13 9 1 9 1 10 9 2
35 15 1 10 9 1 10 0 9 13 16 10 9 13 1 9 1 10 9 4 13 10 0 9 1 9 13 1 10 9 1 9 1 10 9 2
21 13 3 0 16 10 9 13 10 9 0 16 13 10 9 7 9 0 1 10 9 2
15 15 13 10 11 11 11 7 13 1 11 2 11 11 2 2
21 11 11 11 11 2 13 1 13 1 9 1 10 11 11 7 1 10 10 11 11 2
27 10 9 1 9 0 2 1 9 1 13 0 13 1 0 2 15 16 3 13 10 9 16 15 13 1 9 2
59 1 10 12 9 2 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
17 10 9 1 10 11 11 13 10 9 2 8 2 13 1 10 9 2
43 13 10 9 0 1 10 9 1 11 2 10 12 9 2 9 7 9 2 13 3 1 12 9 1 0 7 13 1 12 1 12 8 2 15 16 13 10 9 1 3 1 12 2
73 1 10 9 1 9 11 13 1 10 9 16 3 13 10 10 9 1 10 9 1 11 2 16 13 10 9 0 7 1 13 1 10 9 1 1 13 1 10 9 10 9 1 9 1 10 9 2 9 16 13 1 10 9 2 7 13 10 0 9 0 1 10 11 1 11 1 10 9 1 13 10 9 2
6 13 1 9 1 9 2
32 1 10 9 10 9 0 3 13 0 1 11 2 7 15 13 1 9 3 1 10 11 0 7 1 10 9 1 9 0 1 11 2
11 1 10 9 15 13 1 9 1 9 0 2
20 3 2 12 8 12 2 5 12 2 2 16 13 12 9 0 7 10 9 0 2
20 4 13 1 9 1 11 11 11 11 7 9 2 8 11 11 2 11 7 11 2
14 1 10 9 1 11 13 9 10 9 13 1 11 11 2
21 15 13 11 11 11 7 15 13 1 10 9 1 10 9 1 9 2 9 7 9 2
15 9 0 1 9 0 7 10 9 0 15 4 13 1 3 2
7 0 9 0 1 9 0 2
14 10 9 13 1 12 9 5 7 10 9 1 12 9 2
43 13 1 10 11 1 11 1 12 2 13 10 9 1 9 1 9 7 10 9 1 9 0 2 7 13 10 9 1 10 11 7 11 11 1 11 11 7 10 10 9 1 9 2
57 10 10 9 0 1 11 12 15 13 10 9 2 13 15 10 9 2 10 9 7 13 10 9 2 1 15 11 12 1 11 11 1 11 2 15 13 1 9 9 0 2 7 11 12 1 11 2 15 13 10 9 1 10 9 0 2 2
23 10 9 13 10 9 1 11 7 1 9 1 10 8 8 2 0 9 7 9 0 1 9 2
26 11 13 3 1 12 9 2 12 9 2 2 7 11 0 1 11 13 3 1 12 9 2 12 9 2 2
35 13 12 9 1 9 13 1 10 9 0 1 10 9 0 1 9 8 2 7 3 13 10 9 1 10 9 10 9 15 13 1 9 7 9 2
17 1 10 11 11 1 11 1 11 1 12 13 1 11 12 9 0 2
8 13 10 9 0 1 12 8 2
10 15 13 13 1 10 9 1 9 0 2
36 11 4 13 1 9 1 11 1 11 7 4 13 1 10 9 1 11 12 2 1 12 2 3 1 10 9 1 11 1 11 2 3 13 10 9 2
21 15 3 15 13 13 15 9 2 13 10 9 7 13 10 9 0 2 2 13 11 2
13 3 2 10 9 0 1 10 9 13 11 11 11 2
32 13 1 10 12 5 1 10 9 1 10 9 2 1 10 9 2 3 1 10 2 11 2 11 2 1 9 1 11 1 11 11 2
19 13 10 9 3 0 1 10 11 11 7 1 10 8 9 2 11 11 11 2
20 10 11 12 13 10 9 0 8 1 12 8 2 13 1 10 11 11 11 0 2
16 15 13 1 11 2 9 11 7 11 11 2 11 7 11 2 2
20 10 9 15 13 10 12 1 11 1 12 2 1 10 9 1 12 1 10 11 2
28 13 3 0 1 10 9 1 10 16 15 13 16 4 7 13 10 9 3 1 4 13 1 10 9 1 10 9 2
26 3 3 1 13 1 11 15 13 1 10 9 10 9 1 11 2 16 1 3 12 9 13 1 10 9 2
18 10 15 13 10 9 1 11 2 10 9 1 11 7 10 9 1 11 2
35 10 9 1 9 1 10 9 2 10 11 2 2 10 11 2 2 13 9 1 10 9 1 10 9 0 1 10 0 9 1 11 11 11 11 2
31 11 13 3 3 0 1 11 7 11 16 4 13 1 10 9 0 16 13 16 10 9 0 13 13 15 9 0 1 10 9 2
17 3 3 2 13 10 9 1 11 11 11 2 0 1 11 11 11 2
15 10 9 0 7 9 4 13 9 1 5 2 8 7 5 2
13 10 12 1 11 1 12 13 10 9 1 9 1 11
15 11 13 3 1 3 1 11 10 11 13 1 10 0 9 2
15 3 13 1 10 9 11 11 2 7 1 11 11 1 12 2
19 13 10 9 3 2 11 1 11 7 11 1 11 2 2 16 3 15 13 2
32 15 13 1 10 9 16 13 10 9 1 13 9 13 10 9 7 13 10 9 7 9 1 10 9 8 1 9 1 10 9 0 2
15 10 9 16 3 15 13 3 13 10 9 1 13 10 9 2
20 1 10 9 15 13 9 15 9 13 3 1 10 9 0 3 1 10 9 0 2
14 11 13 1 10 9 1 11 10 12 1 11 1 12 2
21 10 9 13 10 9 0 1 12 1 10 9 11 7 13 10 9 1 12 9 5 2
22 10 12 5 1 15 16 4 13 9 13 9 0 2 3 7 10 12 5 0 13 0 2
31 10 0 9 1 9 0 1 10 9 0 13 1 10 9 0 2 3 7 7 13 10 0 9 1 9 0 13 1 10 9 2
21 15 4 13 15 3 10 9 2 4 13 10 9 7 15 15 13 3 16 13 0 2
21 1 12 13 1 9 2 2 10 9 1 9 0 7 10 9 0 13 10 9 0 2
16 13 10 0 9 2 3 15 16 3 15 4 13 3 10 9 2
20 3 13 10 9 15 13 1 13 1 0 9 10 9 1 10 9 1 10 9 2
12 11 11 13 1 10 9 10 9 2 3 0 2
37 1 10 11 11 11 2 10 9 13 10 9 1 9 7 9 2 1 9 15 10 11 1 11 11 11 13 10 11 1 10 11 1 0 9 1 9 2
14 15 15 13 10 9 1 16 15 15 13 1 10 9 2
22 10 12 1 11 1 12 2 4 13 10 9 11 12 1 11 2 11 12 7 11 12 2
17 11 11 11 2 7 11 11 11 2 13 1 12 1 11 2 11 2
23 1 10 9 1 11 10 9 15 13 1 9 0 1 10 0 8 8 2 9 1 9 2 2
37 11 11 13 12 9 2 12 9 2 11 7 11 2 7 12 9 2 11 2 13 1 12 2 7 11 2 11 2 13 1 10 12 9 1 9 2 2
46 13 10 9 1 10 9 1 10 9 0 1 10 9 1 12 9 2 9 2 7 9 1 9 2 9 2 9 7 9 16 13 10 9 7 9 1 10 9 2 16 13 9 1 10 11 2
20 10 9 15 13 1 10 9 1 10 9 0 1 11 1 10 9 1 11 11 2
41 3 13 1 10 0 9 2 2 11 11 11 11 11 11 11 2 2 2 11 11 11 11 11 11 2 7 2 11 2 11 11 2 2 13 1 10 9 1 10 9 2
24 1 9 1 10 9 0 2 13 1 10 9 1 9 1 10 9 7 1 10 9 2 8 2 2
45 16 15 4 1 13 1 10 11 0 11 15 13 15 9 16 13 10 9 2 10 0 8 0 2 13 1 10 9 7 9 2 16 13 0 13 1 10 10 9 1 10 16 4 13 2
24 1 10 9 2 11 4 1 13 1 11 1 9 1 13 1 10 9 2 1 9 1 9 9 2
12 10 9 13 10 9 1 9 2 3 1 9 2
13 10 0 9 4 13 1 11 2 13 1 10 9 2
38 10 9 3 13 0 9 1 10 9 1 9 2 9 8 16 15 13 1 10 0 9 1 10 9 7 9 1 10 9 2 1 10 9 7 1 10 9 2
18 4 13 10 9 1 9 1 10 0 9 1 10 9 1 13 10 9 2
26 1 9 1 10 9 11 11 2 10 9 15 13 1 2 10 9 1 13 1 10 9 13 1 9 2 2
11 1 10 9 1 10 12 13 10 9 0 2
15 10 9 4 13 1 10 9 1 10 9 1 10 9 7 2
44 1 10 9 1 10 11 11 2 11 12 13 10 9 1 9 1 10 9 1 11 2 15 16 13 10 9 0 1 10 9 0 1 10 9 16 15 13 1 10 9 1 10 12 2
7 15 13 13 3 10 9 2
28 1 9 1 10 9 1 9 7 9 2 11 13 1 9 10 9 0 2 3 1 10 9 0 7 1 10 9 2
27 1 10 9 2 10 9 13 10 9 13 10 9 1 10 9 0 1 10 9 2 11 13 1 10 9 0 2
8 15 4 13 15 3 7 3 2
10 13 9 1 10 9 1 9 1 9 2
41 11 11 2 13 1 10 9 1 10 9 11 11 2 10 9 1 10 9 0 13 13 15 1 10 9 1 10 9 2 8 1 15 16 13 1 10 9 0 1 11 2
22 10 9 16 15 13 12 9 1 10 9 16 10 9 15 13 3 1 10 9 1 11 2
33 11 11 7 11 13 10 9 1 9 13 3 7 15 1 10 9 1 0 9 1 10 15 15 13 9 3 1 10 9 9 7 9 2
13 15 13 3 1 9 1 10 9 11 2 11 2 2
40 10 11 12 1 11 1 12 1 10 11 11 1 11 4 13 9 1 9 1 10 12 9 1 10 11 11 2 12 2 1 9 1 10 9 1 10 9 1 11 2
59 1 10 12 9 2 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
23 10 9 4 13 2 1 10 9 0 2 10 9 1 9 1 10 9 7 10 9 1 9 2
12 10 9 13 1 12 9 1 10 9 0 9 2
23 10 12 1 11 1 12 2 10 9 0 13 1 11 2 1 10 9 1 10 9 1 11 2
37 10 11 4 13 10 9 1 15 1 10 9 1 10 11 16 13 15 13 10 9 1 11 2 10 9 16 3 13 9 1 11 1 13 10 11 11 2
27 15 13 0 9 1 10 9 0 7 1 10 9 1 9 1 10 9 1 10 9 1 9 1 10 9 12 2
42 1 10 11 1 10 11 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
40 11 13 1 10 9 1 9 1 11 0 7 0 9 1 10 0 9 0 2 16 3 13 0 1 10 9 1 11 2 2 13 11 11 2 9 1 9 1 11 2
21 10 9 0 13 1 11 7 9 1 11 7 4 4 13 1 10 0 9 1 9 2
30 13 10 9 1 9 16 13 10 9 1 12 9 0 1 15 9 1 10 9 1 10 9 1 11 7 10 9 1 11 2
28 13 10 9 1 9 0 7 9 1 9 0 2 1 11 2 11 11 2 2 1 12 9 1 9 7 9 0 2
27 13 16 13 10 9 13 1 11 2 11 15 13 1 11 2 7 4 13 1 11 7 11 2 13 3 0 2
30 10 9 8 2 0 15 13 2 16 13 15 1 10 8 8 2 8 8 2 13 13 2 13 2 1 9 8 8 2 2
17 11 11 11 13 10 9 1 9 1 10 9 11 1 10 9 11 2
20 9 1 10 9 0 1 11 11 11 2 1 15 15 13 16 4 13 1 12 2
17 10 11 13 9 0 16 15 13 1 10 9 1 9 1 9 0 2
27 15 13 0 1 13 1 10 9 1 10 9 10 9 2 7 13 1 11 13 10 9 2 16 13 13 0 2
37 16 13 3 12 9 7 0 1 9 2 13 1 10 11 11 11 11 11 11 1 11 2 11 2 13 9 1 9 1 11 11 11 11 7 11 11 2
42 1 11 2 9 1 10 9 1 11 2 13 9 1 10 0 11 1 10 9 2 3 13 10 9 0 1 10 11 11 1 10 9 1 10 9 11 16 13 10 9 11 2
14 10 9 0 13 1 10 9 1 9 1 9 10 9 2
35 10 9 1 9 2 16 10 9 1 9 13 1 9 10 9 7 3 10 9 1 9 0 2 13 10 9 13 1 10 0 9 1 9 0 2
20 16 13 10 9 1 9 2 15 13 10 9 7 13 0 13 1 10 9 0 2
33 11 11 2 9 1 9 0 2 15 13 1 15 1 10 0 9 1 10 9 2 7 3 13 10 9 16 3 13 10 9 2 11 2
25 10 9 1 11 13 1 10 9 12 7 12 2 7 4 13 1 10 9 3 1 10 9 0 0 2
18 10 9 0 15 1 9 7 1 13 3 13 16 4 13 10 0 9 2
36 15 15 13 13 10 9 1 11 1 2 11 1 9 2 2 12 2 2 3 10 9 0 2 3 11 13 10 9 0 2 4 13 1 10 9 2
42 3 13 1 15 15 15 13 7 1 10 9 0 15 13 2 7 13 16 1 15 16 3 4 13 7 13 1 11 4 13 1 9 1 9 1 13 1 3 13 10 9 2
3 10 12 2
30 15 3 13 10 9 3 7 1 10 9 13 15 1 10 9 3 0 1 10 9 11 2 11 11 2 1 11 2 11 2
39 10 9 13 1 9 9 13 1 9 2 1 10 9 3 1 10 9 2 10 9 1 9 0 4 4 13 1 10 9 2 3 2 9 0 7 9 0 2 2
13 13 3 0 7 15 13 10 7 15 9 7 9 2
17 10 9 2 13 1 11 2 13 10 9 1 10 9 7 10 9 2
14 10 9 13 1 12 9 16 13 13 1 10 0 9 2
60 9 0 2 1 10 0 9 1 11 2 7 9 12 9 13 10 9 1 10 0 11 11 11 2 10 9 1 9 16 13 10 0 9 1 9 2 15 13 2 11 11 2 2 2 9 1 9 7 10 9 1 9 13 1 11 2 10 11 2 2
39 13 1 10 9 10 9 2 1 15 1 10 9 2 16 13 3 10 0 9 0 2 1 9 0 16 13 13 10 9 7 13 9 1 10 9 1 9 0 2
11 1 10 9 3 0 13 1 9 10 9 2
21 11 11 11 2 8 11 2 11 2 12 1 11 1 12 2 7 13 10 9 0 2
56 13 1 0 2 1 9 2 1 13 15 9 7 1 13 15 1 13 15 9 2 15 16 13 3 3 1 15 9 2 16 13 10 9 1 10 9 7 16 13 7 13 1 9 10 9 1 10 9 7 10 9 1 10 0 9 2
45 3 2 1 12 2 15 13 10 9 2 13 15 10 11 1 11 2 7 13 10 9 0 1 10 9 1 10 9 1 10 9 2 15 13 10 11 1 10 11 7 11 11 1 11 2
27 11 1 11 13 10 9 1 10 9 1 10 11 1 11 2 1 10 9 1 11 2 11 7 11 2 11 2
11 10 9 1 11 15 13 13 1 10 9 2
25 10 9 0 13 0 2 3 13 3 9 7 10 9 4 13 2 3 10 9 2 10 9 1 9 2
18 10 9 1 10 9 13 10 9 16 13 0 1 10 9 1 10 9 2
35 1 10 9 1 10 9 0 1 12 2 10 12 9 0 3 0 16 4 13 9 1 10 11 3 13 10 12 5 1 10 9 0 1 9 2
32 3 4 4 3 13 2 7 1 3 1 10 9 0 2 7 1 9 3 0 2 13 13 10 10 9 1 3 1 10 9 0 2
21 11 13 10 0 9 1 10 11 1 11 1 11 2 11 2 1 10 9 1 11 2
26 1 9 1 10 9 0 2 4 13 1 10 9 1 11 7 13 3 3 1 10 0 9 1 11 11 2
17 11 2 12 2 11 11 15 13 1 12 1 10 9 1 11 11 2
19 11 13 10 9 1 10 11 11 1 10 0 9 1 10 9 1 11 11 2
33 10 9 13 1 10 0 9 1 10 9 1 10 9 1 9 7 13 16 10 9 1 10 9 4 4 13 1 9 0 1 11 11 2
59 7 15 13 3 3 2 13 16 11 11 11 2 13 3 3 16 10 9 1 9 11 2 3 13 9 0 7 4 13 1 13 1 10 9 10 2 9 1 10 9 1 10 9 1 13 2 2 13 1 10 9 16 15 13 9 1 10 11 2
33 10 9 0 9 4 13 1 10 9 1 9 1 10 9 1 10 9 7 10 9 2 16 10 9 1 10 9 13 0 1 10 9 2
30 1 9 1 15 15 13 13 10 9 13 11 2 11 2 11 7 3 13 10 9 1 10 9 11 12 7 10 9 11 2
6 10 9 0 13 0 2
8 10 9 0 4 13 1 11 2
19 1 12 10 9 11 11 11 13 10 9 11 2 11 1 11 2 11 2 2
59 1 9 2 10 9 0 13 10 9 16 3 4 4 13 1 10 0 9 0 1 10 9 16 13 1 10 9 7 11 2 10 15 2 16 4 4 13 3 11 2 13 3 0 2 1 10 9 1 16 13 10 12 9 10 9 1 10 9 2
30 13 0 9 1 10 2 11 11 11 2 16 15 4 13 1 10 9 1 9 16 4 13 15 1 10 9 1 10 9 2
12 10 9 13 11 2 16 13 10 9 1 9 2
19 1 0 9 2 10 9 4 13 10 9 13 1 10 9 1 9 1 9 2
20 1 10 9 1 11 11 11 15 13 1 9 1 11 11 1 9 1 10 9 2
16 15 13 15 15 15 13 10 0 9 1 10 9 2 11 11 2
11 10 9 1 11 15 13 13 1 10 9 2
28 10 9 1 9 13 1 10 12 5 7 10 9 0 3 0 13 10 12 5 1 10 9 1 11 1 10 12 2
21 13 10 9 1 10 9 0 1 9 2 11 13 1 10 9 13 10 11 1 12 2
34 15 13 16 15 13 1 11 16 13 1 10 9 2 7 13 10 9 3 13 15 16 13 10 9 1 13 10 9 0 1 10 9 0 2
16 1 11 7 11 13 10 0 9 2 13 3 0 1 10 11 2
11 15 13 15 1 10 0 9 3 1 9 2
10 10 9 0 13 0 2 7 13 0 2
20 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 1 10 11 2
18 10 10 9 15 13 0 1 10 11 15 16 15 13 10 9 0 0 2
41 1 9 11 13 1 11 1 10 9 1 10 10 9 1 10 11 11 7 1 10 9 16 9 1 11 7 4 1 13 1 10 11 11 1 10 9 1 10 11 11 2
24 10 9 11 11 11 2 13 1 10 9 1 11 2 11 2 2 9 1 10 9 1 12 9 2
35 10 9 13 1 13 13 1 10 9 13 16 15 13 1 10 9 0 2 7 16 1 10 9 15 4 13 1 10 9 0 7 1 10 9 2
28 1 10 9 15 16 13 13 16 15 13 7 15 13 10 0 9 7 16 10 9 4 13 10 10 9 16 13 2
27 11 15 13 1 10 9 13 1 10 11 11 2 1 10 9 11 2 1 15 15 13 10 9 1 10 9 2
28 1 12 2 10 9 13 1 13 9 1 11 11 2 16 15 1 10 9 0 13 1 10 9 1 10 0 9 2
23 10 11 1 11 11 2 10 1 11 11 7 10 11 1 11 13 15 1 10 9 3 0 2
15 10 9 15 13 10 0 12 1 11 1 10 11 1 11 2
8 7 13 10 9 13 1 9 2
13 15 15 13 10 9 1 10 9 16 13 3 0 2
9 1 10 9 2 11 13 10 12 2
43 10 9 1 10 9 13 10 9 0 1 11 11 2 7 15 1 10 9 15 13 3 1 10 9 13 10 9 11 11 2 15 16 13 10 9 0 15 3 3 4 4 13 2
8 11 13 1 10 9 11 11 2
18 11 4 13 1 13 1 10 9 11 12 2 10 9 9 2 0 2 2
36 0 1 15 2 15 15 13 1 10 9 11 13 10 9 7 9 1 10 9 2 7 10 12 1 11 10 9 1 10 9 4 13 1 11 11 2
46 10 9 2 10 0 9 4 13 1 12 9 2 16 15 13 1 12 9 13 11 2 9 2 11 7 11 2 10 15 13 10 9 1 9 2 1 10 15 13 12 9 16 13 10 9 2
30 1 9 2 15 4 13 9 1 11 7 10 9 1 10 9 11 13 3 1 10 2 9 1 11 2 2 3 13 11 2
17 10 9 4 13 3 3 1 10 9 1 11 1 10 9 1 11 2
21 3 13 10 9 2 13 1 10 9 1 11 1 12 1 10 9 1 10 11 11 2
26 1 10 9 2 13 16 3 1 10 9 16 13 13 16 1 10 9 1 9 13 16 13 1 10 9 2
19 1 11 13 10 11 1 10 11 16 1 12 13 1 10 11 1 10 11 2
36 10 12 1 11 12 2 13 1 13 10 11 1 11 1 10 11 11 2 11 11 2 2 3 1 13 12 9 0 1 10 11 1 10 11 11 2
16 10 11 13 10 9 1 10 9 1 11 2 11 2 11 11 2
20 1 12 10 9 0 13 10 9 1 11 2 16 3 13 1 13 1 10 11 2
5 15 13 1 11 2
42 1 10 11 1 10 11 1 10 11 11 2 11 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 13 1 9 0 7 2 12 5 2 12 5 5 13 9 2
35 1 10 9 0 10 9 4 13 10 9 1 10 9 2 7 3 2 13 1 10 9 7 10 9 13 10 9 1 10 9 1 10 9 0 2
23 15 2 1 9 2 4 13 16 10 9 0 1 9 13 10 9 0 1 15 1 10 9 2
15 11 11 7 11 11 13 10 0 11 1 10 11 2 12 2
26 1 10 0 9 3 10 9 1 11 13 0 1 10 9 0 2 7 3 15 13 10 9 1 15 13 2
59 1 9 1 10 9 1 10 9 10 9 13 10 9 1 11 2 13 3 1 10 9 1 11 1 10 9 1 11 2 1 10 15 13 1 9 2 13 1 9 7 13 9 1 10 9 0 2 11 2 11 2 11 2 11 2 11 7 11 2
27 1 10 11 3 13 11 11 2 1 15 13 0 9 2 7 11 11 1 11 2 1 15 15 13 1 12 2
19 10 9 4 13 1 10 11 7 10 0 9 1 10 9 1 10 11 11 2
11 15 13 1 12 9 1 10 9 1 11 2
32 4 7 4 1 13 16 13 0 7 13 1 10 9 0 1 13 2 7 16 3 4 13 2 13 16 13 3 1 10 9 2 2
21 2 10 9 0 7 0 1 10 9 0 2 3 13 10 9 0 0 7 3 15 2
16 10 9 0 13 1 9 3 1 16 10 9 13 10 9 0 2
37 10 15 13 7 11 15 13 1 11 15 15 13 10 9 1 10 9 1 15 15 2 15 13 7 13 1 11 13 7 13 15 16 3 15 13 0 2
12 1 10 9 15 13 10 9 0 7 10 9 2
22 13 1 9 1 9 16 4 13 1 10 12 5 0 7 1 10 9 1 10 9 0 2
50 1 10 9 15 13 10 9 1 10 9 13 1 10 9 2 9 1 10 9 1 11 2 1 12 9 0 2 15 1 11 7 10 9 16 15 13 1 10 15 2 7 10 9 16 15 13 1 10 9 2
20 10 9 4 13 1 9 0 1 12 9 1 10 9 2 1 12 9 1 9 2
39 1 9 2 13 0 2 0 2 0 2 7 0 2 3 11 15 13 0 1 10 11 2 13 10 9 1 10 9 7 13 9 1 9 1 15 15 15 13 2
31 10 9 3 9 13 11 1 10 9 0 9 1 12 5 8 7 10 9 3 0 13 11 1 10 9 0 9 1 12 5 8
36 10 9 3 0 3 13 1 11 13 12 11 8 2 13 1 11 1 12 2 7 10 3 0 13 1 12 5 8 2 13 1 11 1 12 2 2
14 1 11 11 2 11 2 13 10 9 1 9 1 12 2
8 11 7 11 4 1 13 15 2
57 1 9 1 10 9 11 11 15 4 13 1 13 10 9 1 9 0 1 10 9 2 12 9 2 12 9 2 12 9 2 9 2 9 2 9 1 9 7 9 2 1 15 15 10 9 13 0 1 15 1 10 9 1 10 0 9 2
31 15 13 16 15 13 9 1 10 9 1 9 13 1 10 9 7 13 10 9 0 1 16 13 10 9 7 3 13 0 9 2
31 10 9 7 9 13 10 9 1 10 9 0 1 9 7 9 2 7 1 10 9 1 10 9 1 9 0 1 10 9 0 2
12 7 13 9 1 10 3 0 9 1 11 11 2
15 13 10 9 1 9 11 2 16 15 13 10 12 1 11 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
37 11 13 15 1 10 9 3 0 1 9 1 13 9 0 2 3 16 13 10 9 1 10 9 11 12 7 12 3 4 13 10 9 1 10 9 11 2
33 1 10 9 1 10 9 15 4 13 0 8 2 9 1 9 0 2 1 10 1 11 11 2 11 7 10 11 1 3 1 12 9 2
19 10 9 0 2 13 1 10 9 1 10 11 2 13 9 1 10 9 12 2
19 1 10 9 1 10 11 11 15 13 9 0 1 13 2 1 9 1 9 2
21 13 10 9 0 1 9 0 1 10 11 1 11 2 3 15 13 1 9 1 9 2
19 15 4 13 10 9 0 0 2 16 15 13 1 10 9 0 1 10 9 2
30 10 11 3 3 13 10 9 7 3 13 1 10 11 2 7 3 3 13 16 11 13 10 0 9 1 13 1 10 9 2
27 4 13 7 13 3 1 10 9 1 11 7 1 10 1 11 2 7 15 13 1 15 10 11 11 1 12 2
17 13 10 9 1 13 1 10 9 7 1 10 9 3 3 1 11 2
16 7 3 13 1 10 11 11 2 10 0 9 1 10 9 0 2
29 13 3 1 10 9 0 1 10 9 1 10 11 7 11 3 13 1 0 9 7 3 10 9 13 10 9 3 0 2
73 10 9 7 2 15 1 11 2 13 10 9 0 0 1 9 0 16 15 13 1 9 1 10 9 1 11 11 2 15 9 1 9 1 10 9 1 10 9 15 13 1 13 10 9 1 9 2 9 2 9 2 9 2 9 7 10 9 1 9 0 2 1 0 9 2 16 13 10 9 2 7 9 2
24 2 10 9 1 10 9 2 11 11 2 1 10 13 10 9 13 16 4 13 1 10 0 9 2
19 15 4 13 1 13 13 10 9 16 15 13 9 1 15 3 1 12 9 2
39 15 13 10 9 1 10 9 7 10 9 13 16 13 15 3 0 2 10 9 3 0 2 15 13 1 9 7 3 13 9 1 16 15 15 13 1 10 9 2
14 2 10 9 13 3 10 9 2 10 9 7 10 9 2
9 3 13 1 10 9 0 1 11 2
15 1 10 11 1 11 11 15 13 1 9 7 9 1 12 2
28 1 12 10 9 0 13 10 9 1 10 8 9 16 13 1 10 9 10 9 1 12 9 11 7 2 11 2 2
19 11 13 10 9 13 1 10 9 1 11 1 10 12 9 1 11 1 11 2
20 1 15 9 1 10 9 10 9 13 1 10 9 1 10 9 0 1 11 11 2
9 2 10 11 13 10 9 1 11 2
32 10 9 13 1 10 9 1 11 1 10 11 11 2 7 1 10 13 4 13 1 10 0 9 1 11 2 11 11 2 11 2 2
36 10 0 9 1 10 11 2 1 10 9 2 13 1 10 9 1 11 10 11 2 1 10 9 12 2 15 13 0 1 10 0 9 1 9 0 2
19 10 11 11 4 1 13 2 10 9 11 1 10 9 13 1 10 12 9 2
12 10 9 8 8 1 10 9 13 1 5 12 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
23 7 13 10 9 0 2 10 9 15 4 13 13 1 15 2 7 15 0 3 13 1 9 2
13 10 13 1 10 9 2 4 13 1 9 1 9 2
46 10 11 11 13 10 9 0 1 10 9 1 10 11 11 1 11 2 1 10 9 1 11 11 2 16 13 10 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 8 11 11 2
17 10 9 13 9 0 2 13 10 9 1 10 9 0 7 10 9 2
44 10 12 9 1 11 1 11 2 1 10 9 0 1 10 11 1 11 7 10 11 2 13 1 8 0 2 10 9 0 2 10 9 0 2 10 9 1 9 2 7 10 9 0 2
21 15 1 10 9 13 3 1 9 0 7 2 15 2 4 3 13 1 10 0 9 2
29 16 10 11 11 15 13 2 13 10 9 11 7 13 1 11 16 3 15 13 15 1 10 11 2 16 13 3 9 2
31 1 10 0 9 1 9 0 2 10 9 0 15 13 2 3 3 1 13 2 7 1 13 1 10 9 1 9 0 7 0 2
48 10 9 1 9 4 13 1 12 9 1 9 16 13 10 9 1 12 9 2 7 10 9 4 13 9 1 10 9 2 1 12 9 1 12 9 2 2 15 4 13 1 12 9 7 13 12 9 2
10 13 10 9 1 12 9 2 12 2 2
16 1 10 9 2 11 13 1 10 0 0 9 1 11 1 12 2
30 13 9 1 10 3 9 11 2 9 1 11 12 2 10 9 1 10 11 11 1 11 2 7 9 1 11 11 1 11 2
10 11 13 1 11 11 1 11 1 12 2
74 10 9 1 10 9 1 10 11 7 10 9 13 1 11 15 13 1 10 9 2 1 10 9 1 9 0 2 13 15 1 10 9 1 11 1 11 11 2 9 1 11 16 4 13 1 10 9 1 9 13 1 10 11 7 16 4 13 10 9 1 10 9 1 10 9 1 10 9 1 11 2 11 11 2
56 0 9 0 2 15 16 13 1 10 0 9 7 9 2 10 9 15 13 3 7 0 2 0 15 2 10 9 2 10 9 11 2 7 10 13 0 1 9 8 3 0 2 10 0 9 16 4 13 1 10 9 2 2 15 15 13
27 3 2 10 12 1 11 1 12 2 4 13 10 9 1 10 11 1 10 11 2 7 1 10 0 9 0 2
13 13 1 11 2 13 1 12 1 10 9 1 9 2
13 0 9 7 16 7 15 13 10 9 1 13 15 2
18 1 9 2 11 13 2 1 0 9 2 1 10 0 9 11 1 9 2
20 10 9 15 4 1 13 2 15 13 9 1 9 1 10 9 7 15 13 9 2
11 2 3 15 13 10 9 1 10 9 12 2
17 4 13 1 10 9 1 10 9 1 10 9 1 11 11 1 11 2
4 13 1 11 2
39 1 9 1 10 9 2 11 3 13 16 2 1 9 1 10 9 1 11 0 2 10 9 13 10 9 1 10 2 11 11 2 1 9 1 10 9 0 0 2
28 11 4 13 1 10 11 11 2 3 1 10 9 0 1 10 11 11 13 1 10 9 1 10 9 7 10 9 2
16 2 3 15 15 13 2 2 13 10 9 1 10 11 11 11 2
9 15 13 16 15 4 13 10 9 2
20 9 1 10 9 15 4 13 1 10 9 1 9 1 10 9 1 9 1 9 2
16 13 1 11 10 9 1 11 1 11 7 15 13 9 1 9 2
46 10 9 2 13 1 9 0 1 13 10 9 1 9 1 10 9 2 4 13 1 10 9 2 7 11 11 2 11 8 2 4 13 16 11 13 1 13 10 9 0 1 15 1 10 11 2
28 10 9 1 9 2 10 9 1 10 9 1 9 7 10 9 1 13 10 9 13 9 13 3 1 10 9 0 2
39 1 9 2 10 9 4 13 1 11 1 10 9 2 11 2 2 1 3 10 2 5 2 1 10 9 2 2 16 13 10 15 3 0 1 9 1 10 9 2
40 1 10 0 9 13 3 10 9 13 1 10 11 1 12 1 10 11 2 13 10 2 11 1 10 11 2 7 10 9 1 10 11 1 10 11 11 1 10 9 2
31 16 10 9 1 10 9 13 1 10 9 2 15 4 13 10 9 0 0 1 13 9 0 9 1 9 0 7 9 1 13 2
13 1 11 11 10 9 1 3 13 1 10 12 9 2
15 13 1 10 9 1 10 9 1 9 16 15 15 4 13 2
15 16 1 10 9 1 9 15 13 1 10 9 1 5 12 2
31 9 13 1 10 9 13 1 12 9 0 10 9 1 10 9 13 3 1 10 9 1 10 9 1 10 9 1 9 1 11 2
6 13 12 9 1 9 2
19 1 9 2 10 9 3 15 13 1 9 2 7 11 11 13 10 9 0 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
17 3 13 1 11 2 10 0 9 0 7 0 2 7 15 15 13 2
16 1 10 11 1 12 2 13 12 9 13 1 10 9 1 11 2
23 11 11 11 2 11 2 12 1 11 1 12 2 13 10 9 0 2 11 11 1 9 12 2
31 1 10 9 2 7 13 1 16 10 9 13 1 10 9 13 1 9 0 2 10 9 13 1 9 1 11 11 11 1 11 2
40 10 9 1 10 9 13 1 9 1 11 1 12 2 13 1 10 9 1 10 9 1 10 9 1 11 1 11 7 11 7 10 9 1 10 9 1 11 2 11 2
28 13 10 9 1 13 1 9 1 10 9 16 13 9 1 9 1 11 2 11 7 11 2 15 15 13 10 9 2
17 10 9 0 13 1 10 9 7 10 9 0 1 10 9 1 11 2
31 10 9 1 10 9 12 13 10 9 1 12 9 1 10 9 1 12 9 5 2 1 10 9 0 1 12 9 1 9 5 2
24 13 1 10 9 1 10 11 11 2 12 2 12 2 2 9 1 10 15 13 10 9 1 11 2
28 10 9 15 13 1 10 9 0 0 1 10 9 2 1 10 9 1 9 16 13 7 1 10 9 3 15 13 2
45 1 9 15 15 13 11 11 1 10 9 15 4 13 1 13 10 9 1 9 2 10 9 15 15 4 13 2 15 15 13 1 10 9 2 7 10 9 1 13 15 1 10 9 0 2
22 3 15 13 10 9 1 10 9 1 13 10 9 1 9 7 9 16 15 13 13 15 2
30 10 9 13 3 0 13 10 9 0 2 16 10 9 1 9 3 13 0 7 16 1 10 9 1 9 15 13 0 9 2
7 10 9 13 13 10 9 2
51 10 9 1 9 1 10 2 11 0 2 1 11 13 10 9 1 1 10 12 7 12 1 12 1 9 1 15 13 10 9 0 2 15 15 13 0 1 10 9 1 9 0 1 10 12 1 10 12 1 11 2
55 10 9 0 1 10 9 3 1 9 0 2 1 15 1 9 2 2 13 10 9 16 13 10 0 9 1 12 9 2 13 15 0 1 10 9 2 1 10 9 1 16 10 9 16 3 13 10 9 15 13 1 10 9 0 2
43 10 9 1 10 11 11 1 12 13 10 9 13 10 12 1 11 1 10 9 1 10 11 11 2 13 1 10 9 1 10 9 0 1 11 2 16 13 10 9 1 12 9 2
19 4 13 10 12 1 11 1 12 7 10 9 4 13 1 10 9 1 9 2
7 9 11 2 2 3 13 2
28 10 11 12 1 11 10 9 11 11 1 11 13 10 9 0 13 3 1 10 9 0 11 12 7 10 9 11 2
17 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 11 2
26 1 15 2 13 1 11 11 1 10 9 0 2 7 3 11 15 13 1 13 1 10 9 0 1 9 2
11 7 4 13 1 10 9 2 9 7 9 2
19 10 9 2 11 11 2 15 13 1 7 3 13 9 16 13 1 10 9 2
30 10 9 15 13 1 10 9 0 1 10 9 16 13 0 1 10 9 2 7 16 3 4 13 1 10 9 1 10 15 2
27 10 9 13 0 7 0 2 10 9 0 13 10 9 1 9 13 1 10 0 9 2 13 1 0 12 9 2
49 1 10 9 1 2 11 11 2 2 2 11 11 2 2 1 11 11 7 11 2 3 13 10 9 0 1 10 9 2 1 10 0 7 10 9 2 2 11 11 11 2 1 10 9 1 8 2 11 2
25 1 9 2 1 9 1 12 13 1 9 7 13 16 10 0 9 13 1 10 0 9 1 11 11 2
59 3 0 9 1 10 11 7 1 0 9 0 1 11 11 7 10 11 7 10 14 9 1 9 3 1 10 9 1 10 9 1 11 11 2 11 2 11 11 7 11 2 13 10 0 9 0 2 1 10 11 11 7 1 0 9 1 11 8 2
18 3 1 13 1 10 9 0 2 11 3 13 1 10 9 1 10 9 2
31 15 13 3 1 10 9 11 16 15 13 1 15 0 11 2 2 10 9 1 11 2 13 7 13 1 11 1 9 1 9 2
19 10 9 0 4 13 1 10 0 9 1 10 9 2 13 1 11 1 12 2
20 10 9 0 15 13 1 10 9 1 10 9 2 13 10 9 1 3 13 9 2
19 3 2 13 1 10 9 0 10 0 9 7 9 16 10 9 13 10 9 2
30 1 10 9 10 11 7 11 13 9 0 1 9 0 1 2 9 2 9 2 9 2 9 2 9 2 9 7 10 15 2
19 15 15 13 13 16 13 1 10 9 7 16 13 1 15 13 15 16 13 2
18 11 13 10 9 1 11 2 13 1 10 9 9 1 10 9 1 11 2
16 15 1 10 9 15 13 1 10 9 1 10 9 1 0 9 2
9 10 9 13 0 9 1 10 9 2
49 3 1 9 7 9 13 1 10 9 4 1 13 10 0 9 2 7 13 1 15 3 10 9 0 13 15 2 10 9 13 0 1 4 13 15 1 10 9 0 2 3 13 10 9 1 10 9 0 2
69 1 10 9 3 13 11 11 15 13 10 0 9 2 15 13 1 13 1 11 1 10 9 2 11 15 13 9 1 16 10 13 3 7 13 3 13 10 9 2 10 9 1 11 13 1 10 9 7 15 13 1 10 9 7 11 4 3 2 10 15 15 13 7 10 9 1 10 9 2
25 10 8 1 11 15 4 13 1 12 3 13 1 3 12 9 1 9 0 1 13 7 13 9 0 2
24 11 1 11 13 10 9 13 1 10 9 1 10 9 1 10 11 2 1 11 2 2 11 2 2
9 10 9 1 9 15 13 1 12 2
52 10 13 16 2 10 9 1 9 13 0 1 13 9 10 9 3 13 1 10 9 2 16 10 9 3 13 1 9 2 3 1 0 9 2 10 9 0 1 9 2 13 3 10 9 1 10 9 1 10 3 0 2
18 3 10 11 13 10 9 12 1 0 9 1 10 9 2 10 11 11 2
52 1 15 13 10 9 1 0 9 2 10 9 2 10 9 2 10 9 2 10 9 7 10 9 0 1 11 2 0 1 10 9 7 16 4 4 13 10 9 16 13 13 15 1 10 9 7 13 0 1 10 9 2
28 4 13 9 1 9 1 12 9 2 12 9 4 13 10 9 1 9 7 10 9 1 11 15 4 13 12 9 2
31 10 0 0 9 13 1 9 13 1 10 11 10 11 7 11 2 16 10 9 13 13 9 10 9 2 16 4 13 1 15 2
13 3 0 1 9 1 8 7 8 13 9 1 8 2
20 10 9 13 1 10 9 9 16 13 10 9 2 7 13 9 2 1 10 9 2
13 11 13 15 1 10 0 9 13 1 10 0 9 2
8 10 10 9 13 0 7 15 2
19 15 15 13 1 1 10 9 2 7 3 13 0 9 1 10 9 7 9 2
27 0 9 4 13 1 10 11 2 10 9 16 1 10 9 1 10 9 4 13 1 10 9 10 9 1 11 2
60 13 0 13 16 10 9 3 4 3 13 2 3 16 7 3 13 1 10 0 9 1 9 0 2 1 10 13 11 2 12 3 13 10 9 1 11 2 7 3 10 9 1 9 2 1 15 15 2 13 10 11 11 2 16 3 13 9 1 11 2
14 15 13 3 10 10 9 1 10 9 1 11 1 12 2
27 3 10 9 4 13 1 10 9 3 13 1 9 9 0 1 10 9 0 1 10 9 7 1 9 1 9 2
17 10 9 0 1 10 9 13 1 10 9 12 1 10 9 7 9 2
24 3 15 13 1 11 7 11 1 4 1 13 1 10 10 9 1 10 9 1 11 10 11 11 2
24 16 10 9 1 10 9 13 8 10 9 13 2 7 3 13 0 16 3 15 13 1 10 9 2
41 11 2 11 2 11 13 10 9 0 1 9 7 1 9 13 10 12 1 11 1 12 1 11 2 13 9 1 10 0 2 12 8 2 9 9 1 10 9 11 11 2
28 1 10 9 2 10 9 1 10 11 1 10 11 13 1 10 9 12 2 1 10 3 16 10 9 1 10 9 2
30 10 11 11 13 10 9 1 10 9 0 1 12 9 2 13 1 12 9 2 15 1 12 9 7 10 0 1 12 9 2
12 1 9 2 10 9 15 13 1 11 7 11 2
39 10 9 2 0 1 0 9 7 9 1 9 1 10 11 2 15 13 1 10 11 8 11 11 11 1 12 9 7 13 10 9 1 13 10 9 1 9 11 2
57 10 9 1 9 11 4 13 10 9 0 1 10 9 1 11 1 10 9 1 11 2 7 1 12 10 9 11 1 11 13 10 9 1 11 11 7 10 11 1 10 9 0 10 9 11 1 10 9 2 1 10 9 0 0 1 11 2
8 13 1 10 9 1 10 9 2
22 10 11 11 12 13 0 1 10 9 1 11 2 11 2 1 10 9 11 11 7 11 2
19 10 9 11 11 13 1 10 9 2 16 11 11 13 10 9 1 10 9 2
17 10 9 7 10 9 13 9 1 10 9 7 9 13 1 10 9 2
76 1 13 1 10 9 2 11 4 1 13 9 1 10 9 1 9 1 10 9 2 16 13 13 10 9 7 13 10 9 2 11 15 13 1 10 9 3 13 10 9 2 3 13 10 9 2 10 9 0 7 10 9 1 11 2 3 1 10 9 1 10 9 3 13 2 11 3 4 13 1 13 1 0 9 2 2
28 10 9 13 1 10 9 0 7 16 3 13 3 3 4 7 15 13 10 9 16 13 10 11 11 13 10 9 2
17 13 1 10 9 1 11 1 13 1 10 12 1 11 1 10 12 2
12 11 11 13 10 9 3 3 0 1 10 11 2
10 13 10 9 0 3 0 1 10 9 2
14 10 9 1 10 9 13 1 10 12 7 10 12 9 2
26 1 13 15 15 3 3 15 13 10 9 15 13 7 13 1 12 9 0 2 13 10 9 1 12 9 2
22 11 13 3 11 11 7 4 1 13 9 1 9 0 1 11 11 1 11 2 12 2 2
19 10 9 2 10 11 11 13 1 9 13 1 10 9 0 1 10 0 9 2
46 10 12 11 11 1 11 11 15 13 1 10 9 0 1 11 2 11 2 1 10 12 7 10 12 1 11 1 12 1 10 9 1 10 11 11 1 11 2 11 2 7 10 9 11 11 2
17 15 4 13 2 1 10 10 11 2 2 16 13 9 1 10 11 2
17 10 9 7 2 7 9 16 3 13 3 0 4 13 1 10 9 2
13 1 12 9 1 9 2 13 1 10 9 1 9 2
14 15 13 10 9 3 4 13 9 1 2 11 11 2 2
15 10 11 11 13 10 9 1 10 9 12 1 11 2 11 2
13 1 10 9 1 10 9 9 2 10 9 13 9 2
22 3 13 13 10 9 1 10 9 16 13 10 9 2 3 0 2 1 9 1 0 9 2
17 10 9 13 0 2 13 16 1 16 13 3 13 3 0 8 2 2
22 1 10 0 9 7 3 12 9 0 15 4 13 1 9 3 0 1 10 9 16 13 2
23 10 9 1 15 4 13 1 10 9 1 9 16 10 9 4 13 1 10 0 12 1 11 2
33 1 13 10 0 9 1 10 9 15 3 13 2 13 10 0 9 1 9 0 2 13 1 10 0 9 1 9 1 11 12 1 11 2
24 3 2 10 9 0 13 16 11 11 13 15 1 10 0 9 1 10 9 1 10 11 11 11 2
21 11 13 10 9 1 15 13 10 9 2 1 10 15 15 13 3 2 9 0 2 2
14 11 13 10 9 3 13 2 1 10 12 5 1 9 2
21 10 12 11 11 1 11 15 13 1 11 2 11 11 2 10 12 1 11 1 12 2
23 10 9 4 13 1 12 9 0 1 12 9 10 15 2 1 10 9 1 15 1 12 9 2
28 13 1 9 1 10 11 11 11 1 10 11 11 11 2 13 11 7 11 1 9 0 13 10 9 1 11 11 2
35 11 13 10 9 7 9 0 2 13 1 10 9 1 10 11 11 2 9 1 11 2 1 10 9 1 11 2 15 2 11 7 9 1 11 2
14 13 0 1 11 1 11 2 11 7 11 7 11 11 2
32 10 9 3 13 10 9 1 12 9 2 15 1 9 0 0 7 10 15 2 1 9 0 13 1 10 9 16 13 1 10 9 2
30 10 9 11 12 1 11 1 12 1 10 9 15 13 10 9 1 10 9 1 11 1 11 1 10 9 11 11 1 11 2
21 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
19 10 0 9 1 10 11 11 7 10 9 1 3 15 13 1 10 9 12 2
43 1 10 12 9 13 1 10 9 1 0 9 11 11 1 11 2 3 13 1 12 9 7 3 13 10 9 1 9 0 13 1 10 3 0 9 1 0 9 7 9 1 11 2
48 1 10 0 9 2 11 11 12 7 11 12 2 1 13 10 9 3 1 10 9 0 1 10 9 11 1 10 9 1 9 2 10 9 3 13 3 1 10 9 2 1 10 15 13 10 9 0 2
53 3 2 1 10 9 1 10 9 2 1 10 9 1 11 2 15 13 1 10 9 1 10 9 1 9 13 1 9 0 1 10 9 1 10 9 2 7 0 1 9 2 1 10 0 7 10 9 16 4 13 10 9 2
34 13 1 10 9 0 2 3 2 15 4 13 9 16 13 13 10 0 9 2 16 13 7 3 10 9 1 10 9 1 9 1 10 9 2
50 1 10 9 0 0 15 13 11 11 2 1 9 1 10 11 11 2 11 11 11 2 11 11 2 8 13 2 1 10 9 1 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2
12 1 12 13 10 9 0 1 10 9 1 9 2
29 13 1 10 9 1 10 9 0 2 1 10 9 0 0 7 10 9 0 2 10 0 9 0 3 0 7 10 0 2
15 13 10 9 0 1 10 9 1 10 9 1 11 7 11 2
15 13 1 10 9 15 13 10 9 1 11 11 7 9 0 2
7 2 3 13 10 9 3 2
55 10 9 1 11 13 10 9 0 16 13 9 10 12 1 11 1 12 1 10 9 1 10 0 9 2 1 11 2 1 10 9 1 10 11 11 2 0 2 12 2 2 13 1 10 11 1 10 11 11 1 10 11 11 11 2
75 10 9 1 9 13 16 13 1 10 9 1 9 8 2 0 7 0 1 10 15 1 10 9 2 3 2 1 9 2 13 9 1 15 10 9 3 15 13 1 10 9 1 10 9 0 2 3 2 7 16 13 3 9 0 7 1 9 1 2 1 9 2 10 9 1 10 15 10 9 4 13 10 9 2 2
33 15 15 13 10 9 2 16 8 16 13 1 10 9 1 10 12 1 10 9 1 10 9 1 11 3 13 9 1 13 1 10 9 0
12 10 9 13 13 15 2 7 3 13 10 9 2
15 11 15 4 1 13 10 9 1 9 1 10 9 1 9 2
15 16 13 1 0 9 1 9 1 9 0 4 4 13 11 2
30 3 2 11 13 1 9 1 9 1 11 7 15 13 16 15 3 4 13 10 9 2 7 13 10 9 7 15 13 15 2
25 4 13 9 1 9 1 9 1 10 9 0 1 2 11 11 2 11 11 7 11 11 11 1 11 2
43 1 10 9 1 10 9 1 10 11 11 2 11 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
19 10 9 16 10 9 13 1 9 2 9 7 9 3 9 1 10 9 0 2
61 10 0 9 1 9 1 10 8 9 0 7 10 9 1 10 9 1 10 9 2 15 13 16 3 3 13 1 9 7 9 0 1 13 10 9 1 9 1 10 9 2 7 16 15 4 13 10 9 1 9 0 1 10 9 1 9 1 9 1 9 2
10 11 4 13 1 10 9 1 10 9 2
34 13 9 1 10 9 0 1 10 8 2 16 15 13 10 9 1 9 2 1 15 9 4 7 13 10 9 1 10 11 11 2 2 13 2
22 2 11 11 11 2 9 0 1 9 1 10 9 1 11 2 13 10 9 1 10 9 2
13 13 1 3 0 9 0 1 10 9 0 1 11 2
26 1 10 9 2 10 9 15 13 1 9 0 2 7 3 15 13 3 7 13 0 9 1 9 7 9 2
18 10 9 1 10 9 13 0 1 10 0 9 1 10 9 1 10 9 2
17 7 1 10 9 13 10 9 7 10 9 1 9 0 1 10 9 2
20 9 0 1 10 9 0 2 15 13 1 10 9 7 13 1 10 9 1 9 2
20 1 12 13 10 9 1 10 11 2 3 13 10 9 1 10 9 0 1 9 2
17 1 10 9 2 13 1 11 10 12 1 15 9 16 3 7 13 2
28 10 0 9 1 10 9 0 1 10 9 13 12 9 1 10 11 1 10 0 9 1 9 1 10 9 1 11 2
24 0 9 1 10 9 15 4 13 9 1 10 9 1 10 9 11 11 7 10 9 11 7 11 2
42 12 9 13 10 9 16 10 9 13 1 10 9 2 15 13 1 3 1 10 9 2 13 1 10 9 7 13 1 10 9 2 10 9 13 1 3 10 9 13 10 9 2
31 2 2 2 15 15 4 13 16 1 15 15 4 13 3 3 7 10 9 1 15 1 10 9 13 16 10 9 13 10 9 2
13 10 11 15 13 0 1 0 9 1 9 1 11 2
10 15 13 10 9 7 12 9 1 9 2
16 10 9 1 10 9 13 10 0 9 1 9 2 13 10 9 2
17 10 9 15 13 1 9 1 12 9 2 15 1 9 7 15 1 9
12 10 9 4 13 1 10 9 2 11 11 2 2
41 3 2 13 3 10 9 0 7 0 9 1 9 0 15 16 13 1 10 11 11 1 11 1 13 15 1 9 7 0 2 1 15 15 13 3 13 1 10 9 0 2
11 10 9 0 13 1 9 1 9 1 9 2
12 3 2 10 9 3 13 0 7 3 15 13 2
12 1 3 16 3 13 1 13 15 1 10 9 2
52 0 9 2 13 7 13 1 15 9 1 10 9 2 13 1 9 10 9 15 13 0 2 13 13 2 15 13 1 10 9 1 10 9 7 15 3 13 11 2 10 9 15 13 2 1 9 2 11 2 11 2 2
17 10 12 1 10 0 9 15 13 10 9 1 9 1 10 0 11 2
18 1 10 0 9 13 0 9 13 1 10 9 2 15 1 15 1 9 2
17 10 9 0 1 10 9 15 13 1 10 9 3 0 1 10 9 2
20 10 9 13 1 13 10 9 2 13 2 13 7 13 1 10 9 13 2 3 2
37 1 10 9 2 13 1 10 9 12 2 10 9 1 11 11 11 13 9 1 10 9 1 10 11 11 1 10 9 1 11 2 1 10 15 4 13 2
41 13 10 9 0 1 11 0 2 13 1 11 2 9 2 2 11 2 9 2 2 11 2 11 2 11 2 11 7 11 2 9 2 7 1 10 11 11 2 9 2 2
22 10 9 0 13 16 13 10 9 1 10 9 0 7 15 3 13 15 0 1 10 9 2
25 10 9 1 2 10 11 2 13 11 11 11 2 11 11 2 7 10 9 2 11 2 11 11 2 2
27 16 10 9 13 10 9 1 10 9 1 9 0 7 0 2 15 1 15 4 13 1 9 0 9 1 9 2
28 12 5 11 13 10 9 1 10 9 11 11 1 10 9 1 11 11 1 10 9 5 1 10 11 11 11 11 2
24 13 1 9 1 10 9 1 10 12 3 1 10 9 1 9 13 1 10 9 1 11 11 11 2
36 3 15 13 0 2 1 9 1 9 7 10 9 2 7 10 9 2 1 10 15 1 9 0 2 13 10 9 3 0 7 1 15 15 13 0 2
9 3 13 10 9 1 11 1 15 2
21 11 11 13 10 9 1 10 9 0 16 10 9 3 13 15 15 13 1 10 9 2
33 1 10 9 10 9 15 13 1 10 9 2 3 15 13 10 9 1 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 2
19 13 10 9 1 10 9 1 11 7 10 9 0 1 11 3 1 11 11 2
10 16 13 1 11 13 10 9 1 11 2
40 16 15 13 15 2 16 13 1 10 9 7 16 15 13 10 9 0 7 16 4 13 1 10 9 0 2 16 11 13 0 16 3 1 13 15 0 3 13 0 2
18 11 3 15 13 1 10 9 1 10 11 2 11 2 1 10 9 11 2
29 10 0 9 1 10 12 9 13 16 15 16 13 1 11 3 13 9 2 1 9 15 16 13 1 11 3 15 13 2
24 3 1 10 9 7 10 9 2 10 9 13 10 9 1 9 0 7 0 3 7 3 0 3 2
59 1 9 1 0 2 10 11 11 1 11 11 2 11 2 7 10 11 11 11 11 11 2 11 2 13 1 11 1 10 9 0 1 10 9 2 1 10 9 7 1 11 10 9 13 1 10 9 13 10 13 9 1 10 9 1 10 9 0 2
41 13 1 10 9 1 10 9 1 11 2 1 10 9 1 11 2 7 11 11 2 1 10 9 1 11 2 1 10 9 1 11 7 1 10 9 1 11 2 11 2 2
41 10 9 15 11 13 13 15 1 13 10 9 2 3 13 11 2 7 1 10 9 1 10 9 1 10 11 1 11 1 10 9 1 11 3 16 15 13 11 7 11 2
25 15 13 1 10 0 9 0 1 10 9 1 15 16 13 1 9 1 10 9 2 3 10 9 13 2
25 1 10 9 3 0 2 10 9 4 1 13 15 0 7 1 13 10 9 1 9 0 1 10 9 2
10 10 9 1 9 3 15 13 10 9 2
8 13 10 9 1 9 7 9 2
31 10 9 1 10 11 2 9 11 1 10 11 2 13 13 10 9 1 13 10 9 2 10 9 1 10 9 7 1 10 9 2
11 10 9 13 9 0 1 12 12 9 0 2
14 11 4 13 1 3 1 12 9 1 13 10 10 9 2
10 13 10 9 1 10 11 11 1 11 2
59 10 9 1 10 9 1 10 9 1 10 9 3 3 13 1 10 9 0 2 0 1 15 3 13 10 0 9 0 1 10 13 10 9 1 8 0 1 10 9 0 16 4 13 10 9 1 10 13 9 3 1 10 9 16 4 13 1 9 2
21 1 9 1 10 9 1 11 2 1 9 2 1 11 15 13 12 1 10 12 9 2
43 1 11 7 11 4 13 9 1 9 2 13 3 1 9 2 7 1 9 3 1 11 7 11 2 2 1 9 2 10 9 1 11 1 12 5 2 7 10 9 3 12 5 2
31 1 9 0 2 15 13 1 8 7 13 10 9 0 2 13 1 15 1 9 2 13 10 9 13 1 0 9 1 12 9 2
12 13 0 1 11 2 3 7 1 10 9 0 2
36 10 11 1 10 11 15 13 1 10 9 0 2 1 9 1 10 9 1 10 9 1 10 0 9 1 11 1 10 11 2 11 2 11 7 11 2
27 3 2 10 9 3 13 9 7 13 1 10 9 0 10 9 1 0 9 13 3 0 1 15 1 10 9 2
23 10 12 1 11 1 12 15 13 10 9 0 7 11 15 13 1 10 10 9 1 10 11 2
32 13 1 9 2 13 3 0 7 13 3 9 1 10 9 1 9 2 16 9 1 10 9 4 13 15 1 9 13 1 9 0 2
58 1 9 2 10 9 15 13 10 0 9 1 9 13 1 12 2 15 16 3 13 10 9 0 2 13 1 9 1 10 0 9 1 10 9 7 1 10 9 2 15 3 4 13 1 9 1 9 7 9 1 10 9 3 0 1 11 11 2
36 3 2 16 13 1 11 2 11 11 15 13 1 10 9 1 9 3 1 10 11 11 2 13 15 1 10 15 16 13 1 10 9 1 10 9 2
21 10 9 0 1 10 9 13 2 1 9 2 2 2 3 2 7 2 7 13 2 2
36 11 11 7 11 13 1 10 9 0 3 1 10 9 2 7 16 10 12 9 15 13 2 11 11 15 13 10 9 1 11 7 11 4 13 11 2
38 3 15 4 13 16 7 13 1 9 2 10 9 13 0 2 3 15 13 10 9 1 9 2 7 10 9 1 9 2 3 13 1 10 9 11 1 11 2
9 13 10 9 1 9 16 13 0 2
21 10 11 11 1 11 13 1 11 11 1 11 13 15 1 10 9 1 10 0 9 2
53 16 13 10 9 0 1 10 9 0 7 15 15 13 2 16 10 9 15 13 3 0 2 1 9 2 3 7 13 1 9 1 10 9 3 4 1 13 15 1 13 10 9 1 9 7 1 9 2 0 7 8 0 2
35 10 0 9 13 0 1 10 9 11 11 1 10 9 10 11 1 10 11 2 15 3 4 4 13 3 2 1 10 9 2 1 10 9 0 2
41 9 0 16 15 15 13 0 2 4 1 13 15 16 13 10 9 2 13 3 3 7 3 3 7 0 9 16 13 3 3 13 10 9 2 13 9 0 7 13 9 2
10 15 13 1 10 11 11 2 11 2 2
17 13 1 11 1 10 9 1 9 7 9 3 1 10 9 11 11 2
30 1 10 9 1 9 13 16 13 16 13 10 9 1 10 9 11 2 11 2 11 11 7 10 9 1 11 11 1 11 2
19 16 10 9 1 9 1 10 9 13 0 1 10 1 10 9 1 10 9 2
25 10 9 13 9 1 13 10 9 1 4 13 15 0 2 7 1 10 9 2 13 10 0 9 0 2
57 1 11 11 1 9 2 13 10 9 0 1 10 15 13 10 9 1 8 8 1 10 10 9 2 7 10 9 1 10 15 15 13 9 1 10 9 1 11 1 11 2 3 1 9 1 10 9 7 9 13 1 10 9 1 9 11 2
10 15 13 1 9 2 13 1 12 9 2
43 1 10 9 12 4 13 3 1 10 9 0 1 10 9 11 11 1 10 9 1 11 7 11 2 7 4 13 3 1 13 10 9 0 9 1 10 9 1 11 2 1 11 2
46 1 15 2 1 9 1 10 11 1 11 2 10 9 13 1 10 9 1 9 2 16 13 1 10 12 5 1 10 9 0 1 9 0 2 15 16 13 10 0 7 0 9 1 10 9 2
33 16 10 9 13 10 9 2 9 2 1 10 9 2 10 9 13 10 9 1 10 9 2 7 15 13 15 1 10 9 1 10 9 2
65 1 10 9 13 1 10 9 9 1 10 9 1 10 9 2 10 9 15 13 1 11 9 1 9 0 1 10 9 1 9 1 10 9 0 7 0 1 10 9 1 10 12 12 12 9 1 9 7 1 10 9 1 9 0 1 9 0 0 1 12 9 12 12 9 2
13 1 10 9 15 13 16 13 7 16 13 10 9 2
43 1 10 9 13 16 11 11 13 1 10 9 1 11 11 2 1 13 15 1 10 10 0 9 16 13 1 10 9 7 3 13 13 10 9 1 10 9 1 10 9 0 2 2
20 15 13 9 0 1 10 9 0 1 10 9 1 11 1 9 1 9 7 9 2
12 1 11 10 9 11 13 10 9 1 12 9 2
18 1 10 9 13 10 9 0 11 11 2 13 13 10 9 1 12 9 2
22 10 11 11 13 10 9 1 10 9 1 10 11 11 11 2 13 1 10 11 1 11 2
37 1 9 0 1 10 13 15 15 13 9 16 1 10 9 0 13 10 9 2 10 9 1 9 2 16 8 15 4 13 13 1 10 9 1 10 9 2
28 1 12 2 10 9 0 1 11 13 1 10 9 0 1 12 9 2 9 16 13 9 3 1 10 12 1 12 2
11 11 3 13 9 1 11 1 10 9 0 2
24 1 10 9 2 16 13 10 11 1 11 2 13 13 10 9 1 10 11 11 7 11 11 11 2
16 13 2 1 10 9 2 1 10 15 11 12 13 10 11 11 2
13 11 11 11 13 10 9 1 9 1 10 9 11 2
20 1 10 9 12 5 13 9 2 12 5 9 7 12 5 1 12 7 3 9 2
11 10 9 13 3 10 9 0 7 10 9 2
28 10 9 1 10 9 2 1 9 2 13 15 3 16 10 0 9 1 11 7 3 4 13 3 1 10 9 0 2
6 10 9 3 4 13 2
36 10 9 4 13 10 9 1 1 10 3 12 9 1 9 7 13 0 10 9 2 16 15 13 1 10 9 1 11 2 1 9 2 1 10 9 2
9 13 10 0 11 11 1 10 9 2
15 10 9 4 13 1 11 11 2 11 11 2 8 11 11 2
34 11 11 2 13 10 12 1 11 1 12 2 13 10 9 0 1 9 0 2 13 10 9 1 9 1 11 11 11 1 10 11 11 11 2
14 4 13 3 1 9 0 7 1 9 1 9 1 9 2
41 10 9 2 16 3 13 11 11 11 2 4 13 10 9 1 10 9 2 10 9 2 13 1 10 9 0 2 13 10 0 9 1 10 9 1 3 1 10 0 9 2
18 10 9 1 10 9 11 1 11 11 4 13 10 12 1 11 1 12 2
35 13 1 11 2 11 2 2 1 10 0 7 0 9 0 1 11 12 1 11 2 11 10 11 2 7 11 12 1 11 2 9 10 11 2 2
17 11 11 13 1 10 9 12 13 9 1 9 1 10 9 1 11 2
44 10 9 8 13 1 10 9 1 10 0 9 1 9 2 11 12 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2
23 1 15 2 11 11 2 13 1 10 9 2 15 13 9 1 11 7 13 10 9 1 11 2
29 11 11 11 2 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 13 10 9 1 9 7 0 0 2
7 13 10 9 11 11 11 2
44 13 1 10 11 11 11 1 11 2 4 13 3 0 2 13 10 9 1 13 1 10 9 1 10 15 13 1 13 15 10 9 7 13 3 10 9 1 10 0 9 1 10 9 2
28 1 15 2 10 9 0 4 13 0 1 13 15 9 7 13 1 10 9 1 10 9 0 15 10 9 15 13 2
24 10 0 9 3 1 10 9 4 13 9 1 10 9 1 10 9 7 1 10 9 1 10 9 2
13 11 11 13 10 9 0 1 10 9 1 11 11 2
16 3 13 9 1 15 1 15 2 1 13 3 3 1 12 9 2
20 9 11 2 3 13 1 2 11 11 2 2 13 10 9 0 1 10 11 11 2
20 10 9 1 10 10 9 4 3 13 1 10 9 0 1 13 10 9 7 9 2
31 4 13 1 10 11 11 7 9 1 10 9 11 12 1 12 8 2 13 10 9 8 2 9 1 9 0 7 10 9 8 2
49 1 11 15 15 13 10 9 1 11 2 1 3 12 9 1 9 10 9 1 10 9 4 1 13 15 15 16 15 13 13 10 9 1 10 9 11 13 1 9 7 16 13 1 10 9 1 10 9 2
33 11 11 3 4 13 1 10 11 2 1 15 15 15 13 15 1 10 9 3 0 1 10 9 11 1 10 0 9 2 9 12 2 2
46 10 0 9 13 10 9 11 11 2 1 9 0 15 13 10 9 0 7 0 13 1 9 0 1 10 9 2 3 10 15 9 1 10 0 9 0 1 9 0 1 9 2 9 7 9 2
34 10 9 13 3 3 16 10 9 13 10 11 11 16 13 16 10 9 4 13 3 10 9 16 10 9 0 4 13 10 9 1 10 9 2
34 15 16 3 13 2 1 10 9 2 13 1 3 13 13 16 13 16 3 15 13 13 10 9 2 0 2 0 7 0 2 1 10 9 2
39 15 13 10 9 1 9 1 10 0 9 1 10 11 7 15 13 10 0 9 0 0 1 13 15 1 10 9 2 9 0 2 13 1 10 9 1 10 9 2
54 16 13 15 13 11 0 16 15 13 1 10 9 13 13 1 11 2 15 13 1 10 9 1 9 1 10 13 1 10 9 13 1 10 9 7 3 13 1 13 15 3 15 15 13 1 16 10 9 0 13 10 9 13 8
12 13 0 1 9 0 2 4 13 1 10 9 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
15 15 1 15 2 4 13 15 10 9 0 2 1 15 0 2
58 1 10 9 2 16 13 1 10 9 0 2 15 13 10 9 1 10 11 11 1 11 7 11 2 11 2 1 12 2 1 10 9 1 9 1 10 9 1 12 2 12 7 12 2 10 9 16 10 9 4 13 16 2 3 4 13 2 2
21 10 9 1 10 9 0 9 1 12 2 1 11 7 11 2 13 10 9 9 0 2
16 11 13 10 0 9 2 7 13 9 15 1 10 0 9 0 2
27 10 0 7 0 9 1 10 0 9 1 11 2 13 12 9 1 10 9 11 11 2 1 10 9 1 11 2
16 1 13 15 1 10 9 2 11 13 10 9 1 9 1 9 2
29 10 9 3 13 0 7 1 9 1 11 13 1 10 9 1 15 7 1 10 9 1 12 9 13 13 1 10 9 2
54 15 4 13 1 10 9 1 10 9 1 10 9 1 9 1 10 9 11 13 16 0 9 1 10 9 13 13 1 9 2 0 2 1 10 0 9 1 16 10 0 9 13 2 1 9 2 10 9 1 9 1 10 9 2
27 1 12 2 10 0 9 0 1 3 1 12 9 13 10 11 11 2 16 3 4 1 13 15 11 11 2 2
15 10 9 11 13 3 2 9 2 7 10 9 1 9 0 2
19 13 10 8 2 8 1 9 7 13 1 10 9 1 10 9 1 10 9 2
14 10 9 13 3 0 7 0 2 7 1 10 9 0 2
13 13 13 15 10 0 9 16 4 13 1 10 9 2
8 3 3 4 13 0 10 9 2
21 10 3 0 15 13 1 12 9 7 15 1 0 9 1 12 2 4 13 1 9 2
10 3 13 10 9 0 1 12 9 0 2
22 10 0 9 1 11 15 13 1 12 7 13 10 9 1 12 0 9 8 2 12 3 2
33 1 11 1 12 2 1 9 1 11 2 11 13 10 0 9 1 11 1 12 9 2 1 15 10 9 11 11 2 7 12 9 9 2
18 15 13 2 13 9 1 10 9 2 13 9 7 10 9 1 10 9 2
15 10 15 15 13 10 9 1 9 1 10 9 11 1 11 2
25 1 3 2 10 11 4 13 9 1 10 0 11 1 11 1 12 2 7 1 10 9 0 1 12 2
10 10 9 13 0 7 10 9 13 0 2
36 11 2 8 2 11 13 10 9 7 9 1 11 2 1 10 9 1 11 11 2 9 1 11 2 1 10 9 1 11 2 1 10 9 1 11 2
33 10 9 3 3 15 13 1 10 11 11 1 10 15 13 11 2 7 10 9 1 9 11 13 16 10 9 1 11 2 4 13 3 2
15 3 10 9 1 8 1 8 10 9 13 1 10 12 9 2
52 11 11 4 1 13 10 0 9 1 10 0 9 1 11 16 15 13 2 10 11 1 11 13 15 16 0 1 10 11 11 7 1 10 11 13 1 10 9 1 3 12 9 15 13 1 10 9 1 15 16 13 2
28 16 10 9 13 1 13 15 1 10 9 1 10 9 2 15 13 16 10 9 0 13 10 9 0 3 3 0 2
29 1 9 1 10 9 1 10 9 2 10 0 11 4 13 1 9 0 0 1 11 11 2 11 11 2 7 11 11 2
62 10 9 0 1 10 9 13 1 0 9 2 10 9 1 15 16 15 13 10 9 2 0 2 2 3 13 1 9 1 10 9 0 2 13 1 8 11 1 12 2 10 15 13 16 2 2 10 9 0 3 4 13 1 10 0 9 1 10 9 0 2 2
22 13 10 0 9 1 9 1 10 9 2 7 10 9 1 10 12 9 15 13 1 11 2
16 3 13 10 9 1 10 11 2 15 15 13 1 10 9 0 2
24 1 15 9 1 12 2 10 11 2 12 4 4 13 1 10 9 1 11 1 9 1 0 9 2
56 10 9 1 10 11 11 11 13 10 9 0 1 11 11 11 2 15 13 0 1 10 9 1 10 11 11 1 11 2 7 10 9 4 13 1 10 9 16 13 1 13 15 1 9 13 1 0 9 1 10 9 7 1 10 9 2
48 15 4 13 15 1 10 9 1 10 0 9 1 15 16 13 9 1 10 9 7 2 3 16 3 13 10 0 9 1 10 9 2 3 15 13 13 15 1 15 15 13 7 13 1 10 9 0 2
53 1 9 2 10 9 1 9 1 9 1 9 1 9 1 11 11 2 10 9 15 13 1 9 1 10 13 1 10 9 10 9 2 10 9 16 13 10 9 1 10 10 9 2 9 2 7 9 7 9 1 10 9 2
35 11 13 16 10 9 13 0 2 13 2 15 13 1 10 9 16 15 13 0 7 10 9 15 13 1 10 9 1 9 1 2 9 0 2 2
30 10 9 0 1 10 9 1 10 10 11 11 1 11 11 15 13 1 10 9 1 10 11 2 3 15 13 10 9 0 2
12 2 3 13 10 9 1 10 9 1 10 9 2
9 3 15 2 15 13 11 1 11 2
41 1 9 2 15 13 1 9 10 9 16 13 1 10 9 1 10 9 7 3 1 10 9 16 13 1 10 9 1 9 2 1 13 2 1 9 2 10 9 1 9 2
33 10 9 3 0 15 13 11 2 1 10 15 10 9 4 13 9 1 10 9 1 10 11 13 10 9 1 12 9 0 0 1 11 2
52 1 10 9 10 9 15 13 1 9 1 8 2 9 2 15 1 10 9 7 9 1 10 9 1 9 4 13 3 10 9 1 10 9 7 9 0 2 16 3 15 13 1 9 3 0 1 10 9 1 10 0 2
57 1 10 9 1 8 1 10 13 1 10 9 9 0 1 10 9 1 10 0 9 2 10 11 1 10 11 2 12 2 2 10 9 13 10 9 3 0 7 0 2 1 10 0 7 10 9 2 10 9 3 0 7 0 1 10 9 2
25 11 11 13 10 9 0 16 3 3 13 10 9 1 9 7 2 9 2 9 2 9 7 15 3 2
23 10 9 1 10 9 4 4 13 1 13 9 1 10 9 2 1 13 9 1 9 7 9 2
22 1 12 1 12 13 9 1 10 11 1 11 1 11 11 2 11 11 2 7 11 11 2
16 10 9 1 11 2 5 2 13 10 9 1 9 1 10 9 2
14 1 11 1 12 11 11 13 1 10 9 1 12 9 2
15 10 9 2 1 9 1 10 9 12 2 13 1 12 9 2
36 15 16 3 13 2 9 1 10 9 0 2 13 10 9 1 9 1 10 9 12 2 7 10 9 13 10 9 1 10 0 9 1 10 9 0 2
33 1 10 9 2 10 9 1 11 7 11 3 13 15 15 10 9 13 16 15 3 13 2 7 15 4 13 10 9 1 11 1 11 2
27 10 9 1 9 16 15 13 13 1 12 7 15 3 13 10 9 13 2 10 9 1 10 9 3 13 0 2
36 10 9 9 15 13 1 10 9 7 9 1 16 15 13 10 9 1 9 1 9 3 15 13 2 13 13 2 10 9 1 10 9 1 10 9 2
18 10 9 1 9 2 7 10 3 0 13 9 9 2 7 9 1 9 2
53 1 9 1 10 9 12 2 10 9 13 1 10 9 1 9 16 13 10 9 2 15 13 1 10 9 1 10 0 9 2 1 10 9 9 1 10 9 2 7 3 3 15 13 10 9 1 10 9 1 10 0 9 2
18 1 12 3 13 1 9 10 9 1 8 12 2 8 12 7 8 12 2
25 10 9 13 1 12 9 1 9 2 9 1 9 0 0 2 12 9 0 7 9 13 1 10 9 2
15 15 15 13 1 13 10 0 9 7 10 0 9 1 13 2
50 10 0 9 1 10 11 11 3 13 15 7 15 4 13 15 16 15 13 15 13 1 9 11 1 10 11 7 11 11 1 10 11 2 10 9 10 3 9 1 13 15 1 10 9 16 13 0 9 0 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 5 12 2 1 10 15 12 5 12 13 1 9 0 7 2 12 5 2 12 5 12 13 9 2
7 10 9 13 1 12 9 2
63 3 1 10 0 9 1 10 11 2 10 11 11 13 10 9 0 1 11 2 3 13 1 13 1 10 12 1 11 1 12 2 1 10 9 0 0 1 10 9 1 11 11 2 1 10 9 15 13 10 9 0 11 2 9 1 10 0 11 11 2 11 2 2
17 11 13 10 0 9 0 1 9 13 1 10 11 2 11 1 12 2
32 11 2 11 2 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
34 11 5 11 2 1 9 11 2 1 9 11 2 13 10 9 0 1 10 9 1 10 11 2 13 1 10 9 1 11 2 9 1 11 2
28 10 9 15 13 10 9 1 10 9 11 7 10 9 0 2 1 10 12 9 9 3 1 10 9 1 10 11 2
18 11 13 10 0 9 1 9 1 11 11 2 11 1 10 9 1 9 2
37 1 10 9 1 10 9 11 2 16 4 13 1 10 11 11 1 12 7 12 2 11 13 13 1 11 11 2 9 1 11 7 13 1 9 1 11 2
86 10 9 7 10 9 15 13 1 9 1 3 1 12 0 1 10 9 2 13 1 15 2 16 11 15 13 1 10 9 2 7 13 9 1 13 10 9 2 7 13 10 9 2 1 7 15 13 9 10 9 1 10 9 2 15 10 15 15 13 1 13 9 2 16 10 16 3 15 13 4 1 10 9 1 10 9 0 2 7 1 15 13 1 10 9 2
12 13 1 15 1 10 9 1 9 1 9 0 2
56 11 8 11 11 2 1 11 13 1 2 11 11 2 13 10 9 1 9 2 9 8 3 12 9 0 2 3 10 9 7 10 9 2 2 4 13 1 13 1 10 9 1 9 0 2 1 10 9 1 10 9 1 13 10 9 2
20 10 9 2 9 7 9 15 13 3 1 15 1 10 9 0 1 10 9 0 2
21 13 12 9 0 2 10 9 7 10 9 2 9 0 1 10 11 7 11 2 3 2
35 1 10 11 11 13 10 9 1 16 11 7 11 4 13 2 3 1 10 9 13 1 11 7 11 2 12 9 16 3 13 1 13 10 9 2
7 10 9 4 13 1 12 2
45 3 2 1 10 0 9 1 10 12 1 11 16 15 13 1 10 9 16 13 1 10 11 1 10 11 1 11 2 10 9 1 10 9 2 3 15 4 1 13 10 9 1 10 9 2
25 10 11 1 11 2 9 2 11 11 2 13 10 9 0 1 10 9 1 11 2 1 11 2 11 2
36 10 9 2 3 10 9 0 1 11 2 11 11 2 13 3 0 1 11 9 16 10 9 1 10 9 4 13 3 1 10 9 1 10 9 0 2
51 3 0 2 13 13 10 9 1 10 9 15 10 9 0 13 1 9 1 11 2 13 11 7 10 11 11 2 15 16 4 13 16 10 9 2 11 11 2 4 13 1 10 9 1 9 1 2 9 0 2 2
21 1 9 1 10 9 0 2 4 1 13 9 1 10 0 9 1 9 1 10 9 2
34 1 9 13 10 9 0 1 13 9 2 13 3 1 3 7 13 3 2 9 16 3 1 9 3 15 13 1 10 9 1 10 9 2 2
26 1 15 15 13 10 9 1 10 9 2 3 15 13 13 10 9 1 10 9 0 13 1 10 9 0 2
27 10 0 9 1 9 15 13 1 9 7 9 1 10 9 0 13 1 10 9 3 0 1 10 9 1 11 2
11 10 12 9 0 13 10 9 1 12 9 2
11 13 10 0 9 2 11 11 2 8 2 2
12 3 15 4 13 10 0 9 1 10 11 11 2
17 11 2 15 13 1 13 1 10 9 1 13 10 9 1 10 9 2
47 1 11 15 13 1 10 11 2 9 0 2 13 10 11 2 9 1 9 2 2 10 11 2 10 9 1 9 7 9 2 2 7 10 11 2 9 1 9 1 9 13 1 9 7 9 2 2
27 13 1 11 11 1 11 2 12 2 7 1 11 11 1 10 11 3 1 13 9 1 15 1 10 9 0 2
24 15 13 10 0 9 1 9 2 1 10 9 1 10 11 2 1 10 9 1 10 9 0 0 2
33 9 1 13 10 9 1 13 7 13 9 1 9 13 15 16 13 1 10 9 11 3 16 13 10 0 9 1 10 9 0 7 0 2
34 11 2 11 2 11 2 15 13 1 3 0 9 7 2 11 2 13 9 10 9 0 1 10 9 1 12 9 1 10 9 1 11 11 2
22 1 9 2 4 13 1 10 9 1 10 9 2 3 0 2 7 10 0 9 1 9 2
8 2 1 10 9 3 13 15 2
42 10 9 1 11 13 10 0 9 0 1 10 9 0 0 2 1 10 9 1 10 9 11 7 11 1 10 9 1 10 11 11 2 13 1 10 9 7 9 1 10 9 2
33 4 13 15 10 9 1 9 0 1 11 11 1 10 9 16 13 1 10 9 0 7 10 9 13 16 13 3 0 7 13 10 9 2
13 10 9 13 16 10 9 0 13 0 1 10 9 2
25 1 12 13 10 9 0 11 1 11 11 11 2 13 3 9 1 11 11 1 10 9 11 1 11 2
45 3 2 1 9 2 10 9 1 10 9 1 10 9 0 13 16 15 3 15 13 1 9 1 10 9 2 16 3 13 1 10 9 2 7 16 10 9 1 11 1 10 9 13 0 2
12 13 10 9 10 9 11 11 1 10 9 0 2
34 11 13 10 0 9 1 10 11 11 2 9 16 4 13 3 10 9 15 4 13 7 3 13 7 10 9 1 10 9 13 1 10 11 2
11 15 13 10 9 7 15 13 10 9 0 2
42 3 1 10 9 1 2 11 11 2 11 2 1 12 2 15 13 1 13 9 7 9 1 9 0 1 9 1 9 0 1 10 9 0 2 10 9 0 7 10 9 0 2
27 8 2 8 8 8 8 8 13 10 9 1 9 13 7 13 1 11 1 12 1 11 11 11 7 11 12 2
27 10 9 3 13 15 7 10 9 1 11 11 11 2 11 11 2 15 3 4 1 13 10 9 1 10 9 2
35 3 2 15 13 9 1 9 2 9 0 7 1 10 9 7 9 0 2 1 9 0 2 1 15 16 13 1 9 10 9 11 7 11 11 2
46 13 13 10 9 7 13 9 1 10 9 1 10 9 1 15 15 1 12 13 1 10 11 11 1 11 7 12 13 1 10 9 0 1 10 11 12 13 10 11 11 1 10 9 11 11 2
34 10 9 1 11 15 13 1 9 1 9 2 13 13 1 10 9 1 10 9 16 15 13 1 9 1 9 2 3 1 9 1 10 9 2
12 1 9 2 10 9 4 1 13 15 1 12 2
37 3 13 7 1 12 16 10 9 2 9 1 10 9 2 9 7 9 1 10 9 1 10 9 2 9 1 10 9 7 9 1 10 9 2 15 13 2
38 1 9 0 1 10 9 1 11 2 9 2 10 9 2 13 10 9 0 2 7 1 10 9 0 2 9 15 10 9 0 15 13 1 13 1 10 9 2
39 1 9 1 13 10 9 1 16 4 1 13 3 10 9 3 2 11 3 13 1 10 9 7 9 7 13 13 10 9 1 9 1 10 9 1 10 9 0 2
26 10 9 13 1 10 9 2 1 10 9 2 13 2 13 2 13 7 13 10 9 16 13 1 10 9 2
17 10 9 1 9 13 11 1 11 11 15 13 1 13 1 10 9 2
16 10 3 0 13 3 10 1 11 11 1 11 2 11 11 2 2
39 10 0 9 2 16 15 13 12 9 1 9 2 4 1 13 10 9 1 9 1 10 9 1 9 1 11 7 11 2 15 1 10 0 9 1 10 9 0 2
18 1 12 13 9 1 10 9 0 0 1 10 4 13 1 9 1 9 2
27 15 13 1 10 9 1 12 1 10 9 1 10 9 15 13 11 11 1 11 13 1 10 11 11 1 12 2
21 15 3 13 1 10 0 9 1 10 9 3 10 9 13 9 1 9 1 10 9 2
12 3 13 10 9 0 11 11 11 2 1 12 2
7 4 13 10 9 1 15 2
66 10 9 1 10 9 0 1 10 11 2 11 11 2 13 10 9 1 10 9 1 13 10 9 1 3 12 9 1 9 1 11 2 7 13 16 10 9 13 3 16 10 9 3 15 13 1 10 9 1 10 9 7 3 10 11 13 2 9 0 3 2 7 3 3 2 2
13 3 13 1 10 9 0 0 7 1 10 9 11 2
44 15 4 13 12 9 7 13 12 9 2 1 10 16 15 4 13 12 9 1 9 16 4 13 10 9 1 3 0 16 13 2 1 10 16 13 15 1 10 9 3 0 1 11 2
15 8 1 10 9 2 13 12 10 9 1 10 9 1 11 2
14 4 13 1 12 7 13 10 9 1 10 9 11 11 2
27 11 13 1 10 0 9 2 11 11 2 16 13 10 9 1 10 9 7 15 13 10 9 1 10 9 11 2
6 15 15 4 13 3 2
26 1 10 9 13 1 11 2 11 2 2 16 1 10 3 13 15 1 10 0 9 0 7 0 1 11 2
29 10 11 2 1 9 11 2 13 10 9 0 1 10 9 0 8 10 9 1 9 0 1 9 0 1 9 1 9 2
22 1 9 1 11 2 15 13 1 10 9 1 10 11 2 1 9 9 2 1 10 9 2
35 1 11 11 13 1 10 9 2 1 10 9 12 13 10 0 9 1 10 11 11 13 1 10 9 1 9 1 10 9 1 10 9 11 8 2
26 10 9 1 10 9 7 10 9 0 2 3 7 10 9 2 9 7 10 9 13 0 7 13 1 9 2
30 10 9 0 1 10 11 1 12 15 13 10 12 1 11 1 12 1 13 1 10 0 9 1 10 11 1 10 9 12 2
24 9 1 11 12 10 11 7 1 10 9 13 1 11 11 2 16 13 12 9 0 1 10 9 2
33 4 7 13 16 13 10 9 0 16 4 13 10 9 7 13 15 1 10 9 3 13 7 2 1 9 2 1 11 3 4 13 9 2
13 11 2 3 1 11 2 13 10 0 9 1 12 2
29 15 1 10 9 2 13 11 7 11 2 15 13 1 10 9 7 13 13 15 1 7 13 10 9 1 10 9 0 2
35 1 10 9 1 11 2 11 2 2 11 13 9 7 9 0 1 10 9 1 9 2 13 1 11 2 11 2 11 2 11 2 11 7 11 2
18 13 1 10 9 11 11 1 10 11 11 3 7 13 1 10 11 11 2
24 10 9 1 9 13 13 1 10 9 10 11 2 7 10 9 13 3 10 11 0 1 9 0 2
26 11 10 11 1 10 11 13 10 0 9 1 10 9 0 11 2 13 1 12 1 9 2 9 7 9 2
11 3 15 13 10 11 2 7 13 3 3 2
43 3 2 7 1 13 10 9 10 9 0 3 13 3 11 2 7 10 11 1 11 7 11 2 10 9 0 13 9 1 9 7 9 13 1 9 1 11 11 11 2 11 2 2
37 3 1 10 9 1 10 9 2 13 0 9 16 13 16 10 9 0 13 2 13 2 1 10 9 2 3 1 16 15 4 13 10 9 1 10 9 2
51 1 10 9 1 10 9 0 11 11 11 2 7 1 10 9 1 9 1 11 2 15 4 13 10 0 9 1 10 16 13 9 3 12 9 1 9 2 16 13 13 9 9 1 10 0 9 16 15 4 13 2
21 10 9 9 2 9 15 13 1 11 13 7 13 10 9 1 10 9 1 10 9 2
7 15 13 10 9 1 11 2
31 10 9 1 9 15 13 1 13 15 9 7 9 2 7 3 15 13 1 9 2 9 7 1 10 9 0 1 13 10 9 2
14 1 10 9 13 10 9 1 9 1 10 9 10 11 2
24 10 9 4 13 1 10 9 1 9 0 1 11 2 7 15 13 1 10 11 1 11 1 12 2
32 11 11 13 10 9 1 12 9 2 12 9 2 1 0 9 1 10 9 11 7 10 9 1 11 1 10 11 1 11 1 11 2
42 1 9 1 10 9 0 10 9 4 4 13 1 10 9 0 1 10 10 9 0 2 7 3 15 15 13 9 8 1 11 7 15 15 13 1 11 2 8 2 11 2 2
27 15 4 13 1 9 16 13 15 1 10 9 7 3 13 9 2 7 15 13 1 15 15 7 11 1 15 2
25 10 9 15 13 11 11 12 11 2 7 4 13 1 10 9 11 3 3 3 1 16 15 4 13 2
36 10 8 13 3 16 15 4 13 10 9 1 10 9 1 13 1 9 10 9 0 2 16 4 13 15 1 9 0 1 16 13 1 9 10 9 2
10 11 13 10 9 1 10 0 9 0 2
16 3 4 13 9 1 10 9 2 13 13 1 15 7 1 15 2
4 2 7 3 2
20 11 2 1 9 11 1 11 2 13 10 9 1 10 9 1 11 2 1 11 2
24 10 9 0 1 10 9 0 1 10 9 13 10 11 11 2 1 11 11 2 7 10 11 11 2
29 1 11 2 10 9 1 9 13 10 0 9 1 10 9 1 9 7 15 13 0 10 9 1 9 1 11 1 11 2
12 10 9 13 0 7 0 7 1 9 13 0 2
58 0 13 16 2 1 10 0 9 2 10 9 13 10 9 1 10 0 9 0 13 1 10 9 1 9 7 9 2 1 10 15 15 13 1 15 10 0 9 1 10 9 1 13 15 7 13 1 15 7 1 10 9 3 13 0 9 0 2
20 10 9 13 10 9 15 13 11 11 1 10 9 1 11 11 1 9 1 9 2
29 1 10 9 1 11 11 1 11 2 11 11 13 9 1 10 11 11 1 11 1 12 7 12 2 9 1 10 9 2
17 1 10 9 13 10 9 1 10 9 7 10 9 1 10 9 0 2
14 11 15 13 2 3 15 13 2 15 13 9 1 9 2
23 15 13 1 10 9 0 2 0 2 1 12 9 3 0 7 10 9 1 9 1 10 9 2
13 15 13 1 11 2 9 1 10 9 1 10 11 2
26 11 15 13 16 3 15 13 3 7 12 9 0 2 1 15 16 4 13 9 1 10 9 10 9 3 2
28 10 9 0 13 10 9 1 10 9 15 13 1 9 1 9 16 4 13 9 1 9 0 1 9 0 1 11 2
73 1 10 9 0 1 10 11 11 7 1 10 9 0 7 0 2 1 10 9 1 9 2 9 2 9 2 9 2 9 7 9 2 15 13 10 9 1 13 1 10 2 11 11 1 11 11 2 16 15 13 10 9 12 1 11 1 10 9 2 1 10 9 2 11 11 11 2 1 10 9 1 11 2
11 10 9 1 9 1 9 0 1 10 9 2
8 11 15 13 1 13 10 9 2
21 1 10 9 12 2 10 9 7 9 13 1 9 1 9 1 10 9 10 9 11 2
45 3 13 9 1 9 1 9 1 9 1 11 11 7 3 1 9 1 11 11 3 1 13 10 11 1 11 1 11 1 11 11 7 11 11 2 9 1 10 9 10 11 1 11 2 2
21 0 9 2 13 10 9 16 13 1 15 2 13 10 0 9 9 1 10 0 9 2
23 13 10 9 1 13 9 2 13 7 10 9 13 3 2 7 10 15 16 13 13 0 9 2
63 1 10 12 9 2 10 9 1 11 11 4 0 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
25 10 9 1 11 3 13 10 9 13 9 16 13 0 1 10 9 1 9 1 10 9 7 10 9 2
36 10 0 2 10 1 11 13 1 9 1 10 12 9 7 10 0 2 10 9 13 10 12 9 1 9 16 13 1 10 9 10 11 1 11 11 2
40 11 2 11 11 13 9 1 9 7 13 1 15 10 9 0 1 11 11 1 2 11 11 2 12 2 2 8 7 11 11 2 12 2 8 10 11 2 12 2 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
20 1 3 1 10 9 0 13 9 1 12 9 7 13 0 1 10 9 11 11 2
20 10 9 13 10 9 13 1 10 9 1 11 2 11 2 11 2 11 7 11 2
16 3 13 10 9 1 10 9 0 10 9 1 10 0 9 0 2
32 3 1 13 9 1 9 0 1 9 2 10 9 13 0 9 0 2 1 2 10 9 1 9 1 10 9 2 9 2 9 0 2
27 0 9 1 9 15 13 13 1 10 9 2 7 10 9 0 13 1 10 9 0 13 10 9 2 11 11 2
12 11 11 11 11 13 10 9 7 0 9 0 2
32 3 4 1 13 15 1 10 11 11 2 3 15 1 10 9 2 1 10 9 1 10 9 2 3 0 7 0 2 2 4 13 2
27 10 9 13 10 0 9 1 9 1 11 2 12 9 2 12 9 2 3 10 9 0 2 7 12 9 0 2
47 10 9 3 15 13 1 9 1 12 9 1 10 9 12 2 12 7 12 1 10 9 7 1 10 9 12 2 12 7 12 1 10 9 16 13 10 9 1 10 9 2 1 3 1 11 11 2
33 10 11 11 7 11 11 2 11 11 2 13 10 9 1 9 1 10 9 1 10 11 2 16 15 13 1 11 1 10 9 1 11 2
82 1 11 2 3 15 4 2 13 1 0 9 1 9 1 10 9 2 1 10 9 1 2 9 2 1 10 9 1 16 2 4 13 15 2 1 10 9 2 7 13 9 1 10 9 1 9 2 3 1 16 10 9 1 9 13 1 10 9 1 9 1 11 1 10 9 1 10 9 1 11 4 13 1 12 9 1 9 1 10 9 0 2
27 9 1 13 10 9 3 0 1 10 2 11 11 2 2 13 9 10 9 3 1 10 9 3 0 7 11 2
41 10 9 1 10 9 13 0 1 10 0 7 10 1 10 10 9 0 2 16 13 12 9 1 10 9 1 10 9 2 15 0 1 10 11 2 15 0 7 15 0 2
31 3 2 13 10 9 0 1 9 2 9 7 9 2 7 1 10 9 13 15 0 1 13 15 3 2 2 13 10 0 11 2
18 4 4 13 1 11 1 10 9 0 1 10 9 0 1 11 1 12 2
22 11 11 13 10 9 0 2 13 1 11 11 2 10 0 9 1 12 9 1 11 11 2
17 1 9 2 1 10 0 9 4 13 1 9 0 1 9 1 9 2
46 1 10 9 10 0 9 1 10 9 0 13 15 12 2 3 13 1 9 2 12 2 2 16 13 0 9 1 9 3 0 2 3 11 2 8 8 2 12 2 7 3 8 2 12 2 2
64 1 10 0 9 1 10 9 12 2 10 9 13 10 9 1 10 10 0 9 1 10 9 11 11 11 2 9 15 4 13 1 10 11 11 1 11 7 13 1 10 9 1 10 9 0 1 10 9 1 9 1 13 10 9 1 10 9 1 0 9 1 10 9 2
20 15 15 13 1 13 1 9 1 11 10 9 1 12 7 12 2 15 4 13 2
37 10 9 1 10 9 2 11 11 11 2 13 16 3 1 13 10 9 1 9 0 13 1 11 11 2 16 13 10 9 7 13 16 4 13 10 9 2
35 10 0 9 13 3 15 2 3 7 16 1 9 15 13 13 1 10 9 2 10 9 15 15 13 0 7 13 3 10 10 9 1 10 9 2
29 1 10 9 1 10 9 1 9 3 0 2 10 9 4 13 1 9 0 2 1 10 9 1 13 9 0 1 9 2
29 10 12 1 11 1 12 13 10 9 0 11 11 2 1 10 9 0 2 16 4 0 9 1 10 9 1 10 9 2
17 13 10 0 9 1 10 9 1 10 9 1 10 9 11 7 11 2
14 1 10 9 2 13 11 13 1 10 9 1 11 11 2
19 11 11 2 7 3 11 2 13 10 9 0 13 1 10 0 9 11 11 2
13 10 9 0 3 0 7 1 10 0 9 16 13 2
22 1 10 9 1 10 9 2 10 9 13 10 9 0 1 2 1 10 15 15 13 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
32 10 9 11 11 13 10 9 1 11 1 11 2 11 7 10 9 13 1 9 1 11 2 16 4 13 3 1 10 9 1 11 2
24 10 9 1 10 9 0 0 13 9 0 1 10 9 1 10 9 7 16 10 9 13 3 0 2
24 10 9 0 13 10 9 0 1 9 7 10 9 1 9 2 1 9 10 9 4 13 9 0 2
56 3 13 0 9 1 10 9 1 10 0 9 3 16 11 13 3 10 9 3 1 10 9 1 2 11 2 11 8 11 11 11 2 2 2 7 3 11 11 11 7 10 11 15 4 13 1 10 9 1 11 16 13 10 0 9 2
11 11 7 11 13 10 0 9 1 10 9 2
24 1 9 1 16 15 15 4 13 3 1 9 0 2 15 3 15 4 13 1 9 1 9 0 2
47 10 9 1 10 11 1 11 11 13 10 9 1 9 1 10 15 1 12 10 11 11 11 2 13 11 11 9 1 10 11 2 13 1 10 9 10 9 1 10 9 1 10 11 1 11 11 2
72 1 15 2 1 10 9 13 1 10 9 1 10 9 1 9 9 12 1 11 2 11 11 2 10 9 1 11 11 2 11 11 7 10 9 11 11 13 16 1 9 0 15 13 10 9 1 10 9 0 1 7 13 10 9 1 10 9 2 13 7 10 9 1 10 9 1 9 13 10 0 11 2
33 13 1 10 9 1 9 1 13 15 1 10 9 1 10 9 1 10 9 7 10 9 1 10 9 1 9 0 13 0 1 11 11 2
48 3 15 13 1 9 0 16 13 10 0 9 7 9 2 1 10 9 3 4 7 13 1 10 9 0 1 13 16 10 9 15 13 1 13 1 10 9 7 15 13 1 13 1 10 2 9 2 2
11 1 9 2 11 13 13 7 3 15 13 2
60 1 10 12 9 2 11 11 13 0 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
46 9 13 2 11 2 1 9 2 7 9 13 1 9 2 9 7 9 2 16 13 2 9 2 1 11 7 10 9 1 11 2 16 1 10 9 1 10 9 15 13 10 9 0 9 2 2
23 10 2 9 1 10 11 2 13 10 9 0 16 13 3 1 10 9 2 9 7 0 9 2
26 3 2 10 9 11 2 11 15 9 1 13 9 1 9 16 13 1 12 8 2 12 8 7 12 8 2
16 10 0 9 2 13 1 9 1 10 12 9 1 11 1 11 2
50 10 9 2 3 3 1 10 9 1 10 9 2 10 9 1 10 11 11 13 10 9 1 10 9 3 3 13 1 10 3 13 10 9 0 1 10 11 11 2 13 1 10 9 1 9 1 10 9 0 2
44 15 0 1 16 1 9 1 10 9 1 9 2 16 13 4 1 9 2 13 0 1 10 0 9 0 2 13 0 9 2 16 13 15 10 9 1 10 9 1 9 1 10 9 2
30 10 9 1 10 9 0 0 1 10 9 0 0 13 3 0 2 13 13 1 10 12 5 1 10 12 5 2 9 2 2
39 10 11 1 11 13 10 9 13 1 10 9 1 10 9 1 11 2 16 13 10 9 1 10 9 1 11 2 11 11 2 11 1 11 7 10 9 1 11 2
35 1 15 15 10 9 3 4 13 0 1 3 13 15 10 9 1 9 0 2 1 9 0 16 13 1 10 9 3 9 1 3 13 3 0 2
39 10 9 13 0 2 16 10 9 1 10 9 1 9 1 9 0 13 9 1 8 0 3 0 7 10 9 1 10 9 2 7 13 9 1 10 9 1 9 2
9 13 10 12 1 10 9 1 11 2
11 3 13 9 1 0 9 1 10 9 8 2
15 1 10 0 9 2 1 9 2 11 11 13 10 3 0 2
28 1 10 9 1 10 9 11 15 13 1 10 2 9 1 9 2 13 1 11 11 2 11 1 11 10 9 0 2
22 15 13 1 11 1 11 2 10 9 0 16 4 13 13 13 10 9 13 1 10 11 2
8 3 15 13 1 9 7 9 2
21 15 13 1 11 2 9 1 10 9 11 1 10 9 1 11 7 9 1 10 11 2
18 11 13 10 9 0 1 12 9 1 9 1 9 0 1 10 9 11 2
13 10 9 1 10 0 9 13 1 10 9 12 9 2
57 10 9 1 10 9 1 10 9 1 10 11 4 13 1 13 1 10 2 9 1 10 9 2 9 1 9 7 9 1 10 9 1 11 11 2 13 1 10 9 7 13 13 3 2 2 13 1 11 11 1 10 12 1 11 1 12 2
30 3 2 1 10 9 10 9 0 4 13 1 10 9 3 7 10 9 1 10 12 9 15 13 0 3 1 10 9 0 2
15 10 9 0 4 13 3 1 10 9 2 15 1 9 0 2
18 15 13 1 9 1 10 0 9 7 15 4 13 10 9 1 10 9 2
21 1 10 9 12 15 13 1 10 11 12 9 1 10 9 1 3 1 12 9 5 2
28 10 9 4 13 1 10 10 9 1 9 2 16 3 10 9 4 13 1 10 9 1 9 0 11 3 11 11 2
36 10 9 1 9 7 10 9 1 4 13 10 9 1 10 9 0 13 4 13 1 3 1 15 2 7 10 9 15 13 0 1 9 1 10 9 2
39 10 9 13 1 0 9 1 10 9 1 10 9 2 1 10 9 0 7 1 13 10 9 1 10 9 2 7 10 0 9 0 13 10 9 1 10 9 0 2
45 1 10 0 9 15 13 10 9 1 10 10 9 13 1 10 11 11 2 15 13 0 9 13 1 10 9 7 10 9 1 3 0 9 2 10 15 4 13 1 10 9 0 1 12 2
55 1 9 2 11 2 0 9 1 10 9 1 10 9 2 3 0 7 0 1 9 1 13 15 1 10 10 9 13 1 10 9 0 1 10 9 2 13 13 10 9 1 10 9 1 10 15 4 1 13 10 0 9 1 12 2
34 15 13 1 10 11 11 7 15 13 1 10 11 11 2 11 2 13 7 13 10 0 9 1 9 0 1 11 13 1 11 1 3 9 2
63 2 10 9 0 11 13 3 1 13 1 10 12 9 10 9 1 11 2 11 2 11 2 11 2 11 7 11 1 10 9 1 10 9 1 9 1 10 9 0 11 7 13 10 9 2 1 10 12 2 10 9 1 15 1 10 11 2 11 7 11 1 11 2
79 3 11 4 13 1 10 0 9 1 11 13 1 10 9 1 9 0 2 10 9 1 10 9 1 10 9 2 7 2 1 10 9 2 13 1 12 9 1 10 9 2 1 10 9 10 9 13 1 13 15 3 3 0 15 13 7 1 10 15 10 9 1 10 15 15 13 3 13 1 10 10 9 13 3 16 15 13 0 2
28 15 15 13 1 10 9 10 9 2 11 2 16 13 1 10 9 1 9 2 9 0 7 9 0 1 10 9 2
45 16 10 9 1 10 9 1 10 9 15 13 1 11 10 9 1 9 1 10 9 2 4 13 1 10 9 0 1 9 1 10 11 1 12 2 2 13 3 1 9 1 13 1 15 2
41 10 9 13 3 0 3 16 2 1 10 9 2 13 10 9 1 10 9 0 1 10 9 7 3 1 13 10 9 0 0 1 10 9 2 13 1 10 9 1 9 2
29 1 10 9 1 9 1 0 9 7 9 2 10 9 4 13 10 9 1 10 9 0 2 1 10 9 10 9 0 2
21 10 9 15 13 1 9 1 10 9 0 1 9 1 9 16 13 1 10 12 9 2
3 12 9 2
9 1 10 9 15 13 10 0 9 2
7 13 1 11 2 11 2 2
24 1 9 1 10 9 16 4 13 0 2 13 13 16 10 9 1 10 9 13 1 10 0 9 2
29 10 9 1 10 12 9 13 10 9 1 9 0 2 1 10 9 13 1 0 9 1 10 11 1 11 2 11 2 2
22 3 4 13 1 10 9 8 2 1 10 9 3 0 7 0 0 1 13 9 1 9 2
38 10 9 1 9 1 11 13 9 10 9 13 1 12 12 12 9 1 9 2 7 15 9 13 16 13 10 9 1 9 1 9 2 0 1 13 1 9 2
15 3 2 13 9 1 10 9 0 1 10 9 1 10 9 2
51 10 9 1 10 11 15 13 1 10 0 9 1 15 16 1 10 9 1 9 15 13 2 1 15 3 0 2 11 2 11 2 11 2 11 2 1 15 3 0 2 11 7 10 9 0 2 11 2 11 2 2
9 3 13 10 9 0 1 0 9 2
8 1 10 9 13 3 1 8 2
28 3 15 13 15 4 4 13 15 1 10 9 1 10 12 9 2 7 15 3 7 15 13 1 11 1 9 0 2
29 16 13 3 1 10 9 2 10 9 15 13 13 1 10 11 1 11 2 13 1 10 9 2 15 3 4 13 11 2
10 2 15 3 13 0 9 2 2 13 2
11 10 9 11 1 11 15 13 1 9 0 2
85 13 16 1 9 1 16 10 9 0 13 10 9 0 7 0 2 2 10 9 11 1 11 1 11 2 1 3 2 11 2 2 4 13 10 9 1 9 0 2 10 9 0 13 10 9 0 2 0 7 0 1 10 9 1 10 9 0 2 1 13 10 9 1 10 9 1 10 9 1 9 0 7 1 9 1 10 9 1 0 7 1 0 9 2 2
5 2 13 10 9 2
8 1 15 2 11 11 15 13 2
24 15 13 16 10 0 9 16 15 13 1 10 9 1 10 9 2 13 10 9 1 10 9 11 2
18 1 11 1 9 2 10 9 1 9 13 10 9 0 1 9 1 9 2
37 1 15 15 13 10 3 3 13 9 1 10 9 2 11 11 2 10 9 11 11 2 11 11 2 11 11 2 11 11 7 11 11 11 2 1 15 2
30 1 16 10 9 0 13 2 4 13 0 9 1 10 9 7 1 10 9 1 9 7 9 7 3 13 7 13 1 9 2
33 13 1 10 9 0 2 10 9 4 13 1 13 9 1 10 9 7 10 9 13 10 9 0 1 9 1 10 0 9 1 11 11 2
35 13 10 9 9 1 9 1 11 2 1 15 13 1 10 0 9 1 12 1 9 2 10 9 1 15 11 11 15 13 10 9 1 11 11 2
24 10 9 15 13 10 12 1 11 1 12 2 1 10 11 11 11 2 1 10 9 5 2 8 2
36 3 0 9 2 15 4 13 16 13 16 13 0 7 10 15 0 7 13 16 13 8 0 7 13 3 0 9 7 9 16 3 13 1 10 9 2
44 10 12 9 0 1 11 15 13 1 11 2 11 2 1 10 12 7 10 12 1 11 1 12 1 10 9 1 10 11 11 1 11 11 2 11 2 7 10 11 11 1 11 11 2
62 11 11 11 2 10 9 13 10 9 1 10 9 0 2 1 9 1 10 9 1 9 12 1 11 1 12 13 16 10 0 9 4 13 1 13 1 10 11 1 11 15 1 3 13 10 11 1 11 1 11 2 1 10 9 1 10 0 9 11 11 11 2
23 10 9 1 11 15 13 1 10 9 1 12 5 7 13 1 10 9 0 13 1 12 5 2
34 4 13 10 9 1 12 7 12 1 10 9 1 11 11 2 11 11 7 1 9 1 11 15 13 10 9 1 11 2 11 11 2 2 2
33 10 9 1 10 9 13 1 10 9 0 8 2 9 5 0 2 7 8 2 8 5 9 2 1 9 1 10 9 0 1 10 9 2
26 1 12 2 13 1 10 9 1 11 11 1 2 11 2 2 2 11 13 9 2 7 2 11 9 2 2
14 10 9 1 10 9 13 0 2 5 7 0 2 5 2
14 1 15 15 13 10 9 1 10 9 1 11 7 11 2
20 11 11 13 10 9 3 0 1 10 12 16 13 10 9 0 1 11 2 11 2
28 1 10 9 13 10 9 1 9 0 2 16 13 1 10 9 10 9 1 13 9 13 1 9 1 10 9 0 2
65 7 13 16 4 1 4 7 13 15 10 9 3 10 15 3 2 3 7 10 9 4 13 16 10 9 1 12 9 2 9 11 11 1 12 8 7 9 0 1 12 8 2 3 13 1 9 1 13 1 10 9 0 10 9 1 11 2 16 1 10 9 15 4 13 2
34 10 9 11 11 4 13 16 10 9 4 13 2 10 9 1 0 16 13 3 12 9 0 1 13 10 9 7 15 13 10 0 9 2 2
30 15 4 13 1 10 9 0 2 1 10 12 9 1 9 15 13 0 1 13 1 10 9 3 1 16 10 9 4 13 2
13 12 9 3 2 15 15 13 1 10 9 1 11 2
10 10 9 1 10 9 13 1 12 9 2
20 15 1 10 9 3 0 13 11 11 11 11 2 12 2 2 13 1 11 11 2
10 1 10 9 0 2 15 13 10 9 2
23 11 2 1 13 15 10 9 1 10 9 2 7 1 10 9 1 11 2 13 10 0 9 2
44 1 10 9 1 10 9 1 10 11 11 2 11 9 12 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
18 15 13 1 10 9 12 5 12 12 8 8 12 5 12 12 8 8 2
23 0 13 10 9 0 7 1 10 9 2 11 13 10 9 0 7 10 0 9 2 15 13 2
15 10 9 0 13 12 5 12 2 8 2 12 5 12 2 8
41 1 10 9 2 10 9 0 13 1 10 9 0 7 13 10 9 1 11 2 3 1 11 2 11 2 2 1 10 15 15 13 10 0 11 12 2 15 3 4 13 2
30 15 4 13 9 1 10 9 2 7 10 9 13 0 1 9 2 1 10 9 16 15 13 1 7 13 10 9 10 9 2
40 13 1 10 12 12 9 2 16 15 13 9 1 10 9 11 11 2 13 2 2 10 11 13 10 0 13 1 9 1 12 1 9 1 11 11 11 7 11 11 2
28 10 9 13 10 11 13 10 9 1 10 9 1 9 2 16 13 1 9 1 10 9 3 0 1 10 9 0 2
34 13 1 9 16 10 9 13 1 10 9 1 11 7 11 2 7 1 9 1 3 13 16 13 10 9 1 10 9 1 10 9 1 9 2
25 1 13 10 12 1 11 1 12 2 11 15 13 1 13 1 10 9 1 10 9 11 1 10 11 2
28 10 0 9 13 10 11 16 15 11 11 2 1 9 11 11 11 11 11 2 2 1 3 13 10 9 1 9 2
17 11 13 10 9 7 10 9 1 10 9 1 11 11 2 11 11 2
20 10 9 15 13 1 11 11 2 7 13 0 1 13 10 9 1 10 11 11 2
12 11 11 13 10 9 1 9 1 10 9 11 2
27 7 1 10 0 9 16 13 4 13 10 9 1 10 9 16 13 1 10 9 2 3 13 16 11 4 13 2
27 10 9 1 10 9 1 11 12 7 11 7 11 13 1 9 10 9 1 9 3 0 13 11 12 7 11 2
50 0 10 12 5 1 10 9 13 1 10 9 0 12 0 9 1 11 7 1 10 9 0 12 1 11 1 11 7 10 12 5 15 13 1 10 9 0 12 11 11 0 7 1 10 9 0 12 11 11 2
16 10 9 1 9 1 10 9 13 2 10 9 1 10 9 2 2
21 15 13 0 1 10 9 0 1 10 9 7 9 0 7 0 1 10 9 1 9 2
16 2 13 16 11 11 1 9 13 10 9 0 1 9 1 9 2
17 10 9 1 10 9 15 13 1 13 10 9 3 11 4 7 13 2
26 1 9 2 10 9 4 13 1 10 9 0 2 3 1 7 10 0 9 3 15 13 1 13 10 9 2
23 11 15 13 10 9 1 11 2 7 13 16 2 16 11 13 1 13 15 1 15 2 13 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
16 11 11 13 1 10 9 0 1 10 9 7 10 9 1 11 2
50 10 9 13 1 10 9 1 10 9 1 10 9 2 3 1 8 7 8 2 13 3 2 13 11 2 3 0 11 2 2 7 10 10 9 16 15 13 0 1 9 2 1 11 2 11 2 11 7 11 2
16 10 9 13 1 9 10 9 1 9 0 7 9 1 10 9 2
35 13 16 3 13 9 0 1 3 13 10 9 1 10 9 7 16 10 9 3 4 4 13 1 9 2 7 1 9 1 9 1 9 1 9 2
68 10 9 1 9 2 11 11 2 13 9 1 9 0 2 10 9 15 13 0 1 13 10 9 15 15 13 16 7 15 7 10 9 9 13 0 1 10 9 2 13 3 2 3 10 9 1 9 9 13 10 9 2 16 13 10 9 2 4 13 15 1 9 1 11 7 11 2 2
26 10 9 1 10 9 1 10 9 1 10 9 4 13 10 9 0 1 10 9 0 9 1 10 9 0 2
25 11 13 10 0 9 1 11 11 1 9 2 13 1 12 2 13 1 9 13 1 11 11 7 9 2
15 3 15 13 9 1 9 7 1 9 0 1 13 10 9 2
33 3 13 10 12 1 10 9 16 15 13 1 11 16 13 2 13 10 0 9 3 13 10 0 9 13 1 13 15 9 1 10 9 2
28 1 9 2 11 12 13 13 10 9 1 2 11 1 10 10 11 2 2 16 1 10 9 10 9 13 1 11 2
20 11 13 13 7 13 13 15 1 11 16 15 13 1 4 13 15 1 0 9 2
51 10 12 1 9 1 10 9 0 13 10 9 0 2 10 12 10 9 2 10 12 10 9 2 10 12 10 9 2 3 1 10 9 1 9 2 10 12 10 9 0 7 3 1 10 12 1 9 10 9 0 2
23 11 11 11 2 12 1 11 1 12 2 13 10 9 3 13 1 10 9 1 11 11 11 2
23 2 4 11 1 10 9 1 11 2 11 10 9 1 9 7 11 10 9 13 1 10 9 2
75 11 1 10 11 2 1 10 13 10 9 0 13 1 10 9 1 10 9 2 9 12 2 13 10 9 0 0 2 1 0 9 0 2 3 13 15 9 1 10 9 2 11 11 1 11 11 2 11 1 11 2 2 9 1 11 11 1 11 7 1 11 11 1 11 2 9 1 10 11 1 11 1 10 11 2
15 3 10 9 1 11 2 11 2 7 1 11 2 11 2 2
24 3 3 4 13 1 10 9 0 7 0 7 13 0 16 15 3 15 4 1 13 1 10 9 2
12 3 13 13 15 1 9 7 1 9 1 13 2
20 10 9 1 10 9 0 15 13 1 15 1 10 9 2 15 13 1 11 11 2
13 10 9 1 10 9 4 13 1 10 0 1 11 2
50 10 9 4 1 12 9 13 2 1 9 0 2 1 9 1 0 9 2 12 1 10 9 9 7 9 7 12 1 10 9 9 2 13 1 9 1 10 9 9 7 9 1 9 1 10 9 15 7 9 2
24 10 10 9 13 9 0 2 1 10 9 0 7 9 0 2 16 13 10 9 1 10 12 5 2
14 7 3 7 15 13 3 2 15 13 10 9 1 11 2
8 13 10 9 0 1 11 11 2
41 10 0 9 13 10 9 0 2 15 4 13 1 10 9 1 3 1 12 5 2 7 10 10 9 4 13 1 10 9 8 12 11 1 10 11 13 3 1 10 9 2
25 1 10 9 15 13 1 9 1 10 9 1 10 9 0 7 13 1 9 0 10 9 1 10 9 2
12 13 9 9 1 8 7 8 13 10 9 9 2
19 3 3 2 11 4 13 7 13 2 13 15 15 1 13 13 1 10 9 2
45 3 15 4 4 1 13 10 9 13 8 9 1 11 2 16 13 10 9 1 10 9 1 11 7 11 2 10 9 11 7 10 9 1 10 11 2 1 10 9 1 9 7 10 11 2
34 11 11 13 10 9 0 1 10 13 12 9 1 9 1 10 9 1 3 2 13 10 1 10 9 1 10 11 2 9 2 11 11 8 2
45 1 10 0 9 2 10 9 1 11 13 10 12 5 1 10 12 9 2 13 1 11 2 10 9 13 10 12 5 7 16 13 3 1 10 12 5 1 10 9 1 10 0 1 9 2
14 10 0 9 1 10 11 2 10 9 11 4 13 3 2
22 10 12 1 11 1 12 13 1 10 9 2 11 2 10 9 1 12 9 1 10 11 2
37 1 0 2 10 9 15 4 13 1 10 11 11 0 7 10 9 0 1 11 2 1 10 16 13 1 9 1 10 12 7 10 12 9 1 10 11 2
16 11 11 13 1 11 1 10 9 1 10 9 0 2 12 5 2
104 15 4 13 10 9 1 11 11 13 1 15 1 10 12 9 0 3 0 1 10 9 1 11 16 1 10 12 1 11 7 1 10 9 1 10 11 1 10 11 15 13 1 9 7 9 2 10 9 1 9 1 10 11 1 11 8 2 9 0 1 11 11 2 11 10 11 3 13 10 9 16 13 1 11 11 1 10 9 2 10 11 1 10 11 7 10 11 1 11 2 1 10 8 2 8 9 1 13 2 10 11 1 11 2
67 1 9 1 10 0 9 7 0 9 7 2 13 16 10 9 13 1 13 15 2 13 10 0 9 1 10 9 2 15 13 1 10 0 9 2 3 15 13 9 10 12 1 11 1 10 11 2 1 12 9 1 10 9 1 10 9 7 13 10 9 1 12 9 1 10 9 2
5 2 9 7 9 2
20 11 11 2 11 2 8 12 2 13 9 1 11 11 2 11 7 3 1 11 2
12 11 13 1 10 9 7 15 13 1 16 13 2
24 10 11 12 13 10 9 3 0 7 1 0 9 1 16 15 13 9 1 12 9 1 12 9 2
35 13 1 10 9 11 2 1 10 9 13 0 1 10 9 1 10 11 7 0 1 10 9 0 11 12 2 16 13 1 9 1 10 9 0 2
19 3 15 13 9 13 1 10 9 0 2 1 11 2 1 11 7 1 11 2
14 1 10 9 1 10 9 15 13 10 9 0 1 9 2
48 15 1 10 0 9 1 9 13 1 9 1 10 12 16 15 13 1 13 10 9 1 11 1 10 9 2 1 11 2 1 11 12 2 11 13 16 13 1 10 9 13 1 10 9 1 9 0 2
14 13 1 9 1 9 2 9 2 9 2 9 7 0 2
26 10 9 4 1 13 1 10 9 0 16 2 3 2 15 13 0 1 13 1 10 11 1 13 10 9 2
24 1 9 1 10 9 13 1 10 11 1 11 11 11 11 2 10 9 4 13 1 15 2 3 2
12 15 13 1 10 11 11 1 10 9 1 11 2
5 2 15 15 13 2
20 1 10 0 12 9 15 13 0 9 1 10 9 1 10 9 7 10 12 9 2
42 10 9 0 15 13 3 1 10 9 1 9 1 10 0 9 1 0 9 2 15 1 10 9 7 10 9 1 10 9 4 3 13 15 1 10 9 0 1 10 9 0 2
21 3 2 15 13 10 9 16 3 15 13 7 15 13 1 10 9 1 9 16 13 2
18 0 9 1 10 9 0 2 10 9 4 4 13 1 3 1 12 9 2
11 10 9 4 13 1 3 1 10 9 0 2
29 1 10 9 10 9 13 1 10 0 9 7 15 13 1 10 9 1 10 9 2 13 15 10 9 1 10 9 0 2
27 10 9 1 0 9 2 13 10 9 0 1 10 9 7 13 15 15 16 15 13 1 13 10 0 9 0 2
6 9 3 0 7 0 2
40 15 13 10 9 0 1 10 9 7 8 7 13 10 9 1 13 2 15 13 3 1 9 1 10 9 0 1 10 16 13 10 9 2 11 11 2 3 3 2 2
18 11 11 4 13 1 11 1 11 11 7 13 1 11 11 12 2 12 2
5 2 15 15 13 2
59 10 9 0 2 1 12 9 7 12 9 1 9 16 13 10 9 0 1 12 7 12 5 2 5 1 9 1 10 9 1 10 8 9 10 12 5 16 13 10 9 1 9 1 10 9 0 4 1 13 10 11 8 1 10 9 1 11 11 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
29 1 9 13 11 2 11 2 11 2 11 11 11 11 11 7 11 11 11 11 1 11 11 11 1 10 9 11 11 2
41 15 13 1 10 9 11 11 2 13 11 1 10 9 11 11 2 11 11 2 11 11 2 11 2 11 2 11 2 11 11 2 11 11 2 11 2 11 11 7 11 2
31 10 9 1 10 9 0 3 0 1 10 9 4 4 1 13 10 9 1 10 9 16 4 13 10 9 0 1 10 0 9 2
45 10 9 7 9 13 1 10 9 1 9 2 15 13 9 7 15 13 9 1 13 15 1 16 13 10 9 7 13 1 15 16 4 1 13 10 9 10 9 7 9 15 4 13 11 2
27 10 9 0 11 7 11 13 1 10 9 12 7 12 1 10 9 0 1 9 1 10 9 1 9 3 0 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
26 11 2 3 13 1 9 0 2 13 10 9 1 10 9 1 16 13 10 9 2 7 10 9 4 13 2
50 10 9 13 9 1 10 9 11 1 11 11 7 11 2 12 9 1 11 1 10 11 2 11 1 11 2 12 9 1 10 11 1 10 11 2 12 9 1 10 11 2 7 1 10 9 11 11 1 11 2
73 11 11 11 11 2 11 2 11 2 12 1 11 1 12 2 11 2 11 2 12 1 11 1 12 2 13 9 1 10 11 1 10 11 1 12 9 1 9 16 13 1 12 1 12 7 12 1 12 2 9 1 9 1 10 11 1 10 11 1 12 7 9 1 10 9 0 0 2 12 2 12 2 2
45 10 9 1 10 9 15 13 1 10 9 9 1 10 9 7 9 1 11 11 11 2 7 10 0 9 13 10 9 1 10 9 2 16 13 1 9 1 11 11 2 1 12 1 12 2
15 15 13 16 10 9 1 10 9 3 3 15 13 15 0 2
7 2 3 15 13 16 13 2
17 11 11 13 10 0 9 1 10 9 1 10 9 1 11 1 11 2
19 10 9 13 1 11 1 11 11 1 10 9 2 13 10 11 1 10 11 2
21 10 9 1 10 0 9 2 1 10 9 1 10 9 11 1 11 2 13 1 12 2
16 10 9 13 10 9 1 10 9 0 2 9 0 1 9 0 2
13 16 15 13 10 0 9 3 13 9 0 7 15 2
53 3 2 15 13 10 9 1 10 9 0 1 13 2 0 2 0 7 8 2 8 1 10 9 0 0 2 7 13 1 10 0 9 1 10 9 0 13 1 13 10 9 16 15 13 3 2 1 9 1 10 0 9 2
42 13 1 10 9 1 11 1 11 10 12 1 11 1 12 2 0 9 1 10 11 1 10 11 1 10 11 11 1 10 9 1 9 2 7 1 10 0 9 1 10 9 2
38 3 15 13 1 3 1 12 9 15 10 9 0 2 11 11 1 11 11 2 2 1 10 9 0 2 9 0 2 2 2 11 0 2 7 2 11 2 2
31 10 9 1 16 10 9 4 13 2 13 1 11 11 1 11 2 3 13 0 9 1 10 9 11 2 0 9 1 9 0 2
46 10 9 3 2 10 9 11 11 13 1 11 1 10 9 11 2 3 13 10 9 1 9 16 3 15 13 1 2 11 11 11 2 2 1 15 15 15 15 13 1 13 9 1 10 9 2
33 1 10 9 1 10 9 2 11 2 1 11 2 1 12 2 15 13 0 13 9 1 12 9 7 4 13 1 15 9 1 10 15 2
69 15 3 13 10 0 9 1 13 1 9 1 10 11 11 2 8 2 7 13 15 1 10 12 9 1 9 1 10 0 9 1 10 11 1 9 1 10 9 1 9 0 1 10 9 13 10 3 1 10 9 0 13 1 10 9 1 10 11 2 3 11 3 13 0 1 13 1 9 2
5 15 13 1 11 11
23 1 13 1 11 4 13 1 10 9 1 11 7 13 3 3 8 1 10 9 13 1 11 2
13 13 9 0 16 13 9 1 9 3 3 13 9 2
27 1 9 2 1 11 15 13 16 10 9 15 13 1 10 9 0 1 9 0 2 1 3 10 9 13 0 2
38 1 10 9 12 10 9 1 10 3 1 10 9 1 9 1 11 10 9 11 11 11 15 13 1 0 9 1 16 13 10 9 1 10 9 0 1 9 2
15 10 9 0 1 10 9 11 1 11 11 13 10 9 0 2
10 15 13 1 10 11 0 9 2 11 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
29 10 10 11 11 11 13 1 11 1 0 7 1 11 1 0 1 10 12 9 1 10 11 2 7 1 11 1 0 2
18 2 13 16 10 9 3 3 13 9 1 10 0 9 2 11 7 11 2
38 10 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 1 11 2 1 2 11 2 1 10 9 1 11 2 11 7 9 1 11 2 11 2
18 2 10 9 4 13 13 10 12 9 1 9 0 7 12 9 1 9 2
6 15 13 1 10 9 2
7 10 9 13 10 9 13 2
25 10 9 13 10 9 2 13 1 9 0 1 16 3 4 4 13 3 1 10 9 13 1 10 9 2
25 1 9 2 10 9 1 11 15 13 1 9 1 10 9 15 4 13 1 10 0 9 1 10 9 2
13 10 9 1 9 13 1 12 8 2 2 5 8 2
41 3 2 11 2 11 7 11 13 10 9 2 16 13 1 9 2 10 11 11 1 10 11 2 2 16 15 4 1 13 1 10 9 1 10 11 11 11 2 1 12 2
34 11 2 16 1 12 9 13 10 3 0 1 10 9 1 11 2 13 10 9 1 9 0 1 10 9 2 16 13 12 9 1 10 9 2
31 1 10 0 9 1 10 9 2 1 10 13 0 1 10 9 1 9 2 15 16 15 13 1 9 13 10 9 1 10 9 2
27 11 3 15 4 13 9 16 13 1 10 9 1 0 7 13 1 10 9 16 13 3 0 1 3 13 0 2
16 1 9 1 9 13 10 9 1 11 1 10 11 11 2 11 2
26 1 0 13 3 0 7 10 9 0 1 11 11 11 2 1 15 15 15 15 13 10 2 9 9 2 2
16 13 10 9 3 15 13 10 0 9 2 1 3 10 12 5 2
30 10 9 0 13 10 0 9 0 2 0 2 1 15 15 10 9 1 10 9 4 0 1 9 1 9 7 9 1 9 2
41 11 11 11 13 10 9 1 9 10 12 1 11 1 12 2 7 3 4 1 13 9 1 11 13 10 12 1 11 1 12 2 13 1 10 9 1 10 9 11 11 2
22 15 13 0 9 2 9 13 1 9 7 15 3 13 10 0 9 1 9 1 10 9 2
36 10 9 15 13 1 10 9 11 11 2 13 1 10 9 1 10 9 1 11 11 2 3 4 13 9 1 10 9 0 0 16 13 1 10 9 2
39 11 11 11 13 10 9 0 0 1 10 11 11 13 1 12 2 1 10 9 1 11 11 10 9 13 7 13 1 10 9 11 2 9 1 10 9 10 11 2
29 16 13 10 11 2 13 0 1 13 3 12 9 1 11 2 9 16 13 3 1 10 11 2 9 1 10 11 11 2
31 11 11 13 1 10 9 0 1 10 9 1 10 9 0 2 10 0 9 0 4 13 7 13 1 9 1 10 11 11 2 2
45 10 9 16 13 1 13 10 8 2 0 2 1 10 9 0 13 9 2 3 7 13 15 13 2 3 15 4 13 10 9 1 10 9 1 13 3 10 9 7 13 15 1 10 9 2
22 10 9 1 11 2 13 2 10 9 1 15 1 10 11 1 11 2 15 11 11 11 2
34 11 11 11 11 2 11 1 11 2 12 2 9 0 16 4 13 10 9 1 11 11 2 10 9 1 10 11 1 11 7 10 9 0 2
42 1 13 15 1 9 0 2 10 9 13 10 0 9 1 9 1 10 9 15 13 2 1 15 15 10 9 0 4 13 15 1 10 9 1 9 0 1 9 7 9 0 2
11 15 15 15 13 1 10 9 0 13 11 2
17 3 2 11 13 10 0 9 1 11 1 4 13 1 10 10 9 2
62 11 13 9 0 1 10 9 1 10 9 0 1 13 1 10 9 1 10 11 1 11 7 15 13 1 12 2 9 1 15 15 13 0 1 13 15 1 11 1 10 3 13 1 10 12 9 2 9 1 9 2 15 13 10 0 9 0 13 12 9 3 2
39 13 10 9 1 10 9 1 11 7 1 10 9 1 9 13 9 7 9 1 10 9 0 1 10 11 2 10 9 1 10 11 7 1 10 9 11 2 11 2
18 10 9 1 11 13 10 9 1 9 10 9 1 9 2 9 7 9 2
29 3 13 16 4 13 10 9 1 13 1 15 2 7 13 16 13 2 2 13 10 9 0 1 10 9 1 10 9 2
32 1 10 9 1 10 9 1 12 2 10 9 0 1 9 1 10 9 13 1 5 12 2 7 10 9 0 1 9 13 5 12 2
31 11 1 10 11 2 1 9 2 11 1 10 11 2 13 10 9 16 13 10 9 9 12 1 10 9 1 11 2 11 2 2
9 11 4 13 10 9 1 10 9 2
24 10 15 1 10 9 15 13 1 9 1 10 9 0 1 9 2 0 2 1 9 0 7 0 2
30 1 9 1 10 9 2 15 4 13 1 10 9 0 0 2 13 1 10 9 1 13 9 3 1 10 9 1 10 9 2
33 10 9 3 13 9 1 10 11 3 0 2 1 10 9 0 7 10 9 0 2 16 15 13 13 10 9 1 10 9 1 10 9 2
15 10 9 13 1 12 9 2 12 9 7 12 9 1 9 2
20 2 11 11 2 11 11 2 13 10 9 13 1 11 11 7 13 1 11 11 2
61 10 9 0 11 11 13 1 10 9 16 10 0 9 15 13 10 9 13 1 10 9 1 10 9 0 2 1 10 9 1 9 1 10 9 16 15 9 16 13 13 13 10 9 0 1 10 9 0 1 10 9 1 10 9 7 9 1 10 9 2 2
30 10 12 1 11 2 11 13 10 0 9 1 10 9 12 1 10 9 16 13 1 10 9 1 10 11 11 1 10 11 2
28 11 2 11 7 11 13 1 9 13 1 10 9 1 10 9 2 3 15 4 13 3 1 10 9 1 10 9 2
33 3 2 1 9 2 3 15 13 10 9 1 10 9 7 9 1 13 15 2 3 4 13 3 9 1 13 10 9 1 13 10 9 2
29 1 15 2 1 10 9 0 15 15 13 2 9 0 2 1 15 16 13 10 9 1 10 9 7 3 1 10 9 2
14 1 10 9 0 10 9 1 11 13 1 10 12 9 2
11 10 9 13 9 1 10 9 1 10 9 2
37 10 0 9 1 10 9 0 1 10 9 4 13 1 9 3 7 13 1 9 1 10 9 11 1 11 7 3 15 4 13 9 0 7 1 0 9 2
76 15 4 4 1 13 10 9 2 1 10 0 9 10 11 13 13 15 10 9 7 1 9 1 10 11 11 3 7 1 10 9 2 10 11 4 1 13 9 2 10 9 7 10 9 1 9 0 15 13 1 11 1 12 1 10 0 9 1 2 10 11 2 10 9 1 10 9 1 10 11 11 11 2 3 11 2
7 13 10 9 0 1 11 2
81 1 9 1 10 9 0 2 10 9 13 1 9 1 9 1 0 9 2 10 9 13 10 9 1 10 9 0 7 10 9 0 0 1 10 0 9 1 10 9 2 7 1 9 1 11 11 11 2 3 10 9 1 10 9 13 9 1 9 0 2 1 10 9 10 9 13 9 0 7 0 1 9 0 1 11 1 10 9 7 11 2
25 10 11 2 16 13 1 10 11 2 12 2 1 12 9 1 11 2 2 3 13 1 13 1 11 2
8 1 10 9 15 3 4 13 2
129 10 9 15 13 10 0 7 0 9 2 10 9 1 10 11 11 2 12 2 2 10 11 1 10 11 11 2 12 2 2 10 11 1 10 11 11 2 12 2 2 10 11 1 10 11 11 2 12 2 2 10 11 1 10 11 11 2 12 2 2 10 11 1 10 11 11 2 12 2 2 10 11 1 10 11 11 2 12 2 7 10 11 1 10 11 11 2 12 2 2 1 3 13 1 9 10 0 9 16 13 3 0 1 10 9 2 13 15 3 1 10 9 2 9 7 9 1 9 3 0 2 0 2 0 7 13 1 11 2
5 10 9 13 13 2
18 10 11 11 11 13 10 9 1 9 1 9 1 9 0 1 10 11 2
32 11 11 13 15 1 10 9 2 16 3 1 13 1 10 9 2 3 13 10 9 2 0 1 10 9 16 13 1 10 9 0 2
11 10 16 15 13 3 1 9 13 10 9 2
35 10 9 1 8 3 4 13 15 1 10 9 2 3 7 4 13 15 1 10 9 0 1 13 9 7 9 1 16 13 10 9 1 1 9 2
24 10 9 4 13 15 1 9 1 0 9 1 10 12 9 7 10 9 13 13 1 9 0 0 2
18 13 9 1 9 1 10 9 1 11 7 9 1 10 11 11 1 11 2
7 9 1 10 9 1 9 2
24 11 13 10 0 7 10 0 1 10 12 9 16 4 1 13 10 9 1 9 1 10 9 11 2
32 10 9 13 1 16 10 11 11 13 0 1 13 10 9 0 1 10 9 2 1 0 9 16 10 9 0 13 1 10 9 0 2
17 15 4 13 1 10 9 2 16 15 4 13 1 10 10 9 0 2
25 10 9 13 13 10 9 0 7 13 15 1 10 9 9 1 10 11 13 13 10 9 1 12 9 2
25 10 9 1 9 0 2 0 7 0 2 7 10 9 1 9 7 9 13 10 0 9 0 1 11 2
11 13 1 16 13 1 10 11 11 0 0 2
8 11 15 13 0 1 10 9 2
39 3 15 13 9 1 9 2 7 7 15 13 1 9 15 16 13 2 15 9 0 16 4 13 2 7 16 3 15 13 10 9 2 13 3 15 13 10 9 2
28 10 9 13 0 1 10 9 2 3 16 10 9 1 11 2 11 7 11 15 13 1 10 9 0 1 10 9 2
17 13 1 10 11 1 11 1 10 11 1 9 1 11 2 10 11 2
20 3 4 7 13 3 13 10 9 2 9 2 16 3 13 16 4 1 13 0 2
31 7 10 9 3 0 13 16 15 4 13 9 1 10 0 9 0 16 4 13 1 9 1 10 9 1 12 5 16 4 13 2
8 1 10 9 15 13 11 11 2
25 13 15 1 10 12 9 1 10 9 7 13 10 9 1 10 9 0 1 10 9 9 1 10 9 2
21 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
21 1 10 12 2 10 2 9 2 15 13 1 10 9 1 11 11 7 13 10 9 2
43 10 0 9 13 10 9 1 10 9 2 13 15 1 10 9 0 1 10 0 9 2 13 16 15 13 2 12 2 2 13 1 10 9 3 0 2 3 1 9 13 1 11 2
15 10 9 1 9 0 13 1 10 9 1 1 12 7 12 2
52 11 15 13 1 3 10 9 1 11 3 13 9 1 10 9 7 13 13 10 11 1 3 13 15 2 16 13 16 11 4 13 15 15 13 7 13 16 10 0 9 3 13 11 2 7 15 16 13 13 10 9 2
22 13 1 10 9 0 0 1 11 2 11 1 12 2 7 13 13 1 10 9 1 12 2
14 13 1 15 1 10 9 7 9 0 1 10 9 13 2
28 1 13 1 10 9 10 9 13 10 9 3 0 7 0 13 15 1 10 9 0 15 4 1 13 1 10 9 2
29 10 0 9 1 11 3 13 1 10 9 2 16 13 1 10 9 1 10 9 10 9 7 10 9 1 10 9 0 2
26 13 16 10 9 4 13 10 9 2 16 4 13 10 9 0 1 13 15 1 10 0 9 1 10 9 2
2 11 11
37 13 1 10 9 2 13 10 9 10 9 1 13 15 1 10 9 2 16 3 13 9 2 3 4 13 10 9 7 7 3 13 10 0 9 1 15 2
15 13 10 0 9 16 15 13 1 10 9 0 1 10 11 2
34 1 10 9 13 16 3 13 10 9 1 10 9 2 9 7 9 2 1 9 1 9 1 10 11 11 2 15 13 1 10 12 9 2 2
17 13 1 0 9 2 10 9 3 0 13 10 9 1 13 10 9 2
16 13 3 3 10 9 1 10 9 0 1 10 9 1 10 11 2
9 13 10 9 1 9 1 11 11 2
35 1 10 0 9 0 2 13 1 12 2 13 10 9 11 11 11 1 15 11 1 10 9 0 11 1 10 12 5 1 10 9 7 12 9 2
38 7 3 1 10 13 15 10 9 0 7 1 9 1 10 9 0 1 10 9 2 10 9 4 13 1 9 0 2 9 1 9 7 1 10 9 0 2 2
14 16 10 9 1 9 13 0 2 10 1 9 15 0 2
14 10 9 13 0 2 16 13 1 3 3 9 1 9 2
16 11 7 11 11 4 13 1 10 9 11 1 13 1 10 11 2
22 3 2 15 1 10 12 9 4 13 9 2 10 9 0 0 2 9 7 10 9 0 2
13 1 10 9 10 9 1 10 9 13 10 9 0 2
23 13 9 1 9 0 7 13 10 9 7 10 9 0 1 10 11 1 11 11 7 10 11 2
18 11 2 15 13 1 9 1 10 9 13 16 3 13 9 1 10 9 2
7 9 11 11 2 12 2 2
25 3 13 15 1 10 9 13 1 11 1 10 9 0 1 11 7 11 1 10 9 1 12 7 12 2
39 1 9 1 10 9 1 9 1 10 9 1 11 2 11 3 13 9 1 13 10 10 9 7 9 15 13 2 1 10 15 13 1 12 1 13 11 1 11 2
24 10 9 1 10 11 13 3 0 2 13 1 15 13 10 9 7 13 10 9 1 13 15 9 2
12 13 0 9 1 11 11 1 10 9 1 11 2
29 10 9 0 13 9 7 9 1 3 1 10 12 9 0 1 10 0 9 1 10 9 1 10 3 1 10 0 11 2
26 10 0 9 1 10 9 2 10 9 13 10 9 1 9 1 10 9 1 15 1 13 15 1 9 0 2
30 10 9 0 13 3 1 10 9 2 1 3 12 9 1 10 9 3 0 2 1 12 9 1 10 9 1 10 11 11 2
23 2 3 15 13 2 2 13 16 13 16 10 9 0 4 13 1 0 1 10 9 1 9 2
23 9 0 1 9 1 9 1 9 0 1 9 2 9 1 9 9 7 9 1 9 1 9 2
12 10 9 4 13 1 10 9 12 2 12 2 2
32 7 2 1 9 1 15 2 13 1 9 10 9 1 9 16 4 1 13 3 1 10 9 1 10 9 1 11 11 7 10 11 2
60 16 4 13 9 1 11 1 10 9 2 15 13 15 1 10 9 0 7 1 10 11 11 2 7 13 15 1 10 9 16 15 4 13 1 10 9 1 10 9 1 10 9 2 1 10 16 4 13 12 9 7 10 9 1 9 0 2 11 11 2
24 10 9 1 9 1 9 13 10 9 1 0 9 1 10 9 16 3 13 9 13 1 10 9 2
13 11 11 13 10 9 1 9 9 1 10 9 11 2
15 1 10 12 13 10 9 1 13 1 10 9 1 10 9 2
23 10 9 0 1 10 9 13 10 9 0 1 10 9 0 2 13 1 9 0 7 9 0 2
40 1 10 9 2 10 9 2 9 1 9 7 9 1 0 9 13 10 9 1 10 15 10 9 13 10 9 1 10 9 1 10 0 9 2 3 13 3 7 3 2
13 10 9 4 13 1 10 9 0 1 11 7 11 2
13 10 11 4 13 1 9 10 12 1 11 1 12 2
22 1 13 15 1 16 15 4 13 2 11 11 13 1 10 9 1 7 13 0 7 0 2
68 10 9 1 10 11 1 11 13 10 9 1 15 1 10 9 1 9 0 2 10 9 1 11 13 10 9 2 7 1 10 13 10 9 0 1 10 9 10 9 16 15 13 3 2 10 9 1 10 9 1 9 4 13 1 10 9 1 10 9 9 2 10 9 1 9 3 0 2
13 2 13 10 9 0 9 1 10 9 1 10 9 2
12 10 9 1 9 13 1 12 9 8 9 5 2
20 15 4 0 7 13 1 10 11 1 11 1 16 4 13 1 10 9 1 9 2
67 10 9 1 16 11 15 4 13 1 10 0 9 0 16 13 10 11 11 11 2 13 15 16 13 1 11 1 13 15 16 3 4 8 2 13 10 9 1 11 7 13 10 1 11 2 7 3 2 16 1 10 9 1 10 9 10 9 1 13 1 11 3 13 13 10 9 2
7 13 9 1 10 9 0 2
22 10 9 13 0 2 10 9 15 13 1 10 9 2 13 10 9 7 10 9 15 13 2
19 15 13 1 10 9 0 7 9 1 9 7 9 1 9 1 9 7 9 2
24 13 15 1 10 12 9 16 13 10 0 9 2 16 3 4 13 9 0 7 12 9 9 0 2
11 10 9 9 13 2 2 11 2 11 2 2
20 11 11 13 10 9 1 9 1 10 9 1 10 11 1 10 9 1 10 11 2
25 10 9 1 10 9 13 3 0 2 3 16 10 12 4 3 13 1 10 8 2 9 1 10 12 2
13 11 11 15 13 10 9 1 11 1 2 0 2 2
10 11 7 11 13 2 7 10 9 13 2
51 1 10 9 12 2 11 11 2 10 9 0 1 10 9 0 1 9 2 9 2 13 8 11 11 2 8 8 9 1 11 2 2 1 9 9 2 9 7 13 10 0 9 1 10 9 1 9 1 10 9 2
5 10 9 13 0 2
43 11 13 1 11 16 13 3 10 9 1 10 9 7 2 1 10 13 15 0 1 13 15 2 11 13 1 13 10 9 1 10 9 1 11 2 13 15 16 15 4 13 9 2
13 10 0 9 1 15 13 9 1 9 0 7 0 2
61 3 2 10 12 1 11 1 12 2 10 12 9 1 10 11 11 1 10 11 2 13 1 12 9 2 13 1 9 10 9 1 10 9 1 11 1 11 2 11 1 11 2 1 16 10 9 0 2 13 1 12 9 2 13 10 11 11 1 10 11 2
18 2 13 10 9 1 9 7 9 2 1 10 0 7 9 7 9 0 2
9 10 9 13 0 2 0 7 0 2
18 1 10 9 1 11 2 11 13 10 0 9 0 1 10 11 1 11 2
64 1 13 10 9 1 9 1 9 2 10 12 9 15 13 1 15 9 1 10 9 0 7 1 10 9 16 13 3 1 10 9 1 10 9 1 12 9 7 15 13 10 9 1 10 9 1 10 15 10 9 1 10 9 0 13 2 15 13 10 0 9 0 2 2
50 1 11 2 1 3 15 13 9 0 1 9 0 3 0 1 10 9 9 7 0 1 10 9 9 7 16 4 13 3 0 1 10 9 1 11 2 9 1 9 7 9 0 0 13 10 15 1 10 9 2
17 16 10 9 13 3 0 3 15 13 9 1 9 1 10 0 9 2
47 1 9 1 16 1 10 9 4 13 12 9 1 10 9 0 2 12 7 12 2 7 10 0 9 1 9 13 1 10 12 0 9 2 3 4 13 10 9 0 3 1 10 9 1 9 0 2
43 11 13 3 1 10 9 3 0 2 1 12 9 2 1 10 16 15 4 13 3 11 7 13 10 9 1 11 2 11 7 10 1 11 2 11 1 11 2 9 1 10 9 2
19 10 9 11 2 13 0 1 10 9 1 11 1 10 9 2 11 7 11 2
13 10 9 16 3 4 13 10 9 1 10 10 9 2
39 10 9 1 10 9 0 0 1 10 0 11 11 1 10 9 0 7 10 9 2 11 11 2 4 13 16 1 10 9 15 13 10 9 1 9 0 1 9 2
12 13 1 10 9 1 9 11 2 13 1 11 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
19 9 0 1 10 9 1 10 9 1 10 11 11 1 10 11 1 10 11 2
20 1 10 9 2 11 13 1 10 9 1 12 2 10 2 9 1 11 11 2 2
22 1 10 12 2 4 13 1 9 1 9 1 10 9 0 2 1 9 1 11 7 11 2
19 15 15 13 1 10 9 1 10 9 0 1 10 9 16 13 10 9 0 2
10 13 15 3 16 3 4 13 0 2 2
14 10 12 9 0 1 10 9 13 9 2 9 7 9 2
51 10 9 15 13 1 10 11 1 10 11 11 5 11 2 7 1 3 2 13 10 9 1 10 9 1 9 13 1 10 9 1 10 9 0 1 11 11 2 1 10 11 1 11 7 1 10 11 11 11 11 2
26 10 9 13 10 12 9 0 2 10 9 13 1 12 5 13 1 10 9 7 15 13 3 7 3 0 2
52 11 11 11 2 1 9 2 11 11 11 2 12 1 11 2 12 1 11 1 10 9 0 2 1 12 2 12 1 11 2 12 1 11 1 10 9 0 2 1 12 2 13 10 9 1 9 7 9 0 2 0 2
29 1 9 13 9 9 7 13 1 10 0 9 1 11 7 1 11 1 10 11 1 10 11 7 10 11 11 2 3 2
23 10 9 0 2 11 11 2 2 3 13 11 2 13 10 9 0 1 10 9 1 10 9 2
21 10 9 1 10 10 9 13 1 10 9 15 13 3 1 10 9 13 10 12 9 2
30 9 0 7 15 0 1 10 9 2 9 3 3 0 2 9 0 7 0 2 7 9 9 0 2 1 15 1 9 0 2
23 2 4 13 1 13 15 1 10 9 1 10 9 0 7 1 13 9 1 10 9 1 9 2
28 1 10 9 0 2 10 9 0 13 10 9 1 9 1 10 9 12 1 10 9 12 2 8 12 1 12 2 2
27 10 0 9 13 10 9 1 10 11 11 7 9 1 10 9 0 1 10 11 2 1 10 9 1 10 11 2
56 3 0 9 13 10 9 1 10 9 0 2 3 15 1 10 9 0 1 15 1 10 9 0 2 1 16 2 9 1 10 9 0 2 16 13 1 9 7 3 1 9 1 11 7 10 9 1 10 11 11 2 15 13 10 9 2
32 10 9 0 7 10 9 1 10 12 9 15 13 16 11 4 13 1 10 9 1 11 7 13 2 0 1 9 2 1 10 9 2
12 1 10 9 2 13 3 10 0 9 7 9 2
11 10 9 1 11 15 13 13 1 10 9 2
36 11 7 11 2 9 1 11 2 13 10 9 0 1 10 10 9 2 13 15 9 1 13 1 13 10 10 9 7 10 9 1 10 9 1 9 2
14 9 0 1 13 7 13 9 7 10 10 9 1 9 2
27 10 9 1 12 9 7 12 9 0 13 1 9 10 9 1 10 9 2 16 15 13 0 3 1 12 9 2
15 1 12 13 1 10 2 0 2 10 0 9 0 7 0 2
19 2 7 10 11 11 13 10 0 9 1 10 9 0 9 12 13 1 12 2
11 10 9 13 0 1 10 9 1 9 11 2
8 10 0 9 13 11 11 11 2
17 11 13 10 9 13 1 10 9 1 11 2 9 1 11 2 11 2
29 10 9 3 4 13 10 9 0 2 1 10 0 7 13 1 10 9 1 13 9 2 13 1 10 9 1 10 9 2
24 10 9 13 10 9 1 9 1 10 9 0 1 10 9 7 9 1 10 9 7 1 10 9 2
9 10 9 13 10 9 1 11 11 2
21 11 3 13 10 0 9 2 7 10 9 13 1 10 3 4 13 10 9 1 11 2
5 3 1 10 9 2
18 10 9 13 10 9 0 1 9 12 9 1 10 9 12 1 10 9 2
41 11 3 3 13 10 9 16 15 13 0 2 7 16 3 13 10 9 2 13 10 9 0 2 13 9 0 7 1 9 2 3 7 13 0 9 0 1 10 9 0 2
6 15 13 1 11 11 2
21 3 2 15 13 16 1 12 15 2 13 10 9 1 3 1 12 12 12 1 9 2
58 10 9 4 13 3 1 11 7 13 10 9 0 1 10 9 1 11 16 2 1 3 0 2 13 10 0 9 1 10 9 2 4 3 1 13 12 9 0 9 2 10 9 11 2 12 2 12 2 7 10 9 11 2 0 9 0 0 2
29 10 9 7 10 9 13 0 1 10 9 2 13 9 1 10 9 7 9 0 9 7 9 2 3 16 15 13 0 2
21 3 13 1 10 9 1 11 7 10 9 13 0 2 7 1 10 0 9 1 9 2
9 3 15 13 1 10 9 12 9 2
23 10 9 13 0 7 13 9 1 9 2 16 13 0 9 1 9 2 9 7 9 1 9 2
7 3 0 1 15 16 13 2
43 15 13 10 12 1 11 1 12 2 1 11 2 15 16 13 9 1 10 0 9 1 10 11 1 10 11 2 1 10 9 1 10 9 11 7 1 10 0 9 1 10 11 2
12 13 0 10 9 1 10 3 9 0 11 11 2
5 13 0 1 11 2
27 15 4 1 13 9 16 10 9 15 13 10 9 1 10 11 1 10 9 1 11 11 2 16 13 12 9 2
26 15 13 1 16 10 9 13 3 0 7 16 13 0 13 2 3 7 13 9 7 13 10 9 7 9 2
30 1 10 9 2 10 0 9 15 13 1 9 9 2 7 1 15 16 13 1 10 9 11 2 4 13 10 9 3 0 2
13 11 13 10 9 0 13 1 11 11 7 11 11 2
13 1 9 2 9 1 10 9 4 4 3 13 3 2
45 13 1 16 15 13 1 10 9 10 4 13 1 9 0 1 11 11 2 10 9 13 16 10 9 9 1 16 13 7 3 10 9 16 15 13 3 13 0 13 15 13 10 9 0 2
18 10 0 9 13 2 11 11 2 13 1 9 1 10 11 11 1 11 2
36 11 15 13 3 1 10 9 2 7 10 9 16 13 1 0 2 7 13 3 2 10 9 1 10 9 1 15 15 13 9 1 9 0 0 2 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
16 10 9 0 1 9 2 9 2 9 7 10 0 9 1 9 2
24 1 10 9 1 10 9 2 11 13 10 9 13 15 10 9 1 10 9 16 13 7 16 13 2
29 1 9 1 10 9 13 1 11 2 10 9 13 10 9 0 1 12 9 1 9 7 4 13 1 10 9 9 0 2
19 1 0 9 15 13 13 1 10 9 16 10 9 0 13 10 9 0 9 2
59 10 0 9 4 13 3 1 10 9 0 1 10 0 9 0 2 7 1 10 13 15 2 15 13 1 10 11 1 11 7 1 10 9 1 10 9 2 9 7 9 1 13 10 0 11 1 10 9 2 9 7 9 10 12 1 11 1 12 2
17 1 10 9 1 10 11 11 2 9 1 9 13 9 0 1 11 2
53 10 9 1 9 1 10 9 7 9 1 10 9 1 10 9 1 0 9 1 10 9 13 1 10 9 1 15 2 3 1 10 9 1 15 2 10 9 3 13 16 3 13 10 9 1 10 9 1 9 1 0 9 2
46 10 9 4 13 1 10 9 1 10 9 11 2 7 10 9 1 10 9 1 10 9 10 9 1 3 1 10 9 13 9 1 3 0 9 7 1 10 9 15 13 1 10 9 1 9 2
79 11 13 9 3 3 0 7 10 10 9 1 10 9 1 9 2 11 7 11 2 15 13 0 9 16 3 13 1 10 9 2 1 9 1 10 9 1 9 1 0 9 1 9 13 1 11 2 16 13 10 9 1 4 13 1 9 0 1 10 9 2 7 1 10 9 1 10 9 16 13 10 9 1 9 1 9 7 9 2
21 15 2 13 1 10 9 0 2 13 1 10 9 1 10 9 10 9 1 0 9 2
21 1 13 1 10 12 9 1 10 11 13 10 9 1 9 1 10 9 0 10 11 2
3 2 13 2
22 15 13 10 9 0 7 0 2 3 7 4 13 10 10 9 10 15 0 1 10 9 2
29 3 2 10 0 9 0 0 1 11 4 13 10 9 16 15 4 13 16 13 10 9 1 10 9 0 1 10 9 2
11 4 13 15 1 11 2 16 3 15 13 2
11 11 3 15 13 1 10 9 0 1 11 2
33 15 13 1 0 9 1 10 11 11 11 1 11 1 12 2 7 4 13 10 12 1 11 1 12 1 5 12 3 1 9 7 9 2
33 10 9 13 1 10 9 2 8 10 9 1 10 9 16 13 2 13 0 16 13 1 15 10 9 1 9 1 10 9 0 7 0 2
19 1 10 9 2 10 9 0 3 4 13 0 1 9 0 7 10 9 0 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
20 1 10 9 1 11 1 12 2 11 13 1 13 10 0 9 1 10 0 9 2
25 9 2 2 11 11 11 7 10 9 0 1 11 11 7 11 8 2 9 0 7 9 1 11 11 2
31 15 13 1 10 9 0 13 15 10 9 0 1 13 10 9 0 2 7 16 1 10 9 15 13 7 13 0 1 0 9 2
51 1 9 2 13 0 10 9 7 9 16 15 13 1 10 9 1 9 1 10 9 1 10 9 2 10 9 2 10 9 1 9 4 4 13 1 10 9 16 15 13 1 10 0 9 1 10 9 11 1 11 2
36 1 13 1 10 9 3 0 2 1 3 2 15 13 9 7 9 1 9 13 2 7 1 15 2 13 10 9 0 0 7 13 1 10 9 0 2
20 13 10 9 1 9 0 7 1 9 0 2 12 5 8 2 12 5 8 2 2
15 10 9 13 10 9 0 1 10 11 1 11 10 9 0 2
17 10 9 13 0 2 0 2 3 3 0 2 1 9 7 9 0 2
16 1 10 9 2 15 13 10 0 11 1 11 1 11 1 12 2
19 10 9 4 13 0 10 9 1 9 15 1 10 9 4 13 1 10 9 2
18 11 10 11 13 10 0 9 16 13 1 10 9 1 11 1 10 12 2
88 1 10 9 2 11 11 11 2 1 10 9 10 9 0 7 10 9 0 1 11 2 9 0 1 9 0 2 13 16 10 0 9 16 15 13 1 10 9 1 10 9 1 10 9 0 1 10 9 13 2 9 1 10 9 7 1 10 9 1 9 2 13 1 10 0 9 2 7 10 9 1 10 9 1 10 9 1 10 9 0 2 16 15 13 1 9 9 2
17 10 11 13 0 1 10 9 3 0 1 15 16 13 10 0 9 2
33 10 9 15 13 10 12 1 11 1 11 2 1 9 1 16 10 12 9 13 0 2 1 15 15 10 9 0 15 13 1 10 9 2
13 11 3 13 10 9 1 10 9 0 13 1 12 2
32 4 7 13 16 1 11 10 9 7 9 1 10 9 0 13 16 10 12 0 9 1 9 0 16 13 1 10 9 13 9 0 2
66 1 10 9 15 13 2 1 12 2 11 11 11 2 9 1 11 10 11 2 2 2 2 2 2 1 13 1 10 9 1 10 9 0 1 10 10 9 2 15 4 13 10 9 2 2 2 1 10 9 1 9 3 7 3 1 10 9 2 9 7 3 0 2 2 2 2
38 1 11 11 11 15 13 1 10 9 1 9 0 2 1 10 9 1 10 9 0 1 10 9 2 16 13 10 9 13 1 9 7 10 9 1 10 9 2
49 13 10 9 1 9 3 0 1 11 2 16 13 12 9 1 9 1 10 9 1 9 1 12 9 1 10 9 0 1 11 7 11 2 1 10 9 1 10 11 1 11 1 11 2 1 10 9 0 2
16 11 11 13 10 12 1 11 1 9 1 11 2 11 2 11 2
13 10 9 1 9 13 1 12 13 2 2 9 8 2
37 10 0 9 2 13 1 0 9 1 10 9 2 13 10 9 0 2 9 2 9 7 9 2 16 13 15 1 10 9 1 9 7 9 7 1 9 2
32 10 9 0 1 9 2 12 2 1 9 3 13 10 9 0 16 13 10 9 7 9 1 10 9 1 10 9 0 2 12 2 2
35 10 9 1 9 1 10 11 11 13 3 1 9 1 13 2 13 1 11 2 3 4 1 13 15 3 15 16 4 13 9 0 1 10 11 2
24 10 9 13 10 9 7 3 13 10 9 0 2 7 7 10 9 0 4 13 1 9 7 9 2
32 10 9 1 10 9 13 16 10 9 3 0 3 13 1 10 9 13 10 12 9 7 16 3 4 13 9 1 9 1 12 9 2
25 10 9 2 3 9 1 11 1 10 9 1 10 11 2 15 13 1 10 9 1 9 1 11 11 2
25 13 3 1 9 1 11 2 13 1 0 1 13 10 9 3 2 7 10 9 1 10 9 13 0 2
22 13 10 9 1 9 2 9 2 9 0 2 9 2 9 2 9 7 9 1 10 9 2
23 10 9 4 7 13 10 9 0 7 9 13 1 9 2 16 13 10 9 1 10 9 0 2
26 10 9 1 9 13 1 10 9 1 10 0 9 0 1 13 10 9 1 10 9 7 13 10 9 0 2
8 1 10 9 3 15 13 9 2
33 10 9 1 10 9 13 1 12 9 13 10 9 1 10 9 2 3 7 11 11 11 13 10 11 11 7 11 1 11 10 11 11 2
24 3 1 15 2 1 11 11 11 2 9 1 9 2 13 3 0 1 10 9 1 10 9 0 2
11 9 1 11 13 10 9 1 10 9 0 2
13 10 9 1 10 0 9 3 13 9 7 3 9 2
39 11 3 13 8 2 8 1 10 9 7 15 13 0 9 7 9 2 1 10 9 2 7 13 1 0 9 15 1 10 9 2 13 13 10 9 8 3 0 2
41 1 9 0 2 10 9 0 13 0 7 1 9 15 13 1 10 9 2 1 10 9 1 10 9 1 11 2 0 1 11 2 11 1 10 11 7 11 11 1 11 2
16 10 9 1 10 9 13 10 12 9 2 0 2 0 2 0 2
16 9 9 0 4 13 1 10 9 3 1 10 9 1 10 11 2
12 10 9 0 1 9 1 10 9 1 10 9 2
39 3 1 13 10 9 13 1 11 1 10 0 9 1 11 1 10 9 1 11 2 1 9 13 1 11 1 10 11 11 7 1 11 2 15 16 3 13 11 2
19 10 9 3 0 7 10 9 0 0 2 1 10 0 7 10 9 1 9 2
46 10 9 1 9 4 13 1 10 9 1 9 2 11 11 2 7 10 9 1 9 0 2 11 11 11 2 7 4 13 1 10 11 1 10 11 11 11 11 2 1 10 11 11 11 11 2
22 1 9 3 13 2 11 4 13 1 9 0 1 10 11 11 1 12 1 13 1 11 2
21 13 3 10 9 1 10 9 0 2 11 11 2 11 11 2 11 11 2 11 11 2
60 10 9 1 10 9 11 11 13 3 0 7 15 1 10 9 2 7 3 4 13 10 9 0 1 9 2 13 1 10 9 0 2 1 10 9 1 9 2 9 0 2 9 1 9 2 9 9 1 9 2 9 0 2 9 0 2 7 10 9 2
8 1 10 9 4 13 10 9 2
13 2 13 3 2 7 2 3 2 3 4 13 2 2
25 10 9 15 13 1 11 2 10 11 11 1 10 9 2 13 10 0 9 1 10 9 1 13 0 2
22 11 2 9 2 11 2 13 10 9 1 10 11 1 11 1 10 11 1 11 1 11 2
26 1 9 0 13 1 9 1 10 0 9 7 1 9 12 9 13 13 1 9 10 0 9 1 10 9 2
14 10 9 1 9 3 4 13 1 10 11 11 11 11 2
28 12 2 10 9 0 2 11 11 2 13 16 10 9 0 1 10 9 2 13 0 1 15 16 15 4 13 2 2
9 3 13 10 9 0 2 1 9 2
5 10 9 13 0 2
22 10 9 1 10 9 0 15 13 1 0 9 1 10 9 1 9 1 9 7 9 0 2
59 1 10 12 9 2 11 13 0 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
18 13 15 3 0 2 16 13 1 10 10 9 1 10 9 1 9 0 2
20 15 1 10 9 13 1 10 0 11 11 7 10 9 3 13 10 9 7 9 2
24 1 11 2 10 9 3 15 13 16 3 15 13 1 13 0 9 16 3 13 15 1 0 9 2
12 3 13 13 9 2 15 15 3 13 3 0 2
15 4 13 1 10 0 9 7 15 13 9 7 9 1 3 2
25 1 10 9 1 9 10 9 1 11 15 13 1 9 2 13 9 1 10 9 7 10 9 4 13 2
25 10 9 1 10 9 4 3 13 1 9 1 10 9 7 9 1 0 9 16 3 13 1 9 0 2
10 4 1 13 10 12 1 11 1 12 2
25 10 0 13 10 9 1 9 1 11 2 9 1 11 11 2 3 13 1 10 9 1 9 11 11 2
24 7 13 16 10 9 1 11 11 1 10 11 11 13 0 2 16 11 15 13 3 3 7 3 2
23 1 10 9 1 10 11 11 13 10 9 1 10 9 7 13 9 0 1 10 9 1 11 2
11 10 9 2 10 9 7 10 9 15 13 2
52 10 9 13 16 10 9 1 10 9 3 13 10 9 1 10 9 1 10 9 1 11 2 7 16 3 15 10 9 15 13 1 13 16 13 1 9 7 13 1 9 1 13 9 1 10 0 9 0 1 10 9 2
42 1 10 11 1 10 11 1 10 11 11 2 11 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 4 1 9 0 7 2 12 5 2 12 5 5 13 9 2
60 10 9 11 11 11 13 1 12 10 9 1 13 10 9 0 1 10 9 2 11 11 11 2 7 11 2 9 1 10 15 11 11 11 11 13 1 12 7 12 2 1 2 10 9 1 10 11 11 2 2 1 10 9 2 11 11 11 2 2 2
29 1 11 1 12 13 2 11 11 2 2 1 11 11 2 7 16 2 11 11 2 15 13 1 11 1 10 0 9 2
25 10 9 1 9 1 9 3 3 13 13 1 10 0 9 1 15 9 1 10 9 0 1 10 9 2
13 15 13 1 10 9 1 10 9 1 10 11 11 2
20 13 1 10 9 7 9 16 15 13 0 1 10 9 1 11 13 10 9 0 2
11 15 13 1 10 9 0 1 11 3 0 2
32 1 9 2 11 13 10 9 1 9 2 3 16 13 10 9 1 10 11 11 10 11 1 10 11 11 0 1 10 9 11 11 2
16 15 13 1 11 2 7 13 16 10 9 15 13 1 12 9 2
27 10 9 4 13 10 9 1 10 12 9 1 9 1 10 9 11 11 7 11 11 2 3 13 1 11 2 2
21 11 11 11 2 12 1 11 1 12 1 11 2 13 10 9 0 16 13 1 9 2
28 16 4 13 1 0 9 1 3 1 12 9 2 13 0 13 16 13 10 9 2 13 9 2 0 9 7 9 2
41 1 10 9 1 10 11 2 0 1 10 9 1 11 2 12 5 1 10 8 9 1 11 1 11 7 12 1 10 9 1 11 2 1 10 9 1 11 1 10 11 2
27 1 10 9 2 10 9 1 9 0 1 11 15 13 1 3 1 10 9 1 15 16 13 3 1 10 9 2
20 10 9 0 1 10 9 4 13 1 10 9 1 10 9 0 2 11 11 2 2
25 10 11 11 1 11 8 2 12 15 13 1 11 1 10 12 7 10 12 1 11 1 10 9 12 2
3 4 13 2
29 10 12 9 16 13 1 10 0 9 13 10 9 1 10 9 1 9 13 1 10 9 1 12 2 13 1 11 11 2
46 10 12 1 11 1 12 13 10 9 1 9 0 1 11 2 7 10 9 1 9 1 11 15 13 7 1 10 9 1 12 9 10 11 2 11 7 10 9 1 10 9 4 13 1 11 2
46 10 9 15 13 1 12 9 0 2 10 9 0 2 12 7 12 9 2 2 10 9 0 2 12 5 2 12 5 2 12 5 2 12 5 2 12 5 7 12 5 9 2 7 9 0 2
28 1 13 1 12 11 15 13 1 10 9 1 10 9 1 9 0 16 3 4 13 1 10 9 1 10 0 9 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
49 10 9 1 10 9 13 3 3 1 10 9 0 2 10 9 1 10 9 0 13 1 10 11 11 11 1 11 2 10 9 4 13 1 10 9 15 13 1 10 9 1 13 3 2 10 0 9 0 2
38 3 1 13 10 9 13 1 10 9 7 15 13 2 1 15 16 15 13 15 0 3 1 15 16 13 9 16 3 13 7 9 1 9 16 4 13 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
46 11 11 11 2 1 9 11 11 11 2 13 10 9 0 1 10 9 11 11 13 1 10 9 2 11 11 2 2 16 13 11 2 11 10 9 2 11 2 11 11 7 11 2 11 11 2
35 10 9 13 13 10 9 0 1 9 0 2 3 16 15 9 4 13 1 10 9 7 9 1 9 2 16 3 13 15 9 16 10 9 2 2
18 10 9 13 10 9 0 1 11 2 7 1 10 9 3 15 13 15 2
24 1 10 0 9 1 10 11 10 11 15 13 2 10 9 10 11 2 9 11 7 9 10 11 2
39 10 9 1 16 1 9 15 13 0 9 1 9 1 9 4 4 13 9 2 1 15 15 10 9 4 4 15 13 1 12 9 0 9 1 12 9 1 11 2
24 11 11 3 13 10 9 1 10 9 13 1 10 9 2 1 15 13 10 9 1 10 9 0 2
30 10 8 11 13 1 10 9 1 10 9 2 16 13 10 9 1 10 9 2 2 7 16 15 13 13 12 9 1 9 2
27 10 9 4 13 1 10 9 0 1 10 3 9 11 11 2 3 16 10 9 11 4 13 1 10 11 11 2
52 10 9 15 13 1 10 9 2 13 16 3 4 13 7 10 9 1 10 9 2 16 13 0 2 0 7 0 2 7 16 10 9 15 4 13 1 13 15 16 15 13 7 16 16 15 13 3 3 16 15 13 2
27 10 9 1 9 1 11 13 1 10 9 10 9 0 2 7 3 13 10 9 16 4 13 1 10 0 9 2
18 10 9 11 13 10 0 9 0 1 10 9 1 10 11 1 11 11 2
14 10 12 5 9 0 4 13 1 12 1 11 1 12 2
22 12 9 1 9 0 2 10 11 13 13 15 1 9 7 10 11 13 1 10 11 11 2
14 11 11 2 8 1 11 2 11 2 13 10 9 0 2
21 10 9 1 10 11 7 1 10 11 3 4 4 13 1 11 11 7 1 11 11 2
37 15 13 1 10 9 1 11 2 11 2 11 11 11 11 2 2 2 2 1 10 11 11 2 11 11 2 3 7 10 9 11 11 1 10 0 9 2
16 3 3 4 13 10 9 2 3 10 9 7 10 9 1 9 2
33 10 12 1 11 1 10 9 13 1 9 2 4 13 3 1 10 9 1 11 1 11 8 5 12 10 9 15 13 0 1 11 11 2
13 10 9 4 13 7 0 9 13 1 11 7 11 2
65 11 3 13 1 10 9 9 1 11 11 2 11 11 1 12 2 7 13 10 9 1 10 9 8 9 11 11 2 1 10 15 3 13 11 11 2 10 11 11 2 2 11 11 2 11 11 2 2 11 11 7 11 11 2 11 11 11 2 2 11 11 7 11 11 2
12 15 13 10 9 0 16 13 1 10 10 9 2
44 7 3 13 10 0 9 1 9 7 11 4 1 13 9 1 13 1 10 11 2 10 9 1 10 9 1 9 1 11 11 2 10 9 1 10 9 1 10 9 4 13 10 9 2
36 10 9 13 1 10 9 1 10 9 2 1 10 9 1 10 9 1 10 9 1 9 1 10 9 2 1 10 9 1 10 9 0 7 0 2 2
41 1 16 13 15 2 1 10 11 1 10 11 4 13 1 12 9 0 2 7 1 10 9 1 15 2 16 13 1 10 9 0 1 10 9 2 11 2 11 7 11 2
20 10 9 13 10 9 7 13 10 9 16 13 16 10 9 13 13 1 10 9 2
27 10 9 1 11 15 13 1 13 9 16 3 13 1 11 7 11 2 1 10 9 1 10 9 1 11 11 2
42 1 11 1 11 13 2 10 11 2 2 10 2 11 2 2 10 2 11 2 2 2 10 11 2 7 2 10 11 2 2 3 0 9 3 13 16 13 7 13 10 9 2
34 10 9 0 1 10 9 3 9 2 11 2 13 3 1 12 5 9 7 10 9 15 13 1 11 7 11 16 1 9 13 1 12 5 9
54 16 10 9 4 13 1 9 0 1 10 9 1 12 2 15 13 1 10 9 1 9 1 10 9 1 9 2 13 10 9 0 10 11 1 11 7 10 9 1 10 9 0 7 10 9 0 2 10 9 16 13 10 9 2
31 16 13 10 9 13 0 13 1 13 10 9 7 13 3 2 7 1 0 13 10 9 16 4 7 13 1 10 13 1 11 2
26 3 2 15 15 13 10 12 1 11 1 12 1 9 0 1 10 9 9 0 1 10 9 1 9 0 2
24 10 9 1 10 9 2 1 12 1 12 2 13 10 9 1 9 7 9 0 1 10 9 0 2
28 10 0 9 13 10 9 0 7 0 1 9 2 13 7 1 10 9 1 10 9 1 9 2 1 9 1 9 2
37 12 9 1 9 1 9 2 1 9 0 2 13 1 10 10 9 0 1 10 9 2 13 10 9 0 1 16 10 9 1 11 11 13 1 10 9 2
35 1 10 9 15 13 10 9 1 9 1 10 16 4 13 15 10 9 1 10 9 2 16 10 9 13 16 15 13 1 9 1 9 1 9 2
29 10 9 1 10 9 13 1 12 2 7 13 3 1 9 13 1 10 9 1 10 9 1 10 9 2 10 15 12 2
21 10 9 1 11 7 11 2 11 11 2 13 10 9 1 9 0 1 10 9 9 2
29 10 9 13 9 1 9 0 2 9 1 12 9 1 9 12 5 1 9 1 9 7 9 2 9 1 9 7 9 2
27 15 13 1 10 9 1 10 9 2 3 1 10 9 1 9 2 7 15 3 13 10 9 13 10 8 5 2
10 13 16 13 3 10 9 7 10 9 2
19 1 9 1 10 9 1 11 11 15 13 10 9 1 11 7 10 11 11 2
21 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
24 10 9 13 1 10 11 7 13 1 10 11 12 2 11 2 12 2 0 7 13 1 9 0 2
83 1 13 10 9 1 11 2 13 9 2 13 9 0 7 13 1 0 9 13 1 11 1 13 10 9 2 15 13 13 1 9 9 1 10 10 9 16 15 13 7 13 1 10 9 0 13 9 0 2 2 10 9 1 10 11 11 2 11 1 11 12 2 13 1 9 11 2 1 11 11 2 11 2 11 7 11 2 4 13 1 10 9 2
12 11 11 13 10 9 1 9 1 10 9 11 2
14 13 10 9 1 12 9 2 11 12 2 1 12 9 2
16 10 9 13 0 7 4 13 16 15 15 13 1 10 9 0 2
36 13 10 12 1 11 1 12 1 11 11 11 11 1 11 2 1 9 1 9 2 13 16 10 9 1 9 15 15 13 13 13 7 13 1 9 2
11 15 13 10 9 1 9 16 4 13 0 2
12 2 9 2 2 1 15 15 13 1 15 2 2
12 10 9 0 16 13 2 13 7 13 10 9 2
21 1 9 1 15 15 15 3 13 2 10 9 9 3 13 9 1 10 9 0 0 2
23 10 9 1 10 9 9 11 12 1 11 13 10 9 1 10 9 16 13 12 9 1 9 2
27 13 10 9 1 12 9 1 10 11 11 11 2 8 2 12 9 0 1 11 2 11 12 1 11 1 12 2
31 3 1 13 10 9 2 10 9 13 1 10 9 11 1 10 9 1 10 9 11 2 3 1 10 0 11 2 12 9 2 2
9 11 11 1 11 2 11 2 12 2
12 1 10 9 3 13 10 9 2 13 1 11 2
76 13 1 10 0 9 0 7 1 10 0 9 1 10 9 11 11 2 4 13 1 11 1 12 2 7 9 0 7 9 1 11 1 10 11 11 2 13 15 10 9 1 13 10 9 1 10 9 0 1 10 9 0 1 10 9 1 9 1 10 0 9 1 10 9 2 13 3 1 10 11 11 1 11 1 12 2
20 13 9 1 9 1 10 9 0 2 7 9 1 9 7 9 1 10 9 0 2
44 10 9 13 1 13 9 9 1 10 9 1 9 2 9 7 9 0 2 1 10 9 1 13 10 9 0 1 10 9 1 10 16 3 1 10 9 1 10 9 13 1 10 9 2
21 10 9 4 13 9 1 10 11 13 16 15 4 13 10 9 13 1 10 0 9 2
58 10 9 13 3 7 1 10 9 1 10 9 0 1 11 15 13 10 9 1 10 11 2 1 15 10 9 13 1 10 9 1 9 7 9 1 16 13 16 10 9 15 13 9 15 15 13 1 13 9 7 13 16 10 9 13 1 13 2
28 1 10 9 1 9 1 12 2 10 9 1 10 9 13 3 1 10 12 5 1 10 9 0 9 2 11 2 2
24 11 0 13 10 9 0 1 9 1 9 2 9 1 10 9 1 10 9 2 13 1 10 11 2
29 10 9 1 0 13 15 3 2 0 7 13 1 10 9 1 10 9 3 4 13 9 0 7 3 10 9 3 13 2
26 16 15 4 13 10 0 9 0 1 10 9 7 10 9 2 13 1 10 9 1 0 9 0 7 0 2
17 1 12 13 10 0 9 0 7 1 12 10 2 11 1 11 2 2
78 13 1 16 10 9 15 4 13 10 9 1 9 15 13 1 10 11 1 10 11 1 9 1 13 15 1 12 9 11 13 10 0 9 1 11 1 9 1 11 11 1 9 0 13 10 9 0 10 9 4 13 1 10 9 12 1 10 9 13 3 10 0 9 0 7 3 10 9 13 11 11 9 1 11 1 12 9 2
28 1 10 9 1 10 9 2 10 9 1 9 0 7 10 9 1 9 15 4 13 0 1 9 1 13 10 9 2
9 15 13 13 1 10 9 1 11 2
52 10 9 16 13 10 9 1 9 2 9 1 10 9 13 1 11 7 11 2 4 13 10 9 1 9 1 10 9 1 10 9 1 12 9 2 3 10 9 1 12 9 1 10 9 1 16 10 9 13 12 9 2
10 10 9 13 7 15 13 15 1 15 2
43 13 10 9 1 10 0 9 13 1 10 9 2 3 13 9 0 2 0 2 0 2 0 7 0 2 10 9 1 10 9 7 10 0 9 1 10 9 13 10 0 9 0 2
37 1 11 15 15 13 3 1 10 9 1 0 9 2 0 15 1 13 15 1 10 9 1 10 9 2 1 10 9 0 7 1 10 9 0 1 9 2
15 10 9 15 13 11 2 7 10 0 2 8 2 13 0 2
28 10 11 4 4 13 1 9 1 15 1 10 11 11 7 10 11 11 2 13 1 9 1 11 7 11 11 3 2
10 9 1 9 2 12 8 2 9 8 2
43 10 9 15 13 0 1 10 12 7 12 9 1 11 11 10 0 9 1 10 10 9 2 7 1 12 9 1 10 9 0 3 0 2 10 2 11 2 11 11 11 11 11 2
7 2 10 9 4 13 9 2
19 10 9 2 11 2 1 11 13 3 2 13 2 15 16 13 10 9 2 2
42 1 9 2 13 13 1 10 9 2 11 11 2 11 11 2 2 0 2 7 0 2 16 1 0 9 13 1 9 1 9 7 1 9 1 9 13 9 1 3 13 15 2
35 3 3 15 13 1 16 10 9 0 2 1 10 13 10 9 1 9 1 10 9 2 4 13 2 2 3 13 3 16 13 9 1 10 9 2
18 12 5 13 1 9 0 2 12 5 0 2 12 5 0 7 12 5 0
10 12 5 1 10 9 13 9 1 9 2
16 10 9 0 3 4 1 10 9 7 10 9 1 9 1 9 2
62 1 10 9 0 13 3 12 9 2 10 11 11 13 10 9 1 12 9 16 13 10 9 2 10 9 7 10 9 1 10 9 16 2 13 10 9 0 2 13 2 13 15 2 1 10 9 16 2 1 10 0 9 2 15 13 1 4 13 1 10 9 2
13 13 3 0 15 10 9 13 0 9 1 10 9 2
17 10 9 13 9 1 11 1 11 2 15 13 13 1 9 1 11 2
14 10 9 1 10 9 13 1 9 10 9 1 10 9 2
49 11 11 11 2 13 10 9 2 9 7 0 0 2 9 1 10 9 0 11 2 9 1 10 11 1 10 11 1 11 1 10 9 1 11 1 10 12 0 9 1 10 9 0 13 1 11 11 11 2
24 13 9 1 10 11 11 1 11 11 2 9 7 0 2 1 10 15 13 9 1 12 7 12 2
30 1 10 9 2 10 9 4 13 2 1 15 1 10 9 1 11 2 9 1 9 1 9 7 0 9 1 9 1 9 2
21 3 3 13 10 9 2 7 0 2 9 1 10 9 0 7 10 9 1 10 9 2
12 1 13 10 9 11 15 13 2 7 11 3 2
20 10 9 13 13 3 10 9 0 13 1 10 9 1 10 15 15 13 10 9 2
13 1 10 9 4 13 1 10 9 7 13 1 11 2
15 9 2 9 7 10 9 0 13 0 2 7 13 1 9 2
21 3 10 9 13 9 1 9 5 2 0 1 10 9 0 8 7 8 2 9 2 2
13 1 12 13 1 10 11 1 10 11 7 10 11 2
14 3 15 13 9 1 9 2 3 13 10 9 16 13 2
27 3 1 10 13 1 10 9 15 13 10 9 2 13 12 9 7 12 16 3 13 2 1 10 9 13 11 2
15 10 9 3 0 2 8 0 2 10 9 11 2 10 9 2
14 10 0 9 4 13 16 2 10 9 4 3 13 2 2
24 10 9 13 3 1 16 10 9 13 0 9 2 7 10 9 1 11 15 13 1 16 13 9 2
17 11 2 10 9 2 10 9 2 7 10 9 15 13 3 0 2 2
37 1 15 2 13 15 1 9 2 9 7 1 15 9 2 1 15 16 13 13 15 10 0 9 2 7 3 13 9 1 10 0 9 1 10 9 0 2
18 11 7 11 13 13 10 9 1 9 1 10 13 11 1 9 1 11 2
11 10 9 13 10 9 0 1 12 12 9 2
13 11 13 10 9 2 13 1 11 1 10 0 9 2
36 1 10 9 1 10 9 2 10 9 1 10 11 13 3 0 10 9 1 10 9 1 11 16 13 10 9 7 3 10 9 1 11 13 10 9 2
16 10 9 0 11 13 10 9 1 9 0 16 13 10 9 0 2
25 13 0 10 9 16 10 9 0 3 13 7 1 11 1 12 10 9 13 0 2 1 10 9 0 2
37 10 9 4 13 1 10 9 0 9 16 13 2 12 9 2 2 13 1 16 1 10 9 1 10 11 13 12 0 9 0 7 0 16 4 13 9 2
17 15 13 10 9 11 1 10 9 0 2 16 3 13 1 10 9 2
12 13 9 16 13 9 7 13 9 16 13 9 2
30 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2 11 2
16 10 9 1 10 9 3 13 3 0 9 1 11 1 15 13 2
5 13 3 10 9 2
31 13 4 16 10 9 1 9 3 13 15 0 7 15 3 13 1 9 2 1 15 9 16 4 13 13 1 10 9 1 9 2
26 10 12 9 1 11 13 1 10 9 1 10 9 2 15 4 13 1 13 1 10 9 1 10 11 11 2
43 1 10 9 1 10 9 0 2 10 9 1 9 1 10 0 9 11 13 1 10 9 11 4 13 1 10 9 11 11 11 2 10 0 9 16 4 13 10 9 8 2 0 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
29 10 9 1 11 11 2 1 9 2 11 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
10 10 11 1 11 3 13 1 11 11 2
33 10 9 1 10 10 9 4 13 1 10 9 1 11 2 11 2 7 3 13 1 10 9 10 9 2 10 9 11 7 10 0 9 2
37 16 10 9 0 15 13 7 13 0 15 13 10 9 1 11 3 16 2 16 10 16 15 13 7 13 13 10 9 15 13 10 9 1 11 2 11 2
21 1 12 1 12 13 12 9 1 11 2 3 13 10 9 1 9 2 3 10 9 2
15 1 10 0 9 13 1 10 9 2 11 11 11 11 2 2
30 3 2 3 1 10 9 0 1 10 9 2 11 13 1 10 9 7 1 10 9 2 15 13 1 10 9 1 10 9 2
20 13 1 9 12 9 2 12 9 7 12 9 2 1 12 9 0 1 10 11 2
4 2 15 13 2
35 10 9 1 10 9 13 13 10 9 1 10 9 1 10 16 13 10 9 1 11 1 10 0 9 1 7 10 9 4 13 9 1 10 9 2
31 10 0 9 13 10 9 1 10 0 9 1 10 9 12 1 10 15 10 11 11 1 11 15 13 10 9 1 10 11 11 2
72 10 9 13 3 13 1 11 1 0 9 7 9 1 10 9 1 9 2 7 1 10 9 2 1 0 1 10 9 0 1 10 0 9 0 2 9 2 7 10 0 9 0 7 1 9 1 10 9 1 12 2 10 9 0 1 15 13 0 1 11 11 1 10 9 2 10 9 7 10 0 9 2
26 10 9 7 9 3 15 13 2 1 9 16 13 1 10 9 10 9 0 13 7 1 11 7 1 11 2
8 4 13 15 1 10 9 0 2
35 1 11 1 10 12 10 9 12 1 11 13 12 9 1 10 9 2 10 12 5 1 10 9 13 1 9 0 2 10 12 5 13 9 0 2
54 13 10 9 16 13 1 0 10 0 9 1 9 1 10 9 1 12 2 1 10 16 10 9 11 11 4 7 4 1 13 1 10 9 1 10 9 1 10 9 1 10 9 1 10 13 1 10 9 1 10 9 1 9 2
15 15 13 3 8 7 11 10 9 13 3 3 0 7 0 2
12 10 9 1 10 9 13 10 9 1 11 11 2
33 2 13 15 15 9 1 9 13 1 9 2 15 4 1 16 3 15 13 10 9 0 1 10 11 2 7 3 10 1 10 9 2 2
37 10 9 15 13 16 1 10 11 15 4 13 1 13 10 9 7 10 9 3 7 4 13 9 7 3 15 13 2 7 16 9 1 15 3 4 13 2
49 10 9 1 9 1 10 9 0 15 13 9 1 10 9 1 10 9 1 10 9 11 2 3 16 16 11 13 10 9 1 10 10 9 1 11 2 15 13 0 13 1 10 9 3 0 1 10 9 2
10 13 9 0 1 13 1 15 1 15 2
11 3 13 10 9 16 7 10 9 15 13 2
29 10 9 0 1 9 13 1 11 10 12 9 0 2 15 16 13 10 12 1 12 3 9 1 10 0 9 1 12 2
35 1 9 1 10 9 12 7 9 1 10 12 13 10 0 9 1 10 9 1 9 0 1 10 10 9 2 15 16 13 10 9 1 9 0 2
25 13 10 9 1 10 9 0 1 4 13 10 9 1 10 0 9 7 10 9 13 11 7 11 11 2
28 1 10 9 1 10 9 1 10 9 12 2 1 10 9 12 2 10 9 11 13 10 9 3 0 1 10 9 2
28 10 9 0 15 4 13 1 10 0 9 1 10 9 1 10 9 2 15 4 13 1 11 11 7 13 1 12 2
36 10 9 1 11 0 2 1 10 9 1 11 13 0 1 11 2 7 13 10 9 1 10 9 10 2 1 16 15 13 10 0 9 1 10 9 2
42 1 10 9 12 13 12 9 2 10 11 0 1 11 7 10 9 1 10 9 1 11 2 3 15 13 16 2 3 2 10 10 9 0 13 10 7 10 9 1 9 0 2
8 9 2 11 11 11 2 11 11
59 1 10 12 9 2 11 13 0 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
31 13 1 10 9 1 9 15 10 9 0 11 11 11 13 10 9 1 10 11 11 1 11 1 11 11 1 10 11 2 11 2
11 3 13 0 9 1 9 1 9 1 9 2
28 10 9 0 1 10 9 2 11 2 13 15 1 10 0 7 3 0 9 1 9 0 1 10 9 11 1 11 2
34 11 11 3 3 4 13 10 9 1 10 9 1 10 11 11 11 8 2 13 16 1 11 3 13 0 1 13 1 10 9 1 3 3 2
23 3 2 15 13 10 9 0 1 10 9 7 9 1 10 9 9 1 10 9 1 10 9 2
32 8 13 10 11 11 2 1 11 2 11 2 7 11 2 11 2 2 1 15 9 1 10 15 15 13 10 9 1 11 7 11 2
20 1 9 10 9 0 1 10 9 3 15 13 3 0 4 13 1 11 1 12 2
17 10 9 13 13 9 1 0 9 2 1 3 13 15 1 10 9 2
29 1 0 2 10 9 1 9 1 10 9 0 15 13 1 10 9 1 10 9 0 1 0 7 10 9 1 10 9 2
23 11 13 10 9 2 0 2 2 10 9 15 13 3 7 11 8 15 13 1 10 11 11 2
17 10 9 11 13 1 10 9 1 12 2 3 7 4 13 1 11 2
27 11 11 2 11 7 11 13 0 1 10 9 1 9 7 13 1 16 10 10 9 13 1 10 9 1 15 2
28 11 13 10 9 2 15 13 1 0 7 1 11 1 12 15 13 1 10 11 11 11 11 2 1 10 11 11 2
25 15 13 1 10 9 13 1 10 9 0 2 3 13 1 10 0 9 1 10 9 1 12 7 12 2
37 10 9 13 1 13 0 9 1 10 9 2 1 10 9 2 9 2 9 2 9 2 9 2 9 2 9 2 1 10 15 3 13 9 1 0 9 2
14 10 9 2 10 9 7 10 9 13 1 10 0 9 2
51 10 11 11 3 13 3 12 9 1 9 1 10 9 1 11 11 1 13 3 3 0 7 15 13 1 16 10 0 9 13 10 11 1 11 2 7 15 3 13 1 10 12 9 2 10 9 1 10 9 0 2
16 3 13 7 9 1 15 16 13 10 9 7 10 9 1 9 2
46 11 13 1 9 1 10 9 1 11 10 12 1 11 1 12 1 10 9 0 13 1 10 9 1 11 3 1 10 9 0 1 11 2 1 10 15 10 9 0 13 0 1 12 1 12 2
40 10 9 1 10 9 13 9 13 1 13 1 10 9 2 10 9 13 2 11 1 10 9 2 11 1 11 1 10 9 2 11 11 1 9 7 11 1 10 9 2
60 10 0 9 0 1 9 13 10 9 7 13 9 1 10 9 0 2 13 1 9 1 9 7 9 2 13 1 10 9 1 9 16 15 13 1 10 9 0 2 13 1 9 1 10 9 7 13 1 9 7 9 1 9 1 10 15 1 10 9 2
18 13 13 1 10 9 10 12 1 11 1 10 0 9 1 3 12 9 2
43 13 10 9 11 2 11 7 11 2 10 15 1 11 2 7 10 9 1 9 2 10 9 7 10 9 1 10 11 1 11 2 3 7 10 9 0 1 11 2 10 2 11 2
12 15 13 9 16 10 9 13 13 1 10 9 2
34 10 9 4 13 3 10 0 9 1 13 10 9 1 13 11 11 1 11 2 1 7 15 4 13 1 10 9 11 11 16 13 10 9 2
25 3 13 1 10 9 1 10 9 0 0 2 13 16 10 9 13 0 1 13 10 9 0 3 0 2
38 1 10 9 2 1 10 9 1 10 11 13 1 10 9 1 10 11 7 15 13 10 9 16 13 15 1 10 9 1 11 2 1 10 9 1 10 9 2
3 9 0 2
26 7 3 9 1 10 9 3 13 10 9 2 9 0 1 11 13 1 11 1 15 9 16 13 1 9 2
26 10 9 13 0 2 10 9 13 0 2 10 9 13 1 15 3 9 16 13 7 3 10 9 13 0 2
20 11 11 13 10 9 0 2 13 1 11 2 11 2 10 12 1 11 1 12 2
35 3 2 13 10 9 0 1 10 9 0 2 10 9 1 9 2 13 1 12 2 7 13 10 0 9 0 1 13 12 9 9 1 10 9 2
35 13 1 10 9 0 13 10 9 1 10 9 1 13 1 11 2 1 11 1 12 2 7 10 9 4 13 1 10 0 9 1 10 9 0 2
13 1 10 0 9 3 15 13 10 9 1 9 0 2
16 12 9 4 13 2 15 1 9 0 7 9 1 9 3 0 2
19 10 9 13 10 9 1 10 9 1 10 9 0 2 3 10 9 1 9 2
44 10 11 15 13 1 10 9 0 1 9 15 16 13 10 9 1 10 9 1 9 7 10 9 3 0 1 10 9 0 7 10 9 0 15 13 10 9 1 11 1 10 9 0 2
50 1 10 9 1 10 9 2 3 0 1 10 11 2 13 10 9 1 10 9 1 11 2 15 13 0 1 10 9 1 10 9 2 7 13 1 10 9 11 2 9 1 10 11 2 7 1 10 12 0 2
25 13 10 9 0 1 9 1 10 15 10 9 4 13 1 10 9 7 10 9 1 3 15 4 13 2
15 13 1 10 9 1 10 9 0 1 11 11 1 10 11 2
4 11 11 13 2
13 10 9 1 9 13 1 12 9 2 2 5 5 2
16 11 11 15 13 10 9 2 3 10 9 7 9 1 10 9 2
46 3 2 1 11 1 12 2 10 0 9 1 10 9 1 11 13 13 15 9 0 1 10 11 11 11 1 10 11 1 11 7 11 2 13 1 10 9 10 0 9 0 1 10 9 0 2
65 9 0 7 0 2 9 7 9 2 9 0 1 10 9 0 7 1 10 9 0 2 15 15 13 1 10 9 0 7 13 16 10 9 0 1 8 2 7 1 15 15 10 9 1 10 9 8 2 13 11 2 2 9 1 10 9 2 13 0 2 13 2 13 2 2
41 13 10 0 9 1 9 2 1 9 1 9 2 1 9 1 9 2 1 9 2 1 10 9 12 1 10 12 2 13 2 1 9 7 1 9 1 9 2 1 11 2
90 1 3 1 10 9 2 10 9 13 3 0 2 10 9 13 3 0 7 9 2 10 9 1 9 0 2 7 13 2 7 13 2 1 10 13 1 10 9 2 13 16 4 13 10 9 7 3 10 9 13 1 10 9 1 10 9 1 10 9 2 3 13 10 9 13 7 13 9 7 16 15 13 10 9 2 3 15 13 13 1 16 3 13 1 13 7 13 10 9 2
36 15 13 1 9 1 10 9 0 2 13 1 10 11 0 1 11 11 11 7 11 11 1 11 2 13 10 12 1 11 1 12 16 13 10 9 2
34 1 10 9 1 13 10 9 1 10 9 0 2 7 1 15 16 13 9 1 9 0 2 2 15 13 9 13 1 9 0 1 0 9 2
12 10 9 1 9 13 1 12 9 1 9 0 2
35 11 2 9 2 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
40 15 13 9 1 10 9 1 12 9 1 10 9 1 10 11 11 1 13 9 1 10 9 0 1 10 9 0 1 10 9 1 11 7 10 9 1 10 9 0 2
37 10 9 4 13 3 1 9 1 10 9 1 10 9 0 2 7 16 10 9 16 13 1 9 1 10 9 0 9 4 13 1 10 9 1 10 9 2
13 1 12 15 13 10 9 9 1 9 11 2 11 2
36 11 1 11 2 11 1 11 1 9 2 13 10 9 0 1 10 9 1 11 0 1 10 9 1 10 11 7 1 10 9 0 1 11 2 11 2
23 13 10 9 1 9 16 13 10 9 2 7 13 1 9 10 0 9 1 9 1 10 9 2
17 15 1 10 9 13 15 1 10 12 9 1 10 9 11 2 11 2
20 11 10 11 7 10 11 2 13 1 10 9 7 9 0 1 10 9 11 11 2
51 1 12 9 10 11 8 2 12 13 1 10 9 1 10 9 0 0 1 10 0 9 9 8 1 10 9 0 0 1 16 4 13 10 12 1 11 1 12 1 10 9 1 10 15 15 13 1 10 9 0 2
16 11 13 10 9 1 10 9 1 11 1 11 1 0 11 11 2
23 1 15 16 1 10 9 15 13 2 10 9 1 12 9 13 0 7 15 1 12 13 0 2
25 10 9 1 9 1 9 0 13 1 12 2 16 15 4 1 13 10 9 1 10 11 3 1 11 2
32 10 9 13 16 10 9 13 1 9 1 9 2 13 15 1 10 9 1 9 0 7 1 9 3 13 1 10 9 1 10 9 2
60 10 9 0 13 10 9 1 9 7 9 2 1 3 3 12 9 2 3 16 10 9 0 13 10 9 2 16 15 13 10 9 0 7 10 9 1 10 9 1 10 9 3 15 13 1 10 10 9 13 1 10 9 2 16 13 1 10 9 0 2
19 10 9 2 9 1 10 9 11 11 2 13 10 9 1 9 1 9 0 2
6 11 11 2 9 0 2
40 3 13 13 15 15 3 7 10 0 9 1 11 7 3 15 13 1 15 1 13 10 9 2 16 13 13 1 11 7 13 15 1 10 9 1 10 15 13 15 2
20 1 10 9 0 13 0 13 16 15 15 13 9 1 10 9 0 1 10 11 2
38 10 10 9 1 10 9 1 10 9 4 4 13 1 10 9 0 0 2 3 2 1 0 2 1 10 12 0 9 1 9 10 9 4 13 1 10 9 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
22 1 15 2 13 1 10 9 13 10 9 1 10 9 2 3 7 13 10 9 0 13 2
54 3 3 7 3 13 10 9 1 10 9 1 9 1 9 2 10 9 1 9 2 1 10 9 0 2 13 10 9 0 2 10 9 4 13 1 11 7 10 9 1 10 9 0 2 1 10 10 9 7 15 1 10 9 2
23 13 10 9 0 2 0 2 3 0 2 16 13 10 9 0 7 16 11 13 13 10 9 2
17 10 9 9 4 4 13 3 1 3 0 3 1 10 9 2 0 2
58 10 12 1 11 1 12 13 10 0 9 2 11 2 2 13 1 10 9 1 0 9 1 13 15 1 10 9 1 10 9 7 1 10 9 1 10 9 2 2 13 10 9 1 9 7 13 1 10 9 1 10 9 1 10 9 1 9 2
10 10 0 9 13 1 9 10 9 0 2
20 3 2 10 9 1 12 9 11 4 13 1 10 9 1 9 0 11 2 5 2
14 1 9 1 9 15 13 15 1 10 0 9 1 11 2
20 1 10 9 7 1 10 9 1 13 13 3 1 10 9 1 10 11 11 11 2
35 10 12 1 11 1 12 15 13 10 9 1 9 7 9 1 15 1 9 1 11 7 11 11 1 11 1 15 16 15 13 10 9 1 11 2
38 1 12 4 1 13 1 10 11 1 11 11 2 13 15 10 9 3 1 10 9 1 10 11 1 10 13 15 1 10 9 10 11 11 1 11 1 12 2
31 11 13 10 9 1 10 9 7 15 1 10 9 13 10 9 2 10 15 4 13 0 2 16 3 13 0 15 13 10 9 2
37 1 10 12 0 9 1 10 9 1 15 13 10 9 2 10 9 11 11 13 12 5 2 11 12 5 7 11 4 13 1 9 1 10 12 5 9 2
47 10 9 0 4 13 1 12 0 9 2 10 9 7 9 1 9 2 16 15 13 1 10 9 0 2 9 7 9 16 13 10 9 2 7 10 9 7 9 1 9 16 13 1 10 9 0 2
16 10 9 1 3 9 13 15 1 11 2 11 7 11 2 11 2
15 16 3 13 2 13 1 10 9 1 10 9 1 11 11 2
18 10 9 13 16 10 12 5 13 1 9 1 9 7 12 5 1 15 2
21 11 11 2 11 2 9 1 11 11 2 12 1 11 1 12 2 13 10 9 0 2
20 11 13 10 9 1 0 9 1 9 2 9 7 9 1 10 0 9 1 11 2
9 0 1 11 2 13 3 1 9 2
15 3 2 1 11 12 2 11 13 10 12 9 1 10 9 2
34 1 3 1 12 9 1 9 0 16 13 11 11 0 1 9 1 9 2 11 11 13 10 9 0 13 1 9 1 9 1 9 7 9 2
26 11 4 13 13 9 0 1 10 9 7 10 9 1 11 3 13 13 1 10 9 10 9 1 10 9 2
25 2 1 10 9 13 1 10 9 1 9 1 11 11 2 16 13 10 9 1 9 1 9 0 2 2
57 3 13 10 9 1 12 7 12 2 10 9 1 12 13 3 0 2 16 15 1 12 3 15 15 13 3 2 3 0 13 10 9 1 9 7 13 15 9 1 9 13 15 1 11 1 12 1 11 12 2 7 13 0 16 4 13 2
23 3 16 13 1 10 9 1 10 11 11 2 10 9 13 1 4 13 1 10 9 1 9 2
40 3 2 10 9 13 3 1 15 9 7 9 2 7 13 10 0 9 1 9 7 10 9 1 10 9 2 16 13 10 9 1 15 16 15 13 1 10 11 11 2
17 10 9 13 9 7 3 13 1 10 11 12 1 10 0 9 0 2
28 1 10 9 10 9 11 13 10 9 1 10 9 2 15 13 3 3 1 10 9 1 11 7 13 1 10 9 2
18 10 9 13 3 13 1 10 9 1 9 2 15 13 1 13 10 9 2
18 10 9 13 1 10 9 1 10 9 7 13 9 0 1 9 1 9 2
13 13 15 1 10 9 0 3 0 1 10 12 8 2
5 11 4 13 11 2
33 10 9 13 1 13 1 11 13 11 2 1 10 0 16 1 11 7 11 11 2 10 15 3 15 13 1 13 10 9 1 11 11 2
14 15 4 13 1 10 9 0 1 10 9 0 2 0 2
28 3 1 10 9 7 9 0 11 11 11 2 13 0 9 7 9 1 10 0 9 1 10 9 1 10 9 0 2
16 11 11 13 10 0 9 1 10 9 0 1 10 9 1 11 2
33 15 13 16 10 0 11 11 15 13 9 1 16 13 10 9 0 1 10 15 11 3 4 13 10 9 10 9 15 4 13 10 9 2
21 10 9 1 9 1 11 1 3 1 9 4 13 15 1 10 11 1 10 9 12 2
23 3 4 13 1 9 0 1 10 11 2 11 1 11 11 2 11 7 11 7 10 11 11 2
29 1 10 12 9 1 9 15 13 10 9 1 9 1 3 12 9 1 9 16 13 13 1 9 0 10 9 3 9 2
11 11 16 13 16 4 1 13 10 0 9 2
12 1 9 2 16 13 10 9 10 9 13 0 2
48 13 10 9 2 10 9 1 10 9 7 10 9 1 10 11 2 10 9 13 1 9 0 1 10 9 7 1 10 2 9 2 1 10 9 7 1 10 9 1 11 1 10 9 0 1 10 9 2
15 10 9 13 3 13 1 10 9 1 10 9 1 9 0 2
22 13 1 10 9 16 13 1 13 10 9 2 11 11 7 11 11 13 13 0 10 9 2
23 10 9 13 1 15 3 0 7 10 9 0 2 9 16 15 13 3 0 1 10 0 9 2
10 3 15 13 1 10 11 11 1 11 2
14 13 10 2 9 0 1 9 2 2 1 9 1 9 2
16 10 9 4 13 0 2 4 4 13 9 1 9 2 3 13 2
26 11 11 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 10 9 2 9 7 9 0 2
40 13 2 1 1 10 0 9 2 1 10 9 1 10 10 9 1 9 1 16 11 4 13 9 0 7 3 0 1 9 2 9 7 9 0 1 10 0 9 13 2
12 3 13 10 9 0 1 15 16 13 10 9 2
44 10 9 1 10 9 4 1 13 0 2 16 10 9 13 10 9 1 10 9 1 11 2 12 9 2 7 10 9 11 2 10 9 0 3 13 10 12 9 0 13 1 10 9 2
18 13 7 13 10 9 2 10 9 0 1 10 9 7 10 9 15 13 2
22 13 3 0 7 13 1 10 9 16 15 4 4 13 1 10 9 10 9 7 10 9 2
34 10 0 11 11 2 11 13 10 9 1 0 9 2 3 12 9 3 9 7 10 11 11 7 12 9 3 0 7 10 11 11 2 11 2
48 1 10 9 2 10 9 15 13 1 10 9 2 7 10 11 13 1 9 1 12 2 1 10 9 13 1 11 11 7 11 11 1 9 1 10 11 2 7 11 11 1 9 1 10 11 11 2 2
14 3 2 15 13 10 9 0 2 0 2 11 12 2 2
32 10 9 2 13 1 11 11 2 9 1 11 11 2 13 1 9 0 13 10 9 13 1 10 9 1 11 11 7 13 9 0 2
55 11 10 2 11 2 13 3 1 9 7 9 2 13 1 16 13 1 10 9 0 1 10 11 11 11 7 12 9 1 10 0 9 1 10 9 1 10 9 12 11 1 11 2 13 10 9 12 1 10 11 11 1 11 11 2
46 10 0 9 2 9 0 7 9 0 2 13 1 10 9 2 1 9 0 2 13 15 1 10 9 1 9 0 1 10 15 13 2 1 9 1 9 2 9 3 0 2 9 7 9 2 2
20 15 2 1 10 9 1 10 9 2 13 1 10 9 0 2 9 1 10 8 2
28 1 10 9 1 10 0 9 2 10 11 11 13 10 9 10 12 1 11 1 12 2 1 10 9 11 2 12 2
62 10 9 0 13 1 11 7 11 1 10 9 1 10 9 2 16 10 9 13 1 10 9 1 10 9 2 7 15 13 16 11 2 9 1 11 2 3 1 9 1 11 2 2 13 0 9 7 4 1 13 1 10 9 1 10 11 3 1 3 12 9 2
11 13 1 12 11 11 2 1 10 11 11 2
45 1 9 2 10 9 0 1 10 0 9 4 13 1 10 9 1 11 1 10 9 1 15 16 15 13 10 9 0 7 9 1 9 2 3 7 10 9 0 1 10 9 1 10 9 2
31 10 9 4 13 10 0 9 1 9 16 4 13 0 1 13 1 9 0 1 10 9 2 9 2 7 9 0 1 13 9 2
55 10 0 9 3 13 1 10 9 1 16 13 10 9 2 0 2 1 10 9 1 9 2 1 2 11 2 7 2 10 9 2 2 7 3 1 10 9 1 9 15 13 11 1 10 9 0 1 10 9 2 7 15 3 13 2
7 10 9 4 13 15 3 2
14 13 10 9 0 1 9 0 1 10 9 0 7 0 2
16 16 15 4 1 13 10 9 7 15 9 1 11 0 16 13 2
13 10 9 1 9 13 1 12 8 2 2 9 8 2
18 15 13 1 10 9 1 9 11 12 2 10 15 13 1 10 9 0 2
19 10 0 9 13 10 9 2 1 10 11 11 11 1 10 9 1 11 11 2
25 3 13 1 10 9 16 13 1 10 9 2 7 10 9 16 13 13 10 0 9 7 10 0 9 2
17 10 9 1 9 13 1 9 0 0 1 9 2 1 10 9 0 2
10 10 9 13 1 10 9 1 10 9 2
31 15 13 1 10 9 0 1 10 12 5 2 11 11 1 10 12 5 2 15 3 0 3 10 9 1 9 1 9 1 11 2
43 1 13 10 9 1 3 13 2 10 0 12 9 13 10 0 9 0 1 10 9 2 10 0 12 9 13 10 0 9 0 1 10 9 7 3 3 1 13 10 12 9 0 2
20 10 0 9 13 10 9 2 1 10 9 7 9 3 4 13 10 9 0 0 2
53 2 10 11 7 10 11 4 13 1 10 9 1 2 9 2 16 13 10 9 1 10 9 0 1 10 9 0 11 11 2 8 9 1 10 11 11 7 1 10 11 2 13 3 10 9 0 0 2 11 8 11 2 2
22 10 9 13 10 9 1 10 9 1 10 9 1 11 11 2 15 4 4 13 1 11 2
54 1 10 9 1 9 2 10 9 1 0 9 13 1 10 9 0 7 10 9 1 9 1 0 9 1 10 9 2 9 7 9 1 10 9 2 15 4 13 10 9 1 10 9 0 1 9 7 9 0 1 15 10 9 2
17 3 1 10 12 5 1 10 9 1 10 9 1 11 4 13 3 2
23 10 9 1 10 9 0 4 13 3 1 10 9 11 7 15 13 11 11 11 11 11 11 2
21 1 10 9 0 2 10 0 9 1 9 4 13 10 9 1 9 1 11 1 11 2
11 10 9 13 3 0 2 7 10 9 0 2
26 1 3 1 12 9 2 10 9 7 15 9 13 1 13 15 1 9 7 9 1 9 1 10 9 11 2
19 11 13 10 9 1 10 9 1 10 9 2 7 3 10 9 1 10 9 2
28 10 9 13 10 10 9 1 10 0 9 7 3 15 13 1 15 7 1 15 2 1 10 9 1 9 7 9 2
41 12 1 11 1 12 2 13 10 0 7 12 5 9 1 10 11 1 11 1 10 12 1 11 1 12 1 10 9 1 11 11 7 11 2 9 1 10 16 13 9 2
25 15 13 13 15 2 7 3 13 10 9 1 13 2 13 9 3 3 2 0 1 9 7 9 0 2
25 1 9 13 10 9 1 10 11 2 11 1 15 11 7 10 9 1 9 13 3 1 10 9 0 2
35 10 9 4 13 1 11 12 7 11 2 7 13 10 9 11 11 12 7 12 1 10 0 9 0 7 10 9 11 1 10 0 9 0 12 2
81 1 9 1 12 1 11 1 12 13 10 9 11 1 10 9 1 10 9 1 11 11 1 10 11 1 11 2 11 2 1 9 1 10 0 9 11 7 11 1 11 2 9 1 11 1 11 7 11 1 11 2 12 9 1 11 2 1 10 9 1 10 9 1 10 11 2 16 1 9 10 9 11 15 13 9 1 10 9 1 11 2
68 1 10 0 9 2 10 9 15 13 1 11 15 15 13 10 9 1 11 11 2 10 15 13 7 15 13 2 7 1 10 0 9 15 13 1 11 16 4 1 13 1 10 9 1 9 1 11 11 1 11 1 10 9 7 11 11 7 16 3 13 2 3 13 9 1 10 9 2
35 11 11 11 2 0 7 0 9 2 15 13 1 10 11 1 11 1 13 1 10 11 11 11 11 1 9 1 9 1 10 9 1 10 0 2
9 11 11 15 13 13 1 10 9 2
18 10 9 13 1 10 12 9 1 13 1 15 1 11 1 10 9 0 2
10 3 2 10 10 9 4 3 13 3 2
21 10 9 13 10 0 9 1 13 1 13 15 1 16 0 2 9 1 10 11 2 2
26 15 13 10 9 1 12 12 12 9 1 10 9 2 7 10 9 1 10 11 11 15 13 1 10 9 2
13 1 13 2 3 2 15 13 10 9 0 2 0 2
13 13 10 9 0 1 9 7 15 13 1 13 0 2
47 1 3 10 0 9 1 10 9 13 1 10 9 0 1 10 9 2 4 13 1 13 1 10 9 1 9 2 16 1 9 15 13 13 9 7 13 9 7 10 9 16 13 9 1 10 9 2
20 10 9 4 13 1 9 0 7 0 1 10 9 2 1 0 9 1 10 9 2
26 11 13 3 1 11 11 11 7 11 11 11 1 9 1 9 1 4 13 1 10 9 1 10 12 9 2
31 16 10 9 1 9 0 7 0 13 0 9 1 10 9 0 1 10 9 2 15 13 1 10 9 1 9 1 3 1 9 2
22 7 1 11 1 10 0 9 2 10 9 11 1 11 13 1 0 10 9 1 13 11 2
22 10 9 12 9 13 10 9 0 1 9 1 9 7 9 0 1 9 0 1 9 0 2
43 1 10 9 0 2 13 1 10 9 1 10 3 9 11 11 2 10 9 13 1 9 10 9 0 11 12 7 10 9 1 10 9 1 10 9 0 1 11 13 1 9 0 2
12 7 10 9 13 3 3 2 0 7 3 0 2
21 15 13 3 0 7 3 3 4 13 1 9 1 15 2 3 13 7 13 10 9 2
34 10 12 1 1 11 1 12 2 10 9 11 11 11 13 10 9 1 11 1 9 7 3 10 9 15 13 1 10 9 1 10 9 0 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
23 11 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 10 9 7 9 0 2
15 15 13 9 0 1 10 9 1 9 3 1 10 11 11 2
11 11 11 13 10 0 9 0 1 10 8 2
34 1 10 9 11 4 1 13 1 10 9 0 13 1 10 9 15 10 9 13 1 10 9 0 7 10 9 1 13 10 9 1 9 0 2
15 3 13 15 0 10 9 1 10 9 9 1 13 1 15 2
16 10 11 11 13 10 9 1 9 1 11 1 10 9 1 11 2
35 3 2 15 13 1 9 0 1 10 9 0 1 9 7 13 10 11 1 10 11 2 10 9 1 12 9 16 13 10 9 1 9 1 9 2
40 10 11 1 11 7 10 9 1 11 13 10 9 1 9 7 9 1 9 1 9 7 1 10 9 2 16 13 10 0 9 1 9 13 1 10 9 7 10 9 2
29 15 13 10 9 1 10 0 9 1 9 7 9 1 9 2 10 15 13 10 9 7 9 1 9 13 1 10 9 2
28 10 11 2 12 13 1 10 9 1 10 11 11 12 1 11 11 1 10 15 4 13 7 4 13 11 11 11 2
28 11 11 11 2 11 4 13 1 11 1 12 2 7 13 0 9 7 3 3 1 10 9 1 11 7 11 11 2
7 1 9 0 13 1 11 2
25 10 9 1 11 11 11 11 13 16 10 9 13 0 2 13 1 9 1 3 1 12 9 1 9 2
40 1 9 1 10 0 9 1 10 9 1 11 2 4 13 8 2 9 1 10 11 1 10 11 1 10 11 11 2 3 1 10 9 1 10 9 2 11 11 2 2
31 2 15 4 13 16 1 10 9 15 13 10 9 2 10 9 2 10 9 7 15 15 9 1 9 1 7 15 13 7 13 2
36 10 9 0 15 13 1 9 1 10 9 12 1 9 1 10 9 11 11 2 4 1 13 1 10 10 9 10 11 11 2 13 10 9 1 12 2
16 15 15 13 3 1 10 9 1 9 1 10 3 3 0 9 2
18 9 1 9 0 1 10 9 1 10 11 1 10 9 11 2 9 11 2
38 1 9 2 1 9 7 10 9 1 9 16 15 13 2 15 13 1 11 11 1 10 13 15 10 9 1 10 16 15 13 16 15 4 13 1 11 11 2
18 10 11 11 13 10 0 9 1 10 9 0 2 12 9 13 1 15 2
23 10 9 13 1 9 1 10 9 13 7 1 10 9 1 10 9 1 10 16 15 13 13 2
12 11 11 13 10 9 1 9 1 10 9 11 2
16 10 9 15 13 9 1 9 1 9 1 10 11 7 11 11 2
59 15 3 9 13 0 2 7 1 10 9 1 10 9 0 2 3 9 13 0 2 13 1 16 10 9 1 10 9 1 9 13 12 9 0 1 9 2 10 15 1 10 9 4 13 10 9 1 9 1 9 1 9 1 10 12 9 1 9 2
21 1 15 16 13 10 9 0 2 0 7 0 16 15 13 1 9 1 10 9 0 2
37 11 13 10 9 7 9 0 13 1 10 9 1 11 11 2 9 1 11 2 1 10 9 1 11 2 15 2 11 7 9 1 11 2 15 2 11 2
27 1 13 15 2 4 13 9 1 11 1 10 9 1 10 9 1 11 3 1 10 9 11 11 7 11 11 2
13 10 9 13 3 10 0 9 1 9 7 9 0 2
37 1 15 2 11 13 9 1 11 1 13 1 11 1 11 1 11 11 7 2 11 2 11 11 1 10 11 11 1 10 9 1 9 2 7 4 13 2
20 10 9 13 1 15 10 16 15 13 3 1 10 9 2 7 3 1 10 15 2
13 4 1 13 15 9 2 7 15 13 16 15 13 2
29 7 16 3 13 0 1 10 9 2 15 1 15 13 1 10 9 0 1 13 9 1 10 9 7 10 0 9 0 2
20 2 1 9 1 10 9 0 2 11 4 13 9 0 1 10 9 1 10 11 2
25 10 9 13 9 1 11 2 11 7 11 2 7 4 13 1 10 9 1 9 1 9 0 7 0 2
9 10 9 13 10 9 1 9 0 2
11 15 13 15 9 16 13 10 9 1 11 2
29 11 13 10 9 1 10 9 1 9 0 13 1 12 9 2 11 2 11 2 11 7 11 2 16 13 9 1 11 2
19 11 11 2 15 13 1 10 0 11 2 13 2 2 3 4 13 10 9 2
42 10 9 1 16 15 4 13 1 11 11 13 0 7 0 2 16 11 11 13 10 9 1 10 9 16 13 9 2 7 3 9 7 16 13 1 13 15 1 10 12 9 2
23 11 11 11 1 11 2 10 9 13 13 10 9 7 13 10 11 8 1 10 9 11 11 2
23 1 10 9 2 3 13 2 13 7 13 2 7 3 15 13 1 9 3 12 9 1 9 2
16 1 9 10 9 1 9 0 2 16 15 13 1 10 9 0 2
28 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 11 2
56 10 9 1 10 11 11 3 15 13 1 9 1 10 4 13 1 15 0 13 15 10 9 2 16 10 9 4 13 1 10 9 1 10 9 7 3 13 15 1 15 1 10 9 1 10 0 9 0 16 15 13 1 10 9 0 2
30 10 9 3 0 1 10 11 2 12 2 1 12 9 1 9 1 10 9 0 2 4 13 1 10 9 1 11 2 12 2
21 13 0 1 10 9 1 11 2 7 4 4 13 1 10 9 1 11 7 11 11 2
33 7 3 2 11 11 13 1 10 9 10 9 1 11 11 11 2 10 9 16 13 1 11 11 2 3 13 9 0 1 11 1 9 2
21 10 9 0 13 1 11 11 15 4 7 13 9 3 1 10 0 9 1 10 9 2
69 12 9 3 2 7 1 10 13 10 9 1 3 2 10 9 13 10 9 1 10 15 15 13 10 2 9 1 9 1 10 9 1 9 1 10 10 9 2 16 15 13 10 9 1 9 2 1 10 9 1 16 13 10 9 2 13 1 10 0 9 1 10 9 0 2 1 10 9 2
17 10 9 1 10 9 0 3 13 10 9 1 16 10 9 4 13 2
7 4 13 1 10 12 9 2
60 1 12 2 15 13 1 10 9 12 1 10 9 1 10 12 0 9 1 9 1 10 9 2 12 11 11 11 2 13 1 2 11 11 11 2 7 4 13 1 9 1 10 11 1 10 11 1 10 11 11 2 11 11 11 11 2 11 11 2 2
18 13 10 9 16 13 10 12 9 1 9 2 1 9 16 13 10 12 2
20 15 13 1 11 2 7 1 9 7 9 13 10 10 9 1 10 9 1 11 2
29 13 1 15 16 10 9 13 10 0 9 1 10 9 2 3 16 13 13 15 1 10 9 7 13 10 9 7 9 2
32 10 9 1 10 9 0 13 1 10 9 1 10 9 1 2 2 11 11 2 11 11 2 2 9 16 13 0 1 10 9 0 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
22 1 0 9 1 10 9 2 10 9 9 1 11 11 4 13 10 12 1 11 1 12 2
16 10 9 15 13 13 1 11 11 7 11 11 1 11 2 11 2
29 11 13 16 11 15 13 16 13 16 3 13 1 9 2 7 13 13 1 11 1 16 3 15 13 2 7 1 9 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
9 13 1 9 0 7 9 3 0 2
40 10 9 2 9 2 9 2 9 2 9 2 9 7 9 13 1 10 11 7 1 15 9 1 10 9 0 1 10 9 11 7 3 13 0 1 10 9 1 11 2
26 10 9 2 11 2 4 13 1 10 9 11 7 10 9 0 2 15 1 10 9 8 7 8 2 3 2
34 11 11 13 10 12 1 11 2 3 1 13 10 9 1 3 1 12 9 12 12 9 2 9 1 10 9 11 11 2 3 13 1 9 2
19 1 10 9 2 10 9 0 16 13 10 9 1 10 9 13 10 9 3 2
13 10 9 1 9 13 1 12 8 2 5 5 5 2
27 13 1 11 1 10 9 1 12 9 2 1 10 12 9 4 13 10 9 16 13 1 9 0 7 13 15 2
37 1 9 1 9 2 10 9 3 0 13 10 9 2 7 16 13 10 9 2 10 9 16 13 10 0 9 1 9 1 13 10 9 0 13 10 9 2
30 10 12 1 11 1 12 2 10 9 11 2 11 4 13 9 1 9 1 10 12 9 1 9 2 7 13 1 11 3 2
35 10 9 1 11 11 2 13 1 10 9 1 12 1 10 9 11 11 11 2 13 1 9 10 12 1 11 1 12 2 1 10 9 1 11 2
42 3 3 10 9 13 10 9 1 11 2 3 15 13 10 11 1 11 15 13 3 1 12 9 1 9 1 10 9 0 16 13 3 1 12 9 10 9 1 15 1 11 2
46 11 2 1 9 3 11 2 13 10 9 0 2 13 1 10 9 1 10 9 2 7 10 9 1 10 9 2 9 1 10 9 7 9 0 1 11 2 1 10 9 0 1 10 11 11 2
12 11 2 13 10 9 0 9 1 10 9 11 2
21 15 16 3 15 13 2 9 9 2 7 15 16 3 4 13 15 2 9 9 2 2
40 10 9 11 7 9 11 2 1 9 11 11 11 11 2 16 13 10 2 9 1 10 9 2 2 13 10 9 1 10 9 1 11 2 13 1 10 9 1 11 2
32 10 0 9 13 16 10 9 1 10 11 1 11 11 11 15 13 1 9 1 10 9 1 9 12 1 11 7 10 11 11 12 2
12 13 9 0 16 13 9 0 2 0 2 0 2
25 11 11 11 11 2 11 2 12 2 11 2 12 1 11 1 12 2 13 10 9 7 9 0 0 2
28 10 9 1 10 9 3 4 4 13 1 10 9 1 10 9 2 16 13 15 16 4 13 10 9 1 10 9 2
20 13 16 10 9 4 13 3 1 1 10 9 0 2 1 9 1 13 15 0 2
59 10 9 1 10 9 4 13 1 9 1 16 1 15 15 4 13 10 9 0 7 1 10 9 2 4 13 15 10 9 1 10 9 0 8 2 8 7 3 8 2 3 16 3 3 13 10 9 3 13 7 10 0 9 1 13 7 1 13 2
28 10 11 11 13 1 10 9 1 10 11 11 1 11 7 11 2 10 11 11 2 9 7 9 1 10 11 11 2
21 10 9 13 1 9 10 9 1 11 11 2 1 11 2 3 13 10 9 1 9 2
20 3 10 9 16 15 13 15 13 1 13 15 16 13 7 13 15 10 0 9 2
17 10 9 4 13 1 10 9 1 9 13 1 9 1 10 0 9 2
41 7 1 12 1 13 15 13 1 10 11 1 11 2 10 9 4 4 13 2 3 1 10 10 0 9 1 10 9 1 10 9 11 2 1 9 1 10 11 1 11 2
32 10 9 1 10 9 16 13 10 9 1 10 9 2 10 9 16 10 9 1 9 2 13 10 2 10 9 7 15 13 9 0 2
68 12 1 15 13 11 11 11 2 9 0 1 9 2 7 11 11 2 9 1 9 2 15 0 9 1 10 9 15 13 11 2 7 15 4 13 1 10 9 16 13 1 10 9 1 10 9 1 10 11 10 9 11 11 2 3 4 13 10 9 1 10 2 9 2 11 11 2 2
43 10 11 11 2 0 1 10 9 1 11 11 1 10 11 2 13 10 9 0 0 13 1 10 11 11 1 13 1 10 9 7 5 7 9 1 10 11 1 10 11 1 11 2
43 10 9 1 9 1 10 11 1 11 4 13 10 9 1 12 9 16 13 10 9 16 13 1 10 9 0 1 11 7 13 15 1 10 9 8 2 1 9 1 10 9 0 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
26 1 10 9 1 10 9 0 2 11 13 1 11 1 11 11 1 13 10 9 12 2 12 1 10 11 8
30 10 9 13 10 9 1 11 1 11 2 1 10 12 9 0 2 1 10 0 9 1 9 2 7 13 10 9 1 9 2
22 1 12 2 15 13 10 9 1 9 1 9 16 3 10 9 13 1 10 9 1 11 2
43 2 11 11 2 13 10 9 15 13 11 11 1 12 1 13 9 1 10 9 2 10 9 7 10 9 1 10 9 0 2 1 10 9 13 10 9 3 0 2 0 7 0 2
7 13 9 14 2 12 1 2
28 10 9 2 13 1 10 11 1 10 9 1 9 1 10 11 2 7 13 3 3 1 10 11 8 1 9 0 2
33 10 9 4 13 1 12 7 12 1 10 0 9 11 11 2 11 11 2 11 11 7 11 11 2 15 13 1 13 10 11 1 12 2
43 1 3 13 10 9 1 9 16 3 13 10 9 1 11 2 16 13 16 13 15 2 2 7 15 13 13 10 9 2 13 10 9 1 9 1 3 2 7 3 13 16 13 2
38 3 15 13 10 9 1 10 9 1 10 9 2 1 10 9 16 13 1 9 10 9 9 1 10 9 1 11 1 10 9 1 11 1 13 4 13 9 2
48 1 9 1 10 9 1 10 9 3 1 10 0 9 2 9 2 13 10 9 1 10 9 2 1 10 10 9 1 1 13 10 9 0 1 10 9 2 16 4 13 10 9 3 1 10 9 11 2
22 13 10 0 9 1 10 9 0 2 13 1 10 9 1 10 9 0 11 11 1 11 2
18 15 13 16 10 9 0 15 13 1 15 15 4 13 1 10 11 11 2
11 3 1 10 9 10 9 13 3 1 9 2
25 10 9 13 1 10 9 1 11 7 9 1 11 1 11 1 10 9 11 7 10 9 11 1 11 2
47 0 13 10 0 9 1 10 9 1 9 0 1 13 1 11 2 1 10 9 0 7 0 1 10 9 0 7 1 10 9 1 10 9 13 1 11 11 11 16 13 2 11 1 10 9 2 2
18 1 10 9 2 10 9 13 10 9 0 7 15 4 13 10 9 0 2
17 11 11 13 1 10 9 1 10 9 0 1 11 2 9 1 9 2
25 10 9 1 10 11 7 10 9 0 4 13 1 0 7 0 9 1 9 1 10 9 0 7 0 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
29 1 10 9 15 13 1 9 1 9 1 9 0 0 1 10 9 12 7 12 7 15 13 1 10 9 1 9 0 2
39 1 10 9 1 10 0 9 2 10 9 0 15 13 9 1 10 9 1 10 9 9 11 1 11 11 2 15 1 10 9 13 1 10 9 13 10 9 0 2
16 10 9 13 2 13 10 9 1 10 9 1 9 1 10 9 2
3 13 12 2
27 11 13 10 9 0 1 11 2 7 10 9 13 13 9 1 13 10 9 1 10 9 0 1 12 9 0 2
45 10 9 4 13 3 0 2 3 15 15 4 13 16 10 9 13 1 11 7 11 13 1 9 1 10 9 0 2 15 1 10 9 3 13 1 9 7 9 7 1 3 9 1 9 2
29 2 16 1 11 15 15 13 12 12 7 12 12 9 2 1 15 15 13 1 10 9 0 1 9 2 2 15 13 2
14 10 9 0 13 15 13 1 10 9 1 10 9 0 2
20 1 12 1 12 13 1 10 9 0 1 11 7 13 1 10 9 1 10 9 2
23 1 10 9 0 1 9 1 11 2 10 9 1 12 13 1 12 2 12 9 7 12 9 2
40 1 10 8 0 1 10 11 2 4 13 15 8 16 10 9 4 13 1 10 9 16 15 13 9 1 10 9 0 2 1 10 9 0 7 1 10 9 1 9 2
26 3 2 10 9 1 9 0 2 11 4 13 15 1 10 0 9 0 0 7 0 1 10 9 1 12 2
8 10 9 13 9 1 13 15 2
30 13 1 10 0 9 10 12 2 10 12 1 11 13 10 0 9 1 10 9 2 10 9 15 13 1 10 9 1 11 8
18 11 13 9 7 10 9 13 10 9 12 1 10 11 7 11 11 11 2
38 1 10 9 13 10 9 16 13 9 1 9 10 9 1 10 9 2 16 13 13 15 7 13 1 10 9 1 4 13 1 13 10 0 9 0 1 11 2
12 4 13 1 12 2 1 10 9 11 11 11 2
18 7 15 16 15 13 1 15 13 16 15 13 10 9 2 13 15 13 2
41 11 11 11 2 13 1 12 2 13 10 9 0 13 1 10 9 1 9 11 2 11 2 12 2 7 10 9 11 1 9 2 12 2 2 0 1 10 11 11 11 2
23 10 9 1 11 7 9 0 13 0 7 1 9 3 0 9 2 15 3 0 1 0 9 2
15 10 9 13 10 9 1 10 9 1 10 9 1 10 9 2
10 15 13 12 9 7 11 12 7 12 2
21 13 12 9 0 2 9 0 7 1 9 0 2 9 1 9 2 9 2 8 2 2
42 10 11 11 11 2 13 10 9 1 12 1 10 9 0 2 1 12 10 9 1 10 9 13 13 15 7 13 10 9 1 10 9 1 10 9 11 2 11 7 11 11 2
30 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 5 12 7 10 9 0 1 9 13 5 12 2
30 10 9 3 3 2 11 11 11 13 15 9 2 13 16 10 9 2 1 9 1 10 9 0 1 9 2 13 3 0 2
16 1 10 9 2 1 10 7 15 13 13 13 15 1 10 9 2
25 10 9 13 10 9 1 0 9 1 10 9 1 10 11 7 10 9 1 10 9 0 1 10 9 2
4 13 1 11 2
35 11 11 4 13 10 9 1 9 1 10 9 1 0 9 0 2 7 10 9 1 10 11 11 2 11 11 11 2 4 13 9 1 10 9 2
11 3 13 0 9 0 1 10 9 1 9 2
10 10 9 13 1 12 9 7 12 9 2
25 1 11 3 13 10 9 1 10 9 2 13 9 1 10 0 11 13 15 1 13 1 10 11 10 2
15 13 1 9 1 9 13 9 0 1 11 1 12 7 12 2
37 3 3 2 11 13 1 12 9 0 2 12 9 2 12 9 2 15 0 7 15 9 2 2 7 10 9 0 2 9 2 1 10 11 11 1 11 2
30 1 10 9 13 0 13 1 9 2 8 5 12 1 9 2 8 5 12 2 16 1 9 0 3 13 0 13 9 0 2
21 4 13 1 11 10 9 2 1 11 11 2 3 1 11 7 3 1 11 1 11 2
13 10 9 13 10 9 1 12 12 9 1 10 9 2
34 10 9 1 9 1 9 0 7 10 9 7 9 16 13 1 9 0 1 10 9 1 10 15 13 9 2 3 13 13 1 10 9 0 2
20 10 9 13 15 16 13 2 13 12 9 7 12 13 3 4 13 1 10 9 2
16 10 11 11 2 10 0 9 2 13 10 9 1 9 11 1 8
8 8 9 1 10 9 0 11 2
43 10 9 13 10 0 9 7 13 10 10 9 2 10 9 13 10 16 13 1 3 13 13 2 10 9 13 13 2 7 10 9 13 16 13 2 13 15 10 9 1 10 9 2
15 15 13 9 1 10 9 2 10 9 1 10 9 13 0 2
57 1 10 9 1 10 9 3 3 4 4 13 1 10 0 11 11 12 1 10 8 8 16 13 9 1 15 3 15 15 13 2 3 7 2 1 15 3 13 3 10 9 1 10 9 16 3 4 13 13 15 1 10 9 1 10 11 2
51 13 10 9 16 13 16 11 13 1 10 9 0 1 10 15 13 10 9 16 10 9 1 10 9 11 2 10 11 11 2 15 13 1 10 9 1 9 1 9 13 1 10 9 2 4 3 13 1 10 9 2
27 13 1 10 9 2 7 10 12 1 11 15 13 3 1 10 9 0 2 16 15 13 1 10 9 1 11 2
15 10 9 4 4 13 3 1 11 2 3 1 10 9 0 2
21 1 0 13 1 10 9 1 10 9 1 11 2 11 15 13 1 10 9 1 9 2
12 10 9 8 8 1 10 9 13 1 5 12 2
40 0 9 1 10 9 13 1 10 9 7 10 9 1 10 8 8 16 4 13 1 10 9 2 13 1 10 12 9 1 10 9 7 3 15 13 1 11 2 11 2
36 10 9 16 13 13 3 1 10 12 5 1 10 9 2 10 9 1 10 9 1 10 11 13 0 2 2 13 10 9 0 9 1 9 7 15 2
14 15 13 1 9 10 9 1 3 1 12 9 1 9 2
22 1 10 9 12 13 10 9 1 12 9 1 10 9 1 9 1 12 9 1 9 5 2
22 11 11 11 11 2 12 1 11 1 12 2 2 9 7 9 0 0 1 10 11 11 2
19 1 10 9 2 13 1 11 2 10 9 1 11 11 2 9 1 10 9 2
33 10 9 13 10 9 1 10 9 2 1 15 15 1 10 9 0 1 10 9 0 2 11 11 2 3 7 15 1 10 9 7 9 2
36 10 0 9 1 9 13 10 9 0 1 10 9 2 9 3 1 10 9 3 0 7 0 2 16 13 10 9 2 10 9 1 9 7 10 9 2
16 13 1 11 10 12 1 11 7 10 12 1 11 13 1 11 2
29 10 11 11 15 13 13 1 10 0 9 1 9 7 10 9 1 9 7 13 10 9 0 0 1 10 9 1 9 2
83 7 2 16 10 9 1 10 9 13 1 10 9 1 10 9 1 10 9 0 1 10 9 2 10 9 4 1 13 15 2 1 9 2 1 10 9 1 10 9 10 9 1 9 8 11 11 1 11 2 10 12 1 11 1 12 2 1 10 9 1 10 9 1 11 11 2 9 11 1 10 11 2 3 0 1 10 9 0 2 11 1 11 2
33 1 10 9 1 3 2 7 3 1 10 9 13 2 15 13 9 1 10 9 7 10 9 3 13 13 15 9 7 1 9 7 9 2
13 10 10 9 13 0 2 7 15 1 15 15 13 2
7 10 9 3 15 4 13 2
17 10 11 13 11 2 9 1 10 11 2 13 1 10 9 0 11 2
54 13 10 13 2 11 1 10 11 2 7 2 11 11 2 15 13 1 9 7 9 2 1 15 13 9 2 1 10 15 13 10 9 3 0 1 13 15 10 9 7 1 9 0 15 13 10 9 1 13 15 1 10 9 2
44 2 13 1 10 9 1 10 9 7 1 15 15 13 1 9 1 10 9 2 1 10 9 2 16 13 10 9 13 1 10 9 0 0 8 10 0 9 1 10 9 2 2 13 2
33 10 9 15 13 3 1 10 9 13 1 10 11 11 2 10 9 15 4 13 1 10 9 1 10 9 12 1 10 9 16 13 3 2
27 15 13 10 9 11 12 1 11 7 10 9 11 12 11 1 11 2 3 3 13 2 13 1 13 1 11 2
18 10 0 9 16 13 10 15 0 2 7 1 15 15 12 1 12 13 2
44 10 11 2 1 13 10 9 7 10 9 1 10 9 2 4 13 10 9 1 10 9 2 13 1 10 9 1 16 1 10 9 0 1 10 12 9 1 9 2 10 11 13 0 2
28 10 9 13 9 1 10 9 7 15 13 1 0 9 1 9 2 15 13 7 9 0 9 16 15 13 3 3 2
27 2 11 11 11 1 11 2 11 2 13 10 9 13 1 10 9 11 2 13 3 1 10 9 1 12 11 2
13 3 1 10 9 2 10 9 0 13 10 9 0 2
11 10 9 1 11 15 13 13 1 10 9 2
21 3 13 10 11 11 1 11 11 1 12 2 16 13 10 9 7 9 1 10 9 2
54 11 11 4 13 3 1 10 9 1 10 9 3 1 10 9 0 2 1 10 9 8 8 8 8 8 2 1 10 9 1 10 9 12 7 1 10 9 1 9 2 10 11 13 10 9 1 9 7 13 0 10 9 9 2
36 10 11 1 10 11 13 3 10 9 1 10 9 0 2 13 1 10 9 0 2 1 9 0 1 3 0 9 7 13 9 1 9 1 10 9 2
56 1 11 1 12 2 9 1 15 13 1 10 9 1 10 11 2 13 10 9 1 10 9 7 10 9 0 2 13 1 15 1 10 9 1 11 11 1 10 0 9 0 1 10 11 1 11 1 11 2 10 12 1 11 1 12 2
32 9 2 9 2 9 2 9 0 7 3 9 1 10 9 2 15 13 3 1 10 9 1 10 9 12 1 10 9 1 11 11 2
53 10 9 16 4 13 1 10 9 1 10 9 7 1 10 9 1 9 1 10 9 4 13 10 9 16 4 13 3 2 3 15 13 10 9 1 10 9 7 10 9 13 15 15 13 3 15 15 15 13 1 9 0 2
14 13 0 1 10 9 1 9 1 10 11 1 12 9 2
29 2 11 2 15 13 3 1 10 9 1 11 2 15 13 10 9 0 7 15 13 0 16 15 13 12 9 1 9 2
19 1 9 3 1 10 9 4 13 15 1 10 9 1 9 7 9 1 9 2
11 10 9 1 11 15 13 13 1 10 9 2
36 3 2 13 10 9 1 9 0 7 0 2 10 11 11 2 10 9 13 10 9 0 7 0 1 10 9 2 10 9 7 15 9 1 0 9 2
26 2 11 2 11 13 16 10 9 1 15 13 0 1 10 9 7 16 10 9 7 10 9 13 3 0 2
18 10 9 1 10 8 13 3 15 13 1 10 9 1 8 1 10 9 2
22 13 1 11 11 2 11 11 7 11 11 2 10 9 15 13 1 11 2 11 11 2 2
19 15 13 10 9 1 9 16 4 13 9 1 10 9 1 10 11 1 11 2
42 13 10 9 16 13 1 10 9 0 1 13 2 11 2 13 10 9 1 10 9 2 2 11 11 2 10 11 1 10 11 2 10 11 1 10 11 2 11 2 10 11 2
9 9 0 2 11 11 2 11 11 2
12 10 9 8 1 10 9 15 13 1 10 9 2
13 10 9 13 1 10 0 9 7 10 9 1 11 2
13 15 13 13 1 9 1 10 9 1 10 9 0 2
27 1 2 11 0 2 15 13 16 15 3 13 1 10 9 1 11 2 11 11 10 11 1 15 3 12 9 2
49 1 9 15 13 10 9 11 11 16 13 10 9 0 2 3 13 7 13 7 2 1 10 9 2 11 12 16 1 10 9 13 1 10 9 1 10 9 1 13 1 15 7 10 9 1 13 1 15 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
40 10 9 1 10 9 3 15 13 7 13 10 0 9 1 9 0 2 7 1 9 2 9 2 9 2 9 7 9 2 2 7 10 9 1 9 0 13 3 0 2
8 11 15 13 13 1 10 9 2
32 1 9 3 3 13 10 9 1 9 1 10 9 7 3 13 3 2 7 10 9 13 10 9 16 13 3 7 13 13 10 9 2
28 10 9 13 3 3 12 9 2 7 15 4 13 1 10 9 1 9 1 10 9 1 10 12 9 1 12 9 2
37 1 9 2 10 9 1 10 9 4 13 1 9 0 1 13 10 11 2 12 2 1 0 1 11 2 12 2 2 16 13 3 0 1 10 0 9 2
33 10 0 9 1 10 9 1 10 9 13 10 9 7 11 13 10 0 9 2 10 11 11 2 1 10 15 13 10 9 1 10 9 2
19 1 11 2 9 1 11 2 10 0 9 1 9 1 9 13 2 0 2 2
21 1 10 9 1 12 5 2 10 9 11 11 13 3 10 9 0 7 10 9 0 2
5 15 13 1 11 2
44 10 9 13 9 2 1 3 10 9 13 10 0 9 1 10 9 0 2 16 4 13 10 9 16 13 13 1 10 11 11 1 10 11 3 1 10 0 9 2 1 13 1 15 2
13 10 9 0 16 13 1 10 9 13 1 9 0 2
19 2 4 10 9 13 1 9 16 7 15 13 1 10 9 13 1 10 9 2
46 10 9 2 0 9 2 4 1 13 1 13 0 9 2 7 13 1 11 2 1 9 1 9 7 1 10 9 2 10 9 1 9 16 15 13 0 1 10 9 16 13 10 9 2 11 2
41 10 9 0 1 11 7 1 9 2 11 11 11 2 11 2 2 13 10 9 0 9 1 12 9 2 12 9 2 2 1 9 0 2 16 4 13 1 11 2 11 2
39 11 11 13 13 10 9 1 10 9 1 13 9 0 1 13 10 9 7 13 10 9 1 2 9 1 9 2 7 9 1 9 3 1 10 9 1 9 0 2
23 10 9 16 13 10 9 13 10 9 0 1 10 9 7 9 0 2 15 15 13 10 9 2
8 13 10 9 0 1 10 9 2
23 1 10 9 2 15 13 10 9 1 9 1 11 2 13 1 10 9 1 10 9 1 11 2
47 10 9 4 13 10 9 1 12 5 2 5 1 10 9 1 10 9 7 1 12 5 2 5 1 10 9 1 10 9 2 11 2 1 10 9 3 13 1 9 10 9 1 9 2 0 2 2
9 1 12 9 16 13 13 3 3 2
24 1 10 9 4 13 1 10 11 13 1 13 10 9 1 10 9 1 9 2 13 1 11 11 2
21 13 1 9 12 9 2 12 9 0 7 12 0 2 1 12 9 0 1 10 11 2
18 10 11 13 10 9 1 9 2 3 13 1 9 2 1 10 11 11 2
36 13 1 10 9 1 10 11 2 10 9 1 10 9 13 0 2 1 9 16 13 1 10 12 5 2 11 7 11 11 11 2 7 10 12 5 2
33 10 9 13 1 12 1 13 1 10 9 1 12 9 2 11 7 11 11 2 2 1 12 13 1 13 15 11 11 7 13 1 12 2
20 13 10 9 2 3 13 1 10 9 10 9 1 10 16 4 13 1 10 9 2
43 3 1 15 2 1 9 1 0 7 0 9 2 11 2 1 9 7 9 2 13 1 10 9 10 9 2 16 3 13 10 15 15 2 10 9 2 4 13 7 13 1 15 2
31 10 9 4 13 10 9 2 10 0 9 1 12 4 13 1 10 9 1 10 11 1 11 1 12 1 10 9 1 11 11 2
19 1 12 7 12 15 13 10 9 1 9 16 13 1 9 1 10 9 12 2
41 11 13 1 11 1 12 7 13 3 13 1 10 9 1 10 9 11 1 11 11 7 13 9 1 10 9 0 1 15 1 10 9 0 2 16 13 1 9 7 9 2
35 10 9 12 4 13 1 10 9 1 10 11 1 11 11 10 12 1 11 1 12 7 13 10 12 1 11 1 12 1 10 9 12 2 12 2
25 1 10 0 9 1 9 2 10 9 13 10 9 1 9 1 13 1 10 9 0 1 10 9 0 2
18 11 2 11 11 2 7 11 11 15 13 0 13 1 10 9 1 11 2
23 10 11 11 13 10 9 1 9 9 0 2 13 1 11 11 1 12 1 10 9 1 11 2
10 3 11 7 15 4 13 1 9 0 2
37 10 9 1 9 7 10 9 1 10 9 7 9 13 1 1 10 9 15 13 7 1 10 9 13 1 9 1 10 9 1 10 10 9 16 15 13 2
15 13 10 9 13 3 3 16 13 10 9 7 9 16 13 2
28 13 10 9 1 10 11 11 1 10 12 7 12 9 1 10 9 1 12 7 12 3 2 15 15 4 13 11 2
33 3 15 13 10 9 2 3 3 13 10 10 9 3 7 13 10 9 0 2 15 16 1 10 9 1 10 9 7 10 9 13 9 2
16 1 10 9 15 13 9 0 1 9 13 10 9 1 10 9 2
15 1 2 11 11 2 13 1 11 7 11 7 13 9 0 2
42 1 9 3 0 7 10 0 9 1 9 2 10 9 13 13 1 10 9 1 13 9 1 10 9 2 7 13 1 10 9 3 10 9 15 13 2 2 1 15 13 0 2
7 9 13 9 1 10 11 11
21 11 13 10 9 0 1 9 7 9 2 13 1 11 11 2 11 7 13 1 12 2
9 10 9 15 13 1 10 11 11 2
41 10 9 15 13 1 9 1 10 9 15 10 9 13 1 10 9 7 3 11 13 9 1 10 9 1 9 1 11 11 2 11 11 2 11 7 11 11 2 1 15 2
18 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 11 2
20 10 9 15 13 3 3 0 2 7 1 10 9 15 4 13 11 1 10 9 2
26 10 9 13 1 15 9 16 4 13 7 13 10 9 0 16 13 1 10 9 2 7 15 3 13 0 2
14 13 10 9 0 1 10 9 1 10 2 9 0 2 2
57 10 9 1 10 13 1 9 2 11 11 11 2 13 1 11 11 16 10 9 13 2 3 0 2 15 1 10 0 9 7 1 10 9 1 10 9 1 15 9 9 12 1 11 2 16 15 4 13 15 7 4 13 10 0 9 2 2
33 13 1 10 9 0 1 10 9 1 12 2 10 0 9 2 1 10 0 9 0 1 10 9 2 13 10 9 1 9 1 11 11 2
19 10 9 4 13 1 10 0 9 1 10 9 0 13 1 10 9 1 12 2
27 10 0 8 1 11 1 10 9 9 11 13 15 1 10 9 8 16 1 15 0 13 10 9 1 10 9 2
23 11 13 10 9 0 7 10 9 1 10 9 1 11 2 1 10 9 1 11 2 11 2 2
7 13 10 9 16 4 13 2
17 13 0 2 0 2 0 7 13 13 10 9 1 10 9 7 9 2
13 10 0 9 1 9 13 10 11 11 11 10 11 2
6 15 13 1 11 11 2
36 1 12 2 16 3 13 0 13 10 9 0 11 11 1 10 9 11 7 11 1 11 1 9 7 9 2 13 10 9 1 10 9 11 11 11 2
5 13 0 1 11 2
24 3 1 13 15 1 9 2 11 4 1 13 9 1 10 9 0 1 10 11 11 2 10 12 2
37 1 9 1 10 9 7 10 9 2 13 15 3 16 10 9 1 10 9 16 13 10 9 2 16 10 10 9 1 10 9 1 10 9 13 1 11 2
30 1 10 9 1 10 0 9 2 10 9 13 1 0 9 1 12 9 2 7 10 9 1 10 9 1 9 13 3 0 2
25 16 1 10 9 0 3 15 13 1 13 9 2 13 10 9 13 1 10 11 7 3 13 10 9 2
21 10 9 0 13 0 1 10 9 0 0 1 10 9 1 11 7 10 9 1 11 2
4 3 13 15 2
24 13 1 10 9 13 1 16 13 0 9 16 13 13 15 1 10 9 0 10 9 2 2 13 2
13 13 1 11 1 12 3 0 3 13 9 1 12 2
30 1 10 9 0 1 10 9 12 2 15 10 9 1 10 9 15 13 1 9 0 1 10 9 0 1 9 7 0 9 2
23 1 12 15 13 1 9 1 10 11 11 1 10 11 11 7 15 13 1 11 11 11 11 2
50 10 9 3 0 13 10 9 0 7 9 1 10 9 9 1 11 2 1 10 9 9 1 10 9 0 1 10 9 1 9 0 1 10 9 0 7 10 9 0 2 3 7 10 9 1 10 9 1 11 2
20 1 10 9 1 12 13 1 12 9 2 13 1 12 1 10 9 0 1 12 2
44 1 10 0 9 1 10 9 15 13 10 9 1 10 9 1 10 9 1 9 2 16 13 1 10 9 7 1 10 15 15 13 10 9 2 13 10 9 2 16 13 3 4 13 2
13 11 11 13 10 9 0 1 9 1 11 2 11 2
35 1 11 2 10 9 1 11 13 1 13 10 9 1 11 1 2 10 3 3 2 2 7 10 9 4 13 15 1 10 0 9 1 10 9 2
31 1 10 9 1 12 2 1 9 1 10 11 2 10 9 13 10 9 1 9 0 1 12 9 1 10 12 12 9 13 0 2
56 1 10 9 2 1 10 0 9 7 9 1 10 0 9 1 10 11 2 11 11 2 10 9 2 15 13 1 10 9 10 0 9 1 9 1 10 9 1 12 9 2 13 1 10 9 1 9 2 9 2 9 2 9 7 9 2
19 10 9 13 10 15 1 9 2 16 13 10 9 1 9 1 12 1 12 2
37 10 9 4 13 10 12 1 11 2 10 9 3 1 10 9 1 10 9 0 13 3 1 10 9 1 11 11 2 1 10 9 1 13 3 12 9 2
18 10 0 9 2 10 9 11 11 13 1 10 9 1 11 1 9 0 2
14 1 9 2 11 11 13 0 9 1 13 1 10 11 2
9 10 9 16 13 15 4 13 15 2
24 13 10 9 3 0 16 15 13 1 9 1 9 7 15 13 10 9 1 8 2 8 1 9 2
24 10 9 0 13 15 15 10 10 12 9 3 4 13 2 13 1 10 9 0 1 10 0 9 2
33 11 11 11 2 11 2 1 10 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 2 13 10 9 0 1 10 9 2
13 13 10 0 9 1 3 1 9 1 10 11 11 2
47 1 10 11 11 11 2 10 9 1 9 0 16 13 9 13 10 9 1 13 9 1 10 0 9 1 10 9 1 9 0 1 10 9 0 1 4 7 13 15 1 10 9 1 9 7 9 2
12 11 11 13 10 9 1 9 1 10 9 11 2
18 10 9 1 9 0 1 9 0 3 7 10 9 1 10 9 13 11 2
14 13 10 9 1 10 9 11 3 13 0 9 1 9 2
11 1 12 2 0 1 11 2 13 10 9 2
42 11 2 1 12 9 2 13 1 9 1 9 1 9 1 9 1 10 9 1 10 9 1 10 11 1 10 11 2 10 9 13 1 9 3 13 12 9 13 10 9 0 2
39 1 15 2 1 10 9 2 13 1 10 9 13 1 10 9 16 13 10 9 1 10 9 2 1 9 1 16 15 9 4 13 1 9 7 9 1 10 9 2
22 1 12 4 13 1 10 9 2 11 11 1 10 11 2 2 11 11 1 10 11 2 2
12 3 10 9 4 13 12 9 1 9 1 9 2
11 2 7 3 15 13 3 2 9 1 9 2
21 10 9 4 13 1 9 3 0 1 10 11 11 1 10 11 11 1 11 1 12 2
14 10 9 13 10 0 9 16 11 11 2 2 1 12 2
26 1 12 15 15 13 10 9 1 10 9 1 10 11 1 10 11 7 1 10 11 2 13 15 1 11 2
13 13 3 1 10 9 2 7 1 15 15 13 3 2
16 10 9 0 13 10 9 0 1 10 9 11 1 11 7 11 2
19 10 9 1 10 9 13 12 9 7 10 9 1 10 9 10 12 9 3 2
81 10 12 1 11 1 12 10 9 0 2 10 2 11 11 11 11 2 2 13 10 11 11 1 11 13 10 0 9 0 1 10 9 2 1 12 10 11 1 11 7 11 2 10 12 1 11 1 12 10 11 11 2 11 2 2 10 12 1 11 1 12 10 11 1 11 11 1 11 2 10 12 1 11 1 12 10 11 11 11 11 2
18 13 3 1 12 9 0 2 1 11 3 10 9 11 11 7 11 11 2
15 1 10 9 15 4 13 10 9 1 10 9 0 13 11 2
13 11 7 15 13 10 9 1 13 15 4 4 13 2
21 13 10 9 13 1 10 9 0 7 10 9 0 2 13 3 10 9 7 10 9 2
37 11 11 11 11 2 5 2 13 10 9 1 9 1 9 1 9 1 9 2 1 9 1 11 2 16 15 13 1 13 9 1 9 1 10 0 9 2
21 15 13 13 9 16 4 13 9 1 10 9 2 7 16 15 3 4 13 10 9 2
32 10 9 0 1 11 2 9 1 10 9 12 2 13 10 9 1 9 7 10 9 0 7 13 10 9 16 10 9 13 10 9 2
31 13 10 9 1 9 0 2 1 0 9 2 1 10 15 15 13 10 9 1 9 2 9 7 9 1 10 11 2 12 11 2
36 13 0 10 2 9 2 1 15 16 13 10 9 1 9 16 13 10 9 1 10 9 0 1 10 9 0 1 11 2 9 0 13 1 11 11 2
69 10 9 0 1 10 9 15 13 1 10 0 2 4 7 15 13 2 13 1 10 12 1 10 12 1 11 3 9 1 9 15 13 10 0 9 1 9 1 10 9 1 10 11 2 3 13 1 9 0 7 3 0 9 1 15 13 10 9 2 10 9 1 9 7 10 9 1 9 2
33 10 9 1 15 9 10 9 3 1 10 9 0 4 13 1 10 9 11 11 7 11 11 1 10 9 2 10 11 11 11 11 2 2
29 3 15 1 10 9 1 10 9 13 10 9 7 9 2 10 0 9 7 10 9 1 10 9 2 11 2 16 13 2
69 15 13 2 16 1 9 1 10 11 11 1 11 1 11 11 2 1 12 1 11 2 15 12 2 12 2 16 10 9 13 10 9 1 9 0 4 13 3 1 10 9 1 10 9 1 10 9 7 9 1 10 9 1 10 9 1 10 9 2 3 13 1 10 11 1 11 1 11 2
32 10 10 9 1 9 13 9 1 10 9 0 1 9 1 11 2 7 13 9 1 10 9 1 10 9 1 9 1 9 1 11 2
44 10 9 13 0 7 3 0 2 7 10 9 13 16 3 3 15 13 1 10 9 0 1 10 9 2 7 10 9 4 13 1 10 0 9 1 10 9 1 10 9 1 10 9 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
21 4 13 1 10 11 11 1 11 7 15 13 1 10 9 1 0 9 7 0 9 2
18 3 1 10 9 1 11 15 13 0 3 15 1 10 12 9 1 11 2
21 1 9 15 13 10 9 1 10 9 1 10 9 13 1 11 1 12 2 13 3 2
23 15 13 13 1 10 9 1 12 9 7 13 1 12 5 1 10 9 1 10 9 2 11 2
23 15 4 13 1 11 7 10 9 7 13 3 2 7 16 13 1 10 9 3 2 1 3 2
18 10 9 13 10 0 9 0 7 10 0 9 0 13 10 9 11 11 2
16 1 12 13 1 10 9 0 1 10 11 11 2 1 11 11 2
35 15 13 1 10 9 1 10 9 10 2 11 11 11 2 1 10 15 15 13 1 10 9 1 9 2 13 1 15 10 9 1 9 7 9 2
17 10 9 13 3 1 10 9 1 9 7 9 16 15 13 1 9 2
17 9 0 13 10 9 16 4 13 1 9 0 1 9 10 9 0 2
28 11 3 13 13 1 10 11 11 16 3 13 12 9 7 10 9 1 11 15 13 2 1 15 10 11 1 11 2
32 4 13 15 2 3 2 9 1 9 2 9 1 9 2 7 9 1 9 2 1 10 9 1 9 1 13 10 9 13 0 3 2
44 1 9 0 2 3 15 13 1 16 10 9 13 2 11 13 10 0 9 1 10 9 1 10 9 2 7 10 9 12 1 10 9 2 15 16 15 13 10 9 1 9 3 0 2
17 1 12 15 13 10 9 1 10 9 0 13 1 10 9 1 12 2
35 13 0 10 9 2 13 10 9 1 9 7 9 0 2 13 1 10 9 16 15 13 10 9 1 10 9 1 3 15 15 13 1 10 9 2
64 10 0 9 16 13 1 10 9 1 12 5 1 10 11 11 1 11 11 2 11 11 2 1 10 9 13 2 11 0 12 5 11 2 2 3 15 13 1 10 11 11 1 11 11 12 2 11 11 2 1 10 9 2 9 11 1 8 2 11 2 1 12 5 2
23 1 10 9 1 10 9 10 9 13 1 10 11 15 13 2 3 2 1 10 9 15 0 2
38 10 9 1 16 10 9 0 1 11 15 13 1 9 1 10 9 1 9 2 13 16 1 10 9 1 10 9 10 9 1 11 4 13 10 3 0 9 2
19 15 13 2 13 15 16 15 13 2 13 10 9 7 10 9 13 3 0 2
13 13 0 7 13 3 0 1 11 2 11 7 11 2
10 13 10 9 11 11 7 11 1 11 2
33 3 2 1 0 1 10 9 0 1 9 0 1 10 11 11 2 15 13 9 0 13 1 10 9 1 10 9 0 7 10 9 0 2
13 10 9 1 11 15 13 1 11 2 11 1 12 2
39 1 9 1 12 13 10 0 2 11 1 10 9 1 9 1 9 1 9 2 1 10 15 13 15 1 10 9 0 7 0 7 1 10 9 15 13 10 11 2
8 2 13 10 11 1 10 9 2
21 9 2 10 9 0 1 10 11 11 1 10 11 11 1 11 2 15 13 1 11 2
28 10 9 0 2 12 2 10 9 0 15 13 1 10 9 2 10 9 0 1 10 15 4 13 10 9 1 11 2
28 3 10 9 1 10 11 2 9 3 13 2 7 11 2 9 3 13 2 2 13 10 9 1 9 1 10 9 2
9 13 9 1 11 1 13 10 9 2
41 3 3 7 15 13 10 9 10 9 1 9 15 13 0 7 10 0 9 16 13 0 1 11 13 1 10 9 1 9 1 12 9 10 9 3 0 1 13 10 9 2
51 7 13 1 10 9 1 10 9 2 3 3 13 16 3 13 9 1 13 1 10 9 10 9 2 2 10 9 2 16 13 10 9 2 1 13 15 3 13 15 2 7 12 2 7 12 2 2 13 11 11 2
41 10 11 11 11 11 13 1 9 1 10 9 7 9 1 10 9 1 10 9 13 13 0 9 2 1 9 1 16 10 11 1 11 4 13 10 9 1 10 9 0 2
24 10 9 1 15 1 9 0 2 1 9 2 15 13 1 13 15 1 9 0 2 13 10 9 2
29 10 9 0 16 13 10 9 2 13 1 10 9 0 2 4 13 16 13 10 9 3 0 7 13 1 10 9 0 2
18 10 12 1 11 1 12 2 9 11 2 11 7 11 13 1 10 11 2
39 10 9 1 9 2 10 9 1 11 3 15 13 7 10 9 15 13 1 9 15 10 9 4 4 13 1 10 10 9 1 9 1 13 15 1 13 1 15 2
18 2 1 10 9 15 13 0 2 16 10 9 13 10 9 7 10 9 2
49 1 10 9 2 11 11 13 10 9 1 2 10 0 9 1 0 9 2 1 10 0 9 1 11 11 2 16 13 10 9 1 10 0 9 1 10 9 1 10 11 11 2 11 11 7 10 11 2 2
32 10 9 13 1 10 12 9 7 13 0 1 10 10 9 1 10 9 2 10 0 9 1 10 9 4 13 1 10 11 1 11 2
17 1 9 11 15 13 1 11 7 11 2 1 10 15 13 1 9 2
9 2 10 9 13 2 13 10 9 2
3 9 9 0
38 1 10 9 2 11 11 13 1 10 11 1 11 11 2 7 3 4 13 7 13 10 9 2 9 0 13 1 10 11 11 7 13 2 4 13 1 9 2
51 10 9 0 2 13 1 15 9 1 10 9 12 2 13 1 10 9 1 10 9 13 1 13 15 1 10 9 2 7 10 11 1 11 4 13 1 13 10 9 7 13 1 10 9 10 9 1 13 10 9 2
27 13 10 9 0 1 12 9 2 8 2 0 1 10 9 11 12 8 12 1 10 9 1 9 1 10 9 2
10 10 9 1 9 0 0 13 10 9 2
22 13 10 9 0 2 3 15 13 3 15 16 13 10 9 7 10 9 3 13 15 0 2
26 10 9 2 13 1 13 10 9 1 10 9 2 13 10 9 3 0 1 10 9 2 1 10 9 0 2
9 10 9 13 16 15 13 1 0 2
18 1 0 7 1 11 2 10 9 1 11 13 15 3 3 7 10 9 2
40 3 1 12 9 1 9 1 10 9 1 9 13 7 9 0 2 13 16 15 13 10 9 0 1 10 9 7 13 10 9 0 1 10 9 2 10 0 9 0 2
14 15 13 9 1 10 9 2 11 11 11 2 11 2 2
17 11 4 13 10 9 1 10 11 15 7 1 9 7 9 1 9 2
28 1 10 9 2 10 9 13 15 1 10 0 9 16 13 10 9 1 10 9 1 3 13 1 9 1 9 0 2
50 11 15 4 13 1 9 1 10 9 1 9 0 2 13 1 0 9 1 11 7 11 2 7 13 13 10 9 1 0 9 1 7 15 15 13 10 9 1 9 1 10 12 1 11 12 13 1 10 9 2
26 15 1 10 9 7 9 4 13 1 10 0 11 2 1 11 11 2 11 11 11 2 13 1 10 9 2
22 15 13 1 9 0 7 8 2 0 7 13 1 10 9 1 11 7 1 10 9 11 2
66 1 10 9 2 13 10 0 9 1 10 9 2 13 1 10 9 2 1 10 9 0 2 10 9 7 9 1 10 9 2 2 1 3 13 10 9 1 10 9 0 2 2 2 15 13 10 9 1 10 9 3 16 15 13 10 0 9 16 13 1 9 1 9 7 9 2
31 13 10 9 2 1 9 1 12 11 13 10 9 1 11 11 12 2 1 10 9 1 10 9 2 7 4 13 1 10 9 2
22 13 10 0 9 1 9 2 9 2 13 7 9 0 16 13 10 0 9 1 10 9 2
32 10 11 1 10 11 4 13 10 9 1 11 11 11 11 16 13 3 10 11 1 10 11 2 13 1 10 9 0 1 9 0 2
35 10 9 13 3 1 9 1 11 15 13 1 13 1 10 9 0 2 10 9 3 13 15 1 10 9 3 3 15 13 9 2 9 7 9 2
32 1 10 12 9 13 1 10 10 9 2 13 15 1 0 1 11 2 3 15 13 1 10 9 7 15 13 1 10 9 1 9 2
16 1 15 2 1 9 2 10 0 9 1 9 0 9 1 11 2
46 1 12 15 13 10 9 1 10 9 1 10 9 1 10 9 1 13 10 9 1 10 9 2 16 4 13 1 10 9 2 1 10 0 9 1 10 9 13 1 10 10 9 1 10 9 2
15 13 1 10 9 1 9 0 2 13 10 9 1 9 0 2
12 10 9 8 8 1 10 9 13 1 5 12 2
9 13 1 11 2 9 1 11 2 2
15 16 11 13 1 10 9 3 13 11 2 13 16 13 0 2
43 10 11 1 11 4 13 1 9 10 0 9 0 16 13 1 10 9 1 9 0 13 9 2 1 10 9 2 16 4 13 1 10 9 0 2 4 13 10 9 1 10 9 2
30 1 10 9 3 13 10 9 7 10 9 0 3 4 3 13 3 1 10 9 1 10 9 11 11 1 10 8 11 11 2
36 11 13 1 10 10 9 1 10 9 0 0 2 10 15 13 1 9 0 7 13 1 10 12 1 11 1 12 2 3 15 13 10 0 11 11 2
22 15 4 4 13 1 10 9 7 10 9 16 13 10 9 7 3 13 3 9 7 13 2
13 1 10 9 12 0 10 9 1 9 13 1 11 2
15 11 13 3 10 9 1 9 13 1 2 11 8 11 2 2
27 1 10 9 1 9 2 10 9 13 10 9 1 10 9 2 7 13 10 9 1 9 0 1 10 9 0 2
10 10 9 0 3 16 13 9 0 0 2
36 10 9 13 10 9 0 2 15 16 3 13 1 10 9 2 13 15 1 10 0 9 1 10 9 1 10 9 2 1 3 1 12 9 1 9 2
30 3 3 2 13 16 1 10 9 13 10 11 1 10 9 15 4 13 1 10 9 10 9 1 13 9 16 13 10 9 2
45 1 10 9 0 11 2 11 13 1 10 0 9 7 15 13 1 12 1 10 9 11 2 15 15 13 16 11 2 11 15 13 1 10 9 1 10 9 1 9 1 9 7 9 0 2
17 11 13 10 9 1 10 9 1 11 11 13 1 10 12 5 9 2
9 1 12 4 13 1 11 1 11 2
12 13 13 9 7 10 9 0 3 15 4 13 2
25 10 9 16 15 13 1 9 1 10 9 12 13 10 9 1 9 1 11 13 1 12 7 12 9 2
46 7 3 15 13 10 9 0 2 10 9 15 13 1 9 1 10 9 0 2 1 10 0 9 9 2 9 7 9 0 15 4 13 1 10 11 2 1 0 9 1 4 13 0 7 0 2
14 10 11 12 15 13 1 9 10 12 1 11 1 12 2
13 11 7 8 2 11 13 15 1 10 9 1 11 2
22 1 11 1 10 12 2 13 1 10 9 16 11 4 13 1 11 11 1 10 9 12 2
18 4 13 10 0 9 1 9 2 1 0 9 2 7 10 9 0 0 2
19 10 9 4 13 1 12 1 10 11 1 12 9 7 4 13 1 12 9 2
14 3 2 1 10 9 1 11 3 13 1 9 10 9 2
17 4 13 10 9 1 9 12 1 12 1 9 1 9 1 11 11 2
37 10 9 15 4 13 13 10 9 1 11 11 1 9 1 10 9 12 7 10 9 1 10 11 2 1 9 3 0 7 9 1 9 1 10 9 12 2
6 2 3 13 10 9 2
11 1 15 15 16 15 13 13 16 15 13 2
11 9 2 0 8 2 8 2 8 2 8 2
18 9 1 10 9 0 2 3 15 13 10 9 2 10 9 7 10 9 2
34 10 9 0 13 16 10 9 0 1 10 9 13 1 9 1 10 11 11 1 13 15 1 11 2 7 13 1 9 1 0 9 1 11 2
10 13 1 10 9 8 2 8 7 8 2
25 15 4 13 3 10 9 1 10 9 1 10 9 7 3 4 13 15 10 9 2 3 0 1 15 2
22 10 9 13 0 1 10 9 11 2 10 15 13 9 1 9 1 9 0 1 10 9 2
24 10 9 13 9 1 3 13 10 9 1 13 15 1 9 0 2 1 10 0 9 7 10 11 2
35 13 1 10 9 1 10 9 2 10 15 4 13 2 0 2 1 10 9 16 15 13 0 2 3 16 15 15 4 13 7 13 1 10 9 2
13 10 9 0 13 10 9 1 9 1 10 10 9 2
46 13 16 10 9 3 3 15 13 1 15 0 1 10 0 9 1 9 1 10 9 2 1 9 13 9 2 9 7 9 1 10 9 2 1 15 15 15 15 13 1 0 9 1 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
22 11 13 10 10 9 7 13 3 10 9 1 16 11 7 11 3 15 13 1 10 9 2
38 1 10 9 1 12 9 2 10 9 13 1 10 9 0 7 3 0 0 9 0 1 10 15 15 13 9 13 1 10 9 7 13 1 10 9 1 11 2
20 13 10 11 10 11 1 10 9 2 13 7 13 10 9 7 9 13 9 0 2
29 10 9 16 15 4 13 2 7 16 3 4 13 1 9 1 3 16 13 9 1 10 11 1 11 1 10 10 9 2
20 10 9 15 13 10 11 1 11 1 10 11 11 1 10 10 9 1 10 11 2
38 12 9 3 1 11 11 15 13 1 10 0 9 1 15 13 10 11 11 1 9 0 1 11 11 2 11 4 13 10 9 1 15 16 13 1 10 11 2
36 10 12 1 11 1 10 0 9 2 15 13 10 9 0 1 10 9 1 15 10 9 13 9 0 1 10 9 16 10 9 13 0 1 10 9 2
30 1 10 9 0 13 9 0 1 10 0 9 0 1 10 11 2 0 1 10 9 1 11 2 15 1 10 9 1 11 2
21 1 3 3 12 9 2 10 9 4 13 10 9 8 2 8 2 1 9 1 9 2
54 10 11 1 11 11 13 10 9 1 11 2 13 1 10 9 1 10 11 1 10 11 2 1 10 9 0 1 0 9 1 10 9 1 10 11 2 1 10 9 1 11 2 9 0 1 11 7 11 7 9 0 1 11 2
57 1 10 9 0 2 3 3 13 10 9 0 2 11 11 7 10 9 11 11 2 13 3 10 9 2 11 2 11 7 11 2 10 16 13 10 0 9 0 7 0 2 7 16 13 3 0 9 1 10 9 1 10 9 0 11 11 2
28 10 9 1 10 9 13 1 10 9 1 9 1 10 9 1 11 11 2 3 16 11 13 3 10 3 0 9 2
22 13 1 11 2 11 11 2 10 12 1 11 1 12 2 9 1 11 11 7 11 11 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
20 1 10 11 13 9 7 0 9 1 9 1 10 9 2 3 1 13 1 11 2
28 10 9 1 10 9 15 13 10 0 9 1 9 2 7 15 1 10 9 15 13 1 10 9 7 1 10 9 2
33 0 2 16 3 15 4 13 2 4 4 7 13 15 1 7 10 9 13 1 9 7 3 4 13 10 9 16 4 7 4 13 15 2
11 3 13 9 1 13 2 7 13 3 9 2
69 1 9 2 1 10 9 0 15 4 13 10 9 1 10 9 7 10 9 1 10 9 7 4 7 13 10 9 1 13 10 9 13 1 9 10 9 2 13 13 2 3 9 1 9 2 9 2 13 3 0 2 9 2 7 10 9 2 9 0 2 13 10 9 0 1 10 9 0 2
31 1 10 9 2 13 2 13 1 9 10 9 0 16 15 4 13 1 11 2 13 1 10 9 0 7 10 9 1 9 0 2
18 13 1 10 9 1 10 9 15 13 2 13 15 1 10 9 7 9 2
28 13 9 2 1 10 9 2 1 10 10 9 1 10 9 1 10 9 0 2 10 9 7 10 9 2 12 2 2
60 1 10 9 1 10 0 9 2 13 9 10 0 11 11 11 11 2 3 13 3 1 12 9 1 10 10 9 2 3 1 10 0 9 1 3 1 12 9 1 0 9 2 9 16 13 10 9 1 10 9 13 1 10 9 1 10 9 1 11 2
29 13 10 0 9 1 11 2 12 2 2 15 13 1 10 9 1 9 7 10 9 0 2 0 1 11 11 1 11 2
11 10 0 9 4 3 13 1 9 1 9 2
20 10 9 12 13 15 16 3 9 13 1 10 9 13 1 10 12 1 10 9 2
17 11 13 10 9 0 2 3 15 13 15 1 10 9 1 10 9 2
14 13 9 0 15 4 13 7 4 13 13 15 10 9 2
24 13 10 9 0 7 0 16 15 13 1 13 9 7 3 9 2 9 2 9 7 3 0 9 2
25 13 9 1 9 0 16 13 1 9 0 10 9 2 10 9 2 7 10 9 0 2 10 9 2 2
13 3 15 13 1 10 9 1 11 1 10 11 12 2
22 13 1 9 1 9 1 15 1 10 9 0 3 0 1 10 9 2 10 9 1 11 2
13 11 11 2 11 11 7 11 11 13 9 1 9 2
28 11 11 15 13 1 10 9 1 9 1 10 11 2 9 0 1 10 11 1 10 9 2 7 10 9 7 9 2
27 15 11 2 3 7 3 4 13 1 10 10 9 1 11 3 13 3 0 7 15 4 13 1 3 0 9 2
32 15 1 10 9 0 2 11 11 2 16 13 1 12 1 10 9 2 13 16 11 13 10 9 1 10 15 10 9 3 15 13 2
20 11 15 13 9 8 2 0 2 3 16 10 9 11 13 1 11 7 1 11 2
8 13 1 9 7 13 1 9 2
30 10 9 0 1 11 11 2 13 16 13 0 15 15 13 1 10 9 2 3 16 10 9 3 0 13 1 9 10 9 2
21 13 10 9 1 10 9 1 9 0 1 10 9 1 9 1 9 1 10 9 0 2
31 15 1 10 9 16 10 11 13 13 13 10 9 1 10 16 10 9 4 13 10 9 1 9 1 13 3 1 10 9 0 2
7 15 13 3 1 13 9 2
22 3 13 9 1 16 11 4 13 1 10 11 1 11 3 1 7 11 15 13 1 0 2
21 10 9 15 13 10 0 9 16 2 1 12 2 13 1 9 10 9 1 9 9 2
19 13 9 1 10 11 11 1 10 11 1 12 2 4 13 9 0 1 12 2
22 10 11 2 9 1 10 9 1 11 11 2 9 1 11 11 1 11 2 11 2 11 2
59 3 3 3 3 15 13 16 15 13 16 10 12 9 13 1 13 1 10 9 0 11 11 2 3 7 3 1 10 11 11 7 11 11 1 2 11 2 11 11 2 13 1 13 10 9 1 10 9 1 10 9 1 9 1 10 9 9 11 2
15 1 9 0 2 15 13 9 0 1 11 2 11 7 11 2
14 11 11 13 10 9 1 9 0 9 1 10 9 11 2
5 2 9 7 9 2
25 1 9 1 10 9 2 10 9 11 13 16 11 2 13 15 3 0 1 13 11 7 10 9 2 2
69 3 2 3 3 1 13 15 13 9 2 1 16 15 13 9 0 2 1 10 9 0 0 1 10 9 0 1 9 1 9 15 11 11 15 11 2 13 1 10 9 7 9 1 10 9 0 2 1 10 16 10 9 1 9 13 9 1 10 9 0 7 9 1 10 9 1 10 9 2
28 10 11 11 13 10 9 1 9 1 11 11 2 13 1 10 11 1 10 11 1 11 10 12 1 11 1 12 2
22 13 1 10 9 1 10 0 9 1 13 10 9 1 0 9 3 7 3 1 10 11 2
20 10 9 11 1 9 13 2 9 2 9 2 9 2 9 2 9 7 9 2 2
28 10 9 1 10 9 10 9 11 12 13 1 10 10 9 1 9 2 1 3 13 1 9 2 1 10 9 0 2
54 11 11 11 1 10 11 11 13 10 9 1 2 2 7 9 1 11 0 1 2 11 2 7 2 11 11 11 10 11 2 2 7 13 1 10 9 1 16 11 2 2 1 9 13 3 13 15 1 10 9 1 9 2 2
16 10 9 3 0 2 3 13 0 7 3 13 10 9 1 9 2
43 1 10 11 1 10 11 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
26 1 10 9 10 9 11 11 15 13 1 10 9 1 10 8 1 9 1 9 1 10 9 0 1 11 2
29 16 2 1 10 9 1 11 2 4 1 13 1 10 9 1 11 2 13 1 0 9 10 9 1 11 7 13 0 2
20 13 10 10 9 1 10 10 9 16 13 10 9 0 1 13 13 10 9 0 2
18 3 2 16 10 11 3 4 13 10 9 2 10 9 13 1 13 9 2
11 3 7 10 8 13 9 2 8 13 0 2
11 3 1 9 10 9 3 13 10 9 0 2
51 10 9 1 10 15 15 13 9 13 1 9 0 7 15 13 13 1 10 9 1 10 9 1 11 2 12 5 1 9 1 10 11 11 2 16 13 1 10 9 1 9 1 10 11 2 10 11 7 11 11 2
15 9 0 1 10 9 13 1 10 11 11 11 2 1 9 2
20 11 11 13 10 9 1 9 1 10 9 1 10 11 1 10 9 1 10 11 2
21 15 15 13 1 10 9 0 2 1 11 11 10 9 0 13 1 0 9 10 9 2
74 1 10 9 2 13 10 9 13 1 9 0 1 10 9 11 12 1 11 2 13 1 10 9 13 10 11 12 2 1 10 16 15 13 10 9 1 9 7 9 1 10 9 1 10 9 11 7 10 9 1 10 9 0 1 10 9 1 10 9 0 0 2 8 2 2 13 1 10 9 1 11 1 11 2
40 1 9 1 13 1 10 9 1 9 1 10 9 2 10 9 1 11 15 13 3 13 9 1 9 1 13 10 9 1 10 9 1 10 9 2 13 1 10 9 2
36 10 9 4 13 1 10 9 12 2 1 9 16 13 1 10 9 1 11 11 11 2 9 1 10 9 2 7 11 11 11 2 9 0 1 11 2
20 10 9 0 4 13 1 3 15 9 1 10 9 1 15 2 1 10 12 9 2
22 10 11 11 1 10 11 11 13 10 12 1 11 11 1 10 11 11 1 10 11 11 2
26 15 13 16 1 9 1 10 9 10 9 0 1 11 13 1 10 9 2 13 10 9 0 1 12 9 2
16 11 11 13 10 9 1 10 11 11 1 10 9 12 2 12 2
39 16 13 9 2 13 10 9 0 16 10 9 1 10 11 11 4 13 1 9 0 1 12 1 12 7 10 9 15 13 1 10 9 1 10 11 11 1 12 2
20 10 9 13 1 9 9 0 2 1 9 1 9 1 10 9 0 1 10 9 2
12 7 13 2 2 13 16 3 13 9 1 9 2
17 10 9 1 10 9 0 4 13 1 10 9 1 9 1 10 9 2
32 1 16 15 13 15 2 10 11 4 13 0 1 13 1 12 9 2 12 9 2 5 2 7 13 15 1 9 13 1 12 8 2
48 1 10 11 11 15 13 10 9 0 1 10 9 1 10 9 9 2 8 2 2 16 4 13 15 1 9 2 1 1 10 9 1 10 9 11 16 13 10 9 1 2 11 9 1 9 0 2 2
36 13 11 10 12 1 11 1 12 3 13 10 9 2 13 10 0 1 10 9 1 10 9 2 11 11 11 2 1 15 15 11 4 13 1 0 2
5 10 9 13 9 2
39 10 9 13 0 1 10 9 13 1 10 9 0 0 1 10 9 1 10 11 1 11 1 9 1 10 9 12 2 7 13 3 10 9 1 10 11 1 11 2
33 10 9 13 10 9 1 15 2 7 10 9 2 16 3 15 4 13 1 9 13 0 10 9 16 15 13 1 10 11 1 11 11 2
36 4 13 1 10 9 0 11 1 9 1 11 7 13 10 0 9 1 9 16 15 13 1 10 11 0 2 3 1 15 1 11 2 11 7 11 2
19 10 9 11 13 12 9 2 10 9 0 2 16 13 10 9 1 10 9 2
39 13 7 13 3 12 1 10 9 1 9 1 10 9 11 11 7 11 11 13 2 10 11 2 2 2 10 11 15 11 1 11 2 7 2 10 10 11 2 2
12 10 9 7 9 13 1 10 9 0 11 11 2
23 10 9 1 10 9 0 13 3 0 16 10 0 9 1 10 9 15 13 1 9 1 11 2
12 9 1 10 9 4 13 1 10 9 7 9 2
10 2 1 3 13 10 9 1 10 9 2
21 10 9 4 13 10 12 1 11 1 12 2 7 3 13 0 1 10 12 1 11 2
4 4 13 3 2
17 10 9 13 10 0 9 2 16 15 13 0 1 10 9 1 11 2
22 11 10 11 13 3 1 10 0 9 1 11 2 13 10 9 2 10 9 7 10 8 2
50 1 9 1 15 16 4 13 1 9 0 2 1 10 15 13 0 9 1 9 1 10 9 2 3 2 1 15 1 10 9 1 11 2 10 9 1 10 9 7 10 9 2 2 10 9 15 13 3 0 2
28 11 13 10 9 0 13 1 10 9 1 9 11 11 2 1 10 9 1 11 11 2 9 1 11 11 2 11 2
19 10 9 1 10 0 9 2 9 1 15 2 13 16 10 9 13 3 0 2
28 7 11 3 4 13 1 11 0 15 3 9 7 10 9 1 10 9 15 13 1 0 9 1 10 9 1 13 2
17 11 11 11 11 13 10 12 1 11 1 12 1 10 9 1 11 2
14 3 1 13 9 1 10 9 10 9 13 10 11 11 2
15 3 15 4 13 9 7 9 0 2 8 2 2 9 2 8
40 3 10 9 1 9 1 10 9 15 13 1 9 13 1 10 9 13 10 9 1 9 1 13 2 13 1 10 0 9 13 1 12 9 1 10 9 1 10 9 2
46 10 9 0 13 2 9 2 9 2 9 1 8 8 2 10 9 1 12 9 1 9 2 9 11 1 9 0 2 11 11 12 2 9 12 5 8 7 9 11 12 1 10 9 1 11 2
14 15 13 1 11 2 9 1 10 9 11 2 11 2 2
16 1 10 9 2 10 9 13 10 9 3 1 9 1 10 9 2
40 16 13 10 9 2 16 13 1 3 1 12 9 1 9 1 10 9 2 10 9 13 1 13 1 10 0 12 1 11 1 10 9 0 1 11 1 10 9 11 2
12 10 9 16 13 10 9 1 9 13 10 9 2
18 10 9 3 13 1 9 1 9 1 10 9 2 1 9 13 9 0 2
21 1 10 12 2 10 2 11 2 15 13 1 10 9 1 11 11 7 13 10 9 2
46 15 13 1 8 13 10 9 0 1 10 9 0 7 9 1 9 0 2 3 1 13 10 9 0 1 10 9 7 13 15 9 1 10 9 1 9 2 3 7 13 10 9 1 9 0 2
8 9 13 1 10 11 1 11 12
17 11 2 0 1 10 9 1 10 9 2 15 15 13 1 10 9 2
29 3 12 9 0 4 13 1 11 11 1 9 1 10 11 1 13 10 9 0 3 13 1 10 9 0 1 10 9 2
25 1 10 9 1 12 13 13 9 3 1 4 13 10 9 2 1 13 1 13 10 9 7 10 9 2
23 10 0 9 3 1 11 11 13 10 11 1 10 11 2 15 1 10 0 9 1 11 11 2
26 11 13 3 10 9 1 9 1 10 9 16 3 15 13 11 1 10 9 2 16 10 9 3 3 0 2
31 10 9 2 13 1 11 11 2 9 1 10 11 2 2 4 13 1 10 9 1 10 9 1 10 0 9 0 1 10 9 2
24 10 0 9 4 13 9 1 10 11 1 11 11 7 1 12 13 10 11 1 10 11 1 11 2
21 10 9 1 11 2 10 3 0 7 0 1 10 9 0 1 11 2 13 1 9 2
33 15 13 1 0 9 1 10 11 11 11 1 11 1 12 2 7 4 13 10 12 1 11 1 12 1 5 12 3 1 9 7 9 2
18 13 1 11 11 7 10 14 2 9 11 11 2 11 11 2 11 11 2
32 13 9 1 10 9 1 11 2 10 9 1 11 2 9 1 11 2 10 9 1 11 7 1 9 13 9 1 10 9 1 11 2
18 1 10 9 15 13 10 0 9 0 13 1 10 9 1 10 9 0 2
20 13 3 10 9 2 10 9 13 16 10 0 9 11 11 2 13 0 1 9 2
41 1 1 10 0 9 13 16 10 9 13 1 10 9 16 13 1 10 9 2 9 0 2 3 3 0 2 16 15 13 1 10 9 1 10 9 7 13 2 9 2 2
13 10 9 1 9 13 9 1 0 9 1 10 9 2
16 3 13 3 7 3 4 13 3 13 1 15 16 3 15 13 2
48 10 9 8 2 12 4 4 3 13 7 13 1 10 11 2 13 2 1 13 1 9 13 3 1 10 9 0 2 1 11 2 1 10 9 0 1 11 2 3 13 9 13 1 11 7 11 11 2
12 10 9 13 15 4 13 10 0 9 1 9 2
27 1 10 9 1 10 9 1 11 11 1 11 2 12 2 2 13 7 15 13 3 10 9 0 1 10 9 2
8 11 15 13 13 1 10 9 2
33 1 10 9 1 9 1 10 9 0 0 1 10 11 2 10 8 9 13 16 2 16 10 9 13 3 0 2 3 15 13 10 9 2
29 13 9 13 7 13 1 10 9 1 10 9 1 9 2 9 7 9 0 7 0 1 10 9 1 10 9 1 11 2
22 10 9 0 15 13 1 13 1 10 9 0 2 7 10 9 0 13 9 1 10 9 2
33 11 11 13 1 10 9 1 11 2 7 11 11 13 10 9 1 10 9 1 11 2 15 1 10 9 1 10 9 1 10 9 0 2
21 13 10 9 0 1 10 9 1 13 10 9 1 10 9 0 1 10 15 15 13 2
21 3 2 3 4 13 3 2 16 13 10 9 0 7 10 9 0 2 3 15 13 2
46 15 1 10 9 13 10 9 0 13 11 11 2 1 15 10 9 15 13 10 9 13 9 1 10 11 1 10 11 0 2 9 1 9 0 16 13 1 15 9 7 9 1 10 9 2 2
30 10 9 0 4 3 13 1 9 2 13 13 15 13 1 10 9 0 0 2 2 7 13 1 9 2 13 13 3 2 2
8 11 15 13 13 1 10 9 2
5 13 0 1 11 2
24 1 11 1 12 15 13 1 11 11 1 11 1 13 10 9 11 11 11 11 13 1 11 11 2
24 3 15 13 1 10 9 1 9 1 10 9 0 1 9 1 10 9 12 7 9 1 10 12 2
21 10 9 3 0 13 9 1 10 9 3 16 10 0 9 1 11 11 13 13 9 2
16 10 9 0 15 13 13 3 10 9 7 13 0 9 10 9 2
19 10 11 11 2 7 11 2 11 2 13 10 9 1 10 9 0 1 11 2
38 10 9 13 10 9 7 9 1 10 9 1 10 12 9 13 3 8 10 9 7 13 1 10 9 10 2 0 9 7 9 2 1 10 9 1 10 9 2
13 10 9 1 9 13 1 12 8 2 5 5 5 2
28 10 9 13 1 10 9 1 9 1 10 9 1 10 9 7 10 9 1 10 9 16 13 10 9 1 10 9 2
33 7 10 9 1 11 11 13 16 1 12 9 13 1 10 9 1 10 9 1 10 9 1 13 1 10 9 0 1 10 9 1 11 2
28 1 12 2 1 10 11 1 11 2 11 13 10 0 9 2 7 1 10 9 1 11 7 1 10 11 1 11 2
46 4 13 10 12 1 11 1 10 12 1 10 9 1 11 2 11 11 7 10 9 1 10 9 1 11 2 11 11 2 16 15 13 10 0 9 1 10 9 13 1 9 1 10 9 0 2
28 10 9 1 10 11 13 1 12 2 16 13 10 0 9 2 1 10 15 15 13 1 13 10 11 1 10 11 2
18 11 11 2 11 2 12 1 11 1 12 2 13 10 9 0 1 9 2
15 11 2 9 1 11 2 7 11 2 9 1 11 7 11 2
14 3 13 10 9 13 10 9 2 7 3 13 3 3 2
37 1 13 1 10 9 11 13 1 10 9 1 10 0 9 7 15 13 1 10 9 11 11 2 1 10 15 13 1 10 9 11 11 13 1 10 9 2
33 10 9 15 13 1 10 9 1 9 0 2 1 3 15 13 9 7 11 2 4 13 10 9 0 16 13 1 10 9 12 7 12 2
59 10 11 1 11 2 1 9 2 11 11 2 7 11 1 11 2 1 9 2 11 11 11 2 15 13 1 10 9 11 12 1 11 7 10 9 1 10 11 1 11 11 11 10 12 1 11 1 12 2 1 10 9 1 11 2 0 11 2 2
3 9 11 2
20 9 0 4 4 13 1 10 9 2 7 10 9 1 10 9 4 1 13 15 2
28 10 9 0 4 13 10 9 1 10 0 7 0 9 2 3 1 10 9 1 9 0 0 1 10 0 9 0 2
38 10 0 9 1 9 13 10 2 9 0 1 10 9 2 2 10 9 1 10 9 0 2 7 10 9 1 9 16 15 13 1 10 9 1 9 3 0 2
20 3 1 10 9 0 2 13 9 0 13 1 10 9 1 9 1 10 9 0 2
5 11 15 4 13 2
17 16 13 2 13 10 0 9 1 11 3 13 0 9 0 2 0 2
17 11 11 13 1 11 2 11 9 1 11 11 7 10 9 11 11 2
34 3 13 8 2 9 1 9 2 9 2 9 2 8 2 9 2 9 2 8 2 9 1 9 0 1 10 10 9 7 10 9 1 9 2
16 15 13 1 10 12 1 2 11 11 11 2 2 11 2 11 2
36 13 9 0 2 3 9 2 1 9 1 9 1 15 3 9 2 3 13 9 7 9 13 1 10 9 2 9 2 9 7 3 3 1 10 9 2
19 10 9 15 13 1 9 1 9 16 13 1 10 9 1 10 9 1 9 2
8 10 9 13 10 9 1 11 2
43 13 1 10 9 1 9 1 11 1 11 2 12 2 2 11 11 2 12 2 2 11 11 11 11 2 12 2 2 11 11 11 2 12 2 7 11 11 11 11 2 12 2 2
43 11 11 2 2 11 2 12 1 11 1 12 2 11 11 2 12 1 11 1 12 2 13 10 9 7 9 0 13 9 0 3 1 10 9 0 1 11 1 10 9 1 12 2
61 11 11 2 9 1 10 9 11 11 11 11 2 7 11 11 2 9 1 10 9 11 1 11 2 11 2 2 13 1 9 10 9 1 13 10 11 12 1 10 9 3 0 1 10 16 13 11 12 2 10 11 12 13 10 9 1 10 11 11 2 2
35 10 12 11 11 11 1 11 2 11 12 7 10 11 1 11 1 11 11 3 4 13 10 9 1 9 1 10 10 9 16 13 0 1 13 2
23 13 10 9 2 9 0 7 9 1 9 2 16 15 13 1 10 9 1 9 1 9 13 2
27 3 1 10 9 2 12 2 11 4 13 1 11 1 11 10 9 1 10 9 1 10 9 1 10 9 0 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
14 15 1 10 9 1 9 1 9 0 13 10 9 0 2
31 1 9 0 16 13 2 11 3 3 4 13 10 9 0 2 8 8 16 13 1 13 1 8 7 15 13 10 15 16 13 2
24 13 3 1 12 9 1 7 10 9 4 13 1 16 0 7 1 12 1 12 9 1 13 9 2
32 1 9 1 10 9 15 13 9 0 1 0 9 2 16 13 1 10 9 10 9 7 15 4 13 1 10 9 1 10 9 12 2
12 13 10 0 9 0 16 15 13 2 10 9 2
14 13 3 1 10 9 9 7 1 10 11 11 11 11 2
29 1 9 0 2 10 9 13 10 0 9 0 1 10 11 2 1 10 9 15 13 10 9 2 16 13 10 9 0 2
16 10 9 0 15 13 1 10 9 0 7 10 2 0 9 2 2
25 3 1 11 11 11 13 15 1 10 0 9 1 13 10 9 1 10 9 0 1 9 1 9 0 2
51 1 9 1 10 9 1 9 0 2 10 9 1 11 7 11 15 13 0 2 7 11 15 13 1 10 9 0 2 1 9 0 1 10 9 0 2 0 1 12 2 7 13 10 9 0 0 1 10 11 11 2
15 13 1 10 9 1 10 9 2 3 1 10 9 10 9 2
31 10 9 15 13 10 9 1 11 13 10 9 1 9 1 13 10 9 0 2 13 9 1 9 1 10 9 1 11 7 11 2
19 10 9 1 11 1 10 11 7 11 13 10 9 0 9 0 7 10 9 2
17 1 10 9 4 9 1 11 11 1 0 9 7 9 1 10 9 2
14 3 13 1 15 10 11 11 2 9 1 10 9 11 2
14 10 9 13 15 1 10 3 0 1 15 13 1 11 2
14 1 12 13 10 12 9 1 10 11 1 11 1 11 2
34 10 9 0 15 13 1 10 9 11 11 11 11 2 1 11 2 15 13 16 15 13 1 12 1 10 9 0 7 1 9 1 9 0 2
60 1 10 9 0 2 13 3 1 10 9 1 10 9 7 10 9 11 2 3 10 12 0 9 1 11 11 2 10 0 11 11 7 3 2 10 12 1 11 1 12 15 13 10 9 1 10 9 2 13 3 3 1 11 11 1 9 1 11 12 2
11 10 9 1 10 9 13 1 10 9 0 2
6 10 9 13 3 0 2
16 15 4 13 1 9 0 16 13 10 9 1 9 13 1 9 2
35 10 3 9 2 11 11 11 11 2 13 1 11 11 2 11 11 7 11 11 1 13 9 15 4 13 1 10 9 1 10 9 1 10 9 2
17 13 16 13 1 11 2 1 15 15 3 13 15 1 13 1 11 2
35 12 9 2 12 9 7 12 9 3 1 10 9 7 12 9 2 12 1 12 1 9 2 2 12 9 2 12 9 7 12 9 9 1 11 2
27 1 10 9 2 13 1 10 9 16 15 13 1 9 1 10 9 0 7 15 16 15 13 1 15 3 0 2
34 8 8 13 10 9 1 10 9 1 9 8 8 7 8 8 11 15 4 13 1 9 1 12 9 1 9 0 2 0 2 0 7 9 2
20 10 0 9 2 9 1 11 1 10 11 2 15 13 3 1 9 1 10 9 2
19 11 11 2 11 2 11 13 10 9 0 3 13 1 10 0 9 1 9 2
16 15 13 1 10 11 11 0 2 10 11 11 7 11 11 11 2
2 13 2
22 11 13 10 9 0 1 16 10 9 15 4 13 1 15 0 1 1 10 9 1 11 2
13 10 9 15 4 13 1 10 9 7 1 10 9 2
49 10 9 1 10 9 1 11 11 11 11 7 11 11 2 15 1 10 3 0 9 1 10 11 11 2 13 1 10 9 12 2 16 10 0 9 1 9 11 11 4 13 1 10 9 1 11 11 11 2
17 1 9 2 13 10 0 9 1 15 16 13 1 10 9 1 11 2
39 13 16 10 9 0 0 1 9 0 4 13 15 1 10 9 1 9 0 1 0 9 2 15 13 1 10 9 1 11 2 11 10 9 7 9 1 10 9 2
20 1 10 9 1 11 2 8 2 15 13 1 10 9 2 11 7 11 2 12 2
17 3 1 12 9 0 1 9 7 13 16 10 12 9 0 1 9 2
31 10 9 0 4 13 1 10 9 0 7 11 13 10 10 9 15 4 13 2 1 11 7 10 9 1 10 9 1 10 11 2
18 15 15 13 1 9 1 9 7 10 9 0 4 13 0 1 3 9 2
33 10 9 3 1 10 11 11 1 11 1 13 1 12 9 0 10 9 1 9 0 1 10 9 4 13 10 9 0 1 10 9 0 2
12 3 1 9 10 9 4 4 13 1 10 9 2
13 10 0 9 1 9 13 9 1 10 9 0 0 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
34 1 9 2 11 2 3 13 10 9 1 9 1 9 1 9 1 9 7 10 9 1 10 0 9 0 1 11 2 3 13 9 7 9 2
12 15 4 13 9 1 9 2 13 1 10 9 0
26 10 9 13 11 11 2 10 9 1 10 9 0 9 1 10 9 1 11 11 2 7 10 9 11 11 2
22 1 10 9 13 1 12 9 7 3 10 10 9 15 13 13 10 9 1 11 1 15 2
24 3 13 1 10 9 10 0 9 1 2 11 2 2 16 1 10 9 15 13 1 10 0 9 2
26 1 13 10 12 9 0 3 1 10 9 2 10 1 10 9 7 10 1 10 11 2 3 3 13 0 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
30 1 10 10 9 0 1 10 9 2 11 4 3 13 1 10 0 9 1 11 11 2 10 15 15 13 3 1 10 11 2
12 10 9 1 9 1 10 9 13 1 9 12 2
48 16 10 9 15 13 1 9 7 1 9 1 10 9 0 2 3 1 10 11 1 10 11 7 10 9 1 11 2 10 11 13 3 10 9 1 9 0 13 1 10 9 2 13 3 1 9 0 2
21 1 10 9 10 9 13 1 9 10 9 1 10 9 7 10 9 1 10 9 0 2
12 13 3 7 11 7 11 11 13 13 1 11 2
19 10 9 4 13 1 12 1 10 11 11 1 11 11 7 11 2 11 2 2
20 1 11 1 12 11 11 7 11 11 13 10 9 1 11 1 10 11 1 11 2
39 13 15 10 9 1 10 11 13 1 10 9 1 3 15 2 1 15 1 4 13 1 11 2 9 16 4 13 1 10 8 2 9 2 13 1 10 9 0 2
51 1 10 9 2 10 9 13 1 13 10 0 9 1 10 0 9 1 10 11 1 10 11 7 4 13 1 7 15 1 11 13 1 0 9 2 1 9 0 1 13 16 10 10 9 0 13 1 10 9 0 2
42 1 12 13 10 9 1 10 9 1 10 11 1 11 11 2 11 2 2 1 10 15 13 10 9 0 1 9 1 10 9 1 11 1 11 7 1 10 9 0 1 11 2
32 1 9 1 10 9 3 13 13 10 9 2 1 10 9 1 10 9 0 2 9 7 9 0 2 9 1 9 2 1 10 9 2
13 3 2 13 15 1 10 9 3 0 1 10 9 2
36 10 9 0 2 4 13 9 1 16 1 10 9 1 10 9 7 9 1 9 2 10 9 13 10 9 1 9 7 9 1 10 9 1 9 0 2
27 13 10 9 1 11 1 12 9 2 16 3 4 13 12 5 9 2 10 0 9 16 13 1 10 12 9 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
23 10 9 1 10 11 13 1 10 9 0 9 0 1 7 13 15 16 3 13 1 10 9 2
60 10 0 12 1 11 2 10 9 1 10 11 13 9 1 10 11 11 1 11 2 16 11 1 10 11 2 10 11 7 10 9 11 13 16 13 9 1 9 1 10 9 16 13 1 10 9 10 9 1 13 7 3 10 9 1 9 1 10 9 2
15 15 13 9 1 10 9 1 9 16 3 13 13 10 9 2
48 1 10 9 1 13 1 10 9 1 10 9 1 10 9 0 7 10 9 2 5 13 10 0 9 1 10 16 10 9 4 13 10 9 0 7 0 1 9 2 9 7 9 13 1 10 9 0 2
23 4 13 15 16 10 9 1 11 2 13 10 9 0 2 15 13 1 10 9 1 9 0 2
26 1 12 2 13 1 10 11 1 13 1 11 1 11 11 2 16 3 4 13 1 11 11 2 1 12 2
19 10 9 4 13 3 0 1 15 15 13 10 9 2 13 16 15 13 0 2
12 10 9 1 11 13 0 16 15 13 10 9 2
24 1 10 11 11 11 11 10 9 0 13 11 11 2 13 1 11 7 9 1 11 7 11 11 2
29 13 3 16 15 13 9 1 10 0 9 13 1 10 9 0 2 16 10 9 1 9 13 3 9 7 10 9 0 2
39 10 9 8 7 2 9 0 2 2 13 9 1 10 9 13 1 9 1 10 9 1 10 12 3 10 11 11 1 11 13 10 9 1 10 9 1 9 0 2
12 4 13 1 12 2 1 9 1 10 9 11 2
12 10 9 13 9 7 13 10 9 1 9 0 2
12 10 9 13 13 1 10 0 9 1 10 9 2
29 10 9 4 13 1 11 2 11 2 16 13 2 3 10 9 2 2 13 16 10 9 13 3 10 9 3 0 2 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
19 1 10 0 9 2 15 13 10 9 0 7 15 13 10 12 9 1 12 2
9 2 4 10 9 13 1 10 9 2
8 2 4 13 1 10 11 11 2
34 10 12 13 5 12 1 10 9 1 10 9 8 1 12 8 8 8 2 10 12 0 9 1 9 2 7 13 1 10 9 9 8 8 2
28 15 13 0 2 13 10 10 9 1 9 2 3 1 5 12 2 2 7 3 15 15 13 10 9 1 5 12 2
12 3 4 13 10 9 9 0 1 9 1 9 2
25 3 0 1 12 2 13 9 1 9 16 13 1 11 2 4 13 1 10 9 1 11 1 12 9 2
14 4 13 1 15 1 10 9 3 0 1 10 9 0 2
10 10 9 15 5 13 12 5 3 3 2
15 1 12 13 12 9 2 7 12 13 0 1 9 1 9 2
12 4 13 1 10 15 2 7 3 4 4 13 2
65 10 9 13 15 16 13 9 1 10 9 1 11 11 2 9 1 9 2 1 9 1 10 15 15 13 10 9 9 1 9 1 9 2 13 1 10 9 16 10 0 9 13 1 10 9 1 9 2 1 10 9 15 13 10 9 1 11 2 10 11 0 1 10 9 2
13 10 9 0 13 0 1 10 9 0 1 10 9 2
50 10 9 11 15 13 1 10 9 0 0 2 1 9 3 1 10 9 1 10 11 7 15 13 10 9 2 16 11 2 9 2 13 0 1 10 9 0 2 1 10 9 1 10 9 0 1 9 1 9 2
36 10 9 0 13 1 9 1 10 11 1 10 11 1 11 1 11 1 11 15 13 10 9 1 16 1 12 4 13 7 13 1 10 3 0 11 2
24 16 13 9 2 4 13 1 9 1 10 11 11 11 1 11 2 3 13 10 9 1 10 9 2
22 10 11 11 1 11 13 10 9 0 13 1 11 2 11 2 11 1 10 11 11 11 2
18 15 13 1 10 11 1 11 1 12 7 10 11 11 1 11 1 12 2
15 10 9 0 15 13 0 1 0 9 1 9 1 10 9 2
17 13 10 9 0 1 10 9 1 10 9 1 10 9 1 9 0 2
16 13 1 10 9 1 9 2 8 8 2 1 10 0 9 12 2
32 11 3 13 1 10 9 2 11 2 1 11 11 11 11 11 2 7 13 10 0 9 1 10 9 0 1 12 11 11 11 15 2
31 3 13 10 9 1 10 9 3 4 7 13 10 9 16 15 13 1 10 10 9 1 10 9 2 8 2 9 7 8 2 2
30 10 9 1 11 2 11 11 11 15 13 1 10 9 1 10 9 1 11 2 7 10 9 13 1 0 10 9 1 11 2
46 10 9 13 1 10 9 0 1 10 9 13 8 16 13 1 10 9 0 8 2 8 2 16 13 3 2 10 11 2 2 13 9 1 10 9 0 1 9 0 1 10 15 15 13 11 2
24 10 9 13 10 9 1 12 9 7 12 9 2 7 10 9 13 15 1 12 9 7 12 9 2
12 13 1 11 7 13 1 10 11 1 10 11 2
13 11 13 13 10 9 7 13 10 9 1 10 9 2
18 15 15 13 10 9 1 11 1 10 11 11 10 12 1 11 1 12 2
33 13 10 9 0 16 13 9 0 1 10 9 0 2 0 2 1 16 10 9 15 4 1 13 7 13 1 10 9 16 13 1 9 2
27 1 10 11 11 2 13 10 0 0 9 2 9 7 9 16 13 3 1 10 9 7 1 10 9 1 11 2
23 13 9 1 10 9 7 10 9 2 3 16 13 10 0 9 16 15 4 13 1 10 9 2
30 10 9 3 0 13 2 1 9 0 2 13 1 11 11 2 1 12 8 2 13 15 3 1 10 9 0 1 12 8 2
20 1 11 2 11 13 10 9 9 1 12 2 16 13 1 9 2 11 11 2 2
27 13 10 0 9 0 7 9 1 9 1 10 9 1 11 1 11 2 3 13 1 10 9 1 11 1 11 2
9 10 9 4 13 1 10 0 9 2
36 3 3 2 11 13 10 9 11 11 2 1 0 10 9 1 10 9 13 1 9 0 7 13 8 2 8 2 0 1 10 9 1 10 9 0 2
22 11 13 13 1 11 10 0 9 1 9 1 10 9 0 1 11 7 10 9 1 11 2
35 1 12 11 15 13 1 10 11 1 11 3 2 1 10 9 12 2 13 3 9 1 10 9 0 1 9 0 2 11 2 11 11 11 2 2
33 1 10 9 15 13 1 9 1 9 1 10 9 2 10 9 2 10 9 2 10 9 2 10 9 0 7 9 0 7 10 9 0 2
12 4 13 1 2 11 2 1 10 9 1 12 2
13 3 2 10 9 11 13 13 1 9 7 13 15 2
25 10 9 0 13 10 9 1 9 0 1 10 9 16 13 13 7 13 10 9 1 9 1 9 0 2
26 10 9 13 10 9 3 0 2 7 13 1 10 0 9 1 9 1 10 9 1 10 9 1 9 0 2
30 9 13 7 13 1 11 11 7 16 13 13 7 13 9 1 10 9 0 2 10 9 2 10 9 2 10 9 0 0 2
8 3 2 15 13 1 10 9 2
31 1 13 13 10 9 1 12 1 12 5 8 2 1 15 15 10 9 4 7 13 15 1 12 1 12 9 3 1 10 9 2
27 10 9 0 15 13 1 9 13 1 13 10 9 1 9 7 1 9 16 13 0 10 9 1 10 0 9 2
28 1 10 9 10 12 9 15 13 2 1 10 15 13 0 10 9 0 7 10 9 1 9 0 2 0 7 0 2
40 15 0 15 13 0 1 10 0 9 1 9 1 10 9 0 7 10 9 2 3 1 10 9 1 11 11 16 13 2 3 2 10 9 3 0 1 10 10 9 2
23 1 12 2 10 9 1 11 13 10 9 7 13 10 9 1 11 11 2 10 0 9 0 2
29 1 10 9 7 1 10 9 0 1 10 9 13 2 1 10 9 2 10 0 9 0 1 13 10 9 16 15 13 2
51 3 4 13 10 9 1 10 16 15 13 16 1 9 4 7 13 1 10 9 1 10 9 16 1 15 15 13 10 9 2 7 16 1 15 3 15 13 2 3 15 13 1 13 1 10 9 9 1 10 9 2
29 16 10 9 13 1 0 9 13 1 13 10 9 3 1 13 2 9 1 10 15 10 9 13 10 9 2 13 2 2
14 3 15 13 9 2 13 7 10 9 9 9 13 0 2
33 1 10 9 1 3 2 1 10 12 2 10 9 0 13 1 10 9 1 10 9 0 1 10 11 11 2 13 1 11 11 7 11 2
37 11 13 10 9 1 10 9 1 9 1 10 11 11 11 1 10 9 1 11 2 7 1 10 9 1 12 9 2 4 13 1 10 9 2 11 11 2
35 11 13 7 13 9 1 10 0 9 2 11 11 11 2 2 13 10 9 1 9 10 12 1 11 1 12 1 10 9 0 1 10 11 11 11
23 10 0 9 0 13 1 9 0 1 10 9 2 16 13 1 0 9 1 11 11 1 12 2
15 1 10 9 1 11 11 15 13 10 9 0 1 12 8 2
19 1 10 9 3 0 13 1 10 9 13 10 9 7 10 9 1 10 9 2
7 15 13 1 9 1 9 2
49 1 10 9 1 12 9 2 1 10 15 12 10 9 13 0 1 10 8 2 10 11 7 10 9 13 3 1 12 9 1 9 2 12 9 1 10 9 0 1 10 9 2 9 7 9 1 9 0 2
15 1 10 9 12 13 1 10 11 1 11 11 1 10 9 2
24 3 13 9 0 2 1 9 0 7 0 2 7 3 13 10 8 0 3 10 9 15 13 15 2
37 1 10 9 1 11 1 11 1 12 2 15 13 3 10 9 11 11 11 15 1 10 0 9 13 3 15 4 13 10 10 9 16 13 10 9 0 2
26 15 15 13 1 9 1 10 9 1 10 9 1 10 0 9 1 9 0 7 10 9 13 1 9 0 2
24 15 9 16 4 7 13 13 2 13 10 9 2 13 15 13 10 9 7 13 1 10 9 0 2
24 10 0 9 13 1 10 9 3 1 10 9 1 11 13 10 0 9 0 2 13 1 11 11 2
26 10 9 13 1 9 1 10 9 0 2 10 9 1 10 9 1 10 9 7 15 1 10 1 10 9 2
30 10 9 13 10 9 1 9 3 0 1 16 13 10 9 0 7 0 16 13 1 10 9 1 9 7 9 1 10 9 2
12 11 11 13 10 9 1 9 1 10 9 11 2
34 11 13 10 9 1 3 1 12 9 1 9 3 0 16 15 13 1 10 9 9 0 2 1 10 9 1 10 9 1 11 1 10 9 2
28 1 12 10 0 9 1 10 9 0 1 10 9 4 13 2 15 16 15 13 1 10 0 9 0 1 10 9 2
15 11 11 11 2 11 13 10 9 2 9 0 7 9 0 2
39 7 1 10 13 10 9 15 10 9 0 13 1 1 9 10 9 13 7 13 16 15 13 0 9 2 7 13 10 9 1 10 9 16 13 10 11 1 11 2
14 10 9 13 16 13 9 7 15 13 3 13 10 9 2
22 1 12 2 10 9 0 1 9 1 9 1 11 7 11 1 10 11 13 1 12 9 2
19 3 4 1 13 13 1 15 3 2 16 13 16 15 13 15 2 10 9 2
13 13 10 9 1 9 7 10 9 1 10 0 9 2
6 4 13 1 11 11 2
10 13 9 1 11 11 11 7 1 11 2
14 1 10 9 0 1 12 2 13 10 9 11 11 11 2
22 1 0 9 2 11 11 13 10 9 1 12 2 1 10 15 13 9 15 7 10 9 2
54 1 10 9 1 9 2 11 1 11 13 0 1 10 9 0 2 7 3 0 1 10 9 1 10 9 1 10 9 2 1 15 0 1 10 9 7 9 0 1 11 12 2 3 1 10 9 1 10 9 2 11 1 11 2
34 10 9 1 9 15 4 1 13 13 9 0 7 13 10 9 15 3 0 1 9 1 3 1 10 15 16 13 9 7 10 9 1 9 2
12 10 9 13 3 0 1 10 9 0 7 0 2
16 11 11 2 12 2 13 11 11 2 9 1 9 2 12 2 2
17 3 2 13 1 10 9 11 7 11 2 1 10 9 1 11 11 2
26 10 9 4 13 1 9 10 0 9 16 10 11 11 3 15 13 7 13 9 1 10 2 0 9 2 2
29 10 9 1 12 9 15 13 0 16 11 13 10 0 7 0 9 1 10 9 1 13 9 1 9 0 1 10 9 2
53 10 9 0 13 10 9 0 1 10 9 0 1 10 9 2 1 9 1 13 10 9 0 2 0 7 0 2 16 13 9 0 1 9 7 9 1 9 2 1 9 0 2 13 9 0 1 15 13 1 10 9 0 2
35 11 2 11 11 2 2 11 2 12 1 11 1 12 2 11 1 11 2 3 1 11 2 12 1 11 1 12 2 13 10 9 7 9 0 2
32 1 10 9 15 13 3 16 13 9 1 9 1 10 9 7 16 4 13 1 9 1 9 1 9 2 9 1 9 7 10 9 2
16 15 15 13 10 9 1 10 9 7 10 9 0 1 10 11 2
16 0 9 1 9 0 2 1 15 1 11 16 13 3 9 0 2
15 15 1 15 13 1 10 9 1 10 12 9 1 10 9 2
21 11 13 9 1 9 0 2 11 2 2 10 9 1 0 9 7 9 7 10 9 2
16 2 0 9 1 10 9 12 1 9 1 9 0 9 7 0 2
24 3 1 15 15 13 16 16 13 10 9 15 4 13 3 9 2 7 1 10 9 13 15 9 2
36 1 10 9 15 4 13 2 2 4 4 13 1 10 9 1 9 1 10 9 2 10 9 0 1 10 9 2 7 10 9 0 1 10 9 2 2
10 13 13 9 1 10 11 11 1 11 2
21 3 2 10 9 0 3 13 0 1 9 1 10 9 1 11 7 0 1 9 0 2
31 1 11 13 10 0 9 3 0 1 9 0 3 1 10 11 2 9 16 13 1 10 11 2 11 7 3 10 11 7 11 2
14 10 9 13 10 9 1 9 1 1 12 7 12 9 2
13 1 10 9 1 10 9 11 9 3 2 12 5 2
28 16 15 13 16 10 9 13 10 9 9 7 10 9 9 2 10 12 9 3 4 13 15 10 15 1 10 15 2
8 10 9 1 10 9 13 11 2
36 10 9 0 2 1 10 9 2 0 2 1 10 9 7 1 9 1 10 9 15 4 13 1 10 9 0 2 1 9 7 0 1 10 12 9 2
40 10 10 9 1 9 1 9 0 0 2 0 7 0 3 13 3 7 2 9 0 2 15 10 9 2 7 10 9 1 10 9 1 10 9 0 2 13 1 0 2
19 13 10 9 0 1 13 15 2 3 2 7 1 10 9 9 2 9 0 2
21 13 9 1 10 11 11 11 12 9 0 1 12 7 12 7 9 1 12 7 12 2
35 15 13 1 10 11 0 2 10 9 1 11 2 10 9 1 10 11 1 11 2 10 11 2 10 11 11 7 9 1 10 9 0 1 11 2
7 10 9 3 15 13 2 2
13 11 11 13 1 9 1 10 11 11 11 1 12 2
7 9 0 7 0 1 11 2
16 10 9 0 1 10 15 15 13 2 7 4 13 1 13 15 2
28 1 9 0 13 1 10 9 11 11 11 11 11 2 13 1 10 9 1 11 11 7 3 13 1 11 1 11 2
12 1 15 15 13 2 11 2 2 13 1 11 2
19 15 15 13 3 1 10 9 2 7 3 13 0 9 1 10 9 7 9 2
62 10 9 11 2 11 13 9 0 1 10 15 13 9 0 0 7 0 1 9 1 10 9 0 1 10 9 2 16 4 13 10 0 9 9 2 9 7 9 2 9 3 7 13 1 10 9 11 2 11 7 10 9 11 2 11 2 1 3 13 12 9 2
14 11 13 10 9 7 9 1 10 9 1 11 1 11 2
24 13 10 9 16 13 10 9 7 10 13 3 0 2 10 9 13 3 0 7 10 9 13 0 2
8 10 9 13 1 15 3 0 2
29 15 4 13 3 1 10 9 2 7 3 13 1 10 9 7 15 13 2 1 9 1 10 9 2 1 10 9 0 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
49 1 10 9 1 10 9 2 11 11 15 13 3 0 1 13 1 10 9 1 10 0 9 11 1 9 11 11 11 2 16 13 10 9 1 10 9 1 9 0 16 10 9 4 13 1 10 0 9 2
31 1 10 9 15 10 9 11 13 7 13 2 10 9 13 10 9 1 10 9 1 10 15 13 7 1 10 15 13 10 9 2
35 10 9 13 0 7 13 12 9 0 1 10 9 2 1 10 15 3 3 13 12 2 7 10 0 9 1 12 9 16 13 1 10 0 9 2
67 10 9 0 1 10 9 13 13 2 3 2 1 10 10 9 1 9 16 13 10 0 9 2 10 9 1 10 11 2 16 4 13 1 10 0 9 2 3 0 1 10 9 2 10 9 13 1 10 9 2 10 3 0 1 11 2 10 11 7 15 1 10 3 0 1 11 2
38 3 2 13 0 9 1 16 13 10 0 9 1 10 9 1 10 9 0 1 9 1 10 9 11 11 2 16 13 1 10 9 10 9 1 12 12 9 2
11 10 11 11 1 11 15 13 1 12 9 2
32 10 9 13 10 9 1 10 9 13 1 10 9 1 12 0 9 2 10 11 7 10 11 2 1 9 1 10 9 1 10 9 2
71 3 2 15 15 13 13 2 9 3 1 10 9 2 1 0 9 0 9 1 10 9 2 7 1 10 9 2 1 10 9 1 13 10 9 16 13 10 9 0 7 9 1 9 0 2 3 1 10 9 0 1 1 10 0 9 1 9 0 2 7 10 9 16 4 13 1 10 9 3 0 2
24 10 9 13 15 1 10 9 0 1 10 9 7 13 10 9 9 0 1 9 0 1 10 11 2
38 10 9 4 13 10 9 1 10 9 1 10 9 1 10 11 11 1 10 11 1 11 2 0 11 1 11 2 13 1 10 9 1 10 11 1 10 11 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
20 10 9 1 9 7 11 4 13 15 1 10 9 1 10 9 0 7 10 9 2
17 4 1 13 7 1 0 1 13 9 1 10 9 1 11 7 11 2
10 4 1 13 1 11 7 3 13 0 2
23 10 0 9 1 9 1 10 9 2 13 0 9 16 13 10 9 1 0 9 1 10 9 2
24 10 9 0 4 13 1 10 11 11 2 3 1 10 0 11 2 1 10 9 12 7 3 3 2
35 11 13 13 15 1 10 9 2 7 10 0 9 0 9 1 10 9 1 10 9 2 10 9 7 10 9 2 15 13 1 13 10 0 9 2
15 1 10 0 13 12 0 9 7 1 10 9 13 12 9 2
30 3 16 10 9 13 10 9 7 10 9 0 13 10 9 2 10 9 3 13 1 10 9 0 0 16 13 10 9 2 2
32 10 9 13 10 9 1 9 1 10 9 1 10 9 13 2 9 1 10 9 0 2 2 3 13 1 2 8 2 9 0 2 2
36 1 10 9 0 1 10 11 11 11 7 1 10 9 13 2 9 0 2 2 10 9 4 4 13 1 9 7 10 9 9 15 13 3 1 15 2
17 10 9 15 13 7 13 2 3 15 13 3 9 2 3 1 12 2
21 11 11 2 13 1 10 9 0 1 11 2 10 11 2 2 13 10 9 0 0 2
29 15 13 10 9 1 12 9 13 1 9 2 3 0 10 9 2 7 10 9 1 12 9 1 4 13 3 10 9 2
43 13 1 10 9 15 1 10 9 1 10 9 0 2 10 9 0 13 13 10 9 16 13 1 11 1 10 9 9 1 11 7 11 7 10 3 9 1 10 9 9 1 11 2
20 10 9 13 9 1 10 9 1 9 16 13 16 3 13 15 13 1 10 9 2
25 16 15 13 1 10 9 1 13 15 10 9 1 16 15 13 2 4 13 1 10 9 1 10 9 2
39 11 13 1 11 7 13 10 9 1 15 1 10 9 3 15 13 10 0 9 2 1 15 15 15 4 13 1 10 9 1 10 8 2 9 1 10 0 9 2
52 16 13 1 9 1 4 13 0 1 10 9 2 1 9 1 10 9 16 13 3 1 10 9 1 11 11 2 15 3 13 9 1 10 9 1 11 2 15 15 13 1 10 9 1 16 15 13 1 10 11 11 2
13 4 13 1 10 10 9 7 13 0 1 10 9 2
15 3 13 9 0 13 1 10 11 11 1 11 2 11 2 2
21 9 11 7 11 2 10 9 1 10 9 2 13 10 9 1 9 13 1 10 9 12
14 13 1 9 0 7 13 1 10 9 1 9 1 9 2
41 1 9 1 10 9 2 13 1 11 11 2 13 1 11 2 2 15 15 13 1 10 11 7 15 13 1 16 15 13 1 13 7 13 10 9 2 7 3 13 3 2
11 10 9 13 10 9 1 9 1 11 11 2
13 1 12 2 10 12 9 4 1 13 10 0 9 2
26 1 13 1 12 2 15 13 1 0 9 1 9 0 1 10 11 11 11 1 11 7 11 1 11 2 11
43 10 0 9 11 11 11 4 13 10 9 0 1 16 10 9 8 1 0 9 2 7 10 9 2 3 3 13 1 9 2 7 15 3 4 13 10 9 7 1 13 10 11 2
19 13 11 11 2 13 10 9 1 13 15 3 2 7 10 9 15 13 13 2
32 11 11 13 10 9 0 1 10 11 1 11 1 12 7 13 9 1 12 1 9 1 10 11 11 1 11 2 3 11 1 11 2
16 13 10 9 1 9 3 2 3 0 2 10 12 7 12 2 2
27 1 9 7 0 2 15 13 9 1 9 2 8 2 1 10 9 0 1 10 9 7 9 0 1 10 9 2
5 3 13 10 9 2
13 15 1 0 9 4 13 9 0 2 1 10 9 2
38 10 12 1 11 1 12 2 1 10 9 0 1 10 11 1 10 9 2 11 11 4 13 9 1 10 11 1 10 9 11 1 9 0 1 11 1 12 2
17 1 10 9 12 10 12 5 5 15 13 1 10 9 0 1 9 2
30 16 1 10 9 13 10 9 1 9 9 0 1 0 2 1 10 9 1 10 9 11 2 11 15 13 1 10 9 0 2
16 15 13 10 9 1 10 12 9 0 1 10 15 13 10 9 2
15 13 1 10 9 1 10 9 1 10 9 0 1 10 9 2
23 1 12 15 13 1 10 9 16 15 13 2 7 1 10 15 13 1 15 3 1 10 9 2
36 13 1 12 9 9 1 10 11 1 11 2 13 10 9 1 9 1 9 7 4 13 1 10 9 1 10 11 1 10 9 0 1 11 1 12 2
55 3 1 10 9 9 0 2 10 9 11 3 13 10 9 3 15 13 10 9 0 1 10 9 7 10 9 1 9 1 10 9 0 3 1 10 11 2 10 9 0 7 0 13 10 9 16 1 15 9 13 3 1 10 9 2
13 11 13 10 9 0 1 10 9 1 11 7 11 2
17 1 9 0 2 10 9 0 1 10 9 13 1 12 9 7 3 2
27 13 1 10 9 16 11 11 15 13 1 10 0 9 1 10 0 9 2 1 9 0 7 9 0 1 13 2
43 10 9 0 11 15 4 13 1 10 9 11 1 11 11 7 11 2 10 9 16 13 13 0 9 1 10 0 7 0 9 2 7 13 3 1 10 9 2 3 1 10 9 2
13 10 9 15 13 1 9 7 9 1 10 11 11 2
33 11 13 3 1 10 9 1 10 9 2 0 12 9 1 11 1 12 7 12 2 7 9 0 1 11 7 13 1 10 11 1 11 2
16 4 13 2 3 2 1 15 2 11 2 11 11 7 11 11 2
26 3 15 15 13 11 11 11 2 11 2 1 10 9 1 10 15 10 9 13 10 9 3 1 4 13 2
15 10 9 7 10 9 0 3 13 10 0 9 1 10 9 2
21 13 3 0 16 10 9 15 13 1 10 9 1 11 13 1 10 9 1 10 9 2
24 10 9 13 1 10 9 1 11 11 1 10 11 1 11 2 3 11 13 13 1 10 9 11 12
27 10 9 13 16 10 9 11 15 13 1 10 9 1 11 2 11 11 2 2 1 10 15 3 13 10 9 2
20 11 11 2 12 1 11 1 12 2 11 2 11 2 13 10 9 7 9 0 2
19 13 1 15 16 15 13 13 10 9 1 10 9 7 9 13 1 10 9 2
27 10 9 13 16 10 9 1 10 11 7 10 11 4 13 15 1 10 9 1 13 1 10 9 1 10 9 2
36 1 10 9 1 9 1 10 9 11 1 10 9 1 10 9 2 13 1 9 1 10 9 11 11 10 9 1 9 1 10 9 0 11 2 11 2
10 15 13 1 10 9 13 9 9 0 2
24 13 14 9 1 10 11 0 0 1 9 2 9 1 10 11 1 11 7 11 11 2 8 2 2
9 10 9 0 0 13 10 9 0 2
25 2 10 9 4 1 4 13 1 10 9 1 12 7 12 9 2 2 13 2 11 2 1 9 0 2
10 11 15 13 7 13 16 15 15 13 2
7 15 13 1 10 11 0 2
38 11 13 10 9 7 9 0 2 1 10 9 1 11 2 11 2 9 1 11 2 1 10 9 1 11 2 9 2 11 7 9 1 11 2 1 2 11 2
28 2 11 11 11 11 11 2 13 10 9 1 9 9 2 9 7 9 10 9 13 1 10 12 9 7 12 9 2
32 3 2 1 12 9 1 9 2 13 12 9 1 11 2 1 3 13 1 9 1 12 2 13 1 10 9 1 10 9 7 9 2
29 1 10 9 1 9 11 11 13 1 10 9 1 9 11 11 2 10 9 3 0 1 10 9 11 4 13 1 15 2
19 15 13 16 10 9 8 13 1 10 9 1 10 9 1 13 15 10 9 2
24 1 10 9 1 12 2 11 13 1 10 0 9 0 1 16 13 1 9 0 1 10 9 0 2
12 10 9 13 0 7 0 13 9 1 8 7 8
17 3 1 10 0 9 2 10 9 15 13 3 0 7 13 1 9 2
26 1 10 9 1 9 13 1 10 9 0 15 4 13 9 1 10 10 9 2 1 10 9 7 9 0 2
40 11 11 2 11 2 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 13 9 1 11 1 10 12 1 11 1 12 1 10 12 1 11 1 12 2
23 10 9 0 15 13 1 9 2 13 1 15 10 9 1 10 9 1 9 1 10 9 0 2
37 10 0 9 2 13 10 12 1 11 1 12 2 1 10 9 1 10 9 2 1 10 9 1 11 16 10 11 2 12 3 13 3 1 9 1 9 2
37 1 9 1 10 9 2 11 4 13 1 10 9 1 13 1 10 9 2 7 10 9 13 10 9 7 10 9 15 13 16 3 13 9 1 10 9 2
25 10 9 13 10 9 1 13 10 9 0 7 13 15 16 13 10 9 1 9 0 1 10 9 0 2
26 10 9 9 1 11 10 11 15 13 0 1 13 10 9 1 10 9 1 9 0 1 9 1 10 9 2
11 1 10 9 13 10 1 10 9 1 9 2
11 10 9 1 9 13 10 11 11 11 11 2
14 10 0 9 2 12 5 2 13 9 1 10 11 11 2
29 14 3 13 16 10 9 16 15 13 10 9 1 9 13 0 1 3 1 10 9 2 1 10 9 7 1 10 9 2
36 13 9 1 10 9 0 11 11 11 11 11 11 2 3 1 8 2 9 1 10 11 11 7 2 3 2 9 1 10 11 11 11 2 11 2 2
42 1 10 15 2 4 13 16 10 9 1 9 2 16 4 1 4 13 10 9 10 9 1 9 13 0 2 4 1 13 0 1 10 9 0 1 10 9 16 13 10 9 2
57 16 13 3 2 10 11 2 1 10 11 11 2 10 9 1 12 9 13 15 1 10 9 16 3 13 1 10 9 2 1 15 15 13 10 11 1 11 7 10 11 2 10 9 13 10 9 16 13 10 9 10 0 9 2 10 12 2
37 15 16 13 1 10 9 0 9 3 13 10 13 9 1 10 9 1 10 9 2 7 10 9 1 13 1 10 9 1 9 1 10 9 9 1 9 2
10 10 9 1 9 15 13 1 12 9 2
43 10 9 0 2 13 1 10 9 1 11 2 11 1 10 11 7 11 3 2 10 12 0 9 15 13 1 10 11 11 11 7 10 0 9 13 1 10 11 11 11 11 11 2
21 11 13 10 9 1 11 2 1 10 9 1 11 2 9 0 1 11 2 10 11 2
55 1 11 1 12 2 13 16 10 9 13 2 2 2 2 3 3 0 1 10 9 1 9 0 2 7 3 3 0 2 2 13 10 9 1 10 9 0 1 10 9 16 13 1 0 9 0 1 10 9 1 11 7 10 9 2
13 11 11 1 11 15 13 1 10 9 12 1 12 2
14 10 9 11 13 10 9 10 9 13 3 0 7 0 2
18 15 13 2 1 9 0 2 10 9 1 10 11 2 10 12 1 11 2
23 10 9 13 2 3 2 10 9 0 1 10 3 0 1 10 9 7 10 9 1 10 11 2
29 15 13 3 7 3 1 10 9 1 9 7 4 13 15 1 10 9 1 10 10 9 0 1 10 16 13 10 9 2
36 1 12 2 1 12 9 1 9 2 10 9 11 13 16 10 9 0 3 13 9 7 16 13 10 9 1 13 10 9 1 11 11 1 10 11 2
22 10 9 13 10 9 1 3 12 9 7 10 9 1 10 9 4 4 13 1 9 0 2
32 13 10 0 9 1 13 15 1 10 9 1 10 11 11 2 7 3 15 13 1 10 9 0 1 9 2 16 13 15 3 0 2
42 1 10 0 9 1 10 9 13 10 9 1 10 9 7 9 10 2 9 0 2 2 7 10 9 1 10 9 7 9 1 10 9 11 7 1 10 9 7 9 1 11 2
22 3 1 13 15 1 10 10 9 2 3 11 11 13 15 1 15 7 3 15 13 15 2
37 3 1 10 9 1 10 9 10 11 2 11 12 13 13 15 10 0 9 1 11 11 2 3 1 10 0 9 1 10 9 1 10 11 1 10 11 2
22 3 4 1 13 10 0 9 1 9 2 15 16 15 13 13 1 9 1 9 1 9 2
31 10 9 2 13 1 9 11 2 4 13 1 10 9 1 0 9 1 9 1 11 2 7 4 13 1 0 9 1 9 0 2
27 3 13 5 2 0 9 1 11 2 11 7 15 2 2 9 0 1 9 1 9 7 9 2 7 11 8 2
21 10 9 13 16 10 9 1 11 4 13 3 1 10 9 13 1 11 1 10 9 2
12 10 9 7 10 9 13 1 15 9 1 11 2
60 15 2 13 1 10 0 9 1 13 1 10 9 7 1 10 9 1 2 9 2 2 10 9 2 9 13 1 10 9 1 11 2 11 11 2 13 3 3 0 13 10 0 9 7 3 0 10 9 1 10 9 1 10 9 7 9 1 10 9 2
20 10 9 2 1 10 0 9 2 3 13 9 2 13 1 10 9 1 10 9 2
57 13 1 16 10 9 1 9 0 13 2 8 2 7 2 8 2 1 10 9 1 10 9 1 9 0 2 15 13 12 8 12 8 2 8 2 8 2 8 2 8 2 8 2 8 2 7 8 8 8 8 2 8 2 1 10 11 2
23 16 10 9 13 9 1 9 2 1 9 2 10 9 4 13 10 9 0 13 10 9 0 2
21 10 12 1 11 1 12 4 13 0 9 1 10 11 2 1 9 1 11 1 11 2
4 7 15 13 2
30 10 0 9 7 9 0 0 7 0 1 11 13 1 11 1 12 2 13 1 10 9 0 11 11 1 9 1 10 11 2
28 15 13 0 2 7 13 10 9 3 0 1 9 0 1 9 1 9 1 12 9 1 11 1 16 15 13 9 2
18 10 11 13 10 0 9 0 13 1 11 11 2 1 10 9 1 12 2
22 1 15 9 10 8 13 10 9 15 0 2 1 9 1 10 9 16 13 1 9 0 2
31 1 12 2 4 13 1 8 9 1 13 10 9 1 9 1 9 1 10 11 11 1 11 2 1 9 1 10 11 1 11 2
31 10 9 0 1 10 9 16 3 13 13 0 1 10 9 1 9 2 13 1 13 10 9 0 1 15 0 2 0 7 0 2
10 10 9 13 4 1 13 1 10 9 2
7 3 13 1 10 9 0 2
10 10 9 13 3 0 16 13 1 9 2
41 1 10 9 3 1 10 9 2 11 13 1 10 9 15 13 13 0 1 10 9 2 7 3 4 13 1 10 11 11 2 3 7 13 1 9 1 10 9 1 9 2
37 10 9 3 0 1 10 9 13 0 1 1 13 10 9 10 9 3 2 1 9 10 9 13 1 10 9 0 16 9 7 9 15 15 13 1 3 2
90 1 10 9 2 1 10 9 0 2 10 11 1 11 2 9 1 10 9 0 2 13 1 10 9 11 12 16 13 1 13 10 9 2 1 15 15 15 15 13 2 13 16 10 9 1 10 9 13 1 10 9 0 7 0 2 16 13 10 9 7 9 1 11 2 10 9 1 10 9 0 1 10 11 7 10 9 1 10 10 9 0 1 10 9 1 9 1 10 11 2
8 11 15 13 13 1 10 9 2
23 10 9 3 13 10 9 7 13 9 1 10 10 9 1 10 9 1 10 9 1 10 9 2
21 8 2 7 13 1 9 16 10 9 2 3 1 11 15 13 1 10 9 1 11 2
11 11 13 10 9 1 13 10 9 1 11 2
20 1 15 2 11 15 13 13 1 10 9 7 3 1 10 11 2 10 9 0 2
16 1 15 13 0 10 9 1 10 9 2 7 15 13 3 0 2
39 1 10 9 2 15 13 1 10 9 0 3 0 16 13 1 10 9 0 0 1 12 2 13 1 11 11 2 16 4 13 1 10 9 1 12 9 1 12 2
20 10 12 9 15 13 1 10 9 1 13 15 2 9 1 10 11 1 9 2 2
18 13 1 15 1 12 9 2 16 13 13 15 3 1 9 1 10 9 2
24 1 10 11 11 2 10 11 0 13 1 10 9 1 9 2 9 2 7 9 0 1 10 9 2
86 10 9 1 10 9 1 11 2 11 7 11 2 13 1 10 9 0 1 10 9 0 2 7 13 1 11 2 15 13 1 10 0 9 1 13 10 9 7 13 10 0 9 2 16 15 13 1 3 1 12 9 1 9 2 13 10 9 7 9 7 10 9 1 9 1 9 16 13 10 9 1 10 11 2 7 15 3 15 13 1 0 9 1 10 9 2
23 11 11 11 2 13 12 1 11 1 12 1 11 2 11 2 2 13 10 9 1 9 0 2
24 13 10 0 9 1 11 2 10 9 1 10 9 4 13 15 1 10 9 1 10 11 7 9 2
33 1 13 10 11 11 4 13 1 10 9 1 11 2 3 13 1 10 11 11 7 11 2 10 9 13 1 10 11 1 11 1 11 2
46 1 10 9 12 10 9 2 1 10 9 0 2 15 13 1 15 1 11 7 0 9 1 10 9 13 15 1 10 9 1 11 12 2 1 16 4 13 1 10 9 1 10 11 1 11 2
26 10 9 4 4 13 12 9 13 15 3 0 10 9 1 12 9 13 1 10 9 11 11 11 1 12 2
15 13 10 9 1 10 15 13 1 11 1 9 1 10 9 2
21 10 9 0 11 11 13 10 9 13 2 11 11 1 10 11 2 1 10 0 9 2
40 15 15 13 1 10 9 2 10 9 1 10 12 5 9 4 13 1 10 9 0 0 2 16 1 9 4 13 15 0 16 10 9 0 1 11 13 1 13 15 2
39 1 15 16 1 10 9 15 13 2 7 1 13 3 0 2 10 9 3 13 16 1 10 9 7 15 15 13 9 1 16 10 9 13 7 4 13 10 9 2
38 11 11 13 1 0 9 1 12 1 10 0 9 1 11 11 7 10 9 1 9 1 11 11 2 1 9 10 9 1 11 13 16 15 13 1 10 9 2
56 1 9 1 12 7 9 1 12 2 15 13 10 9 1 9 1 10 9 1 10 9 1 10 9 11 11 7 11 11 2 1 10 9 11 1 11 11 7 11 11 2 3 13 11 11 2 11 11 2 11 11 7 10 0 11 2
26 1 13 10 9 4 13 10 0 9 1 0 9 0 2 0 7 0 1 10 11 1 11 7 11 11 2
15 10 9 13 15 0 2 7 13 9 10 9 1 10 9 2
18 7 11 15 13 1 10 9 7 13 13 15 1 9 1 10 10 11 2
21 10 11 11 15 13 10 12 1 11 1 10 12 1 10 9 1 10 9 1 11 2
12 3 2 11 13 0 16 11 15 13 1 11 2
13 10 11 1 11 13 1 12 9 13 1 9 0 2
29 3 1 10 9 11 11 13 3 10 9 1 10 9 1 11 11 7 13 3 10 9 0 1 13 9 1 10 9 2
32 4 13 1 10 9 1 9 1 10 9 1 10 11 2 1 9 1 11 11 2 11 11 11 2 11 1 11 7 11 10 11 2
21 1 10 9 10 9 13 1 9 10 9 0 1 13 1 9 3 0 1 10 9 2
25 11 15 13 9 1 16 15 3 13 10 9 1 11 2 7 16 10 9 15 4 13 1 10 9 2
25 1 10 11 2 1 10 11 1 11 2 13 10 9 0 1 10 11 1 10 11 1 10 9 0 2
10 1 10 9 12 2 12 13 10 9 2
40 9 1 15 2 1 9 1 15 1 11 11 2 0 1 9 0 2 15 4 13 1 9 10 0 9 1 9 2 9 7 9 1 10 10 9 0 1 10 9 2
18 10 9 0 1 10 9 0 2 7 10 9 1 10 9 0 13 0 2
50 1 9 2 16 3 10 9 13 10 9 1 10 11 11 1 10 11 1 11 1 10 12 7 12 1 11 1 12 1 10 9 1 10 11 1 11 11 1 11 15 13 16 10 9 1 11 13 3 0 2
36 11 11 11 2 1 10 9 1 10 9 11 11 7 11 1 10 11 7 11 11 2 11 11 2 13 10 9 15 4 13 1 12 1 9 0 2
19 10 9 4 13 1 12 7 8 15 4 13 1 3 3 1 12 12 9 2
32 1 9 1 10 0 9 11 13 10 9 1 9 0 1 11 2 13 1 12 9 0 1 9 1 10 12 0 7 13 10 9 2
35 10 9 13 13 10 9 16 13 1 10 9 1 10 9 3 7 10 9 0 15 13 1 11 10 9 1 9 1 10 9 7 10 9 0 2
6 13 10 9 1 11 2
20 15 16 10 9 13 11 11 4 13 1 13 1 10 9 2 1 10 9 0 2
24 11 2 10 9 2 13 10 0 9 2 13 10 9 16 13 16 13 10 9 0 1 0 9 2
32 4 7 13 10 9 0 1 10 11 7 15 13 1 10 9 1 10 9 2 1 15 13 1 10 9 1 8 9 2 2 13 2
11 10 9 4 13 10 12 9 1 9 0 2
41 1 9 2 15 4 13 1 10 9 1 10 12 1 11 1 12 1 10 9 11 2 11 2 13 1 9 0 1 10 9 11 11 2 13 10 9 1 10 9 0 2
17 10 9 0 13 11 11 2 15 15 13 1 10 0 9 1 9 2
20 1 10 9 10 9 4 13 3 0 7 3 0 2 13 1 10 9 10 9 2
25 1 10 0 9 1 9 13 10 9 1 11 1 10 11 11 1 11 11 2 15 4 13 1 11 2
32 10 9 0 1 10 9 7 10 0 9 13 1 10 9 10 9 3 0 2 15 4 13 3 3 1 10 9 2 9 9 2 2
35 4 3 13 1 10 9 15 4 13 1 9 1 10 0 9 1 10 9 1 10 9 7 15 4 4 13 1 10 9 2 1 10 9 0 2
34 13 10 9 0 1 1 9 0 7 15 1 10 9 1 10 11 1 9 2 7 1 10 9 11 11 13 1 11 1 10 11 1 11 2
27 10 0 9 1 10 9 13 1 10 9 2 7 1 10 9 1 9 13 10 9 1 10 9 1 10 9 2
23 11 2 3 1 11 11 2 11 11 7 11 11 13 15 1 10 12 9 0 1 10 9 2
38 10 9 9 1 10 9 15 13 1 3 1 10 12 5 8 7 1 9 1 9 13 0 15 15 13 9 0 3 1 12 5 8 1 12 2 12 5 8
14 10 9 13 3 0 1 10 9 0 1 10 9 11 2
31 13 10 9 0 16 15 13 1 9 15 0 1 10 9 0 1 10 9 1 11 1 9 1 9 16 13 12 1 10 9 2
10 3 11 11 4 13 1 11 1 12 2
6 13 1 11 1 12 2
27 2 13 0 15 9 1 9 7 1 9 0 2 3 7 1 9 0 1 10 9 1 10 11 2 2 13 2
13 10 9 1 9 13 1 12 8 2 2 9 8 2
22 1 10 9 12 4 13 1 10 9 0 11 2 1 9 0 2 1 9 1 10 9 2
27 15 1 10 9 0 1 10 9 13 15 13 0 13 10 9 1 10 9 2 1 10 13 10 9 1 15 2
19 11 11 13 10 9 1 9 16 15 13 1 11 2 1 10 9 1 11 2
15 1 12 13 10 0 9 1 3 1 12 9 11 2 11 2
17 1 9 2 13 3 10 9 0 15 16 13 10 9 1 10 9 2
12 13 10 12 1 11 1 12 1 11 2 11 2
30 11 2 9 1 11 11 13 1 10 9 1 10 9 1 11 2 11 13 1 11 1 12 7 13 1 11 1 12 11 2
5 3 13 1 9 2
35 15 1 10 9 3 0 13 1 10 9 1 12 2 3 1 10 9 0 2 16 3 13 0 1 10 9 2 1 9 1 16 15 4 13 2
33 13 3 3 10 9 0 1 13 10 9 1 9 16 3 13 10 9 0 7 1 13 10 9 1 0 9 1 10 9 1 10 9 2
21 10 9 1 9 0 7 0 16 13 10 9 1 0 9 7 9 1 10 0 9 2
21 10 9 11 13 0 1 9 1 11 16 13 16 3 13 15 1 10 9 1 11 2
9 15 13 1 11 2 11 11 2 2
32 10 9 13 1 12 1 10 9 1 11 2 16 13 1 10 9 10 9 11 12 1 10 9 0 1 10 9 11 12 1 11 2
18 11 11 11 11 2 8 11 1 10 11 2 11 2 11 2 12 2 2
31 4 13 2 2 10 9 1 10 9 12 3 13 1 10 9 0 2 7 1 10 9 13 10 9 1 9 1 12 9 0 2
19 1 12 4 13 9 0 1 10 9 2 3 1 9 0 7 3 1 9 2
55 13 1 10 9 1 10 9 1 11 7 11 2 1 10 9 1 10 9 1 11 2 10 11 7 11 2 1 10 15 1 10 9 1 11 11 1 11 7 11 7 1 10 9 1 10 9 1 9 1 11 7 9 1 11 2
12 13 10 9 1 10 9 2 9 7 10 9 2
17 13 10 0 9 9 2 13 9 13 15 9 7 3 4 13 9 2
22 1 11 2 10 9 1 9 7 10 9 2 0 2 1 10 9 13 9 1 10 9 2
41 1 10 9 0 2 1 10 9 13 1 10 9 1 10 9 1 11 7 11 2 10 9 3 0 13 10 9 7 13 3 0 10 9 2 1 15 15 13 10 9 2
19 11 13 1 12 9 1 10 12 15 4 13 15 7 13 9 1 10 12 2
23 10 0 9 1 10 9 15 13 1 10 9 12 2 13 15 1 13 1 10 9 3 0 2
26 10 9 4 13 9 0 1 9 1 10 9 1 10 9 0 7 13 1 10 9 12 1 10 11 12 2
15 13 12 9 10 11 11 1 10 11 1 12 7 1 12 2
31 10 11 2 9 0 2 13 10 9 7 9 16 15 13 1 10 9 1 10 9 1 9 2 0 1 9 2 9 7 9 2
23 13 3 3 13 13 10 9 7 13 15 1 0 9 1 15 16 3 15 13 2 13 9 2
18 10 9 3 4 13 1 10 9 2 10 9 1 9 7 10 9 0 2
29 10 3 9 1 10 9 0 0 1 10 9 2 11 11 2 13 1 12 10 9 13 2 11 1 9 1 9 2 2
18 10 9 13 0 3 16 13 10 0 9 1 9 0 1 10 9 0 2
69 10 9 1 10 9 1 9 13 0 9 1 10 9 1 9 13 1 11 2 3 16 1 10 9 1 9 10 9 13 13 0 9 1 9 1 9 1 9 13 1 9 1 9 1 9 1 9 2 3 1 10 0 9 0 1 9 3 15 13 0 2 7 0 2 9 1 10 9 2
51 3 3 10 9 0 13 10 9 0 2 1 0 7 0 9 1 10 9 0 7 1 10 9 0 2 13 1 9 1 13 1 10 9 12 2 9 0 2 9 1 11 2 11 1 11 2 11 1 11 2 2
15 0 1 12 11 1 11 2 13 0 9 2 9 7 0 2
12 11 11 13 10 9 1 9 1 10 9 11 2
17 3 13 16 1 11 11 3 13 10 9 1 10 9 2 11 2 2
13 11 11 13 10 9 1 9 0 1 10 9 11 2
28 11 2 9 2 7 10 9 1 9 1 9 7 9 0 13 0 9 7 9 7 10 9 1 9 7 9 11 2
20 13 10 9 0 1 10 9 2 7 4 13 1 13 10 9 0 1 9 0 2
16 10 9 13 10 9 1 9 7 15 13 13 1 10 9 0 2
45 10 9 13 13 11 11 2 0 9 1 10 9 2 1 10 15 4 13 10 9 13 1 11 11 1 10 9 13 13 1 9 16 1 9 13 1 10 9 1 10 9 1 10 9 2
29 1 9 13 10 9 16 13 16 11 13 1 9 1 10 9 11 11 2 10 15 13 1 10 9 12 1 10 12 2
35 13 1 11 2 1 11 11 7 11 2 1 10 9 13 9 7 9 1 10 9 1 7 10 9 15 13 0 7 4 13 7 13 1 9 2
16 15 13 1 10 0 9 1 10 9 1 10 9 11 7 11 2
15 10 9 15 13 10 12 1 11 1 12 1 10 9 0 2
22 3 13 1 10 9 0 2 1 10 15 15 15 4 13 10 9 3 0 1 10 9 2
32 13 10 0 1 10 9 16 2 9 1 11 2 10 0 9 2 13 1 10 9 1 9 2 1 10 11 11 7 10 11 11 2
37 10 9 1 10 11 13 3 1 10 11 1 11 7 1 10 9 1 11 2 7 13 13 10 9 7 3 0 9 1 10 9 0 13 1 10 9 2
14 10 9 1 11 11 13 10 9 13 1 11 1 11 2
25 11 11 11 13 9 1 10 9 1 10 9 1 10 9 1 11 2 1 10 11 1 10 11 11 2
21 4 13 0 9 3 0 7 0 7 3 15 13 1 11 3 1 9 7 1 9 2
30 10 9 1 10 15 13 11 16 13 10 9 1 11 13 2 10 9 1 10 9 0 11 7 10 9 1 11 1 11 2
18 4 1 13 9 0 2 13 1 9 13 1 10 9 1 10 9 0 2
12 13 1 10 9 1 11 1 11 1 10 9 2
14 11 11 13 10 9 1 9 1 10 9 1 10 9 2
56 11 13 15 16 15 13 1 9 1 11 8 11 11 11 2 10 9 0 1 10 15 10 9 13 10 9 16 13 10 9 1 9 1 10 9 7 13 1 9 1 10 9 0 13 9 2 10 9 15 13 7 13 1 10 9 2
12 13 10 9 1 13 1 15 10 9 3 0 2
7 10 9 13 10 9 0 2
11 9 7 9 13 1 10 9 2 3 0 2
35 13 13 3 2 7 10 9 3 13 10 9 0 1 12 2 9 3 0 13 10 9 15 13 10 9 1 9 1 10 9 0 1 10 9 2
56 15 13 10 9 1 10 2 0 9 2 1 10 9 1 9 9 1 10 9 1 10 9 2 9 16 15 13 1 10 9 0 1 10 9 0 1 10 9 2 10 9 1 12 9 13 1 10 9 1 10 9 2 1 10 9 2
63 10 9 13 1 9 0 2 1 11 1 11 2 1 10 9 13 1 10 9 7 10 9 1 13 13 10 9 1 10 9 1 10 9 0 1 10 9 2 16 13 10 9 0 7 0 9 2 3 7 3 10 9 7 9 1 10 9 7 1 10 9 0 2
24 3 1 10 9 1 9 2 1 11 13 10 9 11 11 2 10 9 11 7 10 9 10 11 2
49 10 9 3 2 10 9 11 2 9 0 1 10 11 2 13 10 9 7 13 16 15 13 1 10 0 9 15 10 9 1 10 9 13 1 2 10 9 0 2 15 4 13 1 13 1 10 9 2 2
26 13 1 10 9 1 10 9 2 1 10 9 1 10 11 11 7 10 11 1 10 11 11 1 10 9 2
40 15 3 1 11 2 1 12 2 13 9 1 10 9 0 2 7 10 9 11 15 13 7 15 13 1 9 1 10 9 0 2 1 13 1 10 9 1 10 11 2
12 10 0 9 13 1 10 12 1 11 1 12 2
7 13 1 9 0 1 11 2
28 1 3 1 12 9 2 10 12 1 11 2 15 13 1 10 0 9 1 10 9 2 3 15 13 1 12 9 2
46 10 0 9 11 2 11 13 10 9 16 13 1 10 9 1 10 11 1 9 1 10 12 0 9 0 1 11 2 11 11 2 11 11 2 7 11 11 11 11 2 11 11 11 11 2 2
26 3 1 12 2 11 11 11 13 1 0 9 1 10 9 2 11 10 11 2 1 11 11 8 11 11 2
24 4 13 9 1 10 9 0 1 10 11 1 11 7 4 13 10 9 1 10 9 1 10 9 2
14 1 10 12 9 15 13 13 1 11 7 13 10 9 2
17 10 9 1 10 9 4 13 11 15 1 10 9 3 0 1 11 2
43 10 9 1 9 4 13 1 1 10 9 1 10 9 1 10 9 2 10 15 3 15 13 3 2 13 1 10 9 1 9 1 9 2 9 1 9 2 9 7 9 1 9 2
63 1 10 12 9 2 10 9 1 11 11 13 0 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 9 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
39 1 10 9 1 10 11 1 11 1 11 11 1 11 1 10 12 2 13 12 9 7 12 9 1 10 9 2 7 10 9 1 12 5 1 12 9 1 12 2
34 10 9 13 3 1 10 0 9 0 1 9 7 10 9 0 13 2 16 13 9 7 9 13 10 9 1 9 1 9 0 7 15 0 2
9 15 13 3 1 10 10 9 0 2
15 1 10 9 2 11 4 1 13 11 2 10 9 3 0 2
56 11 4 13 10 12 1 11 1 12 9 1 10 9 1 12 9 16 13 1 11 2 11 7 11 2 11 11 11 2 13 1 11 2 2 11 2 11 2 2 11 11 11 2 11 2 2 11 2 11 2 7 11 2 11 2 2
29 1 10 9 2 4 7 13 16 11 13 16 11 13 1 11 1 12 2 3 13 1 10 9 3 0 2 11 11 2
44 10 9 13 15 1 10 9 1 10 9 0 2 1 10 9 1 10 9 13 0 10 9 1 10 11 1 9 2 10 9 0 2 11 11 11 2 9 1 11 11 2 11 2 2
52 10 9 3 0 1 10 9 0 2 1 10 9 1 10 9 0 2 10 9 1 9 1 9 2 10 9 1 9 13 1 9 0 7 10 9 0 1 10 9 0 2 4 13 15 1 9 1 10 9 3 0 2
29 13 9 1 10 0 2 9 0 2 3 1 10 11 1 9 2 10 11 0 7 10 11 1 11 16 13 1 9 2
41 3 15 13 10 9 1 10 9 1 10 11 11 1 9 1 10 11 1 11 2 9 1 9 0 16 1 10 9 4 13 1 10 0 9 1 9 1 10 9 0 2
16 11 11 11 13 1 11 2 11 2 10 12 1 11 1 12 2
32 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2 9 2 11 2
51 10 9 1 10 9 13 16 15 13 10 0 9 0 2 7 16 3 13 9 1 10 12 9 16 1 10 9 15 4 13 1 9 0 2 1 10 9 11 11 2 1 10 11 1 11 11 7 11 1 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
40 0 9 4 13 10 9 2 1 1 9 10 9 1 11 1 10 11 2 11 11 11 2 7 10 11 1 11 11 1 10 11 2 11 11 11 2 2 11 2 2
19 10 9 1 10 9 13 1 10 0 9 1 9 1 10 15 10 12 13 2
35 3 1 12 9 1 9 15 13 1 10 9 1 11 2 16 13 1 1 10 9 1 10 9 1 12 9 2 13 13 1 11 7 1 11 2
17 10 9 15 13 3 13 1 10 13 15 0 1 13 10 9 0 2
16 11 11 11 13 1 11 11 1 11 10 12 1 11 1 12 2
35 1 9 2 10 9 11 1 10 9 0 2 13 10 9 0 1 10 15 1 10 12 9 2 9 16 3 3 15 13 16 10 9 4 13 2
24 10 9 4 3 13 1 10 0 9 11 2 10 15 3 4 13 15 3 1 10 9 1 12 2
54 3 2 4 13 16 10 9 13 0 1 15 16 13 10 0 11 2 3 15 13 10 9 0 1 10 9 1 13 10 9 0 1 10 9 7 9 1 9 0 1 10 9 0 2 1 10 16 15 13 10 9 1 9 2
28 2 10 11 11 2 2 2 11 11 2 2 13 10 9 13 1 10 9 1 10 11 11 1 10 9 1 9 2
40 4 13 1 11 11 11 1 10 9 1 10 0 9 2 11 11 11 2 16 15 13 10 9 0 7 10 9 0 1 10 9 1 13 10 9 1 9 3 0 2
53 11 11 2 3 1 10 9 0 1 13 1 11 11 11 1 10 9 1 10 9 1 11 7 4 13 10 11 2 13 10 9 0 13 1 15 0 1 10 9 1 11 11 11 2 11 2 1 10 9 0 1 12 2
62 1 9 2 16 1 10 9 15 15 13 10 9 2 10 9 13 1 9 1 9 3 1 10 0 9 2 7 3 3 10 9 15 13 1 9 0 2 1 10 9 0 7 0 1 10 9 2 2 15 13 10 9 1 16 10 9 13 3 0 7 0 2
19 11 1 11 15 13 10 9 1 13 10 9 1 11 11 2 1 9 0 2
24 3 1 10 9 4 13 9 1 10 11 1 12 7 12 2 7 9 1 11 1 12 7 12 2
28 10 9 4 13 15 15 2 13 1 10 9 1 10 9 7 15 13 1 13 2 7 13 10 9 7 10 9 2
19 11 4 13 3 1 10 9 12 1 10 9 1 9 2 2 11 11 2 2
10 3 10 9 15 13 1 8 7 8 2
50 11 2 3 1 10 0 9 0 7 0 1 10 9 0 2 13 10 9 1 10 9 7 9 1 10 9 0 2 0 1 10 9 1 11 7 10 11 2 9 0 2 1 11 2 9 1 10 9 2 2
10 15 13 0 3 15 13 1 10 9 2
22 10 9 1 10 9 13 1 10 9 2 13 1 12 9 0 1 10 0 9 1 9 2
25 10 9 1 10 9 15 13 1 12 16 13 10 9 1 9 0 1 10 9 1 10 9 1 9 2
37 15 2 13 1 10 9 2 15 13 10 9 1 10 9 1 3 2 13 15 1 10 9 1 10 15 13 11 11 2 11 11 2 7 11 11 2 2
16 3 1 13 1 10 9 2 10 9 13 11 2 11 2 11 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
22 4 13 1 10 9 0 0 11 10 12 1 11 1 12 3 1 10 9 11 2 11 2
13 11 3 15 13 1 15 7 4 13 1 10 9 2
24 10 9 1 9 1 9 15 4 1 13 1 11 11 11 11 1 10 9 1 11 11 1 12 2
62 10 9 4 13 1 10 3 0 9 0 11 11 2 15 4 13 1 11 1 11 1 12 1 9 0 7 9 9 2 7 15 13 10 10 9 9 1 13 1 10 9 1 11 2 16 3 4 13 1 10 9 1 10 9 7 10 9 1 13 10 9 2
57 10 9 3 0 7 15 16 13 11 13 2 1 15 9 2 1 13 16 10 9 1 9 16 13 9 1 10 9 0 2 3 7 10 9 16 15 13 3 7 3 2 7 1 10 9 10 9 13 0 2 4 9 1 10 9 0 2
37 13 12 9 1 10 9 2 10 9 12 13 10 3 0 2 13 1 9 0 1 10 9 13 7 4 13 9 1 10 9 0 1 15 7 12 9 2
20 3 13 10 9 2 13 16 13 0 2 10 9 15 13 7 3 13 1 3 2
17 10 9 1 10 9 0 13 16 13 10 9 13 1 2 11 2 2
7 13 10 9 1 9 0 2
19 11 13 10 9 1 12 9 1 9 1 9 0 1 10 9 1 10 9 2
7 10 9 0 13 3 0 2
30 15 13 1 12 9 1 10 9 1 12 2 15 1 12 7 10 15 1 12 2 16 13 10 9 1 13 10 9 0 2
36 3 15 13 10 9 11 11 11 11 7 10 11 11 1 10 11 7 10 9 2 9 1 10 11 1 10 11 2 10 11 11 7 10 11 11 2
38 10 9 1 11 11 13 10 9 7 10 11 11 13 3 1 10 0 9 16 13 1 10 11 11 11 7 15 13 3 10 11 1 13 11 13 10 9 2
30 1 10 9 2 16 13 1 9 1 12 9 2 13 10 9 1 9 10 9 1 9 1 10 9 0 11 1 10 11 2
18 3 1 10 9 2 11 13 10 9 0 1 10 9 1 13 1 11 2
31 13 1 16 1 10 9 11 11 13 10 9 0 13 1 11 2 4 13 10 9 2 1 10 9 7 15 1 10 0 9 2
19 1 10 0 12 9 13 1 11 7 1 11 3 13 1 10 9 11 11 2
89 3 3 13 0 10 9 0 1 10 9 1 10 9 1 9 2 13 15 13 10 9 1 10 9 2 2 10 9 1 10 0 9 1 10 9 4 13 7 4 13 10 9 1 10 9 1 10 9 1 10 9 2 13 15 15 3 3 3 13 15 10 9 0 7 10 9 2 7 16 13 10 9 13 1 10 9 16 15 13 1 10 9 1 10 9 1 10 9 2
19 7 3 1 10 11 13 10 0 9 0 0 9 1 10 11 2 10 9 2
25 10 9 1 9 2 11 11 2 13 1 10 9 9 0 7 1 10 9 10 9 0 1 10 9 2
17 10 9 4 13 9 1 13 1 10 9 0 1 10 9 1 9 2
42 1 9 13 3 1 10 9 1 9 0 11 2 11 13 16 10 9 4 13 1 10 0 9 1 11 1 10 9 1 10 9 2 11 11 2 1 10 16 15 0 13 2
10 9 0 7 9 0 1 10 0 9 2
12 11 13 9 1 10 9 2 1 9 0 2 2
40 10 9 15 13 1 10 9 0 2 13 15 1 10 9 3 3 0 1 10 10 9 1 11 2 13 15 1 10 9 0 7 0 1 10 9 0 1 10 9 2
24 10 9 4 13 1 10 9 2 1 10 9 1 10 11 7 10 0 9 2 1 11 1 12 2
34 10 9 15 13 1 9 1 10 9 0 2 7 1 9 1 9 1 9 7 9 2 9 7 9 2 9 1 10 9 0 1 10 9 2
21 10 9 7 9 0 1 10 9 15 13 9 1 10 9 7 0 9 1 10 9 2
9 2 1 15 13 1 13 1 9 2
16 1 12 15 13 9 1 9 7 10 9 1 10 9 1 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
31 3 1 10 9 1 9 2 10 11 13 1 10 9 9 2 10 9 1 9 2 12 9 0 13 1 9 7 10 0 9 2
11 13 0 9 7 10 0 9 1 9 0 2
19 11 13 10 9 13 1 10 9 1 9 1 10 9 7 9 1 10 9 2
19 1 10 9 1 10 9 1 12 2 13 11 11 2 0 9 1 10 9 2
16 10 9 11 13 1 10 9 10 9 1 10 9 1 10 9 2
23 13 16 10 9 13 10 0 9 1 9 0 16 15 13 10 9 0 7 9 1 10 9 2
22 1 9 2 13 16 10 9 4 13 12 9 1 10 9 2 3 10 9 7 10 9 2
30 10 9 9 0 1 12 5 9 2 12 5 9 2 7 9 0 1 3 10 10 9 2 12 12 9 7 12 9 2 2
19 15 3 13 7 15 3 13 13 2 3 2 15 8 8 7 15 8 8 2
27 10 11 11 13 10 9 0 1 12 2 13 1 11 11 2 13 1 10 9 1 10 0 9 1 11 11 2
45 3 1 16 15 13 1 13 10 9 2 10 9 1 9 2 11 11 2 13 16 1 10 9 0 2 13 10 9 1 0 9 7 9 16 4 13 1 11 1 10 9 1 9 2 2
30 7 16 3 15 13 2 1 10 9 15 13 1 10 9 1 9 1 10 9 16 13 15 7 3 13 1 16 15 13 2
66 11 11 2 11 2 11 2 12 1 11 1 12 2 2 13 1 2 11 2 2 13 10 9 1 9 0 0 16 13 3 10 9 1 11 5 12 1 10 11 11 2 11 11 11 2 3 1 10 9 11 11 11 9 15 13 1 10 9 1 10 9 1 10 9 12 2
27 10 9 4 13 1 9 15 13 1 13 2 1 15 13 10 9 0 7 0 1 9 0 7 0 1 9 2
3 13 3 2
13 3 12 1 10 9 13 1 10 9 1 9 0 2
12 13 9 1 10 9 0 1 10 9 1 12 2
20 15 13 11 11 11 2 2 16 13 10 9 1 10 9 1 11 11 7 11 2
26 1 0 2 13 10 9 7 13 15 16 13 0 1 15 1 10 9 1 10 9 1 11 1 10 11 2
33 10 9 7 9 13 1 3 9 1 10 9 13 1 11 7 10 16 4 13 16 15 13 16 13 10 9 1 9 2 1 9 2 2
14 3 3 2 13 1 10 9 1 16 15 13 10 9 2
19 3 13 1 11 2 3 4 13 3 1 11 7 13 1 15 1 10 9 2
19 13 15 15 3 16 1 9 13 0 16 10 9 13 1 3 1 12 9 2
19 13 1 10 9 1 9 7 9 0 2 9 1 10 9 1 9 15 13 2
14 1 0 2 10 9 15 13 1 10 9 1 12 9 2
17 12 1 11 1 12 2 13 10 8 9 0 16 13 1 9 0 2
28 16 10 9 13 1 10 9 0 2 11 13 16 15 13 1 10 9 0 2 13 1 10 9 1 10 0 9 2
33 11 13 10 11 12 2 1 13 12 9 1 9 1 9 1 10 9 0 16 13 1 9 1 10 9 1 13 15 10 9 1 9 2
12 10 9 13 1 13 10 9 0 1 10 9 2
23 3 15 13 10 0 9 1 10 11 1 10 9 1 11 2 1 9 1 10 9 1 8 2
7 13 1 9 1 9 0 2
31 10 9 13 1 10 11 1 11 2 3 11 1 11 2 11 7 11 2 2 4 10 9 13 1 10 11 1 11 7 11 2
19 10 9 1 11 2 1 10 10 9 2 4 13 1 9 1 10 9 0 2
24 1 12 15 13 1 13 1 11 2 11 2 2 3 13 9 1 10 9 1 9 1 9 0 2
60 10 9 1 10 11 11 2 11 11 2 4 13 3 16 15 13 10 2 0 9 2 13 9 1 9 1 10 9 7 4 13 16 15 13 16 10 9 13 16 3 4 13 9 1 2 9 7 9 2 2 7 3 4 13 0 1 10 9 0 2
12 13 9 0 1 9 0 0 1 10 9 11 2
15 10 9 15 13 3 7 11 13 10 9 1 11 1 12 2
9 15 13 15 16 13 7 15 9 2
56 1 15 15 13 1 16 15 13 10 9 2 4 1 13 1 9 10 9 1 10 9 11 8 5 12 2 16 13 9 16 13 13 10 9 1 9 0 2 9 0 1 9 16 1 10 9 15 13 1 9 1 9 7 9 9 2
16 10 9 13 3 1 10 9 1 10 9 7 10 9 1 9 2
49 11 3 15 13 3 0 7 10 9 1 10 9 1 0 9 7 13 16 10 9 16 13 10 9 1 9 13 1 0 13 7 2 10 9 1 16 10 9 1 11 13 3 1 11 13 3 15 2 2
13 1 10 9 15 4 13 1 10 9 1 10 9 2
19 3 1 9 2 10 9 4 13 1 10 9 0 1 11 11 7 11 11 2
22 1 10 9 2 11 11 2 13 10 0 9 1 9 1 10 9 2 16 15 13 0 2
15 1 9 2 13 15 1 10 9 0 1 9 1 11 11 2
21 10 9 4 13 1 10 9 1 9 2 11 11 2 1 10 9 1 10 9 0 2
25 11 11 11 11 2 3 13 1 11 2 13 10 12 1 11 1 12 2 13 10 8 2 9 0 2
12 1 10 9 1 12 15 13 3 1 12 9 2
21 10 9 3 0 15 13 10 9 13 10 1 13 1 10 9 1 13 10 9 0 2
61 1 10 9 15 13 1 10 9 13 16 10 9 13 1 10 9 1 9 1 9 2 7 1 9 10 9 2 9 1 11 1 12 2 4 1 13 15 1 10 0 9 13 1 10 9 2 10 12 1 11 1 12 2 13 1 10 9 1 10 9 2
27 1 10 11 9 10 0 9 15 13 1 10 11 2 1 12 1 12 2 13 1 11 7 9 1 0 9 2
42 13 1 10 9 3 13 9 1 10 9 1 13 1 10 9 2 1 13 15 1 10 0 2 9 2 11 2 15 15 13 1 15 1 4 1 13 1 15 1 10 9 2
27 10 11 11 1 11 11 2 11 2 13 10 9 3 0 1 9 0 2 13 9 0 1 9 1 10 11 2
18 15 13 1 10 9 3 0 1 10 11 1 10 11 1 11 7 11 2
34 10 0 9 2 11 11 2 4 13 2 13 3 0 10 9 1 13 9 2 9 1 9 2 7 1 0 2 13 9 1 10 9 0 2
53 15 13 1 9 1 13 1 10 9 0 2 11 11 2 13 1 10 11 2 2 16 10 9 1 10 9 11 11 2 11 2 13 10 9 7 13 12 9 1 10 9 2 13 15 16 13 10 9 1 10 9 11 2
31 7 10 0 9 1 9 13 1 10 9 0 1 10 9 1 10 11 1 11 2 13 15 1 10 12 9 7 13 12 9 2
40 3 13 1 11 2 16 13 15 1 10 9 2 16 15 13 10 9 16 15 13 3 1 10 9 2 7 10 9 16 3 13 1 10 0 9 13 1 10 9 2
18 10 9 1 10 9 0 13 10 9 0 3 13 1 11 2 11 2 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
38 1 11 11 2 11 13 10 11 11 11 2 10 0 9 13 1 11 11 2 11 1 10 9 2 11 1 11 9 12 2 7 1 10 9 1 10 9 2
12 13 9 1 10 11 2 1 10 9 1 11 2
70 9 1 11 13 3 7 13 2 1 9 2 1 10 0 9 13 1 16 15 13 3 13 15 2 11 13 10 9 13 2 2 10 9 1 10 9 15 13 16 13 15 16 15 4 13 7 13 1 10 9 1 11 7 13 10 9 1 10 11 1 10 11 16 13 10 9 1 11 2 2
20 13 16 15 13 1 10 9 0 7 3 3 2 9 1 15 15 13 3 9 2
48 1 10 9 13 9 1 10 0 9 1 10 11 11 11 2 11 11 2 10 9 1 10 9 11 2 10 9 11 11 2 11 11 1 11 2 10 9 11 11 11 7 10 9 10 9 11 11 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
29 13 1 10 9 1 10 3 0 2 11 11 2 13 1 10 0 9 7 15 13 13 1 10 9 1 11 7 11 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
61 7 1 9 10 9 2 9 2 4 13 10 9 0 1 13 1 13 1 10 9 8 10 9 0 1 10 11 11 2 10 11 11 11 2 10 11 11 1 10 11 2 13 13 1 10 9 1 10 9 10 9 1 10 9 7 10 9 1 10 9 2
28 11 11 2 12 2 12 2 13 10 9 2 11 2 9 0 2 13 9 1 10 2 11 11 11 1 11 2 2
54 10 9 0 13 16 10 9 15 13 1 11 2 11 7 1 10 9 11 1 10 11 1 10 11 7 1 10 15 15 13 10 9 1 9 2 9 2 1 10 9 0 9 1 10 9 0 8 9 0 7 9 1 9 2
23 10 0 9 1 9 3 13 10 9 1 10 9 0 7 9 1 10 9 1 11 7 11 2
19 10 9 1 9 13 1 12 8 5 5 5 2 12 8 5 8 5 2 2
23 13 10 9 0 4 13 15 3 10 9 0 1 13 1 10 15 15 4 13 10 9 0 2
12 3 13 1 13 16 3 13 15 4 13 15 2
8 1 9 2 10 9 4 13 2
18 10 9 16 15 4 13 13 15 2 7 3 10 9 3 15 4 13 2
24 1 10 0 9 10 9 15 13 3 0 7 0 2 1 10 9 1 13 10 9 1 10 9 2
15 13 10 0 9 1 9 7 15 16 3 13 15 15 13 2
19 3 7 3 2 1 12 2 10 9 13 10 8 1 11 3 1 10 11 2
16 11 3 4 13 9 0 7 9 1 9 1 13 9 3 0 2
17 7 2 1 13 10 9 0 13 9 13 1 9 10 9 0 8 2
41 10 9 13 1 12 5 1 10 12 5 1 10 9 0 7 12 5 1 10 9 0 13 15 1 10 11 11 11 11 10 10 12 5 1 10 9 0 1 10 9 2
8 10 9 1 9 13 5 8 2
15 10 9 2 1 10 9 2 13 1 10 9 1 10 9 2
48 10 9 13 1 10 9 1 10 9 1 10 9 11 11 2 0 13 7 16 8 4 7 13 1 10 9 11 11 2 12 2 2 16 15 13 1 9 0 16 15 13 1 8 1 10 0 9 2
44 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 13 10 9 1 10 11 1 11 11 1 11 7 9 7 8 2 9 1 10 9 1 9 1 9 7 10 9 0 2
15 1 10 9 2 10 9 0 13 3 9 1 9 1 13 2
22 15 4 13 15 2 10 9 0 2 10 0 9 2 10 9 0 2 7 10 9 0 2
32 10 11 1 11 1 11 2 11 2 11 1 11 1 11 2 13 10 0 9 1 9 1 11 1 10 11 13 1 11 2 11 2
15 13 10 9 1 10 9 16 15 13 2 13 15 1 15 2
31 10 9 0 1 10 9 3 7 10 9 1 9 4 13 15 1 10 10 9 1 10 9 2 5 2 1 10 9 1 9 2
34 10 9 1 10 9 13 0 9 2 16 3 10 9 0 1 9 7 9 0 13 1 10 9 1 10 9 1 10 9 1 10 9 11 2
13 15 13 1 9 2 11 2 11 2 7 11 11 2
26 15 13 10 9 16 13 12 9 2 13 3 1 10 9 0 2 0 1 9 2 16 13 12 9 3 2
14 10 9 0 13 1 11 13 11 11 7 9 11 11 2
22 1 10 9 3 1 12 9 13 1 12 9 1 9 2 1 10 9 0 1 12 9 2
46 10 9 1 10 9 1 12 9 0 1 10 9 15 4 13 13 1 3 1 12 0 2 1 3 1 12 9 2 1 10 9 2 7 0 9 7 9 2 10 15 13 7 13 10 9 2
7 2 11 11 8 8 0 2
11 15 13 0 2 11 2 11 7 11 2 2
20 10 9 13 13 1 10 9 13 3 1 9 10 9 1 10 9 7 10 9 2
11 3 10 9 1 12 9 13 15 16 13 2
13 4 1 13 12 5 1 10 9 1 9 16 13 2
17 10 9 1 11 2 11 7 11 13 10 9 1 10 10 9 0 2
13 11 13 1 9 10 9 3 0 1 10 0 11 2
16 1 15 16 13 9 2 4 13 15 1 10 0 9 10 9 2
18 11 13 15 1 10 12 9 1 15 4 13 3 10 9 0 1 11 2
29 3 15 13 1 10 9 10 15 15 13 12 9 3 0 7 1 10 10 9 1 10 9 2 9 16 13 3 0 2
41 1 12 2 10 9 0 0 1 12 9 13 1 12 9 2 1 15 12 13 10 9 0 2 12 10 9 2 12 10 9 2 12 15 2 12 15 7 12 3 13 2
23 10 11 11 11 2 11 2 13 15 1 10 12 9 0 0 1 10 11 1 10 11 11 2
8 11 15 13 13 1 10 9 2
13 3 7 11 13 3 2 9 0 1 15 9 2 2
17 10 9 13 10 9 1 11 7 13 10 9 1 3 1 12 9 2
15 16 13 10 9 15 13 9 7 9 2 9 7 9 2 2
26 13 1 10 11 11 2 13 10 9 2 1 10 12 9 2 7 1 9 4 13 1 9 1 10 9 2
28 1 11 1 10 9 2 11 13 1 10 9 0 10 11 11 3 1 15 1 10 9 1 9 3 0 1 11 2
42 10 9 0 1 10 9 15 13 1 10 9 13 1 10 9 11 11 2 11 2 11 2 2 16 13 1 10 9 1 9 1 10 0 9 1 10 9 2 11 11 2 2
21 15 13 1 12 2 13 10 0 1 13 15 1 9 1 10 9 1 10 11 11 2
39 3 2 10 9 13 0 10 9 1 10 9 12 1 10 16 15 13 1 10 9 0 1 13 15 1 10 9 1 9 1 10 9 3 0 1 13 10 9 2
29 1 11 1 12 13 1 10 11 11 1 11 11 1 11 2 1 10 13 10 9 0 7 13 1 15 1 11 11 2
15 13 13 1 13 16 10 9 13 1 10 11 11 1 9 2
33 10 9 1 10 9 1 11 11 15 13 0 1 9 7 9 1 10 12 9 1 9 2 9 1 10 16 13 0 10 9 0 0 2
16 10 9 2 3 1 9 0 2 13 10 9 13 1 10 9 2
32 10 9 1 10 9 12 2 13 10 9 1 12 9 1 10 9 1 12 9 5 2 1 10 9 0 1 12 9 1 9 5 2
26 11 13 10 9 9 12 1 11 2 10 9 0 1 10 9 7 13 10 9 1 4 13 3 1 15 2
19 3 13 10 9 1 10 9 0 1 10 9 1 11 2 3 1 10 9 2
25 3 0 2 1 10 0 9 4 13 10 9 9 1 10 9 16 15 13 10 9 16 13 11 11 2
16 10 9 1 10 11 4 13 3 1 10 9 1 11 7 9 2
19 11 13 16 13 4 13 1 10 9 7 16 13 3 1 10 9 1 9 2
35 3 4 13 0 9 1 13 15 10 9 16 13 1 9 1 10 9 1 11 2 11 7 11 7 3 13 2 1 10 13 1 11 1 11 2
12 1 10 9 13 10 11 1 10 11 1 11 2
22 10 9 13 1 10 9 16 13 3 15 3 9 13 2 9 2 9 7 1 15 9 2
36 4 13 1 15 1 10 9 1 9 2 13 10 9 0 1 10 9 7 13 1 12 10 0 9 1 10 9 0 2 10 9 1 9 7 9 2
42 0 1 10 11 8 11 11 2 1 11 1 12 2 11 13 1 10 9 1 12 9 1 9 1 10 11 16 13 1 9 1 9 7 1 9 0 1 9 1 10 11 2
43 1 9 2 10 0 9 1 10 9 12 2 12 2 1 10 9 1 10 0 9 16 3 15 13 1 10 11 1 11 2 13 10 9 1 10 9 10 12 1 11 1 12 2
31 1 10 9 15 15 13 3 1 13 10 9 1 9 2 1 10 9 2 7 9 2 4 15 13 3 10 9 1 10 9 2
27 10 9 0 1 13 10 9 13 1 10 9 1 9 2 7 10 9 13 16 0 9 13 0 1 10 9 2
56 1 10 9 12 7 12 2 10 9 1 10 9 4 13 3 0 2 13 1 10 9 1 10 9 7 10 9 2 3 7 1 10 9 1 10 9 0 7 0 13 1 10 9 0 7 10 9 1 10 11 7 10 9 1 11 2
23 1 10 9 1 9 1 10 11 11 1 11 2 4 13 10 9 1 0 9 1 10 9 2
21 10 1 10 9 4 13 1 10 11 11 7 13 10 0 9 0 1 11 1 11 2
26 13 1 10 9 1 11 2 4 9 2 11 11 2 2 15 16 13 9 1 15 13 9 1 10 9 2
32 11 13 10 9 7 9 0 2 1 10 9 1 11 2 11 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
12 10 9 1 11 11 15 13 13 1 10 9 2
21 13 1 10 9 1 12 9 10 9 13 12 8 12 9 7 15 13 1 12 9 2
42 10 9 0 7 0 2 0 7 0 1 10 9 13 10 9 13 1 10 9 16 13 3 4 13 10 9 1 9 2 4 13 15 1 15 9 1 3 12 9 1 9 2
24 13 0 16 10 9 13 10 7 10 9 1 10 9 1 13 10 9 1 10 9 1 9 0 2
27 11 13 10 9 1 11 2 15 1 9 3 0 2 10 9 1 13 1 11 1 10 0 9 0 1 9 2
12 10 9 4 13 13 10 12 9 1 9 0 2
19 12 7 12 1 11 2 1 9 1 10 9 1 10 11 7 1 11 11 2
15 10 9 13 10 9 1 10 9 3 13 0 9 1 9 2
7 10 9 13 11 1 9 2
50 10 9 2 10 9 2 10 9 7 10 9 13 3 13 1 10 9 2 1 9 1 10 10 9 3 15 13 10 9 7 10 9 2 12 9 3 0 7 13 0 1 10 9 7 10 15 1 10 15 2
14 10 0 9 13 10 9 0 1 10 11 1 10 11 2
13 13 10 0 9 1 11 0 1 9 1 10 11 2
24 11 2 10 9 0 2 1 10 15 13 10 11 11 2 13 0 0 7 13 3 1 10 9 2
19 11 11 2 9 1 9 2 13 10 9 1 9 0 2 1 10 9 11 2
19 1 9 2 10 9 1 11 13 1 10 9 13 16 10 9 1 9 13 2
17 10 9 1 9 1 10 9 2 13 10 9 1 10 9 1 11 2
17 11 11 11 12 13 9 1 10 9 0 3 1 11 11 11 12 2
19 10 9 16 15 13 1 10 9 1 10 11 4 7 13 3 1 15 9 2
10 4 3 13 1 9 0 7 1 9 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
58 10 9 3 1 10 9 2 10 9 11 11 13 1 11 11 11 15 9 2 2 13 7 10 9 15 13 1 10 9 2 7 16 10 9 13 10 9 16 13 11 11 1 12 2 10 9 15 13 1 10 9 1 9 1 0 9 2 2
26 13 16 1 3 10 10 9 2 10 9 15 13 1 11 2 3 16 10 9 1 9 0 13 10 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
15 1 9 9 9 1 10 11 11 2 13 9 1 10 9 2
18 1 10 9 1 10 11 11 11 2 11 1 9 13 10 9 3 0 2
23 10 9 1 11 2 10 11 1 11 2 1 9 2 13 10 9 13 1 11 11 1 12 2
70 15 15 13 1 16 1 10 9 15 13 12 9 2 16 13 1 10 9 8 1 10 9 12 2 1 10 9 0 2 15 4 13 1 10 0 9 2 7 1 10 11 11 1 11 2 11 11 2 10 9 12 7 12 1 11 1 12 2 1 10 9 0 1 10 9 2 11 11 2 2
20 13 10 9 2 7 3 4 1 13 16 15 13 16 13 9 7 16 13 9 2
22 10 9 0 13 3 9 2 7 3 4 4 13 10 9 1 9 1 9 1 10 9 2
17 1 10 9 10 9 1 10 9 13 0 7 1 9 0 3 0 2
13 10 10 9 1 10 9 13 0 1 10 9 0 2
25 1 10 9 1 13 10 0 9 3 7 3 1 10 9 2 13 0 9 1 9 1 9 7 9 2
26 13 3 16 13 1 13 10 9 2 13 9 0 7 0 3 4 13 12 0 9 0 7 10 11 11 2
38 10 0 9 13 10 9 0 1 10 9 1 9 1 9 9 1 10 9 1 10 0 9 0 2 1 9 1 9 1 11 11 1 10 9 1 9 0 2
12 3 3 13 2 15 13 13 3 1 12 9 2
14 13 0 4 13 1 10 9 1 9 1 9 1 15 2
9 11 11 13 9 1 10 9 0 2
11 10 9 13 15 7 10 9 13 3 3 2
34 1 11 11 1 11 11 13 1 11 2 7 13 10 9 1 10 9 2 7 3 1 10 9 2 13 1 10 9 10 9 1 10 9 2
29 1 13 10 9 1 9 0 7 10 9 1 9 1 10 9 2 10 9 4 13 9 0 1 10 9 1 10 9 2
10 15 13 1 15 8 10 9 1 9 2
4 13 1 11 2
15 1 9 1 13 0 7 0 4 13 10 9 1 10 9 2
22 10 11 1 11 1 10 11 1 11 13 15 1 10 9 0 1 10 9 0 1 11 2
8 13 10 0 9 1 0 9 2
14 3 13 0 10 9 7 2 1 0 2 10 10 9 2
20 10 9 0 1 11 11 11 15 13 1 10 9 1 10 0 9 0 7 0 2
32 3 15 4 13 1 10 9 1 15 0 16 4 13 10 9 1 10 9 1 9 2 3 7 3 13 13 3 9 1 10 9 2
12 3 13 1 11 11 2 11 11 7 11 11 2
30 2 11 13 1 10 9 1 10 9 16 13 13 1 10 2 9 2 11 11 1 10 0 9 2 2 13 10 0 9 2
29 10 11 1 11 13 3 10 9 1 15 1 10 9 16 13 1 10 9 3 1 7 15 13 10 9 1 11 12 2
8 10 9 1 10 11 1 11 2
9 4 13 10 0 9 1 10 9 2
14 3 13 1 11 11 1 10 9 10 11 1 11 11 2
6 13 1 9 1 9 2
25 0 9 15 13 1 10 9 2 16 3 13 15 1 10 0 9 1 9 1 10 9 1 10 11 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
18 3 13 10 9 1 10 9 2 7 1 10 9 1 13 1 10 9 2
44 11 11 15 13 1 10 9 1 13 1 10 12 1 11 2 3 1 7 10 9 0 4 4 7 13 15 1 10 9 10 9 13 1 9 1 9 13 1 10 9 1 10 9 2
34 11 2 9 1 10 9 7 10 9 2 13 1 11 2 11 2 7 13 10 9 1 12 9 2 13 10 9 10 9 0 11 11 1 8
17 8 10 12 9 13 9 1 10 9 1 9 0 1 11 2 11 2
27 1 12 9 13 1 11 11 2 10 9 13 1 10 9 0 1 10 9 1 9 0 3 13 1 10 9 2
50 4 13 3 0 1 10 9 7 15 13 1 15 1 13 15 16 13 15 10 9 2 10 9 0 1 10 9 13 15 16 15 13 2 7 1 15 2 16 15 4 13 10 9 0 2 7 10 0 9 2
38 3 1 13 3 1 11 7 1 13 1 10 9 1 10 9 2 10 9 15 13 1 10 9 1 9 9 1 10 9 2 9 7 9 0 1 0 9 2
12 10 9 15 13 13 15 1 9 7 13 15 2
12 10 12 5 1 10 9 13 1 10 9 0 2
33 15 13 13 7 13 2 1 15 15 13 0 13 15 10 9 0 16 13 3 13 15 1 10 9 1 10 9 7 13 1 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 8 2
28 1 10 12 7 12 9 1 10 9 1 10 11 2 13 10 9 16 3 13 9 1 10 11 1 10 9 0 2
19 3 11 11 13 10 2 9 8 2 1 10 9 3 0 1 10 11 11 2
6 4 13 1 10 11 2
30 1 10 9 2 10 9 12 12 12 13 1 3 1 15 1 10 9 1 9 1 10 9 2 3 1 9 1 9 0 2
31 13 10 9 0 1 11 10 9 1 10 0 9 3 4 13 7 13 10 9 0 1 0 9 7 3 13 1 10 9 11 2
10 4 13 1 10 9 0 1 12 9 2
15 10 9 1 9 0 13 10 16 13 10 9 1 10 9 2
27 10 9 13 2 10 9 1 12 9 10 15 13 1 10 9 2 13 0 1 10 9 2 2 1 4 13 2
37 1 10 9 12 10 9 0 4 1 13 1 10 9 2 7 3 1 10 9 1 10 9 0 1 10 9 12 15 13 3 10 9 7 9 1 9 2
24 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 1 10 11 2
22 11 13 10 9 1 9 1 15 16 13 0 1 13 10 9 1 0 9 1 10 11 2
46 13 1 15 16 1 9 1 11 11 7 1 10 9 11 11 2 13 13 10 9 1 10 9 0 7 1 9 8 1 10 9 13 11 11 11 2 2 10 11 1 11 1 11 2 2 2
19 11 11 13 10 9 1 11 2 16 13 10 9 0 7 0 1 10 9 2
13 10 0 9 2 12 2 15 13 1 9 1 12 2
14 1 0 10 9 3 0 3 7 13 10 9 1 9 2
37 10 9 4 13 1 10 9 1 9 1 10 9 1 10 9 7 10 9 16 13 3 0 2 15 13 9 3 7 3 4 13 15 3 1 10 9 2
41 0 1 10 9 0 1 9 1 9 7 9 1 11 2 11 11 11 2 10 11 13 10 2 9 0 2 1 13 1 10 9 1 9 1 9 2 9 7 9 0 2
22 1 9 10 9 1 9 3 13 0 7 10 9 7 9 4 4 13 1 11 3 0 2
18 13 9 1 10 9 1 11 2 11 1 11 1 12 7 11 1 12 2
6 13 10 12 9 13 2
10 10 9 4 4 13 1 10 0 9 2
60 1 10 0 9 1 10 16 10 9 13 0 2 10 9 0 4 13 3 3 1 12 9 8 2 16 13 9 0 1 10 9 1 9 1 10 9 2 1 1 9 9 1 9 2 9 0 2 9 0 2 10 9 11 11 7 9 1 10 9 2
21 11 7 11 15 4 13 1 3 1 10 11 7 11 13 10 9 1 9 1 12 2
13 13 13 10 0 9 1 10 9 1 10 11 11 2
10 4 13 1 10 11 11 1 9 0 2
39 13 15 1 10 9 1 3 9 1 10 9 2 1 10 15 15 4 13 9 1 9 0 2 7 4 13 13 1 9 0 1 10 9 1 9 1 9 0 2
41 1 9 1 10 9 2 10 9 11 7 3 9 0 1 10 11 2 11 4 13 15 2 2 3 2 2 11 2 4 13 9 1 10 9 0 2 1 10 9 0 2
11 10 9 4 13 1 9 1 9 7 9 2
27 3 15 13 1 10 9 10 9 1 10 11 1 11 11 11 2 16 15 4 13 1 11 16 13 10 9 2
36 15 13 1 9 15 10 0 9 2 15 13 1 10 9 2 11 2 3 1 10 9 2 7 2 15 13 16 15 13 10 9 0 1 10 9 2
8 13 9 0 1 10 9 0 2
14 13 10 9 1 9 1 9 2 0 2 9 7 0 2
21 15 13 1 0 2 7 1 9 1 13 2 9 1 10 9 2 2 1 9 0 2
34 2 13 16 10 9 1 10 9 4 4 13 1 10 9 0 7 10 9 2 7 13 10 9 16 10 9 4 13 16 13 10 9 2 2
35 10 12 1 11 1 12 2 10 11 11 1 11 7 10 9 1 11 11 11 13 1 10 9 10 9 1 9 2 13 15 1 10 9 11 2
27 1 12 15 13 10 11 1 10 9 1 9 1 11 2 1 10 15 11 11 1 11 13 10 2 9 2 2
22 10 9 13 1 10 9 7 13 7 3 13 9 1 16 3 4 13 9 1 10 9 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
41 10 12 1 11 1 12 2 13 3 9 1 10 11 2 15 13 16 11 4 13 10 9 1 12 9 1 10 8 8 8 0 1 10 9 0 1 12 9 1 9 2
25 1 11 2 10 11 13 9 1 10 9 0 1 11 2 9 16 13 1 10 13 15 1 10 9 2
29 11 2 11 2 11 11 11 13 9 1 10 11 11 11 7 9 1 11 11 11 1 10 9 7 1 11 11 11 2
11 15 13 10 9 1 10 9 0 1 11 2
15 2 13 16 11 13 10 9 2 7 15 3 13 13 0 2
32 1 10 9 1 10 9 1 12 2 10 9 0 1 9 1 10 9 13 1 9 12 2 7 10 9 0 1 9 13 9 12 2
43 3 15 13 9 7 3 10 0 9 3 15 13 2 3 7 15 4 13 1 10 9 16 4 13 2 15 16 13 16 3 13 10 9 3 0 2 1 15 10 0 9 2 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 12 2
16 11 15 13 1 11 11 16 13 10 9 16 13 10 11 11 2
54 16 11 1 11 13 10 9 1 9 0 16 13 9 8 1 9 0 7 13 1 10 9 16 13 2 13 2 7 13 9 0 1 9 2 3 13 9 1 16 10 9 13 10 8 2 8 7 9 1 9 1 10 9 2
27 1 10 9 13 3 15 1 10 9 0 3 0 1 15 15 13 9 1 9 1 13 3 1 12 12 9 2
9 13 10 9 0 1 10 9 0 2
21 11 13 3 13 2 7 13 10 9 1 10 9 13 15 16 4 4 13 1 15 2
13 13 9 1 10 9 0 1 11 2 11 2 11 2
38 3 2 1 10 9 1 13 10 9 0 1 10 9 1 10 9 2 13 16 13 10 9 1 9 1 9 1 10 9 10 9 1 9 0 1 10 9 2
19 10 9 1 11 1 9 0 13 10 9 3 0 1 9 0 1 9 0 2
43 10 9 1 11 4 13 1 15 1 3 0 1 10 9 1 11 2 15 15 4 1 7 10 9 0 13 1 10 9 0 2 9 3 0 2 9 1 0 9 7 9 2 2
23 10 9 1 9 13 10 9 1 10 9 0 9 2 16 15 13 3 0 1 10 9 0 2
82 9 2 9 2 9 2 9 2 9 0 2 9 2 9 2 9 0 2 9 2 9 2 9 2 9 2 11 2 2 9 2 11 2 9 2 2 9 2 9 2 2 9 2 10 9 10 0 1 0 2 9 0 2 9 2 9 2 2 9 2 12 9 2 2 9 2 9 2 2 9 2 9 2 9 2 9 2 9 2 9 2 8
31 13 10 0 7 3 0 9 1 9 0 1 10 9 1 12 9 1 9 0 2 12 1 9 0 7 12 9 1 12 9 2
43 11 11 2 11 11 2 12 2 13 10 9 0 0 2 16 4 13 10 0 9 1 10 9 1 9 2 3 9 2 9 2 9 7 9 2 3 1 10 9 1 10 9 2
11 13 13 10 9 1 10 9 1 10 9 2
16 15 13 1 9 0 7 13 10 9 0 1 10 1 10 11 2
49 15 13 2 1 10 9 2 1 10 9 3 0 1 13 10 9 1 10 9 1 11 1 11 2 15 13 1 12 9 7 12 9 2 9 1 13 3 2 2 13 3 1 10 9 1 10 0 9 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
14 10 9 1 9 13 16 10 9 15 13 1 10 9 2
11 10 9 13 3 1 10 9 1 10 9 2
59 1 10 12 9 2 11 13 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 9 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
16 15 13 10 9 1 9 2 4 15 13 10 9 1 10 9 2
35 1 9 0 1 10 9 0 1 10 11 13 0 13 10 9 2 0 9 0 2 2 2 0 9 0 11 11 13 3 9 0 1 11 2 2
41 1 9 2 10 9 1 10 11 1 11 11 7 11 11 11 13 0 1 10 9 16 13 10 9 1 11 11 11 11 7 13 13 10 0 9 1 10 11 11 11 2
15 10 12 13 9 0 1 9 7 9 0 13 9 1 9 2
39 1 10 9 1 10 9 2 10 9 0 1 9 0 3 15 13 1 9 7 9 2 1 10 9 1 10 9 7 10 9 7 15 1 10 9 7 10 9 2
41 1 9 2 15 13 3 1 9 1 9 0 1 0 9 2 1 10 15 15 13 0 9 1 9 2 16 13 10 9 2 7 1 15 16 13 10 9 2 3 0 2
27 11 2 3 1 13 7 13 10 9 1 11 11 2 15 13 10 12 1 11 1 10 9 0 1 11 11 2
16 10 9 13 3 0 2 13 10 10 9 7 10 9 0 0 2
19 10 9 0 1 9 13 12 2 3 16 10 9 13 0 1 10 9 0 2
25 10 9 13 10 9 0 1 11 11 2 13 9 1 10 11 2 11 2 2 11 2 11 7 11 2
17 13 10 9 1 9 1 13 10 9 7 10 9 7 9 1 0 2
31 10 9 15 13 12 9 1 9 16 13 1 10 11 11 12 1 9 1 10 11 1 10 11 1 10 11 11 11 1 12 2
32 11 11 12 13 10 9 1 10 0 9 1 11 11 11 2 7 13 1 9 1 11 11 11 2 7 10 9 1 11 11 11 2
31 15 16 3 13 12 7 3 9 16 13 1 10 3 12 9 1 10 9 1 12 3 13 0 2 13 15 16 13 10 11 2
30 0 9 3 13 3 7 13 10 9 16 13 1 10 9 3 0 7 10 9 2 16 13 13 10 9 0 2 2 13 2
62 1 10 12 9 2 10 9 1 11 13 0 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
20 10 9 4 13 0 7 13 10 9 1 10 0 9 7 4 13 1 9 0 2
32 3 3 2 11 4 13 16 2 1 3 2 10 9 13 9 1 10 9 3 0 2 16 4 13 10 9 0 2 10 11 2 2
8 11 15 13 13 1 10 9 2
13 1 10 9 13 10 9 1 10 11 1 11 11 2
21 3 15 13 16 10 9 16 13 13 0 1 10 9 3 1 3 9 2 11 11 2
38 3 2 10 9 13 10 9 1 12 9 2 7 1 10 9 15 13 12 2 13 1 10 9 1 10 9 1 3 2 16 3 4 13 15 0 1 9 2
16 3 15 13 10 0 9 8 9 1 10 12 9 1 11 11 2
38 1 10 9 0 2 10 9 0 13 0 7 4 4 13 1 9 0 2 0 2 9 2 8 2 1 10 9 1 10 0 9 7 10 9 15 4 13 2
15 10 9 13 1 12 2 12 2 12 2 12 7 12 9 2
13 13 1 10 9 2 15 13 1 10 9 1 11 2
23 13 1 10 9 0 8 2 12 7 8 2 12 2 3 4 13 3 7 1 10 9 0 2
17 10 9 4 4 13 1 12 9 2 1 10 9 12 2 1 11 2
23 11 11 4 4 13 1 10 9 16 13 1 10 9 1 11 2 3 7 4 4 13 3 2
85 10 9 0 13 1 10 9 12 16 10 11 1 11 7 11 2 11 2 13 10 9 1 10 11 11 1 10 11 11 1 11 11 1 11 7 11 2 11 2 2 13 1 10 9 1 10 9 13 11 11 10 9 1 10 9 0 0 1 10 9 1 10 9 16 13 1 9 10 9 0 1 10 9 0 1 10 9 7 10 9 0 1 10 9 2
8 15 13 12 9 1 9 0 2
30 10 9 13 1 12 11 7 10 9 13 1 11 1 12 2 16 10 9 3 13 9 1 10 12 1 11 1 10 9 2
24 7 15 1 9 1 16 11 0 3 13 10 9 1 10 11 7 13 10 9 0 2 10 9 2
33 3 3 2 1 10 9 12 2 10 9 4 13 1 0 9 2 8 2 1 11 2 15 1 10 9 1 11 1 10 9 1 11 2
24 1 10 11 1 10 11 10 9 13 10 9 1 10 9 1 11 2 11 7 10 9 1 11 2
33 10 2 11 11 11 2 4 13 1 15 1 10 12 9 3 0 1 10 9 7 9 7 15 15 13 10 9 0 1 10 9 0 2
8 13 0 1 10 11 1 11 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
28 10 9 0 2 9 1 10 9 0 2 11 11 2 4 13 10 12 1 11 1 12 1 10 9 1 12 9 2
28 1 9 15 13 1 10 9 7 1 0 1 10 9 1 9 0 1 9 0 7 1 10 9 1 10 0 9 2
22 10 9 1 10 9 13 11 11 11 2 7 13 1 10 9 1 11 7 11 2 11 2
23 11 13 10 9 1 10 9 1 10 11 2 1 10 9 1 11 2 11 7 11 2 11 2
23 3 0 2 10 9 13 13 10 11 11 7 13 10 9 1 10 9 1 12 1 10 11 2
24 3 2 7 1 13 10 9 1 10 9 2 13 10 9 1 9 7 10 9 13 1 11 11 2
21 10 9 1 9 4 4 13 1 10 0 9 1 10 9 0 16 13 1 10 9 2
25 11 13 10 9 16 3 15 13 1 9 0 7 9 2 16 3 13 10 16 10 9 1 9 0 2
50 10 9 13 1 10 11 1 11 1 11 7 10 9 13 10 9 1 10 9 0 1 9 1 10 9 0 1 11 2 1 9 1 10 0 9 1 10 9 0 11 8 11 2 13 1 10 9 1 11 2
32 10 9 1 9 7 9 13 0 1 13 10 12 9 16 13 1 10 9 1 9 2 10 9 0 7 10 9 0 1 13 15 2
22 2 3 13 15 10 0 9 16 10 9 7 9 1 11 13 1 15 1 10 0 9 2
25 10 0 9 1 10 9 3 4 13 9 1 9 2 1 9 7 1 0 9 1 13 1 0 9 2
22 11 13 1 9 1 11 1 10 9 12 1 10 9 11 1 10 9 0 11 8 11 2
11 1 9 1 10 9 13 12 9 0 0 2
19 13 1 10 9 1 11 11 16 10 9 4 13 7 13 3 1 10 9 2
28 1 9 0 13 9 10 9 0 11 11 2 15 3 3 13 1 11 2 13 1 10 9 1 11 2 3 13 2
29 10 9 1 11 15 13 0 2 7 10 9 13 10 9 13 16 15 13 1 10 9 15 13 1 9 1 13 15 2
42 10 9 1 9 2 13 9 1 10 9 0 16 15 13 1 9 3 1 13 16 4 0 7 15 13 10 0 9 1 10 9 0 2 9 7 9 2 7 10 9 0 2
45 13 10 12 9 13 1 10 9 2 1 10 9 0 2 10 9 1 10 9 2 10 9 13 10 9 7 9 1 10 0 9 1 10 9 11 11 2 7 10 9 0 1 10 9 2
63 1 9 1 10 0 9 2 10 9 1 10 9 4 1 13 15 1 9 1 10 0 9 2 11 13 3 13 16 10 9 9 13 10 9 2 11 3 4 13 7 13 1 10 9 2 11 13 10 9 1 11 7 11 13 16 10 9 13 1 11 1 13 2
21 1 9 1 10 9 2 13 10 9 2 9 7 9 1 10 11 1 9 0 9 2
16 3 2 13 10 9 1 9 0 7 13 1 9 1 10 9 2
53 10 9 15 4 13 1 10 9 1 9 1 10 9 2 7 1 10 13 15 15 13 10 9 13 1 9 1 10 9 2 7 3 10 9 1 9 9 1 10 9 2 11 2 11 11 2 11 2 7 2 11 2 2
44 3 13 9 2 1 10 9 0 9 1 10 9 13 1 9 0 2 3 16 13 10 9 0 1 10 9 0 2 16 10 9 13 3 9 1 10 9 1 9 0 1 10 9 2
13 15 13 10 9 1 12 9 7 9 1 10 9 2
31 13 16 13 9 1 10 9 0 2 7 16 1 10 9 1 9 13 3 10 9 0 13 9 13 7 13 16 3 3 13 2
20 3 13 10 0 9 1 10 9 2 7 3 1 9 3 13 9 1 0 9 2
32 1 9 2 1 9 1 10 9 2 11 11 13 3 1 10 9 1 10 9 1 10 0 9 16 13 10 9 0 13 11 11 2
25 10 9 11 11 13 1 12 9 0 1 10 9 1 10 0 9 1 10 9 1 2 9 0 2 2
36 13 10 9 1 10 9 1 12 9 7 13 2 3 2 10 9 1 13 10 9 16 3 9 4 13 1 10 11 11 1 15 9 1 10 9 2
13 10 9 1 10 9 1 11 2 11 13 12 12 2
35 1 3 10 9 1 10 9 2 16 13 1 10 9 0 1 10 9 1 10 9 0 1 10 9 2 3 7 10 9 1 10 9 3 0 2
39 10 11 11 1 11 2 1 9 10 11 11 11 2 13 10 0 9 1 9 1 9 0 0 16 4 13 1 10 9 1 9 0 1 15 9 1 10 9 2
14 11 11 11 13 3 1 10 9 1 11 11 1 12 2
7 10 9 13 10 9 0 2
9 10 11 4 13 1 9 1 12 2
27 10 9 1 10 9 2 10 9 7 9 1 10 9 2 13 1 10 9 2 13 1 10 9 1 13 15 2
33 11 11 2 10 9 0 1 11 1 10 11 0 2 13 10 0 9 13 15 1 10 9 1 10 9 7 9 3 0 1 10 9 2
30 10 11 7 3 10 11 13 1 1 10 9 1 11 11 7 3 13 15 16 13 10 11 2 10 12 9 1 9 3 2
21 10 9 1 10 9 0 13 16 2 3 15 4 13 10 9 0 1 10 9 2 2
21 1 10 9 1 12 15 15 13 1 11 10 9 1 12 9 2 13 10 12 9 2
19 10 9 1 11 13 10 9 0 16 4 13 9 1 1 12 1 12 9 2
23 10 11 11 11 13 3 1 9 1 10 11 11 11 2 13 3 1 10 9 1 11 11 2
25 10 9 0 9 4 13 9 1 9 3 0 9 1 9 1 11 1 9 2 9 2 7 9 9 2
21 1 11 3 13 1 10 9 2 10 9 15 13 1 13 1 2 10 11 11 2 2
21 10 9 1 10 9 2 11 11 7 11 11 2 13 10 0 9 1 10 0 9 2
39 10 9 4 13 1 9 1 9 1 11 2 0 3 1 10 9 1 11 2 7 11 2 1 9 13 11 2 0 15 1 10 11 7 1 9 1 11 2 2
44 10 9 11 11 2 1 10 9 11 11 2 1 10 9 11 2 11 2 4 13 1 10 9 1 11 7 11 1 10 0 7 10 9 1 11 2 13 10 9 1 10 9 11 2
50 3 2 13 16 11 13 10 9 0 15 10 9 13 1 15 3 13 9 2 11 15 13 1 10 9 1 10 9 0 2 10 15 15 13 11 1 10 9 15 11 11 2 13 13 3 10 9 1 9 2
57 2 3 2 13 2 2 10 9 16 13 1 3 2 10 9 1 15 13 0 3 12 9 0 1 10 0 12 9 7 10 9 2 3 15 4 13 10 9 13 1 10 9 2 10 9 0 7 13 15 16 15 13 1 10 9 2 2
40 11 2 11 2 1 2 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2 11 2 1 2 11 2
23 13 10 9 3 1 10 9 16 13 9 1 10 11 11 1 11 2 15 16 13 10 9 2
32 10 9 1 9 13 10 9 1 11 2 15 16 13 13 7 13 10 9 0 2 1 11 15 4 13 3 13 1 12 9 2 2
29 10 9 1 11 1 9 0 13 1 10 9 15 13 3 13 1 10 9 1 10 9 0 1 11 7 10 9 0 2
33 11 13 10 9 7 9 0 2 13 1 10 9 1 11 11 2 9 1 11 2 1 10 9 1 11 2 11 7 9 1 15 11 2
20 13 3 2 3 15 4 13 15 3 3 9 7 4 13 10 9 1 9 0 2
44 4 13 10 9 0 1 10 9 2 13 1 12 2 7 1 11 1 10 11 2 10 9 1 10 9 1 11 1 10 9 0 2 13 1 12 1 9 1 11 1 10 11 2 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
12 1 10 9 0 15 13 10 9 7 10 9 2
22 3 13 10 9 1 10 9 1 9 1 10 9 1 10 9 1 12 2 11 12 2 2
16 1 12 13 1 10 11 11 11 11 7 13 10 9 1 9 2
47 10 9 15 4 13 3 1 2 11 2 11 2 1 10 9 1 10 9 1 12 3 15 13 3 10 9 0 2 13 13 9 7 9 1 10 9 0 7 13 15 15 1 9 1 10 9 2
8 10 9 0 13 1 12 9 2
21 1 10 9 1 12 2 10 9 13 1 12 9 2 12 9 7 12 9 8 0 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
42 10 9 13 1 13 1 10 9 9 9 1 9 16 15 13 1 10 9 16 13 10 9 16 15 13 1 3 1 10 9 7 3 13 10 0 1 13 3 1 10 9 2
31 10 9 2 1 10 13 15 2 15 13 1 10 9 0 7 1 10 9 7 15 1 9 13 9 7 9 2 9 7 9 2
23 10 11 1 11 4 13 3 10 9 1 11 1 10 9 1 0 9 0 1 10 10 9 2
15 11 1 11 2 10 0 9 1 9 16 13 3 1 11 2
17 12 9 3 2 1 10 12 2 12 2 13 1 10 11 11 11 2
26 11 13 0 1 16 10 9 2 1 9 1 9 2 15 4 13 10 9 1 13 9 1 10 0 9 2
18 13 10 9 3 0 1 10 9 7 13 1 10 11 13 10 10 9 2
15 11 11 11 2 11 2 11 2 12 1 11 1 12 2 2
13 4 13 7 13 10 9 1 10 9 1 9 11 2
30 10 9 0 13 4 13 1 10 9 1 2 11 11 2 10 9 1 13 1 10 9 16 13 15 16 13 2 1 3 2
27 15 13 1 10 9 0 9 1 10 9 1 9 7 9 16 13 10 9 1 9 1 10 9 0 1 11 2
21 1 10 9 12 10 9 13 10 0 9 2 1 10 9 1 10 9 1 10 9 2
24 10 9 1 11 13 10 9 0 0 2 13 1 10 9 1 11 7 10 9 1 11 2 11 2
47 3 15 13 16 4 13 7 16 13 4 13 1 10 9 2 1 10 9 2 16 10 9 13 1 11 1 12 2 10 9 13 11 11 11 2 10 9 0 1 11 11 2 7 3 1 11 2
19 13 10 9 11 1 10 11 1 10 9 13 1 10 9 1 11 1 12 2
19 11 11 13 1 12 1 9 1 9 7 11 11 13 9 1 9 1 12 2
28 15 4 13 15 1 9 0 2 0 1 10 9 1 9 0 2 3 13 0 7 13 1 0 9 1 10 9 2
22 3 13 16 10 11 11 13 3 1 10 10 9 2 13 13 1 10 9 1 10 9 2
13 1 9 3 13 9 16 10 9 13 0 7 0 2
20 10 9 4 13 1 10 9 1 12 9 1 11 2 15 4 13 1 11 11 2
45 1 10 9 1 9 0 2 10 9 3 4 13 13 9 1 15 16 1 9 15 13 2 7 13 3 10 9 12 1 11 1 10 9 1 13 10 9 1 11 16 3 4 13 3 2
69 10 9 1 10 9 15 13 1 9 1 10 9 12 2 16 10 9 1 9 1 9 0 0 1 10 9 11 11 2 0 1 15 1 0 9 1 10 9 2 1 9 1 10 9 1 10 9 2 13 13 10 9 1 0 9 7 15 1 9 2 15 1 9 7 3 10 9 0 2
54 15 16 3 13 3 1 11 11 13 2 13 1 10 0 9 0 10 9 2 7 13 16 10 9 1 10 9 2 1 15 13 1 10 9 0 2 13 2 0 2 16 2 4 13 9 7 1 10 9 1 10 9 2 2
36 13 1 9 1 4 13 0 1 11 2 3 16 13 3 9 0 2 7 1 11 2 16 13 1 10 0 9 2 4 13 2 13 3 10 9 2
20 10 2 9 1 9 0 2 13 10 9 0 1 10 9 7 10 9 1 9 2
18 10 9 13 10 9 0 1 9 12 9 1 10 9 12 1 10 9 2
15 1 10 9 2 15 15 4 1 13 3 1 11 1 11 2
25 1 9 1 13 10 9 0 7 9 1 13 10 9 0 2 3 10 11 0 13 3 1 10 9 2
12 13 10 9 0 7 10 9 0 1 9 0 2
30 0 1 12 9 2 11 13 9 1 10 9 1 10 0 9 1 9 1 10 9 9 1 10 9 1 10 9 7 9 2
21 13 16 1 15 9 1 10 9 4 13 1 10 9 0 2 10 9 7 10 9 2
18 1 11 1 12 2 10 11 11 4 13 12 9 1 10 9 1 9 2
20 10 9 2 1 10 9 11 11 11 2 11 1 11 2 11 11 2 12 2 2
54 1 10 9 10 11 1 10 11 11 1 11 11 4 13 1 10 3 9 11 11 11 1 9 0 1 10 9 1 10 9 0 1 10 9 1 10 12 1 11 1 12 2 4 13 1 10 7 3 13 10 12 1 11 2
15 10 9 4 13 3 1 13 15 1 9 13 1 10 9 2
14 11 2 13 10 9 1 9 0 0 1 10 9 11 2
17 11 14 2 13 10 9 1 11 11 1 12 1 13 9 1 11 2
14 1 10 9 7 13 1 10 11 11 12 10 0 9 2
29 3 15 13 10 8 3 0 13 1 15 1 10 9 1 0 1 10 9 2 13 9 1 15 11 11 7 11 11 2
74 1 9 1 10 9 11 11 2 0 9 1 9 1 10 9 0 2 7 16 1 15 15 13 10 9 0 2 2 1 11 13 10 9 1 16 10 9 0 3 4 4 13 1 10 9 1 9 1 10 11 7 16 2 1 10 9 2 4 13 10 2 9 1 10 9 2 1 9 1 10 9 0 9 2
22 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 11 2
17 13 1 12 7 12 9 2 1 16 13 15 7 12 1 10 9 2
22 11 13 1 10 9 0 2 13 15 0 1 2 2 10 9 1 2 10 0 9 2 2
15 3 1 11 1 12 2 11 13 10 9 1 10 9 0 2
19 10 9 1 10 9 1 11 15 13 0 2 1 9 2 1 10 9 0 2
9 13 1 10 9 0 1 10 9 2
28 10 11 1 11 1 11 11 2 11 2 2 13 15 16 13 1 0 9 1 9 2 1 12 9 7 12 9 2
72 10 0 9 3 1 10 9 11 13 3 1 11 11 2 1 10 11 11 11 11 1 11 1 12 7 10 0 9 1 10 9 1 10 11 11 11 3 1 11 11 1 11 1 12 2 13 15 10 0 9 16 10 11 11 13 1 9 11 2 3 15 13 1 11 2 1 0 3 1 10 9 2
30 10 9 0 15 13 3 3 2 16 10 9 0 13 9 1 9 1 11 2 15 16 13 9 1 10 0 9 1 9 2
8 1 0 9 13 13 10 9 2
26 1 9 2 15 13 3 1 13 1 9 1 10 9 2 11 7 11 2 13 16 3 13 9 1 13 2
11 15 13 1 11 2 1 10 11 11 11 2
19 1 9 1 10 11 11 2 0 1 10 9 0 1 10 11 1 10 11 2
21 7 15 9 13 16 10 9 1 10 9 3 13 15 7 13 3 1 10 9 0 2
49 1 11 2 11 2 11 2 11 7 10 9 1 10 9 4 13 10 9 1 8 2 9 7 9 2 7 7 10 11 2 11 12 7 11 9 13 10 8 5 1 9 1 10 9 0 7 10 9 2
37 10 11 13 1 9 1 10 11 1 11 11 2 13 1 10 11 12 1 15 1 10 10 9 1 4 13 9 0 1 10 9 1 10 11 11 11 2
24 10 9 2 9 13 1 10 9 2 8 2 13 9 1 10 9 0 15 13 5 10 9 0 2
20 10 9 16 13 0 2 15 13 1 9 0 2 10 9 2 13 9 13 0 2
19 1 9 1 11 1 10 12 13 10 9 0 13 11 2 11 2 11 11 2
24 13 1 10 11 1 12 7 10 9 1 9 15 13 1 10 11 11 2 1 9 1 12 9 2
34 15 3 13 13 0 9 1 10 9 1 10 9 7 1 10 9 2 13 15 1 13 0 9 7 13 0 9 2 9 1 10 15 13 2
26 1 10 9 10 9 13 1 10 9 1 10 9 0 1 11 13 11 2 3 13 3 1 15 1 11 2
24 7 3 1 10 9 1 11 2 11 11 2 1 12 9 2 16 13 10 0 9 1 10 9 2
16 1 11 13 11 2 11 2 11 11 7 11 2 13 1 11 2
58 1 11 10 9 7 10 9 1 10 9 13 9 1 10 11 11 2 9 16 15 13 1 10 9 16 3 13 1 10 0 12 9 7 16 13 10 9 1 9 1 10 11 16 15 13 1 10 12 1 11 7 10 12 1 11 1 12 2
37 9 3 13 10 9 0 1 10 13 10 10 9 13 1 10 9 0 2 1 15 10 1 3 13 9 0 7 9 0 1 10 9 0 7 1 11 2
5 10 9 4 13 2
15 10 9 0 16 13 1 9 13 3 0 7 13 3 0 2
12 10 9 1 9 1 10 9 13 1 5 12 2
19 1 10 12 9 0 1 10 9 0 1 9 2 3 12 13 1 10 9 2
30 1 13 15 1 9 0 1 0 1 10 13 10 9 1 10 11 2 11 13 10 9 1 10 9 1 9 1 10 11 2
18 11 11 13 10 11 11 2 7 11 11 11 13 15 0 1 10 9 2
21 11 11 2 13 10 9 1 9 11 1 10 9 11 2 16 13 1 10 9 11 2
21 3 15 13 10 9 1 11 11 2 3 10 1 11 2 13 1 10 9 1 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
14 10 9 16 13 10 9 13 9 3 1 10 9 0 2
19 1 10 9 1 10 9 1 11 11 2 15 13 1 15 1 10 9 0 2
36 10 9 1 9 15 13 1 9 3 1 10 9 2 3 16 15 4 13 10 0 9 1 10 9 1 9 1 10 9 7 10 9 0 1 9 2
33 1 10 9 0 3 0 16 13 11 15 13 10 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 11 7 11 11 11 2
29 15 8 13 16 13 9 1 9 7 3 15 13 1 13 2 16 13 10 9 3 0 7 13 0 8 1 13 9 2
29 10 11 1 10 11 13 2 1 0 2 0 2 1 9 1 10 9 2 1 10 9 1 9 7 1 10 0 9 2
21 10 9 0 13 16 10 0 9 0 1 9 0 3 1 11 4 4 13 1 9 2
18 15 3 2 1 9 2 13 3 0 7 10 15 2 7 13 10 9 2
8 13 9 1 10 9 11 11 2
28 10 9 1 10 10 9 7 1 10 9 13 1 10 9 0 10 11 2 7 1 10 9 3 13 9 0 10 2
27 10 9 1 9 7 9 0 2 1 10 9 0 2 13 0 1 13 1 10 9 1 10 9 1 10 9 2
18 10 9 1 11 13 9 0 3 13 1 9 1 9 1 13 0 9 2
26 10 11 13 10 9 1 9 13 1 9 2 7 11 13 1 10 9 1 10 9 0 13 1 11 11 2
10 10 11 13 10 9 1 9 3 0 2
36 10 0 9 1 10 9 0 3 13 13 7 3 0 9 2 10 11 11 1 10 9 1 11 2 10 11 1 10 11 2 2 4 13 1 9 2
12 11 11 13 10 9 1 9 1 10 9 11 2
17 1 9 13 10 9 1 13 16 10 9 15 13 16 13 1 9 2
24 10 0 9 15 13 1 10 9 1 15 11 2 10 9 0 2 4 13 16 10 9 13 0 2
51 10 11 1 11 1 10 11 1 10 11 11 2 13 1 12 2 15 13 1 9 7 9 16 4 13 2 0 9 1 10 9 2 9 7 9 2 1 10 9 7 10 9 7 1 10 9 1 10 9 0 2
21 10 9 13 0 16 4 13 1 3 2 1 10 9 0 3 9 7 10 9 0 2
55 1 10 9 1 10 9 0 0 10 9 13 0 1 10 9 2 1 16 4 13 1 12 1 10 9 2 16 15 13 1 10 9 1 11 1 13 15 1 10 9 1 10 9 1 10 11 11 2 3 15 13 1 10 9 2
24 10 9 1 11 7 11 2 1 10 15 15 13 2 13 1 10 9 10 12 1 11 1 12 2
67 10 0 9 1 10 9 0 2 11 2 11 1 11 2 11 2 11 2 11 2 11 2 11 0 2 11 0 2 11 2 11 2 11 7 10 0 9 1 10 11 4 1 13 1 10 9 1 9 0 3 0 9 1 10 11 2 11 2 10 11 2 10 11 7 10 11 2
15 10 9 8 0 1 11 2 3 1 10 9 7 0 9 2
77 9 1 10 11 1 10 11 1 11 2 4 13 1 9 1 11 11 2 1 9 2 7 11 10 11 2 1 9 2 2 11 11 1 12 3 1 9 2 10 9 1 10 9 13 16 13 1 10 0 7 0 9 1 9 1 15 13 11 11 2 11 11 2 11 11 7 11 11 7 10 9 1 9 1 11 11 2
20 13 1 9 10 9 7 10 11 2 3 7 10 9 13 9 7 9 3 0 2
26 1 10 11 1 11 2 15 13 10 9 2 16 10 9 11 15 13 13 9 0 1 10 9 0 0 2
43 15 13 10 0 9 1 12 9 2 1 10 9 10 9 0 1 10 9 7 13 1 10 9 7 10 9 1 10 9 7 1 10 9 10 9 7 10 9 0 1 10 9 2
41 10 12 1 11 1 12 2 10 9 9 4 13 1 9 1 10 9 1 10 9 1 10 11 11 11 2 9 1 10 9 2 2 7 13 1 10 9 1 10 9 2
22 1 12 7 12 2 11 13 1 3 1 12 9 10 9 1 10 9 1 13 1 11 2
15 1 3 10 9 1 10 9 15 13 3 0 1 10 9 2
27 1 10 9 1 10 9 1 9 2 1 9 1 10 9 12 2 13 10 9 2 10 9 16 3 13 15 2
34 9 16 13 10 9 3 13 7 1 10 9 16 13 13 16 13 15 3 7 3 2 1 10 9 2 7 10 9 3 3 13 1 15 2
18 1 10 9 10 9 1 9 15 13 15 1 9 7 1 9 1 9 2
21 3 4 13 1 10 9 1 10 9 1 11 2 9 1 11 2 1 10 9 11 2
17 13 10 9 12 1 10 0 9 7 10 9 16 15 13 1 11 2
35 1 10 9 16 13 10 9 11 11 4 4 4 13 1 9 0 7 9 1 9 0 16 3 4 4 4 13 1 9 1 9 1 10 9 2
40 10 9 1 10 11 15 13 2 1 15 2 16 13 9 1 9 0 1 10 15 13 12 7 3 9 2 13 10 9 0 16 13 4 13 10 9 1 10 9 2
12 13 10 9 12 3 3 3 10 9 13 0 2
25 11 13 2 13 13 10 9 1 10 9 2 13 1 10 9 3 0 1 10 9 1 10 9 0 2
13 10 9 13 10 0 9 1 10 9 1 10 9 2
27 1 12 10 9 0 11 1 11 15 13 3 0 1 11 2 10 9 0 7 1 10 9 1 11 7 11 2
26 11 13 3 1 11 11 11 7 11 11 11 1 9 1 9 1 4 13 1 10 9 1 10 12 9 2
10 11 0 13 10 9 1 10 9 11 2
8 11 15 13 13 1 10 9 2
24 13 10 0 9 2 7 3 13 13 15 1 10 8 2 8 2 13 10 9 1 12 5 9 2
42 3 15 13 10 9 15 1 13 10 9 3 2 1 10 9 7 0 2 7 15 15 13 3 2 3 15 13 10 8 0 1 9 9 7 3 15 13 1 10 9 2 8
48 16 4 13 10 9 1 9 2 4 4 13 1 11 1 10 9 2 13 10 9 7 3 13 1 3 1 12 9 1 15 2 15 4 13 1 13 15 1 10 9 13 1 10 0 9 1 11 2
18 10 9 13 1 10 9 0 16 13 9 3 1 9 0 1 10 9 2
5 15 13 1 11 2
52 10 11 13 2 16 13 2 1 10 9 0 1 12 9 2 12 8 12 2 2 13 11 12 11 2 9 11 11 13 1 12 8 12 8 1 8 2 12 8 1 9 7 10 15 13 1 10 9 1 12 9 2
36 1 3 2 10 9 16 13 13 10 9 7 13 1 11 2 16 13 12 9 1 12 9 7 16 13 3 9 3 1 10 9 7 3 1 15 2
19 1 11 13 1 10 9 1 9 4 13 15 10 9 1 9 1 0 9 2
26 10 9 13 3 12 9 2 10 9 0 3 1 9 1 9 2 7 10 9 9 1 15 7 1 9 2
16 10 9 4 13 1 10 9 1 10 0 1 2 10 9 2 2
35 10 9 1 13 1 15 1 10 9 1 9 3 0 2 4 13 10 9 0 1 13 2 13 10 9 1 13 10 9 16 13 1 10 9 2
17 10 9 7 10 9 1 10 9 12 7 12 13 1 9 0 9 2
13 10 9 0 4 13 9 1 10 3 1 10 9 2
9 13 1 11 2 11 2 1 12 2
42 11 13 1 10 9 1 10 9 2 13 0 7 10 9 3 3 13 1 15 2 13 9 0 1 13 9 0 2 13 10 9 0 7 0 13 9 0 1 0 9 2 8
22 10 9 0 13 3 10 9 1 10 9 0 7 10 9 1 10 9 13 1 10 9 2
20 11 11 11 2 13 1 11 11 2 13 10 9 16 15 15 13 1 15 9 2
26 13 1 12 2 10 9 1 9 1 11 11 12 4 13 1 11 11 7 13 1 9 2 9 7 9 2
34 13 1 11 11 11 2 13 1 11 1 2 11 11 2 1 11 11 2 12 2 2 13 1 2 11 2 7 2 11 11 2 1 11 2
30 1 10 9 1 10 9 2 10 9 1 10 9 2 15 13 1 10 9 0 1 10 9 1 10 9 1 10 9 0 2
43 10 9 1 10 9 1 10 9 11 13 1 10 9 16 10 11 4 13 13 1 10 12 1 10 12 1 11 1 9 1 9 2 1 15 15 10 9 15 13 1 10 9 2
24 13 10 0 9 15 16 13 1 10 9 1 10 11 11 1 10 9 1 12 1 12 5 0 2
47 4 13 1 10 9 0 1 11 2 11 2 1 10 9 0 1 10 9 11 2 9 1 11 11 2 12 9 1 10 9 1 11 7 12 9 1 10 9 1 11 2 10 9 1 10 11 2
17 10 12 0 1 10 9 7 10 12 0 0 13 1 10 0 9 2
29 1 9 0 7 1 13 10 9 1 9 1 10 9 1 9 2 10 9 3 13 1 10 9 2 7 1 9 0 2
29 10 9 1 10 0 9 13 1 10 11 1 11 11 2 10 0 9 1 10 9 0 11 11 2 1 10 9 12 2
26 15 13 10 11 16 13 7 10 9 13 1 10 1 10 9 2 3 13 7 3 1 10 9 3 0 2
27 1 10 9 0 1 9 0 2 11 13 10 9 1 12 9 5 16 13 9 1 10 9 1 11 1 11 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
11 3 2 11 3 4 13 10 9 3 0 2
32 1 10 0 9 13 3 0 0 9 1 10 9 1 10 9 0 1 2 10 9 1 10 9 2 7 0 9 13 1 9 11 2
25 11 11 2 10 9 0 1 9 1 11 1 11 11 2 4 13 10 9 3 1 10 11 1 11 2
50 11 7 11 2 1 9 0 2 2 11 3 7 1 10 9 0 0 2 13 10 9 1 11 2 11 11 2 13 1 10 9 1 10 9 0 2 3 13 11 7 11 2 1 10 9 1 10 11 11 2
29 1 10 9 0 1 9 0 7 0 2 10 9 4 13 1 10 9 9 1 10 9 1 10 11 11 1 11 12 2
42 10 9 16 13 4 13 10 9 1 3 7 13 10 9 0 1 10 9 1 10 10 9 2 3 4 13 10 9 16 15 13 2 7 13 15 16 13 1 10 0 9 2
5 15 13 9 0 2
37 1 9 1 10 9 2 1 12 10 9 4 1 13 10 9 1 10 11 7 2 3 2 1 10 9 0 2 13 13 15 3 0 7 15 3 0 2
27 15 3 13 7 13 10 9 0 7 3 0 9 1 9 1 10 9 2 16 10 9 13 3 13 10 9 2
23 10 9 13 1 10 9 1 10 9 2 2 11 2 1 9 7 2 11 2 1 10 9 2
20 2 13 0 16 3 1 10 9 1 10 1 10 11 15 13 9 1 10 9 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
65 1 10 9 15 4 13 9 7 9 1 10 9 1 10 9 2 1 15 15 10 9 15 4 13 3 12 9 2 13 10 9 1 10 9 1 10 15 3 13 10 9 0 7 13 1 9 10 9 16 13 1 10 9 1 9 1 10 9 2 16 3 4 13 15 2
28 13 1 10 0 9 1 10 11 1 10 11 11 2 10 9 2 11 2 4 13 1 9 0 1 11 1 12 2
54 3 1 15 2 13 11 2 10 9 1 11 2 2 3 0 1 9 2 7 11 3 11 2 10 9 11 1 10 9 11 2 3 13 1 11 2 2 15 4 1 13 1 11 1 13 10 11 1 13 2 13 10 9 2
58 7 3 2 10 9 0 1 10 9 1 9 2 4 13 10 12 1 11 1 12 1 10 11 1 11 2 3 13 11 1 11 2 2 13 1 9 16 1 13 13 0 13 1 9 13 1 9 1 9 2 9 7 9 1 9 1 9 2
60 1 10 9 10 9 1 9 0 4 13 10 9 0 7 1 10 13 9 3 13 1 10 9 1 10 9 2 13 16 10 9 0 15 13 10 0 9 1 10 9 7 3 1 10 9 2 16 3 2 1 9 3 2 13 0 1 10 9 0 2
22 13 3 0 16 10 9 1 10 9 0 13 1 13 10 9 3 0 1 10 15 9 2
16 16 10 9 13 0 10 9 13 3 1 1 10 9 1 9 2
40 1 10 9 1 9 16 13 9 1 10 9 1 10 9 1 11 2 10 9 13 1 13 9 1 10 9 1 10 9 1 10 9 7 16 13 1 2 11 2 2
23 10 9 0 13 1 10 0 9 1 10 9 9 2 13 1 10 9 2 13 1 10 9 2
21 1 10 11 1 12 2 13 1 11 2 11 2 13 9 1 11 1 9 1 9 2
21 10 9 13 13 1 10 9 11 2 11 2 13 1 10 9 11 11 11 2 11 2
32 10 9 0 1 9 1 10 11 13 15 16 3 9 4 13 2 16 11 7 11 3 4 13 10 9 1 9 1 10 0 9 2
41 10 9 1 9 15 13 7 15 13 1 13 10 9 1 10 9 1 11 2 13 1 10 9 2 16 4 13 9 1 10 9 1 9 0 1 10 9 1 10 9 2
51 10 9 16 15 13 9 0 0 13 13 3 9 1 10 9 1 10 9 9 2 13 3 10 9 1 10 9 1 11 1 3 1 10 9 11 2 7 3 2 3 13 10 9 11 1 10 9 1 9 0 2
27 10 9 3 13 15 7 10 9 1 11 11 11 2 11 11 2 15 3 4 1 13 10 9 1 10 9 2
60 3 3 2 10 9 13 16 3 15 13 10 9 1 9 7 16 3 4 1 13 1 10 9 9 1 0 2 9 1 10 9 2 13 1 10 9 7 9 1 10 9 2 1 15 15 1 10 9 1 10 9 15 13 10 9 1 0 2 9 2
21 10 9 15 13 10 12 1 11 1 12 7 15 13 3 10 12 1 11 1 12 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
49 13 10 2 8 2 2 3 15 13 10 9 0 1 9 2 13 10 9 0 1 13 1 10 0 9 1 10 9 0 7 13 10 9 0 1 10 9 2 1 10 9 1 10 9 7 13 9 0 2
27 10 9 1 10 9 0 13 10 9 13 1 10 9 2 13 1 10 9 0 11 11 11 7 11 11 11 2
36 1 10 11 11 3 4 4 1 13 9 1 10 10 11 7 1 11 11 2 16 3 13 1 10 9 1 11 16 10 9 13 1 10 9 0 2
49 11 11 2 3 13 1 2 11 2 2 10 9 16 13 1 10 9 7 10 9 3 1 10 9 1 10 9 2 13 1 10 9 0 16 4 13 1 10 9 2 9 16 13 10 9 1 10 9 2
54 1 10 9 1 11 11 11 2 10 9 1 9 15 4 13 1 11 1 11 11 1 10 9 1 12 7 16 4 13 1 9 1 11 11 2 11 13 1 10 9 15 9 1 9 1 9 1 11 11 2 13 9 11 2
32 15 13 1 9 0 1 10 9 0 0 7 13 3 1 10 9 0 1 10 9 1 9 0 13 1 10 9 1 10 9 0 2
29 10 9 13 10 9 1 10 0 9 1 9 0 1 10 9 0 1 10 11 2 16 15 13 1 9 7 15 13 2
76 10 9 1 12 1 10 9 0 11 1 11 2 15 13 10 9 13 1 10 9 11 11 7 11 11 1 11 1 10 9 13 1 11 2 9 1 9 7 9 2 1 10 9 1 12 9 1 10 9 13 2 13 15 10 9 0 1 12 9 2 1 10 9 1 13 15 15 4 13 10 9 1 11 3 0 2
43 15 13 1 10 9 1 9 0 7 0 2 16 3 13 0 1 10 9 8 7 16 3 13 1 10 9 1 10 0 9 0 2 16 15 13 15 1 15 1 10 0 9 2
43 3 15 1 15 2 3 11 2 11 7 11 2 13 10 9 3 0 1 9 0 2 16 3 11 2 11 2 11 7 11 13 1 10 9 1 10 9 3 0 1 9 11 2
22 1 10 11 11 11 7 10 9 1 10 11 2 10 9 15 13 1 11 11 11 11 2
25 15 13 1 9 0 1 9 1 9 11 11 7 11 2 13 1 9 1 10 9 2 13 10 9 2
13 3 1 10 9 10 9 1 9 0 13 10 9 2
71 13 1 10 11 0 1 10 9 0 1 10 9 0 1 9 0 2 1 10 9 1 11 7 1 10 9 1 11 2 15 13 1 10 11 1 10 9 11 1 10 9 1 10 9 1 10 11 7 9 1 10 9 0 15 13 1 10 9 1 10 9 0 1 10 15 13 9 10 9 11 2
25 10 12 9 0 4 13 1 11 7 1 10 11 11 2 1 3 10 9 11 13 0 1 10 9 2
10 10 9 4 13 1 2 11 11 2 2
15 1 11 13 10 15 11 2 11 2 2 9 0 1 11 2
13 3 13 1 12 9 16 15 13 1 10 15 2 2
21 1 15 15 13 1 10 9 0 2 11 9 7 11 9 2 7 13 2 13 2 2
20 13 16 13 9 16 3 4 13 10 9 2 7 10 9 4 13 1 10 9 2
29 1 10 0 9 13 1 10 9 15 13 10 9 1 13 10 9 13 1 11 2 7 13 10 9 1 10 9 12 2
6 10 9 1 10 9 2
15 1 12 2 11 15 13 1 11 1 13 1 10 9 0 2
12 3 10 11 15 13 3 16 3 10 9 13 2
45 1 12 2 15 13 1 10 0 9 1 13 9 1 10 9 0 1 11 7 1 12 4 13 9 1 11 11 1 10 11 11 11 11 11 2 16 13 10 9 1 10 9 1 11 2
17 3 13 1 10 9 13 10 9 0 2 13 1 9 0 7 0 2
23 10 9 1 9 1 10 9 1 10 12 1 11 1 12 15 13 1 10 9 1 10 9 2
24 13 10 9 1 13 10 9 1 11 11 1 10 9 2 13 10 9 0 1 13 1 10 9 2
44 10 9 4 13 1 13 1 10 9 1 15 1 10 12 9 2 1 10 9 1 10 9 2 10 9 0 4 13 15 1 9 7 3 4 4 13 1 10 9 1 10 9 0 2
21 11 11 2 11 11 1 9 2 13 10 9 1 9 1 9 0 13 1 11 11 2
47 10 9 0 1 11 11 2 11 11 2 13 10 9 1 13 1 10 11 11 2 3 1 10 11 13 1 13 1 10 0 9 2 10 11 11 11 2 2 15 1 10 0 9 1 11 2 2
20 11 11 13 10 9 2 11 10 11 11 11 2 1 10 9 1 10 0 9 2
49 10 9 0 11 11 13 10 9 0 7 1 9 1 11 2 2 11 2 2 13 1 2 11 2 11 11 7 11 11 11 2 2 12 2 2 7 13 3 1 9 0 1 2 11 2 2 12 2 2
22 10 9 4 3 13 1 10 9 1 11 2 15 1 10 9 0 1 10 9 1 11 2
18 10 9 1 10 9 1 10 9 13 10 9 1 10 9 7 10 9 2
5 12 9 1 9 2
70 11 11 12 3 13 10 9 1 10 9 0 1 10 9 1 9 1 9 1 9 11 11 2 11 11 11 13 11 11 11 11 11 11 12 2 11 11 2 10 9 13 1 8 13 1 11 11 13 1 11 11 12 2 15 4 13 3 0 1 10 9 0 1 16 13 1 11 1 12 2
62 0 16 13 9 1 10 9 1 10 9 7 9 2 7 15 3 13 16 13 0 2 7 3 0 2 13 15 16 10 10 9 1 9 13 1 10 11 2 0 9 1 9 2 0 9 2 0 9 1 9 2 13 0 1 13 1 10 0 9 1 9 2
51 1 10 9 1 11 2 10 9 13 1 2 11 11 11 2 11 2 7 11 11 11 2 11 2 2 3 0 1 10 10 9 0 2 13 1 9 0 1 2 9 2 9 1 9 2 9 2 9 7 9 2
16 10 9 13 0 2 0 9 0 2 2 1 12 1 0 9 2
62 15 3 13 10 2 9 2 0 1 10 9 0 13 10 9 0 1 10 9 7 9 1 9 0 2 11 11 2 16 15 13 2 0 2 1 16 10 0 9 0 1 10 11 15 2 13 1 10 9 0 7 1 10 9 1 9 1 10 10 9 2 2
51 0 2 3 13 9 16 13 10 9 0 3 2 16 3 13 10 9 2 3 2 3 9 13 10 9 1 10 9 11 1 10 9 7 1 10 9 0 1 10 9 2 16 13 10 9 1 10 9 1 9 2
51 1 11 1 12 11 11 2 9 1 10 9 1 11 11 1 10 11 1 11 11 2 13 1 11 1 9 1 10 11 11 11 2 11 11 11 2 2 7 10 9 10 11 13 1 2 9 0 7 0 2 2
22 1 10 0 9 13 10 9 2 1 10 16 2 1 13 2 13 1 10 9 1 9 2
21 1 11 2 10 9 13 15 3 9 1 10 9 2 13 1 10 12 9 1 9 2
11 2 3 13 3 1 10 9 7 10 9 2
21 2 10 11 7 10 11 4 13 9 0 2 2 4 13 10 9 2 11 11 11 2
26 3 10 9 1 9 4 13 1 10 10 9 2 1 9 15 3 15 4 13 9 1 10 0 9 0 2
29 13 3 10 9 2 7 2 1 10 9 1 16 9 9 13 3 0 2 13 10 9 1 10 9 0 11 7 11 2
12 3 1 0 3 15 4 13 1 10 9 0 2
20 3 0 2 15 13 1 11 7 15 13 3 4 13 1 10 9 1 10 9 2
26 10 9 2 9 11 2 4 13 10 9 1 10 9 1 11 13 10 11 2 16 13 1 12 7 12 2
8 2 16 15 15 13 1 11 2
7 13 10 9 7 13 15 2
35 1 10 9 1 11 11 2 11 11 2 10 9 1 11 11 2 10 9 1 11 11 7 1 10 11 0 2 11 13 10 0 9 1 9 2
16 10 9 13 10 9 9 2 16 10 9 3 13 13 10 9 2
23 13 10 9 7 10 9 1 10 0 9 1 9 1 10 9 1 11 7 11 13 3 13 2
43 8 2 11 11 13 10 9 1 10 9 0 1 11 11 2 13 1 10 9 1 10 9 2 1 10 9 1 11 11 11 1 3 3 1 10 9 1 10 9 1 10 9 2
19 11 11 13 10 9 1 9 0 1 10 9 11 1 10 9 1 10 11 2
8 13 10 9 9 5 7 1 8
33 13 1 10 9 2 10 9 7 9 13 1 10 0 9 0 1 10 1 10 9 1 10 0 7 0 9 1 9 0 7 9 0 2
47 11 11 2 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 0 16 15 13 1 9 0 7 1 10 9 1 10 11 11 1 10 11 1 11 7 1 10 9 1 9 1 11 2
18 1 15 15 13 10 9 1 10 9 7 10 9 0 1 10 9 0 2
19 10 9 1 9 13 10 9 11 11 2 2 10 9 3 0 1 10 9 2
21 10 9 0 15 13 1 10 9 1 9 2 1 10 9 2 10 11 7 10 11 2
39 10 10 9 1 15 0 0 4 13 1 9 3 0 7 1 9 3 0 2 16 10 9 4 13 9 13 1 2 9 2 2 2 9 2 7 2 9 2 2
31 10 12 1 11 2 1 11 2 15 13 2 0 1 11 2 1 10 10 9 1 12 9 2 1 10 9 1 10 9 11 2
32 15 13 16 1 10 13 1 10 9 9 1 10 11 11 2 0 1 10 11 11 2 15 4 13 1 10 11 2 3 13 9 2
35 1 0 2 3 1 12 9 1 9 1 10 9 2 11 11 2 15 4 13 1 9 1 10 12 1 9 1 10 0 9 1 10 0 9 2
31 10 9 1 10 11 3 13 10 9 0 1 12 9 2 10 8 8 0 7 10 9 1 9 1 11 11 2 1 10 9 2
17 10 11 1 11 4 13 10 9 0 7 1 9 1 10 0 9 2
16 3 1 10 12 5 1 10 9 13 1 10 9 1 9 0 2
50 10 9 13 10 9 0 0 0 1 10 9 0 1 11 1 16 4 13 1 12 2 15 3 4 4 13 1 9 0 1 10 9 7 9 1 9 0 1 9 0 2 13 1 10 9 2 1 0 9 2
10 13 9 2 9 2 9 7 9 0 2
22 11 15 13 2 7 13 13 15 2 16 13 13 10 9 0 2 7 13 13 1 11 2
20 10 9 1 10 11 11 4 13 1 9 7 10 9 0 13 3 0 1 9 2
19 10 9 11 2 11 11 2 11 2 11 7 11 13 10 9 1 10 11 2
33 10 9 15 13 1 11 1 12 1 10 9 1 10 9 1 10 9 1 11 11 2 11 2 11 10 11 2 2 13 1 11 11 2
37 11 3 13 10 9 1 10 9 1 11 1 13 10 9 1 11 11 1 10 11 2 7 15 13 3 13 1 10 11 11 1 12 1 11 1 12 2
32 11 11 15 13 1 10 0 9 1 9 1 15 9 1 10 9 0 7 16 13 1 12 1 12 9 1 10 9 1 10 9 2
32 3 2 13 10 0 9 1 9 1 0 9 16 15 13 1 13 10 9 2 7 9 1 9 2 2 13 1 10 9 1 9 2
20 13 1 9 10 9 0 1 11 2 13 9 0 1 10 9 1 12 1 12 2
14 1 15 11 11 13 13 1 10 9 0 1 10 9 2
16 13 1 15 16 10 9 1 10 9 1 9 15 13 10 9 2
23 10 9 1 10 9 13 3 0 2 13 1 9 2 9 7 10 9 13 13 1 0 9 2
18 10 9 13 10 9 1 10 9 7 16 3 15 13 1 10 9 0 2
16 11 11 2 5 2 13 10 9 0 16 13 10 9 0 11 2
8 9 0 0 2 8 12 2 2
13 10 9 13 10 0 9 1 13 1 11 1 12 2
28 4 13 3 0 1 10 9 0 1 11 13 10 9 0 1 10 9 10 9 1 10 0 9 16 15 13 0 2
43 15 1 15 16 15 13 13 2 1 10 9 2 0 16 13 9 1 9 16 3 3 3 13 1 0 9 1 10 12 11 7 11 12 2 16 15 4 13 10 15 1 9 2
13 1 12 1 12 13 9 2 9 1 10 9 0 2
32 1 9 1 11 1 10 9 0 2 11 11 13 3 1 12 9 2 16 13 3 9 1 10 9 0 2 7 3 13 10 9 2
42 1 9 3 0 7 10 0 9 1 9 2 10 9 4 13 1 10 9 1 13 9 1 10 9 2 7 13 1 10 9 3 10 9 15 13 2 2 1 15 13 0 2
32 3 13 13 1 9 1 11 1 10 9 1 10 9 1 10 9 1 9 0 11 11 13 1 13 1 10 9 1 12 11 11 2
11 1 13 1 10 9 10 9 3 13 0 2
15 13 9 1 10 9 11 11 2 3 3 13 1 10 9 2
47 13 10 9 15 1 9 0 7 1 10 9 2 13 1 15 10 9 1 10 9 1 10 9 1 9 2 13 10 9 13 1 10 9 1 9 7 9 1 10 9 1 13 10 9 1 9 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
13 13 10 9 1 10 9 3 1 13 15 1 15 2
37 10 9 0 2 3 1 10 11 1 11 2 10 11 2 13 10 9 1 10 9 0 1 10 9 1 13 1 10 9 1 10 9 0 1 10 9 2
28 13 1 9 3 0 16 13 1 15 1 10 9 1 10 0 9 0 13 15 10 9 16 3 13 9 1 9 2
69 10 9 1 10 9 13 1 13 10 9 0 1 10 11 2 10 9 1 10 9 0 3 0 1 10 9 0 1 10 9 2 10 9 16 15 13 3 1 10 9 0 2 2 0 2 2 1 13 1 13 10 9 3 0 1 10 0 9 16 4 13 1 10 11 1 10 9 0 2
6 10 9 13 15 0 2
17 1 10 12 9 1 9 13 3 1 11 2 13 1 10 0 9 2
20 10 9 11 7 11 13 1 12 9 0 7 12 2 12 1 10 9 2 9 2
31 13 10 9 13 9 1 9 1 9 2 7 1 13 10 9 15 13 1 10 9 7 13 15 16 0 9 15 13 1 9 2
22 10 9 1 9 4 13 13 3 9 1 9 16 13 10 9 1 9 0 9 1 9 2
38 13 1 10 0 9 5 8 10 12 9 5 8 16 12 1 10 0 9 15 13 10 9 1 12 9 3 9 1 10 9 2 1 13 10 0 12 9 2
20 10 0 9 1 11 11 1 13 15 10 9 1 10 9 0 1 10 0 9 2
13 3 15 13 1 13 10 9 11 1 10 9 11 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
20 10 9 13 1 9 1 9 0 7 15 4 13 9 1 9 1 10 9 11 2
38 10 9 1 10 9 15 13 1 0 9 1 11 1 9 1 10 9 2 11 2 1 12 2 10 9 3 1 10 9 1 10 9 0 2 11 11 2 2
50 13 1 10 9 13 1 10 9 1 9 1 10 11 2 10 11 2 11 12 7 11 2 11 7 2 3 3 2 1 12 2 15 13 1 9 0 2 13 9 1 9 1 9 1 11 11 7 11 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 8 2
39 10 9 13 1 10 9 1 10 9 0 2 1 10 9 1 10 9 10 9 2 16 1 10 9 0 1 10 9 15 4 4 13 1 10 9 1 10 9 2
9 10 9 13 0 2 0 7 0 2
8 10 9 13 13 15 1 11 2
17 1 10 9 2 11 13 16 11 15 13 3 1 15 1 10 9 2
15 11 11 13 10 9 1 11 2 13 10 9 12 1 11 2
36 3 4 13 10 9 1 13 10 9 2 7 3 15 4 13 0 1 13 10 9 1 10 9 2 15 7 15 13 7 3 13 15 13 10 9 2
30 10 9 0 13 0 7 13 10 9 2 10 9 2 10 9 0 2 9 0 2 10 9 2 9 0 7 10 9 0 2
20 1 10 9 15 13 10 9 0 2 1 9 2 13 7 3 1 10 0 9 2
26 10 12 9 13 1 10 0 0 9 1 10 11 1 11 2 11 2 2 10 9 13 0 1 10 11 2
30 1 10 9 13 10 0 9 0 2 1 9 0 2 16 13 0 9 1 10 9 0 1 10 9 7 10 9 1 9 2
14 10 11 13 3 10 9 2 7 10 9 3 4 13 2
37 10 9 1 10 9 1 10 9 2 13 1 10 9 1 9 1 10 9 2 4 13 10 9 1 10 9 2 1 9 1 10 9 7 10 9 0 2
23 13 12 9 1 9 2 0 2 0 2 0 7 12 9 1 9 16 15 13 1 10 9 2
15 9 1 10 9 11 1 10 11 1 10 11 11 1 11 2
23 9 1 16 10 9 13 1 10 0 9 1 9 1 10 9 1 9 1 12 9 1 9 2
16 1 10 9 2 10 9 13 10 9 7 10 9 1 10 9 2
6 15 15 4 13 1 8
34 15 1 15 13 10 9 0 11 11 16 15 13 1 11 7 16 13 9 2 10 9 13 10 11 16 15 13 1 10 9 1 10 9 2
6 11 11 13 10 9 0
32 13 10 9 1 11 2 9 1 9 2 11 2 11 11 2 11 7 11 2 7 10 9 1 11 11 2 9 1 11 7 11 2
21 13 1 10 9 1 10 9 1 10 15 15 13 2 10 9 13 0 1 12 9 2
23 10 9 2 13 1 10 9 0 0 2 13 1 10 9 10 9 1 10 9 11 11 11 2
21 3 13 9 1 4 13 15 1 9 1 15 2 15 3 15 13 13 10 0 9 2
18 11 13 10 9 8 1 10 9 11 0 1 10 9 1 10 9 11 2
8 1 10 9 2 11 13 3 2
15 1 10 9 2 11 13 9 11 1 9 2 3 1 9 2
13 10 0 9 1 10 9 13 1 10 9 1 12 2
12 10 12 1 11 1 12 10 9 13 11 3 2
52 10 9 13 12 9 15 3 0 1 10 9 1 10 9 13 10 9 1 10 9 7 1 9 0 7 15 1 10 15 15 13 1 10 9 1 10 9 1 10 9 12 1 10 9 1 10 9 1 10 9 0 2
33 3 1 13 15 1 10 11 11 11 11 2 11 13 1 9 1 12 1 10 9 11 11 2 13 1 10 9 13 3 1 11 11 2
17 15 13 10 9 1 9 1 10 9 1 10 9 2 3 3 3 2
23 10 9 1 10 9 8 11 11 4 13 1 13 1 10 9 0 1 16 13 1 10 9 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
25 10 9 13 1 10 9 0 1 10 11 2 13 15 1 10 9 1 9 2 9 7 9 1 9 2
35 13 1 10 9 2 1 10 9 1 10 9 13 2 10 9 0 1 4 13 10 9 13 1 5 12 1 9 1 12 1 5 12 1 12 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
7 13 12 9 1 9 0 2
39 3 13 10 9 1 10 9 16 2 1 10 9 1 10 9 2 15 13 1 15 1 10 3 0 7 0 1 10 9 0 1 11 7 10 9 0 1 9 2
36 10 9 1 9 2 13 1 10 9 1 9 1 10 11 2 13 10 9 2 10 9 7 10 9 1 10 11 2 0 1 10 9 0 1 9 2
57 11 15 13 10 0 9 1 10 9 0 1 13 10 0 9 1 10 9 0 1 11 2 1 15 15 11 15 13 2 1 10 9 1 10 0 11 2 2 13 1 9 1 10 9 2 7 15 3 4 13 1 10 9 1 13 2 2
4 11 11 11 2
27 10 9 1 9 13 0 1 10 9 7 10 9 1 10 9 0 7 0 7 13 1 9 10 9 1 9 2
7 13 10 9 1 9 0 2
16 10 11 11 1 10 12 13 12 9 0 0 2 13 0 9 2
9 2 10 9 3 13 1 10 9 2
34 10 9 15 13 1 12 7 10 9 3 13 10 9 1 10 11 1 4 1 13 10 9 3 13 2 3 1 11 2 1 10 9 0 2
20 13 1 9 7 10 9 0 13 10 11 11 1 10 11 11 11 1 11 11 2
83 9 7 9 0 1 11 2 13 10 9 0 1 10 9 2 16 15 13 1 10 9 1 16 9 0 0 13 10 9 0 16 13 10 9 0 13 13 10 9 1 10 9 0 15 13 10 9 0 2 1 9 1 10 9 1 13 10 9 0 16 15 13 2 3 13 10 9 1 10 9 2 10 8 2 9 2 9 2 9 2 9 0 2
24 1 10 9 1 9 16 13 9 2 10 9 9 13 1 10 9 7 15 13 1 10 9 0 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
45 1 10 9 13 10 9 1 13 9 1 11 2 1 10 9 1 10 15 11 13 10 9 1 15 2 2 16 13 10 9 9 1 10 13 10 9 7 15 13 1 10 9 1 9 2
31 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 9 12 2 7 10 9 0 1 9 13 9 12 2
54 1 10 9 0 13 1 9 1 10 9 1 9 13 11 11 2 11 2 12 2 2 12 2 7 3 3 9 1 10 9 1 11 1 11 7 11 2 3 7 9 1 9 9 0 1 10 11 1 11 3 1 10 11 2
23 10 9 1 13 10 9 0 0 4 13 3 3 10 9 2 1 15 15 15 13 0 9 2
31 10 9 2 1 10 9 2 11 2 13 1 10 9 10 9 0 16 15 13 10 9 1 10 9 1 9 1 10 9 12 2
29 10 9 0 2 4 4 13 10 11 11 11 12 1 12 8 2 13 1 9 9 2 15 4 4 13 1 10 9 2
30 1 12 2 11 4 1 13 1 9 0 1 10 9 1 10 11 11 7 1 9 11 13 7 4 1 13 1 12 9 2
4 10 9 13 2
11 10 9 15 13 1 11 2 11 7 11 2
44 1 10 9 0 1 10 9 1 9 0 9 1 10 9 1 10 9 1 9 10 9 1 9 0 13 10 9 0 1 10 9 1 9 1 9 1 10 9 1 10 9 1 9 2
16 10 9 1 11 2 1 9 0 2 15 13 3 1 10 9 2
32 1 10 9 10 9 11 2 11 11 13 1 9 11 2 12 2 13 3 1 15 1 10 9 1 10 9 7 10 10 9 0 2
17 2 11 2 13 7 13 13 2 9 2 9 7 9 1 11 2 2
7 11 11 4 13 10 9 2
12 10 0 9 1 11 1 13 9 1 10 9 2
8 13 0 9 1 10 0 9 2
44 1 10 9 2 15 1 10 9 7 9 16 13 10 11 13 0 9 1 10 9 2 13 3 9 1 10 9 2 9 1 10 9 7 9 0 1 11 2 2 7 10 9 0 2
29 10 9 0 7 0 2 3 3 15 13 10 9 0 2 7 3 15 13 1 10 9 1 10 9 16 13 13 9 2
27 1 11 1 12 2 15 13 1 10 9 1 9 1 10 11 1 11 2 7 11 11 4 13 1 10 9 2
29 13 10 9 2 3 15 1 9 0 2 10 9 1 9 0 13 9 2 7 13 0 9 1 10 9 7 10 9 2
7 15 4 13 10 9 0 2
45 10 9 0 13 10 2 9 1 9 0 2 1 11 1 10 9 1 10 9 0 7 10 2 0 9 2 16 13 1 9 1 10 9 0 1 9 1 11 2 8 2 2 1 11 2
16 10 0 9 3 13 1 15 7 1 10 0 9 2 15 13 2
20 10 9 13 3 10 9 0 1 10 9 0 2 3 3 15 13 10 9 0 2
28 10 9 13 1 9 0 2 13 3 1 10 9 10 9 1 10 11 1 11 2 13 1 10 9 1 10 9 2
26 3 13 0 10 9 0 1 10 11 11 2 7 9 1 10 9 2 7 10 9 1 10 11 1 11 2
18 0 2 10 9 13 0 2 3 1 10 11 1 10 11 7 10 11 2
26 3 2 1 12 10 0 11 1 10 9 13 9 1 11 2 4 13 9 1 10 9 16 8 10 9 2
34 1 9 1 10 9 1 10 9 2 10 11 13 1 10 9 1 13 1 10 11 11 1 8 0 1 10 0 9 1 10 9 11 11 2
35 1 9 1 10 9 13 1 13 3 10 9 7 3 13 10 9 10 11 1 11 2 1 10 15 13 10 0 9 1 10 9 2 12 2 2
33 11 1 10 11 2 9 7 1 9 0 2 13 10 9 1 10 9 1 11 1 11 1 11 2 16 15 4 13 1 9 10 9 2
30 3 1 10 9 2 9 11 11 13 2 11 2 10 9 3 0 1 10 15 11 13 10 9 0 7 11 13 10 9 2
62 1 3 16 1 10 9 4 13 15 10 9 0 1 10 12 1 11 1 12 1 10 9 0 0 7 0 12 9 13 1 10 0 9 7 1 9 9 0 2 9 7 9 2 9 0 2 9 1 9 0 2 9 7 10 9 1 9 0 1 12 9 2
26 10 9 11 11 13 10 9 0 1 9 0 7 9 1 9 1 9 0 1 9 7 1 9 7 9 2
18 10 9 1 10 9 13 1 10 9 1 12 1 12 9 7 12 9 2
33 10 9 13 1 10 9 16 13 10 11 11 1 11 7 16 15 13 9 9 1 10 9 13 1 10 11 11 1 11 2 11 2 2
49 3 2 11 13 0 1 10 9 1 9 1 2 9 1 10 9 2 2 10 12 5 1 9 7 13 1 9 2 7 2 10 11 11 2 2 10 8 2 8 2 0 9 0 1 10 9 0 11 2
11 4 13 1 9 10 12 1 11 1 12 2
6 2 15 13 10 9 2
50 2 10 9 1 10 9 1 9 0 7 8 2 8 2 1 10 9 1 9 2 13 0 1 10 9 16 15 13 1 9 1 12 9 2 9 1 10 16 2 15 13 2 3 3 13 9 1 10 9 2
16 3 0 10 11 11 11 13 0 9 1 10 9 1 9 0 2
15 15 13 16 13 1 10 9 0 3 0 1 10 9 0 2
42 13 1 9 1 9 1 11 1 12 2 13 1 10 9 1 11 1 11 2 7 2 1 9 2 16 13 10 9 1 9 1 11 2 13 1 9 10 12 1 11 12 2
41 11 4 13 1 10 9 2 2 3 13 15 1 10 9 1 11 7 1 10 9 2 16 3 4 13 1 15 1 10 9 1 10 9 0 7 10 1 10 9 2 2
12 15 13 10 9 1 12 9 13 1 10 9 2
8 1 9 13 1 9 1 9 2
32 11 11 13 1 12 10 9 1 9 0 1 11 1 11 16 10 9 2 1 10 9 1 10 9 0 11 11 2 13 10 9 2
32 3 11 13 9 1 10 11 11 1 10 11 1 11 2 3 11 11 1 11 1 10 11 2 10 15 13 1 10 9 1 12 2
39 15 1 10 9 2 1 12 8 2 13 10 9 0 0 7 0 7 15 13 1 9 1 10 9 9 12 2 7 10 9 4 13 0 7 10 9 3 13 2
43 1 10 9 15 13 1 9 0 2 1 10 0 9 1 13 10 9 1 10 9 0 15 15 4 1 13 1 9 1 9 7 9 1 10 3 4 13 1 9 3 3 13 2
15 1 10 9 11 11 13 10 9 1 10 9 1 12 2 2
21 15 13 1 11 2 11 2 11 2 11 2 11 7 10 9 1 11 2 11 2 2
14 15 13 12 9 1 10 9 7 10 9 1 12 9 2
10 13 10 9 1 9 7 1 9 0 2
27 15 15 13 1 0 9 9 1 10 0 9 2 1 0 9 0 7 1 9 0 16 3 13 1 13 0 2
43 10 9 4 13 1 11 11 11 8 2 10 9 13 10 9 11 11 11 2 10 9 8 1 12 9 1 10 9 8 8 12 9 2 9 9 0 2 9 11 12 7 8 2
29 10 9 1 10 9 15 13 1 10 9 0 8 2 16 13 2 0 2 2 7 8 2 16 13 2 0 9 2 2
20 1 10 9 15 13 10 9 9 2 10 9 1 10 9 2 11 1 11 2 2
20 11 13 7 4 13 1 11 7 11 16 15 13 15 1 10 9 1 10 9 2
34 10 9 1 9 0 2 3 13 11 2 3 13 10 9 1 12 9 1 9 0 2 15 16 13 10 12 5 1 10 9 1 10 9 2
27 1 10 9 1 11 11 16 13 10 9 1 10 11 1 11 1 12 15 4 13 15 1 10 9 1 11 2
39 10 9 2 10 0 9 13 11 10 11 2 13 3 12 9 7 3 13 1 10 9 1 11 1 10 9 13 1 9 1 10 9 1 9 0 1 10 9 2
11 1 10 9 15 13 10 0 9 1 11 2
27 11 11 3 13 10 9 0 1 11 7 11 2 7 15 3 13 13 16 3 13 9 7 9 1 10 9 2
14 1 9 1 0 9 2 10 9 13 10 9 11 12 2
51 11 7 11 2 10 9 1 10 9 2 2 16 13 15 1 10 9 13 1 11 1 10 12 9 13 2 4 13 1 10 0 1 10 9 0 16 0 1 10 1 10 9 13 1 13 15 1 10 9 0 2
4 13 1 11 2
12 1 11 2 3 15 13 10 9 1 10 9 2
22 10 9 7 15 4 1 13 1 10 9 7 13 1 2 16 15 13 2 10 9 2 2
9 10 9 15 13 1 9 1 13 2
51 1 10 9 0 12 7 12 2 10 9 0 1 9 0 13 1 10 9 1 10 9 2 13 10 9 1 9 0 7 0 9 1 9 1 9 2 13 1 10 12 5 1 10 9 0 9 1 10 11 11 2
14 9 1 9 2 1 3 0 9 2 3 0 7 0 2
21 13 10 9 1 10 9 2 3 13 3 7 13 10 9 1 13 10 9 1 9 2
21 13 10 9 1 9 1 9 2 10 9 4 13 3 12 9 0 3 1 10 9 2
12 10 11 13 10 9 7 13 9 1 10 9 2
35 10 11 2 12 4 13 1 10 9 3 1 16 11 11 4 4 13 7 13 1 12 13 1 13 3 10 9 1 10 9 11 11 2 12 2
16 1 9 13 11 2 7 1 9 2 11 7 11 13 1 11 2
12 3 13 0 13 15 13 9 0 7 9 0 2
31 10 9 1 10 9 3 4 4 13 1 9 0 7 9 1 10 9 2 1 11 11 7 11 11 1 10 9 3 1 9 2
35 1 10 9 1 9 0 15 15 13 1 10 9 0 1 10 9 2 7 10 9 3 4 13 1 10 9 1 12 5 1 10 9 1 9 2
14 11 11 13 1 13 10 9 10 9 1 10 11 11 2
13 1 13 1 12 15 13 3 7 1 10 0 9 2
43 1 10 9 1 10 9 1 10 11 11 2 11 11 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 13 1 9 0 7 2 12 5 2 12 5 5 13 9 2
18 1 10 10 9 1 9 16 4 13 1 11 15 4 1 13 1 15 2
15 1 15 13 10 9 12 16 13 10 11 11 7 10 9 2
36 10 9 13 13 1 13 10 9 1 10 9 16 10 9 4 13 1 10 9 7 2 1 15 2 13 10 9 1 10 9 16 3 13 10 9 2
39 10 0 9 13 9 0 0 2 1 0 12 2 10 12 9 7 13 1 10 9 1 10 9 2 15 13 13 10 12 9 0 1 10 9 13 9 1 9 2
26 1 10 9 2 10 9 1 9 0 13 10 0 9 1 10 11 2 13 15 1 10 9 7 10 9 2
41 1 10 12 1 10 9 2 10 9 1 10 9 0 0 1 9 13 1 10 9 1 10 9 2 13 1 9 1 9 10 9 7 9 1 10 10 9 1 9 0 2
18 1 12 15 13 10 9 1 0 9 13 11 1 11 2 2 12 2 2
20 13 3 0 10 9 1 9 0 1 9 0 2 1 1 8 2 8 7 8 2
36 1 10 12 1 11 1 12 7 10 12 1 11 1 12 13 1 9 0 1 10 9 1 11 11 2 7 16 11 11 1 11 13 1 10 9 2
37 10 9 13 3 0 1 10 9 1 10 9 2 1 10 9 3 0 1 10 9 1 11 7 1 10 9 0 1 10 9 1 11 11 7 11 11 2
29 15 13 16 11 3 13 1 10 9 16 13 9 2 0 2 1 0 9 1 9 2 1 10 9 1 10 9 0 2
13 10 0 9 1 10 9 13 0 2 12 5 2 2
3 2 9 2
31 10 0 9 13 10 12 1 11 1 12 2 16 11 4 13 1 10 9 11 16 13 10 9 16 13 10 9 1 9 0 2
25 16 13 1 10 11 1 9 1 9 2 13 10 9 2 9 1 11 1 16 15 13 1 10 11 2
16 1 12 2 13 10 9 1 10 0 9 1 10 9 1 11 2
6 11 11 11 2 8 2
29 10 11 2 11 3 13 10 9 1 10 9 1 9 2 3 1 0 9 0 1 9 7 9 1 9 0 10 9 2
70 10 9 1 9 1 10 11 11 13 16 15 13 4 4 1 13 10 2 11 11 2 2 16 13 13 9 3 3 1 10 9 0 1 9 0 2 2 1 10 9 3 15 13 9 7 10 9 0 1 9 4 13 1 10 9 1 10 9 2 13 16 10 11 1 10 9 13 1 11 2
51 1 10 9 1 10 9 0 7 10 9 2 11 4 3 13 13 12 9 1 13 1 10 9 10 9 1 10 9 0 7 13 1 9 1 10 9 1 11 2 16 13 10 9 1 9 1 10 11 11 11 2
17 1 12 4 13 10 9 1 9 1 11 11 1 10 9 0 0 2
40 13 10 0 9 16 15 1 10 9 1 10 16 4 13 15 13 16 4 13 10 9 3 0 16 7 3 3 13 1 11 2 1 10 9 1 13 10 15 3 2
30 10 9 7 9 1 10 11 4 13 1 15 7 10 9 0 2 3 16 10 9 1 10 11 3 4 13 1 3 0 2
18 10 9 13 3 0 1 10 9 9 7 13 10 9 1 10 9 9 2
26 0 2 13 1 9 7 3 15 4 1 13 2 13 13 1 9 7 3 13 9 1 13 1 10 9 2
25 10 9 13 1 10 11 2 11 1 11 11 2 1 12 2 1 10 0 9 13 1 10 9 0 2
15 1 12 9 1 9 2 13 1 10 9 1 9 2 9 2
10 13 10 9 1 11 2 2 1 13 2
53 1 10 9 0 13 10 9 1 9 1 0 9 2 1 10 15 13 10 11 1 10 11 2 16 15 13 1 10 11 1 11 2 2 3 13 13 0 9 1 9 1 9 0 2 13 10 0 9 0 1 9 0 2
15 10 9 3 15 13 2 7 11 15 13 3 13 1 9 2
24 13 0 1 10 9 0 1 11 11 2 1 10 9 11 2 9 1 10 9 0 1 11 2 2
18 10 9 0 4 13 1 10 9 1 10 9 16 13 9 1 10 9 2
11 13 12 9 16 3 4 13 1 10 9 2
37 1 11 1 12 2 10 11 1 11 1 11 11 13 10 11 11 11 11 11 10 15 15 13 1 10 9 0 1 11 11 2 10 9 1 10 11 2
32 1 12 2 11 13 1 10 9 2 11 11 11 2 11 2 2 1 11 8 11 11 2 1 10 9 2 2 11 11 11 2 2
50 1 10 0 9 13 9 1 0 9 1 9 7 15 13 10 9 0 7 10 9 2 7 1 10 9 15 13 10 9 2 10 9 0 7 10 9 7 13 9 3 2 0 2 0 2 0 2 8 2 2
28 15 1 10 9 13 9 1 9 2 9 2 1 9 1 9 2 7 13 15 15 13 1 10 9 1 10 9 2
17 10 9 13 12 9 2 7 13 1 10 9 0 1 10 11 11 2
15 10 9 0 13 1 12 9 1 9 0 2 8 5 2 2
42 10 9 13 1 10 9 13 10 9 1 12 9 2 10 9 1 11 11 2 11 2 7 11 11 2 11 2 13 10 0 9 1 12 9 2 11 2 11 2 12 2 2
74 3 13 15 1 10 9 1 10 9 2 13 3 16 13 10 9 1 10 9 7 10 9 1 10 13 9 2 1 10 9 1 10 9 7 10 9 15 4 13 1 10 9 2 1 10 15 13 15 15 13 10 9 16 10 9 13 0 1 10 9 2 7 7 3 10 9 13 15 4 13 1 10 9 2
47 2 10 9 16 13 13 1 10 9 0 7 13 10 9 3 0 15 1 10 11 7 1 10 9 2 7 15 13 10 11 2 10 11 7 10 11 7 15 4 13 10 9 2 2 13 11 2
24 7 2 3 1 10 15 2 13 10 10 9 16 3 13 0 7 16 13 10 9 0 7 0 2
14 11 13 1 10 9 1 10 9 13 1 10 0 11 2
23 13 0 9 1 13 10 11 2 15 1 10 9 0 2 13 9 1 10 9 1 0 9 2
11 10 9 1 11 15 13 13 1 10 9 2
8 11 15 13 0 1 10 9 2
24 13 1 10 9 1 10 9 1 11 11 1 10 9 1 11 2 13 3 1 10 9 1 11 2
19 15 13 1 12 9 1 9 0 1 10 9 1 11 2 9 1 10 9 2
12 13 9 11 2 15 7 10 9 3 15 13 2
40 1 15 15 4 13 16 10 9 13 10 9 0 2 2 1 10 9 2 0 2 2 1 10 9 1 9 7 1 10 9 2 7 13 1 10 9 1 10 9 2
22 10 9 0 2 13 3 10 9 0 2 9 1 10 9 1 9 7 9 1 10 9 2
38 10 9 2 16 13 9 1 10 11 11 11 1 10 9 1 11 11 10 12 1 11 1 12 2 13 1 10 9 1 11 11 7 1 10 11 11 11 2
41 10 11 11 1 10 9 0 13 12 9 2 12 1 12 2 1 10 12 12 12 9 16 10 9 1 9 0 9 13 12 9 2 12 1 12 2 1 10 12 9 2
9 1 10 9 0 13 10 0 9 2
41 10 9 0 13 1 10 9 1 11 13 1 15 2 3 1 10 9 0 1 11 7 10 9 1 10 11 11 2 11 2 10 9 0 7 9 1 10 11 11 2 2
28 10 9 16 15 13 13 10 9 11 2 15 13 3 13 9 1 10 9 7 13 16 15 15 13 1 10 9 2
26 10 9 0 13 0 2 0 2 0 7 0 2 8 8 8 9 2 0 2 0 2 0 0 1 0 2
35 15 15 13 1 10 0 9 0 0 2 12 2 2 7 13 1 10 9 0 1 10 9 0 2 13 1 10 11 11 2 7 10 11 11 2
55 1 10 9 1 0 9 2 3 1 11 2 13 12 1 10 9 2 11 2 11 2 11 2 11 10 11 2 11 10 11 2 11 7 11 2 2 3 1 10 9 7 10 0 9 1 10 9 1 9 2 9 7 9 0 2
22 11 13 1 10 9 0 13 1 11 2 11 2 11 11 2 3 11 2 11 11 2 2
19 11 11 2 10 9 1 2 11 11 11 2 2 4 13 1 13 10 9 2
56 10 9 2 13 1 12 2 13 2 15 1 10 9 16 10 9 13 1 10 9 2 2 1 11 2 15 13 10 9 1 10 9 1 10 16 15 13 10 9 1 10 9 11 11 2 8 2 2 15 13 2 0 2 1 11 2
55 10 9 1 11 4 13 1 9 1 9 9 2 16 3 13 9 0 2 1 9 1 10 11 1 11 7 11 2 1 9 1 11 2 11 2 7 11 2 11 2 2 7 1 10 9 1 10 11 11 1 11 2 11 2 2
6 13 12 9 1 12 2
7 15 13 13 0 1 11 2
7 10 9 15 13 3 3 2
10 13 1 10 9 1 10 11 11 11 2
55 1 10 9 11 7 10 9 9 2 11 7 11 13 16 15 1 10 15 13 1 10 9 13 9 1 10 9 16 15 13 0 2 7 13 1 10 9 2 16 15 13 15 0 13 16 10 9 4 13 1 9 1 10 9 2
20 10 12 9 3 13 10 9 1 9 1 9 0 1 10 9 13 11 11 11 2
12 10 0 9 1 10 9 15 13 1 9 0 2
32 10 11 11 2 11 2 12 2 13 10 9 2 0 1 10 9 0 1 10 11 11 2 16 3 13 10 9 1 9 1 9 2
21 3 7 15 1 10 9 7 10 9 3 2 1 10 9 2 10 9 13 10 9 2
44 11 11 11 2 8 12 1 11 1 12 2 2 13 10 9 0 1 9 0 2 0 2 16 3 1 10 9 2 9 1 10 11 11 2 13 15 1 10 0 9 1 10 9 2
40 1 12 13 1 13 9 1 9 2 7 1 12 10 9 15 13 1 9 1 9 2 13 1 10 11 1 10 11 2 15 1 9 0 15 4 7 13 1 12 2
9 4 13 10 12 1 11 1 12 2
9 10 9 1 9 13 0 12 9 2
28 1 10 9 2 10 9 13 1 9 10 9 0 7 3 10 9 0 16 13 1 13 3 10 9 1 9 0 2
27 10 9 1 10 9 15 4 13 1 12 1 10 12 9 1 10 9 2 15 4 4 4 13 1 10 9 2
36 0 9 0 1 10 0 9 0 2 4 13 1 9 7 9 1 9 0 3 10 0 9 13 10 9 1 10 2 9 2 16 1 15 15 13 2
76 1 10 9 2 10 9 11 11 2 1 10 0 11 1 11 2 2 3 4 13 10 12 1 11 1 12 16 10 9 4 4 13 1 9 1 10 9 9 0 11 1 10 9 7 10 9 1 0 9 0 1 10 3 2 13 10 9 7 16 10 9 7 10 9 13 3 13 10 9 1 9 0 1 9 0 2
17 3 16 13 1 9 7 1 9 2 15 3 0 2 3 10 9 2
10 10 9 0 0 13 10 9 0 0 2
25 15 13 9 1 10 9 1 10 9 1 10 9 1 11 1 10 11 1 10 9 1 11 1 12 2
36 10 9 3 13 9 5 12 1 9 0 2 1 15 15 13 10 0 9 3 0 1 12 2 7 15 1 10 10 9 9 1 11 1 10 9 2
47 15 13 1 10 9 7 15 15 13 2 7 3 11 13 1 11 11 1 10 9 1 10 9 0 1 9 1 9 2 13 15 3 0 2 11 13 9 7 9 1 10 9 7 13 10 9 2
18 11 3 13 10 9 1 10 9 0 7 13 1 10 9 1 10 9 2
17 10 9 3 2 10 9 1 10 9 13 16 10 9 13 3 0 2
20 13 10 9 1 16 10 9 1 10 16 3 13 13 2 3 2 1 9 0 2
25 10 9 9 3 13 3 0 1 16 0 2 3 1 0 9 2 16 9 7 9 13 10 0 9 2
20 1 9 2 1 10 9 1 9 3 13 0 13 9 0 1 9 1 12 8 2
5 13 9 1 11 2
47 10 9 13 10 9 1 12 5 5 2 1 10 9 12 5 5 4 13 1 9 2 7 10 9 1 12 9 2 1 10 9 1 9 1 12 8 2 5 5 2 1 9 0 1 12 2 2
10 11 11 13 10 9 7 13 10 9 2
18 10 9 0 1 10 9 0 13 2 2 1 2 10 9 7 10 9 2
31 10 9 0 1 10 9 13 1 12 5 0 2 12 5 0 0 2 12 5 1 10 9 7 12 5 1 12 7 3 9 2
29 10 0 11 11 11 4 13 1 10 9 12 1 10 11 11 1 11 2 1 10 0 11 1 10 11 1 10 9 2
16 11 0 13 10 9 1 9 1 10 9 11 1 10 9 11 2
20 10 9 12 1 11 1 12 15 13 10 0 9 1 9 1 10 9 1 9 2
48 1 10 9 1 10 9 1 11 2 10 9 13 0 9 16 13 10 9 1 11 2 15 13 9 7 9 0 7 16 15 13 13 1 10 9 1 9 2 13 0 7 13 15 9 1 10 9 2
28 10 9 13 10 9 1 9 1 9 1 10 9 0 16 13 10 9 0 1 9 0 13 10 9 0 1 9 2
45 1 9 1 9 2 10 9 13 1 10 10 9 1 10 9 0 1 13 10 9 0 1 10 9 3 4 0 2 9 0 1 9 2 9 1 9 2 9 1 10 9 7 10 9 2
37 1 12 9 13 1 9 0 1 10 9 1 12 9 15 4 4 13 16 13 9 2 3 12 9 4 13 1 10 9 1 12 5 1 10 9 0 2
21 15 13 1 10 9 1 10 9 11 2 3 13 1 10 10 9 1 10 9 0 2
40 10 9 0 1 10 0 9 1 11 13 10 11 10 0 9 1 9 1 10 9 0 9 1 11 2 1 10 9 1 15 1 10 9 8 1 10 11 11 12 2
24 1 10 9 0 1 11 2 10 11 13 1 10 9 1 9 1 13 13 10 9 1 10 9 2
11 10 9 13 10 9 0 1 0 9 0 2
28 10 9 7 9 11 11 13 16 13 2 11 11 11 11 11 2 11 2 16 13 10 9 3 0 1 10 9 2
15 10 9 1 11 13 1 10 0 1 10 11 1 10 9 2
27 10 2 1 10 9 2 0 9 0 4 13 10 9 10 11 11 2 12 2 2 1 11 11 7 11 11 2
19 10 9 1 10 0 9 7 10 9 1 9 13 10 9 0 1 10 9 2
83 10 9 13 10 9 2 16 10 9 13 13 7 13 10 9 0 2 13 1 10 9 0 16 13 10 9 1 10 9 2 9 7 9 0 1 10 9 2 15 4 13 1 10 11 11 1 11 7 11 1 10 11 2 11 11 2 15 1 10 9 15 13 1 11 11 1 10 9 2 15 16 15 13 0 13 10 9 7 13 10 0 9 2
27 10 0 7 0 9 13 10 9 1 9 1 10 0 9 16 13 10 9 1 9 1 10 9 1 10 9 2
29 11 13 13 1 10 9 13 1 10 11 2 7 16 15 13 13 10 9 1 10 9 0 13 10 9 13 1 11 2
70 1 10 9 2 10 9 13 10 9 1 9 16 4 13 15 1 10 9 0 2 9 2 9 2 9 2 9 8 2 9 9 2 10 9 2 10 11 2 2 16 13 10 9 0 1 10 9 2 13 10 9 1 9 1 9 0 2 0 7 0 2 1 10 16 13 9 1 10 9 2
22 1 10 9 1 10 11 2 3 11 13 1 11 1 11 7 13 1 10 9 1 9 2
11 2 15 4 13 16 3 4 13 10 11 2
6 2 15 13 10 9 2
27 13 10 9 0 1 10 9 16 10 9 13 16 10 9 13 9 7 16 13 15 13 10 9 1 10 9 2
29 11 13 10 9 0 7 0 1 10 9 0 1 9 7 9 3 0 7 3 0 1 11 2 1 3 1 12 8 2
32 16 10 9 13 1 11 2 10 12 1 11 1 12 13 3 1 10 9 1 9 0 2 1 10 13 10 9 1 10 9 2 2
12 13 1 10 9 0 2 11 11 2 11 2 2
47 11 2 15 13 1 10 9 1 3 1 10 9 2 3 13 3 10 9 1 0 2 13 9 1 15 3 0 1 9 0 2 7 1 9 13 9 0 1 10 9 1 10 9 1 10 9 2
21 1 10 12 3 10 9 1 11 2 11 11 13 11 15 13 1 13 15 1 15 2
19 3 13 10 9 1 2 9 2 2 1 9 1 10 12 1 11 1 12 2
30 15 13 1 13 10 9 7 15 4 1 13 10 9 2 1 10 15 15 15 13 1 10 0 9 2 13 10 9 8 2
42 10 8 8 0 13 9 3 0 1 9 2 13 1 9 7 13 1 10 9 1 9 0 7 10 9 0 0 2 1 9 7 10 9 13 3 1 9 1 1 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
32 1 9 1 12 2 16 15 13 10 9 0 1 11 7 10 11 2 10 9 1 10 11 11 13 12 11 1 10 11 11 11 2
10 11 11 13 10 9 9 1 9 0 2
8 3 13 9 1 9 7 9 2
27 3 11 11 2 10 9 1 11 16 13 9 7 9 0 2 15 13 1 10 9 0 1 13 10 9 11 2
14 15 13 10 9 3 7 10 9 16 15 13 3 3 2
18 10 0 9 13 10 9 13 1 10 9 11 11 2 0 1 11 11 2
19 1 15 15 13 15 2 7 1 15 10 9 2 3 4 1 13 10 9 2
17 13 10 0 9 7 10 10 9 1 13 7 13 0 7 0 9 2
9 1 13 1 10 9 1 10 11 2
38 10 11 2 12 4 4 13 7 4 3 13 1 10 11 1 11 11 7 3 1 10 11 11 1 11 1 11 7 1 10 9 1 10 11 11 1 11 2
21 13 9 1 10 11 1 11 1 11 11 7 13 9 1 11 11 1 10 11 11 2
42 3 2 13 13 10 9 1 9 1 10 9 13 15 1 9 7 1 10 9 1 9 1 4 13 1 10 11 10 9 1 10 0 9 1 9 0 2 7 4 13 9 2
34 13 10 12 0 9 11 11 12 2 11 11 2 11 11 12 2 11 11 2 11 11 12 2 11 11 2 7 11 11 12 2 11 11 2
29 7 10 9 4 1 13 1 10 9 1 10 9 0 2 3 1 7 15 15 13 2 7 3 1 10 9 1 9 2
13 13 1 11 2 11 2 10 12 1 11 1 12 2
35 13 0 1 10 9 2 11 11 2 1 10 9 1 9 1 9 2 10 12 5 1 10 9 1 10 9 1 11 11 3 13 0 1 9 2
27 10 9 13 10 9 1 10 15 10 9 0 1 9 2 0 2 9 7 15 2 15 13 1 13 9 0 2
40 16 10 9 1 10 9 1 10 9 4 13 1 12 2 10 9 3 13 9 1 10 9 1 10 9 1 12 2 1 9 1 10 9 0 11 11 7 11 11 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
13 9 1 10 9 1 11 13 9 1 10 0 9 2
22 11 11 11 11 11 13 10 9 1 12 13 1 10 9 0 1 10 9 1 11 11 2
25 15 13 16 11 13 10 9 1 10 12 9 2 7 1 9 13 12 2 1 10 10 9 7 9 2
13 10 9 1 10 9 1 10 9 1 9 13 0 2
17 1 9 1 10 9 0 2 13 12 9 1 9 2 0 7 0 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
29 1 12 10 9 15 4 13 7 15 4 13 10 9 2 7 10 9 0 1 12 3 13 3 0 1 10 9 9 2
18 4 13 1 9 1 11 11 2 11 11 11 2 11 11 7 11 11 2
21 4 13 13 1 10 12 10 11 7 4 13 3 0 1 10 9 1 9 16 13 2
6 3 15 4 13 9 2
34 13 1 10 9 1 10 9 1 10 9 1 10 9 2 9 1 11 2 1 9 0 2 10 9 11 13 0 1 9 1 10 9 2 2
5 15 13 1 11 2
12 10 9 1 9 1 10 9 13 1 5 12 2
18 3 4 13 10 9 1 9 0 16 11 11 13 1 9 1 10 12 2
23 1 10 9 3 15 13 10 9 0 1 10 13 1 10 9 15 2 3 2 0 9 12 2
41 13 1 11 2 11 2 11 2 2 13 10 9 0 16 13 10 9 1 11 1 10 9 2 13 1 9 1 9 2 1 10 9 2 1 10 9 1 10 9 11 2
73 13 0 10 9 16 13 10 9 1 10 15 4 13 15 10 9 16 13 10 15 16 13 10 9 9 2 7 10 9 13 0 9 2 1 0 9 2 3 7 9 7 9 2 13 3 0 10 13 15 1 10 9 1 9 1 9 7 9 2 13 1 9 2 9 7 11 2 13 15 1 9 0 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
28 10 9 1 0 9 2 7 9 11 2 13 10 9 1 10 9 1 10 15 10 9 13 0 9 1 9 0 2
11 10 9 0 1 10 9 13 1 11 11 2
44 1 9 1 10 9 1 12 2 10 0 9 1 9 7 9 11 11 13 10 9 0 1 11 2 11 12 2 10 9 0 2 1 10 9 11 1 10 9 1 11 11 2 11 2
26 3 2 11 11 4 13 1 10 9 10 9 15 1 10 9 1 9 7 1 10 9 1 10 9 0 2
17 10 9 13 10 0 0 9 2 7 10 9 1 11 13 4 13 2
15 4 13 1 11 1 11 1 10 12 2 13 1 11 11 2
16 1 10 0 9 16 15 13 15 16 4 13 15 13 1 15 2
21 9 3 3 0 7 15 13 15 16 3 13 9 16 13 0 2 7 4 13 3 2
14 1 10 9 1 12 2 13 12 9 13 1 10 11 2
9 10 10 9 13 9 0 2 11 2
21 10 9 1 9 1 12 9 3 13 10 9 1 9 1 9 7 15 1 12 9 2
6 13 13 9 7 9 2
43 11 11 2 13 10 12 1 11 1 12 1 11 2 11 11 2 2 13 10 12 1 11 1 12 1 11 11 2 2 9 0 1 11 2 13 10 9 2 9 7 9 0 2
43 3 15 4 13 11 11 1 11 2 1 3 13 16 10 9 3 0 1 11 11 12 4 13 1 9 1 10 9 1 10 11 2 2 13 1 10 9 7 15 4 13 2 2
21 13 9 2 3 7 9 1 9 2 7 10 9 13 3 0 7 3 13 9 0 2
6 3 15 4 13 2 2
22 1 10 9 13 1 10 9 1 11 2 15 1 10 15 2 11 11 2 11 11 2 2
11 1 10 9 1 9 2 15 4 13 15 2
36 1 10 9 1 9 2 10 9 1 11 11 13 10 9 16 13 10 9 1 10 9 1 15 2 16 13 1 10 9 0 16 4 13 1 3 2
66 1 3 1 10 11 11 2 1 10 9 1 10 9 2 1 9 1 12 8 2 9 8 1 9 7 9 0 1 12 8 2 2 13 1 10 9 15 1 10 9 1 10 9 2 15 13 3 9 3 2 7 0 2 1 10 9 2 1 10 0 9 2 1 12 9 2
27 1 12 4 1 4 13 9 0 1 10 12 11 7 1 12 1 12 13 10 9 1 10 9 1 10 11 2
39 10 9 1 9 13 13 0 1 15 15 3 13 10 9 1 10 9 0 3 16 13 10 9 1 10 9 0 2 1 10 9 3 0 1 10 9 3 0 2
24 1 10 9 2 13 10 9 1 10 9 1 13 1 11 2 10 9 4 13 1 10 11 11 2
26 15 13 1 11 1 9 1 11 1 13 10 9 1 10 9 1 11 7 13 1 11 11 1 9 0 2
24 10 9 1 10 9 1 9 11 15 13 7 13 10 9 0 7 10 9 0 1 10 9 0 2
12 11 13 10 9 0 1 10 9 1 11 11 2
26 1 10 9 2 16 4 13 9 1 9 1 9 0 2 11 13 16 15 7 15 15 13 1 10 9 2
28 10 9 13 1 10 9 13 1 10 9 12 1 0 9 2 9 12 1 12 9 7 9 12 7 12 1 9 2
24 1 11 2 10 9 13 1 10 12 9 1 9 2 9 15 3 4 4 13 1 10 0 9 2
38 10 9 1 10 9 1 10 9 13 3 13 1 10 9 1 11 1 10 0 9 1 11 11 11 9 2 15 13 3 2 1 2 15 13 3 0 2 2
23 1 9 0 2 10 12 1 11 2 10 9 4 13 3 1 9 1 10 11 1 10 11 2
9 15 4 13 13 15 0 9 0 2
5 15 13 12 5 2
56 10 9 1 13 15 3 15 13 1 13 10 9 15 1 12 9 13 2 10 11 2 1 15 3 0 1 10 15 13 2 10 11 2 2 10 15 13 1 10 9 0 13 1 10 11 11 7 13 1 10 11 1 11 1 11 2
14 10 9 13 1 10 9 1 10 9 0 2 11 11 2
24 1 9 2 10 9 1 10 9 1 10 11 11 13 10 9 1 2 9 0 2 16 15 13 2
57 12 9 3 2 10 12 1 11 1 12 2 10 9 13 9 1 13 10 0 9 2 10 15 4 13 1 11 11 2 1 10 9 13 10 9 10 9 13 1 10 9 11 7 11 11 11 2 0 7 1 10 9 1 10 9 11 2
39 13 1 12 9 10 11 11 11 11 2 10 0 9 1 10 9 1 10 9 9 2 7 1 10 12 9 10 11 11 11 11 2 0 9 0 1 9 0 2
25 13 10 9 0 1 10 11 2 9 0 2 11 2 11 2 11 2 9 2 9 7 9 1 15 2
11 1 3 13 15 10 9 16 13 10 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
18 10 10 9 1 10 9 15 13 1 9 9 1 10 9 1 10 9 2
17 10 9 15 13 13 10 10 9 1 10 9 2 10 9 13 0 2
8 1 11 9 2 15 13 3 2
11 1 10 9 13 10 9 11 11 1 11 2
32 1 10 9 0 1 10 9 1 10 9 10 9 15 13 16 10 9 1 9 13 9 15 10 9 1 10 9 13 9 1 13 2
12 10 9 0 13 10 9 0 16 13 1 9 2
50 1 10 9 2 15 13 10 9 2 7 10 9 1 10 11 13 0 2 13 15 1 11 2 15 13 10 9 0 7 0 1 10 2 10 9 0 7 0 15 13 10 10 9 2 7 15 1 10 9 2
15 10 9 13 0 16 16 13 9 4 13 1 10 11 0 2
16 10 9 15 13 9 1 11 2 13 10 9 1 0 9 0 2
69 11 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 10 9 0 16 13 9 0 3 1 13 10 9 1 0 11 11 1 10 3 9 0 1 10 11 11 1 10 11 11 2 11 11 2 7 16 15 15 13 13 15 3 1 13 10 11 11 2 15 15 11 13 2
12 1 10 9 2 11 4 13 1 11 1 12 2
37 1 10 12 9 2 1 13 10 9 2 13 1 10 11 11 11 11 3 13 10 9 1 9 2 13 3 10 0 9 1 10 9 7 1 9 0 2
51 1 9 2 10 9 0 13 10 0 9 0 2 10 9 1 10 9 4 13 1 10 9 1 10 9 1 9 1 9 2 9 7 9 2 7 1 0 9 1 9 16 2 0 1 10 9 2 13 0 9 2
30 1 15 9 2 10 9 0 13 3 0 7 10 9 0 2 7 13 3 1 9 2 16 4 13 0 2 0 7 0 2
19 3 2 16 13 10 9 11 2 10 9 4 13 9 16 13 10 0 9 2
28 1 15 13 10 9 1 10 9 2 1 10 9 2 1 10 9 2 15 13 1 10 9 0 2 10 9 0 2
18 10 9 1 10 11 13 10 9 1 10 9 0 1 11 2 12 2 2
43 10 11 13 10 9 1 10 9 1 10 9 0 1 11 1 10 8 9 1 9 11 11 11 7 10 12 9 1 9 1 0 9 2 13 1 10 9 1 10 0 9 0 2
28 4 13 10 9 1 10 0 9 16 4 13 1 11 1 13 10 0 9 1 10 15 15 4 13 2 11 11 2
39 11 11 13 1 10 0 9 1 11 1 11 1 11 1 11 11 11 11 1 11 1 10 3 11 1 11 11 11 2 3 11 2 10 12 1 11 1 12 2
39 10 0 9 13 9 1 11 1 12 1 10 11 2 12 2 3 1 10 9 11 11 1 10 15 15 13 10 9 12 7 10 9 11 16 13 3 10 9 2
23 3 1 13 1 10 9 9 2 10 9 1 10 9 13 9 1 9 1 10 9 1 9 2
30 10 9 1 11 13 10 9 1 10 9 1 13 16 13 3 10 9 0 7 0 1 10 9 16 13 7 13 10 9 2
43 15 13 10 9 1 10 15 11 13 10 9 1 10 9 1 10 13 2 10 9 1 9 11 11 2 11 1 11 2 13 11 2 7 3 10 0 9 11 13 1 11 0 2
40 1 15 2 16 15 13 9 7 15 13 3 13 10 9 2 7 3 15 13 3 16 10 9 0 7 0 3 15 13 1 10 9 2 3 1 10 9 1 11 2
25 3 2 10 9 0 4 13 2 15 15 13 1 10 9 1 11 1 13 10 0 9 1 10 9 2
45 1 10 9 1 10 11 15 4 13 9 11 1 10 9 1 11 7 11 2 11 2 11 2 2 16 13 9 1 10 9 1 10 9 1 11 7 3 1 10 9 1 10 9 11 2
40 16 10 9 0 1 9 2 10 9 1 11 11 11 11 2 3 13 10 9 1 10 9 1 9 11 11 2 4 13 15 1 10 9 1 9 1 10 9 9 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
45 16 1 10 0 9 15 15 13 1 10 9 0 1 10 9 0 2 1 10 11 3 15 13 3 2 3 16 10 9 1 10 9 15 13 3 1 10 9 0 7 1 10 9 0 2
8 2 15 13 10 0 9 0 2
27 3 2 2 1 15 4 13 10 9 1 10 0 12 9 16 10 11 13 16 3 13 9 10 12 0 9 2
19 1 9 15 3 3 13 3 2 7 15 3 0 13 4 15 7 13 3 2
27 1 9 2 10 12 5 1 10 9 13 1 10 9 1 9 2 3 7 10 12 5 0 1 10 1 9 2
9 15 3 4 13 9 1 10 9 2
32 11 13 1 12 7 0 1 10 9 1 9 11 11 11 2 13 15 1 10 9 9 1 10 9 0 1 9 1 9 1 9 2
19 15 13 10 9 1 9 0 2 12 9 1 9 7 12 9 1 9 0 2
19 15 13 1 10 9 0 2 1 11 11 2 11 2 11 7 1 10 9 2
24 10 9 13 9 1 11 2 16 4 13 1 10 9 1 11 1 15 13 10 9 0 7 0 2
18 2 13 0 1 10 11 7 13 15 16 13 10 11 2 2 4 13 2
25 13 1 10 9 1 11 2 1 10 9 1 11 2 1 10 9 1 11 7 1 10 9 1 11 2
19 10 9 4 13 1 10 9 11 11 7 11 2 8 2 1 11 2 11 2
28 3 4 13 10 11 1 10 11 11 1 11 2 16 13 1 9 1 9 0 2 12 9 7 10 9 0 0 2
13 2 10 9 4 13 13 10 12 9 1 9 0 2
16 10 11 11 13 3 10 9 0 7 0 2 12 1 12 2 2
7 10 9 13 0 1 9 2
38 1 10 9 3 13 10 9 7 9 16 13 3 0 1 13 10 9 1 10 9 1 10 11 7 10 9 4 13 2 7 3 2 3 0 1 15 13 2
49 9 1 11 1 11 7 10 11 1 10 11 1 11 11 7 10 11 7 11 11 11 1 11 11 13 1 10 9 3 0 7 3 2 0 2 2 3 0 1 10 9 1 10 9 1 10 9 0 2
39 15 0 3 13 1 10 9 1 9 11 12 1 11 2 15 2 1 10 9 1 10 9 1 10 9 0 0 1 11 15 13 1 13 11 7 13 10 9 2
38 16 10 9 13 0 1 10 10 9 1 10 9 2 10 9 0 1 10 9 0 4 13 1 10 9 1 10 9 1 9 0 1 9 11 2 8 2 2
21 15 13 1 9 2 7 13 1 11 2 7 3 1 10 9 1 9 1 11 11 2
23 13 1 10 11 1 10 11 2 7 10 9 0 15 13 3 1 10 1 10 9 1 11 2
22 4 13 1 0 9 16 13 1 9 0 1 10 9 7 0 7 0 1 10 9 0 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
30 13 16 10 9 1 10 9 13 0 1 10 9 7 15 1 15 1 13 15 1 13 10 9 16 15 15 13 1 9 2
10 13 3 13 15 1 11 3 1 15 2
38 1 10 9 2 10 9 11 13 1 11 3 7 10 9 1 10 9 11 11 13 1 10 11 2 1 10 12 9 1 10 9 2 9 0 1 10 9 2
20 10 9 13 3 10 9 1 10 10 9 2 15 16 11 13 13 1 9 3 2
11 15 13 1 9 7 13 1 10 15 13 2
20 1 10 9 2 11 4 1 13 10 9 3 16 11 4 13 1 10 9 11 2
39 3 13 9 1 10 9 0 2 16 3 15 4 13 2 7 4 13 3 3 10 9 0 1 10 9 0 2 7 3 15 0 7 10 9 15 13 10 9 2
12 11 11 13 10 9 1 9 0 1 11 11 2
14 11 13 1 12 9 2 12 9 7 12 9 1 9 2
9 13 10 0 9 0 0 1 11 2
49 10 9 1 10 11 7 11 4 13 1 10 9 13 1 11 1 11 1 12 9 7 10 9 13 16 10 9 1 9 16 13 1 12 9 13 3 1 10 9 1 10 13 1 10 10 9 1 11 2
28 10 9 15 13 11 13 10 9 1 10 9 1 10 9 2 1 10 9 1 9 0 7 0 7 10 9 0 2
18 15 13 16 13 15 3 12 9 10 9 1 10 9 0 7 10 9 2
32 11 2 11 11 2 11 2 12 2 11 2 12 2 13 10 9 0 2 9 1 9 7 9 1 10 0 9 1 10 9 12 2
21 16 15 13 2 10 9 1 10 9 9 1 13 7 10 9 13 9 1 10 9 2
36 3 15 13 10 9 1 9 13 10 9 2 7 13 10 9 1 9 1 10 9 11 16 13 10 9 1 10 9 1 9 0 1 10 9 11 2
19 1 10 10 9 1 11 2 15 13 1 10 9 1 10 15 13 12 9 2
29 10 9 11 11 2 11 11 2 11 11 7 11 11 3 15 13 1 10 9 1 13 1 10 9 7 13 10 9 2
68 2 13 16 10 9 13 9 0 1 9 1 10 9 1 10 9 16 13 7 16 1 10 0 9 16 13 13 15 1 15 16 13 10 9 15 13 1 10 9 7 1 10 9 2 16 3 15 13 1 9 9 1 10 9 1 10 9 2 16 3 4 13 9 2 2 13 11 2
24 15 15 13 9 1 16 3 13 10 9 7 10 0 9 13 10 9 1 10 9 1 10 11 2
16 1 9 0 2 10 9 13 1 0 9 7 0 9 1 13 2
29 10 12 1 11 1 12 2 10 9 13 10 9 1 10 11 11 1 11 0 2 3 1 10 11 11 11 11 11 2
25 1 10 9 13 10 9 0 1 10 9 0 7 3 13 13 10 9 1 9 7 15 13 1 11 2
29 10 12 1 11 10 9 4 13 1 10 12 11 1 9 1 10 9 1 11 11 0 1 10 10 9 1 10 9 2
98 10 9 13 1 11 15 13 1 9 1 10 9 1 2 11 7 11 2 10 9 15 13 1 10 9 2 2 11 11 2 1 9 1 9 7 9 2 2 10 11 2 9 7 9 1 9 2 2 10 9 2 3 10 9 3 13 3 10 9 2 2 11 11 2 3 0 7 8 2 8 2 2 11 2 10 9 1 10 12 7 12 9 2 7 11 2 9 7 9 1 10 9 1 10 9 0 2 2
54 10 9 1 10 9 1 10 9 1 9 1 10 9 13 16 10 9 0 1 9 0 4 1 13 8 5 2 8 2 12 2 1 9 2 12 9 1 9 13 10 9 7 15 13 3 1 10 9 1 13 3 10 9 2
7 11 11 4 13 1 11 2
20 1 10 9 2 11 13 0 2 13 1 10 0 9 7 1 9 1 4 13 2
30 1 0 10 9 4 13 0 1 15 13 10 0 9 1 10 9 3 7 13 1 12 9 13 1 10 9 1 10 9 2
6 13 0 1 10 0 2
16 1 12 2 13 10 9 0 1 10 9 1 11 11 11 11 2
9 4 13 1 10 9 1 9 0 2
36 11 2 1 9 11 2 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 1 11 2 11 2 1 10 9 1 11 7 9 1 11 2
11 10 9 1 11 15 13 13 1 10 9 2
23 3 3 1 4 13 10 0 9 2 10 9 13 1 9 1 10 0 9 2 1 0 9 2
11 10 9 1 10 11 11 13 8 8 15 2
9 3 13 9 1 10 9 1 11 2
29 10 9 0 1 11 13 10 3 9 1 10 11 7 15 13 1 10 12 9 1 9 1 11 11 2 13 10 9 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
21 10 12 1 11 1 12 13 13 15 1 9 1 11 2 11 2 7 13 1 9 2
35 10 9 0 2 3 1 9 2 1 9 8 2 8 13 1 9 8 2 13 10 0 9 1 9 1 0 8 8 2 16 3 4 1 13 2
17 11 4 13 10 9 0 0 1 10 9 1 10 9 0 1 9 2
16 10 9 1 10 9 1 10 9 2 13 10 9 1 10 11 2
46 11 11 11 2 11 2 3 13 1 10 9 11 11 7 11 11 2 11 11 2 12 1 11 1 12 2 8 2 12 1 11 1 12 2 2 13 10 9 0 1 9 0 7 1 9 2
26 3 2 15 15 13 10 12 1 11 1 12 1 9 0 1 10 9 9 0 1 10 9 1 9 0 2
30 11 13 10 9 7 9 0 2 1 10 9 1 11 11 2 9 1 11 11 2 1 10 9 1 11 7 9 1 11 2
36 10 9 0 7 0 13 9 1 10 9 1 9 2 9 1 10 9 2 2 16 15 13 1 13 10 9 0 7 0 1 10 9 1 10 9 2
12 11 4 13 1 3 10 9 1 10 9 0 2
23 15 10 9 1 11 1 10 1 11 13 2 3 1 10 9 1 11 1 12 2 9 0 2
28 13 0 1 9 9 10 12 1 11 2 7 3 13 10 9 12 1 11 7 15 13 1 10 9 1 11 11 2
32 11 11 11 2 12 1 11 1 12 2 11 2 11 2 12 1 11 1 12 2 11 11 2 11 2 13 10 9 7 9 0 2
17 11 2 13 10 9 0 1 9 0 0 1 10 9 1 10 11 2
40 10 9 1 9 8 2 11 2 1 9 1 11 1 10 11 7 10 11 2 11 2 15 13 1 13 10 9 1 9 0 0 1 11 2 11 1 9 11 2 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
71 1 10 9 1 3 11 1 11 3 4 13 9 1 9 1 9 2 3 0 1 0 2 15 3 3 13 9 1 9 1 10 9 2 1 9 1 10 9 11 11 11 2 1 9 2 11 11 2 7 11 1 11 2 11 2 10 15 4 13 10 0 9 1 9 1 10 9 1 9 0 2
60 12 9 4 13 0 7 15 4 13 9 2 1 10 9 0 2 1 9 1 10 9 0 1 12 9 2 15 0 7 15 0 2 13 10 9 1 11 1 11 2 11 2 2 1 10 9 11 2 12 2 4 13 9 1 10 11 11 1 11 2
22 13 3 0 7 13 1 10 9 16 15 4 4 13 1 10 9 10 9 7 10 9 2
44 10 9 1 10 11 2 15 13 1 13 15 1 10 9 7 1 13 10 9 1 9 0 7 10 9 1 13 10 9 1 9 2 13 1 10 9 2 13 10 9 1 9 0 2
13 4 13 10 9 16 15 15 13 9 7 9 0 2
12 1 10 9 0 13 10 12 9 11 11 11 2
71 10 9 2 11 11 2 13 1 10 9 1 10 0 11 1 11 2 13 1 13 10 9 1 9 1 10 9 12 2 7 13 1 13 15 1 12 1 10 9 2 16 15 13 0 2 11 11 1 11 2 9 0 1 11 2 7 11 11 1 11 2 9 0 1 10 9 1 11 1 12 2
18 9 0 1 9 0 2 1 9 0 7 9 1 9 2 13 1 12 2
38 10 9 1 10 9 1 9 1 10 0 9 15 13 10 12 1 11 1 12 2 3 3 15 13 10 9 11 11 10 12 1 11 1 12 1 11 11 2
26 10 11 11 13 10 9 13 10 0 11 1 10 9 1 11 1 10 9 1 11 11 2 11 2 11 2
46 13 10 9 16 10 9 11 10 11 2 11 11 10 11 7 11 11 15 13 1 10 9 1 13 10 9 1 10 9 2 7 16 15 1 10 9 15 13 10 15 13 1 10 0 9 2
22 10 9 0 1 11 11 15 13 1 10 9 0 11 11 12 1 15 0 11 13 12 2
15 13 1 10 9 2 9 13 1 9 0 2 7 10 9 2
9 2 2 2 13 10 9 2 2 2
16 16 15 13 0 2 10 9 4 13 1 10 9 1 10 9 2
13 0 7 0 2 13 9 2 7 3 13 10 15 2
42 2 15 2 10 9 1 11 2 13 10 9 0 3 1 11 11 7 13 13 15 1 15 16 13 13 10 11 2 2 13 11 11 2 9 1 10 9 2 11 11 2 2
35 10 9 0 1 10 9 4 13 7 13 1 12 9 0 2 10 15 1 10 15 13 10 9 0 1 9 2 9 2 9 7 9 1 9 2
48 10 9 11 13 0 16 10 9 4 13 7 10 9 1 10 9 7 10 9 2 16 3 11 4 13 2 15 13 13 1 10 9 1 13 15 1 3 2 7 13 13 1 10 9 1 10 9 2
12 10 9 1 9 1 10 9 13 1 5 12 2
30 10 9 4 13 1 10 9 11 1 10 11 1 12 3 3 1 11 11 2 1 13 1 10 15 10 9 13 10 9 2
42 3 2 1 10 11 1 11 2 10 11 15 4 13 10 9 1 10 2 0 2 9 2 13 13 1 10 9 7 9 1 10 9 13 10 9 7 9 1 9 3 0 2
18 11 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
26 1 10 9 1 10 9 0 10 9 13 13 10 9 1 9 0 1 13 10 9 7 13 13 10 9 2
35 11 1 9 15 13 1 10 9 3 0 2 7 13 3 1 16 11 11 13 10 9 1 11 12 2 7 10 9 4 7 13 1 10 9 2
29 15 1 15 2 10 0 9 2 13 10 9 1 11 1 10 9 15 9 11 7 10 9 13 1 11 11 1 11 2
38 15 13 1 10 11 13 10 9 0 1 16 3 13 10 13 9 7 13 3 1 10 12 9 2 16 3 13 1 9 1 9 16 13 9 7 13 9 2
22 13 10 12 1 11 1 12 1 11 1 11 2 11 2 13 9 1 10 9 11 11 2
15 10 0 9 15 13 8 11 1 10 9 1 11 7 11 2
36 13 9 0 7 9 1 9 0 16 13 13 10 9 1 11 2 9 1 9 1 9 16 13 13 9 0 1 0 9 13 1 9 1 9 2 2
20 1 10 10 4 9 1 11 13 10 9 7 3 13 10 9 1 9 1 11 2
47 1 9 0 15 13 9 1 10 9 0 2 3 1 10 0 9 2 3 1 10 9 0 1 10 9 2 1 10 0 9 7 9 7 0 1 10 9 0 2 3 3 4 13 15 10 9 2
14 10 9 3 15 13 3 3 1 10 9 1 10 9 2
40 10 9 13 3 10 9 1 9 1 0 9 1 11 2 13 10 9 3 0 10 16 13 1 10 9 12 1 11 2 11 2 2 8 1 10 9 10 11 11 2
25 1 10 9 2 11 13 16 11 2 16 1 10 9 13 3 12 9 2 13 10 9 0 1 11 2
24 1 10 9 4 13 10 11 2 10 9 1 0 9 0 1 13 10 9 0 1 9 1 9 2
52 10 9 1 10 9 3 1 10 9 13 1 10 9 0 7 0 2 3 10 9 15 13 1 9 0 16 3 15 13 1 10 9 1 10 9 2 3 15 13 10 9 2 1 3 13 15 1 10 10 9 0 2
22 16 10 9 0 4 13 3 2 15 13 3 16 10 9 1 9 13 10 9 1 9 2
14 1 0 9 15 13 10 9 2 13 1 10 9 0 2
27 3 3 10 9 13 1 9 2 10 9 1 9 7 9 1 9 13 0 7 13 10 9 1 9 7 9 2
29 1 15 1 12 4 13 9 2 10 9 13 1 10 9 1 10 11 2 16 3 13 7 10 0 9 7 0 9 2
19 1 10 9 2 10 9 3 13 10 0 9 1 10 9 0 1 10 9 2
39 10 9 1 10 9 0 7 10 9 1 9 1 9 1 10 9 0 13 10 9 1 9 13 1 10 11 11 7 13 1 9 1 10 10 9 0 1 11 2
38 1 9 2 16 10 9 13 1 0 9 2 0 2 2 15 13 1 10 9 1 9 0 2 10 9 1 9 1 9 0 2 1 9 1 9 0 0 2
32 3 1 10 11 1 10 9 12 13 0 10 9 11 2 8 2 8 2 8 2 8 2 7 11 2 8 2 5 2 8 2 2
36 10 9 1 10 11 13 10 9 0 2 10 9 2 11 2 8 13 10 9 1 13 1 10 9 1 9 7 13 15 4 1 13 1 10 9 2
25 1 11 2 1 10 0 7 1 10 0 11 2 10 9 13 10 0 9 0 2 13 1 10 9 2
20 10 9 0 0 13 15 1 10 9 2 3 10 9 2 16 13 3 10 9 2
21 11 11 11 13 10 9 0 13 1 11 2 11 2 1 12 7 13 1 9 0 2
39 11 11 2 11 2 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 10 9 0 2 1 0 9 1 10 9 0 0 1 10 9 0 7 0 2
15 10 11 1 11 13 1 10 11 11 11 12 9 3 9 2
16 10 0 9 0 1 10 9 13 11 11 2 13 1 12 8 2
14 10 9 13 1 10 9 0 1 10 15 13 10 9 2
27 10 9 1 10 9 13 1 10 9 11 2 0 2 7 11 2 9 0 2 2 1 9 1 10 9 0 2
26 3 2 10 9 13 0 1 13 7 13 1 10 9 1 10 9 2 15 16 3 13 1 11 2 11 2
56 10 9 1 9 15 13 1 15 1 10 9 7 9 0 1 10 9 2 9 1 9 2 9 1 9 2 9 1 9 2 8 2 13 1 10 9 0 2 1 10 9 1 9 2 0 1 10 9 1 10 9 7 10 9 2 2
57 10 9 1 9 0 1 9 0 2 7 10 0 9 0 2 13 10 0 9 1 10 9 13 2 1 10 9 0 0 2 7 3 11 13 1 10 0 9 1 10 9 1 10 9 0 2 1 15 1 10 9 0 7 1 10 9 2
15 10 9 0 13 2 9 2 9 2 9 2 9 7 9 2
9 15 13 1 9 1 10 9 12 2
31 3 7 2 1 10 15 1 10 9 15 13 9 1 9 16 13 10 9 7 13 13 10 9 1 9 0 1 10 9 0 2
27 1 12 15 13 1 0 2 10 9 1 9 1 10 9 1 10 9 12 1 10 9 2 13 15 1 9 2
31 11 13 16 13 11 11 11 15 2 13 1 10 9 2 1 10 9 2 13 10 9 1 9 16 13 1 10 9 1 11 2
35 1 10 0 9 1 15 15 13 10 9 0 11 11 11 2 9 0 16 4 13 9 1 9 2 9 2 9 0 7 9 0 2 1 15 2
15 13 3 16 16 13 1 10 9 4 13 10 9 3 0 2
14 13 10 12 1 11 1 12 16 4 13 12 1 12 2
39 13 10 9 0 1 9 1 10 9 1 10 9 0 7 10 9 1 10 9 0 2 1 10 9 1 9 7 9 2 13 10 9 7 10 9 2 3 2 2
17 11 13 10 9 1 9 1 9 2 13 1 10 9 11 11 11 2
45 11 2 3 4 7 13 15 2 13 10 9 13 1 10 2 9 2 1 10 9 1 11 11 2 9 1 9 1 10 15 13 10 2 9 2 1 11 11 7 15 13 0 9 3 2
22 13 13 10 9 1 12 1 10 13 15 10 11 11 11 2 13 1 13 9 1 9 2
12 13 13 16 1 3 1 3 13 0 13 9 2
10 7 3 13 9 1 10 9 3 0 2
34 3 1 10 0 9 2 9 2 9 2 9 7 9 13 13 10 9 2 1 15 15 15 4 1 13 1 10 0 9 0 1 9 0 2
13 3 15 13 15 1 13 2 13 10 9 1 13 2
13 10 0 9 13 1 9 16 4 13 1 10 9 2
9 7 3 15 13 10 9 3 3 2
23 10 9 15 13 1 10 11 2 11 2 11 2 11 7 1 10 9 1 9 1 10 9 2
39 10 9 1 9 1 15 9 1 10 0 9 2 16 13 3 3 1 10 9 1 10 9 2 1 9 3 0 1 15 9 1 10 9 0 2 1 0 9 2
32 11 1 10 9 13 10 9 1 9 0 2 10 9 15 4 13 1 13 9 1 9 0 2 1 9 0 7 9 0 7 0 2
8 11 15 13 13 1 10 9 2
46 10 9 4 13 1 12 1 10 2 11 11 1 10 9 2 1 10 3 9 1 11 11 2 11 11 11 2 15 13 1 11 1 12 1 10 11 0 1 10 9 2 10 9 11 11 2
21 10 9 15 13 1 10 9 0 2 7 10 9 1 9 1 10 9 1 9 2 2
16 7 10 0 9 1 9 1 10 9 13 9 0 1 0 9 2
21 10 11 3 4 13 16 2 1 9 1 11 2 13 10 9 1 11 11 1 11 2
3 11 13 2
40 1 9 0 2 10 9 13 0 9 1 9 7 9 2 9 1 9 2 9 3 0 7 9 9 9 2 1 10 16 10 9 1 9 13 1 9 13 10 9 2
18 1 15 10 9 13 10 9 2 10 9 2 2 9 2 1 10 9 2
66 13 0 16 10 0 9 1 10 9 0 1 10 15 15 13 0 2 7 10 9 1 10 9 1 9 2 13 1 9 1 11 11 2 13 15 1 10 9 10 9 1 10 12 1 11 1 12 1 10 9 1 1 11 2 2 4 13 10 9 1 10 9 1 10 9 2
7 3 13 1 10 11 11 2
55 3 2 15 13 1 10 9 10 9 1 0 9 1 9 0 1 10 9 2 11 11 2 7 12 9 2 11 11 2 2 7 10 9 1 9 0 2 13 9 1 10 9 1 9 2 11 11 2 11 11 7 11 11 2 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
23 1 10 9 3 15 4 13 10 9 7 2 7 10 9 0 16 3 15 4 13 9 0 2
26 9 0 7 0 2 1 9 0 1 10 9 0 1 10 9 3 1 9 0 2 1 15 10 9 2 2
30 13 3 0 1 15 7 13 1 13 10 0 9 1 3 13 10 9 2 7 15 13 1 10 9 1 10 9 1 9 2
54 1 10 11 4 13 16 15 13 10 9 1 13 10 9 2 2 1 13 15 1 10 9 16 10 9 13 10 0 9 1 13 10 0 9 1 10 9 2 1 10 16 15 13 13 10 0 9 0 1 10 16 13 2 2
54 11 13 16 10 9 1 10 11 13 1 10 2 3 0 9 1 10 9 2 7 13 16 2 16 3 10 9 15 13 9 1 10 9 16 13 2 16 13 0 2 2 4 7 13 15 16 4 13 10 9 1 10 9 2
44 10 9 0 13 16 10 9 13 3 2 16 3 15 13 10 9 7 10 9 2 16 10 9 0 13 16 10 9 13 1 9 1 10 9 0 1 10 9 0 1 9 1 11 2
76 1 10 9 2 15 15 13 1 9 7 13 1 15 10 0 9 1 10 11 1 10 11 3 11 2 13 3 1 13 15 1 9 2 9 2 9 2 9 7 0 9 2 13 3 9 16 13 1 9 0 7 16 13 13 1 9 1 10 9 1 11 11 2 9 2 2 11 1 11 2 11 11 7 11 11 2
45 1 15 3 13 0 10 9 1 10 9 0 7 10 9 0 1 10 9 2 7 16 13 10 0 9 0 1 10 10 11 2 1 10 9 2 10 11 2 1 10 9 1 10 9 2
28 13 9 1 9 0 7 9 1 10 11 1 10 11 11 7 9 0 1 10 11 11 2 1 10 11 1 11 2
33 13 10 9 1 9 1 10 12 9 1 10 9 1 9 1 11 11 2 8 9 1 9 2 9 0 7 9 1 0 9 0 2 2
27 3 1 10 9 2 10 9 16 13 7 13 1 10 9 1 10 0 9 4 13 1 10 9 1 10 9 2
16 1 0 9 13 10 9 1 9 1 9 2 11 8 8 8 2
18 10 9 13 10 9 0 1 9 12 9 1 10 9 12 1 10 9 2
36 1 9 2 3 1 13 1 12 10 9 3 15 13 7 4 13 7 15 4 13 16 10 9 0 1 11 3 4 13 1 10 9 12 7 0 2
17 12 9 3 3 4 3 13 2 7 10 9 4 13 1 10 11 2
18 13 10 9 9 2 9 1 9 1 9 0 1 10 9 1 11 11 2
23 4 13 12 9 7 7 4 13 10 9 7 15 4 13 1 10 9 0 1 15 16 13 2
34 3 2 11 4 4 13 10 9 1 10 9 1 10 11 1 11 2 2 10 9 1 11 2 2 1 10 0 9 1 10 11 1 11 2
10 15 13 1 10 9 7 15 15 13 2
14 1 10 9 12 3 13 12 9 1 12 1 12 9 2
34 10 9 13 10 11 11 1 9 1 10 11 2 3 16 11 11 11 13 1 10 0 9 10 11 1 11 1 10 11 11 1 10 11 2
39 1 10 9 1 11 7 15 1 10 11 2 13 1 10 11 7 0 1 10 11 10 9 1 11 15 13 1 10 9 1 12 9 1 10 9 1 10 9 2
28 1 0 9 1 9 2 10 9 13 12 9 16 3 13 15 1 10 9 2 13 10 9 7 13 9 1 9 2
15 4 4 3 13 10 9 0 2 3 10 9 1 10 9 2
37 1 10 10 9 0 7 2 7 0 2 10 9 0 1 10 9 2 13 1 10 9 11 11 2 13 16 10 9 15 13 7 13 7 13 10 9 2
30 10 9 0 13 10 0 9 0 2 0 2 1 15 15 10 9 1 10 9 4 13 1 9 1 9 7 9 1 9 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
24 10 9 1 9 0 13 10 11 10 11 2 11 2 11 2 11 1 10 11 7 11 1 15 2
13 10 9 1 10 9 13 0 1 10 1 10 9 2
26 3 2 16 10 11 11 13 1 10 11 11 11 12 7 15 13 10 9 2 11 15 13 1 13 15 2
10 3 3 2 3 10 9 4 13 11 2
33 1 12 2 10 9 0 0 2 10 11 11 1 10 11 11 2 13 1 11 11 1 10 9 11 7 9 2 13 9 1 10 9 2
21 10 11 11 2 11 2 13 10 9 1 10 9 2 11 2 1 10 9 1 11 2
67 10 9 3 0 7 16 13 9 1 9 1 10 9 1 10 9 13 11 11 2 9 1 11 11 8 11 11 11 11 11 11 2 9 0 13 1 10 0 11 2 7 1 10 9 1 9 2 9 2 13 7 13 1 9 1 10 9 12 1 10 9 3 0 10 11 11 2
30 7 15 4 13 16 4 7 13 9 1 3 13 10 0 9 1 10 9 2 7 10 0 9 1 10 9 1 10 9 2
13 1 10 9 2 13 13 1 10 9 1 10 9 2
59 1 10 12 9 2 11 13 13 1 10 12 5 0 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
23 0 9 15 13 3 1 10 9 2 0 1 13 1 10 9 1 9 7 0 1 10 9 2
20 1 3 1 9 1 10 9 12 2 10 9 13 10 9 1 10 9 1 11 2
32 1 9 2 13 10 9 1 10 9 2 13 10 9 1 10 9 2 10 9 1 10 9 1 11 7 10 11 11 1 11 11 2
41 1 11 1 12 2 1 9 1 10 9 1 10 9 13 1 11 2 1 10 15 10 9 1 11 4 13 1 10 9 1 11 2 11 13 1 4 13 1 13 15 2
23 13 1 10 9 1 10 9 2 10 9 13 1 12 5 1 10 0 9 1 10 12 5 2
64 10 0 9 1 11 7 11 13 10 0 9 1 10 11 16 4 13 10 9 1 13 10 11 2 1 9 16 13 3 9 1 10 9 1 10 9 1 9 0 16 4 13 10 9 0 9 7 16 13 1 9 1 10 0 9 1 10 9 2 1 11 7 11 2
19 1 12 13 1 11 11 11 1 11 1 15 2 8 2 2 1 11 12 2
10 15 13 1 10 9 1 10 9 11 2
26 11 13 1 10 0 9 0 1 9 1 11 1 11 1 11 7 3 13 12 9 3 1 11 1 11 2
52 1 0 7 1 10 11 1 10 11 11 1 11 2 10 9 15 13 3 3 1 10 9 2 10 9 13 1 10 12 9 16 13 1 11 7 3 13 10 9 2 7 1 10 9 7 1 10 9 16 15 13 2
36 3 13 1 10 9 7 10 9 13 1 10 9 3 7 13 1 10 9 16 13 1 10 9 7 13 15 16 10 9 15 13 16 3 15 13 2
31 11 13 3 10 9 1 10 9 7 1 10 9 1 10 9 2 11 2 11 1 9 2 10 11 1 11 1 10 9 2 2
10 4 13 1 9 1 10 11 1 12 2
44 10 9 13 1 10 9 1 9 0 1 10 11 0 1 9 1 10 9 12 7 13 10 9 1 11 11 1 0 9 2 10 9 2 10 9 1 10 9 7 10 0 9 2 2
56 1 11 10 9 13 1 9 16 3 13 1 10 9 0 1 10 9 0 2 3 9 11 11 1 10 11 2 9 0 2 13 13 9 1 10 9 1 9 0 0 11 11 1 15 13 15 10 9 0 1 11 11 2 8 2 2
14 4 7 13 3 9 1 9 1 10 9 1 10 9 2
29 10 9 2 16 13 1 9 1 11 11 2 13 10 9 0 2 15 16 13 1 11 1 13 10 9 1 10 9 2
24 1 10 9 2 12 1 12 9 0 4 13 10 9 1 9 1 9 13 1 10 9 1 11 2
18 10 11 11 13 1 10 9 11 1 13 1 10 9 7 13 10 9 2
18 7 10 9 3 13 3 0 7 10 9 15 15 15 13 1 15 2 2
9 10 9 15 13 1 0 9 0 2
25 11 11 11 2 11 2 11 2 12 1 11 1 12 2 2 13 1 11 11 2 13 10 9 0 2
6 13 0 1 9 0 2
37 10 9 9 13 11 11 11 11 13 13 9 1 10 9 1 13 1 10 9 1 9 0 1 10 9 2 11 11 11 2 7 4 13 1 10 9 2
25 1 0 2 3 1 12 9 2 16 13 10 12 1 12 1 10 9 0 1 11 2 1 10 9 2
22 10 9 1 9 1 10 9 13 1 5 12 9 2 1 10 9 13 1 10 0 9 2
44 7 2 3 16 10 9 13 1 13 10 9 0 2 9 1 9 2 2 10 9 13 1 13 9 0 3 10 9 15 13 1 9 0 1 9 1 0 9 1 9 1 9 0 2
15 13 10 9 1 9 1 10 9 1 10 16 3 4 13 2
42 11 11 4 13 1 11 2 3 7 15 13 1 10 9 13 10 9 1 10 9 1 11 2 1 10 9 16 13 9 0 1 10 9 8 10 0 12 1 11 1 12 2
31 13 10 9 0 1 9 1 12 2 7 3 1 9 1 9 4 13 1 10 12 5 9 1 10 11 11 1 11 1 12 2
11 10 9 1 10 9 1 9 13 11 11 2
20 4 13 13 15 16 13 15 16 13 15 10 5 7 4 13 16 13 9 0 2
7 1 10 9 15 13 0 2
22 10 9 3 0 0 3 13 1 10 9 13 10 11 11 1 11 2 1 9 1 12 2
27 11 11 7 1 10 9 1 11 11 2 11 11 11 11 11 2 1 9 1 10 12 5 9 1 11 11 2
22 1 10 9 1 10 9 1 9 10 9 0 1 10 9 13 1 10 9 1 10 9 2
34 1 10 0 9 2 1 9 1 10 9 16 11 13 1 10 9 2 3 13 16 15 13 1 10 11 11 1 10 12 1 11 1 12 2
19 11 11 11 2 11 2 12 1 11 1 12 2 13 10 9 7 9 0 2
41 9 2 15 13 1 10 9 0 1 13 2 9 0 2 9 2 9 1 9 2 9 1 9 0 2 9 0 7 0 2 9 2 9 1 9 1 9 2 9 0 2
5 13 0 1 3 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
22 9 1 10 9 13 1 9 4 13 2 12 2 1 9 1 10 9 1 10 9 0 2
34 3 13 10 0 9 16 13 1 10 9 13 12 9 1 9 0 2 7 3 13 0 13 15 1 10 1 10 11 11 7 10 1 11 2
25 11 13 10 9 7 10 9 1 10 9 1 10 0 9 2 16 13 1 10 9 1 11 1 11 2
59 13 16 10 9 1 11 13 15 1 10 9 16 13 10 9 1 10 9 1 10 9 2 10 11 2 11 13 1 11 1 9 1 10 9 1 11 2 10 9 2 16 13 15 1 11 2 9 1 10 9 2 16 13 1 11 1 10 9 2
26 11 13 10 9 1 9 0 1 10 9 1 11 1 10 9 1 11 2 11 2 1 10 9 1 11 2
10 1 10 9 15 13 1 10 9 0 2
35 10 9 1 10 9 1 9 1 9 15 13 13 9 1 12 9 2 15 1 12 9 3 13 10 9 2 16 15 13 1 9 7 9 0 2
38 13 16 9 1 10 9 1 9 0 7 9 0 13 1 9 2 1 15 15 15 15 4 13 10 9 2 10 9 2 10 9 2 10 9 0 2 8 2
46 11 13 1 15 1 13 10 11 11 1 10 9 11 11 1 10 9 1 9 1 9 1 10 9 1 11 7 2 3 2 13 9 0 3 1 10 9 1 11 11 11 7 1 11 11 2
17 10 9 1 10 9 1 11 13 3 0 2 1 12 1 12 9 2
49 10 9 13 10 9 1 10 9 0 2 3 10 11 11 11 2 11 2 2 1 9 1 10 9 1 9 1 10 11 11 2 10 9 16 3 13 1 10 9 1 10 11 11 1 10 11 11 11 2
22 10 9 4 13 15 1 15 7 15 3 13 16 3 13 1 10 0 11 1 10 11 2
22 9 0 16 13 12 9 0 2 12 1 15 1 11 2 7 13 12 9 1 10 9 2
31 10 11 16 13 10 9 1 10 9 13 11 4 7 4 13 1 10 11 1 9 1 11 2 13 3 10 9 1 9 0 2
35 10 12 1 11 1 12 2 10 11 11 1 9 1 10 11 11 13 1 11 7 1 10 9 1 9 1 10 13 15 13 1 10 9 0 2
35 10 0 9 0 1 15 9 1 10 9 4 13 1 10 9 11 1 11 11 2 16 13 1 13 10 9 1 10 11 11 1 13 1 3 2
16 1 11 13 10 9 1 10 9 1 10 9 1 9 1 9 2
11 13 15 1 13 15 2 7 1 13 15 2
15 10 11 4 4 13 1 9 7 3 13 1 10 0 9 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
40 10 9 0 15 13 3 1 10 9 1 10 9 12 9 2 2 11 11 2 2 2 11 11 2 7 2 11 11 2 2 10 9 16 13 10 9 1 10 12 2
18 3 13 1 10 0 9 10 9 1 10 0 11 15 13 10 9 0 2
37 3 2 10 9 13 0 1 10 11 1 11 1 11 1 11 11 7 11 2 13 15 11 1 11 1 11 2 2 1 10 9 1 9 1 10 9 2
28 3 15 13 9 1 10 9 1 10 11 11 7 10 11 11 2 10 0 9 3 0 2 3 13 1 11 11 2
14 10 9 16 13 1 9 16 13 10 9 1 10 9 2
25 1 9 2 11 13 0 1 13 1 10 9 0 2 0 2 16 13 10 9 0 1 10 9 0 2
22 10 0 9 16 15 13 13 1 10 9 16 13 9 2 9 1 8 7 8 2 8 2
10 13 1 10 9 0 1 11 2 11 2
17 3 13 9 1 10 9 1 10 9 1 10 2 9 1 9 2 2
6 15 15 13 1 9 2
36 2 1 10 9 1 10 9 0 2 4 13 10 9 1 9 1 11 16 13 0 7 3 0 7 16 4 3 13 9 1 10 9 2 2 13 2
55 1 10 9 0 10 9 15 13 10 9 0 2 10 9 1 10 9 0 7 15 13 16 15 13 10 0 9 1 10 9 1 12 2 16 1 15 1 12 2 7 16 15 4 13 1 10 9 1 10 9 1 9 1 9 2
46 4 13 1 11 11 7 4 13 12 9 2 11 2 12 1 11 1 12 2 5 12 1 11 1 12 2 2 15 11 2 12 1 11 1 12 2 7 11 2 12 1 11 1 12 2 2
37 1 9 1 16 1 10 9 1 10 9 3 13 9 2 15 13 1 0 9 7 15 1 9 13 1 10 9 1 10 9 16 13 1 9 1 15 2
22 11 1 11 11 13 10 9 1 9 1 9 1 10 9 1 10 9 11 11 11 11 2
32 10 9 0 15 13 1 10 9 2 1 10 9 2 3 10 9 13 0 7 15 13 10 9 1 13 10 9 1 10 9 0 2
7 9 0 2 0 7 0 2
19 11 13 10 9 0 1 10 9 1 11 2 9 1 11 2 1 12 9 2
7 2 3 13 9 10 9 2
30 1 9 1 10 9 2 10 9 1 10 9 0 1 10 9 1 9 0 7 10 9 1 10 9 0 13 0 9 3 2
46 1 10 9 2 10 9 0 13 1 10 9 1 10 11 1 11 2 13 1 10 9 1 10 11 11 2 7 1 10 11 11 11 11 11 11 2 11 2 3 13 1 11 1 11 11 2
33 1 11 12 2 12 2 11 15 13 1 10 0 11 1 13 12 11 1 10 9 16 10 13 10 9 8 1 9 1 10 11 11 2
28 1 12 10 9 11 1 11 13 1 11 13 10 0 9 2 0 1 13 3 2 1 10 9 2 1 10 9 2
59 1 10 12 9 2 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
13 10 0 9 3 13 0 2 15 4 7 13 15 2
17 3 3 15 13 3 3 10 9 2 7 13 3 10 9 1 13 2
22 3 12 9 3 3 15 13 11 11 7 3 13 10 9 1 13 1 10 11 11 11 2
19 3 13 11 7 13 10 0 9 13 1 10 11 1 10 9 7 10 9 2
11 10 9 15 13 1 10 9 7 15 13 2
36 13 16 13 16 13 15 2 10 9 1 11 2 15 13 1 13 10 9 1 9 8 13 10 9 16 15 13 1 13 16 13 0 1 10 9 2
22 1 10 12 10 9 13 10 9 1 12 9 1 10 9 0 1 12 9 1 5 5 2
21 13 10 0 9 1 10 0 9 7 1 10 9 1 9 8 13 9 7 9 0 2
17 11 4 1 13 9 3 13 1 9 13 1 11 1 13 10 9 2
16 1 9 1 13 15 13 1 13 15 2 7 1 13 9 0 2
39 0 1 5 8 13 10 9 1 15 2 4 13 13 10 9 7 9 1 9 2 15 13 7 4 1 13 3 2 15 9 10 9 7 9 1 13 15 3 2
25 10 9 13 1 10 9 1 10 9 1 15 1 10 9 2 3 16 13 1 13 15 1 10 9 2
31 1 11 12 2 9 1 12 2 7 11 12 2 11 13 11 2 1 10 9 0 1 11 11 2 1 9 0 1 9 0 2
10 10 9 1 13 1 9 2 11 2 2
17 13 10 9 3 0 1 10 9 1 12 9 2 11 2 12 2 2
18 10 9 13 10 9 0 1 5 12 9 1 10 5 12 1 10 9 2
12 3 2 12 9 1 9 13 1 12 9 0 2
15 15 13 10 9 11 7 12 9 2 11 7 11 11 0 2
17 10 9 13 13 10 9 3 0 2 7 13 13 15 1 10 9 2
13 1 10 9 1 12 2 13 12 9 1 12 9 2
24 13 0 1 10 9 0 16 13 10 9 0 1 10 9 1 16 13 3 7 3 10 9 0 2
12 15 3 4 13 3 10 9 2 2 13 11 2
12 11 13 10 9 1 12 9 1 9 1 9 2
72 13 10 9 0 1 10 15 15 13 1 10 9 1 10 9 1 10 11 13 10 9 1 10 9 7 13 1 10 9 1 10 11 2 10 9 2 3 0 2 11 11 1 11 2 7 13 1 10 9 1 11 1 16 13 10 9 0 2 10 9 11 2 1 10 9 1 9 1 13 10 9 2
78 13 10 9 3 0 2 16 15 13 1 10 9 1 16 10 9 13 10 9 1 9 1 10 9 0 2 3 7 10 9 0 1 10 15 15 13 2 10 11 11 12 2 8 2 12 2 13 3 3 10 9 2 7 10 0 9 3 1 10 9 1 10 0 11 2 11 2 2 9 0 2 13 10 9 1 10 9 2
15 10 9 0 1 10 9 2 13 13 1 10 9 1 11 2
66 2 15 13 1 10 11 10 0 9 1 10 9 7 10 9 0 4 13 1 10 9 2 16 13 9 2 3 0 2 2 4 13 11 2 16 13 1 10 9 16 2 13 2 2 16 2 13 1 10 9 2 7 16 2 4 1 13 7 13 10 9 1 10 9 2 2
40 10 9 1 10 9 13 13 15 3 1 10 11 2 3 16 1 10 9 1 11 11 15 4 13 9 1 10 9 15 13 1 10 9 7 10 9 1 10 9 2
37 10 9 13 4 4 13 3 1 12 1 12 8 3 1 10 9 1 10 9 0 2 11 2 1 9 1 16 10 9 4 13 1 10 9 3 0 2
17 15 4 13 3 3 1 10 9 1 11 11 1 10 11 11 11 2
25 13 16 13 1 3 4 13 16 10 9 1 9 13 1 9 2 7 1 3 13 3 13 7 9 2
17 10 9 4 13 1 9 1 10 12 1 10 12 1 11 1 12 2
22 10 9 13 1 10 9 1 9 0 3 3 13 9 2 7 3 13 0 13 10 9 2
44 10 12 1 11 1 12 13 1 10 9 1 9 0 0 7 13 3 10 9 1 11 1 12 2 1 11 1 10 9 13 10 9 7 13 10 9 0 13 10 9 1 11 11 2
37 15 13 13 10 9 1 10 9 2 16 15 13 3 1 10 9 2 7 4 13 1 10 9 1 10 9 7 10 9 1 9 0 3 1 10 9 2
10 1 12 15 13 10 9 1 10 11 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
19 10 9 4 13 1 10 0 9 1 10 0 9 1 9 1 11 11 11 2
20 3 13 7 1 0 9 2 3 3 4 7 13 15 1 11 16 13 10 9 2
29 1 13 1 12 13 1 9 0 1 10 9 0 1 9 2 13 3 1 10 9 2 1 4 15 13 1 10 9 2
34 4 13 1 11 1 2 11 2 11 2 11 2 11 1 11 2 11 11 2 11 11 7 11 11 7 13 1 11 2 11 7 11 11 2
15 1 10 9 10 9 13 13 10 9 1 12 1 12 9 2
40 10 9 4 1 0 13 10 9 1 10 9 0 13 1 10 9 1 15 10 0 9 1 10 9 2 12 5 2 4 13 1 9 0 2 9 0 7 10 9 2
27 1 10 12 9 1 11 2 11 13 3 7 3 0 16 1 10 9 13 10 9 7 1 10 15 2 15 2
26 1 10 9 1 10 11 1 10 11 2 11 2 11 15 13 1 10 11 16 11 11 2 15 13 9 2
28 1 10 9 10 9 13 10 0 11 1 10 9 16 15 13 1 10 9 2 15 13 1 15 7 13 10 9 2
41 10 9 13 10 9 1 9 16 13 0 1 13 2 0 9 2 2 9 0 1 9 2 9 2 7 9 2 1 9 1 13 15 3 1 10 0 9 1 9 0 2
25 10 9 0 1 9 1 11 2 11 2 2 4 13 1 11 7 13 9 1 10 9 1 11 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
28 1 9 2 13 10 9 1 9 0 9 1 9 1 10 13 1 10 9 13 1 9 7 3 1 2 8 2 2
26 13 10 0 9 1 10 9 1 9 7 15 1 9 1 10 9 0 2 7 10 9 13 10 10 12 2
20 15 15 13 16 13 13 1 13 2 13 10 9 7 15 13 13 15 1 15 2
26 11 1 11 13 1 10 9 8 5 9 2 2 8 5 9 1 2 2 16 15 13 1 9 1 9 2
20 15 13 15 10 9 2 3 7 3 1 10 9 2 4 13 16 13 10 9 2
41 10 9 2 16 13 3 0 1 0 2 13 10 9 7 15 13 3 13 3 15 16 15 13 13 2 10 9 1 10 8 2 10 9 0 16 4 13 2 10 9 2
25 10 9 1 9 0 15 13 2 13 7 13 13 15 16 13 10 9 1 10 9 0 1 0 9 2
22 15 13 1 11 11 2 15 15 13 7 13 16 15 15 13 3 16 13 1 10 9 2
19 9 3 0 7 3 0 9 1 10 9 7 1 10 9 0 16 15 13 2
12 10 9 1 9 13 1 10 9 1 10 9 2
16 3 13 1 15 10 9 1 16 10 9 3 13 1 10 9 2
38 13 1 13 7 13 10 9 1 10 16 4 13 10 9 16 15 13 2 9 1 9 2 1 9 0 7 9 0 1 9 2 10 9 15 9 1 11 2
27 3 3 13 0 2 13 10 0 9 7 13 10 0 9 2 7 4 13 10 9 1 15 0 2 10 9 2
45 4 13 10 9 0 1 10 11 11 11 1 10 11 2 11 2 12 2 12 2 7 1 10 11 11 1 11 11 2 11 2 1 12 2 1 10 15 13 9 1 10 11 1 11 2
27 2 15 13 10 0 9 2 7 10 0 9 13 3 0 2 13 1 9 16 13 1 9 16 3 13 9 2
23 11 2 13 1 11 2 11 2 11 2 11 11 11 2 2 9 1 10 9 1 10 9 2
11 10 9 13 10 9 3 0 1 10 9 2
30 13 16 16 13 1 11 3 13 3 3 7 10 11 7 10 11 2 15 13 10 0 9 1 15 3 4 13 0 3 2
17 15 13 1 10 9 16 15 13 10 9 3 0 1 10 9 0 2
76 3 13 3 9 1 10 9 1 16 15 13 2 10 9 1 9 3 3 2 10 9 2 9 1 10 9 2 7 13 3 10 9 1 10 9 0 7 1 10 9 0 16 15 13 1 10 9 2 10 9 1 9 2 10 9 0 2 10 9 0 0 2 10 9 13 1 10 9 2 12 9 1 11 11 2 2
49 10 9 1 10 11 1 11 13 1 10 9 2 9 1 11 13 0 1 10 9 1 10 9 0 2 3 11 2 1 10 15 3 15 13 13 1 10 9 0 1 10 13 15 3 10 9 1 11 2
17 11 11 11 2 16 13 10 9 1 12 2 13 10 12 9 0 2
39 1 10 9 1 11 2 11 2 11 7 11 10 9 1 9 1 10 9 13 2 11 2 11 2 11 7 11 1 8 1 8 7 10 11 1 8 1 12 2
34 3 1 12 15 13 10 9 0 1 10 0 9 2 7 3 13 1 10 9 12 7 15 13 10 9 7 4 9 1 13 15 10 9 2
25 10 0 11 15 13 1 10 12 7 3 13 12 9 0 15 13 1 13 2 10 9 1 9 2 2
31 10 9 9 13 10 16 15 13 1 10 9 1 10 12 0 9 2 3 7 10 9 13 1 10 9 0 13 10 9 9 2
34 1 10 11 11 11 11 13 10 9 0 1 12 9 0 2 1 10 9 12 5 12 13 0 1 9 7 12 5 12 13 0 1 9 2
33 10 9 13 1 0 9 7 1 11 15 13 2 10 9 13 1 10 9 0 2 10 9 0 7 0 9 15 13 10 9 1 11 2
32 11 11 13 10 9 0 13 7 13 1 11 11 16 13 1 0 9 10 12 1 11 1 12 1 10 9 11 11 7 10 11 2
21 1 12 4 1 13 9 1 9 13 1 10 9 3 1 10 9 1 9 1 9 2
20 10 9 4 13 1 10 9 11 11 11 1 10 2 0 0 9 0 0 2 2
46 10 9 0 13 1 10 9 3 3 7 10 9 1 10 9 2 7 10 9 2 3 13 7 10 12 1 12 2 1 10 0 9 0 1 10 9 0 2 13 11 1 9 1 9 0 2
17 3 7 13 11 3 13 9 1 13 1 11 16 13 1 10 11 2
32 10 9 0 13 10 9 1 9 1 12 9 7 12 11 2 12 9 2 1 9 1 12 9 7 12 9 2 12 9 0 2 2
46 3 15 13 9 1 10 9 2 1 10 9 1 10 11 1 11 16 13 16 2 10 9 0 13 2 1 9 2 12 9 1 10 9 1 12 9 2 1 13 10 9 7 10 9 2 2
12 15 15 13 1 13 10 9 0 2 11 2 2
25 10 9 13 15 0 2 0 1 10 9 2 9 1 10 9 16 15 13 1 10 9 7 15 13 2
39 10 9 16 13 1 10 9 1 2 9 12 2 13 3 11 11 11 16 13 3 13 0 10 11 11 1 11 1 11 3 15 13 10 9 1 9 1 9 2
33 1 10 9 12 7 13 1 10 0 9 1 10 0 9 11 11 2 11 11 15 13 0 1 10 9 13 1 10 9 7 10 9 2
51 10 0 9 1 10 9 0 16 13 1 10 9 10 11 1 10 9 12 7 16 4 13 1 9 1 9 2 4 13 3 1 10 9 1 11 2 11 11 7 10 9 1 10 9 0 2 11 11 11 11 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
19 10 9 1 9 15 13 1 10 9 0 2 1 0 16 15 13 9 0 2
30 13 1 10 9 1 10 15 10 9 13 10 9 2 13 1 10 9 1 10 3 7 1 10 9 1 11 2 11 11 2
16 1 10 9 1 11 13 12 9 1 9 2 16 13 1 11 2
16 13 10 9 0 16 15 13 10 10 9 1 10 9 1 11 2
15 16 13 12 1 12 9 1 9 15 13 1 10 9 0 2
15 15 13 10 9 13 10 9 7 10 10 9 13 15 9 2
7 10 9 13 1 12 9 2
33 0 9 1 0 1 10 9 3 1 10 9 2 13 1 10 9 0 2 7 16 13 9 0 1 8 1 10 9 7 1 10 11 2
30 10 9 13 2 1 10 0 9 1 10 15 0 2 0 9 1 10 9 1 10 9 1 10 0 9 1 10 9 12 2
33 10 9 4 13 1 10 3 11 11 1 11 2 3 11 1 11 1 11 2 7 10 11 11 1 10 11 7 10 11 2 11 2 2
22 13 10 9 11 2 13 1 10 9 9 7 16 15 13 1 15 9 2 13 10 9 2
42 13 1 10 9 1 9 16 13 1 11 1 10 9 2 11 10 11 2 2 7 3 4 13 3 16 10 9 0 2 11 11 2 15 13 1 10 9 15 3 7 3 2
9 3 13 12 9 7 10 9 2 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
26 3 2 13 9 0 1 11 1 11 11 2 7 1 9 13 10 9 1 9 1 11 1 10 11 11 2
23 13 15 1 10 9 3 0 1 10 9 2 13 1 3 1 10 9 0 7 10 9 0 2
46 1 10 0 9 15 13 1 10 0 9 2 13 12 9 1 3 12 9 1 9 1 9 2 15 16 13 1 10 12 9 1 9 15 13 1 13 1 10 0 9 1 11 1 10 11 2
16 1 10 9 13 9 1 2 11 11 2 7 2 10 11 2 2
9 10 0 9 9 13 11 11 11 2
11 3 2 10 9 4 4 13 1 13 9 2
23 10 9 15 13 11 11 2 9 0 2 7 13 10 9 12 9 0 1 10 9 1 11 2
12 10 9 0 4 13 10 12 1 11 1 12 2
33 15 9 13 13 16 1 10 9 3 15 4 13 1 10 9 0 2 7 1 10 9 0 2 1 10 16 15 13 10 9 13 3 2
44 1 15 2 10 9 1 10 9 2 11 11 11 2 9 1 10 0 9 13 1 10 9 2 16 10 9 11 11 3 13 9 1 10 9 7 16 3 15 13 1 10 9 0 2
29 13 10 9 1 13 10 9 1 9 0 2 2 1 13 1 9 16 3 15 4 13 9 7 3 4 13 9 2 2
19 11 15 13 1 11 16 13 0 2 7 11 13 10 9 1 16 13 0 2
9 13 10 9 0 1 10 12 9 2
59 3 15 13 1 13 1 13 10 9 2 1 10 9 2 2 1 9 0 2 1 9 1 9 7 9 0 1 9 2 7 10 9 1 9 13 9 8 7 1 12 8 1 10 16 13 10 9 1 9 0 2 10 9 13 1 12 0 2 2
25 13 1 9 1 11 2 11 2 11 2 11 11 2 11 11 2 7 11 11 13 1 11 1 12 2
20 10 11 9 9 13 10 9 1 9 1 11 16 13 1 10 9 0 1 9 2
23 1 12 10 9 4 13 1 10 0 9 1 9 0 2 10 11 11 1 10 0 12 9 2
37 11 11 11 2 11 2 11 2 12 1 11 1 12 2 2 2 3 13 1 11 11 2 13 10 9 0 1 10 9 0 1 11 2 13 1 11 2
37 10 9 11 13 9 1 15 1 10 0 9 1 10 8 2 11 2 1 10 9 1 10 3 0 9 11 2 11 2 9 0 7 10 9 3 0 2
22 1 10 9 0 1 12 2 10 9 1 10 3 13 0 0 4 13 3 1 10 9 2
20 1 9 2 10 9 13 1 9 1 10 9 0 2 10 9 1 10 9 0 2
29 11 11 11 2 0 11 2 13 10 9 0 0 1 8 8 13 1 11 1 12 2 0 1 11 9 2 11 11 2
25 10 9 1 10 9 2 16 3 15 13 10 9 2 13 10 9 0 13 1 16 13 10 9 0 2
18 10 15 13 10 10 9 16 13 0 2 13 9 0 16 15 13 0 2
74 3 1 9 2 0 9 1 10 9 13 10 9 1 0 9 1 10 9 2 1 10 9 11 2 11 11 7 11 2 2 11 2 11 11 7 11 2 2 11 2 11 11 7 11 2 2 11 2 11 11 7 11 2 2 11 2 11 11 7 11 2 2 11 2 11 11 7 11 2 2 11 11 2 8
58 10 9 4 13 2 3 1 9 0 2 1 10 9 2 1 10 11 11 1 11 2 13 1 11 1 11 7 11 2 16 13 10 10 9 1 10 0 11 11 2 1 10 9 9 1 10 11 1 10 11 2 15 10 9 13 4 13 2
30 15 13 13 10 9 1 9 0 2 3 0 2 13 1 13 3 9 13 3 1 9 0 2 13 10 9 1 10 9 2
21 13 10 9 1 11 7 10 0 9 1 9 2 11 8 11 2 11 2 12 2 2
34 1 10 9 3 1 10 9 13 2 10 9 3 4 13 0 2 1 10 9 4 1 13 3 9 1 13 10 9 1 3 9 7 9 2
7 3 8 10 9 1 15 2
28 3 13 1 15 1 10 9 1 10 9 2 13 0 1 15 10 9 2 10 11 1 10 11 2 0 1 11 2
32 1 9 1 16 10 9 1 11 13 10 0 9 1 10 9 2 10 9 4 13 1 12 1 10 9 1 10 11 11 1 11 2
5 15 13 1 11 2
22 13 13 2 15 3 13 10 9 0 1 10 9 11 2 16 4 7 13 3 15 13 2
21 10 9 1 10 9 3 3 15 13 2 13 16 1 15 1 10 9 0 2 0 2
29 10 12 1 11 1 12 2 13 1 10 11 11 11 1 10 9 1 10 0 9 9 1 10 11 8 8 1 11 2
17 13 1 10 9 13 11 13 1 10 9 1 11 2 11 2 11 2
16 10 9 13 3 10 9 7 13 10 9 0 1 10 9 0 2
5 15 13 1 11 2
20 11 13 16 10 9 13 0 1 10 9 1 10 9 2 7 13 1 15 0 2
20 10 9 1 11 4 13 1 10 11 7 10 9 1 13 9 1 10 9 0 2
5 10 9 13 3 2
47 1 10 9 10 9 3 0 13 10 9 2 16 1 10 0 9 1 9 13 4 13 2 3 1 13 3 3 10 9 7 13 0 9 16 15 13 13 0 9 16 13 1 10 9 1 9 2
50 1 12 2 10 9 1 11 2 11 4 4 13 1 2 9 2 1 12 9 1 10 9 1 9 0 2 11 2 11 11 11 2 3 1 10 9 13 0 2 16 13 10 9 1 10 9 1 12 9 2
27 10 9 1 9 0 13 15 9 0 7 0 7 8 2 3 16 10 9 0 13 3 10 9 1 10 9 2
35 7 15 3 9 1 9 2 10 9 1 10 9 2 16 3 1 10 9 16 15 13 3 2 15 4 1 13 7 13 10 9 1 10 9 2
23 11 11 13 10 9 0 16 13 11 11 2 11 8 11 8 11 11 2 1 12 7 12 2
4 13 10 9 5
26 10 9 15 13 1 12 9 1 16 10 9 4 13 2 3 10 9 1 10 12 1 9 1 10 9 2
23 15 4 13 9 1 0 9 1 11 11 2 11 7 11 11 11 1 13 15 10 9 0 2
20 13 16 11 13 10 0 9 0 0 2 15 13 1 15 1 10 9 3 0 2
78 10 9 1 9 13 10 0 9 1 9 2 10 9 0 2 13 1 10 9 1 10 9 2 4 13 15 2 1 10 10 10 9 7 1 10 15 15 15 15 13 7 13 16 15 13 0 7 0 1 13 2 2 9 16 4 13 13 10 9 2 13 10 9 2 13 10 9 2 13 10 9 7 13 9 1 10 9 2
43 1 15 2 10 9 1 10 9 13 13 10 9 0 7 1 11 1 10 11 2 11 1 11 2 2 13 1 12 3 1 10 9 7 1 10 1 11 2 11 1 11 2 2
29 13 1 12 9 1 10 11 1 11 1 10 11 1 11 1 11 2 1 10 15 13 12 9 7 12 9 1 9 2
7 10 9 13 10 9 0 2
32 10 9 0 13 1 2 13 10 9 0 2 0 2 0 2 0 2 0 2 0 2 16 13 7 13 10 9 7 10 9 2 2
12 1 9 13 1 10 11 7 10 9 1 9 2
22 1 9 1 13 1 10 9 2 15 4 13 1 10 9 1 10 9 0 1 10 9 2
37 10 9 13 10 9 1 0 9 0 1 9 1 9 1 12 2 7 3 1 10 0 9 1 9 1 9 2 1 12 9 1 9 13 10 0 9 2
36 3 13 10 9 1 9 13 1 10 9 1 9 8 2 15 16 13 1 10 9 16 13 1 10 9 1 10 11 11 2 12 9 1 12 13 2
9 1 10 9 2 10 9 4 13 2
43 13 1 10 9 1 10 9 1 11 10 12 1 11 1 12 2 13 1 9 1 10 11 11 1 11 1 12 7 13 10 9 1 11 1 11 1 10 11 11 11 1 11 2
14 1 10 9 1 9 0 2 15 15 13 2 9 2 2
28 10 9 13 10 9 2 11 1 10 11 2 1 10 9 1 9 11 11 11 11 7 13 9 1 10 9 11 2
24 11 13 1 11 15 1 11 7 11 13 13 15 1 15 2 15 13 10 9 7 13 10 9 2
52 1 9 9 2 11 13 0 3 1 9 8 9 1 10 9 0 1 11 7 11 2 13 10 9 0 1 13 15 1 10 9 1 9 1 10 0 9 2 13 15 1 10 9 1 10 0 9 1 10 9 0 2
13 10 9 13 1 10 9 1 11 2 9 1 11 2
32 10 9 1 9 3 13 3 0 2 3 7 15 4 1 13 1 9 1 10 9 7 15 4 1 13 1 10 8 1 10 9 2
3 2 9 2
29 1 10 9 1 10 9 1 10 9 1 10 0 9 2 10 9 13 10 9 0 2 12 9 0 1 11 1 12 2
22 1 10 0 9 11 13 10 0 9 13 1 10 9 12 16 15 13 3 1 10 9 2
49 10 9 13 10 9 7 3 10 9 4 13 1 15 1 10 9 1 10 9 0 2 1 10 0 9 1 11 1 10 9 1 10 9 1 10 9 1 11 11 1 15 1 10 0 9 1 10 9 2
53 3 2 11 11 4 13 16 1 10 9 1 9 10 9 13 15 7 1 0 9 16 0 13 13 0 1 13 15 1 10 9 13 1 10 9 0 2 1 10 9 1 16 10 9 15 13 7 10 9 13 1 13 2
26 13 1 3 13 1 10 9 2 15 13 1 13 10 9 1 10 9 0 1 9 16 3 15 13 0 2
23 1 16 13 1 10 9 2 13 15 3 0 1 3 1 10 9 0 7 0 1 10 9 2
18 1 10 0 9 13 10 9 1 11 2 11 2 11 11 7 11 11 2
20 13 1 12 7 12 1 11 11 11 2 15 13 1 12 9 13 1 9 0 2
25 13 10 9 0 1 10 11 11 2 3 13 3 10 12 5 1 10 9 16 15 13 1 10 9 2
24 1 10 9 15 4 1 13 7 1 9 10 15 4 13 1 13 1 11 7 13 0 1 15 2
30 3 13 16 10 9 4 13 1 9 1 10 9 1 10 11 1 11 11 1 11 2 10 15 13 0 1 10 11 0 2
17 10 9 2 2 11 2 2 4 13 1 10 9 1 10 9 12 2
45 10 9 11 11 2 12 2 12 1 0 9 1 9 2 8 2 15 13 1 10 0 9 0 16 13 10 9 2 13 12 9 7 13 10 9 0 1 12 9 1 9 1 10 9 2
25 15 13 10 9 1 10 9 7 9 2 3 1 10 9 1 10 9 7 13 3 0 3 4 13 2
72 10 9 12 1 10 9 1 9 1 15 9 7 9 13 10 9 1 10 9 11 7 11 11 2 9 1 5 2 1 10 13 15 1 4 13 1 12 9 10 9 12 9 2 9 2 1 10 9 8 5 12 16 13 10 9 0 2 1 4 13 15 1 10 9 15 4 13 3 1 10 9 2
11 1 10 9 4 13 1 10 9 1 9 2
22 11 1 9 1 10 11 11 1 12 9 2 4 1 13 1 11 11 7 1 11 11 2
21 10 9 1 10 9 13 13 10 9 1 9 9 1 10 0 9 13 1 10 9 2
17 1 10 9 10 9 0 15 13 3 1 10 9 1 10 11 11 2
29 1 11 1 12 1 12 2 10 11 13 1 11 7 10 11 9 1 9 2 9 2 9 2 7 9 1 10 9 2
31 3 1 10 0 9 1 10 9 2 15 9 13 2 16 13 1 11 7 11 11 2 16 10 9 13 9 0 1 10 9 2
10 11 11 1 10 9 0 1 10 9 2
43 10 9 15 13 1 10 0 9 0 1 9 1 10 9 0 2 7 15 13 3 0 1 10 9 7 13 3 10 9 1 10 9 1 16 11 4 13 1 10 9 1 9 2
16 10 9 13 10 9 16 13 1 10 10 9 1 13 10 9 2
13 13 1 11 2 11 2 10 12 1 11 1 12 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
11 13 13 10 12 9 1 10 9 1 11 2
7 13 1 9 1 10 9 2
8 3 3 13 9 7 9 0 2
6 13 15 9 3 13 2
16 3 1 10 9 12 2 10 9 1 10 9 13 10 9 0 2
22 13 13 15 9 1 10 9 0 1 10 15 10 9 2 11 11 2 4 4 7 13 2
41 10 9 1 10 9 0 13 10 9 1 1 10 9 2 13 16 10 9 0 13 10 12 5 1 10 9 1 10 9 1 9 7 10 12 5 1 10 9 1 9 2
8 1 11 10 9 4 13 1 2
16 13 2 1 9 1 9 2 15 13 1 10 9 1 10 9 2
28 10 9 15 13 3 16 13 1 11 1 10 9 1 9 0 2 1 15 15 13 1 10 9 11 1 10 9 2
10 13 9 0 13 1 11 1 10 9 2
10 7 3 13 1 9 1 10 9 0 2
11 15 13 1 12 9 9 1 10 11 11 2
15 1 10 9 2 10 9 3 13 9 1 9 1 15 0 2
10 10 9 0 13 10 0 12 1 9 2
44 3 2 10 9 1 11 15 4 13 1 10 0 9 1 9 1 10 0 9 0 7 0 13 1 10 9 2 3 16 15 13 1 9 1 10 0 9 0 1 10 9 1 11 2
40 10 11 1 11 7 10 9 1 11 13 10 9 1 9 7 9 1 9 1 9 7 1 10 9 2 16 13 10 0 9 1 9 0 1 10 9 7 10 9 2
26 10 9 8 13 0 1 10 9 0 2 7 1 9 10 9 0 1 10 9 0 7 10 0 9 0 2
25 10 9 16 10 9 16 15 4 13 2 15 13 1 10 9 2 3 13 16 13 0 1 10 9 2
25 13 1 10 9 2 10 0 9 15 13 1 13 1 9 7 4 13 13 1 10 0 9 13 11 2
32 10 9 3 4 4 13 1 10 11 11 2 13 0 2 1 10 9 11 2 9 1 9 2 13 1 10 9 0 1 10 9 2
22 15 13 13 15 3 9 16 3 13 13 9 2 7 13 0 15 9 16 13 10 9 2
36 10 9 1 9 7 9 1 9 0 1 9 0 7 0 2 15 13 1 10 9 2 10 9 2 9 2 7 1 10 9 1 10 2 9 2 2
61 11 11 13 1 10 9 15 13 2 0 7 0 2 7 10 13 3 1 10 12 9 15 0 1 13 10 9 2 13 16 10 9 0 1 11 3 13 1 10 9 1 9 2 7 3 15 13 1 10 9 1 10 9 9 1 10 9 1 9 0 2
47 1 11 7 1 9 2 16 15 13 2 10 9 2 10 9 7 13 1 15 13 7 1 15 3 2 1 10 9 1 10 11 7 10 9 1 10 11 2 1 16 10 9 15 13 16 13 2
29 1 10 9 2 10 9 3 10 9 13 10 9 13 1 9 1 9 1 10 9 1 10 9 13 1 9 1 9 2
24 13 10 9 10 9 1 2 11 11 2 7 10 12 0 9 1 9 0 3 13 0 1 15 2
8 15 13 1 11 7 10 11 2
16 13 0 2 16 13 10 9 1 11 11 1 11 11 1 12 2
28 13 1 12 7 13 1 0 9 1 11 11 1 12 2 10 9 1 10 9 4 13 1 11 11 11 1 12 2
17 10 9 0 1 10 11 13 1 9 1 10 9 13 1 10 9 2
5 10 9 13 0 2
41 10 9 1 9 0 2 0 4 4 13 7 13 1 9 0 2 1 10 8 0 2 7 1 9 0 2 1 10 9 13 1 9 0 7 10 9 0 8 8 2 2
22 13 3 10 9 1 10 9 0 1 11 2 1 10 15 15 13 9 1 11 7 11 2
40 15 13 2 15 15 13 1 10 0 9 2 13 1 9 2 3 0 7 3 3 3 1 10 9 7 10 9 2 15 4 13 13 1 10 10 9 1 10 9 2
29 13 3 1 10 11 10 9 1 10 9 1 10 9 1 10 9 0 13 11 11 11 2 1 9 1 13 10 9 2
21 15 13 1 10 12 1 10 11 1 11 1 10 9 2 10 9 0 1 10 9 2
19 11 4 13 2 10 9 0 7 10 0 9 8 2 0 13 1 9 0 2
36 13 10 9 0 10 9 0 1 10 9 7 10 9 1 10 11 2 3 7 1 10 9 0 7 10 9 16 4 13 1 15 9 1 10 9 2
13 11 1 10 9 2 11 1 10 9 2 7 11 2
26 13 1 10 9 1 10 9 2 11 13 9 0 1 12 1 10 0 9 0 2 11 2 11 7 11 2
59 1 10 12 9 2 11 13 0 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
17 10 11 11 11 13 10 9 11 11 13 7 13 1 11 1 12 2
3 13 0 2
9 1 3 0 13 1 10 9 0 2
76 1 10 0 9 1 10 9 1 11 1 11 2 11 11 2 8 1 11 1 11 11 11 2 13 16 16 13 10 9 1 10 9 1 10 9 9 0 4 13 1 10 9 1 10 9 0 1 9 1 11 1 10 9 1 9 1 9 0 0 16 13 13 10 9 1 9 7 13 10 0 9 1 10 10 9 2
18 2 1 10 9 0 15 13 10 9 3 3 0 7 0 2 10 9 2
33 10 9 15 13 1 9 1 10 9 1 12 1 11 7 13 10 9 13 1 10 9 11 0 1 10 1 9 1 11 11 7 11 2
53 10 9 1 13 10 11 2 12 11 4 13 1 12 1 10 9 1 13 10 9 16 13 10 9 1 9 1 9 1 10 11 11 2 12 7 10 9 11 1 10 1 11 11 11 2 12 11 7 11 2 12 11 2
27 11 11 13 10 0 9 1 11 11 11 2 12 2 2 1 11 11 1 11 2 7 10 9 2 11 11 2
17 10 9 15 13 1 10 9 11 2 3 10 9 0 7 15 0 2
29 1 10 9 15 13 10 10 9 16 10 9 0 1 10 9 13 1 9 0 7 16 3 1 10 9 4 1 13 2
8 13 15 15 4 13 1 15 2
18 10 9 1 9 7 9 4 13 10 9 3 13 1 10 0 9 0 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
18 1 13 1 9 15 13 1 10 9 11 3 15 13 11 7 11 11 2
18 9 2 13 10 9 7 3 13 2 15 4 13 1 9 0 1 9 2
14 3 4 4 13 10 9 11 10 12 1 11 1 12 2
65 1 10 9 2 4 4 13 1 9 10 9 16 13 10 9 0 1 9 1 10 9 1 9 0 2 15 16 13 13 10 9 1 9 0 7 15 13 1 10 9 1 10 11 2 12 2 3 7 15 1 10 9 1 10 9 1 10 9 2 1 10 9 1 11 2
60 10 11 13 1 9 9 1 13 9 0 1 10 11 11 2 1 11 1 10 11 2 1 10 9 1 9 1 10 11 2 11 11 2 11 2 9 11 11 2 11 2 11 7 11 2 2 1 11 2 1 11 2 1 11 7 1 10 11 11 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
16 11 13 16 10 9 1 11 3 13 10 2 9 9 2 0 2
21 10 9 15 4 13 1 10 9 1 9 1 10 9 1 10 9 0 1 10 9 2
17 13 10 9 1 10 9 10 9 1 9 1 11 11 11 11 11 2
24 11 13 1 12 10 0 9 1 10 9 1 10 0 11 0 2 1 10 12 5 9 1 12 2
19 10 11 1 11 2 7 1 0 11 2 4 13 1 10 9 1 10 9 2
13 11 13 10 9 1 9 0 7 13 1 10 9 2
9 10 9 1 11 13 1 12 9 2
23 11 11 2 8 11 2 12 1 11 1 12 2 13 10 9 1 9 2 9 7 9 0 2
26 3 10 9 0 3 15 4 13 1 10 9 1 10 0 9 11 11 2 16 3 13 10 9 1 9 2
20 0 9 0 13 10 9 11 11 2 15 13 1 10 9 1 11 12 1 11 2
15 1 9 4 13 10 9 1 10 16 15 4 13 1 9 2
10 3 4 1 13 10 9 1 10 9 2
13 10 9 15 13 1 11 1 12 1 10 9 0 2
33 7 2 1 9 1 9 1 10 9 2 10 9 4 13 10 2 9 1 9 2 3 13 10 9 3 0 1 10 9 7 10 9 2
21 13 3 10 9 0 1 10 9 7 10 9 13 10 9 1 10 9 1 10 9 2
32 4 13 10 9 16 13 15 10 9 1 10 9 10 9 1 10 9 2 7 4 1 13 16 10 9 2 9 2 13 3 3 2
31 11 11 11 2 11 2 2 12 1 11 1 12 2 11 2 11 2 12 1 11 1 12 2 11 13 10 9 2 9 0 2
18 11 13 1 11 7 13 0 9 1 10 9 1 11 2 13 1 12 2
59 10 11 1 11 2 1 9 2 11 8 2 7 11 1 11 2 1 9 2 8 8 11 2 15 13 1 10 9 11 12 1 11 7 10 9 1 10 11 1 11 11 11 10 12 1 11 1 12 2 1 10 9 1 11 2 0 11 2 2
28 13 11 11 1 11 2 9 1 10 9 11 11 7 11 2 11 11 4 13 1 10 9 16 13 10 9 0 2
16 1 10 0 9 4 13 1 10 0 9 1 10 11 11 11 2
27 1 12 1 12 11 11 13 1 10 11 1 11 1 9 1 9 0 2 9 1 10 15 13 1 11 11 2
17 13 3 10 9 0 2 1 9 8 2 7 10 12 9 3 0 2
31 10 9 16 10 9 1 11 13 10 9 1 10 9 0 7 1 10 9 0 13 10 0 9 1 9 3 0 1 10 9 2
21 1 10 9 1 10 9 2 11 13 10 9 1 10 9 1 11 2 11 11 11 2
32 13 10 9 11 2 13 10 9 11 7 2 1 13 15 1 11 2 13 1 10 9 1 11 2 11 7 10 9 1 11 11 2
23 15 13 13 1 9 1 10 0 9 7 10 11 13 15 1 15 1 13 1 10 11 11 2
48 16 1 15 15 13 16 15 13 1 15 2 15 4 13 10 9 1 9 1 15 13 0 1 16 13 0 16 3 4 13 10 9 1 10 9 1 10 9 1 9 2 9 16 1 15 15 13 2
27 3 2 10 9 4 1 4 13 2 16 3 3 4 13 1 0 9 13 1 10 9 1 9 0 1 11 2
30 10 2 11 1 10 11 11 2 3 13 2 10 11 1 10 11 2 2 13 1 10 9 12 13 10 0 9 1 11 2
34 3 13 15 1 10 9 2 11 2 1 12 9 2 4 13 1 10 12 9 2 2 10 9 3 1 3 1 10 9 1 10 9 2 2
36 1 10 9 1 11 15 13 8 1 9 1 10 8 1 9 2 1 7 15 13 10 9 2 3 7 3 12 9 3 1 10 9 0 1 13 2
4 13 15 0 2
30 3 15 13 10 9 1 10 9 1 11 7 11 7 10 9 1 11 7 11 11 7 11 1 10 9 1 11 7 11 2
38 12 13 10 9 1 9 1 10 9 12 13 1 11 2 11 2 11 2 3 13 10 9 0 1 10 9 3 3 15 13 2 8 2 13 1 10 9 2
72 9 1 12 9 13 1 10 11 1 10 11 11 2 10 0 9 0 1 11 15 13 1 15 9 1 10 11 11 2 1 9 1 10 9 1 9 2 13 13 12 9 1 9 2 10 9 1 3 12 9 1 9 13 3 1 9 10 9 1 10 11 1 11 2 7 1 10 9 1 12 8 2
31 10 0 11 15 4 13 15 2 13 1 10 9 1 9 1 10 9 2 4 13 10 9 0 7 10 9 0 1 10 9 2
45 16 4 13 2 15 15 4 13 1 10 9 7 15 4 13 16 13 9 1 10 9 16 4 7 13 15 7 16 16 13 10 12 1 10 9 1 10 12 3 13 3 16 13 15 2
15 4 13 1 12 1 10 11 11 1 11 1 10 9 9 2
42 10 9 13 1 10 9 0 1 10 9 1 10 9 1 12 2 16 4 13 1 10 9 0 1 11 7 11 7 10 9 1 10 9 0 2 16 4 13 10 9 0 2
60 1 10 12 9 2 11 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
31 10 9 1 9 13 1 12 13 9 1 12 2 3 10 10 9 0 13 1 10 0 9 2 12 9 1 10 9 1 11 2
47 1 10 0 7 0 9 1 11 11 10 11 1 10 11 2 9 1 10 9 1 10 11 13 1 10 9 1 10 11 1 13 15 1 10 9 2 1 13 15 9 7 13 15 1 9 0 2
40 10 9 15 13 3 0 7 10 9 0 1 10 9 0 2 13 3 1 10 0 9 1 9 1 15 9 1 10 9 7 1 10 0 9 1 10 9 2 11 2
49 13 0 16 10 9 4 13 1 11 12 1 11 2 3 16 10 9 0 1 11 15 13 3 3 1 10 9 1 10 9 1 10 9 13 3 1 10 9 1 11 7 1 10 9 1 13 9 0 2
14 13 16 10 9 1 9 15 4 13 10 9 3 0 2
23 0 2 13 1 10 9 16 3 1 13 10 9 15 13 1 3 2 7 13 1 11 11 2
14 4 13 1 12 7 13 9 1 10 9 0 0 11 2
58 10 3 9 1 10 0 13 10 9 2 11 12 1 11 2 10 15 13 13 1 10 9 1 10 9 1 10 0 9 2 7 10 0 11 12 1 11 2 10 9 1 2 11 1 11 2 11 8 13 0 3 1 13 1 10 9 0 2
47 10 0 9 1 9 15 13 13 9 1 10 11 1 11 11 13 1 10 9 0 1 10 11 11 2 13 1 10 9 1 9 1 10 9 1 11 2 11 7 1 9 1 10 9 1 11 2
18 4 7 13 10 9 1 10 9 2 3 13 15 13 7 3 15 13 2
16 10 9 13 3 1 10 9 7 13 9 0 1 10 11 11 2
17 10 12 1 11 10 0 15 11 15 13 1 11 16 13 10 9 2
33 15 1 10 9 13 10 9 7 10 9 1 9 1 11 2 3 1 10 9 7 10 9 2 2 13 10 9 1 9 1 9 9 2
61 7 13 3 10 9 16 1 15 15 13 16 10 11 1 11 3 13 10 9 7 15 3 10 9 1 10 9 0 1 9 1 13 10 9 1 13 9 1 10 9 7 13 1 10 9 16 13 4 1 9 3 13 15 0 7 1 4 13 0 9 2
13 1 9 2 10 9 13 1 10 9 11 7 11 2
23 1 10 9 3 15 13 1 10 9 0 1 10 9 1 10 9 16 15 13 1 10 9 2
14 11 15 13 1 10 9 7 13 1 12 1 10 9 2
8 13 11 11 10 9 11 11 2
35 3 15 13 1 10 9 1 11 11 1 11 2 7 1 11 12 1 10 11 2 3 10 9 0 13 10 9 1 10 9 13 1 10 11 2
22 10 9 15 13 1 13 3 10 12 1 11 1 12 2 1 10 9 9 0 1 11 2
27 10 9 0 1 10 11 13 10 9 1 10 9 0 1 11 11 2 16 13 16 13 13 2 13 9 2 2
19 11 11 11 2 13 10 9 3 13 1 13 1 11 11 1 11 7 11 2
15 10 9 1 11 4 4 13 7 10 9 13 10 9 9 2
23 3 15 13 1 9 1 11 2 16 10 0 7 0 11 13 3 3 15 9 1 10 9 2
23 1 3 16 1 10 9 1 10 9 2 10 9 13 1 9 2 9 1 10 9 11 9 2
18 3 15 13 1 10 9 0 11 1 10 9 16 13 3 1 10 9 2
20 10 9 8 1 0 13 9 1 13 1 10 9 2 10 9 7 10 9 0 2
27 2 11 1 11 2 13 10 9 1 10 9 0 1 11 10 11 2 13 1 10 9 7 0 9 11 11 2
24 1 10 12 1 11 1 12 2 11 11 2 10 9 0 0 3 0 1 11 2 13 12 9 2
16 10 9 11 13 16 10 9 15 4 13 1 10 13 10 9 2
39 10 9 13 10 9 1 9 1 10 9 0 1 10 9 1 3 9 1 4 13 1 10 9 7 3 16 10 9 13 1 9 0 16 15 13 1 9 0 2
27 3 11 12 13 13 11 1 13 15 2 7 13 11 1 12 16 15 13 1 9 0 1 10 11 1 11 2
7 10 9 13 1 9 0 2
27 1 12 2 10 11 11 1 10 11 13 10 0 9 1 10 0 9 1 10 9 1 10 9 1 10 9 2
16 15 4 13 9 13 1 15 1 11 11 7 10 11 1 11 2
25 11 13 16 10 9 1 9 13 9 1 9 16 13 3 0 1 10 9 1 10 9 1 9 0 2
29 15 13 16 2 1 10 9 1 11 2 10 9 15 13 1 13 10 9 1 10 9 1 10 9 1 10 0 9 2
26 10 9 1 10 9 13 11 11 7 10 9 2 11 11 2 15 13 1 10 9 1 10 9 1 9 2
28 13 3 10 9 10 16 15 13 9 1 9 0 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2
25 10 9 11 11 13 10 9 16 10 9 1 10 9 1 10 9 0 2 3 15 4 13 3 2 2
7 13 1 0 2 4 13 2
30 10 11 0 16 13 12 9 1 10 9 4 13 1 11 2 11 11 2 11 7 10 11 11 10 12 1 11 1 12 2
9 13 3 0 7 13 1 9 0 2
39 3 2 1 12 10 9 13 1 4 13 1 9 0 7 16 10 9 3 10 9 15 13 1 10 9 13 2 11 15 11 11 2 2 10 9 13 10 9 2
15 1 10 0 9 13 3 13 1 10 0 9 11 2 11 2
27 1 9 1 10 0 9 1 9 2 4 13 1 10 9 1 9 1 10 9 0 1 10 9 2 11 11 2
20 11 11 2 10 11 1 11 2 13 10 9 0 9 1 10 9 1 10 11 2
34 10 9 1 9 4 13 1 13 10 9 0 9 1 10 9 1 9 0 13 2 9 1 9 1 0 9 0 7 1 3 9 1 9 2
27 1 10 9 1 11 11 13 3 1 10 9 1 0 7 0 9 2 1 10 9 1 11 2 11 7 11 2
30 10 11 1 11 13 10 9 1 11 1 12 2 1 15 15 15 13 1 10 0 9 0 13 1 11 1 10 9 12 2
8 3 4 13 15 1 4 13 2
23 10 0 9 0 1 10 9 0 15 13 1 12 7 13 1 10 9 0 0 1 10 9 2
20 16 13 9 0 7 15 13 9 15 3 1 9 2 15 13 1 10 0 9 2
24 10 9 13 10 0 9 1 9 1 10 9 1 9 16 15 4 13 1 10 9 0 1 11 2
38 10 9 1 11 11 13 10 9 1 10 9 1 10 0 9 1 9 7 9 2 1 10 9 1 9 7 9 2 13 7 13 15 1 9 7 9 0 2
47 10 9 1 10 9 12 1 11 11 13 16 2 10 9 13 10 9 1 9 2 13 10 9 16 15 4 13 1 10 9 16 3 4 13 1 9 7 10 9 16 15 13 1 10 9 2 2
15 15 13 1 11 1 10 12 7 1 10 9 13 12 9 2
15 15 9 13 16 11 11 13 10 9 0 1 12 9 0 2
11 11 11 2 1 9 2 13 0 10 9 2
38 13 16 15 13 0 1 16 15 4 13 13 10 9 1 10 9 1 10 9 7 13 15 1 10 9 2 1 15 1 10 9 16 11 13 1 10 9 2
35 10 9 4 13 10 9 1 12 9 1 10 9 11 11 2 1 9 8 7 8 7 1 0 9 2 9 0 7 0 1 10 12 8 2 2
18 1 13 1 11 3 1 9 7 3 3 1 10 4 13 2 11 13 2
19 13 10 9 16 15 13 1 10 9 1 10 2 9 1 10 0 9 2 2
43 16 11 13 2 11 13 10 9 1 10 9 1 13 10 9 0 2 1 15 1 10 9 13 1 10 11 2 9 1 10 0 9 2 2 7 0 2 13 1 13 10 9 2
22 10 9 11 13 10 9 13 1 10 9 1 10 9 1 10 9 0 1 10 0 9 2
20 1 12 10 11 13 10 9 1 10 9 9 12 12 2 1 10 9 11 12 2
28 10 9 13 0 7 10 9 1 10 9 3 3 0 2 15 13 11 2 15 13 10 9 7 15 13 10 9 2
20 10 9 1 10 9 3 13 0 2 16 13 9 16 3 13 10 9 1 15 2
25 11 3 13 1 15 0 3 7 1 15 3 2 13 3 0 2 10 9 1 10 9 1 11 11 2
38 10 12 1 11 13 10 9 1 10 9 11 11 7 10 9 1 10 9 1 13 15 1 10 9 1 11 11 2 16 3 13 10 9 10 12 1 11 2
41 1 13 1 10 9 1 10 9 11 2 13 10 9 1 9 7 13 1 9 1 10 9 11 2 11 11 12 2 10 15 4 13 1 9 1 9 1 10 3 13 2
16 10 9 13 10 9 0 1 5 12 1 5 12 1 10 9 2
31 10 9 1 10 9 15 13 1 10 0 9 1 10 12 2 1 12 9 2 13 1 0 9 1 10 9 1 10 9 11 2
37 1 9 2 1 10 9 1 10 9 1 10 9 0 0 4 4 3 13 2 10 9 0 4 13 1 9 7 2 1 0 9 2 4 4 3 13 2
17 16 10 9 15 13 4 13 10 9 3 7 13 10 9 1 9 2
23 1 10 9 10 9 1 10 9 2 15 4 13 1 10 9 0 1 10 9 1 10 9 2
33 13 3 1 10 9 1 9 7 9 3 0 13 1 11 11 1 10 11 12 2 13 9 1 11 11 2 11 11 7 11 11 11 2
32 1 13 16 10 9 0 3 15 13 2 15 13 1 12 9 9 0 2 12 1 10 9 7 10 10 12 10 12 1 10 9 2
34 10 9 1 13 1 11 11 11 1 10 9 1 12 2 1 10 9 13 9 0 16 13 13 10 9 1 10 9 2 3 13 1 11 2
38 9 3 0 13 9 1 9 2 0 1 9 1 9 7 9 0 2 9 1 9 1 9 1 9 0 1 9 1 0 9 0 7 9 1 9 1 9 2
32 10 9 3 3 2 16 11 13 9 1 11 2 12 2 12 2 2 11 15 13 1 10 9 0 7 3 1 9 1 11 11 2
18 3 2 13 1 10 0 9 1 9 2 9 7 9 1 10 11 11 2
30 3 3 10 9 3 15 13 10 9 2 1 10 15 4 1 13 10 9 0 2 10 9 1 9 2 1 12 1 12 2
34 11 7 11 1 10 11 13 10 9 1 10 9 1 11 2 13 1 10 8 1 10 9 2 1 10 9 2 7 1 10 11 1 11 2
18 1 15 15 15 13 16 15 15 13 1 3 3 10 12 12 9 0 2
23 7 11 11 13 16 11 3 13 10 9 1 13 16 13 10 9 1 9 1 10 9 11 2
49 0 1 10 9 2 10 9 4 13 10 0 9 0 2 9 1 10 9 1 9 1 9 0 1 12 9 2 1 10 9 1 1 10 3 10 12 1 12 1 10 9 2 1 9 0 7 0 2 2
33 13 10 9 15 13 16 13 10 9 2 1 10 9 11 1 10 9 11 2 13 1 10 9 11 7 11 7 11 2 9 1 11 2
41 10 0 9 13 10 9 10 9 0 13 1 15 1 10 9 1 9 1 11 13 1 11 11 2 10 9 16 3 4 2 13 2 1 11 1 10 11 11 11 2 2
16 1 9 2 8 9 7 8 0 2 16 13 9 1 10 9 2
18 10 9 13 10 9 0 7 0 2 7 3 13 9 16 0 9 13 2
23 10 11 13 1 10 9 0 1 12 9 2 13 1 12 9 2 16 15 13 1 12 9 2
22 11 13 10 9 3 1 11 11 11 2 11 11 1 3 12 1 15 13 10 0 9 2
15 7 1 10 9 11 12 2 11 8 5 0 2 13 0 2
12 13 10 9 2 11 11 4 13 1 10 9 2
44 1 10 0 9 15 13 10 9 1 10 12 0 9 1 11 1 10 15 13 0 1 10 0 9 2 16 10 9 4 13 15 0 1 9 13 1 10 9 7 9 1 10 9 2
36 4 13 0 1 10 9 0 8 12 2 13 1 12 10 11 11 8 12 7 1 10 9 0 8 12 13 9 1 10 11 8 2 12 1 12 2
28 10 11 2 12 1 11 1 12 2 13 10 9 0 13 3 1 13 10 9 1 10 9 1 0 9 0 0 2
30 1 10 9 2 10 9 13 0 1 9 0 2 10 11 2 2 10 9 15 4 13 1 9 1 11 1 10 9 0 2
13 15 13 1 12 5 1 10 9 9 2 11 11 2
17 10 9 15 13 1 10 9 12 1 10 9 1 10 9 1 9 2
40 10 9 3 4 1 13 15 1 11 2 7 10 12 1 11 1 12 2 3 10 9 3 1 10 0 9 1 10 9 2 15 13 16 10 9 4 13 1 11 2
22 11 13 10 9 1 9 1 10 9 11 16 13 13 1 10 9 1 9 1 9 0 2
36 15 9 13 16 15 13 1 10 9 1 10 11 7 1 10 0 11 7 16 10 9 4 13 15 16 3 15 13 1 13 1 2 10 9 2 2
21 1 10 9 13 11 11 2 10 14 9 1 11 16 13 1 9 1 10 0 9 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
32 15 13 1 10 9 1 3 1 12 9 1 10 9 1 12 9 11 11 11 1 11 2 16 3 15 13 10 9 0 0 0 2
30 15 13 0 1 10 9 1 11 7 15 15 13 1 11 11 16 15 13 10 9 1 9 1 10 15 13 1 12 9 2
6 10 9 13 1 9 2
55 1 13 10 9 10 9 1 10 11 1 10 11 1 10 11 1 10 11 2 9 10 9 1 11 11 11 2 7 1 10 9 1 11 11 2 9 1 10 9 2 13 1 10 9 1 10 9 16 13 10 9 1 10 9 2
40 15 2 13 1 10 0 9 1 9 1 9 13 16 3 13 10 9 1 10 9 1 10 9 2 9 5 9 2 2 15 13 1 10 9 3 0 1 10 9 2
101 10 12 9 13 13 11 2 11 2 10 11 2 11 2 10 11 2 11 2 10 11 2 11 2 10 11 2 11 2 11 1 10 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 10 11 2 10 11 2 11 11 2 10 11 2 11 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 11 2 10 11 2 10 11 2 11 11 7 10 11 2
25 10 9 2 1 10 16 13 10 0 9 1 10 0 9 2 15 13 10 9 1 10 12 1 11 2
33 1 15 2 10 9 1 11 3 3 4 8 4 1 13 1 9 2 1 15 15 3 13 1 9 0 1 10 3 13 3 10 9 2
25 10 9 13 15 1 10 9 1 10 9 1 10 9 2 16 13 1 10 9 10 9 1 0 9 2
20 13 1 10 9 0 15 13 9 2 10 15 13 11 7 10 11 1 11 11 2
21 10 11 1 10 11 15 13 1 11 1 11 2 3 1 10 9 1 11 2 11 2
19 3 2 10 0 9 13 10 9 3 0 7 0 2 1 15 1 10 9 2
34 10 9 13 1 9 1 10 11 1 11 11 2 10 9 0 7 10 9 0 2 13 13 2 1 10 10 9 1 9 0 1 10 11 2
65 13 10 9 1 3 9 0 0 2 12 2 13 15 1 10 9 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 7 12 7 3 13 13 10 0 9 1 10 9 0 1 10 9 12 2
24 10 9 0 15 13 3 1 10 9 1 9 2 15 16 13 10 9 0 13 1 10 9 0 2
40 15 13 3 13 1 10 9 1 10 11 2 1 15 9 1 10 0 9 16 13 1 10 9 1 10 9 1 10 9 1 10 9 2 1 9 1 11 7 11 2
26 15 13 1 11 1 9 0 2 13 7 10 9 15 13 13 9 1 10 9 2 1 9 15 13 3 2
26 13 3 10 12 9 2 13 15 1 15 1 15 1 9 0 2 9 1 10 12 1 11 1 12 2 2
21 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
10 10 9 1 9 15 13 1 10 9 2
27 11 2 11 2 0 1 1 12 5 2 15 13 1 10 9 2 10 9 0 0 2 13 1 10 0 9 2
26 1 9 1 10 9 2 16 13 1 12 2 13 10 9 1 9 0 11 11 2 11 11 7 11 11 2
21 1 13 10 9 2 9 1 11 3 4 13 10 0 9 0 2 10 11 11 11 2
18 13 9 1 11 1 10 9 1 11 2 11 2 11 2 11 7 11 2
54 10 9 1 10 9 2 11 11 11 11 2 4 13 10 11 3 1 10 0 9 0 2 11 11 2 9 3 1 10 9 1 10 9 1 9 0 1 10 16 15 13 10 9 0 1 13 10 9 1 9 1 10 11 2
12 3 0 2 16 13 15 1 9 1 10 9 2
10 10 9 11 4 3 13 1 12 9 2
27 15 2 1 10 3 16 10 10 0 9 1 11 2 4 13 1 11 11 7 11 11 2 9 1 10 9 2
27 10 9 1 9 0 1 10 11 12 2 12 13 1 10 12 2 3 1 3 1 10 10 9 1 10 9 2
26 1 10 9 0 1 11 7 10 11 13 1 12 9 0 2 1 10 15 15 13 10 9 0 1 9 2
19 11 13 10 9 13 1 10 9 1 11 2 11 1 10 9 0 1 11 2
39 10 9 0 2 11 11 2 13 10 9 1 9 0 1 10 9 11 16 15 13 1 11 2 3 7 1 9 7 1 10 9 1 11 2 3 4 4 13 2
17 13 16 15 13 3 0 1 10 9 1 15 10 9 1 10 9 2
19 11 11 11 2 11 2 13 1 11 2 10 11 10 12 1 11 1 12 2
31 1 9 1 9 2 10 9 1 11 4 13 10 9 0 1 10 9 0 2 13 13 2 10 9 1 9 1 9 3 0 2
11 11 2 11 3 4 1 13 1 10 9 2
26 4 13 15 1 10 9 7 9 1 10 9 1 1 10 9 1 9 2 3 1 10 9 1 10 9 2
30 1 10 9 2 10 9 0 13 13 10 9 1 9 1 10 9 2 7 10 9 13 2 1 9 0 2 13 10 9 2
45 11 11 11 13 1 10 9 0 0 10 12 1 11 1 12 1 10 9 11 1 10 9 8 12 8 13 1 10 11 11 1 11 2 11 2 13 9 1 10 9 11 11 1 9 2
52 1 10 9 0 2 10 0 9 1 9 13 10 9 1 9 1 10 9 7 1 9 13 7 13 10 9 1 10 9 7 13 0 13 16 4 13 1 10 9 1 10 9 2 10 4 9 15 13 3 0 9 2
17 1 10 9 15 13 10 9 2 10 9 2 10 9 7 10 9 2
29 10 9 1 9 4 13 1 13 10 9 2 10 9 13 1 10 9 7 11 13 9 1 11 1 10 9 1 9 2
13 1 9 13 9 1 10 0 9 7 10 9 0 2
12 10 9 13 16 11 13 10 9 1 13 15 2
43 10 0 9 8 13 0 1 10 9 0 0 7 4 13 3 1 10 9 0 1 9 1 9 7 9 13 10 9 0 9 1 10 9 7 1 9 1 10 9 1 10 9 2
10 13 16 13 15 9 3 0 1 11 2
17 9 0 7 11 11 2 11 11 1 10 11 11 2 11 11 11 2
24 13 10 9 11 11 1 0 9 2 1 11 11 13 1 12 9 0 2 0 2 0 7 0 2
41 1 10 9 11 1 10 9 1 10 9 0 7 0 1 10 9 11 2 10 9 16 15 13 1 9 3 0 1 10 11 7 10 11 3 15 13 1 9 3 0 2
3 9 11 11
44 10 9 4 13 1 10 9 13 1 10 9 11 1 10 9 1 10 11 1 9 7 9 1 10 9 0 2 16 13 1 12 9 13 1 10 9 1 10 9 1 9 1 9 2
48 10 9 13 1 10 9 0 1 10 3 11 1 11 7 11 11 11 2 11 7 13 1 9 1 10 9 2 10 9 2 10 9 1 10 9 1 10 9 1 11 11 2 7 10 11 11 11 2
25 16 10 9 13 1 10 9 0 3 13 15 16 13 1 10 9 0 7 10 9 0 1 10 9 2
35 1 10 11 11 2 1 12 9 15 13 10 9 2 7 1 15 15 13 1 12 9 2 1 9 0 2 16 13 15 7 13 15 10 9 2
15 13 1 11 11 15 13 1 9 1 10 9 0 1 12 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
44 10 9 0 1 10 0 9 2 10 9 1 11 2 4 13 1 10 9 1 11 11 11 7 1 10 0 9 11 11 1 11 2 15 15 13 1 10 9 1 9 1 10 9 12
28 8 9 0 13 1 10 9 1 11 13 9 1 9 1 10 9 11 7 10 9 1 10 9 1 10 9 0 2
37 1 9 1 15 2 10 9 0 1 10 9 1 11 11 4 13 3 7 13 1 10 0 9 1 9 2 1 9 1 9 2 16 3 13 1 12 2
5 10 9 13 0 2
15 10 9 15 4 13 1 10 9 1 10 9 1 11 11 2
39 10 9 1 9 13 15 1 10 12 9 16 13 10 9 1 10 11 2 13 1 10 9 1 11 2 1 10 9 1 10 9 0 1 11 2 1 10 11 2
11 11 11 13 1 10 11 11 1 10 11 2
20 1 10 15 15 13 10 9 0 13 1 10 9 2 13 1 10 9 7 9 2
53 1 9 1 15 2 15 13 10 0 9 1 9 0 2 7 1 10 9 0 15 13 9 1 10 9 1 9 0 7 9 1 10 9 0 1 9 0 2 13 13 10 11 1 15 3 9 1 15 16 4 13 0 2
10 11 11 13 1 10 9 1 10 9 2
16 15 13 1 13 9 1 10 9 7 3 13 15 13 10 9 2
13 1 0 2 10 9 13 1 8 13 13 3 0 2
19 13 9 0 1 9 2 9 1 10 9 7 9 0 2 1 11 7 11 2
20 1 12 2 11 13 9 0 7 9 1 10 9 1 9 2 11 2 1 11 2
29 3 13 0 10 9 7 9 0 2 16 13 9 1 9 1 10 9 1 9 7 1 9 10 9 0 1 10 9 2
53 10 11 13 10 9 1 10 11 2 11 11 1 10 11 11 2 2 9 1 10 11 11 7 1 10 11 1 10 11 2 11 1 11 11 11 2 2 16 13 1 12 7 12 7 15 4 13 1 10 9 11 11 2
37 3 1 9 1 10 9 12 0 9 1 9 13 1 10 9 1 10 9 16 13 0 7 13 15 1 10 9 7 1 10 9 9 0 1 10 9 2
19 11 2 2 11 2 1 9 2 13 10 9 0 1 9 1 9 11 11 2
27 1 10 12 10 9 0 2 11 11 2 13 1 10 9 1 11 1 10 11 11 11 11 1 10 0 9 2
16 10 9 15 13 1 0 9 0 10 9 10 15 1 10 15 2
28 12 9 1 11 1 11 2 12 1 10 9 1 11 1 11 2 7 10 12 9 3 1 10 9 1 10 12 2
16 3 1 10 12 5 1 10 9 13 1 10 9 1 9 0 2
22 15 13 1 10 9 10 9 13 1 9 0 1 9 0 16 13 10 9 1 11 13 2
25 1 9 2 10 0 9 1 10 9 2 11 2 3 13 10 9 0 1 10 11 11 1 11 11 2
13 10 9 15 13 1 10 9 3 1 10 9 0 2
35 10 9 1 10 11 11 11 13 10 9 1 9 13 1 10 11 1 10 11 1 11 2 7 10 9 3 4 13 16 10 9 13 1 11 2
23 13 9 0 1 10 0 9 11 11 11 2 3 0 7 15 2 7 3 2 7 3 0 2
27 1 10 9 1 10 0 9 2 15 13 1 10 13 10 3 0 2 11 2 2 13 15 7 13 9 0 2
20 10 0 9 13 7 13 10 9 1 9 0 1 8 2 13 1 11 11 11 2
32 15 13 0 1 10 9 0 3 0 2 3 16 15 4 13 9 1 10 9 1 9 16 4 13 10 9 0 1 10 9 0 2
28 10 9 0 1 10 12 9 0 7 10 0 9 0 13 7 13 10 9 1 10 9 1 10 9 0 2 0 2
22 15 1 10 9 15 4 13 1 10 9 1 10 9 7 1 10 9 1 10 9 0 2
21 3 4 1 13 15 1 10 9 7 3 15 13 10 9 16 15 13 10 9 15 2
10 11 13 1 11 7 11 2 11 11 2
20 10 9 13 0 7 10 9 13 0 1 9 0 7 9 16 13 1 10 11 2
38 3 15 13 9 2 1 9 0 1 10 9 2 1 10 9 1 10 9 2 1 15 15 15 13 10 9 0 2 15 15 13 10 9 7 13 10 9 2
66 16 13 3 15 15 4 1 13 1 0 9 15 9 1 10 0 9 1 9 2 10 9 1 9 7 9 16 13 10 9 13 2 10 9 1 10 9 15 2 3 3 2 3 13 7 9 1 9 0 2 7 16 13 1 9 0 10 9 16 10 4 13 1 10 9 2
19 10 9 0 1 10 9 0 13 10 12 1 11 10 9 0 1 10 9 2
19 3 15 13 10 9 1 10 9 1 10 11 15 13 1 9 11 7 11 2
26 15 16 3 4 13 1 10 9 0 13 10 9 1 10 9 16 13 1 11 11 2 1 10 0 9 2
62 9 1 10 11 1 11 11 2 12 2 2 1 10 15 13 1 12 7 12 2 1 10 11 1 11 11 2 12 2 2 1 10 15 13 9 1 12 2 7 1 10 11 1 11 11 1 11 11 2 12 2 2 13 10 9 1 10 11 11 1 11 2
43 11 13 10 9 1 10 0 9 2 11 15 13 3 16 11 15 13 16 13 10 9 1 10 9 9 2 7 15 15 13 7 15 4 13 7 13 13 10 9 1 10 9 2
35 15 7 10 9 0 7 9 4 13 1 10 9 11 1 10 9 1 9 1 10 9 1 10 11 1 11 2 11 2 11 2 11 11 2 2
24 10 11 11 2 11 12 2 2 10 9 1 12 9 2 13 9 1 10 9 0 1 10 9 2
23 1 10 9 12 2 13 1 10 9 11 11 11 16 13 1 11 11 1 10 9 11 11 2
11 1 10 0 9 2 10 9 13 5 12 2
21 1 10 9 0 2 9 9 7 9 9 2 4 13 9 1 11 2 9 1 11 2
34 10 9 11 1 10 0 9 13 0 1 10 9 1 10 9 0 2 1 10 9 16 13 1 10 9 1 9 7 10 9 1 10 9 2
22 13 1 10 9 1 10 9 2 10 9 13 10 9 1 9 7 10 0 9 1 9 2
27 11 13 16 3 13 1 9 2 3 7 15 13 1 9 16 13 1 2 13 1 9 1 10 9 0 2 2
6 4 13 1 12 9 2
29 15 13 1 10 9 3 0 7 0 2 15 4 4 3 13 7 4 13 9 1 10 9 2 10 11 1 11 2 2
23 3 15 13 10 9 9 1 11 2 9 1 11 2 3 15 13 3 10 9 1 12 9 2
32 3 13 10 11 1 11 3 13 10 0 9 0 2 7 1 0 9 13 0 9 1 10 9 11 11 1 12 2 12 2 12 2
38 10 9 0 1 10 9 13 1 12 9 1 15 4 13 1 10 11 11 11 11 2 11 11 1 11 2 2 10 0 9 0 1 10 11 11 1 11 2
10 13 15 1 10 9 3 0 1 11 2
42 16 10 9 11 13 1 10 11 2 15 13 10 9 1 9 13 2 11 2 13 13 10 9 2 15 13 15 13 10 9 1 10 11 7 10 9 1 10 9 11 2 2
8 11 15 13 13 1 10 9 2
23 10 0 9 1 10 9 0 15 13 1 12 7 13 3 3 1 10 9 0 1 10 9 2
21 10 9 13 10 0 9 7 9 11 11 2 0 9 9 1 10 9 8 8 8 2
11 10 9 1 11 15 13 13 1 10 9 2
23 10 12 13 1 10 9 3 0 7 1 15 15 3 0 7 10 12 1 10 9 3 0 2
32 1 11 2 13 10 9 2 3 15 13 1 11 10 9 11 11 16 13 1 11 7 11 11 13 3 13 1 9 1 10 9 2
26 13 10 0 9 16 13 10 9 1 11 11 2 10 9 1 15 2 11 2 13 13 15 1 10 9 2
9 2 10 9 13 10 0 9 2 2
39 9 1 15 2 10 9 1 11 11 15 13 1 9 7 15 13 10 9 2 3 7 11 2 3 1 10 9 1 9 13 10 9 1 10 9 1 10 9 2
33 13 2 3 1 12 2 10 9 0 1 10 9 1 10 11 1 11 2 15 3 3 4 13 1 10 9 1 11 11 1 10 9 2
14 13 10 9 15 13 10 9 1 10 9 2 11 11 2
29 13 1 10 9 1 11 11 1 10 9 1 10 9 9 1 10 9 2 13 15 1 11 7 1 9 2 12 2 2
20 4 13 16 13 10 9 7 3 15 4 13 10 9 1 11 7 10 9 0 2
31 9 3 0 7 9 1 13 10 9 2 10 9 15 15 13 1 10 0 7 15 13 10 9 1 10 9 7 9 1 15 2
27 3 1 10 9 2 13 0 10 9 1 10 9 1 13 15 10 9 1 10 9 1 10 9 1 10 9 2
34 1 10 9 1 10 11 2 11 2 11 7 11 11 2 13 10 9 1 10 9 15 10 11 15 13 3 7 15 13 3 1 10 9 2
14 7 13 16 2 16 4 13 15 2 15 3 15 13 2
11 10 12 13 1 10 9 1 11 7 11 2
9 3 1 10 9 1 10 9 0 2
32 10 9 3 13 10 9 1 9 1 9 2 16 15 15 13 2 13 10 9 1 9 2 3 4 13 10 9 0 1 10 9 2
31 10 9 1 9 0 13 10 9 13 3 10 0 9 1 10 9 1 9 1 0 9 0 7 10 9 1 10 9 0 0 2
37 15 13 15 10 9 1 10 11 11 2 11 2 10 11 2 9 2 1 11 2 11 2 11 11 2 10 0 9 7 9 1 10 9 7 10 9 2
10 13 3 13 1 9 1 9 0 0 2
6 15 13 1 10 11 2
29 13 0 16 15 13 1 13 1 9 1 10 9 11 1 11 8 9 7 9 0 1 11 7 11 13 1 10 9 2
25 1 10 9 1 10 11 13 2 0 1 3 9 2 10 9 11 2 3 13 9 2 9 7 9 2
14 10 9 13 1 12 9 4 13 1 10 9 11 11 2
47 11 11 13 10 9 1 11 1 9 7 9 13 1 11 11 11 11 1 9 1 11 11 11 16 15 13 10 12 1 11 1 12 7 16 13 1 9 1 11 11 2 11 11 7 11 11 2
22 1 9 2 13 10 9 0 7 13 15 1 9 7 9 0 13 1 9 1 9 0 2
13 13 1 9 13 7 13 10 9 0 1 9 0 2
15 9 1 15 1 0 1 13 1 15 10 10 9 16 13 2
12 10 9 1 9 1 10 9 13 1 5 12 2
13 13 12 9 5 1 9 7 12 9 5 1 9 2
62 1 9 2 10 9 0 2 9 7 0 2 3 15 2 1 10 9 13 10 9 1 12 9 1 9 2 9 7 9 2 16 13 16 10 9 15 13 1 13 7 13 10 9 1 10 9 1 10 9 2 1 4 7 13 15 1 13 7 13 10 9 2
27 1 10 9 2 10 9 1 9 15 13 1 10 9 1 9 2 9 2 16 15 4 13 13 9 1 9 2
29 3 1 4 13 2 7 1 9 1 10 9 2 11 15 13 1 11 15 15 3 4 13 9 1 10 9 2 11 2
20 10 9 11 13 10 12 1 11 1 12 1 11 2 11 2 1 10 9 0 2
21 10 10 9 11 11 11 3 4 13 12 5 1 10 9 1 15 1 10 9 0 2
20 11 13 10 9 1 10 8 1 11 2 1 11 2 9 0 1 10 9 0 2
18 1 10 9 0 7 10 9 0 2 10 9 15 13 3 1 10 9 2
35 1 15 2 10 11 13 10 9 0 2 10 9 0 2 10 9 0 7 9 2 10 9 0 0 7 9 1 10 9 7 1 10 9 0 2
26 1 10 9 1 10 9 1 9 13 11 1 0 9 9 1 11 1 10 9 1 9 1 10 9 0 2
40 1 10 9 2 13 1 10 0 9 0 7 13 1 10 12 9 0 13 1 10 0 9 2 1 10 0 9 1 11 2 3 13 10 9 7 13 1 9 0 2
11 11 11 11 13 10 9 1 9 1 12 2
24 1 10 9 13 10 9 1 9 15 4 13 7 13 1 9 1 10 0 9 1 10 9 0 2
60 10 9 13 15 2 10 9 13 1 10 9 1 10 9 0 2 10 9 7 9 1 10 9 1 9 0 16 15 13 1 9 9 0 7 3 2 1 12 2 10 9 1 10 9 1 10 9 11 11 2 16 13 9 1 10 9 0 1 11 2
37 10 11 13 10 9 0 3 0 1 11 2 13 10 9 0 1 12 9 1 9 2 13 1 3 15 13 10 0 9 1 10 9 0 1 10 9 2
39 10 9 13 15 1 10 9 3 0 1 10 9 1 10 9 2 16 13 1 10 9 0 0 13 10 9 1 10 0 1 10 15 13 1 10 9 1 11 2
7 1 11 13 0 9 0 2
16 11 13 0 2 0 1 9 7 3 0 1 9 1 10 9 2
40 10 9 7 9 3 13 13 10 9 1 10 9 7 9 0 1 10 9 1 10 9 1 9 2 10 9 7 10 9 1 10 11 7 10 9 0 1 10 9 2
45 1 10 9 4 13 9 1 10 9 1 11 11 2 11 11 2 11 11 7 11 11 2 11 2 7 3 4 13 10 9 1 4 1 13 1 10 9 1 9 7 1 9 3 0 2
25 11 13 10 0 9 3 0 15 13 10 9 1 10 11 1 3 3 1 10 9 1 11 11 11 2
25 1 9 10 9 15 13 1 10 13 10 11 1 11 12 9 11 11 2 13 1 9 8 11 11 2
41 3 15 13 12 9 1 9 1 10 11 1 10 11 1 11 2 10 9 15 13 1 10 11 1 11 2 13 1 0 9 1 9 1 10 0 9 1 10 9 12 2
26 3 13 15 16 13 1 1 1 10 9 7 3 1 10 9 1 10 9 7 1 10 9 1 10 9 2
27 11 13 10 0 9 1 10 9 1 10 9 7 10 9 2 10 9 13 9 0 1 10 9 1 10 9 2
24 15 15 13 1 9 0 2 3 15 13 1 10 9 1 11 0 1 15 15 13 10 11 11 2
12 10 9 1 11 11 15 13 13 1 10 9 2
4 13 1 11 2
13 10 9 13 10 9 1 10 9 1 0 9 0 2
16 3 3 2 10 9 2 9 2 4 4 13 1 10 0 9 2
17 10 12 1 11 1 12 15 13 10 9 1 10 9 12 7 12 2
33 11 13 1 10 9 1 10 9 0 12 2 9 12 1 10 9 2 9 12 1 10 9 2 7 1 10 9 1 10 9 11 11 2
24 11 11 4 13 1 10 9 1 10 11 11 7 3 13 3 0 1 16 13 1 9 1 9 2
20 15 1 10 9 7 9 1 11 11 2 11 13 9 1 10 9 0 7 0 2
18 1 10 9 12 10 9 11 13 10 9 2 11 11 11 11 11 2 2
25 10 9 13 10 0 9 0 16 13 10 9 0 2 13 1 10 9 1 10 9 0 2 7 13 2
33 10 11 13 10 9 15 13 10 9 1 9 13 1 10 9 0 1 10 0 9 2 9 1 11 11 2 9 1 11 11 2 11 2
22 13 10 12 1 12 9 1 9 1 10 9 2 7 16 10 9 13 3 1 12 9 2
42 1 12 11 13 10 0 9 1 13 10 9 1 0 9 1 11 11 2 3 15 13 1 13 10 9 1 11 2 10 9 16 13 10 9 0 1 10 13 1 11 11 2
19 1 13 10 9 1 10 9 0 2 11 13 10 9 0 0 1 10 9 2
33 15 13 1 9 16 13 15 10 9 1 9 1 10 9 0 16 13 0 7 15 13 9 1 13 10 15 1 10 9 1 10 9 2
17 10 11 11 11 13 10 9 1 9 1 11 1 10 9 1 11 2
32 1 12 2 11 11 13 1 10 9 1 9 10 9 1 9 1 10 9 1 11 11 11 2 13 1 10 9 1 10 8 0 2
23 1 12 13 3 1 11 11 1 10 9 11 11 11 11 2 13 1 11 2 13 9 0 2
21 10 9 15 13 3 1 9 7 0 1 10 15 13 10 9 0 13 7 10 9 2
41 7 10 9 13 3 10 9 0 1 10 9 1 15 3 13 3 3 0 2 7 16 13 9 2 3 10 9 13 0 7 3 7 3 9 2 7 9 1 10 9 2
23 13 10 9 0 16 13 10 9 1 12 9 1 9 2 0 2 13 1 9 1 12 9 2
25 10 9 0 1 10 15 4 13 15 10 9 13 9 2 9 2 9 7 9 2 9 7 9 2 2
24 10 9 1 11 11 11 13 15 1 13 9 3 3 1 10 9 1 9 1 3 1 10 9 2
20 13 1 11 2 4 13 1 15 1 10 9 1 10 9 0 1 9 1 11 2
18 11 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
81 1 10 9 2 10 9 1 10 11 11 11 4 13 16 10 9 3 4 13 0 1 13 10 10 9 0 1 10 9 11 11 2 2 15 15 4 13 1 10 9 1 9 2 11 11 2 1 10 4 15 13 1 10 9 1 12 9 10 9 13 1 10 11 7 10 9 1 9 2 1 9 1 10 9 1 10 9 0 1 11 2
20 10 9 1 10 9 3 13 0 2 7 10 9 1 11 3 1 15 13 0 2
27 1 10 9 2 10 9 1 9 0 1 11 15 13 1 3 1 12 9 1 10 16 13 3 1 10 9 2
24 1 10 9 12 2 10 9 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
20 4 13 1 13 1 10 0 9 3 1 11 2 16 13 1 9 1 10 9 12
87 13 10 9 1 9 2 15 1 9 7 1 9 2 16 3 15 13 1 12 9 1 10 9 0 7 16 13 1 9 12 9 1 9 0 2 1 9 1 9 3 15 4 13 15 2 1 9 0 1 10 9 0 1 10 9 7 13 1 10 9 0 3 2 10 9 13 0 7 15 15 13 10 9 1 10 9 1 10 15 15 13 2 3 1 10 9 2
28 10 9 3 0 3 13 10 11 2 11 11 2 2 13 1 12 2 9 16 11 3 13 15 1 10 0 9 2
17 10 9 1 10 9 4 13 1 10 9 1 11 15 11 1 12 2
16 10 9 13 1 10 9 1 11 11 2 0 9 11 1 11 2
23 11 13 10 0 9 1 10 9 7 1 11 15 13 1 10 9 1 10 9 1 11 11 2
13 1 9 15 13 10 9 1 10 9 1 9 0 2
29 15 1 10 0 9 13 10 9 0 7 10 0 7 0 9 1 9 0 1 10 13 15 1 9 0 1 9 0 2
22 1 10 9 1 11 2 4 13 1 0 9 2 13 11 11 2 11 11 7 11 11 2
38 1 0 9 1 10 9 16 13 10 11 11 11 11 11 2 15 13 0 9 16 13 1 10 9 2 13 1 0 7 0 9 7 10 0 7 0 9 2
32 9 1 10 11 1 11 2 10 11 1 11 0 2 10 11 11 0 2 4 1 4 13 1 9 1 10 9 1 9 0 0 2
12 11 11 13 10 9 1 9 1 10 9 11 2
35 1 10 0 9 1 10 9 2 11 13 1 10 9 0 3 13 10 9 1 9 9 13 1 10 9 1 10 9 0 11 11 7 11 11 2
55 1 9 1 10 9 2 10 9 0 13 10 9 1 10 9 1 10 9 0 2 10 15 13 1 10 9 1 12 12 12 9 2 1 10 9 1 10 11 2 9 16 15 13 1 12 12 12 9 1 10 10 9 1 9 2
17 10 9 15 13 1 10 0 9 2 13 9 10 9 0 1 11 2
23 10 9 1 9 16 13 1 10 9 1 9 1 11 13 8 11 11 11 1 11 11 11 2
5 10 9 3 0 2
17 13 1 11 1 12 2 13 3 9 3 1 16 10 9 4 13 2
18 10 9 15 13 1 10 9 7 3 13 2 13 10 9 1 10 9 2
25 11 13 1 11 11 2 11 2 11 1 11 2 11 1 11 2 11 11 2 11 11 7 11 11 2
9 4 13 3 1 9 1 10 9 2
12 1 10 3 11 11 4 13 1 9 1 11 2
14 16 15 13 1 9 0 2 10 9 13 13 12 9 2
35 1 10 9 0 1 3 1 12 12 9 1 9 0 1 11 2 10 11 13 9 1 9 1 9 16 13 9 0 2 0 7 0 1 9 2
30 15 1 10 0 9 1 10 15 4 13 15 10 9 1 10 9 0 13 1 10 9 1 10 9 0 7 10 9 0 2
14 10 9 13 2 10 9 15 13 1 0 9 1 9 2
26 10 9 1 9 15 13 10 12 1 11 1 12 1 10 9 1 10 9 11 7 10 9 1 11 11 2
28 1 9 2 1 0 9 2 4 13 2 3 1 3 4 13 1 10 0 9 16 13 3 10 9 1 10 9 2
11 12 11 13 10 9 1 11 7 10 9 2
10 15 13 1 11 2 11 1 10 11 2
12 1 10 9 10 9 13 9 1 10 9 11 2
24 1 10 9 2 11 15 13 1 13 10 9 1 12 9 0 1 9 16 13 1 12 1 9 2
20 1 0 9 2 10 9 1 10 9 3 4 13 1 10 9 1 10 0 9 2
27 10 9 1 10 9 13 1 10 9 7 10 9 1 10 9 13 7 3 10 9 1 9 16 15 4 13 2
19 1 9 1 10 9 12 2 11 13 10 9 1 9 0 0 7 11 11 2
38 7 3 11 11 13 16 13 10 9 0 1 11 2 10 9 0 2 11 3 15 13 2 7 13 0 15 3 15 13 1 10 9 13 1 10 9 0 2
29 10 9 1 9 13 1 10 9 1 11 2 1 10 9 2 10 11 11 2 2 1 10 9 1 10 9 1 11 2
26 11 4 13 2 3 3 3 1 9 2 1 10 12 9 1 9 2 9 1 15 10 9 15 13 13 2
70 8 2 2 10 9 13 1 16 10 9 13 10 0 9 7 1 15 3 13 10 11 2 2 13 2 10 9 1 9 1 10 9 1 11 2 8 11 11 2 13 10 9 13 1 10 9 1 9 1 10 9 2 11 11 2 1 10 9 1 10 0 9 1 11 11 1 11 1 9 2
31 1 10 9 11 13 3 1 13 10 0 9 1 10 9 0 7 0 1 15 13 10 9 0 1 11 11 1 11 1 12 2
27 11 15 13 1 13 10 9 1 9 1 13 7 16 13 10 9 16 15 13 0 1 10 9 0 1 9 2
14 1 12 13 10 9 0 1 10 0 9 0 0 0 2
24 3 2 10 11 13 13 3 10 9 1 11 11 2 10 9 16 13 1 9 0 7 1 9 2
14 13 1 10 9 0 13 15 1 10 9 16 13 13 2
59 10 9 15 13 0 2 16 1 10 9 15 13 1 15 2 10 9 16 13 10 9 2 1 10 9 2 3 13 16 10 9 13 1 10 9 16 13 16 1 10 9 3 15 13 2 7 11 11 4 1 13 1 12 7 12 9 10 9 2
28 15 13 3 1 10 9 0 10 0 9 2 10 11 11 2 16 15 13 13 10 9 10 12 9 1 10 9 2
52 1 10 9 4 13 1 10 9 11 11 11 1 13 15 1 10 9 1 11 11 2 3 13 1 9 1 12 3 10 9 11 11 11 15 13 1 10 9 2 16 3 13 12 9 2 3 16 11 13 10 9 2
34 11 2 11 11 11 11 13 10 11 1 11 11 1 12 7 13 10 9 1 13 9 1 11 2 15 3 4 4 13 1 11 11 2 2
31 1 12 9 1 9 0 1 3 9 2 10 9 4 4 4 3 13 1 9 0 2 3 1 10 9 0 1 10 1 12 2
6 3 1 9 7 9 2
18 10 9 15 13 1 15 3 9 2 13 1 10 10 9 1 10 9 2
12 4 13 3 2 12 5 2 1 10 9 0 2
17 3 1 16 10 9 4 13 10 9 13 1 12 9 1 10 9 2
22 4 13 1 10 9 1 10 0 7 0 9 1 10 9 1 9 1 10 11 11 11 2
20 4 13 3 1 10 9 1 9 7 13 3 13 10 9 1 9 1 10 9 2
19 1 13 2 15 13 1 10 9 1 10 9 11 7 9 1 10 9 13 2
28 10 9 13 0 7 13 9 2 10 9 1 10 9 13 10 9 1 10 9 3 7 1 10 9 7 9 0 2
30 1 10 9 2 11 13 1 10 11 11 1 11 7 11 11 2 0 1 11 11 2 8 9 1 10 11 11 1 11 2
35 4 1 13 10 9 1 10 11 8 7 13 10 9 16 3 13 9 1 10 9 7 15 13 0 7 0 9 1 10 9 7 1 10 9 2
49 11 11 2 8 12 1 11 1 12 2 13 10 9 1 9 0 2 9 7 9 1 9 2 3 13 1 4 13 10 9 1 11 11 12 7 3 3 1 13 10 9 1 10 9 1 9 0 11 2
35 13 10 9 16 13 1 10 9 1 10 11 2 13 10 11 1 10 9 1 10 16 15 13 1 10 9 16 4 13 2 7 10 9 13 2
27 1 10 0 9 1 10 9 2 1 12 2 11 13 13 10 9 1 9 2 1 15 16 13 9 7 9 2
38 10 12 9 13 1 9 13 10 9 1 10 9 2 1 10 9 7 1 10 9 0 2 13 1 10 9 0 16 13 10 10 9 0 1 10 0 11 2
7 10 9 0 13 12 11 2
27 11 11 4 13 1 10 9 8 2 12 0 2 1 10 13 12 9 1 10 15 13 10 0 9 1 9 2
11 4 13 1 10 9 1 10 9 1 9 2
29 7 1 15 13 12 9 2 10 0 15 0 1 9 2 9 2 8 7 10 0 15 0 1 10 9 1 10 9 2
58 3 2 10 9 0 13 1 10 9 1 11 11 2 9 1 10 9 1 11 11 11 2 3 13 1 9 10 9 1 9 1 10 9 1 11 2 7 10 9 1 10 9 0 1 10 9 1 9 7 1 9 1 10 9 1 10 9 2
36 11 11 11 1 11 7 11 2 12 1 11 1 12 2 2 12 9 1 11 2 12 9 1 11 2 12 9 1 11 11 7 12 9 1 11 2
28 1 11 2 11 2 11 7 11 13 10 9 12 2 12 7 12 2 3 2 1 10 9 1 10 9 10 11 2
36 10 9 1 11 3 13 10 0 9 15 4 13 1 10 9 1 11 9 3 7 4 13 1 15 7 1 10 9 1 13 1 10 9 3 13 2
17 1 9 2 15 4 13 10 9 1 9 7 9 1 3 12 9 2
37 1 10 9 0 1 10 9 2 3 13 9 1 10 9 1 11 2 1 15 15 4 13 1 9 0 9 1 10 9 0 1 10 9 1 10 11 2
25 1 10 9 1 12 2 11 11 13 10 9 7 13 10 0 9 1 10 9 0 1 10 9 0 2
24 10 9 13 13 9 12 1 9 0 2 13 9 0 1 9 0 2 9 0 2 7 9 0 2
38 10 9 13 1 11 11 13 1 10 9 10 9 0 1 9 1 2 11 11 7 11 2 16 2 8 9 1 13 0 9 2 15 13 12 9 1 11 2
70 10 9 1 9 1 11 4 4 13 1 10 9 0 9 1 9 1 12 7 13 10 0 9 1 10 9 1 11 1 10 9 1 11 2 13 1 10 9 1 10 11 7 11 2 1 10 9 1 11 7 11 2 16 13 1 10 9 0 1 11 7 11 16 15 13 1 15 1 11 2
24 10 0 9 2 9 3 0 7 0 9 2 13 1 10 11 11 10 9 0 1 13 10 9 2
20 15 4 13 10 12 9 16 13 10 9 1 10 9 7 13 15 10 0 9 2
27 1 10 0 9 15 13 10 9 1 10 9 2 1 10 9 0 1 11 7 11 11 11 2 9 1 11 2
11 9 0 1 10 9 1 10 9 1 11 2
28 15 13 16 10 9 1 10 9 15 13 10 9 1 10 9 2 7 3 3 4 13 1 10 9 1 9 2 2
32 10 9 0 3 3 13 10 9 13 15 1 10 9 1 1 10 9 3 2 7 16 3 13 9 1 9 7 9 1 0 9 2
32 10 11 11 13 10 9 1 9 1 10 9 11 2 13 1 11 1 9 11 1 11 1 12 7 1 11 1 9 1 9 11 2
15 13 1 10 9 0 2 9 7 1 10 9 1 10 11 2
22 10 9 1 10 9 11 13 1 9 0 2 13 0 9 1 11 11 7 10 9 0 2
39 3 13 9 1 9 7 9 2 3 4 7 13 2 13 2 13 10 9 1 0 9 2 9 2 9 2 7 0 9 16 13 1 9 3 0 2 3 0 2
27 10 0 9 4 13 9 1 9 0 2 9 16 13 1 13 1 9 1 10 11 11 1 11 11 1 12 2
19 13 10 9 13 10 9 1 10 9 2 13 10 9 1 10 0 9 0 2
31 10 0 9 15 13 1 9 1 9 2 0 9 1 9 2 9 1 9 0 2 7 1 10 9 0 2 3 0 2 11 2
41 10 9 2 13 10 9 1 9 0 2 0 2 0 2 0 2 0 7 0 2 13 1 10 9 0 1 9 0 3 13 1 9 1 10 9 1 12 9 1 9 2
16 1 10 0 13 12 9 1 9 1 10 9 1 11 2 11 2
17 1 10 9 15 13 9 2 9 2 9 7 9 1 10 9 0 2
41 11 4 1 13 1 10 9 2 3 10 9 13 0 2 7 1 10 9 2 13 10 9 1 9 16 13 10 9 1 13 10 9 1 9 16 3 4 13 1 9 2
8 3 13 1 10 9 1 11 2
38 1 10 9 1 9 2 13 1 9 2 9 1 9 2 2 15 13 10 0 9 1 10 9 7 9 16 13 13 1 10 0 9 16 13 10 3 9 2
35 10 9 1 9 1 9 13 1 10 9 1 13 10 9 2 7 10 9 16 15 13 13 10 9 12 9 2 1 10 12 1 10 9 12 2
50 13 3 15 16 10 9 0 15 13 1 9 7 3 13 9 16 13 10 9 1 10 9 1 10 2 9 2 16 15 13 1 9 7 2 13 10 9 2 16 13 1 10 9 10 9 0 1 10 9 2
48 10 9 7 10 9 2 8 5 8 1 9 2 13 10 9 0 1 12 1 9 0 7 0 0 7 0 1 11 11 2 7 0 1 11 11 11 2 11 11 11 2 11 11 7 11 11 15 2
22 11 11 11 2 13 8 8 10 9 1 9 9 0 1 12 2 13 1 11 11 11 2
37 7 2 1 10 8 2 9 1 13 10 9 1 9 12 2 13 10 9 0 1 10 9 0 0 2 15 16 15 13 3 1 10 9 1 12 9 2
9 13 10 9 7 13 10 0 9 2
32 1 13 1 10 9 11 13 13 15 3 1 10 12 5 1 9 1 10 9 0 1 10 9 2 15 9 15 15 13 1 13 2
5 1 9 13 0 2
25 15 15 13 10 9 0 1 10 9 1 15 7 9 1 11 13 10 9 3 7 4 13 10 9 2
47 10 9 13 10 9 1 12 9 5 2 10 15 12 9 5 4 13 1 9 2 2 10 9 1 12 9 2 7 10 9 1 9 13 1 12 8 2 9 5 2 1 9 0 1 12 2 2
27 10 9 1 10 9 13 1 9 0 1 9 3 0 2 16 13 10 9 1 10 9 7 10 9 1 9 2
9 15 13 0 1 9 1 10 11 2
19 2 13 3 1 9 16 13 9 0 1 15 16 15 4 13 2 2 13 2
34 15 13 10 0 9 1 11 7 1 10 9 2 4 13 1 13 10 0 9 1 11 11 11 2 13 15 1 10 0 9 1 10 9 2
35 13 0 1 16 4 13 1 10 9 1 10 9 7 16 1 9 1 16 15 13 1 10 9 15 3 1 15 16 13 2 15 4 13 0 2
60 1 10 12 9 2 11 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 9 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
48 7 10 9 1 11 3 4 13 10 9 0 2 8 9 1 10 9 2 13 13 15 16 13 15 1 10 9 2 15 7 13 13 15 1 10 10 9 1 11 7 4 1 13 15 15 1 9 2
12 1 12 13 9 1 10 9 11 1 9 0 2
11 1 10 9 2 15 3 3 13 10 9 2
28 13 10 9 1 9 0 13 1 10 9 2 3 1 10 9 1 9 2 9 0 2 9 1 9 7 9 0 2
16 15 13 1 10 9 16 3 4 13 3 10 9 1 10 9 2
30 10 9 13 0 1 9 1 9 2 10 9 13 15 16 13 2 3 1 13 9 2 4 13 15 1 10 15 1 9 2
19 10 9 13 13 15 13 1 9 7 3 15 13 10 9 1 13 10 9 2
12 16 15 13 13 9 1 10 9 15 15 13 2
16 15 13 1 10 0 9 1 9 13 1 9 1 10 11 11 2
32 3 0 2 7 2 13 2 10 9 3 13 9 1 13 15 10 9 1 10 9 1 10 9 2 10 13 0 7 10 9 0 2
13 0 9 4 13 7 13 1 9 1 10 9 0 2
51 1 15 9 1 10 9 1 12 7 12 2 11 13 10 9 0 1 9 0 2 7 15 15 13 16 13 9 1 10 9 1 10 9 0 2 10 9 0 1 10 9 0 7 10 9 0 13 1 10 11 2
22 11 11 2 4 13 10 9 1 10 9 1 10 10 9 2 1 10 9 1 10 9 2
11 13 1 0 9 10 9 7 9 0 0 2
22 13 16 10 9 15 13 1 11 7 1 10 9 15 4 13 1 15 16 13 1 9 2
3 9 0 2
60 1 10 12 9 2 11 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 9 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
21 1 9 2 10 12 1 11 1 12 13 10 0 9 16 15 13 1 3 0 9 2
9 1 10 9 15 13 10 9 0 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
19 15 13 1 11 11 2 10 9 16 4 1 13 10 9 1 9 1 9 2
14 13 10 0 9 1 10 9 7 3 13 3 0 9 2
47 4 4 13 1 10 9 11 12 11 11 1 11 11 1 10 9 1 9 11 2 11 2 7 9 2 9 12 5 11 1 11 11 11 11 11 1 10 11 11 1 9 1 11 2 1 15 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
85 13 1 10 9 1 10 9 1 11 2 11 2 7 11 2 11 2 2 1 10 9 1 11 2 11 2 7 11 2 11 2 11 2 2 1 10 9 1 11 2 11 2 2 1 10 9 1 11 2 11 2 2 1 10 9 1 11 2 11 2 1 10 9 1 11 2 1 2 11 2 7 1 10 9 1 11 2 11 11 7 11 2 11 2 2
12 13 0 13 10 9 0 1 4 13 10 9 2
60 1 10 12 9 2 11 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
36 10 9 16 13 9 0 3 15 4 13 1 9 0 2 7 16 10 9 0 16 13 13 10 0 9 3 13 10 9 2 16 3 4 13 9 2
20 2 10 11 2 13 10 0 9 0 7 10 9 10 9 1 10 11 11 2 2
23 10 9 13 10 9 16 4 13 1 10 9 0 0 7 0 2 1 10 9 0 7 0 2
35 10 9 13 1 10 9 0 1 15 1 10 9 0 3 1 10 9 0 2 1 15 15 15 13 16 3 13 10 9 0 1 10 11 11 2
18 10 9 1 10 9 7 1 10 9 13 0 1 10 9 1 10 9 2
18 10 9 3 13 8 7 16 13 9 15 13 3 3 2 0 1 9 2
13 3 15 13 1 10 9 1 9 7 10 10 9 2
27 1 10 9 0 1 10 9 1 9 2 10 12 5 13 0 1 12 7 10 12 5 13 0 1 12 9 2
25 15 13 10 9 0 1 10 9 1 10 9 13 1 9 1 11 1 10 9 1 11 11 1 11 2
33 1 12 13 10 9 2 4 1 13 1 9 1 10 9 0 1 11 2 11 7 11 2 7 1 13 1 10 9 1 10 9 0 2
24 3 13 1 11 1 10 9 1 11 11 11 2 1 10 9 2 11 11 11 2 2 12 2 2
18 13 1 10 0 9 10 12 1 11 1 12 13 1 10 11 1 8 2
24 10 9 13 13 2 1 10 9 0 7 0 2 1 12 9 0 0 2 1 9 9 2 9 2
16 13 10 0 9 16 13 1 10 9 1 9 7 1 10 9 2
44 1 10 11 12 3 1 9 13 1 10 9 0 1 10 11 2 2 3 11 13 10 11 12 1 11 11 13 10 9 0 7 13 1 10 9 3 1 16 10 9 13 3 0 2
13 11 11 13 15 1 10 9 16 10 9 13 13 2
54 10 9 4 4 13 1 9 1 10 9 1 9 1 10 9 2 13 1 9 1 10 0 11 1 10 11 2 10 8 9 1 10 11 11 11 11 2 7 10 0 13 1 9 11 11 2 1 10 9 1 11 11 2 2
12 10 9 7 9 0 13 10 9 0 7 0 2
39 3 2 10 12 1 11 11 13 1 11 2 11 11 7 11 11 1 10 11 1 10 9 1 16 3 13 9 1 9 1 10 9 7 11 4 13 10 9 2
19 10 9 4 13 1 12 1 10 11 1 12 9 7 13 0 1 12 9 2
12 13 3 1 11 11 2 3 13 10 0 9 2
29 1 12 2 10 12 0 9 0 1 10 9 1 9 2 13 16 13 9 1 10 9 1 9 1 10 9 4 13 2
60 1 12 13 1 10 9 11 11 8 8 8 1 10 0 9 0 10 9 13 3 12 9 1 10 15 10 9 12 13 1 10 9 1 13 1 10 11 11 7 11 11 11 1 11 2 1 3 1 10 12 13 1 10 9 11 11 11 1 11 2
5 13 1 11 11 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
36 7 3 15 13 1 9 1 16 13 1 10 0 9 0 1 11 2 3 13 9 1 10 9 1 7 15 13 7 10 9 0 16 13 10 9 2
19 1 9 3 13 10 9 1 10 16 13 1 15 15 15 13 1 13 15 2
83 10 9 2 13 1 10 9 0 1 10 9 0 1 10 9 1 10 11 2 3 12 2 2 10 9 1 9 1 11 7 1 10 9 1 11 2 2 8 2 2 3 7 10 9 1 9 1 10 9 1 9 16 4 13 1 10 9 11 2 8 2 2 13 1 9 10 9 1 9 0 9 1 10 11 2 16 15 13 1 12 7 12 2
10 10 9 7 9 1 10 9 13 0 2
11 1 12 2 11 4 13 9 0 1 11 2
26 11 2 11 2 11 13 10 9 1 9 1 10 2 11 11 11 11 11 2 1 10 9 0 1 11 2
21 4 3 13 2 9 12 2 13 15 15 10 9 1 10 9 7 10 9 0 9 2
33 10 9 15 13 1 9 1 10 9 1 13 1 10 9 1 9 1 10 9 1 10 9 2 10 9 13 16 10 9 13 3 0 2
29 15 13 13 1 10 9 1 9 0 1 11 8 8 11 11 8 8 11 2 10 9 0 1 11 11 7 11 11 2
32 10 9 4 13 1 9 2 12 9 2 12 9 2 12 9 2 10 11 1 8 2 12 9 2 12 9 2 12 9 7 9 2
58 10 9 1 9 16 13 10 9 0 13 13 10 0 9 1 9 1 9 1 10 9 2 16 1 10 9 15 13 1 9 1 9 1 9 2 1 15 1 10 16 10 9 13 10 16 13 10 9 0 1 16 10 9 4 13 10 9 2
28 10 9 4 13 1 12 9 2 0 2 1 9 0 2 9 7 9 2 2 7 0 2 9 0 2 9 2 2
13 7 11 1 11 11 13 1 10 9 1 10 9 2
22 3 13 1 11 11 15 1 10 12 0 9 1 10 9 7 1 10 0 1 9 0 2
4 13 1 11 2
6 13 1 15 4 13 15
21 15 13 13 15 9 7 9 0 7 13 0 1 13 10 9 1 9 1 10 9 2
18 11 13 1 11 1 10 12 9 1 10 9 1 13 9 1 10 9 2
12 10 9 2 3 7 1 10 9 1 10 9 2
2 13 12
13 2 9 2 9 10 11 2 12 1 11 1 12 2
27 1 12 10 9 13 10 9 11 7 13 1 11 2 3 13 10 9 7 1 9 13 10 9 1 9 0 2
20 11 11 13 10 9 1 10 9 1 9 1 11 7 10 9 1 9 1 11 2
21 1 10 9 0 13 0 16 10 9 4 13 0 1 10 9 7 10 3 0 9 2
41 1 10 9 0 13 0 13 2 1 9 0 2 1 9 7 0 2 9 7 9 0 2 8 1 9 2 3 13 2 1 10 9 3 0 2 0 9 7 0 9 2
57 9 7 3 11 2 1 9 2 8 2 1 9 0 2 9 2 1 9 2 9 2 13 10 9 1 11 2 13 1 10 9 3 1 10 9 1 11 7 1 11 2 1 3 12 9 1 10 9 1 11 7 1 12 9 1 11 2
18 1 10 9 1 12 2 1 12 9 2 4 13 10 9 1 9 0 2
58 10 9 15 13 7 13 10 9 1 9 0 2 0 7 0 2 16 16 15 4 13 10 9 0 2 16 16 15 13 12 9 7 15 15 2 7 9 7 13 13 2 0 13 10 9 0 2 2 7 3 13 1 13 15 1 10 9 2
56 1 10 9 12 7 1 10 0 9 1 10 9 1 10 11 2 10 11 11 11 1 9 1 10 9 11 1 15 2 13 1 0 9 3 1 12 9 0 2 10 9 0 3 1 10 9 1 11 2 0 9 0 1 10 9 2
75 1 9 1 10 9 2 15 13 10 9 1 10 11 11 1 11 11 2 1 9 7 1 10 9 1 12 9 2 1 10 9 11 1 10 11 1 11 2 10 12 1 11 1 12 2 1 10 15 15 13 10 9 0 7 0 1 11 11 1 10 9 2 15 13 10 9 13 7 15 13 1 13 10 9 2
16 1 3 13 0 1 9 2 15 13 3 1 9 0 1 9 2
44 3 15 13 16 10 9 3 0 2 1 9 0 2 3 13 9 0 0 1 10 15 1 15 1 9 2 7 16 13 10 9 1 2 13 9 1 9 2 2 16 13 10 9 2
20 1 10 9 1 10 11 15 13 9 1 2 2 9 1 9 1 0 9 2 2
48 3 0 2 16 3 13 10 9 10 9 0 9 1 10 9 1 11 2 13 1 9 3 2 0 2 1 13 0 2 13 10 9 16 1 10 9 13 1 10 9 0 15 13 16 13 1 13 2
16 3 10 9 13 10 9 1 13 15 7 13 15 1 10 9 2
29 13 9 1 9 0 1 11 7 11 11 2 15 1 10 9 1 11 2 7 13 10 9 1 9 7 1 9 11 2
38 3 2 10 9 1 0 9 7 10 9 1 13 9 13 10 9 0 2 13 10 9 1 11 2 15 15 2 3 2 1 9 0 13 1 9 1 9 2
22 2 2 2 15 3 13 10 9 0 2 4 4 13 1 10 9 0 13 1 9 2 2
43 10 0 9 13 16 11 11 2 9 1 11 2 1 10 13 13 1 11 7 10 9 15 13 1 11 11 1 12 1 10 9 0 1 11 1 10 9 1 10 9 11 11 2
40 13 10 9 2 16 3 13 10 9 1 9 7 1 9 2 2 1 4 4 13 1 10 9 1 10 9 13 1 10 9 0 0 1 10 12 1 11 1 12 2
33 3 13 1 10 11 1 12 2 7 3 13 1 10 9 7 9 0 16 4 13 9 2 1 10 9 1 10 11 11 2 11 11 2
21 4 1 13 10 12 9 16 13 2 16 13 16 13 10 9 1 9 2 2 13 2
11 1 15 13 10 9 11 1 13 1 11 2
40 1 10 9 13 1 10 9 0 1 11 1 10 9 2 10 9 1 11 2 9 1 11 2 13 16 3 13 2 10 10 9 13 1 10 9 0 1 9 2 2
16 1 10 9 13 10 9 1 10 9 1 9 0 7 9 0 2
46 10 0 9 13 10 11 16 13 0 7 16 13 13 1 10 11 11 16 13 10 9 16 13 1 11 11 2 10 9 1 12 9 16 13 1 9 7 1 9 13 10 9 0 1 11 2
27 10 12 11 11 1 11 11 1 11 15 13 1 11 2 11 2 1 10 12 1 10 12 1 11 1 12 2
33 10 9 15 13 1 10 9 0 1 9 0 2 13 10 9 1 10 9 16 15 13 3 2 9 2 9 2 9 2 7 15 2 2
42 10 11 11 11 11 13 10 9 0 13 1 10 9 1 10 9 11 1 12 9 1 11 11 2 1 10 9 1 11 2 2 11 2 7 11 2 11 2 2 10 11 2
23 1 12 13 1 11 7 10 9 1 10 9 12 0 13 1 10 0 9 1 13 10 9 2
5 15 13 1 11 2
11 4 13 1 9 0 1 10 9 7 9 2
16 2 9 13 10 9 1 11 11 2 2 13 10 11 1 11 2
52 10 9 7 9 13 3 10 9 1 9 1 10 9 1 9 1 9 1 9 13 3 1 10 9 1 10 9 2 10 9 1 10 9 1 10 9 1 10 9 7 10 9 1 10 9 1 9 15 13 9 11 2
9 10 9 4 4 13 1 9 0 2
17 10 9 3 15 13 1 13 10 9 0 7 1 13 10 0 9 2
26 15 13 9 1 10 9 15 11 13 1 10 9 11 11 2 15 1 10 9 13 1 10 3 0 9 2
31 10 9 0 2 0 1 10 9 2 13 10 9 1 10 9 1 15 2 10 12 9 1 0 1 10 12 9 1 9 2 2
20 10 12 1 11 2 10 9 13 10 9 1 10 11 2 13 1 10 9 9 2
52 10 9 4 13 10 12 1 11 1 12 7 10 9 13 1 11 11 13 1 12 9 1 11 11 2 11 11 2 13 11 1 10 11 2 11 1 11 2 7 11 11 11 11 2 10 11 9 11 1 11 2 2
12 13 3 0 10 9 13 11 13 1 11 11 2
32 13 1 10 0 9 1 10 9 2 4 13 15 1 10 9 1 12 9 0 2 10 9 0 2 10 9 0 7 10 9 0 2
41 1 9 1 16 10 9 13 0 7 3 13 9 1 9 3 15 15 4 13 1 10 0 9 1 10 9 8 10 0 9 2 3 15 13 1 10 9 1 10 9 2
16 11 11 11 11 13 10 9 1 9 1 9 1 11 2 11 2
39 1 12 9 13 1 10 9 7 13 10 0 9 2 15 16 15 13 1 13 2 3 1 11 2 1 3 13 10 9 1 9 16 15 13 1 10 10 9 2
7 11 13 3 7 15 13 2
48 3 1 10 9 1 9 2 10 9 0 1 9 4 4 13 1 13 0 9 1 9 2 0 1 9 1 0 9 7 9 1 9 2 9 2 1 10 9 1 10 9 1 9 0 1 9 0 2
19 13 10 11 11 11 1 11 1 12 2 7 4 1 13 10 9 0 0 2
27 3 11 2 11 2 11 7 11 13 10 0 9 2 13 1 10 9 10 11 11 1 11 11 7 10 11 2
22 10 9 13 16 3 3 15 13 7 15 13 1 11 16 15 13 1 10 9 7 13 2
57 11 13 13 10 9 1 10 11 0 3 13 0 9 2 15 3 1 15 16 4 13 1 9 1 3 2 3 7 4 4 13 3 10 9 4 13 1 3 1 3 1 10 9 1 9 1 16 4 13 1 10 0 9 13 10 9 2
13 10 9 1 12 9 13 1 12 1 12 9 3 2
40 10 9 13 2 1 10 9 2 9 1 10 9 7 9 1 9 2 10 9 2 0 2 2 10 9 1 9 1 10 15 15 13 13 10 9 1 10 9 0 2
17 13 1 10 9 1 10 9 2 10 9 0 13 16 13 9 0 2
43 1 9 0 2 10 9 1 11 2 13 3 1 10 9 1 11 2 11 7 10 9 1 11 2 11 2 13 10 9 0 1 13 9 1 10 9 7 9 1 10 9 0 2
61 1 11 1 12 10 9 2 13 1 10 9 2 13 9 1 11 1 10 9 1 11 1 10 9 1 11 12 1 11 15 13 10 9 1 10 9 2 7 3 1 3 13 15 1 11 7 1 11 2 1 12 2 7 13 10 9 1 9 7 9 2
42 1 10 9 1 10 9 2 15 13 10 9 0 1 11 1 11 1 9 1 12 7 13 1 9 0 15 1 10 0 9 1 9 13 1 10 9 0 1 10 10 9 2
30 13 1 3 1 15 10 9 1 10 9 2 9 1 9 1 9 2 9 1 9 2 9 0 7 9 1 10 9 0 2
15 3 2 10 9 4 13 9 1 9 1 10 11 11 0 2
44 11 2 11 1 10 11 2 13 10 9 1 9 1 10 9 1 0 9 11 2 4 13 1 10 9 0 1 11 10 9 12 1 11 1 12 2 1 10 9 0 1 12 9 2
45 10 9 1 10 9 13 10 9 1 10 9 13 1 10 9 1 11 1 10 9 1 10 9 15 13 10 11 11 11 11 7 10 9 0 16 13 1 11 13 1 0 11 1 11 2
13 13 9 0 7 15 13 1 9 1 10 3 9 2
27 11 13 0 10 9 7 13 1 13 10 9 3 0 7 10 9 7 13 1 12 9 3 1 10 11 11 2
9 10 9 1 10 9 13 11 11 2
12 10 9 1 9 1 10 9 13 1 9 12 2
24 10 9 1 10 9 15 13 3 1 12 9 2 3 3 1 10 9 1 9 0 1 10 9 2
43 10 9 1 10 0 9 13 10 9 1 10 9 0 1 12 9 1 9 0 2 1 10 15 15 13 1 10 12 9 0 16 13 1 9 1 3 1 12 9 10 9 11 2
12 15 13 9 1 10 9 0 1 10 9 0 2
12 11 13 3 9 2 7 3 15 13 1 9 2
28 10 9 9 10 9 1 10 9 16 13 1 10 9 7 16 13 10 2 9 0 0 2 1 13 10 9 0 2
8 2 2 2 10 11 2 2 2
42 10 9 13 0 1 10 12 9 2 3 13 9 1 9 1 10 9 15 15 13 1 10 9 1 9 0 2 0 9 1 10 9 2 0 9 7 9 1 10 9 0 2
39 11 12 3 13 1 10 9 2 1 0 9 2 1 10 9 0 1 11 2 7 10 9 1 10 9 0 1 11 11 7 11 11 2 1 10 9 1 12 2
21 10 9 0 13 3 0 7 0 2 13 1 10 9 7 9 1 10 9 1 9 2
30 1 10 9 1 10 9 9 1 10 11 11 1 11 2 10 9 13 10 9 0 1 10 11 11 1 10 9 0 0 2
41 10 9 13 10 9 0 1 9 1 9 16 13 10 9 1 9 7 10 9 1 10 9 2 2 3 0 2 2 13 11 2 1 10 9 1 10 16 13 9 0 2
31 10 9 3 13 10 9 1 15 16 15 13 12 2 7 3 13 3 0 13 10 9 1 9 16 13 10 9 2 10 9 2
18 7 10 9 13 1 11 11 2 10 9 16 15 13 1 13 15 9 2
27 10 9 4 13 1 3 9 1 10 9 9 1 9 0 7 0 7 15 1 10 10 9 1 10 11 11 2
30 13 12 13 10 9 0 10 15 13 9 3 0 16 13 10 9 2 9 0 2 9 0 2 7 10 9 0 7 9 2
25 1 12 4 13 1 10 0 9 2 0 1 10 9 2 1 10 11 1 10 11 1 10 11 11 2
21 15 1 10 9 3 0 1 10 9 13 10 9 1 11 11 1 11 7 10 9 2
27 15 13 1 10 9 1 9 3 0 1 15 2 10 9 0 7 0 13 0 7 13 7 2 1 9 0 2
35 13 1 10 9 2 10 3 9 11 11 2 1 10 9 1 10 9 1 11 1 11 1 12 2 12 9 3 3 2 1 12 2 13 9 2
37 10 0 9 1 10 9 13 2 10 9 11 2 10 9 11 2 9 1 9 0 1 12 9 2 2 10 9 11 2 10 9 11 11 1 10 11 2
9 1 10 9 3 0 13 10 11 2
26 3 10 9 1 10 9 1 11 2 11 13 13 1 10 9 1 9 7 10 9 1 10 9 1 9 2
77 1 13 13 10 9 1 10 9 1 10 9 0 1 10 9 1 11 2 3 1 10 11 2 11 13 1 10 9 13 1 10 9 1 10 9 7 15 13 1 10 0 11 2 1 10 9 1 11 2 3 4 13 1 10 9 0 1 10 9 7 15 13 13 1 9 13 10 9 1 10 9 1 9 0 1 11 2
19 10 9 13 0 7 0 7 10 9 10 9 7 3 9 1 15 16 13 2
14 3 13 16 13 3 9 0 7 0 2 12 8 2 2
30 13 9 1 0 9 1 9 7 9 7 13 9 1 9 1 9 0 7 0 2 15 16 13 16 3 13 0 9 0 2
18 10 9 13 10 9 0 7 1 15 15 4 13 15 1 10 9 0 2
69 16 7 10 9 4 13 3 1 10 9 1 10 9 1 10 9 2 3 10 10 9 13 1 10 0 9 1 9 2 11 1 10 9 13 3 10 9 1 9 7 9 1 9 0 2 1 13 1 10 3 9 1 9 1 9 0 7 9 0 16 13 10 9 1 10 2 11 2 2
33 1 10 9 2 10 9 0 1 10 9 0 3 13 1 9 1 13 1 10 9 1 10 9 2 3 13 7 10 9 7 9 3 2
18 10 9 13 10 9 0 1 5 12 9 1 10 5 12 1 10 9 2
59 13 10 9 1 10 9 1 10 9 0 1 9 1 10 9 0 0 7 1 10 9 1 10 9 1 9 2 13 9 1 10 9 0 1 10 9 0 10 0 1 9 2 13 16 10 9 0 1 10 9 3 13 15 3 16 13 10 9 2
17 3 15 13 1 9 0 13 10 9 1 10 9 11 11 2 11 2
10 11 3 13 1 11 11 1 11 11 2
23 15 13 1 13 10 9 1 10 9 7 15 13 0 1 10 9 1 11 2 3 13 9 2
41 10 9 1 10 9 13 0 16 15 13 0 7 1 15 16 15 13 3 2 1 9 1 10 9 1 10 9 1 9 2 7 13 3 0 16 15 13 1 10 9 2
24 3 15 13 0 3 13 1 10 9 0 0 2 7 13 1 9 1 10 9 1 9 1 9 2
20 7 10 9 3 0 1 10 9 15 13 2 3 1 11 11 2 1 11 11 2
23 7 3 2 1 9 1 10 9 1 10 9 1 10 9 2 4 13 3 10 9 13 3 2
18 11 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
23 3 4 13 10 9 2 7 15 13 1 10 12 5 1 9 0 2 3 13 15 1 9 2
16 13 3 0 1 10 9 1 9 1 9 2 7 15 7 15 2
19 11 11 2 11 2 12 2 13 10 0 9 0 0 7 9 1 10 9 2
25 11 11 4 13 1 11 11 11 1 11 7 13 1 11 11 7 11 11 2 12 2 12 2 8 2
12 10 0 9 13 10 0 9 1 12 9 11 2
28 10 9 15 13 1 11 2 13 15 10 9 1 13 10 9 1 0 1 13 15 1 11 1 9 1 10 9 2
34 10 9 1 10 9 13 13 15 3 1 12 2 7 4 1 13 15 1 11 2 16 10 0 9 1 9 0 13 10 9 11 7 11 2
21 2 13 3 15 13 2 3 1 10 9 1 11 2 3 1 10 0 9 1 11 2
16 4 13 9 1 10 9 0 1 11 2 11 2 11 7 11 2
8 10 9 3 4 13 1 9 2
81 10 9 13 10 9 1 12 9 2 1 10 9 1 9 3 0 1 10 9 1 10 12 9 1 9 2 13 10 9 0 7 10 9 1 9 1 10 9 1 10 9 1 11 2 10 9 1 10 9 1 10 11 1 10 11 7 1 11 11 7 10 9 0 1 10 12 9 2 3 1 10 9 1 11 2 11 2 11 7 11 2
25 1 10 9 0 7 1 13 10 9 2 11 13 10 9 1 10 9 1 10 9 7 10 9 0 2
16 3 1 16 11 11 13 10 9 1 11 13 15 2 4 13 2
23 15 13 0 9 0 1 9 1 9 7 1 15 10 9 13 10 9 13 1 10 9 0 2
5 3 3 13 15 2
9 13 0 7 0 13 3 1 9 2
14 13 9 1 9 1 9 1 10 12 1 11 1 12 2
43 15 13 1 10 9 2 1 15 15 10 9 2 1 10 15 15 3 4 1 13 2 10 9 2 2 15 13 16 16 11 7 15 4 13 0 13 15 3 9 13 10 9 2
17 1 10 9 1 11 2 10 9 1 0 9 0 13 1 12 9 2
21 11 7 11 13 10 9 0 1 10 15 13 10 9 0 2 9 1 10 11 11 2
10 11 15 13 13 1 11 1 10 9 2
26 11 13 10 9 3 1 10 11 1 15 13 7 4 13 0 1 10 11 1 11 1 10 9 1 11 2
53 1 11 1 12 1 10 12 1 11 1 12 2 10 9 16 13 1 9 1 11 4 13 15 9 1 9 1 10 9 1 11 7 1 0 9 13 3 1 11 1 11 1 11 11 10 0 9 0 1 12 9 0 2
62 1 0 9 10 9 11 11 4 13 10 0 9 1 10 11 11 2 11 1 9 7 12 2 12 9 1 10 16 15 13 1 9 1 10 12 9 1 9 2 10 9 1 10 0 9 2 1 10 9 7 12 9 1 10 0 9 16 13 1 10 9 2
36 10 9 1 10 11 11 15 13 1 10 9 9 1 10 11 11 2 3 13 13 1 11 11 1 10 9 1 10 0 9 1 16 13 10 9 2
7 10 9 1 9 4 13 2
16 10 9 13 10 9 1 9 0 2 10 9 2 3 15 0 2
53 13 9 1 10 9 1 10 9 0 3 3 1 10 9 1 11 11 2 7 1 10 10 9 2 11 13 16 2 10 9 4 13 3 3 2 9 1 16 10 9 1 9 13 10 9 1 9 1 10 9 0 2 2
21 1 10 9 12 13 10 9 1 12 9 1 10 9 0 1 12 9 1 9 5 2
96 15 1 10 0 9 13 10 11 11 7 10 9 11 10 9 0 16 3 13 9 1 10 9 0 16 13 1 10 9 1 10 9 2 3 7 3 13 9 1 10 9 0 1 11 2 11 2 16 13 1 10 9 9 2 3 9 7 9 1 10 9 0 11 11 16 13 9 1 10 9 1 11 1 2 10 9 1 11 2 13 1 10 9 0 15 13 10 9 0 1 10 9 0 1 11 2
57 1 9 1 10 9 1 10 12 9 1 10 9 1 11 13 3 1 11 1 12 10 9 7 9 4 13 1 10 9 16 15 13 7 13 1 10 9 1 10 0 9 2 10 15 13 3 9 4 13 1 10 9 0 1 11 11 2
13 1 15 2 13 10 9 1 10 0 9 2 11 2
10 13 9 1 10 9 1 11 7 11 2
17 1 10 10 9 9 13 10 9 16 13 10 12 9 3 7 3 2
32 10 9 13 1 9 16 4 13 1 13 1 9 0 13 0 1 13 7 13 1 9 0 10 9 0 1 13 10 9 3 0 2
41 13 1 13 10 9 7 3 1 13 12 5 1 9 1 9 1 13 10 9 1 10 9 3 15 13 7 3 15 13 13 10 9 1 3 3 4 15 13 1 9 2
41 3 1 10 0 9 13 4 1 13 1 2 9 2 13 16 3 10 9 0 1 10 9 1 10 9 7 9 0 1 10 10 9 13 1 10 9 1 10 0 9 2
31 10 0 9 2 13 1 11 2 12 9 3 3 2 13 10 9 1 2 10 0 2 2 11 2 10 12 1 11 1 12 2
16 1 9 15 4 13 10 9 13 1 10 9 1 5 7 9 2
19 13 9 1 10 3 9 0 11 7 11 11 2 7 9 1 11 11 11 2
30 13 10 9 1 10 9 0 7 3 3 13 1 10 9 2 2 4 13 1 13 15 7 13 10 9 1 13 15 2 2
14 10 9 13 13 15 1 10 9 1 9 1 10 9 2
46 10 0 9 1 9 9 0 13 1 0 9 1 10 9 1 12 2 1 10 9 1 11 11 2 10 9 11 0 9 1 11 11 16 13 10 9 1 10 9 9 1 10 9 8 0 2
7 13 12 9 1 10 9 2
33 10 9 1 9 1 11 13 3 0 1 9 7 10 1 10 9 1 11 2 4 1 13 1 3 1 12 9 1 9 1 10 9 2
23 10 9 15 15 4 13 11 1 11 12 9 3 2 3 1 13 15 3 13 10 11 11 2
49 10 9 13 1 10 9 1 8 2 1 9 1 10 9 0 2 13 1 9 1 10 9 11 11 7 11 2 1 15 15 13 3 10 9 16 13 10 11 1 11 1 10 11 1 10 11 1 11 2
43 7 1 10 9 10 9 11 11 13 10 9 1 9 1 10 9 1 10 0 9 11 2 7 10 9 1 10 9 1 10 10 9 1 10 9 2 11 11 2 11 11 2 2
43 15 13 10 9 1 10 12 5 10 9 11 11 2 15 13 10 9 1 10 12 5 1 10 9 1 10 9 1 9 1 9 2 16 7 3 3 10 12 5 13 10 9 2
20 1 12 2 13 10 9 1 9 0 2 9 9 2 1 10 9 0 1 11 2
12 13 1 10 9 1 9 0 16 13 10 9 2
46 1 10 9 1 12 10 11 11 15 13 3 2 4 7 13 10 0 9 1 10 0 9 15 1 11 7 11 2 7 1 9 1 10 9 2 13 10 3 1 10 9 1 0 9 0 2
52 13 1 10 9 11 1 11 10 11 11 1 10 9 13 2 11 2 2 12 2 2 1 9 1 11 11 2 10 15 3 1 10 9 13 10 9 1 9 1 9 0 2 10 15 15 4 13 1 9 1 9 2
49 1 10 9 1 11 13 10 9 0 1 9 0 1 10 9 1 10 9 0 2 13 10 9 1 10 9 0 1 12 2 1 9 1 11 11 13 1 11 11 2 11 11 7 11 11 2 1 15 2
29 16 10 9 1 11 1 11 13 10 9 0 1 13 1 10 9 12 2 12 2 11 13 1 15 1 10 9 0 2
30 1 10 9 10 11 11 13 1 10 0 9 10 9 1 10 9 0 1 10 11 11 2 3 9 1 10 11 1 11 2
21 11 13 10 9 7 9 0 1 10 9 1 11 2 9 1 11 2 1 12 9 2
23 10 9 2 16 4 1 13 9 1 10 0 9 11 11 2 13 10 9 12 1 10 9 2
17 1 9 1 9 15 4 13 0 2 1 9 1 10 9 13 0 2
33 16 13 10 0 9 16 10 9 13 1 11 11 11 12 2 11 11 11 11 11 2 11 11 12 3 13 10 9 0 1 10 9 2
26 10 11 11 13 10 9 1 9 0 13 1 10 9 11 12 9 12 1 10 9 0 1 10 9 0 2
23 11 11 11 2 11 11 2 11 2 12 1 11 1 12 2 13 10 9 0 1 9 0 2
9 13 1 10 9 1 11 7 11 2
15 1 12 13 1 10 11 11 2 1 10 15 13 12 9 2
36 10 9 2 7 9 2 13 10 9 0 2 1 15 1 10 9 1 10 9 0 2 7 3 1 15 13 1 10 13 2 9 1 10 9 2 2
10 10 0 9 15 13 0 1 10 8 2
23 3 15 13 10 9 1 10 9 0 2 0 2 7 3 1 10 9 3 0 2 11 11 2
15 10 9 1 10 9 1 9 3 13 10 9 1 10 9 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
28 15 8 4 13 1 10 9 1 9 15 16 15 13 1 10 0 9 1 9 7 10 0 9 1 13 10 9 2
32 11 11 2 10 9 1 11 13 10 9 1 10 9 11 1 10 9 11 11 2 10 9 1 9 1 11 13 1 10 9 12 2
10 3 2 1 13 10 9 1 11 11 2
30 1 10 9 1 12 9 2 13 10 9 0 1 4 13 1 10 9 1 10 12 9 16 13 10 12 9 1 10 11 2
16 2 11 11 11 2 11 11 11 11 7 11 11 11 11 2 2
14 15 4 13 1 9 1 10 9 0 1 11 7 11 2
41 10 11 11 1 11 12 2 1 10 15 13 1 9 10 11 10 11 2 13 10 9 0 13 1 10 3 11 11 1 11 2 3 2 11 11 1 11 11 11 2 2
53 15 13 1 10 9 0 3 1 9 2 3 1 9 2 3 1 9 0 2 3 1 9 0 1 10 8 2 9 7 1 10 9 2 1 10 9 0 2 13 1 13 10 8 2 9 2 3 3 3 13 10 9 2
34 2 11 11 2 2 1 9 2 2 9 0 2 2 13 10 9 1 10 9 7 9 0 11 11 2 8 9 1 10 9 0 11 11 2
7 13 13 0 1 11 11 2
27 13 10 9 1 10 9 1 9 0 7 0 1 13 3 10 9 1 9 1 10 9 1 13 1 10 9 2
47 13 3 2 16 10 9 11 1 11 2 13 9 1 11 11 11 2 15 1 10 9 1 10 9 1 11 13 1 13 10 0 9 1 9 11 7 10 9 11 11 2 9 1 10 9 0 2
16 15 13 10 11 2 1 10 9 1 11 7 1 9 1 9 2
40 10 9 1 10 9 13 1 10 9 11 11 11 2 9 1 10 9 1 10 9 11 11 15 13 1 10 11 11 11 11 1 10 9 1 10 9 12 7 12 2
38 13 0 1 9 0 1 10 15 13 13 3 1 12 9 0 2 16 1 10 9 13 12 0 2 4 1 13 3 1 12 9 2 3 1 12 9 0 2
33 10 9 0 13 13 10 9 0 3 0 1 11 1 10 0 9 2 7 15 1 10 0 9 1 10 9 0 1 9 7 9 11 2
31 10 11 4 13 3 1 10 9 1 12 13 11 11 11 2 11 2 0 1 11 11 11 11 7 10 11 1 10 11 11 2
21 10 9 13 10 9 0 2 1 12 9 1 9 7 12 1 9 2 13 12 9 2
31 3 2 11 13 1 9 0 10 1 11 2 1 9 1 10 15 13 10 9 1 10 9 2 11 2 11 7 11 2 2 2
36 15 4 13 1 10 0 9 0 1 10 9 1 11 1 3 1 10 9 1 10 9 13 1 10 0 9 1 13 15 1 11 1 10 9 0 2
20 3 2 4 13 10 9 1 9 1 9 1 9 0 2 10 9 0 1 9 2
33 1 9 1 10 10 9 0 1 9 1 11 2 11 2 10 9 13 0 1 9 1 9 0 2 7 3 2 15 13 10 9 0 2
6 13 7 3 13 0 2
18 10 11 11 1 11 13 10 9 1 9 1 10 11 11 11 1 11 2
21 15 13 16 4 4 13 1 10 9 1 13 1 11 2 10 9 3 0 1 11 2
26 10 9 13 13 10 0 9 1 10 9 1 9 1 9 16 10 9 0 1 10 11 3 4 3 13 2
33 10 9 1 9 1 10 11 11 2 3 1 9 1 10 9 2 13 1 10 9 0 0 13 10 0 9 1 10 9 1 10 9 2
46 1 10 9 2 15 10 9 1 10 9 0 1 10 9 7 10 9 1 9 1 9 2 10 9 0 2 4 4 13 1 9 7 9 1 10 0 9 1 10 2 9 2 1 10 9 2
29 10 11 13 10 0 9 1 9 7 10 12 2 11 7 13 10 9 1 12 9 2 12 9 2 1 10 9 0 2
34 10 9 1 12 7 12 13 1 15 2 2 10 9 1 10 9 13 3 10 9 7 10 9 2 15 13 1 9 1 10 9 1 9 2
37 4 13 10 0 9 1 10 9 1 10 9 1 9 1 10 9 1 11 2 0 1 10 9 1 10 11 16 15 13 3 1 10 9 1 10 9 2
39 1 9 2 10 9 1 9 0 16 3 4 1 13 15 3 1 12 9 1 10 9 2 13 12 9 10 9 1 10 11 12 2 12 9 7 12 9 2 2
24 11 15 13 1 12 9 2 8 2 1 0 8 2 2 1 10 15 12 13 10 9 1 9 2
20 10 9 13 0 9 7 9 2 7 13 9 1 10 9 3 1 10 9 11 2
13 4 13 9 1 9 1 0 9 1 10 9 0 2
33 1 13 9 1 9 2 11 13 16 10 9 1 11 13 3 10 0 9 7 10 9 1 11 2 7 3 13 1 10 9 3 0 2
14 11 13 10 9 1 9 13 1 11 1 10 9 12 2
18 15 13 1 9 1 10 9 1 11 11 1 11 1 10 9 1 11 2
16 10 11 1 11 11 11 7 11 11 1 10 11 11 1 11 2
16 1 15 13 9 1 10 9 1 11 1 9 1 11 1 12 2
53 3 4 13 1 10 9 1 9 1 10 11 11 11 1 10 8 11 7 10 8 11 1 15 2 1 7 1 12 13 15 1 10 0 9 1 9 1 10 11 11 11 11 2 9 1 10 15 13 1 12 1 12 2
45 10 9 3 13 10 9 1 10 9 0 2 3 7 1 9 0 2 13 1 10 9 1 10 9 1 10 9 1 11 2 3 10 9 1 10 9 15 13 1 10 9 1 12 9 2
37 10 9 1 10 9 13 10 9 2 13 0 2 7 1 11 11 10 9 1 11 13 0 7 3 4 7 4 13 15 1 15 3 16 13 10 9 2
16 2 3 2 3 15 13 1 15 2 13 15 16 3 15 13 2
11 10 9 1 10 9 13 10 9 1 11 2
22 1 9 12 9 0 13 16 15 4 1 13 10 9 1 10 9 16 3 3 15 13 2
25 10 9 1 10 9 0 13 1 11 11 11 7 11 11 4 13 2 7 4 4 13 1 11 11 2
13 10 0 9 0 13 11 2 11 2 11 7 11 2
19 10 16 13 1 8 13 16 3 13 10 8 0 1 11 7 1 10 9 2
32 11 11 2 11 1 11 11 2 13 10 9 0 1 10 9 0 11 13 1 9 13 0 1 9 0 2 9 7 9 1 9 2
20 11 4 13 1 10 0 9 1 10 11 1 12 2 13 10 12 5 9 0 2
18 10 0 9 1 10 9 13 1 10 9 13 1 8 9 1 11 11 12
18 1 10 9 3 15 13 1 10 0 16 13 10 9 1 10 9 12 2
18 11 11 15 13 1 10 9 2 10 0 9 1 9 7 10 9 0 2
20 15 13 16 1 11 11 10 9 3 13 9 1 10 9 7 13 16 13 0 2
21 3 0 7 0 16 13 10 15 1 13 7 3 15 4 13 2 3 1 10 3 2
75 16 11 9 13 10 0 9 1 8 16 3 13 13 10 9 2 9 16 13 1 16 10 9 0 11 9 1 10 9 0 1 9 1 10 9 2 2 10 9 1 10 9 1 9 1 9 13 10 9 0 2 10 9 15 13 3 1 10 9 2 13 10 10 9 1 9 2 7 10 9 1 0 0 2 2
59 1 10 12 9 2 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
17 15 13 1 3 1 10 0 11 7 3 13 13 15 1 16 13 2
45 10 11 11 1 11 13 10 9 0 13 1 10 9 1 11 2 11 2 13 10 9 1 9 1 10 9 1 10 9 1 9 0 1 10 11 11 11 1 10 11 11 11 2 11 2
19 1 10 9 12 13 10 9 0 2 11 8 9 2 3 3 1 11 11 2
18 10 9 0 13 1 0 2 9 1 10 9 0 13 1 10 9 11 2
19 4 7 13 15 10 9 1 12 9 16 15 15 13 10 9 1 10 9 2
42 13 3 1 9 2 9 2 9 2 9 2 11 2 9 1 9 2 9 13 1 9 2 9 0 2 9 2 9 0 1 9 2 9 2 9 1 9 1 9 7 9 2
15 13 1 11 1 9 0 16 10 8 11 13 9 1 9 2
46 13 0 16 2 1 9 2 10 9 1 9 0 3 13 1 11 2 7 3 3 9 16 15 13 1 9 0 1 9 2 13 1 9 16 10 0 9 1 10 9 0 0 13 9 0 2
20 13 1 11 1 12 1 10 9 1 10 9 0 2 1 10 16 13 10 9 2
18 10 9 13 10 9 16 13 10 9 1 10 9 7 9 1 10 0 2
34 10 9 0 11 11 2 1 9 1 10 9 11 13 13 9 1 10 9 0 1 11 2 13 1 10 9 10 9 0 1 11 7 11 2
43 10 9 0 13 1 16 1 10 13 10 9 1 11 15 13 10 9 1 9 0 1 11 2 13 1 0 9 10 9 1 9 1 10 9 9 16 15 13 0 1 10 9 2
18 3 15 13 9 3 9 1 9 0 2 9 2 9 2 9 7 9 2
17 11 13 10 9 7 11 13 10 9 1 10 9 1 11 1 12 2
47 10 9 1 9 1 10 9 1 9 13 1 10 9 2 7 1 9 1 10 9 15 13 9 1 12 11 11 13 1 10 9 1 12 9 2 16 10 9 13 1 10 9 0 1 10 9 2
35 10 9 1 11 11 1 11 15 13 1 10 9 1 9 1 11 0 1 10 9 1 11 1 11 7 1 15 1 10 9 1 10 11 11 2
33 10 9 0 11 10 11 13 0 1 13 10 9 1 11 7 10 9 11 1 11 2 16 13 1 11 1 11 7 3 13 1 11 2
37 7 3 10 9 1 10 9 3 4 13 0 9 1 15 9 1 10 9 2 1 12 15 13 10 9 0 0 2 10 16 3 15 13 1 10 9 2
16 1 10 9 11 1 11 13 10 9 7 15 13 1 10 9 2
48 13 10 9 1 16 11 15 13 10 9 1 11 1 11 7 16 15 13 10 9 7 1 10 9 15 13 2 15 16 13 10 10 9 7 1 10 0 9 13 10 9 1 11 7 1 10 9 2
38 10 9 13 10 9 16 13 10 9 1 10 9 0 7 10 9 0 2 16 13 10 9 1 10 9 1 9 0 7 2 7 1 10 9 1 10 9 2
35 1 10 9 3 15 15 9 10 9 1 11 2 10 9 1 11 11 2 13 1 11 11 11 7 13 1 10 11 1 11 1 11 1 11 2
33 10 9 2 13 1 11 11 11 2 13 1 12 2 16 16 10 9 2 1 9 0 2 13 1 12 7 13 9 1 11 11 11 2
13 9 7 9 1 10 9 16 15 13 1 10 9 2
14 1 9 13 9 0 7 13 9 7 13 1 10 9 2
39 11 11 11 2 11 2 10 11 2 12 2 9 0 16 13 1 10 2 9 0 2 1 11 1 11 13 10 9 13 1 10 11 11 1 11 2 11 2 2
17 10 9 0 15 13 1 10 9 1 11 11 12 2 11 11 11 2
20 10 9 0 1 10 9 11 13 10 9 2 13 1 10 9 1 10 9 0 2
25 10 9 3 15 13 7 15 13 1 10 9 0 1 10 9 16 13 1 9 0 7 9 9 0 2
44 1 9 3 4 7 13 10 9 1 10 9 1 9 1 10 0 9 2 7 1 10 9 1 10 9 0 1 10 9 1 10 9 2 13 15 1 15 1 10 9 0 1 11 2
15 15 13 16 11 15 13 1 11 13 10 9 1 11 11 2
28 1 12 10 9 4 13 2 7 1 3 10 11 1 11 4 13 15 1 10 9 3 0 1 10 9 1 11 2
13 15 13 12 9 1 10 9 11 1 12 7 12 2
43 16 10 9 1 11 11 2 11 11 4 13 1 10 9 2 10 10 9 4 13 1 10 9 1 9 11 11 2 16 15 13 1 9 0 3 3 1 10 9 1 10 9 2
11 1 10 9 13 10 9 9 0 2 9 2
42 10 9 13 9 1 10 9 1 10 9 7 3 1 12 2 1 9 1 10 9 1 9 16 13 1 10 9 1 11 2 15 13 1 9 9 0 1 11 7 10 9 2
24 15 13 13 10 9 0 1 9 16 13 10 9 0 7 3 15 13 9 1 10 13 10 9 2
36 10 9 1 10 9 13 16 10 9 11 13 3 2 1 9 7 9 16 13 16 3 13 10 9 1 13 15 1 10 9 16 7 13 10 9 2
22 11 11 2 8 8 2 2 11 1 10 11 12 2 11 12 2 2 9 7 9 0 2
19 15 13 1 10 9 1 10 11 11 1 10 9 1 11 2 11 11 11 2
21 13 0 7 9 1 10 0 9 0 10 11 11 1 10 10 0 9 2 12 2 2
27 1 9 0 13 16 13 10 10 9 7 13 10 0 9 1 9 7 9 1 9 2 15 1 9 7 0 2
19 10 9 1 10 9 13 10 9 1 10 9 11 11 11 11 11 11 11 2
20 10 9 0 11 11 13 12 9 1 12 2 10 15 4 13 1 9 1 11 2
18 13 1 10 9 1 10 9 2 7 1 10 9 15 13 1 9 0 2
8 11 13 10 9 0 1 12 2
18 13 1 9 7 10 9 0 13 10 11 1 11 1 10 0 9 0 2
15 3 1 10 9 13 9 3 1 10 9 11 7 10 9 2
28 10 9 3 13 1 0 9 13 1 10 11 11 3 13 9 1 10 0 9 1 10 9 16 15 13 10 9 2
19 1 15 10 9 1 11 1 10 0 9 1 11 13 10 0 9 1 9 2
9 11 11 15 13 13 1 10 9 2
4 13 1 11 2
25 3 15 13 0 16 16 13 10 9 15 13 10 8 7 16 13 10 9 1 9 1 9 1 0 2
14 10 0 9 0 13 0 9 7 10 0 9 1 9 2
13 15 13 1 11 1 10 9 0 13 1 10 9 2
39 3 1 9 1 10 11 1 11 11 2 11 10 0 9 7 11 11 9 3 13 1 10 9 1 9 7 1 9 1 9 1 11 7 11 9 13 16 13 2
59 11 4 13 10 9 1 9 1 10 9 3 0 3 7 3 1 11 2 9 1 12 7 12 9 1 9 0 3 13 0 13 1 10 9 2 10 9 2 13 10 9 2 13 15 1 9 1 10 8 2 8 7 13 13 10 9 1 9 2
35 13 3 1 10 11 11 1 10 11 11 1 11 12 1 11 11 2 11 2 8 2 7 13 1 10 11 12 1 11 2 11 2 8 2 2
27 3 13 10 9 0 2 1 9 1 11 11 2 10 9 7 0 9 1 10 9 1 10 9 0 11 11 2
14 10 9 13 3 0 7 0 1 10 0 7 10 9 2
24 1 10 9 13 10 9 1 10 9 2 10 9 0 2 10 9 0 7 10 9 1 12 9 2
23 2 11 2 13 3 3 10 9 0 1 10 9 1 0 2 0 7 0 2 2 13 11 2
29 3 2 1 7 15 13 1 8 7 8 1 9 1 10 9 8 2 11 11 15 2 13 2 3 1 9 3 9 2
27 1 10 9 12 2 11 2 3 1 10 9 1 9 2 13 10 0 9 2 1 10 9 0 1 11 11 2
34 3 10 9 0 15 13 1 11 7 15 13 13 11 2 4 13 15 13 10 9 2 7 3 13 0 1 10 9 2 3 13 1 12 2
5 11 13 1 9 2
27 3 2 13 1 10 9 3 0 7 3 4 13 13 9 0 1 15 1 15 2 16 10 9 13 3 0 2
20 9 10 1 9 2 9 0 2 7 10 9 1 9 0 1 9 13 13 0 2
19 10 9 1 10 9 13 1 11 11 2 9 7 9 1 8 2 7 9 2
17 5 12 1 10 12 9 3 13 1 10 9 12 2 13 10 12 2
13 15 13 10 9 1 11 7 10 9 13 1 11 2
43 1 10 9 2 1 11 1 12 2 11 11 2 11 2 13 10 9 1 13 7 13 9 1 10 9 1 11 2 16 1 3 4 13 10 9 1 11 2 7 1 9 0 2
21 13 3 0 7 15 1 10 9 1 11 12 16 3 15 4 13 1 16 15 13 2
5 13 9 7 9 2
25 13 9 1 9 2 9 7 9 2 7 4 13 1 10 9 0 15 13 1 15 9 1 10 9 2
27 1 10 9 16 10 9 1 10 9 13 10 9 1 9 1 9 16 2 13 10 9 2 4 13 9 0 2
15 10 9 1 9 13 3 1 10 9 1 9 1 9 0 2
32 10 11 11 1 11 1 9 4 4 13 1 11 7 9 2 13 9 13 1 10 11 11 1 11 2 1 10 9 1 12 9 2
66 16 11 3 15 4 13 7 16 4 13 1 9 10 9 2 3 13 9 2 3 13 10 9 1 10 9 7 9 3 3 2 16 13 16 10 9 13 13 10 12 8 7 15 13 1 10 9 1 10 9 13 3 13 15 10 9 1 10 9 16 13 1 10 0 9 2
8 10 9 13 16 15 4 13 2
33 15 13 10 9 1 10 15 4 1 13 15 10 9 0 2 10 9 13 10 9 2 9 1 9 2 10 9 1 9 1 10 9 2
72 10 0 9 1 10 11 11 12 2 12 13 0 2 3 7 10 9 4 4 13 1 13 10 9 16 13 15 3 1 10 9 1 15 7 13 16 15 13 3 1 10 9 11 10 9 7 15 1 9 1 13 10 9 16 13 15 0 1 15 1 10 11 11 16 1 10 9 1 10 9 0 2
29 3 1 10 9 0 15 13 2 1 10 9 11 11 2 10 9 1 10 11 2 9 1 9 1 10 9 0 2 2
36 11 13 16 10 9 4 13 1 13 1 9 1 9 1 16 13 16 10 9 3 3 4 4 13 1 9 1 9 13 1 10 0 9 1 9 2
54 1 10 9 3 3 15 13 10 9 1 9 0 2 9 0 2 7 15 1 9 0 2 9 0 2 2 7 3 10 9 0 1 9 2 9 1 9 7 3 10 9 1 9 3 15 13 9 7 10 9 1 9 0 2
24 10 2 11 11 11 2 13 10 9 0 1 12 5 5 5 7 10 9 1 12 5 5 5 2
34 10 9 0 3 3 13 9 0 2 9 4 13 16 3 1 10 9 1 10 9 1 10 11 11 13 9 1 10 9 1 13 10 9 2
14 10 0 9 1 10 9 4 13 1 11 11 1 12 2
7 15 13 1 11 2 11 2
43 1 10 11 1 10 11 0 2 10 9 13 9 2 3 0 1 10 9 0 2 4 13 1 9 0 2 0 2 10 9 2 15 1 10 9 1 10 11 2 7 1 11 2
40 10 9 1 9 0 7 9 0 1 11 13 3 9 1 9 1 9 1 10 9 2 13 7 4 13 1 10 9 10 9 1 10 9 0 1 13 16 13 13 2
22 15 13 1 10 9 7 11 0 1 3 2 1 10 9 1 3 7 1 10 9 1 3
18 3 2 10 9 13 1 10 9 1 9 7 9 13 1 9 3 0 2
17 1 12 2 11 13 10 9 0 7 3 4 13 9 1 12 9 2
21 10 9 0 1 12 2 13 10 0 9 0 13 1 9 1 10 13 9 1 11 2
35 11 12 11 13 9 13 3 1 11 2 11 2 11 2 11 2 11 2 11 2 0 11 2 11 2 9 1 11 11 7 9 1 11 11 2
67 2 15 13 0 16 15 16 4 13 13 2 1 10 9 2 10 9 1 10 9 2 0 2 2 1 10 9 7 1 10 9 1 9 2 3 13 9 16 15 13 9 2 2 13 11 11 2 9 1 10 9 9 2 16 13 1 9 2 9 7 9 2 8 2 1 11 2
63 1 10 12 9 2 10 9 1 11 11 4 13 1 10 12 5 9 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
33 1 10 9 2 10 9 1 10 9 4 13 1 10 9 1 10 0 9 16 13 10 12 1 11 1 12 1 15 9 1 10 11 2
40 1 10 9 4 13 15 1 10 9 1 10 9 0 2 7 10 9 13 0 1 10 9 7 3 3 1 10 9 0 2 16 13 0 13 9 0 1 0 9 2
24 11 13 10 9 0 2 0 1 12 9 13 10 12 1 11 2 13 10 0 9 7 9 0 2
47 1 10 9 1 10 11 1 10 11 15 13 1 10 9 2 13 15 1 9 1 10 9 1 12 1 9 1 10 9 16 13 1 10 9 0 1 3 2 13 10 9 1 9 1 10 9 2
5 15 13 1 11 2
17 10 0 9 1 9 1 9 2 9 7 9 13 10 9 1 11 2
55 13 9 0 1 10 9 1 11 7 11 16 15 13 1 9 13 1 10 11 11 1 9 1 10 9 12 2 16 13 1 12 9 0 16 15 13 1 10 9 1 11 2 11 1 11 2 11 11 1 11 7 11 1 11 2
9 1 11 13 1 10 9 1 11 2
15 1 9 2 13 0 16 15 13 9 3 1 10 9 0 2
10 10 9 1 12 13 1 12 12 9 2
15 1 10 9 12 13 1 12 9 2 13 1 10 9 0 2
17 13 1 9 1 10 9 1 10 9 1 11 1 10 9 1 12 2
27 3 1 15 2 15 13 10 9 1 10 9 0 1 10 9 7 1 10 9 0 1 10 9 1 10 9 2
38 11 11 13 1 10 9 7 10 9 0 9 1 9 7 13 1 10 9 2 1 10 9 1 10 9 0 2 10 9 1 9 0 1 10 9 1 9 2
21 10 9 13 16 10 9 3 13 10 9 1 9 1 13 10 9 1 10 11 12 2
37 1 11 1 12 2 11 13 10 9 1 12 9 7 0 1 15 1 10 9 1 11 2 10 11 11 2 9 16 15 13 10 9 0 1 10 11 2
28 10 9 1 10 9 4 13 0 2 1 9 1 16 10 0 9 0 4 13 1 9 10 9 0 1 10 9 2
11 13 9 0 1 10 11 1 11 1 11 2
54 10 9 1 9 3 13 10 9 1 10 9 3 1 9 1 10 12 5 2 16 1 10 9 10 9 15 13 1 10 9 0 16 1 10 13 15 13 10 9 1 9 0 2 7 3 0 7 0 13 10 9 1 9 2
35 15 13 16 13 10 9 7 10 9 2 3 13 10 9 0 7 9 3 0 1 9 1 13 15 10 9 2 2 13 10 9 1 10 9 2
28 10 9 1 11 13 10 9 16 13 10 0 9 1 10 9 2 11 11 2 7 3 13 9 1 10 1 3 2
22 10 9 15 13 1 9 7 15 13 9 2 7 10 9 4 13 3 2 13 10 9 2
45 1 10 9 2 9 13 0 13 0 13 0 2 13 3 12 9 1 9 2 2 0 2 7 2 13 2 2 7 13 12 9 2 12 9 2 0 2 7 12 9 2 13 2 2 2
50 1 15 15 13 10 9 0 2 3 2 1 9 2 9 0 7 0 2 9 0 7 0 1 2 9 0 0 2 2 2 13 10 9 1 10 9 2 2 7 9 16 3 4 7 13 1 10 9 0 2
37 11 11 11 11 2 11 2 11 2 11 1 12 2 11 2 11 1 12 2 13 10 9 2 9 7 9 0 1 0 9 1 10 11 7 10 11 2
6 10 9 1 10 11 2
24 1 12 10 11 13 13 15 1 10 11 11 13 10 9 1 11 1 9 1 10 9 11 11 2
21 13 1 10 9 1 13 9 1 9 7 1 13 10 9 1 10 9 0 7 0 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
79 1 10 9 1 10 9 0 1 10 9 1 10 9 2 13 1 11 1 12 2 10 9 1 11 11 11 13 10 9 1 10 9 1 10 9 1 11 11 1 13 2 10 9 0 1 13 9 2 7 13 10 0 9 1 10 0 9 1 10 9 2 11 11 2 1 9 2 0 1 10 9 2 1 9 2 9 7 9 2
21 11 1 11 2 15 13 10 14 11 10 11 2 3 15 13 10 9 0 11 11 2
12 4 13 7 13 1 2 9 1 9 0 2 2
13 15 13 10 9 1 10 9 1 9 7 10 9 2
39 10 1 10 9 13 0 1 10 12 1 11 1 12 1 15 4 13 1 11 10 9 1 10 9 0 11 1 11 2 1 0 9 1 10 9 11 11 11 2
32 3 13 1 13 9 1 11 1 10 9 1 9 1 10 9 1 11 11 2 10 9 0 7 3 0 16 3 13 1 10 9 2
21 11 13 10 9 1 10 9 7 0 7 15 13 10 9 7 15 4 13 10 9 2
13 7 3 15 13 1 10 9 16 15 13 10 9 2
30 1 9 1 11 2 10 9 13 2 10 9 0 1 9 0 2 16 13 10 9 0 13 7 13 1 15 1 10 9 2
59 1 10 12 9 2 11 4 13 1 10 12 5 0 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
15 1 9 13 0 9 2 3 7 3 0 2 1 10 9 2
43 10 9 3 2 11 11 4 13 1 10 9 1 10 11 11 11 2 1 9 1 11 11 2 9 0 2 15 4 13 10 9 7 9 1 11 11 1 10 9 0 1 11 2
38 13 10 9 1 10 9 0 2 3 15 13 10 0 9 1 10 9 2 3 9 1 10 9 1 10 9 16 15 13 1 10 9 16 13 10 9 0 2
27 1 10 11 1 11 10 9 2 1 10 9 1 10 11 11 2 4 13 1 11 7 10 9 0 4 13 2
34 10 9 1 11 15 13 1 10 12 1 10 9 1 11 11 2 15 16 13 16 1 11 10 9 13 1 9 7 10 9 1 10 11 2
23 10 15 2 13 11 11 11 2 13 10 9 1 9 0 2 1 9 1 10 0 9 11 2
29 10 9 13 1 10 9 0 10 9 0 16 13 1 10 9 7 13 10 9 1 13 1 10 9 0 1 10 9 2
14 11 13 1 10 11 11 1 10 11 11 11 1 12 2
30 10 0 9 0 13 3 0 1 13 1 10 9 0 1 10 9 2 1 9 2 15 13 10 9 0 7 10 0 9 2
34 1 10 9 2 15 13 3 16 13 10 9 0 1 11 7 11 2 10 15 15 13 2 16 13 10 9 1 10 9 2 1 10 9 2
25 1 9 1 10 12 5 1 10 9 7 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
51 10 12 1 11 1 12 12 1 10 9 4 13 1 10 9 0 11 11 2 11 2 13 12 11 1 10 9 2 13 10 12 9 3 1 9 1 10 11 11 3 7 11 4 3 13 12 3 1 10 9 2
50 10 9 1 10 9 13 2 2 15 1 10 9 7 9 13 1 10 9 13 1 10 9 0 2 2 7 15 13 10 9 1 10 9 0 1 10 9 1 10 9 0 2 16 15 13 1 10 9 13 2
24 11 13 10 9 7 9 0 1 10 9 1 11 2 9 1 11 2 11 11 2 1 12 9 2
28 10 11 11 11 11 2 3 13 1 11 11 2 13 10 9 1 9 1 11 2 1 10 9 1 11 2 11 2
36 10 9 1 11 13 1 13 10 9 13 10 9 11 2 15 13 13 1 11 2 1 13 16 13 10 9 2 16 15 13 15 10 9 1 11 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
23 11 13 10 9 13 1 10 9 13 1 10 9 1 11 11 1 10 9 0 1 11 11 2
4 13 12 9 2
10 3 4 4 1 13 16 13 1 11 2
33 10 9 1 9 13 1 10 9 1 10 9 0 1 9 2 0 11 2 15 13 1 12 9 1 11 2 10 12 5 9 1 11 2
20 15 13 16 10 9 1 9 13 10 0 9 1 9 1 10 9 7 10 11 2
13 13 1 10 9 16 13 9 1 10 9 1 9 2
58 12 9 0 2 1 10 11 11 5 12 2 8 12 2 2 10 9 11 11 13 10 9 1 10 9 7 10 9 1 16 10 2 9 1 9 0 2 3 13 10 9 1 10 9 2 7 3 10 9 16 2 13 10 0 9 0 2 2
8 3 2 13 0 0 1 12 2
25 15 13 11 11 2 13 10 0 9 1 10 9 11 11 2 13 1 12 1 10 11 1 10 9 2
61 10 0 9 13 10 0 9 0 1 10 9 2 7 13 15 1 10 9 16 4 13 3 9 7 9 1 10 9 1 10 0 9 2 2 13 11 11 11 2 9 1 10 9 11 10 11 2 0 9 0 13 10 9 7 9 1 10 9 1 11 2
14 2 1 3 1 10 3 9 3 15 15 13 13 9 2
30 11 13 1 11 1 9 1 11 13 1 11 11 7 13 3 1 11 11 2 9 1 11 7 9 2 1 11 11 0 2
13 1 10 9 13 10 9 0 7 4 7 13 15 2
17 1 12 10 9 13 1 9 1 10 11 11 1 11 1 10 11 2
16 1 10 9 8 4 13 1 10 0 9 1 10 11 11 11 2
23 1 15 2 15 13 10 9 1 10 9 2 9 3 1 16 1 11 15 13 10 9 0 2
38 10 11 1 10 11 2 3 2 11 11 7 11 1 10 11 2 13 10 9 9 0 16 15 13 1 10 9 0 1 10 11 2 1 10 9 1 11 2
61 1 15 2 10 9 4 13 1 9 1 3 1 10 0 9 1 9 1 10 9 11 7 11 11 11 2 3 15 3 15 13 1 11 16 16 13 16 10 9 0 13 1 10 9 2 1 10 9 0 2 13 1 9 1 9 7 1 9 1 9 2
12 13 9 1 9 0 2 0 7 13 12 9 2
31 1 10 0 9 1 10 9 0 1 12 7 10 9 1 10 12 1 11 1 12 2 11 13 10 0 9 1 10 9 0 2
19 11 11 1 10 11 11 1 11 11 2 13 16 2 13 9 1 10 9 2
10 13 10 9 0 1 11 1 10 11 2
10 10 9 1 11 11 15 13 1 12 2
26 1 12 1 12 2 11 13 10 0 8 9 2 11 11 11 11 2 13 1 11 11 2 11 11 2 2
81 11 11 1 11 7 11 11 1 11 2 10 11 1 11 11 2 11 2 12 1 11 1 12 2 11 2 11 11 2 12 1 11 1 12 2 13 10 9 1 11 1 9 1 9 11 1 9 16 1 10 13 9 15 13 1 9 0 1 11 7 9 1 12 1 12 7 9 9 1 11 1 12 1 12 1 10 9 1 10 9 2
16 3 10 9 13 13 1 12 9 2 12 9 0 7 12 0 2
30 7 16 3 13 10 12 9 1 3 9 2 3 0 2 10 9 3 7 13 10 9 0 13 1 10 0 9 16 13 2
30 11 11 11 13 10 9 1 10 9 1 11 11 16 15 13 1 9 1 10 9 11 1 10 9 11 1 10 9 12 2
33 1 10 9 2 10 9 1 9 15 13 1 9 0 2 16 13 10 9 0 1 9 1 9 1 10 9 1 10 9 1 10 9 2
43 1 12 13 1 11 11 10 0 9 0 2 11 11 2 7 10 0 9 13 10 9 1 12 1 10 11 11 1 11 2 11 2 13 1 10 9 1 10 9 1 10 9 2
14 4 1 4 13 7 13 1 10 9 1 10 12 9 2
28 1 10 0 9 0 15 13 1 11 7 11 10 0 9 2 1 10 15 15 13 1 11 16 4 1 13 15 2
21 1 10 0 9 15 13 10 9 16 15 4 13 2 1 9 0 1 3 0 9 2
13 13 10 12 1 11 1 12 1 11 2 11 2 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
28 10 9 13 10 9 3 0 1 11 1 12 2 7 15 13 3 12 5 1 3 1 10 9 1 11 1 12 2
12 1 10 11 3 15 13 10 9 1 10 9 2
21 13 10 9 11 1 10 9 2 1 9 13 7 10 9 13 0 1 10 0 9 2
19 11 11 13 10 9 1 9 0 1 10 9 11 1 10 9 1 10 11 2
19 15 13 1 15 1 10 9 16 13 2 10 9 1 10 0 9 0 2 2
36 11 2 11 13 10 9 7 9 0 2 1 10 9 1 11 2 11 2 9 1 11 2 1 10 9 1 11 2 11 2 11 7 9 1 11 2
52 3 13 9 1 9 1 10 9 0 2 10 9 3 15 13 1 9 7 3 1 10 9 2 7 10 0 9 13 10 0 9 1 9 1 10 13 15 1 10 9 1 10 9 16 13 15 16 13 1 10 3 2
19 3 15 13 10 9 1 10 9 0 7 9 9 1 10 11 1 10 11 2
16 3 2 10 9 0 15 13 2 11 1 11 7 1 11 2 2
31 10 11 11 11 13 1 10 9 10 9 1 0 9 0 7 1 12 13 10 3 0 2 4 3 13 1 10 11 11 11 2
28 10 9 13 16 9 1 10 11 13 1 9 1 9 1 9 15 13 13 10 9 16 13 2 9 2 3 13 2
15 13 10 9 3 0 1 10 9 11 7 11 11 1 11 2
29 15 15 13 1 10 11 2 12 2 7 1 9 1 11 2 11 13 13 1 10 9 2 16 11 15 13 10 9 2
10 3 3 13 13 10 9 1 10 11 2
49 10 9 1 9 13 10 9 0 2 7 10 9 1 9 3 7 10 9 0 2 12 9 1 9 2 15 1 10 9 3 0 1 10 9 1 10 9 1 10 9 12 2 13 1 15 10 9 0 2
28 11 2 15 13 10 9 13 1 10 9 0 2 15 13 3 3 2 7 13 1 11 1 10 9 1 10 9 2
9 11 13 10 9 1 10 9 0 2
7 3 13 9 16 13 9 2
18 15 13 10 9 1 11 7 13 10 9 1 9 2 9 1 10 9 2
47 10 0 9 13 10 11 2 12 2 16 13 1 10 9 1 10 11 2 12 1 11 11 2 7 13 1 10 9 13 11 2 11 2 10 9 1 11 11 7 10 9 1 10 11 2 12 2
35 10 9 0 1 13 10 9 13 13 10 9 1 9 16 13 1 10 9 1 10 9 13 1 10 9 0 1 10 9 15 13 10 0 9 2
39 10 9 1 10 11 2 11 11 2 13 16 10 11 11 13 1 10 11 7 16 4 13 1 10 9 0 2 4 13 15 3 1 10 9 1 10 9 0 2
13 15 13 1 10 9 1 11 1 10 9 1 11 2
17 16 15 13 9 1 10 9 2 11 15 13 2 7 13 10 9 2
19 3 3 13 15 1 10 3 0 9 0 2 7 3 10 0 9 1 13 2
22 15 13 1 10 0 9 1 9 3 0 1 11 7 10 9 0 1 10 11 11 11 2
5 13 1 9 0 2
29 16 10 9 3 13 0 2 10 9 2 9 2 13 10 15 16 2 13 2 1 10 9 7 13 1 13 10 9 2
9 15 13 7 4 1 13 1 12 2
24 13 10 9 0 1 10 9 1 11 2 3 3 1 11 16 13 10 9 1 9 7 15 13 2
28 10 9 1 0 9 1 10 9 13 13 1 10 9 1 11 2 1 3 15 4 13 1 10 3 12 1 15 2
30 16 10 9 1 10 9 16 13 1 10 9 7 1 10 9 0 7 0 2 3 4 13 7 10 3 0 9 1 9 2
38 1 3 13 10 3 0 9 0 1 10 11 0 1 10 9 0 2 1 10 11 1 10 11 7 3 9 1 10 11 11 1 10 11 11 7 11 11 2
13 10 9 1 9 13 1 12 13 2 2 9 8 2
31 10 9 13 10 9 0 1 10 9 3 0 1 10 9 0 2 2 3 13 2 0 1 13 7 1 15 15 13 2 9 2
20 11 11 13 10 9 1 9 1 10 9 1 10 9 1 10 9 1 10 11 2
30 1 10 9 1 10 9 1 10 9 0 13 1 11 7 1 13 12 9 13 1 10 11 11 3 13 10 9 1 12 2
9 13 10 9 0 1 13 10 9 2
15 11 11 11 13 10 9 0 13 10 12 1 11 1 12 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
14 2 10 9 7 10 9 13 10 9 1 10 9 0 2
23 10 9 13 10 9 1 13 10 9 1 10 15 4 0 2 13 13 2 13 1 9 0 2
22 1 10 9 13 1 9 9 0 7 13 10 9 1 13 9 0 1 10 9 1 11 2
26 10 9 4 13 15 1 0 9 0 1 16 10 13 10 9 15 3 0 1 4 13 1 9 0 0 2
24 10 9 0 4 13 0 1 10 9 0 2 1 15 15 10 9 0 13 1 10 9 1 9 2
54 1 10 9 1 10 9 4 13 2 13 3 13 10 9 2 7 15 13 10 9 1 10 9 0 1 10 9 2 16 13 1 13 15 2 0 2 1 9 2 9 7 9 1 9 13 1 10 9 0 2 0 7 0 2
9 10 9 4 13 15 1 10 9 2
20 1 0 9 10 9 1 10 9 2 11 11 2 13 3 16 10 9 13 0 2
16 10 9 1 10 9 13 1 10 9 1 10 15 2 9 2 2
22 11 13 11 1 2 10 0 9 1 0 9 2 7 15 13 0 1 10 9 7 9 2
28 13 3 0 7 0 2 16 13 10 9 13 13 1 15 1 10 9 2 15 13 10 9 15 0 1 10 9 2
27 15 13 1 10 9 12 13 1 11 13 1 11 11 10 12 1 11 1 12 7 13 1 10 9 11 11 2
19 1 10 9 2 13 10 9 1 9 0 1 9 1 11 0 1 11 11 2
26 15 13 1 9 7 15 9 16 4 13 13 16 15 13 16 13 10 9 1 10 9 3 4 13 15 2
16 10 9 3 13 0 2 7 10 9 7 10 9 15 15 13 2
13 15 1 10 9 16 13 1 10 9 13 9 0 2
29 11 12 13 0 9 1 11 1 10 9 11 2 7 4 7 13 15 1 12 1 4 13 9 0 1 11 7 11 2
31 13 1 10 9 0 1 10 9 2 15 13 1 13 9 0 1 10 9 16 15 13 2 7 3 1 9 1 9 1 9 2
28 11 11 2 7 13 10 9 11 2 11 2 11 2 13 10 0 9 0 13 10 12 1 11 1 12 1 11 2
44 3 15 2 13 10 9 1 9 10 0 9 1 11 1 11 7 11 9 16 13 1 0 9 2 7 13 10 9 1 11 1 11 1 3 13 3 1 10 0 9 1 10 12 2
22 10 9 1 10 0 13 1 12 5 8 2 7 10 9 1 10 9 13 1 12 5 8
61 1 9 1 10 9 0 2 10 9 13 0 1 10 9 1 10 9 2 10 9 3 13 10 12 5 8 7 10 0 3 13 1 3 1 12 5 8 10 9 3 0 13 1 11 13 1 12 5 8 2 1 11 11 2 10 12 1 11 1 12 2
30 11 11 11 2 11 2 12 2 2 13 10 9 0 2 9 0 7 9 2 13 1 10 9 1 10 9 1 10 9 2
67 7 16 1 10 9 4 13 1 13 1 10 9 1 10 0 9 1 10 11 11 1 11 2 1 10 9 4 13 15 3 3 1 13 10 9 3 3 13 1 10 11 11 1 11 7 1 9 1 15 13 1 10 9 7 9 10 0 0 9 2 11 11 11 11 11 11 2
6 13 0 1 10 9 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
19 7 1 9 1 10 9 2 10 9 4 13 10 12 5 2 13 10 9 2
41 10 9 7 10 9 4 13 1 10 9 1 10 9 2 4 13 1 10 9 0 1 10 9 1 11 0 1 10 9 1 11 10 12 1 11 2 16 3 15 13 2
28 1 12 2 11 13 1 10 9 1 11 1 13 16 15 13 10 9 0 1 11 11 7 13 0 1 10 9 2
26 1 10 9 1 12 13 1 10 12 9 0 1 9 1 11 2 3 13 1 13 15 1 11 7 11 2
30 3 3 2 10 9 1 11 11 13 10 9 0 0 2 16 10 9 0 1 10 9 15 13 1 10 9 1 9 0 2
11 15 15 13 2 7 15 13 1 0 9 2
38 10 11 11 13 15 15 13 10 9 1 10 1 2 11 11 11 2 1 9 1 15 1 10 9 1 11 1 10 9 11 9 1 11 1 11 11 11 2
18 10 9 13 11 11 11 2 0 9 1 9 2 9 2 9 7 9 2
23 10 11 1 11 13 10 9 1 9 1 12 8 8 12 8 2 12 5 8 12 5 2 2
45 3 7 3 10 9 13 9 0 0 2 15 13 1 9 3 1 4 13 1 9 7 1 9 0 15 4 4 13 1 10 9 1 9 2 1 13 9 2 9 1 9 7 9 0 2
29 10 9 1 9 13 3 10 9 1 16 10 10 9 13 1 10 0 9 2 7 13 9 0 1 13 1 10 9 2
19 1 9 1 10 11 1 11 1 12 10 9 1 10 9 13 10 12 9 2
37 10 9 3 0 2 15 3 10 12 5 9 2 7 4 1 13 16 9 0 7 10 10 9 0 2 15 1 10 0 9 8 15 13 7 15 13 2
26 10 9 4 13 10 0 9 2 1 12 2 1 12 9 1 10 9 1 15 1 10 9 1 10 9 2
12 10 9 3 4 4 1 13 15 2 2 13 2
7 1 15 15 13 12 9 2
25 9 0 7 0 1 10 9 0 1 10 9 0 2 10 9 0 15 13 1 10 9 1 10 9 2
30 1 9 1 10 9 12 13 0 9 1 9 0 1 10 9 2 2 9 11 2 11 2 9 11 7 11 2 11 2 2
17 10 9 15 13 1 10 9 1 10 9 0 1 15 1 10 9 2
34 10 9 0 1 10 13 10 9 1 9 0 7 13 10 9 7 9 2 1 15 15 1 10 9 2 13 10 9 1 10 9 3 0 2
25 10 9 0 13 15 15 13 11 11 1 12 1 10 9 1 10 9 1 10 11 11 12 1 11 2
54 9 2 11 10 11 11 13 1 10 0 9 10 9 1 10 9 1 13 1 10 9 12 9 1 10 9 13 1 10 9 1 10 9 1 10 9 13 1 16 10 9 1 10 9 7 10 9 3 15 13 1 13 9 2
26 11 15 13 16 15 13 1 10 9 1 10 9 1 11 1 10 9 9 7 1 9 15 13 1 13 2
21 11 3 13 0 9 2 1 9 1 16 10 0 9 13 3 1 9 1 13 15 2
46 1 12 11 11 13 10 0 9 1 9 1 10 9 11 2 1 10 9 15 13 10 0 9 2 2 10 9 4 13 1 10 0 9 1 10 9 1 9 1 9 1 9 1 10 9 12
34 11 11 4 13 1 10 9 11 1 12 1 13 11 11 2 13 15 1 9 1 11 11 2 3 1 4 13 1 10 9 0 11 11 2
8 15 13 0 2 0 2 0 2
26 2 1 9 15 13 10 15 0 2 7 3 13 1 13 15 1 10 9 2 2 13 1 10 9 9 2
60 2 10 9 13 10 11 10 9 1 11 11 2 15 13 10 9 1 10 11 1 10 9 7 9 10 9 13 10 9 0 1 10 8 8 2 8 2 8 8 8 2 7 10 2 8 1 10 9 2 2 16 13 10 9 1 8 9 1 13 2
21 10 9 0 13 1 10 9 13 10 9 2 7 10 9 13 1 9 1 10 9 2
16 1 10 9 0 13 10 9 2 10 9 7 9 1 10 9 2
46 10 11 1 10 11 1 11 1 11 2 1 9 12 1 11 1 12 2 13 10 9 1 16 10 11 11 1 10 11 4 13 9 1 10 11 11 1 10 11 7 1 10 9 1 11 2
8 11 15 13 0 1 10 9 2
70 1 10 9 2 10 9 1 10 9 15 13 1 9 10 9 1 9 1 9 1 11 11 2 11 11 11 2 11 11 7 11 11 2 3 1 10 0 9 0 1 10 15 1 10 9 16 13 10 9 1 10 9 2 7 16 10 9 0 13 1 9 1 10 9 10 9 13 10 9 2
15 13 10 0 9 1 9 7 9 1 9 1 3 0 9 2
11 10 9 1 11 15 13 13 1 10 9 2
14 1 15 13 1 0 9 10 4 13 15 1 10 9 2
14 1 12 7 12 2 13 1 10 9 0 1 11 11 2
26 16 3 15 13 2 15 13 1 10 0 9 1 10 13 7 10 9 13 1 10 9 0 1 10 9 2
33 10 9 12 11 11 2 1 9 2 11 12 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 1 10 11 2
13 10 9 3 0 13 1 9 0 1 10 9 0 2
29 1 10 9 2 3 2 15 13 10 9 2 11 11 2 1 10 9 0 16 13 10 9 1 10 9 1 10 9 2
36 10 9 15 13 3 1 9 1 10 9 13 1 11 1 11 7 11 11 2 13 1 11 11 2 11 11 2 11 11 7 11 11 2 1 15 2
7 1 0 2 13 0 9 2
10 15 13 1 10 11 11 1 10 11 2
27 1 12 2 11 13 0 1 11 11 7 11 11 10 9 11 11 11 2 9 1 9 7 3 3 9 2 2
15 13 13 1 10 9 3 7 10 9 1 9 13 3 0 2
49 10 9 2 11 15 13 1 10 9 2 7 13 16 13 16 4 4 13 10 0 9 2 9 2 16 3 1 4 4 13 10 9 2 13 10 9 0 16 15 13 10 9 1 13 1 9 1 9 2
27 3 2 3 1 13 1 10 9 1 10 9 1 9 2 15 1 10 9 1 15 2 13 1 10 11 11 2
37 3 13 16 1 10 9 15 13 1 10 9 1 10 9 0 13 1 9 0 2 3 7 1 10 9 7 9 1 10 9 1 9 0 2 8 2 2
47 13 1 10 9 1 10 0 9 1 10 9 3 0 13 1 11 13 1 10 9 7 3 1 10 11 2 10 9 13 10 9 0 0 13 1 10 9 1 10 9 1 11 11 1 11 11 2
29 10 0 9 2 13 3 2 7 10 9 3 2 4 13 10 9 1 13 16 13 0 3 7 13 10 9 1 9 2
28 3 2 10 8 11 2 13 16 10 9 8 2 8 7 8 2 13 2 1 10 9 1 10 9 13 1 9 2
8 13 10 9 1 12 9 8 2
57 2 10 9 1 10 9 2 15 1 10 0 2 2 10 9 1 10 9 2 10 1 10 9 2 2 10 9 1 10 9 16 15 13 2 10 9 1 10 9 1 11 11 16 13 10 9 1 10 9 16 3 13 1 15 9 13 2
34 10 9 4 4 13 3 1 9 0 2 16 4 13 12 2 13 1 10 12 1 9 1 9 2 10 0 9 7 15 13 1 10 9 2
21 1 0 2 15 13 0 1 10 9 13 1 10 9 1 9 2 16 13 1 13 2
21 13 0 16 15 15 13 1 7 10 9 16 13 1 9 9 3 13 1 10 9 2
76 1 10 9 4 13 9 0 1 2 11 10 11 11 1 11 2 2 2 11 11 11 15 11 11 2 2 10 3 0 1 10 9 2 2 2 11 2 2 7 3 9 1 9 3 0 2 13 15 2 11 2 2 10 0 2 11 11 15 2 7 10 0 2 11 11 2 1 10 15 15 13 10 9 1 11 2
13 10 11 11 13 10 9 1 10 9 1 10 9 2
41 10 9 3 1 10 9 4 13 9 1 10 9 1 10 9 2 10 9 2 9 7 9 16 13 0 2 7 10 9 1 9 7 9 0 16 13 9 1 10 9 2
38 7 3 13 1 10 9 12 16 13 10 0 9 1 9 1 10 13 1 10 9 11 11 3 13 1 11 11 2 13 1 13 1 11 1 10 9 8 2
14 3 10 0 9 13 13 15 1 10 9 1 10 9 2
13 4 13 15 1 10 9 3 0 1 10 9 0 2
12 13 1 12 7 12 9 1 9 2 3 0 2
20 10 11 11 13 10 9 0 16 13 13 10 9 0 1 10 9 0 7 0 2
24 15 13 1 10 9 1 10 9 1 9 1 10 9 2 7 1 13 2 15 4 13 10 9 2
16 10 0 9 15 13 2 11 11 2 2 11 11 2 12 2 2
18 10 9 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
52 1 9 1 10 0 9 1 10 9 7 10 9 13 3 10 9 1 10 9 13 1 10 9 0 1 10 9 2 10 1 10 9 2 10 1 10 9 1 11 7 10 9 1 10 11 13 1 10 9 1 11 2
4 13 1 13 2
44 13 0 9 1 10 9 1 10 9 0 2 7 15 1 10 3 0 7 13 1 0 9 1 10 9 13 10 9 1 12 9 1 11 1 11 16 13 10 9 1 11 2 11 2
29 1 10 9 1 10 9 2 10 0 9 4 13 1 13 10 9 0 1 15 7 13 1 10 0 9 16 13 11 2
33 3 1 10 9 0 1 10 9 1 9 1 10 11 11 1 11 12 1 11 2 10 9 15 13 1 13 9 1 10 9 1 12 2
40 1 10 9 2 10 9 4 13 15 1 10 3 9 1 10 9 1 9 2 3 1 16 13 10 0 9 0 1 13 10 9 1 10 9 2 9 2 9 2 2
10 13 9 0 1 11 11 7 11 12 2
73 1 10 9 1 9 8 2 0 2 11 2 2 15 4 1 13 7 1 13 10 9 0 16 4 8 10 9 1 10 9 1 10 9 2 3 1 12 1 10 9 0 2 1 3 13 15 1 13 1 10 9 12 1 3 13 1 10 9 1 11 11 11 2 3 13 1 2 10 9 1 9 2 2
22 1 10 9 2 10 9 3 13 1 10 9 1 9 10 12 9 2 13 11 11 3 2
8 10 11 1 11 3 13 3 2
21 10 0 9 13 1 11 1 12 7 10 9 15 4 13 10 12 1 11 1 12 2
21 10 9 0 0 7 9 0 2 11 11 2 13 10 9 1 9 0 1 10 9 11
10 3 13 10 11 12 7 10 11 12 2
40 3 13 10 9 16 13 10 9 0 2 7 10 11 11 2 11 11 2 7 10 11 1 10 11 11 2 11 11 2 13 10 9 0 1 10 9 1 10 9 2
10 3 11 13 10 9 1 11 1 12 2
16 15 13 3 1 10 9 9 2 9 7 0 1 10 9 0 2
18 1 9 0 2 10 9 1 11 4 13 1 12 9 1 9 7 9 2
35 1 9 2 11 13 10 12 1 11 1 12 2 1 12 10 9 2 1 10 9 1 9 13 1 10 9 1 11 1 10 9 0 11 11 2
22 10 9 4 13 1 13 10 3 0 9 1 10 11 2 10 9 0 13 10 12 9 2
10 10 9 13 0 7 13 10 15 9 2
52 13 3 4 13 7 3 13 2 1 15 3 15 13 9 1 15 16 4 13 3 3 2 15 16 3 15 13 13 16 15 4 13 3 1 10 9 1 7 15 13 10 9 1 10 9 7 1 10 9 16 13 2
19 1 11 2 11 11 13 10 0 9 1 9 3 1 9 1 10 0 9 2
18 13 9 1 9 9 2 9 7 9 2 9 2 9 7 15 1 9 2
74 10 9 1 10 9 15 13 1 10 9 1 16 10 9 4 13 1 10 9 1 9 7 10 9 3 13 0 9 1 10 9 2 9 0 2 4 13 1 10 9 1 10 9 2 13 9 0 7 10 9 3 0 1 10 9 1 9 1 9 16 13 0 9 1 10 0 9 1 10 9 16 15 13 2
44 10 9 0 16 13 10 9 0 13 9 0 1 9 0 3 0 2 9 0 2 9 0 2 0 7 0 2 9 1 9 2 9 2 9 1 10 9 0 7 9 1 10 9 2
10 11 11 13 1 10 9 1 11 12 2
22 1 3 1 10 9 1 9 2 11 13 3 1 11 1 12 9 1 9 1 9 13 2
11 10 0 9 13 1 10 11 10 8 11 2
20 1 12 2 13 10 9 1 11 16 13 1 10 9 1 13 9 1 10 9 2
9 1 10 9 12 13 1 12 9 2
20 13 0 16 10 9 13 3 1 12 9 1 13 10 9 1 9 1 10 9 2
9 10 9 13 10 9 7 10 9 2
45 10 9 1 10 9 15 13 1 10 9 1 10 11 1 10 11 11 2 9 16 3 15 13 1 13 12 9 7 16 3 4 13 1 11 1 9 1 9 1 9 1 10 10 9 2
31 10 9 0 2 11 4 13 1 0 9 1 10 11 1 10 9 1 9 1 12 1 10 11 1 11 1 10 11 1 11 2
26 1 10 9 0 2 11 13 1 10 9 1 13 16 10 9 1 9 15 4 13 7 13 1 10 9 2
23 13 9 7 9 7 15 13 1 9 1 9 2 1 9 1 9 15 13 1 9 0 2 2
34 10 9 1 10 9 1 11 2 9 1 10 12 5 9 0 2 3 15 13 1 9 1 11 1 12 1 10 9 1 10 9 1 9 2
18 10 9 11 13 10 9 1 9 0 13 9 0 7 0 1 10 9 2
25 10 9 1 11 15 13 1 0 9 10 12 1 11 1 12 1 11 2 3 15 13 1 10 9 2
26 10 9 15 13 3 1 10 9 2 1 11 0 15 13 2 11 2 1 10 9 13 7 13 1 9 2
39 13 1 11 16 13 1 10 11 1 11 2 7 15 13 10 9 7 10 9 13 3 1 16 11 13 10 9 1 13 15 2 13 1 11 1 11 1 12 2
33 10 9 0 2 3 13 1 10 9 1 9 11 2 13 10 9 1 9 16 13 1 9 1 10 9 1 9 2 13 3 1 9 2
22 13 3 0 13 1 10 9 2 13 9 0 7 13 9 16 13 1 10 9 7 9 2
37 9 1 10 11 11 1 11 1 11 0 2 11 2 2 16 13 9 1 10 11 11 1 11 11 2 11 2 2 1 10 15 13 9 1 12 9 2
16 10 9 13 1 10 9 0 1 10 0 9 7 13 3 0 2
14 1 10 9 0 15 13 9 1 9 2 11 11 2 2
33 1 10 9 1 10 12 10 9 1 9 0 1 10 9 1 10 9 13 1 12 9 7 10 9 0 1 10 9 13 1 12 9 2
8 11 13 3 0 1 10 9 2
51 13 1 10 9 3 1 11 13 10 9 0 1 10 9 7 9 1 11 1 12 9 2 10 9 2 10 9 0 1 10 9 0 7 1 10 9 1 13 15 10 9 13 1 10 9 2 3 1 10 9 2
7 3 4 13 10 9 0 2
27 15 13 2 1 15 2 1 10 9 1 10 9 0 1 10 9 7 10 9 1 10 9 0 1 10 9 2
19 13 2 9 1 10 9 2 2 9 9 2 1 10 11 1 10 11 11 2
8 13 10 10 9 1 9 0 2
23 3 3 2 11 13 10 9 2 13 1 11 2 1 10 0 9 2 16 3 15 13 11 2
5 7 3 13 0 2
22 11 11 11 13 10 0 9 9 1 10 9 0 1 11 11 11 7 4 13 1 12 2
45 1 15 13 10 9 1 9 1 9 0 16 13 10 9 0 3 0 7 0 1 10 9 0 1 3 1 10 9 2 13 1 9 0 2 10 15 13 1 9 7 10 9 7 9 2
31 1 10 9 1 9 2 10 9 0 13 16 11 13 9 1 10 9 7 13 10 9 1 9 1 10 9 16 13 3 3 2
57 16 10 0 9 1 10 9 15 13 16 0 9 15 13 1 10 9 1 11 2 4 13 15 1 9 1 0 9 16 3 13 0 9 15 13 10 9 2 7 13 3 0 1 13 1 9 16 10 9 4 13 1 10 9 1 11 2
23 3 10 9 3 0 7 15 15 13 16 1 10 9 1 11 13 0 10 9 1 10 11 2
12 10 11 4 13 1 0 9 13 1 10 11 2
30 10 9 7 10 9 0 1 0 9 13 10 9 1 9 7 1 9 2 9 0 1 10 9 1 10 9 1 10 9 2
53 1 11 1 12 15 13 16 10 0 9 0 1 9 0 1 0 9 2 10 11 11 12 4 13 1 4 13 1 9 0 1 10 9 2 1 9 1 16 10 9 3 13 15 3 0 16 10 9 11 11 2 12 2
84 10 9 0 16 13 1 10 9 1 10 9 3 13 15 7 10 0 11 1 11 2 13 1 10 9 1 9 0 7 0 2 1 10 15 15 13 0 10 11 11 1 11 1 11 2 10 11 11 1 10 11 1 11 2 11 11 2 8 2 10 11 8 1 11 11 1 11 2 10 9 1 10 11 11 1 10 11 1 10 11 2 8 2 8
46 1 15 9 2 12 7 12 1 9 13 1 10 9 1 11 1 2 9 1 9 2 1 10 9 2 1 9 1 10 9 1 10 9 1 10 9 1 10 11 2 3 13 1 10 9 2
17 10 9 15 13 10 9 2 13 12 9 7 13 10 9 16 13 2
17 16 9 1 9 13 16 13 10 9 2 10 9 13 13 10 9 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
19 10 9 13 11 11 2 0 1 11 2 7 11 11 11 2 0 1 11 2
9 13 9 1 10 9 1 9 13 2
16 3 3 1 10 9 1 10 9 1 10 9 2 11 4 13 2
32 10 9 1 13 9 0 1 9 3 0 15 13 1 9 1 10 9 0 12 2 12 1 9 1 10 9 1 12 1 12 9 2
25 13 9 16 13 1 13 10 9 1 10 9 2 13 1 10 9 2 13 1 9 3 3 1 9 2
24 1 9 2 1 10 9 2 1 11 2 11 7 11 2 3 1 10 9 1 10 9 13 0 2
8 3 13 1 10 9 1 11 2
29 10 9 0 3 0 13 11 2 12 2 2 11 2 12 2 2 11 2 12 2 7 11 11 7 11 2 12 2 2
63 1 10 12 9 2 10 9 1 11 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
47 10 9 2 13 1 9 1 10 9 13 1 10 9 1 10 9 2 10 11 1 11 2 2 13 3 1 10 9 1 11 11 2 9 1 9 7 10 9 0 1 10 9 1 10 9 0 2
29 11 12 13 10 9 3 0 1 3 1 10 9 2 3 16 13 0 1 11 12 1 9 0 2 7 3 13 0 2
31 10 9 0 1 10 9 2 1 10 3 1 10 9 0 1 1 13 1 15 2 1 10 9 0 2 10 9 0 7 0 2
30 10 9 1 15 13 1 10 9 1 10 9 1 9 1 9 2 9 1 10 15 13 2 1 10 9 1 13 1 3 2
13 1 10 9 2 13 1 10 9 1 10 9 0 2
17 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 11 2
24 13 3 1 10 9 2 11 11 2 2 13 1 12 9 2 9 2 9 1 9 7 9 0 2
25 1 10 9 2 10 0 9 1 11 12 1 10 9 1 10 9 13 10 9 1 10 9 1 9 2
20 10 9 1 10 9 11 13 1 10 9 10 9 1 10 9 1 9 7 9 2
35 10 9 13 1 10 9 10 11 1 10 9 1 11 1 10 9 16 13 2 13 10 9 7 10 9 2 13 1 11 7 1 10 9 2 2
20 10 9 1 10 9 15 13 1 0 9 2 9 7 2 7 9 1 9 2 2
11 1 3 4 13 10 15 13 1 10 9 2
17 10 9 0 2 9 1 16 15 13 0 2 3 13 15 1 0 2
24 10 10 9 1 10 9 13 11 11 2 11 11 2 11 11 7 10 9 1 11 11 1 11 2
45 10 0 9 1 13 10 9 1 10 9 2 16 10 9 13 0 1 13 2 13 1 10 9 10 9 1 11 11 1 10 11 1 11 1 9 1 11 11 2 16 13 1 10 9 2
20 1 13 10 9 11 13 10 9 13 1 9 1 10 9 1 9 2 11 2 2
26 1 10 9 13 10 9 2 16 13 10 11 11 7 10 9 1 10 9 1 10 9 1 9 1 9 2
20 11 11 13 10 9 1 9 1 10 9 1 10 11 1 10 9 1 10 9 2
25 11 13 1 10 9 0 1 9 1 11 2 15 16 15 13 13 1 10 9 1 11 1 15 13 2
19 13 0 1 11 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2
43 1 9 1 10 9 1 10 11 2 10 11 7 10 9 1 10 9 1 10 9 1 10 11 2 1 10 9 1 10 9 2 10 11 2 10 9 2 11 2 7 10 9 2
10 1 10 9 15 13 1 9 1 0 2
35 10 9 1 9 7 9 15 13 1 10 15 0 2 10 1 10 9 8 2 0 7 9 15 9 4 1 13 1 10 9 1 10 9 0 2
27 10 9 13 13 10 9 0 1 9 1 10 9 2 1 10 9 1 10 9 16 15 13 1 10 9 0 2
19 15 13 1 9 1 15 1 10 9 0 1 10 9 1 10 9 1 9 2
18 11 13 1 10 9 13 2 1 10 9 1 10 9 7 1 10 9 2
24 10 9 1 9 13 1 10 9 1 10 9 1 10 9 2 10 9 7 10 9 16 15 13 2
37 10 9 16 13 1 10 0 9 1 10 11 16 10 9 11 11 13 1 11 13 10 9 10 9 2 1 10 9 1 11 2 1 12 9 1 9 2
11 13 1 9 3 1 9 1 10 9 0 2
41 1 10 9 1 3 10 9 2 1 10 0 9 2 9 1 9 1 10 9 1 9 7 10 9 1 0 9 1 9 11 2 13 0 1 10 0 9 0 0 0 2
45 1 10 9 4 13 0 9 1 10 9 2 10 9 2 10 11 7 10 9 2 7 3 15 3 0 1 10 9 2 10 11 1 9 2 10 11 2 10 9 7 10 10 9 0 2
73 13 0 1 10 9 16 13 2 7 15 1 10 9 0 13 16 15 1 15 2 13 10 9 15 16 15 13 13 3 0 2 7 3 15 13 10 9 16 4 13 16 13 15 1 3 2 13 3 0 2 15 15 15 13 1 15 2 1 15 13 15 1 10 0 8 8 8 16 4 13 1 11 2
24 10 9 4 13 15 0 2 3 1 2 9 0 2 2 2 7 3 13 0 1 10 9 0 2
12 3 4 3 13 1 10 9 1 10 9 12 2
34 10 9 1 11 3 13 10 9 1 10 10 9 16 15 13 1 10 9 0 1 10 9 13 1 10 9 0 1 9 13 1 10 9 2
8 1 10 9 13 10 9 11 2
29 11 11 11 11 13 10 9 1 11 11 13 1 10 0 9 0 1 10 9 3 2 7 3 3 0 16 10 9 2
33 13 1 10 9 0 1 11 2 15 13 1 10 9 1 10 9 1 12 1 13 10 9 11 1 10 12 2 13 1 10 9 11 2
17 3 13 9 0 2 3 13 10 9 1 10 9 0 1 10 9 2
36 1 9 1 10 9 1 12 13 1 10 9 1 11 2 10 9 1 9 13 1 12 12 9 2 12 5 2 7 12 12 9 2 12 5 2 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
21 1 10 11 2 11 11 12 13 10 9 7 10 9 1 9 1 9 1 11 12 2
12 13 1 10 11 2 11 1 11 11 7 11 2
69 11 11 1 11 2 13 3 11 7 1 12 1 11 2 2 11 11 1 11 1 9 2 2 13 10 9 0 13 1 11 2 11 2 1 12 1 9 1 11 7 3 3 1 9 2 0 2 1 10 11 11 2 1 11 11 1 10 11 11 2 7 11 11 7 1 10 11 0 2
25 13 1 9 1 10 9 7 15 13 2 10 9 13 0 2 3 7 13 10 9 1 9 7 0 2
34 10 9 2 16 13 10 9 1 10 9 0 2 15 13 1 3 13 1 10 9 2 16 15 13 1 13 7 13 1 9 1 10 9 2
43 1 13 1 10 9 2 7 13 10 9 1 10 9 7 16 10 9 3 13 1 10 9 2 7 13 16 15 13 15 16 4 13 10 9 2 15 13 1 10 9 1 11 2
8 13 10 9 1 9 3 0 2
27 13 10 15 16 13 1 10 9 1 9 2 3 1 9 13 10 9 1 10 9 16 13 1 10 9 13 2
7 13 10 9 1 11 11 2
38 11 11 2 13 10 12 1 11 1 12 1 11 2 13 10 12 1 11 1 12 1 11 2 4 13 1 9 7 0 9 1 10 9 0 1 9 11 2
15 15 13 9 7 9 1 0 9 1 13 16 3 4 13 2
21 10 9 0 15 13 1 9 0 1 10 0 9 1 10 11 2 1 9 0 9 2
11 10 9 3 0 13 15 1 11 11 11 2
11 11 13 10 0 9 1 10 9 0 0 2
53 1 11 1 10 11 2 16 13 10 9 0 2 15 15 13 10 9 1 10 9 0 16 13 1 10 9 1 11 11 11 1 11 1 9 1 10 11 1 13 15 9 1 10 9 2 7 3 1 9 7 1 11 2
14 10 9 13 10 9 1 10 9 4 13 1 15 0 2
11 10 9 13 10 9 0 1 0 9 0 2
28 13 1 10 11 1 11 1 12 2 16 15 13 3 7 15 13 1 11 1 13 1 10 9 0 1 10 9 2
31 13 3 1 12 9 13 10 9 16 4 7 13 1 10 9 1 11 7 3 3 3 13 2 7 16 7 3 13 10 9 2
21 10 11 15 4 13 1 10 9 1 10 9 11 2 9 0 1 10 0 11 11 2
18 10 11 13 10 9 0 1 12 9 2 10 9 4 4 13 1 11 2
19 10 9 1 9 1 11 2 11 13 10 9 1 9 0 1 10 9 1 9
40 1 10 9 2 10 9 13 1 10 9 1 9 2 13 1 10 9 0 2 2 13 1 10 9 1 10 9 9 2 1 10 9 1 8 2 8 1 10 9 2
40 11 2 13 1 3 4 4 13 1 11 2 13 13 10 9 1 9 2 15 16 13 1 11 7 11 2 15 13 13 15 1 4 13 1 9 1 10 0 11 2
37 10 9 0 1 11 11 13 15 1 10 12 9 1 10 9 1 10 11 2 13 1 10 9 1 10 11 2 1 10 9 10 9 0 1 10 11 2
6 2 3 13 1 9 2
29 1 10 9 13 10 9 0 1 9 0 2 3 15 15 4 13 1 10 9 1 10 9 7 10 9 1 9 0 2
22 15 13 1 10 11 1 11 1 12 9 1 11 1 10 11 2 12 7 11 2 12 2
33 10 9 4 13 1 9 2 9 7 9 1 10 9 2 7 15 13 1 10 9 1 11 1 12 2 16 4 13 1 10 9 0 2
17 1 10 9 2 15 13 1 10 0 9 8 2 7 1 9 0 2
8 10 9 7 10 9 3 13 2
13 10 9 1 10 9 13 3 1 15 1 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
34 1 10 9 13 1 11 2 3 13 9 1 10 9 11 2 13 3 10 9 1 10 9 1 10 9 1 9 7 9 2 1 15 2 2
40 1 0 7 15 1 10 9 1 10 11 15 13 15 1 10 9 1 9 2 7 10 0 9 1 10 9 13 1 10 9 1 10 11 12 2 10 12 1 11 2
30 10 9 0 13 10 9 1 10 9 0 16 13 16 10 9 4 13 1 9 0 2 7 13 10 9 1 9 3 0 2
33 10 10 9 1 11 3 13 0 1 10 11 11 1 10 9 1 9 1 9 1 11 2 10 15 4 13 10 12 1 11 1 12 2
30 3 2 10 9 11 12 13 10 9 10 12 1 11 1 12 2 13 15 1 10 9 10 12 1 11 1 10 0 9 2
23 1 12 11 7 11 13 1 9 16 13 10 9 13 1 11 1 9 1 10 11 11 11 2
13 10 9 13 15 1 15 16 1 9 13 10 9 2
30 10 9 13 13 10 9 1 9 15 16 13 10 9 1 0 9 1 9 7 16 3 13 1 10 0 9 1 10 9 2
12 13 10 9 0 2 0 7 1 10 9 0 2
14 10 9 13 1 10 9 0 1 10 13 13 1 12 8
31 10 11 11 13 15 1 10 12 0 9 15 4 4 13 1 10 9 1 10 9 3 1 10 11 11 7 1 10 11 11 2
5 15 13 1 11 2
15 13 10 9 7 10 9 0 1 10 0 9 0 1 11 2
30 13 9 1 9 10 9 0 7 0 16 13 1 10 9 1 9 0 7 9 0 16 13 1 10 9 7 9 1 9 2
8 2 9 1 9 1 10 9 11
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
28 10 9 1 10 9 13 10 9 0 2 1 9 0 9 3 15 15 13 1 0 9 3 1 10 9 1 9 2
32 11 13 1 10 9 2 2 10 9 8 13 9 0 2 3 0 2 16 13 10 9 0 2 1 15 10 9 1 10 9 0 2
25 3 1 10 9 13 10 9 0 2 10 15 4 13 1 10 9 1 10 9 3 15 13 10 9 2
14 10 9 1 9 3 13 1 10 0 9 1 10 9 2
27 15 13 9 0 1 13 9 0 2 0 7 0 1 10 9 2 1 9 0 1 10 0 9 1 10 9 2
21 13 12 9 2 13 12 7 13 12 2 13 12 9 7 13 12 2 13 12 9 2
56 11 4 13 1 9 1 10 9 16 13 13 3 3 10 9 1 10 9 2 11 1 10 11 2 11 1 10 11 2 11 11 2 11 2 11 2 11 2 1 10 9 1 10 9 2 1 10 9 1 9 2 0 2 1 11 2
27 10 9 0 2 1 9 2 13 12 9 1 0 2 13 1 9 1 15 9 1 10 9 0 1 10 9 2
59 10 9 0 13 15 1 10 9 0 9 3 0 7 0 2 15 13 1 9 1 9 2 13 10 9 1 0 9 0 1 10 9 2 10 16 15 13 3 0 2 3 15 13 1 10 9 1 9 0 2 9 7 9 1 9 1 9 0 2
13 4 3 13 1 15 1 10 9 0 1 10 9 2
21 10 9 13 12 9 2 7 10 9 13 10 9 1 9 10 12 1 11 1 12 2
36 1 10 9 12 13 1 13 10 9 0 11 10 9 1 10 11 2 9 2 7 13 10 9 0 1 9 1 9 16 13 10 11 1 10 11 2
4 10 0 9 2
9 13 13 1 10 9 2 7 13 2
14 10 9 0 13 16 1 10 9 13 3 1 12 9 2
46 10 12 1 11 1 12 10 9 4 13 1 10 9 0 1 9 8 2 5 2 3 1 10 0 9 1 9 2 1 10 9 1 10 9 1 10 9 2 15 15 13 3 1 10 9 2
25 10 9 0 16 13 10 9 13 10 9 0 7 2 1 10 9 0 2 13 3 1 12 9 0 2
18 10 9 0 1 10 9 13 10 12 5 1 10 9 0 1 10 9 2
10 11 11 4 4 13 1 0 9 0 2
50 9 16 13 9 1 10 11 11 1 10 11 2 13 1 10 9 11 2 1 10 9 0 1 10 11 2 9 3 15 4 1 13 10 9 0 1 9 2 13 1 10 9 10 0 9 7 10 0 9 2
36 13 15 2 9 1 11 11 2 13 10 9 1 9 7 9 0 13 1 11 2 16 13 1 10 9 13 7 13 10 9 1 9 1 10 11 2
11 4 13 1 10 9 0 1 10 9 12 2
24 3 2 13 9 1 9 2 9 2 9 2 9 1 9 2 9 1 9 1 9 7 8 0 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
13 10 9 13 10 9 3 0 1 10 9 1 11 2
21 10 13 10 0 7 0 9 2 7 15 13 1 10 9 1 10 12 9 1 9 2
47 10 11 4 13 1 13 3 1 5 12 9 1 10 9 0 1 10 9 7 4 13 3 1 5 12 9 1 9 1 9 15 4 4 13 1 13 10 9 0 2 9 7 10 9 1 9 2
9 3 13 11 7 10 11 1 11 2
24 13 15 9 2 3 15 13 15 13 15 16 13 1 10 9 1 10 9 0 1 11 7 9 2
19 11 13 10 0 9 0 7 9 0 1 9 2 7 1 3 15 13 9 2
49 10 0 9 2 11 11 11 11 11 11 2 4 13 7 10 9 1 11 13 1 12 2 13 15 1 10 0 11 11 1 11 1 10 11 2 1 15 15 10 9 13 3 9 1 10 11 1 11 2
11 15 13 1 11 11 1 10 11 7 11 2
46 10 0 9 13 9 1 15 1 10 9 1 10 9 0 1 11 2 13 10 0 9 0 1 11 3 1 10 9 1 10 9 7 13 10 9 0 0 2 1 10 9 0 0 7 0 2
17 10 0 9 13 1 10 10 9 1 10 9 2 9 7 9 0 2
11 15 13 10 9 7 3 15 13 10 9 2
39 10 9 13 10 9 0 1 10 9 7 4 7 13 15 3 16 10 9 1 9 1 9 1 10 9 1 10 9 7 1 10 9 1 10 9 4 13 9 2
39 10 9 13 13 15 1 10 11 2 1 11 7 10 9 1 11 1 11 7 11 2 7 13 9 1 10 9 1 10 9 1 10 11 7 10 9 1 11 2
107 1 10 9 3 0 1 12 15 13 12 1 10 12 9 1 9 13 1 10 11 11 2 10 11 11 2 12 2 1 10 12 13 2 12 9 1 10 9 0 2 8 1 12 2 8 1 12 7 8 1 12 2 2 12 0 9 1 10 9 0 2 12 7 12 2 1 12 9 1 10 12 9 1 10 9 7 12 11 11 2 12 7 12 2 2 9 16 13 1 10 9 1 10 0 9 7 1 10 15 11 9 0 1 10 9 0 2
44 10 9 0 7 0 2 1 10 9 1 10 9 0 7 0 2 10 9 0 2 10 9 1 10 9 2 10 9 1 9 7 10 9 0 2 13 1 16 10 9 13 9 0 2
20 1 10 9 2 13 11 10 9 1 10 9 7 3 4 13 1 11 1 12 2
16 7 3 11 3 13 10 9 2 13 10 0 9 1 10 9 2
15 3 2 10 9 15 13 1 10 9 1 10 9 1 11 2
15 10 9 15 13 1 11 2 12 2 7 11 2 12 2 2
16 7 3 2 15 13 10 9 2 15 4 13 15 15 1 15 2
35 1 11 1 12 2 12 9 4 13 1 10 9 1 9 2 1 11 1 12 2 9 1 9 0 13 1 10 9 7 13 1 10 10 9 2
23 10 0 9 0 13 1 11 2 1 11 7 11 11 7 13 15 10 9 0 1 10 9 2
42 1 10 9 0 9 1 9 13 0 1 12 1 10 9 1 13 9 0 2 12 9 0 2 12 9 0 2 7 16 15 13 1 10 9 0 13 13 1 0 12 9 2
84 10 9 1 15 11 1 10 8 13 3 2 1 9 2 13 10 9 1 11 1 15 4 13 1 11 2 11 2 11 7 11 1 10 13 16 10 9 7 9 16 10 8 13 3 2 1 9 0 2 1 10 9 11 11 2 13 1 11 11 2 10 11 2 2 13 9 1 10 9 2 11 2 1 11 2 2 4 13 10 9 1 9 0 2
30 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 5 12 7 10 9 0 1 9 13 5 12 2
51 10 9 11 13 16 16 3 13 10 9 0 0 1 10 9 1 9 7 13 15 0 1 10 9 3 0 2 13 0 16 10 9 13 10 9 1 10 9 2 1 9 1 10 9 9 1 9 1 10 9 2
19 4 7 13 16 10 9 4 13 1 11 11 2 9 1 9 1 11 11 2
14 1 10 9 13 10 9 13 1 9 0 2 11 11 2
22 11 11 4 13 1 12 2 1 10 9 1 10 9 1 11 11 11 1 11 2 11 2
11 15 13 16 15 13 16 4 13 1 9 2
28 10 9 13 10 9 1 10 9 1 9 1 11 2 7 10 9 1 10 9 1 10 9 1 0 9 1 11 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
9 10 9 0 4 7 13 15 0 2
48 10 9 0 1 10 11 1 11 2 11 11 2 13 9 3 16 10 9 3 3 4 13 10 9 0 1 10 9 1 10 9 0 2 1 10 16 15 13 1 10 11 11 7 1 10 11 11 2
6 13 12 9 1 12 2
25 1 15 2 15 13 1 10 9 0 1 16 13 10 9 7 13 16 3 15 13 1 9 0 0 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 9 2
23 10 0 9 1 10 9 15 13 13 1 9 0 2 3 15 4 13 10 0 9 7 9 2
14 3 15 13 16 13 1 10 9 0 2 3 15 4 2
28 15 13 10 9 1 16 10 9 4 4 13 1 10 9 1 13 3 1 10 9 1 10 9 2 1 3 0 2
34 3 3 13 9 1 10 9 0 1 10 9 9 2 3 7 4 13 3 1 9 1 10 9 12 2 9 1 10 15 4 10 0 9 2
14 13 10 0 9 1 9 0 1 10 15 15 13 9 2
19 3 3 2 15 13 1 10 9 1 11 2 1 10 9 1 11 7 11 2
62 10 9 1 12 7 12 1 13 10 9 0 2 16 13 1 11 11 10 9 0 9 1 10 10 9 0 2 13 10 9 2 7 10 9 0 13 1 10 9 1 10 9 0 2 1 10 11 11 2 4 13 1 13 16 10 9 3 3 4 13 15 2
9 2 13 3 1 15 1 15 2 2
54 11 3 11 13 10 9 0 1 10 9 1 9 1 11 11 2 15 1 10 9 1 11 11 7 3 15 1 10 9 1 10 9 0 1 11 11 2 9 1 9 1 10 11 11 2 10 9 1 11 7 10 9 0 2
61 11 11 13 16 15 3 15 13 1 2 0 9 2 7 2 13 0 1 10 9 2 1 9 2 2 1 9 1 10 9 1 10 9 1 11 10 11 2 11 11 11 2 15 13 1 10 9 1 2 13 1 9 2 16 13 10 2 9 0 2 2
21 3 13 12 2 9 1 10 9 2 13 1 11 7 11 2 11 2 11 11 8 2
8 13 7 13 11 11 1 11 2
20 7 15 3 9 13 16 13 9 7 9 1 13 15 16 13 15 2 2 13 2
55 3 2 10 9 15 4 13 1 10 2 9 8 2 0 2 2 13 1 10 9 16 13 10 9 1 10 9 1 10 9 1 10 9 11 1 10 11 1 10 9 0 2 1 10 9 16 13 3 1 10 9 1 10 11 2
45 13 1 10 9 1 10 9 1 11 3 15 13 10 0 9 1 10 9 2 2 13 10 9 2 15 13 13 2 10 0 9 2 7 3 0 2 1 11 11 2 10 9 1 11 2
22 3 1 10 9 1 13 1 10 9 2 2 13 0 4 7 13 16 3 1 13 9 2
14 11 13 10 9 1 11 12 7 12 1 11 1 12 2
30 13 13 15 1 10 9 0 1 10 11 11 1 10 9 2 12 2 7 10 9 16 13 1 10 9 0 7 10 9 2
21 1 9 0 10 9 4 13 1 10 13 9 0 2 1 9 2 9 7 1 9 2
34 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 11 2 1 10 9 1 11 7 9 1 11 2 11 2 11 2
26 10 11 1 10 11 7 9 1 10 11 1 10 11 13 10 9 0 13 1 10 9 1 9 1 9 2
10 10 0 9 13 12 9 7 12 9 2
10 15 13 15 13 10 9 1 11 11 2
39 1 10 9 0 2 13 1 11 1 9 1 9 1 10 9 11 11 11 2 1 15 13 1 11 16 13 10 9 0 1 10 15 13 13 1 10 9 0 2
11 15 13 1 9 0 2 9 1 12 2 2
14 10 0 9 1 9 1 15 4 13 10 9 1 15 2
31 1 10 9 0 1 10 9 0 2 1 10 16 13 10 3 0 9 2 13 13 10 9 1 10 9 16 13 13 10 9 2
38 10 9 1 11 11 13 9 1 10 9 11 11 1 10 9 1 11 2 11 2 13 3 1 10 9 0 0 1 10 9 1 10 11 2 9 11 2 2
6 0 16 3 15 13 2
11 7 1 15 10 9 7 9 13 3 0 2
27 10 12 1 11 1 12 2 13 1 10 9 1 10 9 7 5 12 9 1 9 1 10 11 1 11 11 2
30 10 9 13 15 1 10 9 0 1 10 11 11 2 4 13 1 10 9 1 10 11 11 1 10 12 1 11 1 12 2
9 1 9 2 9 0 2 1 0 2
17 1 11 1 10 9 12 2 13 1 9 7 15 13 1 10 11 2
20 15 13 10 9 7 9 2 3 15 13 10 0 9 1 10 9 1 10 9 2
51 16 15 13 16 10 9 7 10 9 13 10 9 2 15 13 3 0 2 7 2 1 13 2 10 9 7 10 9 13 0 7 4 13 1 10 9 2 16 13 3 13 3 1 15 16 1 11 13 9 2 2
24 1 12 10 9 1 9 11 2 11 13 10 0 9 16 15 13 1 10 11 11 1 10 9 2
33 10 9 4 4 13 3 1 10 9 1 11 2 13 10 0 9 1 9 1 10 9 9 1 9 1 10 9 0 1 12 9 9 2
12 10 9 11 13 15 1 10 9 1 10 11 2
51 10 9 4 13 1 10 12 5 2 10 9 1 10 12 5 2 10 9 1 10 12 5 2 10 9 1 10 12 5 2 10 9 1 10 12 5 2 7 10 10 9 2 1 10 9 2 1 10 12 5 2
41 10 9 16 13 10 9 1 10 9 1 10 11 13 13 9 1 10 9 7 10 9 1 10 9 2 13 15 16 10 9 15 13 1 9 1 10 9 1 10 9 2
25 10 9 13 9 1 10 10 9 0 2 0 2 0 2 0 16 13 1 10 0 9 0 1 11 2
27 15 4 13 1 10 9 1 9 13 1 10 9 7 10 9 7 2 1 10 9 2 10 9 1 10 9 2
10 3 2 13 10 0 9 1 12 9 2
10 13 10 8 13 1 10 9 1 11 2
54 10 9 13 1 10 9 12 12 9 1 9 0 7 12 12 3 13 1 10 9 2 16 7 10 9 13 9 1 12 12 9 1 9 2 1 10 9 1 12 7 12 12 9 1 9 15 13 1 10 9 1 10 9 2
29 11 4 13 1 10 9 0 1 11 2 7 1 3 9 13 1 10 9 1 10 12 9 2 3 1 10 9 13 2
24 9 1 10 9 2 0 7 3 2 16 13 1 10 9 1 11 13 2 10 9 7 9 0 2
13 10 9 0 1 10 9 1 11 11 13 12 9 2
17 13 10 9 0 1 10 9 1 11 1 11 2 0 7 3 0 2
10 1 10 9 3 0 1 10 9 13 2
25 9 1 9 0 13 3 1 10 9 16 13 3 1 12 9 2 1 9 1 10 9 1 9 0 2
24 10 9 15 13 1 10 8 2 9 1 10 9 0 11 2 11 11 2 11 11 7 11 11 2
19 10 12 15 13 10 9 3 13 0 9 0 2 13 10 9 0 7 0 2
13 4 13 1 12 7 13 1 10 11 11 1 11 11
7 2 1 15 13 10 9 2
25 11 11 11 11 2 2 11 2 2 13 1 12 7 13 10 9 1 10 9 0 11 11 1 11 2
62 10 9 13 9 1 10 9 1 3 2 11 2 1 10 9 0 1 11 2 16 10 9 0 2 16 15 13 1 10 9 1 11 2 0 1 11 7 10 9 2 16 13 1 11 2 13 3 1 10 9 1 10 9 12 2 1 10 9 1 10 11 2
28 10 9 1 10 9 13 16 2 3 1 0 9 2 10 12 1 11 1 12 15 13 1 10 9 1 10 9 2
18 15 13 1 12 9 0 3 13 1 12 9 1 9 7 1 12 9 2
9 11 7 11 13 1 13 10 9 2
19 15 13 1 10 9 2 7 1 10 9 4 13 1 9 1 13 1 11 2
55 10 12 1 11 10 11 11 1 9 13 1 12 9 0 2 12 9 7 12 9 2 1 9 1 10 9 0 1 11 1 11 2 16 13 12 9 1 9 0 7 16 13 1 10 9 2 2 11 1 10 9 1 11 2 2
14 13 1 10 9 0 1 10 16 10 9 13 10 9 2
12 10 9 2 9 2 13 1 10 9 1 13 2
15 10 10 9 4 7 13 3 1 10 9 13 1 11 11 2
29 3 2 1 10 9 12 2 13 10 0 9 13 11 1 11 2 1 9 1 10 11 11 11 2 9 1 10 9 2
8 2 13 16 10 9 13 0 2
31 11 11 15 13 1 10 9 1 9 0 2 0 0 2 13 1 10 9 1 10 9 2 11 11 11 2 1 9 1 9 2
10 16 13 3 3 4 13 2 0 13 2
30 11 13 4 15 13 1 10 9 7 10 9 0 1 10 9 7 9 16 1 10 9 4 13 9 1 10 9 0 2 2
17 10 9 1 10 9 15 13 10 9 1 2 10 11 1 11 2 2
10 11 4 13 10 12 1 11 1 12 2
25 10 9 1 9 13 10 0 9 1 10 9 2 16 13 3 1 9 1 10 9 2 9 7 9 2
20 1 10 9 0 2 11 0 4 13 10 9 1 9 1 10 9 7 10 9 2
38 11 1 11 4 13 10 11 11 16 13 10 9 0 1 10 11 11 9 1 10 9 16 15 13 1 10 11 11 11 1 11 2 1 10 0 9 0 2
45 10 9 1 10 11 0 13 1 10 9 0 7 1 10 9 1 10 9 13 1 10 9 0 1 10 11 1 11 11 2 11 2 2 10 9 0 16 13 10 9 1 10 9 2 2
15 3 15 13 1 10 9 1 10 9 11 7 10 9 0 2
41 7 3 7 15 13 15 13 2 1 10 9 3 15 4 13 1 13 2 7 1 10 9 1 9 2 16 4 13 15 16 15 4 13 3 2 3 13 1 13 15 2
32 11 11 2 1 11 2 11 2 4 13 3 1 4 13 10 9 0 1 9 16 15 4 13 10 0 9 7 10 9 3 0 2
15 1 9 1 10 9 2 13 10 9 1 9 0 0 0 2
47 10 9 1 13 1 10 9 10 9 1 10 9 0 13 10 9 1 11 2 10 0 9 1 13 13 1 10 9 1 9 0 1 10 9 0 7 0 2 13 1 9 10 9 8 10 9 2
21 10 9 3 8 10 9 1 3 1 12 9 2 12 9 2 13 1 9 0 9 2
44 10 9 2 9 1 9 2 13 10 9 1 9 1 10 9 0 2 16 3 3 15 13 1 10 9 7 1 10 9 1 9 2 7 3 4 13 15 1 4 13 1 9 0 2
20 11 11 2 8 12 1 11 1 12 2 11 2 13 10 9 1 9 0 0 2
20 10 11 11 11 2 11 2 11 2 13 10 9 0 13 1 10 9 1 11 2
29 10 9 3 13 0 9 1 10 9 7 3 3 1 10 9 1 10 0 9 2 11 11 11 2 13 10 9 12 2
31 1 10 9 2 11 13 1 15 1 10 9 1 10 9 1 9 1 10 13 10 9 1 10 9 7 13 15 1 10 9 2
49 11 13 1 10 9 2 0 2 7 2 0 2 1 10 9 2 3 1 11 11 7 11 11 2 16 13 16 10 9 7 10 9 13 9 1 10 9 7 4 4 13 1 9 1 9 0 7 0 2
15 11 11 13 10 0 9 1 9 1 11 2 12 2 11 2
23 0 9 1 10 9 0 13 9 1 10 9 0 0 7 15 1 10 9 13 1 9 9 2
56 1 10 9 13 1 9 13 10 9 1 10 11 1 10 11 2 15 1 10 0 9 1 10 9 2 7 10 9 1 10 9 11 2 16 13 10 9 1 10 12 9 7 10 9 1 10 0 9 1 10 9 2 10 11 2 2
11 13 1 9 7 10 0 9 13 11 11 2
8 15 4 13 0 1 9 0 2
47 1 11 1 12 2 10 9 13 10 9 0 1 9 2 1 15 10 9 1 12 9 2 5 1 10 9 1 12 9 2 7 10 9 1 12 9 2 5 1 10 9 1 12 2 12 9 2
23 1 9 2 11 13 3 0 1 11 11 2 10 0 9 2 16 4 13 13 1 10 9 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
39 11 11 13 10 9 0 1 10 9 1 9 1 9 7 8 2 11 11 11 2 1 15 1 9 1 9 1 9 2 1 9 0 2 1 9 1 9 8 2
8 13 10 12 1 11 1 12 2
27 3 2 11 2 3 16 13 1 11 2 13 10 12 9 7 13 16 10 16 3 15 4 4 13 13 15 2
29 13 1 11 1 10 9 12 1 11 9 7 13 10 0 9 1 11 2 7 4 13 1 11 11 3 1 12 9 2
4 13 1 9 2
20 11 11 11 2 11 2 11 11 2 12 1 11 1 12 2 13 10 9 0 2
14 1 11 2 10 9 4 13 1 10 9 11 2 8 2
35 11 2 1 10 9 1 9 2 11 7 10 9 11 2 4 7 13 3 1 11 11 7 1 10 9 1 16 3 13 1 9 10 0 9 2
24 10 9 1 10 9 15 13 1 9 2 13 1 10 9 1 9 1 11 7 10 9 1 9 2
16 1 13 10 9 1 9 2 10 9 0 3 13 10 9 0 2
35 1 10 9 1 10 9 1 13 12 9 1 9 2 10 9 13 1 10 9 1 13 15 10 0 9 1 9 1 10 9 1 10 9 12 2
15 10 9 1 9 7 9 13 3 16 15 13 1 10 9 2
12 13 9 0 1 10 9 13 1 8 2 8 2
10 13 10 9 0 1 9 1 10 11 2
21 1 11 1 12 4 13 1 10 12 5 11 2 5 2 2 12 5 11 1 11 2
30 1 10 9 1 12 1 15 1 10 9 0 10 9 13 3 2 1 13 9 1 10 9 1 10 9 1 10 9 0 2
38 10 9 13 10 9 1 13 1 10 12 9 0 1 10 9 2 11 11 2 11 11 2 11 11 7 11 11 2 1 10 0 9 1 9 11 1 12 2
12 1 9 13 1 10 9 0 1 2 11 2 2
115 10 9 15 13 1 10 9 1 9 1 10 11 11 1 10 9 1 10 11 1 9 2 13 15 1 10 9 1 0 9 1 9 0 7 0 2 1 9 1 9 0 13 1 8 0 1 10 11 2 1 15 15 10 9 13 1 0 9 10 9 1 9 2 0 7 3 0 2 3 10 9 0 13 1 9 0 16 15 13 1 10 9 2 13 15 10 0 9 1 9 0 2 9 2 9 2 9 2 2 7 1 10 9 0 16 15 13 1 9 1 10 12 8 8 2
34 10 9 3 0 7 1 10 9 3 0 2 13 10 1 13 10 9 0 1 10 9 1 10 0 1 10 9 1 10 9 1 10 9 2
27 1 10 9 2 11 15 13 3 1 11 3 1 4 15 13 15 0 7 13 11 10 16 15 13 1 11 2
28 3 2 1 15 8 10 9 15 13 1 3 7 15 13 1 10 9 1 10 9 11 2 1 10 9 1 11 2
50 1 0 9 4 13 15 16 9 2 8 9 7 9 0 0 2 9 1 9 2 9 0 7 9 2 13 1 16 10 9 13 3 3 1 12 9 1 9 1 9 0 1 9 0 7 2 7 0 2 2
50 11 11 2 9 0 16 13 1 11 10 9 2 13 16 11 13 1 9 0 7 1 9 0 2 13 15 2 1 10 9 2 1 15 1 10 9 2 15 1 9 0 2 13 9 0 0 1 10 9 2
21 10 9 3 13 1 10 9 1 10 9 11 7 10 9 2 11 11 1 11 2 2
39 15 3 9 1 10 9 13 16 10 0 9 13 1 10 0 9 1 10 9 15 4 13 1 13 10 9 2 7 3 13 0 9 13 1 9 1 10 15 2
14 15 13 1 10 11 11 2 13 1 11 11 1 12 2
18 1 12 2 13 10 0 9 2 11 1 10 9 2 1 11 2 11 2
33 10 9 1 10 9 13 10 9 0 1 9 0 13 1 12 2 13 1 11 11 7 13 1 11 1 11 2 11 11 7 11 11 2
12 1 0 9 10 9 0 15 13 1 10 9 2
28 3 2 1 10 9 1 10 9 1 10 11 2 4 13 16 1 10 9 13 1 10 9 1 10 9 1 9 2
12 11 11 13 10 9 1 9 1 10 9 11 2
20 1 10 9 12 7 1 9 1 10 11 12 2 11 13 10 0 9 0 0 2
27 11 2 1 10 3 7 10 12 9 2 13 1 11 2 11 2 9 1 10 9 7 1 10 9 1 9 2
30 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 5 12 7 10 9 0 1 9 13 5 12 2
52 11 11 4 13 1 16 10 9 13 1 10 9 0 1 10 11 2 2 1 10 9 9 1 13 10 9 0 16 13 15 1 10 9 1 10 9 7 1 10 9 2 16 13 1 0 9 8 10 9 0 2 2
11 11 4 7 13 10 9 1 3 12 5 2
18 11 11 13 1 9 0 2 1 0 9 2 16 4 13 1 12 9 2
34 1 9 1 10 9 2 1 12 2 15 13 1 10 9 10 9 1 9 0 1 12 8 2 7 9 1 9 0 1 12 7 12 8 2
11 11 13 9 1 10 9 0 1 10 9 2
30 1 10 9 12 2 3 1 10 0 9 2 13 1 10 9 1 11 11 2 7 1 10 9 1 11 11 2 8 2 2
8 11 15 13 13 1 10 9 2
30 9 1 9 2 9 2 9 1 9 7 9 0 4 13 10 9 1 9 2 9 7 9 1 11 1 11 7 11 11 2
28 11 11 2 10 9 0 9 1 10 9 10 11 2 13 10 0 9 7 13 9 1 10 9 1 10 12 9 2
19 3 13 10 0 9 0 1 10 9 11 11 13 1 10 9 0 11 11 2
18 3 0 9 1 9 2 7 13 3 0 7 10 9 3 13 3 0 2
3 1 9 2
36 1 15 2 13 0 16 15 11 15 13 7 15 13 0 1 10 9 16 13 10 9 7 16 13 3 2 1 9 2 16 13 0 7 0 9 2
98 11 7 11 13 10 9 2 10 9 11 2 13 10 9 2 11 2 9 1 10 11 11 1 10 9 1 10 9 9 11 12 2 11 1 11 2 0 9 1 10 9 2 9 7 9 1 10 9 2 10 0 11 12 2 11 2 9 1 11 11 1 11 2 9 1 11 7 11 2 11 2 9 1 11 2 11 2 13 1 11 11 1 11 2 9 1 11 2 7 11 2 9 0 2 0 9 0 2
37 1 13 1 10 9 1 11 2 10 9 13 10 9 1 12 9 0 2 1 10 0 9 1 10 9 0 13 3 1 10 9 2 7 10 0 9 2
47 9 0 7 0 1 12 1 12 9 1 0 7 1 12 1 12 9 0 2 1 12 1 12 9 1 0 10 15 2 1 9 0 0 16 13 1 10 0 9 0 1 10 9 1 10 9 2
48 10 9 13 10 0 9 16 15 13 1 13 10 9 2 10 9 2 9 1 10 9 2 13 1 9 0 2 16 4 13 15 7 13 15 2 13 1 9 0 7 2 1 10 9 2 3 0 2
10 4 13 10 9 0 1 10 9 0 2
43 13 10 9 1 11 11 2 12 2 7 1 10 9 1 11 13 2 10 9 1 11 11 1 11 2 13 3 1 11 1 11 2 10 9 1 11 11 2 11 1 10 11 2
36 13 3 1 10 9 0 1 10 0 9 1 10 9 2 7 10 0 9 1 10 9 13 1 10 9 1 10 11 11 13 10 9 1 10 9 2
22 16 10 9 4 1 13 10 9 1 15 9 1 10 9 2 11 3 4 13 10 9 2
9 1 12 13 1 10 11 1 11 2
4 13 3 0 2
24 10 9 0 11 11 11 13 10 9 1 10 9 1 10 9 1 10 9 0 2 3 0 2 2
29 11 1 10 11 2 13 10 9 0 1 10 11 2 1 10 9 1 12 9 0 1 9 1 9 3 7 10 9 2
45 1 9 1 10 9 1 10 12 11 13 1 10 9 11 11 7 10 0 11 11 2 12 2 1 10 11 2 0 13 9 0 1 11 7 13 1 10 9 2 16 3 13 0 9 2
17 10 9 0 2 9 13 10 11 1 11 7 15 13 3 1 11 2
24 11 2 12 2 15 13 1 9 7 3 13 1 12 9 0 1 16 10 9 15 13 1 12 2
23 10 0 9 13 10 0 9 1 9 0 2 9 2 9 2 9 7 9 1 9 3 0 2
9 13 15 10 9 7 10 9 0 2
18 10 9 1 10 9 0 0 2 9 2 2 4 13 3 1 10 9 2
21 1 12 2 16 13 1 9 1 11 11 2 11 2 11 11 7 11 11 11 11 2
17 11 11 11 2 8 11 11 2 11 2 12 1 11 1 12 2 2
16 10 9 1 9 0 15 13 1 11 10 12 1 11 1 12 2
14 2 15 13 9 0 2 7 3 10 9 2 2 13 2
50 10 11 1 10 11 1 10 9 1 9 1 11 12 13 10 9 1 10 9 1 10 9 2 3 13 1 10 9 0 2 13 9 0 0 1 10 2 11 2 2 10 9 0 1 10 11 1 10 9 2
26 1 9 2 10 0 11 13 10 9 1 9 0 1 12 9 2 11 11 11 2 11 11 7 11 11 2
38 15 3 15 13 1 10 9 0 2 7 15 13 0 1 13 10 9 2 3 7 10 9 7 9 16 13 1 10 9 13 9 1 9 2 13 10 9 2
33 11 11 11 11 2 11 2 12 1 11 1 12 2 13 10 9 1 9 0 16 13 3 1 10 11 11 2 3 15 13 1 9 2
25 10 9 13 15 0 7 10 1 10 9 0 1 9 2 7 3 0 7 15 1 9 0 9 8 2
12 10 9 4 13 13 10 12 5 1 9 0 2
14 1 12 13 1 9 2 1 15 11 2 11 7 11 2
56 13 2 1 11 1 12 2 10 0 9 1 9 1 13 10 9 1 9 1 10 9 2 1 0 10 9 1 10 9 1 9 7 1 9 2 1 10 15 3 15 13 15 2 7 15 1 10 9 1 10 9 1 10 0 9 2
21 1 10 9 16 13 10 9 2 11 13 10 9 1 10 9 1 2 11 11 2 2
17 13 15 1 10 9 0 0 1 11 11 11 1 10 11 11 11 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
27 7 3 2 10 9 1 11 7 11 13 1 10 9 0 2 16 13 10 9 1 13 9 2 9 7 9 2
42 3 1 13 12 0 9 1 10 9 1 9 2 1 11 7 11 2 2 10 9 3 13 13 1 10 9 0 1 11 2 13 10 0 9 7 10 0 9 1 11 11 2
16 3 2 4 13 1 10 9 12 9 7 4 13 15 1 15 2
11 10 9 1 12 7 12 9 13 1 9 2
12 10 9 13 4 13 10 12 9 1 9 0 2
45 1 16 1 11 1 10 12 10 9 4 13 1 10 0 9 1 9 11 2 15 15 15 13 1 10 9 2 10 9 13 1 15 7 10 9 15 13 15 3 13 1 15 15 13 2
78 10 9 0 15 13 1 10 9 1 10 9 0 2 1 10 15 13 10 11 2 9 1 10 12 9 2 13 3 1 2 8 2 2 2 10 11 2 9 0 1 9 2 2 10 9 2 9 1 9 2 2 10 11 2 9 0 2 2 7 10 9 2 12 9 1 9 1 3 12 9 13 1 10 9 7 9 2 2
26 10 9 1 10 9 13 16 10 9 1 11 1 11 7 1 11 13 10 0 9 0 1 10 9 0 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
5 10 9 0 13 2
50 10 9 3 0 15 13 3 1 10 9 1 10 9 1 10 9 2 1 9 2 8 15 13 1 10 9 1 9 2 8 15 13 1 10 9 1 9 0 2 8 15 13 1 10 9 1 9 0 2 8
10 10 0 9 13 10 9 11 1 11 2
14 7 1 15 15 13 1 10 9 0 2 16 13 13 2
11 10 9 13 10 9 0 1 10 9 12 2
20 15 13 1 11 2 9 1 10 9 11 11 7 11 3 1 11 2 11 2 2
18 16 10 0 9 2 11 2 15 13 3 0 2 3 13 1 15 13 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
35 3 2 13 1 10 9 1 13 9 1 9 7 9 0 1 9 1 10 9 0 16 2 13 10 0 9 0 1 15 16 4 1 13 2 2
35 10 9 11 11 15 13 13 1 11 1 10 9 1 10 9 0 2 3 13 1 13 1 12 9 16 4 4 13 1 10 9 1 10 9 2
17 11 13 10 9 1 10 9 11 11 1 10 9 13 1 11 11 2
5 1 9 0 0 2
39 3 1 10 9 0 1 10 9 13 13 1 9 3 0 10 9 0 1 11 11 2 13 1 12 2 1 10 15 15 13 0 9 1 10 9 12 7 12 2
10 10 0 9 13 1 10 11 1 11 2
23 13 10 9 13 15 10 15 1 9 7 13 15 10 9 1 9 3 7 15 13 10 9 2
40 15 15 13 1 11 13 1 3 1 10 9 1 10 9 2 13 9 3 1 10 9 0 2 9 1 9 0 1 10 9 0 2 16 13 1 13 10 0 9 2
8 1 15 15 13 3 12 9 2
44 1 10 9 1 12 11 4 13 1 10 9 1 10 9 2 7 1 9 1 10 9 1 12 13 10 9 11 2 11 7 11 2 9 2 1 10 9 7 13 10 9 11 0 2
10 15 13 1 10 11 11 1 10 11 2
21 1 15 13 9 0 1 10 9 0 0 1 10 9 2 1 11 11 7 11 11 2
15 10 9 1 9 15 13 3 3 0 1 13 10 11 11 2
25 10 9 4 4 13 1 10 11 7 2 1 9 1 11 11 2 1 3 1 12 9 1 10 11 2
67 10 9 1 11 11 7 11 2 16 13 10 9 0 2 2 3 13 1 11 11 2 13 10 9 1 9 0 16 13 3 1 10 11 1 12 1 12 7 1 12 1 10 9 7 3 9 1 13 2 1 10 9 1 9 0 1 11 7 1 10 9 1 11 1 11 11 2
33 10 9 1 10 9 0 15 13 1 10 0 9 2 13 1 10 9 1 10 9 13 1 10 9 1 10 9 0 2 16 13 9 2
62 10 12 1 11 1 12 11 11 11 7 11 1 11 4 3 13 1 10 11 1 11 1 11 12 1 11 2 9 1 11 1 11 2 16 15 4 13 2 7 9 11 11 2 15 13 1 10 9 0 7 0 1 10 9 1 10 9 2 11 1 11 2
22 1 9 0 13 1 11 1 9 1 9 2 13 1 10 9 1 10 9 13 1 11 2
44 13 10 9 7 13 1 10 15 1 9 1 10 11 2 1 11 7 3 13 11 2 3 13 10 9 2 3 13 1 12 9 2 13 1 12 3 9 1 10 9 0 1 11 2
31 13 0 9 1 9 7 9 1 13 7 13 10 11 11 7 10 11 2 7 1 0 9 13 9 2 9 2 9 7 9 2
10 2 2 10 9 13 10 9 1 9 2
12 1 15 1 10 9 13 10 9 1 10 9 2
11 15 13 10 0 9 1 10 10 9 2 2
15 3 13 9 1 10 11 1 10 11 1 11 11 1 12 2
19 10 11 11 1 11 13 10 0 9 1 11 1 9 2 9 7 9 0 2
30 10 9 0 13 0 1 10 9 1 9 0 2 3 13 1 10 9 2 7 10 9 1 9 1 10 9 1 10 11 2
17 13 1 11 11 11 11 11 12 7 1 11 11 11 11 12 11 2
35 9 1 9 13 10 9 1 9 1 9 2 9 7 9 3 1 9 1 10 9 1 9 0 7 13 1 9 0 1 9 1 9 7 0 2
16 3 15 13 16 1 10 9 1 13 10 9 3 15 13 15 2
27 15 13 1 10 9 0 7 0 0 2 13 13 2 1 10 9 7 1 10 9 0 2 1 9 0 2 2
32 1 10 9 2 10 9 1 10 9 13 10 10 9 0 9 1 10 9 7 10 9 1 9 1 10 9 3 15 13 3 0 2
55 13 1 9 7 15 13 1 10 8 2 8 1 11 1 10 16 15 13 16 4 13 10 9 7 16 15 13 1 9 1 10 9 1 10 16 13 10 9 3 7 13 0 10 9 1 10 9 7 3 4 4 13 10 9 2
30 11 2 1 9 1 9 0 1 16 13 10 9 1 12 2 13 1 10 9 10 9 1 10 0 9 0 2 11 11 2
17 10 11 11 4 13 1 11 1 10 0 9 1 10 11 2 11 2
27 3 13 9 0 1 11 11 11 1 12 5 2 11 11 12 5 2 11 11 12 5 7 10 11 12 5 2
33 10 9 1 10 9 0 4 13 1 0 16 15 4 13 1 3 10 9 1 10 0 9 1 15 7 1 3 10 9 4 3 13 2
61 10 9 2 10 9 0 1 10 9 2 3 4 13 1 11 11 2 16 15 15 13 1 10 9 2 7 11 13 9 1 10 9 1 10 9 7 15 13 1 3 0 1 10 9 16 13 10 9 0 2 13 16 11 15 13 15 7 3 4 13 2
15 15 13 10 9 13 1 9 2 15 13 3 10 11 11 2
88 9 0 0 1 10 9 1 9 4 13 10 9 0 1 10 9 2 10 9 1 9 0 2 10 9 1 9 1 10 9 3 7 10 0 9 1 9 16 4 7 13 1 10 9 1 9 1 9 1 13 10 9 2 9 9 7 11 2 7 1 9 1 16 13 10 9 2 9 1 9 1 10 9 2 9 1 10 9 1 9 1 16 3 13 0 2 8 2
25 3 13 7 1 10 12 1 11 15 3 13 13 10 9 1 10 9 2 1 10 9 1 10 9 2
20 7 16 10 12 9 13 9 1 10 11 11 2 11 13 9 1 11 10 9 2
39 10 9 15 13 1 10 9 0 1 11 2 9 16 1 10 9 15 13 1 15 1 10 12 9 16 13 1 10 9 1 11 2 10 0 9 12 1 11 2
42 11 11 15 4 13 3 1 9 0 2 3 16 11 11 4 13 10 9 1 10 9 1 11 2 11 2 11 11 2 11 11 2 11 2 11 2 11 2 11 7 11 2
48 1 10 9 1 9 2 11 2 11 2 11 2 11 7 11 2 10 9 0 13 1 9 7 9 0 2 4 13 2 16 13 0 2 1 9 0 16 13 10 0 9 1 10 9 1 10 9 2
34 11 2 15 13 2 13 1 11 2 7 13 2 16 13 0 1 13 15 1 10 9 1 10 9 7 1 10 3 1 15 1 15 2 2
22 10 9 1 10 9 13 10 9 1 9 2 9 2 9 2 9 2 9 0 7 9 2
11 10 9 13 1 10 1 10 9 1 9 2
20 11 13 10 9 7 10 9 0 0 2 1 11 7 11 2 11 2 11 2 2
18 10 9 1 10 9 1 12 9 2 1 9 1 1 12 9 1 0 2
9 10 9 0 0 13 10 0 9 2
31 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 9 12 2 7 10 9 0 1 9 13 9 12 2
20 10 9 4 13 9 9 1 9 0 1 12 1 10 0 9 1 9 0 0 2
19 9 3 3 13 1 10 9 1 11 2 11 2 2 1 10 15 13 9 2
23 1 3 2 10 9 13 7 10 9 1 9 4 7 13 2 3 7 3 2 1 9 0 2
26 2 11 11 11 11 11 2 2 15 3 13 10 9 2 13 10 9 16 10 9 15 13 1 10 9 2
16 3 14 1 10 9 1 11 10 9 13 3 0 7 3 0 2
29 1 10 9 1 10 9 2 0 1 9 1 9 2 10 9 11 13 10 9 0 9 0 7 9 2 9 1 9 2
18 11 11 2 9 1 10 11 2 13 10 9 1 10 11 1 10 11 2
13 3 15 15 13 16 3 4 13 15 7 16 13 2
21 0 9 1 10 9 13 10 9 1 10 9 0 16 13 2 7 10 9 1 9 2
15 3 3 4 13 1 10 9 1 9 1 10 9 3 0 2
17 1 0 9 2 0 13 10 9 1 9 0 10 9 13 9 0 2
42 11 2 1 9 2 15 13 9 15 13 0 9 1 10 9 11 7 13 10 9 1 10 9 1 11 8 11 11 2 15 15 13 1 10 9 7 3 9 0 1 11 2
27 10 11 13 1 10 9 0 13 1 10 11 2 7 13 9 1 10 11 11 11 11 1 10 9 1 12 2
43 1 10 9 1 10 9 1 10 11 11 2 10 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
23 10 9 13 13 1 10 9 7 10 9 1 9 1 10 9 12 1 10 9 11 11 11 2
13 2 3 13 15 1 15 13 2 7 1 15 0 2
13 11 13 10 9 0 1 9 0 1 10 9 11 2
41 1 10 11 1 11 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
51 13 10 9 1 10 9 1 10 9 1 10 15 15 13 10 9 2 11 15 13 0 1 10 9 2 10 9 11 11 2 1 15 3 13 3 1 13 15 2 7 15 13 13 15 13 10 9 1 10 9 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
27 1 9 2 4 3 13 1 10 9 1 9 1 4 13 9 1 10 9 0 2 3 13 10 9 1 11 2
6 11 11 2 9 2 2
27 15 13 1 10 9 13 1 10 9 15 13 1 13 10 11 1 10 9 1 10 9 0 2 13 9 0 2
26 15 13 10 9 1 9 1 9 2 1 9 7 1 9 2 7 3 3 1 10 9 1 9 7 9 2
12 10 9 2 1 15 9 2 13 1 9 0 2
10 13 10 11 11 11 1 9 1 15 2
36 1 9 2 13 1 15 2 13 7 13 9 7 9 1 10 9 2 1 10 9 13 3 9 2 3 13 0 16 13 10 9 13 1 10 9 2
6 10 9 13 3 0 2
24 10 9 1 9 13 3 13 10 9 1 9 1 10 0 9 1 15 1 10 8 1 10 9 2
9 4 13 1 10 9 0 1 12 2
48 10 9 1 10 9 4 13 15 2 16 15 13 2 9 1 10 9 11 2 3 15 13 10 9 0 1 9 16 13 1 10 9 1 9 0 2 13 10 9 9 2 9 2 9 7 9 2 2
39 1 15 1 10 9 16 13 1 10 9 1 10 9 2 11 11 2 1 10 15 13 1 10 9 11 11 2 2 15 13 1 9 1 10 9 1 10 9 2
17 10 9 15 13 13 1 12 1 12 9 7 3 15 13 7 13 2
48 16 3 15 4 13 10 9 0 2 10 9 1 9 13 13 1 10 9 2 1 13 1 10 12 9 1 9 0 2 7 13 16 10 9 4 13 10 9 1 2 9 1 0 9 1 9 2 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
22 15 13 1 10 9 7 3 4 13 15 2 7 9 0 7 9 1 9 2 2 13 2
14 10 0 9 13 1 9 1 12 2 16 13 12 9 2
12 15 13 10 9 1 10 9 2 15 13 2 2
26 11 11 13 9 1 9 1 10 9 1 12 2 13 10 0 9 1 10 9 2 0 1 10 9 0 2
15 10 9 0 13 10 9 1 11 11 7 11 15 13 0 2
38 2 15 4 13 10 0 9 1 10 9 2 10 0 9 1 9 2 9 1 16 15 3 13 0 7 3 15 4 13 10 15 16 15 13 2 2 13 2
27 10 12 1 11 1 12 3 15 13 10 9 1 10 0 9 2 11 11 7 10 9 1 10 9 1 9 2
13 13 12 11 1 11 2 13 10 1 0 9 0 2
18 10 9 0 13 12 5 8 12 5 8 7 10 9 13 1 12 8 2
25 10 9 13 10 9 7 9 3 0 2 16 15 13 1 10 9 3 0 2 4 13 15 3 0 2
15 9 0 2 9 1 10 9 0 1 10 9 1 10 9 2
61 1 3 2 11 13 3 3 12 9 1 9 7 1 10 9 1 9 4 13 1 10 9 0 1 11 2 1 10 9 1 11 2 1 10 9 1 11 1 11 2 3 13 10 9 1 10 9 0 7 0 16 15 13 10 9 0 7 10 9 0 2
16 13 1 9 1 9 10 9 1 11 2 0 11 2 11 2 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
28 1 13 10 9 1 11 2 4 13 1 13 1 11 10 9 0 13 10 12 1 11 0 1 10 9 1 11 2
17 11 11 2 13 10 9 1 9 0 9 1 10 9 1 10 9 2
35 10 9 0 2 13 13 1 9 0 2 1 10 16 13 1 10 11 2 11 2 13 10 9 1 10 9 11 2 13 1 10 9 1 11 2
18 16 13 1 11 11 8 11 2 10 9 1 3 9 1 10 11 11 2
29 3 1 12 13 10 9 1 13 1 15 10 9 2 10 9 1 9 7 10 0 11 16 10 9 7 9 0 13 2
37 10 9 1 10 9 2 1 9 2 13 2 13 10 9 10 9 1 10 9 2 13 1 10 0 9 2 7 16 11 13 1 10 9 1 10 9 2
23 10 0 9 1 11 2 1 9 2 13 1 3 12 9 1 10 9 1 10 9 1 11 2
11 15 13 10 9 0 7 10 9 1 9 2
19 11 15 13 9 2 7 2 1 9 1 15 2 15 13 13 1 10 9 2
11 1 15 2 10 9 13 10 9 1 9 2
41 11 11 15 13 3 1 10 11 2 11 2 10 9 1 9 0 13 1 11 2 7 1 15 13 1 10 9 2 16 4 1 13 1 10 9 0 13 1 10 11 2
12 1 10 9 1 11 15 4 13 10 9 0 2
133 11 1 11 11 7 11 13 10 9 1 12 1 11 1 11 7 13 10 12 1 11 1 12 1 11 1 11 2 9 0 1 10 11 1 11 2 12 9 1 11 1 11 2 11 1 11 2 9 0 1 11 1 10 11 7 9 0 1 10 11 2 9 1 10 11 1 11 2 9 1 9 7 3 1 9 1 10 9 1 11 12 7 11 12 2 9 7 9 0 1 10 9 1 11 2 9 1 10 11 1 9 1 11 12 7 1 11 11 2 9 7 9 0 1 10 9 1 9 2 9 1 10 11 1 11 2 9 1 10 11 1 11 2
13 10 9 1 9 13 1 12 8 2 5 9 5 2
26 1 10 9 2 13 1 10 9 11 2 8 1 11 11 2 11 7 10 9 7 9 1 9 11 11 2
11 9 1 10 0 9 0 1 10 15 0 2
28 15 15 13 1 13 1 10 9 2 1 16 11 11 2 10 9 2 1 10 15 11 13 13 15 2 15 13 2
12 13 10 12 1 11 1 12 1 11 2 11 2
33 1 9 1 12 2 13 1 11 3 2 1 0 7 13 9 2 4 13 1 11 11 11 1 13 1 10 9 1 10 12 1 11 2
11 10 10 9 13 1 10 11 11 13 9 2
19 10 9 2 13 1 11 11 2 13 10 0 9 15 1 9 1 1 9 2
26 10 9 13 13 7 13 10 9 16 13 15 1 10 9 1 10 9 0 2 15 16 1 11 13 15 2
29 13 1 10 9 12 1 10 11 1 11 1 12 9 1 11 1 10 12 2 13 10 12 5 9 0 13 1 11 2
10 10 9 4 4 13 1 10 9 0 2
28 10 9 1 10 9 0 13 10 9 0 2 16 15 1 10 9 2 13 16 3 13 10 9 1 13 10 9 2
14 3 13 10 9 2 7 13 13 10 9 1 10 9 2
26 10 12 5 1 10 9 15 13 1 10 9 1 10 8 9 0 7 10 12 5 1 15 1 10 9 2
11 3 13 10 9 1 10 9 7 10 9 2
20 10 9 13 3 0 7 3 15 13 1 10 9 1 10 9 16 4 13 2 8
42 3 1 3 10 9 13 1 12 1 11 1 10 12 2 10 9 1 10 12 5 2 7 1 13 1 11 4 1 13 10 9 1 13 10 9 16 13 13 3 12 9 2
25 1 12 13 9 1 11 7 13 1 11 1 13 10 0 9 1 12 2 13 1 11 12 9 3 2
18 1 10 9 0 2 10 9 15 13 13 3 1 10 9 1 10 9 2
32 10 9 13 16 10 9 13 3 0 2 10 9 15 13 1 10 9 2 13 3 0 2 7 10 9 3 13 3 0 7 0 2
15 13 10 9 1 10 9 1 12 9 7 10 9 1 12 2
21 10 0 9 1 10 9 0 2 13 16 13 1 0 9 16 13 1 10 8 0 2
16 9 0 2 13 15 0 7 1 3 10 9 13 1 10 9 2
25 13 13 2 16 1 10 13 10 9 10 9 13 12 7 12 2 3 15 4 13 1 10 9 0 2
22 1 10 9 1 9 1 12 5 2 1 10 15 15 13 10 9 1 9 1 12 5 2
25 10 9 0 2 10 0 9 0 9 3 13 9 1 13 10 9 1 10 9 0 1 10 9 0 2
16 10 9 1 11 2 11 7 11 1 10 9 3 3 4 13 2
12 3 13 9 10 9 11 7 11 13 1 11 2
43 1 10 9 1 10 13 1 10 9 11 2 10 9 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 13 1 9 0 7 2 12 5 2 12 5 5 13 9 2
36 1 10 9 1 13 10 9 0 2 7 3 10 9 0 2 10 11 1 11 13 12 9 0 2 10 9 0 10 11 7 10 9 0 1 11 2
57 1 9 1 10 9 1 10 9 1 10 9 2 15 13 10 9 16 4 13 0 1 10 9 2 3 13 10 9 2 9 0 2 9 2 9 2 7 9 1 9 1 10 9 2 9 2 4 13 15 0 7 3 15 1 15 2 2
19 1 11 2 16 13 10 9 0 2 7 3 0 1 10 9 1 10 9 2
11 3 3 15 13 10 9 1 10 0 9 2
31 1 15 10 9 4 13 1 13 15 1 15 3 0 10 9 13 2 3 16 10 0 9 1 9 0 15 13 15 13 0 2
41 3 13 1 11 1 12 7 10 9 13 1 9 13 1 10 9 2 12 9 3 1 4 15 13 10 9 0 7 10 12 1 11 13 1 10 9 1 10 11 11 2
8 3 13 3 0 7 11 11 2
5 3 13 3 0 2
11 10 9 0 12 7 10 9 0 12 12 2
25 13 1 11 2 11 10 12 1 11 1 12 2 13 1 11 2 11 11 10 12 1 11 1 12 2
17 9 2 9 7 9 1 9 1 10 9 0 2 10 9 0 2 8
9 10 9 1 9 13 11 7 11 2
23 4 13 1 9 10 9 2 7 10 9 3 13 7 1 12 15 13 1 10 9 1 9 2
32 13 9 3 0 7 16 13 9 2 16 13 9 7 9 16 13 15 13 7 10 9 13 15 0 7 13 1 15 1 13 15 2
40 1 10 0 9 2 10 9 7 9 13 0 2 1 10 9 0 1 12 12 9 0 2 9 1 9 2 2 13 1 10 9 3 1 12 9 16 13 10 9 2
33 10 9 4 13 1 10 9 1 9 0 7 11 11 2 3 13 1 13 1 9 1 9 2 13 10 9 0 1 10 9 1 9 2
35 15 13 0 10 9 15 13 0 7 13 0 2 3 13 10 9 1 9 16 13 0 7 10 9 15 8 1 10 9 0 9 7 10 9 2
20 16 13 10 9 2 10 9 0 16 13 10 9 8 13 1 10 9 0 0 2
22 1 12 10 11 11 1 11 2 11 13 10 9 1 11 2 11 1 10 11 1 11 2
30 3 2 1 10 9 13 0 13 10 9 1 10 9 1 10 9 2 1 10 9 0 13 1 10 9 1 10 12 9 2
10 10 9 1 11 2 11 4 13 9 2
19 10 9 3 0 3 15 13 2 7 3 15 13 1 10 9 1 10 9 2
35 10 11 3 13 9 2 7 10 9 2 10 0 9 11 11 2 13 1 10 9 1 9 1 12 2 15 16 13 1 11 1 10 0 11 2
11 1 9 2 13 10 0 9 1 10 9 2
15 16 10 9 13 9 7 9 2 3 15 13 9 7 9 2
51 1 10 9 2 16 10 9 13 0 2 15 3 13 10 9 1 10 9 0 16 13 2 16 2 16 4 13 2 3 3 1 9 0 1 10 12 1 12 4 13 16 11 4 1 13 10 9 1 10 9 2
60 9 1 10 9 16 13 1 9 2 10 9 13 1 9 0 11 11 7 10 9 11 11 13 13 3 2 16 10 9 1 9 13 10 12 9 2 1 10 0 7 15 13 1 10 9 1 10 9 0 7 10 9 1 9 1 9 1 12 9 2
44 10 9 0 16 13 9 1 10 9 1 0 9 13 1 10 9 1 9 1 9 4 13 16 15 13 3 9 7 2 3 2 15 13 1 13 9 15 4 4 13 3 1 9 2
42 10 9 13 1 10 9 16 1 9 1 16 11 2 11 13 3 7 10 9 1 13 10 9 2 10 11 13 1 10 9 2 1 10 10 9 10 9 0 1 9 2 2
21 15 15 13 1 9 1 10 8 1 13 1 10 11 1 13 10 9 7 10 9 2
47 13 0 13 16 10 9 13 10 9 1 11 7 11 7 1 10 9 12 0 9 1 9 4 1 13 10 9 1 15 1 10 9 7 15 13 1 10 0 9 13 1 10 0 9 1 11 2
28 1 10 9 1 10 9 11 13 13 16 10 9 4 13 1 1 9 2 1 10 9 1 16 13 0 1 15 2
30 3 2 13 10 9 16 13 1 11 1 9 1 10 9 11 11 2 15 13 10 9 1 9 1 10 9 1 11 11 2
21 1 10 9 1 9 10 9 4 13 0 2 1 9 13 1 9 2 0 9 2 8
32 13 1 10 9 16 2 1 12 2 13 1 9 1 10 9 1 10 9 11 10 9 2 1 10 9 1 9 1 10 9 0 2
21 11 11 13 10 9 13 1 9 1 13 9 7 9 1 10 9 1 9 0 11 2
8 3 13 16 13 13 10 9 2
7 13 1 10 9 1 12 2
33 1 9 2 10 9 0 13 10 0 9 0 8 2 0 1 10 9 0 8 1 10 9 0 2 1 1 10 9 7 8 5 12 2
14 13 1 10 9 1 11 1 10 11 11 1 10 11 2
18 1 12 13 10 0 9 2 1 10 9 11 2 3 13 1 11 11 2
73 10 9 2 1 10 9 1 10 11 11 1 11 2 15 4 13 2 1 10 9 2 3 1 10 9 1 10 11 11 1 11 1 11 1 11 1 10 9 2 10 9 1 10 9 1 9 1 10 11 11 2 2 13 3 1 11 7 13 1 10 11 1 11 1 9 1 10 9 0 1 10 11 2
31 1 9 1 9 10 9 1 11 13 10 11 1 10 11 2 11 1 9 13 12 7 1 9 13 12 13 1 9 1 9 2
29 15 13 9 1 10 9 10 9 2 16 13 1 9 0 10 9 1 11 1 10 11 2 11 7 11 2 1 15 2
14 1 10 9 0 2 13 9 1 10 9 11 7 11 2
18 11 2 9 0 2 9 1 10 9 1 11 2 1 9 2 11 2 2
19 3 13 10 9 0 1 11 2 11 2 7 10 9 1 11 2 11 2 2
11 11 4 13 1 10 9 3 0 1 11 2
39 2 11 13 10 9 1 9 0 16 13 3 0 1 13 1 10 9 1 9 2 9 0 7 10 3 9 1 10 9 0 1 10 9 2 2 13 11 11 2
27 11 2 12 2 2 9 1 9 1 9 1 10 11 11 7 11 2 11 7 11 1 10 9 1 10 9 2
49 3 16 10 9 1 9 1 10 9 1 10 9 1 9 0 13 1 10 9 1 10 9 1 9 0 1 9 1 10 9 2 3 3 4 10 9 13 10 9 3 16 13 10 9 16 13 10 9 2
5 13 1 10 9 2
7 10 9 13 0 1 15 2
39 13 13 10 9 1 12 9 2 1 15 16 13 1 10 9 0 2 7 10 9 1 10 9 15 13 16 16 13 9 1 10 9 4 7 13 10 12 9 2
32 9 1 11 2 13 10 11 11 11 11 7 11 1 10 9 2 3 10 9 0 0 3 0 1 10 9 1 10 12 1 11 2
33 3 4 13 15 3 1 4 13 1 9 2 1 16 13 1 10 9 3 2 3 10 9 0 2 3 0 7 3 0 2 1 9 2
12 10 10 9 13 1 11 11 1 3 15 13 2
21 13 9 1 10 2 11 11 11 2 11 11 2 2 7 9 1 10 11 1 11 2
34 10 9 0 2 10 9 1 9 2 10 9 7 10 9 1 10 11 2 12 13 10 9 13 1 11 11 1 10 9 1 11 2 11 2
33 1 13 1 10 9 7 1 10 10 9 1 10 12 2 13 1 10 0 9 1 9 1 10 11 11 2 13 10 9 1 11 11 2
15 1 10 9 13 10 9 16 3 15 13 1 10 9 13 2
56 1 10 9 2 10 9 4 13 1 10 9 1 10 9 0 2 9 2 10 0 9 2 12 9 2 9 2 9 1 9 2 9 0 2 0 9 2 1 10 9 2 3 7 10 9 1 9 1 9 1 9 7 9 1 9 2
11 10 9 1 11 15 13 0 1 10 9 2
35 13 1 10 9 1 12 0 9 2 13 2 10 9 13 1 15 15 13 1 9 2 7 11 2 10 9 13 1 15 15 13 1 9 2 2
38 1 10 9 1 11 1 10 11 1 11 2 10 9 3 4 13 1 10 9 2 4 13 1 0 1 9 1 10 9 12 1 10 9 0 1 11 11 2
20 10 9 16 13 1 11 13 13 15 1 9 13 1 10 9 1 10 9 0 2
26 1 10 9 12 10 9 13 9 1 0 9 2 1 15 15 15 13 1 10 11 1 11 1 10 9 2
6 15 13 13 10 9 2
23 11 11 11 13 15 1 10 9 3 9 1 10 9 1 10 9 1 10 11 2 11 11 2
12 1 12 13 10 9 1 10 9 1 0 9 2
25 3 2 13 12 9 0 2 1 15 2 10 0 11 2 2 13 1 11 11 7 13 1 11 11 2
46 3 4 13 1 10 0 9 1 12 2 12 7 12 2 13 3 10 0 9 1 11 2 1 12 9 1 10 12 9 1 11 7 15 1 3 12 9 1 13 12 9 1 10 0 9 2
31 10 9 1 9 16 13 1 10 9 13 10 9 1 9 16 15 13 3 0 1 10 9 7 15 13 10 9 0 3 3 2
11 11 11 2 8 2 13 10 9 9 0 2
34 1 10 9 1 9 1 3 2 13 10 0 9 16 13 15 1 11 7 16 2 3 2 15 13 7 13 1 10 0 9 1 10 11 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
64 10 9 1 10 11 0 4 13 10 9 1 10 9 7 4 13 16 13 10 9 0 2 3 7 2 1 15 2 10 9 2 2 11 11 2 2 13 1 9 1 10 9 2 11 2 13 9 1 9 1 9 1 13 10 9 1 11 2 7 3 13 1 15 2
19 10 9 11 13 10 9 13 1 13 10 9 2 13 3 10 9 3 0 2
26 1 9 1 10 9 1 10 9 0 2 4 1 13 10 9 2 13 10 9 1 10 0 9 1 9 2
13 13 1 10 9 10 0 9 2 8 7 13 9 2
43 9 7 9 0 1 11 13 16 10 9 13 10 9 1 9 1 10 9 2 1 0 1 10 9 1 9 0 1 10 11 7 11 2 1 15 15 13 9 16 13 10 9 2
40 10 11 11 11 11 11 13 10 9 1 10 9 1 11 3 1 10 0 2 9 2 7 10 9 1 10 9 1 11 1 10 9 7 10 9 2 1 9 2 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
38 10 11 11 1 11 11 2 11 2 13 1 9 1 11 12 0 9 0 1 9 0 1 10 11 2 11 11 1 10 11 11 2 1 11 2 11 2 2
34 1 9 1 10 9 15 13 10 9 1 9 1 9 7 0 2 3 1 10 11 1 9 3 15 13 9 1 10 9 1 10 9 2 2
18 3 15 13 1 12 9 2 8 2 1 13 1 12 9 2 8 2 2
25 10 9 12 9 1 11 11 2 11 13 10 9 1 12 9 13 1 10 0 9 11 11 2 11 2
12 1 12 4 13 1 10 9 0 1 10 9 2
5 10 12 13 0 2
4 13 1 11 2
27 10 0 9 7 11 1 10 11 13 1 10 0 9 1 11 2 3 4 13 1 10 0 9 1 13 11 2
35 1 9 0 1 10 9 1 11 15 13 10 9 0 1 9 1 10 9 2 7 13 0 10 9 1 10 9 1 10 10 9 0 1 9 2
30 3 13 13 16 11 13 9 0 2 7 3 4 7 13 3 13 10 9 0 2 16 13 1 15 1 10 9 3 0 2
32 3 4 13 10 12 1 11 1 12 2 13 16 10 9 13 13 1 10 9 0 2 15 13 1 13 1 10 9 7 4 13 2
28 10 9 13 1 10 12 9 16 13 11 16 13 1 11 2 10 9 2 9 7 0 16 13 10 9 16 13 2
11 10 11 15 13 10 9 1 10 0 9 2
24 3 3 2 16 10 12 9 13 9 0 2 11 7 11 15 13 10 9 3 0 1 10 9 2
51 1 9 0 1 10 9 0 13 10 11 2 9 1 9 16 15 13 1 9 1 9 2 9 2 9 7 9 0 2 10 9 2 10 10 9 1 9 0 1 9 0 16 15 13 1 0 9 1 0 9 2
40 10 9 4 13 1 10 10 9 1 9 2 13 1 12 9 0 2 1 10 2 11 11 11 2 1 10 0 9 1 10 2 11 11 2 2 10 9 3 0 2
15 15 13 2 1 10 9 0 1 10 9 0 1 10 9 2
12 11 13 10 9 1 9 0 1 10 9 11 2
35 13 10 9 1 9 7 3 3 13 1 10 11 2 13 3 7 15 13 1 10 0 9 15 3 13 1 13 9 1 10 11 11 1 9 2
10 15 13 1 10 0 9 3 1 9 2
17 1 13 10 0 9 1 9 16 13 1 10 9 15 13 9 11 2
48 3 13 1 10 9 11 2 10 11 11 7 10 11 11 2 2 1 10 9 11 2 11 7 11 2 2 1 10 9 11 2 11 7 10 11 11 2 7 1 10 9 11 2 11 2 8 9 2
22 11 13 1 9 1 10 9 10 12 1 11 1 12 2 13 1 10 9 1 10 9 2
9 3 15 15 13 13 1 10 9 2
30 10 9 1 9 0 1 11 1 10 11 2 13 1 10 9 1 10 9 1 11 11 2 13 10 9 0 1 9 0 2
11 3 1 13 1 10 9 0 13 1 9 2
83 10 9 13 1 10 9 7 1 10 9 1 10 9 0 11 7 11 11 13 1 10 11 3 13 10 0 9 2 13 11 11 11 2 11 11 11 2 11 11 7 11 11 11 7 1 10 9 1 9 13 10 0 9 1 10 9 2 11 11 2 16 13 13 1 0 10 9 1 10 9 1 10 9 2 13 1 10 9 0 1 10 9 2
27 10 9 1 11 13 12 9 0 2 10 12 1 11 2 13 1 10 9 11 11 1 10 9 1 11 11 2
25 10 9 13 10 9 1 10 12 15 13 11 2 13 15 1 11 2 12 2 7 11 2 12 2 2
19 1 10 0 9 2 10 9 0 4 13 1 11 2 7 3 0 1 11 2
16 10 0 9 13 1 10 9 0 11 11 3 13 9 1 11 2
8 1 10 9 4 13 10 9 2
34 1 9 1 10 9 1 12 2 11 4 13 10 9 1 10 9 1 10 11 7 15 4 13 1 10 11 11 11 10 9 1 10 9 2
16 11 2 0 9 1 10 9 2 3 13 10 9 1 9 0 2
9 0 1 15 13 13 11 1 9 2
20 10 3 0 2 9 3 0 13 15 16 13 16 10 9 7 10 9 15 13 2
15 10 9 0 15 13 1 10 9 1 10 0 1 12 9 2
28 10 9 0 11 13 10 9 16 3 15 13 15 7 10 9 13 1 10 9 2 1 15 15 3 15 13 3 2
36 1 10 9 3 13 10 9 1 9 15 13 2 1 10 9 1 12 10 9 2 0 1 11 1 9 11 11 11 2 1 10 9 1 11 11 2
19 11 13 13 2 1 13 16 10 9 4 13 1 10 0 9 13 1 11 2
18 10 9 1 11 13 0 9 1 9 16 13 16 10 9 13 3 0 2
22 11 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
20 13 1 10 9 7 13 15 8 13 15 7 15 2 16 15 13 9 7 9 2
25 15 13 1 10 9 13 15 3 7 10 2 9 1 10 9 2 2 3 13 16 13 10 9 11 2
19 1 9 2 10 9 13 16 13 0 13 7 13 10 9 1 11 10 11 2
17 10 9 11 11 4 13 1 3 12 9 2 12 9 2 1 9 2
16 1 13 15 2 15 13 7 15 13 16 15 13 3 1 3 2
14 1 10 9 1 12 2 13 12 9 13 1 11 11 2
49 1 10 11 11 1 10 9 15 13 10 9 3 0 1 9 1 0 9 2 8 9 7 9 2 16 13 10 9 1 10 9 0 1 11 0 2 10 9 0 7 0 13 10 0 9 1 10 9 2
22 3 15 13 10 9 13 1 10 9 0 1 9 1 9 16 3 13 13 1 0 9 2
9 15 13 10 9 1 11 1 12 2
37 3 3 1 10 9 1 10 9 0 2 11 4 13 10 9 1 12 9 2 12 1 10 9 0 7 9 8 7 12 1 10 9 0 7 9 8 2
14 16 13 2 3 13 10 9 1 10 9 0 1 11 2
18 10 9 13 4 1 13 2 3 2 10 9 1 9 1 9 1 9 2
32 10 9 2 13 1 10 9 1 9 11 2 13 10 9 1 13 3 2 13 10 9 0 1 11 2 11 7 10 9 1 11 2
13 13 0 1 10 9 2 1 9 1 9 0 0 2
23 9 1 10 9 0 11 11 2 13 1 10 9 0 9 1 10 9 0 1 10 9 12 2
11 10 9 1 10 9 1 10 9 13 0 2
33 1 10 9 2 1 15 1 9 1 9 0 2 10 9 1 10 9 1 9 0 7 0 13 10 9 0 1 10 9 1 10 9 2
11 10 11 1 11 13 10 0 9 1 9 2
28 7 13 16 3 1 10 9 10 9 1 10 11 1 10 9 11 13 1 10 9 0 1 13 10 9 2 0 2
25 3 1 10 9 1 11 1 10 11 3 13 10 9 0 7 0 1 10 9 7 10 9 1 11 2
7 11 3 13 13 15 9 2
26 10 9 0 16 15 13 13 1 1 12 5 9 1 9 2 7 10 9 3 1 12 5 9 1 9 2
21 9 1 10 9 1 10 9 0 2 2 12 2 13 10 9 3 0 1 10 9 2
14 1 9 1 9 15 13 1 10 9 0 7 0 9 2
68 10 9 1 9 4 13 15 10 9 0 1 10 9 0 2 16 13 3 1 12 9 0 1 13 9 1 9 3 13 2 1 9 13 10 9 3 0 7 1 13 0 1 13 9 1 10 9 1 10 9 2 7 1 9 1 15 15 13 1 10 9 7 15 13 1 10 9 2
12 15 13 1 12 9 2 11 2 11 7 11 2
67 10 11 11 1 11 1 10 9 12 7 11 11 11 1 11 1 10 9 12 13 10 9 0 16 1 10 9 15 4 13 1 9 1 11 1 9 1 10 9 0 13 1 10 9 0 1 10 9 1 11 11 2 11 7 13 9 1 10 11 11 11 7 1 10 11 11 2
18 10 9 0 1 10 9 13 0 2 4 1 13 15 3 1 10 9 2
13 11 13 1 11 11 1 16 11 4 13 10 9 2
9 15 13 16 15 13 1 10 9 2
34 2 3 9 2 16 4 7 13 3 10 9 1 16 10 11 2 13 11 2 13 10 9 1 10 9 16 1 12 9 4 13 10 9 2
34 10 9 1 11 11 1 9 1 10 9 12 13 15 1 10 9 1 10 9 2 13 1 13 10 9 1 15 9 7 9 1 11 11 2
24 13 10 9 2 10 0 9 2 1 10 15 3 13 2 10 9 2 1 9 2 11 7 11 2
15 7 1 3 13 9 0 2 1 10 0 9 1 13 15 2
34 10 9 13 10 9 13 2 9 2 7 2 9 0 2 7 13 3 1 13 1 10 9 0 16 2 3 2 13 10 9 1 10 9 2
21 15 13 10 9 7 15 13 1 9 2 3 13 15 7 13 0 10 9 1 9 2
37 10 9 15 13 1 9 1 11 13 1 9 0 3 13 1 10 9 1 2 11 11 11 11 2 2 13 9 1 9 15 3 0 7 10 0 9 2
30 3 2 10 9 15 13 1 10 0 9 7 1 12 13 1 3 1 12 9 2 1 15 15 13 0 13 10 9 0 2
23 3 1 11 11 13 9 1 10 9 1 9 13 10 11 1 10 15 3 13 9 11 11 2
12 9 13 1 10 9 2 12 1 11 1 12 2
24 13 1 10 9 1 10 9 1 10 11 1 11 1 3 3 12 9 1 9 1 11 1 12 2
22 7 10 9 0 15 4 13 1 10 9 0 2 1 10 9 11 2 11 7 10 11 2
18 10 9 3 4 13 1 9 16 13 10 9 1 9 1 10 9 0 2
21 10 9 3 13 15 9 16 10 11 11 13 11 1 10 11 2 11 11 11 2 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
24 13 1 10 11 11 11 11 10 9 1 11 2 12 2 7 9 2 12 2 3 13 10 9 2
42 1 12 13 1 10 9 1 11 0 7 3 13 1 15 1 11 11 1 11 11 7 11 11 2 7 1 11 1 11 11 11 11 2 9 1 10 15 13 1 0 9 2
25 1 10 9 13 10 9 0 2 13 1 10 3 9 7 9 1 9 13 1 10 9 9 2 9 2
12 1 9 15 13 1 9 16 13 1 1 11 2
14 10 10 9 3 15 13 1 10 11 8 11 11 12 2
25 1 12 13 10 9 0 7 1 12 13 1 10 9 10 9 1 9 1 10 11 1 11 1 12 2
18 11 13 9 1 10 11 1 11 1 13 1 10 11 11 1 10 9 2
29 10 9 11 4 4 13 1 9 0 1 11 2 11 2 11 11 2 11 11 2 11 2 11 11 2 11 7 11 2
17 13 13 1 11 2 3 13 12 9 2 3 1 9 1 10 9 2
42 3 15 4 1 13 1 13 15 13 7 3 13 2 7 3 15 13 1 9 2 1 9 2 1 9 7 3 1 9 2 13 3 4 1 13 1 10 13 1 10 13 2
11 13 9 1 10 9 1 10 9 0 11 2
67 13 13 1 10 9 16 4 1 13 1 10 11 11 1 10 11 7 1 0 1 10 9 2 15 4 13 1 10 9 1 10 9 7 1 9 13 1 10 9 1 7 15 13 1 10 9 8 10 9 15 13 1 10 9 7 13 10 10 9 7 9 1 15 16 15 13 2
40 10 9 13 0 16 15 13 1 9 1 9 13 1 9 2 1 9 2 9 9 8 7 9 1 0 9 1 9 2 1 9 2 9 1 10 9 11 11 2 2
31 15 15 13 1 10 9 11 11 2 15 15 13 1 9 7 13 2 1 15 15 9 1 10 9 1 11 13 10 9 0 2
13 10 9 1 9 13 1 12 8 2 2 5 12 2
41 10 9 0 13 13 12 9 13 1 10 9 1 11 2 10 0 1 15 13 1 10 11 11 2 9 1 10 9 2 11 2 2 3 7 10 0 9 1 10 9 2
42 11 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 11 2 7 10 0 11 1 11 15 13 7 13 2 13 1 11 0 7 13 1 10 9 1 15 2
19 10 9 13 1 9 10 9 0 2 10 9 1 9 7 10 9 1 9 2
17 10 9 13 10 9 1 10 9 1 11 2 1 10 9 1 11 2
17 10 11 11 11 15 13 3 1 10 9 1 11 11 1 10 9 2
14 10 9 3 15 13 1 10 9 1 11 7 10 9 2
9 1 9 2 13 9 0 1 11 2
16 10 9 1 10 9 13 10 9 1 9 1 10 12 9 0 2
17 13 10 9 0 0 2 8 2 2 16 3 13 1 10 9 0 2
26 13 10 9 1 10 9 2 3 16 15 13 1 10 9 1 10 9 15 13 10 0 9 1 10 9 2
94 1 10 9 2 10 11 4 13 1 9 0 7 0 1 10 9 1 9 1 8 8 2 7 10 9 0 1 9 1 10 9 2 10 9 0 7 10 9 0 2 13 10 9 0 0 2 15 16 13 16 1 10 0 9 1 9 2 10 0 9 1 10 9 15 13 0 2 7 16 10 0 9 0 15 13 1 9 3 0 2 0 1 12 9 1 9 1 10 9 1 10 3 0 2
50 13 3 1 10 9 0 1 10 9 3 13 10 15 7 3 1 10 9 3 0 1 15 2 11 13 10 9 0 7 13 10 9 0 0 1 10 9 1 10 9 1 10 9 7 15 15 13 1 3 2
9 15 13 13 1 10 9 3 0 2
49 11 11 13 3 16 3 13 2 1 12 13 10 9 1 9 1 11 11 7 15 8 1 13 10 9 1 10 9 1 10 15 15 4 4 13 10 9 7 15 13 16 13 3 0 2 0 7 0 2
64 10 9 1 11 2 10 9 7 10 0 9 1 10 9 1 9 7 1 9 3 1 11 2 11 2 11 2 11 2 11 2 13 1 10 9 0 1 11 11 1 9 1 10 0 9 1 9 1 13 15 1 10 9 1 13 1 10 9 1 10 9 0 3 2
32 1 9 1 10 0 9 2 4 1 4 13 1 10 0 9 1 11 11 2 15 16 2 3 2 13 1 16 4 1 13 9 2
26 1 10 9 0 2 10 9 1 9 1 9 15 4 13 1 9 1 10 9 1 10 9 0 7 0 2
46 13 1 10 9 1 10 16 15 13 2 13 2 2 10 9 1 10 9 4 13 0 1 10 12 7 12 9 7 3 13 10 0 13 2 3 4 1 13 10 0 9 1 10 9 2 2
56 11 8 10 9 0 13 1 11 11 11 1 10 0 9 13 1 9 1 11 11 11 1 10 9 0 1 11 11 16 15 13 10 12 1 11 1 12 7 16 13 1 9 1 11 11 2 11 1 11 2 11 11 7 11 11 2
20 10 9 2 3 1 0 2 0 7 0 2 13 9 0 3 1 10 9 3 2
37 1 4 13 10 9 1 10 9 2 11 13 1 11 2 13 16 11 15 13 7 15 13 16 13 13 15 2 7 13 1 10 9 15 3 15 13 2
12 10 9 13 0 9 2 13 13 1 10 9 2
37 1 12 13 3 9 1 10 9 0 1 10 9 0 1 11 2 16 13 3 1 10 9 1 9 11 7 13 1 12 1 10 9 1 10 9 12 2
37 10 9 0 13 1 10 11 11 1 10 9 11 11 13 10 12 1 11 1 12 2 16 15 13 10 9 2 13 15 3 9 7 10 9 1 9 2
39 10 9 0 2 10 9 2 10 9 0 2 10 9 2 10 9 0 7 10 9 2 1 10 15 4 7 13 10 11 2 10 9 7 10 9 1 10 9 2
30 10 9 13 1 3 9 13 1 10 9 8 1 10 9 7 13 9 1 10 9 1 10 8 2 8 2 1 10 9 2
26 11 1 11 11 2 12 2 2 10 0 0 9 1 9 2 4 13 10 9 1 9 7 10 9 0 2
34 9 1 10 9 10 9 13 10 9 0 1 10 0 9 2 7 1 10 0 9 4 7 13 16 13 10 9 1 10 3 0 0 9 2
27 13 10 9 1 10 9 0 1 10 9 11 2 13 3 1 11 2 3 9 3 4 13 10 9 11 11 2
16 10 9 4 13 1 10 9 1 11 11 2 1 12 7 12 2
17 13 10 9 1 9 7 1 9 0 7 13 1 10 9 1 9 2
23 15 13 1 10 11 1 11 2 10 11 1 11 11 7 1 11 7 1 10 11 1 11 2
18 10 9 1 9 10 15 0 2 13 1 9 10 9 3 13 3 0 2
28 10 9 0 13 10 9 1 12 5 1 10 11 1 11 11 2 13 1 10 9 0 1 10 11 11 1 11 2
40 10 9 1 10 11 11 13 13 1 11 1 10 9 1 10 9 1 11 2 11 7 11 2 16 11 13 15 2 7 13 1 10 9 0 1 10 9 1 9 2
24 1 12 2 15 13 11 1 9 1 10 9 2 11 11 1 11 2 9 2 11 11 2 2 2
7 1 12 13 10 11 11 2
18 3 15 13 1 13 10 9 1 11 2 10 9 0 7 10 9 8 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
33 10 9 3 0 13 1 10 9 1 11 2 1 15 10 8 11 11 15 13 10 9 0 2 2 7 11 11 13 1 10 11 11 2
55 1 11 2 11 13 10 9 1 10 9 16 13 10 0 9 1 13 10 9 1 9 1 9 1 10 12 1 10 12 0 9 1 9 1 11 2 15 16 16 13 2 15 13 1 10 9 1 10 12 5 1 9 1 12 2
25 11 11 11 2 11 1 10 11 2 9 1 11 2 12 2 2 9 0 2 0 1 10 11 0 2
11 4 13 1 11 11 13 1 10 0 9 2
17 10 9 0 15 13 0 7 0 9 0 1 10 13 1 10 9 2
48 10 11 11 1 11 11 13 10 9 0 1 10 9 1 10 9 0 13 1 10 9 1 11 11 2 3 3 1 10 9 9 1 10 9 2 1 10 9 1 10 11 8 2 12 2 11 2 2
20 10 9 0 4 13 1 10 9 11 11 1 10 9 0 11 2 11 7 11 2
15 15 13 3 1 9 0 2 7 15 13 7 13 1 9 2
33 13 9 1 9 1 10 9 0 13 9 2 9 2 9 2 9 7 9 0 2 7 13 10 3 0 7 1 9 0 1 10 9 2
23 1 9 1 10 9 2 10 9 11 13 4 1 13 15 7 13 15 1 9 1 10 9 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
49 4 13 10 9 1 15 11 13 9 1 9 0 1 9 3 1 10 11 11 1 10 11 2 11 2 1 10 9 1 1 11 7 10 11 1 11 1 10 9 1 10 11 1 1 11 2 11 11 2
20 10 9 0 15 13 13 1 10 0 9 1 9 2 1 15 15 15 13 0 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
13 1 9 1 12 15 13 10 0 9 0 1 11 2
33 15 13 16 1 10 9 15 13 10 12 5 1 10 9 1 9 0 1 11 7 15 13 10 9 0 1 10 12 5 1 10 9 2
33 3 13 9 1 10 11 11 2 10 9 1 9 1 11 2 1 3 13 9 1 11 11 11 2 11 11 2 11 11 7 11 11 2
26 3 1 13 10 9 0 2 10 9 15 13 2 1 9 1 9 2 1 9 1 10 9 7 10 9 2
30 10 9 15 13 1 11 1 12 2 13 15 10 9 0 12 16 13 10 9 0 2 10 12 1 11 1 10 0 9 2
21 13 10 9 0 1 9 1 10 9 16 13 10 9 1 9 1 9 3 3 13 2
21 10 8 1 10 9 0 2 3 1 10 12 5 2 4 1 13 1 10 12 5 2
23 13 1 10 9 2 11 13 13 7 13 10 9 2 13 12 9 1 15 9 1 12 9 2
33 1 10 9 0 15 13 10 9 0 1 10 15 13 9 7 9 1 10 15 13 10 9 1 10 0 9 16 15 13 1 10 9 2
22 13 1 10 9 7 10 9 0 1 10 11 11 11 2 4 13 1 10 11 1 11 2
65 4 13 10 9 1 10 15 3 13 13 9 2 11 13 13 15 1 10 9 1 10 9 2 1 10 13 1 11 4 13 1 10 9 1 10 9 1 10 9 2 11 11 2 15 3 15 13 1 10 9 16 15 13 1 11 2 10 9 16 15 13 1 10 9 2
49 1 10 9 10 9 1 10 11 1 10 11 11 13 16 10 9 0 2 0 7 0 3 13 0 3 7 3 13 0 1 13 9 7 13 1 15 3 2 0 16 15 13 3 0 1 13 10 9 2
18 10 9 13 1 10 9 5 12 1 10 9 0 2 1 9 1 12 2
25 10 15 13 1 10 9 1 9 11 2 16 1 10 9 15 13 1 10 9 1 10 9 1 11 2
19 11 11 11 2 13 10 12 1 11 1 12 2 11 2 13 10 9 0 2
32 1 10 9 2 10 9 1 10 15 10 9 1 10 11 15 13 1 10 9 1 11 13 16 10 11 15 13 3 3 1 11 2
8 1 10 9 4 13 15 9 2
25 15 15 13 1 9 0 2 9 2 2 9 0 2 9 1 9 0 2 9 2 9 7 0 11 2
22 13 0 7 10 9 13 10 9 1 10 9 0 2 10 15 15 13 3 1 10 9 2
20 1 10 9 0 1 10 11 11 0 2 10 9 0 4 13 7 13 1 11 2
47 10 10 9 3 13 3 2 15 1 13 15 1 10 9 0 1 10 9 1 11 2 9 11 2 16 13 7 13 10 9 2 3 10 9 7 9 0 1 10 2 9 2 13 1 9 0 2
17 9 1 9 2 9 2 15 13 0 9 1 10 0 9 1 9 2
23 1 9 1 11 2 10 9 0 13 1 11 11 13 1 12 9 2 12 9 7 12 9 2
22 10 9 3 0 13 10 9 1 9 1 10 9 0 1 11 12 1 10 9 1 11 2
16 1 10 9 11 13 3 2 13 10 0 9 1 10 9 2 2
18 12 8 12 9 2 0 2 3 0 2 3 0 2 3 0 2 0 2
25 10 9 1 11 4 13 1 9 1 10 9 2 16 13 10 9 0 1 9 1 10 9 1 11 2
60 11 13 1 12 9 1 10 8 11 2 4 13 1 10 9 1 10 9 0 2 1 15 10 11 1 11 2 16 13 1 3 1 10 9 11 11 2 13 1 10 9 11 2 10 9 1 11 11 7 10 8 11 3 13 10 9 1 10 9 2
36 10 9 11 2 10 9 0 13 11 11 1 11 11 1 11 2 13 10 0 9 0 1 9 0 0 1 15 15 3 13 10 9 1 11 11 2
8 8 9 10 0 9 1 11 2
33 1 10 9 2 11 15 4 13 1 10 9 0 1 11 2 13 10 11 1 11 7 10 9 1 10 9 1 13 3 1 12 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
17 10 9 15 13 1 10 11 11 16 13 10 9 7 10 9 0 2
14 15 13 1 11 2 11 2 11 7 11 2 7 11 2
60 1 10 9 2 10 9 1 9 2 11 11 2 13 10 0 9 1 3 1 12 9 2 1 10 9 1 10 9 1 8 9 1 10 9 2 7 13 16 10 9 0 3 1 10 9 0 13 2 13 10 10 9 0 1 7 15 15 13 2 2
48 10 9 4 13 2 7 1 9 1 9 2 11 11 13 1 10 11 11 11 2 13 15 3 1 10 0 8 1 11 11 1 13 1 10 9 7 1 10 9 13 12 9 1 12 9 1 9 2
63 1 0 2 3 1 12 12 9 0 1 3 1 12 9 1 15 9 1 10 9 15 13 1 9 2 16 10 11 1 11 11 13 1 10 9 0 1 10 11 12 1 11 1 10 15 15 13 10 11 2 10 11 1 11 7 10 11 11 1 14 2 9 2
22 10 9 1 11 13 10 9 0 1 10 9 0 3 0 1 11 2 13 1 12 2 2
15 11 7 10 9 15 13 13 1 10 9 0 7 3 0 2
30 1 9 4 13 3 1 10 0 9 1 9 7 1 10 13 15 1 10 0 9 1 10 11 11 2 13 3 10 9 2
12 10 9 1 10 9 13 1 10 9 11 11 2
28 15 15 13 13 3 1 10 9 2 16 1 10 11 11 15 13 10 9 1 9 1 9 3 0 1 10 9 2
21 10 9 15 13 1 11 11 2 9 0 9 7 9 0 2 7 15 13 1 11 2
11 11 15 13 1 10 9 1 11 7 11 2
28 10 9 13 1 9 0 1 10 9 0 7 0 1 9 1 9 0 2 9 1 9 7 9 0 1 10 9 2
101 1 10 9 1 10 15 4 13 13 11 2 10 11 2 12 2 2 10 9 1 10 9 2 12 2 2 1 11 11 2 11 2 12 2 2 1 11 2 11 11 2 12 2 2 1 11 2 11 2 11 1 11 2 12 2 2 1 11 11 2 10 9 1 11 2 12 2 2 1 11 11 2 11 11 7 10 11 1 10 11 2 12 2 2 1 10 9 1 11 7 10 11 2 12 2 2 1 11 11 11 2
66 1 12 2 1 9 1 10 11 1 11 1 11 11 11 2 13 9 1 11 1 10 9 1 10 9 1 10 9 0 1 11 11 2 11 2 1 9 1 9 0 2 9 1 9 2 9 0 1 13 10 9 11 2 7 9 1 9 1 10 9 7 9 1 10 9 2
16 10 11 11 11 2 11 11 2 11 11 11 2 8 12 2 2
17 10 0 9 0 13 1 10 9 1 10 3 13 11 2 1 12 2
29 10 12 1 11 2 1 11 1 10 11 2 13 15 0 2 15 16 13 1 10 9 0 7 10 9 1 12 9 2
10 0 2 0 7 15 3 9 0 13 2
28 1 10 9 3 10 9 0 11 7 10 9 1 15 3 13 2 4 13 3 9 1 9 0 1 10 9 0 2
43 10 9 1 9 7 10 9 13 12 9 1 9 16 13 1 10 0 9 2 1 10 9 1 9 13 10 9 1 10 9 16 15 13 10 9 1 10 9 7 16 13 13 2
10 10 9 1 9 1 9 13 1 9 2
10 11 13 0 10 9 1 10 0 9 2
13 2 11 11 11 11 12 13 10 0 9 1 15 2
15 1 10 9 12 13 1 10 9 1 12 9 2 11 2 2
31 3 2 15 13 10 9 1 9 0 1 10 9 8 1 9 13 0 1 10 9 0 2 7 15 13 3 1 13 15 9 2
70 7 15 1 10 9 0 3 0 13 10 9 11 11 11 2 15 1 12 13 2 10 11 11 13 1 10 9 1 11 2 10 15 13 1 16 10 9 0 2 12 2 10 9 0 0 13 1 10 9 0 1 9 2 1 10 9 1 0 1 12 9 1 9 13 1 9 1 9 0 2
24 16 13 10 9 1 10 9 2 13 9 0 1 10 9 7 1 10 13 10 9 13 1 11 2
23 0 1 10 11 11 1 11 1 12 2 15 0 13 1 10 9 1 10 9 0 1 11 2
9 11 11 15 13 13 1 10 9 2
21 10 9 1 11 13 11 1 11 2 13 1 11 1 10 9 1 11 2 1 11 2
10 4 1 4 13 1 10 11 1 11 2
28 11 1 11 2 11 2 3 1 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 9 0 0 2
36 10 9 13 10 9 1 9 1 9 2 13 1 9 1 10 9 2 9 2 9 2 9 1 9 2 7 9 1 9 0 1 11 11 1 11 2
32 3 1 15 10 9 13 2 7 1 9 1 10 9 8 10 9 0 4 1 13 9 1 10 9 0 16 13 10 9 1 11 2
4 10 9 13 2
33 15 1 10 9 13 10 9 0 2 7 10 15 15 13 1 10 9 1 10 9 0 1 10 9 1 10 9 1 10 9 1 9 2
92 10 12 1 11 1 12 9 1 9 1 10 9 7 9 7 1 10 9 0 1 13 1 15 16 3 13 13 7 13 2 13 1 11 13 15 1 10 10 9 1 11 2 13 1 10 3 0 9 7 13 15 10 9 1 10 15 16 2 1 10 7 10 9 2 15 13 1 13 10 9 15 15 13 2 16 13 10 9 1 10 9 16 13 10 9 2 13 10 9 1 9 2
13 10 9 1 9 13 1 12 13 2 2 5 5 2
15 10 9 3 0 13 10 9 2 13 1 10 9 11 11 2
30 13 1 10 9 1 10 9 1 10 9 1 10 9 0 1 10 9 7 9 1 10 9 0 2 9 15 13 1 12 2
66 1 15 9 1 10 9 1 9 1 10 2 11 1 10 9 2 2 1 9 3 13 10 2 11 2 2 1 10 0 9 1 9 1 10 0 9 16 15 13 1 10 10 9 2 1 13 10 9 2 10 9 7 10 9 2 3 15 4 13 1 10 9 1 10 9 2
18 1 10 9 13 3 1 12 9 1 10 0 9 1 9 1 10 9 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 13 1 9 0 7 2 12 5 2 12 5 5 13 9 2
20 10 9 4 13 1 10 9 11 11 2 16 3 13 10 9 0 1 10 9 2
23 9 7 9 15 13 1 10 0 9 11 2 3 1 9 3 13 1 10 0 9 1 11 2
31 1 9 1 16 10 9 1 11 13 10 3 0 1 10 11 11 10 9 1 10 9 13 3 7 3 0 1 10 10 9 2
43 16 4 13 11 2 10 9 0 1 9 0 2 10 9 1 9 0 4 13 1 9 1 10 3 1 12 9 1 10 9 0 10 9 1 11 2 11 16 13 13 12 9 2
14 10 9 0 4 13 9 1 9 9 1 10 9 0 2
20 0 1 12 9 1 9 2 11 13 1 10 11 11 11 11 1 11 2 11 2
26 3 1 10 9 1 11 2 11 1 11 11 15 11 2 13 1 13 9 1 9 1 10 9 1 9 2
19 10 12 1 11 1 12 12 9 13 16 10 9 0 13 1 10 9 11 2
40 10 9 13 1 10 9 1 13 10 9 0 1 10 13 11 11 2 3 1 0 9 2 10 9 0 13 1 10 9 1 10 11 1 10 9 0 1 10 11 2
31 11 13 15 1 10 10 9 16 13 1 11 2 15 0 2 16 15 13 1 10 9 1 10 9 0 1 10 9 1 9 2
21 10 9 1 9 13 13 1 11 1 10 9 1 0 9 1 9 1 13 10 9 2
27 11 11 2 1 9 2 9 0 0 2 11 8 2 13 10 9 1 9 0 13 1 10 0 9 1 11 2
11 13 10 9 1 9 8 7 10 9 8 2
37 11 11 13 10 9 0 3 2 16 13 10 9 1 9 0 7 13 10 9 1 10 0 9 1 10 9 1 11 1 9 1 10 9 10 9 0 2
28 1 9 1 10 9 2 10 9 13 1 11 2 11 2 7 13 1 11 1 10 13 10 0 11 11 1 12 2
40 15 13 3 1 10 9 16 15 4 13 1 9 1 10 0 9 1 10 9 1 10 11 7 10 11 7 3 1 10 9 7 9 1 10 9 15 15 15 13 2
44 10 9 15 13 3 0 16 15 13 16 10 9 3 13 10 9 4 13 11 2 11 7 11 2 7 16 13 10 9 1 9 16 8 10 9 0 1 12 9 1 10 9 0 2
33 1 10 9 1 10 11 1 10 11 2 3 4 13 10 9 1 12 7 12 9 2 15 13 10 12 9 1 9 7 10 12 9 2
8 10 9 0 4 13 1 11 2
8 10 0 9 15 13 10 11 2
9 13 9 1 10 9 0 11 11 2
14 1 10 9 3 1 11 13 15 10 9 0 11 11 2
14 15 13 0 1 13 15 1 10 9 0 1 10 12 2
29 4 13 10 12 1 11 1 12 1 9 1 10 9 1 11 11 7 13 10 9 1 10 9 1 10 9 11 11 2
14 10 0 9 1 9 15 13 1 10 9 1 13 11 2
32 10 9 11 15 13 1 11 2 11 16 11 13 12 9 7 13 1 10 9 3 11 13 1 10 0 9 2 10 11 11 11 2
24 9 1 10 9 2 7 3 10 9 2 13 16 13 9 1 10 9 1 9 1 10 11 0 2
39 1 10 9 1 11 2 10 9 16 15 4 13 1 10 9 1 9 4 4 13 2 3 13 2 1 9 2 2 2 16 13 9 0 7 1 10 0 9 2
25 4 13 10 12 1 11 1 12 1 13 10 9 1 11 7 11 16 3 4 4 13 1 10 9 2
33 7 1 13 13 1 10 0 9 2 11 15 13 10 9 1 10 9 2 15 15 13 1 15 7 13 10 9 1 13 15 10 9 2
46 10 9 1 10 9 0 1 11 1 9 1 11 2 11 2 4 13 10 9 1 10 9 1 10 9 1 10 9 1 10 16 4 13 0 1 13 15 1 10 9 1 10 9 16 13 2
58 11 11 13 3 10 9 1 10 9 0 11 11 16 13 1 10 0 9 2 7 3 2 3 4 13 15 1 13 3 16 10 11 11 13 3 1 12 9 7 3 2 9 13 1 9 1 13 1 10 9 13 1 10 9 1 10 11 2
24 10 11 1 11 13 9 1 9 13 1 11 11 1 10 12 7 12 2 7 3 15 4 13 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
36 11 13 10 9 0 1 10 9 1 11 11 2 15 13 3 1 10 11 11 7 9 1 11 11 2 10 2 11 2 1 3 1 12 12 9 2
39 10 9 13 15 1 10 9 3 13 1 10 9 0 1 10 11 11 2 7 15 4 13 9 1 9 0 7 9 2 11 11 2 7 9 2 11 11 2 2
18 15 13 1 10 13 15 10 12 9 1 10 9 1 10 9 0 11 2
42 10 9 1 10 9 1 10 9 7 10 11 11 13 16 1 10 9 0 15 13 10 9 13 1 10 0 9 13 1 10 9 0 2 10 0 9 1 10 15 13 0 2
29 13 9 1 10 9 1 11 1 10 9 12 7 3 13 1 11 11 1 10 9 1 11 15 11 13 12 1 12 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
53 10 9 13 1 11 2 9 1 11 2 3 13 13 1 10 9 1 10 11 1 11 11 13 3 10 9 1 10 9 0 1 11 11 2 9 3 9 1 10 9 0 1 10 9 9 1 10 11 1 0 12 9 2
32 1 3 0 2 11 13 16 13 9 1 13 2 3 1 10 9 1 10 9 1 10 9 1 11 2 1 10 9 11 7 11 2
16 10 9 13 10 9 0 13 10 9 1 9 0 1 10 9 2
5 13 0 1 11 2
30 10 9 1 11 7 9 13 0 1 10 9 1 10 9 1 15 15 13 10 9 0 11 1 10 9 0 1 10 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
31 10 9 0 15 13 1 9 3 0 1 2 9 2 9 2 9 2 9 2 9 0 2 9 2 9 2 9 0 7 9 2
7 3 4 13 2 1 3 2
12 10 10 9 13 1 9 1 3 1 12 9 2
6 1 0 2 12 9 2
6 3 3 0 1 9 2
20 11 11 11 2 3 13 1 11 11 11 2 13 10 9 0 1 11 2 11 2
23 13 9 1 10 11 1 11 1 10 11 1 10 11 7 1 10 11 11 1 11 11 11 2
38 3 2 13 16 10 9 13 3 0 1 10 13 2 1 9 1 10 11 1 9 2 10 9 1 10 9 1 9 0 13 7 3 13 10 9 1 9 2
30 3 2 11 13 1 10 9 1 11 1 12 1 10 9 1 12 9 2 15 15 4 13 1 9 1 9 1 10 9 2
23 1 15 1 10 9 4 7 13 15 3 13 9 0 7 13 15 3 1 10 9 1 11 2
17 10 9 8 13 10 0 9 8 2 7 1 9 3 0 7 0 2
28 10 9 1 11 1 10 11 2 3 13 3 0 2 7 3 15 13 1 15 1 10 9 1 10 9 1 11 2
30 10 9 7 9 1 11 2 13 1 9 10 12 1 11 1 12 2 13 10 0 9 1 9 1 10 9 1 10 11 2
32 10 9 0 1 10 11 11 13 10 9 1 12 9 11 2 7 10 9 4 13 1 10 11 1 11 7 11 1 11 1 12 2
7 15 13 10 9 1 9 2
10 10 9 1 0 9 0 13 11 11 2
16 13 1 10 11 1 10 11 1 10 9 1 11 11 1 11 2
46 10 9 13 10 9 1 10 9 2 3 13 1 10 9 1 10 9 11 11 2 11 13 10 0 9 2 11 13 1 11 1 13 15 10 9 1 11 2 11 13 10 9 1 11 11 2
17 1 10 9 1 9 2 11 13 13 3 10 0 9 13 1 9 2
16 15 13 1 10 9 1 11 3 1 10 9 1 10 11 11 2
34 10 9 1 10 15 15 13 10 9 13 12 9 2 15 4 13 1 10 9 7 9 1 10 9 1 9 13 1 10 9 1 10 9 2
11 13 10 9 1 13 10 11 1 11 11 2
72 16 1 15 15 13 15 2 1 3 7 13 10 9 0 2 13 1 13 1 10 9 1 15 1 10 9 16 13 1 9 1 10 0 9 0 7 16 2 1 9 2 15 13 1 10 9 1 10 9 1 10 9 0 7 10 9 1 10 11 11 9 2 12 9 0 10 9 1 13 10 9 2
19 11 13 10 9 7 13 10 9 1 12 9 2 13 3 1 10 9 0 2
28 10 9 3 1 13 9 1 9 12 7 9 12 1 12 12 9 3 1 13 15 1 10 9 1 10 9 12 2
34 1 13 10 11 2 1 12 13 10 9 0 1 10 9 1 11 2 4 10 3 13 7 13 1 9 1 10 9 1 10 11 1 12 2
35 10 2 9 2 1 10 9 13 4 13 1 10 9 1 11 11 7 11 11 2 1 10 11 11 11 8 11 1 10 11 11 1 11 11 2
4 13 1 11 2
21 15 13 1 10 9 3 0 2 10 9 0 7 0 2 7 10 9 1 10 9 2
26 13 1 15 10 9 13 13 16 13 1 10 9 0 1 9 1 10 9 1 11 10 9 13 10 9 2
9 11 13 10 9 1 10 9 12 2
24 10 9 13 1 10 9 1 11 11 2 3 15 13 9 2 16 13 1 10 9 1 10 9 2
18 13 10 9 0 7 1 9 0 16 13 1 12 7 12 9 1 9 2
7 10 9 10 9 13 0 2
38 10 9 0 1 10 9 2 11 11 2 15 13 1 10 9 0 11 11 2 15 15 13 0 1 10 9 1 9 1 10 9 1 10 12 1 10 12 2
52 10 9 0 13 10 9 16 3 13 10 9 1 10 9 10 12 9 16 10 9 11 11 2 16 15 13 1 3 12 9 1 10 9 2 13 10 9 16 13 10 9 1 9 7 9 16 15 13 10 12 9 2
38 11 3 13 1 12 1 12 1 11 1 10 9 0 1 10 0 9 2 7 1 10 9 13 11 11 2 10 0 9 1 9 1 10 11 11 2 11 2
40 1 10 9 3 13 1 9 0 2 3 13 10 9 1 10 9 2 11 1 10 11 2 11 13 10 9 2 11 9 1 10 9 2 2 3 1 11 11 11 2
32 3 2 1 10 9 1 10 9 2 10 9 1 11 13 10 9 1 9 16 15 13 1 10 9 13 7 13 10 9 3 0 2
23 13 1 9 1 0 9 1 11 11 1 11 7 13 9 0 1 11 12 1 10 9 0 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
19 1 10 0 9 2 11 15 13 1 10 9 1 10 9 3 0 1 11 2
8 1 10 9 0 13 3 0 2
73 1 10 9 13 1 10 0 11 11 2 7 1 10 16 13 10 0 8 2 11 11 2 7 10 0 9 2 11 11 2 11 8 8 11 1 12 2 2 10 9 13 10 0 9 0 1 10 9 1 10 9 1 10 0 9 0 2 3 9 0 1 9 2 7 10 9 1 10 9 1 10 9 2
13 3 13 3 15 13 10 9 1 10 3 0 9 2
11 1 12 15 13 1 10 9 11 11 11 2
21 11 11 1 11 13 10 9 7 9 1 10 11 11 1 10 9 1 11 2 11 2
65 1 15 11 15 4 13 9 1 11 11 2 11 2 11 7 11 11 2 7 3 4 13 0 9 1 10 9 2 3 1 10 11 10 11 2 11 10 11 7 3 10 12 9 0 16 15 13 3 1 10 9 11 1 11 2 3 1 10 9 11 11 7 10 11 2
27 10 9 1 9 0 11 11 2 16 13 10 9 1 10 9 0 2 13 3 1 13 9 1 10 9 0 2
22 10 9 3 3 13 1 10 9 2 16 15 13 16 13 10 9 1 12 5 3 9 2
27 11 13 3 10 0 9 0 1 10 9 2 7 11 10 9 0 9 1 10 9 1 10 9 1 10 9 2
20 13 1 10 9 11 11 1 12 2 11 11 1 12 7 10 11 11 1 12 2
21 1 9 2 12 13 9 0 7 10 9 13 1 9 0 2 11 2 11 12 2 2
17 7 11 3 13 9 7 9 1 13 10 9 0 1 10 9 0 2
34 15 13 16 10 0 9 1 9 1 10 9 1 10 9 16 3 15 13 16 13 9 2 4 13 1 10 0 9 0 1 10 9 0 2
18 15 13 10 9 1 7 15 13 3 7 3 15 13 1 9 1 9 2
44 16 11 11 2 1 9 2 13 13 3 1 10 9 12 9 13 1 9 1 9 13 1 12 12 9 2 15 13 1 16 15 13 10 9 16 13 3 1 10 9 10 10 9 2
9 13 3 9 4 13 1 10 9 2
31 11 11 15 11 11 11 11 2 12 2 2 4 13 1 15 1 10 9 2 15 16 13 10 9 1 10 11 1 10 11 2
28 1 10 9 1 10 11 11 1 12 2 10 9 4 1 13 10 9 1 10 9 1 10 9 0 1 10 11 2
24 11 11 2 16 13 1 11 2 13 10 9 2 7 11 2 10 9 2 15 13 13 1 9 2
60 13 16 1 10 9 0 2 3 13 1 11 2 15 13 10 9 16 3 13 10 9 2 9 2 9 2 9 7 9 2 7 13 16 10 10 9 16 13 9 1 9 2 9 2 9 2 9 7 9 2 1 15 2 4 13 9 1 0 9 2
30 9 1 10 9 0 2 10 9 1 9 0 1 10 11 11 2 2 15 2 2 2 13 15 1 10 9 0 3 0 2
20 7 3 13 3 2 10 0 9 1 10 11 1 10 11 2 13 10 9 0 2
3 11 11 11
24 13 12 9 0 1 10 9 1 9 2 10 0 2 10 14 2 0 2 10 0 7 10 0 2
30 10 9 13 0 1 10 13 10 0 9 1 10 9 11 0 13 15 1 10 0 9 1 10 11 2 1 10 11 0 2
25 10 9 1 11 2 11 16 13 10 0 9 13 11 2 9 7 11 1 10 9 0 1 10 9 2
33 1 0 13 9 7 9 1 10 9 2 1 15 15 10 9 15 13 1 10 9 0 1 9 11 11 2 1 10 12 9 1 9 2
20 10 9 13 10 9 1 10 9 11 7 1 15 15 2 13 3 0 1 9 2
24 1 9 2 13 16 15 13 2 3 3 2 1 10 9 1 11 2 2 11 7 10 9 2 2
40 9 0 1 11 7 9 0 1 10 11 15 13 1 10 9 1 9 13 1 10 9 1 2 10 11 2 2 1 10 9 1 11 1 11 2 1 12 7 12 2
28 10 9 0 13 13 0 2 15 15 13 1 10 9 1 10 9 13 1 10 9 0 7 10 9 1 12 9 2
19 10 9 1 9 1 10 9 4 13 3 1 10 12 1 11 1 10 12 2
29 3 1 13 1 11 1 10 9 1 10 8 2 13 9 1 10 9 3 15 13 10 9 1 10 9 1 10 9 2
8 10 9 13 13 1 12 9 2
19 1 10 9 4 13 1 10 9 0 2 13 3 1 10 9 1 11 11 2
21 10 9 15 13 3 1 10 9 7 10 9 13 1 9 1 10 9 1 12 9 2
75 13 1 10 2 9 1 9 3 0 7 0 10 9 4 13 1 10 9 0 1 10 0 9 1 9 1 9 7 9 1 10 9 1 9 2 16 7 3 13 1 0 9 1 0 9 1 10 9 1 9 2 2 2 11 13 11 2 13 1 10 9 0 1 9 2 2 11 11 2 2 1 11 11 2 2
28 4 13 1 10 9 12 5 12 8 9 9 7 12 5 12 2 9 9 2 7 9 1 10 9 1 12 8 2
32 11 15 13 1 10 9 2 7 1 10 0 9 1 11 1 10 9 2 3 2 13 1 10 9 7 13 10 9 1 10 9 2
20 11 11 11 2 9 0 2 13 10 9 13 1 10 9 11 2 9 11 2 2
20 10 9 1 10 11 13 9 1 15 1 11 1 11 2 1 9 1 11 2 8
18 3 1 10 9 1 12 2 10 11 11 4 13 1 9 7 0 9 2
25 3 0 9 2 15 4 13 10 9 0 1 10 9 7 10 9 9 2 3 0 9 7 9 0 2
37 7 3 2 1 12 1 10 9 1 11 15 13 10 9 16 1 0 13 0 1 10 9 1 10 9 1 10 9 1 10 9 1 10 15 13 0 2
13 13 10 9 0 7 13 10 9 0 7 10 9 2
17 10 9 13 3 1 9 1 15 0 9 1 9 1 9 7 9 2
32 1 9 2 9 13 10 9 0 0 13 3 1 10 12 5 1 9 0 1 9 1 9 0 1 12 9 13 1 10 9 0 2
25 10 9 13 10 9 1 9 2 10 9 1 10 9 1 11 13 0 3 7 3 1 10 1 11 2
17 9 4 4 13 1 10 9 1 10 9 0 11 12 11 1 12 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 9 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
13 1 12 13 11 7 13 1 11 1 10 9 11 2
23 15 13 1 15 1 10 9 0 13 1 11 11 11 1 9 3 1 9 7 1 10 11 2
18 4 13 10 9 0 1 10 9 0 2 10 9 9 7 10 9 0 2
52 3 2 10 11 1 11 11 4 13 1 10 10 9 1 15 1 10 9 1 9 1 9 2 0 1 11 1 11 7 11 1 10 11 2 9 3 0 1 15 16 13 10 9 1 9 1 10 9 1 9 11 2
55 12 9 3 1 10 9 16 4 13 1 10 9 2 13 0 13 1 9 0 0 1 10 9 2 9 0 0 1 9 1 9 1 11 11 7 9 16 13 0 1 13 9 0 1 12 7 12 9 0 2 10 5 12 2 2
31 10 9 13 10 9 1 9 7 10 9 1 13 7 13 9 7 9 1 16 4 13 9 1 9 0 7 1 9 1 9 2
33 1 13 15 1 10 11 1 11 11 10 9 8 2 9 2 10 9 4 13 1 9 3 1 10 9 13 1 10 9 1 11 11 2
11 3 15 2 1 11 2 10 9 15 13 2
26 13 10 9 0 1 12 9 2 12 9 5 2 2 1 9 1 10 9 1 12 9 2 12 9 2 2
26 10 9 1 10 9 1 10 9 13 0 13 15 1 10 9 1 13 10 9 1 9 1 10 11 11 2
13 3 1 15 9 2 13 1 11 1 10 9 0 2
32 10 12 9 7 10 10 0 9 2 3 1 11 11 2 13 3 13 1 10 9 1 10 9 7 1 10 9 1 10 11 11 2
38 11 11 1 11 2 11 11 2 11 2 12 1 11 1 12 2 2 3 13 1 11 2 13 10 9 0 16 13 1 10 11 1 10 11 12 1 11 2
34 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 10 9 0 2 16 15 13 1 13 3 1 9 7 3 1 10 9 2
14 13 9 1 10 11 1 11 2 3 15 13 1 12 2
15 11 11 13 1 10 9 1 9 12 2 12 1 12 9 2
27 10 9 0 1 10 9 1 9 2 3 13 1 10 9 0 1 9 7 9 2 15 13 1 13 10 9 2
12 10 9 4 13 1 10 9 0 1 10 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
32 11 1 12 13 10 9 1 0 9 2 11 11 2 2 16 13 16 11 4 13 10 9 7 13 10 15 9 16 10 4 13 2
6 13 12 9 1 9 2
17 3 13 10 9 1 10 11 1 10 11 7 10 11 11 11 11 2
49 10 9 13 10 0 9 1 10 9 1 10 9 0 13 10 9 1 10 9 0 2 15 16 15 4 13 1 10 9 1 10 9 7 10 9 1 10 9 1 10 9 0 2 13 0 9 1 9 2
21 13 10 9 0 1 9 2 7 15 1 10 9 16 15 13 4 13 1 9 0 2
42 10 9 1 9 2 16 13 1 3 1 12 9 1 11 7 3 1 12 9 1 11 2 13 16 10 9 1 10 9 0 13 1 13 10 9 1 9 0 1 10 9 2
14 1 10 0 9 1 10 12 8 4 13 3 1 9 2
27 1 10 9 1 10 12 2 3 13 10 9 13 1 10 9 1 13 10 9 0 2 0 1 10 10 9 2
29 13 10 12 9 1 11 1 10 9 1 11 1 9 1 10 11 11 2 12 1 11 7 10 11 11 12 1 11 2
38 1 9 0 2 10 9 15 13 1 10 9 2 11 11 2 2 2 11 11 11 11 2 2 2 11 8 11 2 2 2 11 11 2 7 2 11 2 2
37 10 9 0 13 10 9 1 10 0 9 1 10 9 1 10 9 11 1 9 1 10 9 1 11 2 16 13 10 9 1 9 0 15 13 10 9 2
22 10 9 13 13 1 10 9 1 11 2 11 2 7 13 9 7 9 1 11 1 12 2
7 10 9 13 3 10 9 2
24 10 11 11 11 13 10 9 13 1 9 0 0 1 9 2 13 1 9 0 1 10 9 0 2
22 10 9 1 9 4 13 1 10 9 2 13 3 10 9 1 10 9 1 11 7 11 2
45 10 9 1 10 11 11 13 0 1 10 9 11 2 7 13 9 1 10 9 1 10 11 1 9 1 11 11 11 11 1 11 2 10 11 11 16 4 1 10 9 2 1 10 11 2
6 2 15 13 1 11 2
19 15 13 1 12 1 10 0 9 2 1 10 15 4 13 9 0 1 12 2
23 11 3 13 1 9 1 10 9 9 7 9 1 9 0 7 0 16 13 1 13 10 9 2
12 13 10 9 1 11 1 10 9 7 0 9 2
41 10 9 13 0 1 13 13 3 1 10 9 0 1 9 0 2 8 2 7 3 9 1 10 9 1 9 0 13 11 11 16 13 10 11 11 1 9 1 9 0 2
9 13 1 9 0 3 1 10 9 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
18 10 9 13 10 9 9 1 9 12 3 1 10 9 12 1 10 9 2
43 11 13 10 9 9 12 1 10 9 1 11 11 2 11 11 2 13 1 12 1 10 9 0 1 11 2 16 1 10 9 13 10 9 9 3 13 11 11 7 3 11 11 2
21 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
15 10 9 1 10 9 15 13 13 10 0 9 1 9 9 2
21 10 9 11 11 11 13 10 9 0 1 10 11 1 11 11 16 13 3 12 9 2
47 9 1 10 8 7 10 9 13 1 10 9 0 2 16 15 13 10 0 9 1 10 9 1 10 16 4 13 10 9 1 10 9 2 2 1 9 1 10 9 16 13 10 9 1 9 0 2
21 13 10 9 1 10 9 1 11 11 7 1 10 9 13 13 15 12 5 1 3 2
16 13 13 1 10 9 2 10 9 1 9 2 7 15 13 0 2
18 11 13 10 9 13 1 10 9 1 10 11 1 10 9 0 1 11 2
10 13 1 10 9 9 2 9 7 9 2
22 1 10 9 12 2 13 1 10 9 0 1 11 11 2 7 13 10 9 1 12 9 2
12 13 12 9 1 10 9 1 10 9 1 9 2
23 12 1 10 12 9 1 11 11 4 13 1 10 9 1 10 0 9 1 9 1 10 9 2
54 11 13 1 3 9 1 10 11 7 10 9 15 4 13 1 12 9 1 13 15 16 10 9 0 13 13 1 11 7 3 1 10 9 11 2 15 16 13 1 10 11 16 3 13 0 10 9 7 10 0 9 1 11 2
14 3 13 9 3 0 9 10 9 7 9 1 10 9 2
24 10 9 1 10 8 4 13 15 13 9 1 10 9 9 0 1 12 5 9 7 12 5 9 2
16 3 15 13 3 13 1 10 9 1 11 1 10 9 1 12 2
12 10 9 1 9 4 13 1 12 9 1 9 2
18 1 12 13 1 13 1 11 2 3 13 1 9 0 1 10 9 0 2
22 13 1 11 1 12 2 7 1 12 7 12 13 9 1 10 9 1 10 9 1 11 2
18 16 11 7 11 13 10 0 9 0 2 11 3 13 1 9 1 11 2
20 1 12 11 13 1 10 9 10 0 9 1 10 8 11 13 1 10 11 11 2
36 10 9 1 10 9 13 1 10 9 12 1 10 11 11 11 2 12 1 11 1 11 12 2 16 16 10 9 1 10 9 13 1 10 9 12 2
26 11 11 11 2 12 1 11 1 12 2 11 2 2 3 13 1 11 11 2 13 10 9 7 9 0 2
100 11 13 0 9 7 9 2 9 1 10 15 3 15 13 10 11 1 11 2 11 7 11 2 12 2 2 11 1 11 2 12 2 2 11 1 10 9 1 11 2 12 2 2 11 2 11 7 11 2 12 2 2 11 10 9 2 12 2 2 11 7 11 2 12 2 2 11 1 11 2 12 2 2 11 1 11 2 12 2 2 11 1 11 2 11 1 9 2 0 2 12 2 2 11 1 11 11 2 12 2
33 10 9 3 0 2 11 11 11 2 15 4 13 1 10 9 1 10 11 1 11 2 7 13 15 1 3 12 9 13 1 10 9 2
29 3 13 13 16 9 0 1 3 13 10 9 0 2 7 13 2 13 16 4 13 0 7 3 13 1 15 13 15 2
30 13 9 1 10 9 7 13 2 15 2 16 3 13 9 0 7 3 0 9 1 9 2 9 4 13 15 1 10 9 2
12 3 13 11 1 11 2 11 11 7 10 11 2
14 15 1 9 4 13 2 10 9 2 1 10 11 11 2
16 1 9 2 4 13 9 1 10 3 15 0 9 1 10 9 2
23 10 11 11 12 13 10 9 1 10 11 11 1 10 9 0 13 1 11 1 10 9 0 2
19 13 1 10 9 0 2 10 9 0 1 10 0 9 13 10 9 1 11 2
62 1 10 12 9 2 10 9 1 11 13 0 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
16 13 3 9 1 9 2 8 8 8 8 8 8 15 8 2 2
37 10 9 1 9 0 13 10 16 15 13 1 10 0 2 9 2 2 16 4 13 1 2 9 2 2 16 15 13 1 10 11 11 11 2 11 2 2
13 1 12 1 12 2 13 10 9 1 12 1 12 2
34 1 15 1 10 9 2 10 9 15 13 1 10 9 1 10 16 15 13 1 9 9 1 9 0 2 9 0 7 0 1 10 10 9 2
78 10 9 13 1 9 1 10 9 1 10 9 0 2 11 11 11 2 15 13 1 10 9 1 13 15 1 9 8 13 10 9 0 1 13 10 9 0 1 10 9 0 2 1 15 10 9 11 11 13 10 9 1 12 12 9 1 9 1 10 9 2 13 13 2 12 12 9 3 1 15 13 1 10 9 1 10 9 2
15 3 2 13 1 13 9 1 10 9 1 9 2 13 13 2
32 13 11 2 9 1 9 2 7 11 2 11 2 2 10 9 1 10 9 0 13 1 10 9 1 15 15 4 13 1 9 0 2
21 11 11 13 10 9 1 12 9 13 1 11 15 13 10 9 1 13 15 1 9 2
25 13 16 15 4 1 13 10 9 1 10 9 7 15 13 10 9 2 2 13 10 9 1 10 9 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
22 7 10 9 15 13 7 15 13 1 11 3 9 3 0 1 13 15 13 10 9 0 2
58 10 9 4 3 13 1 13 10 9 1 13 9 7 9 2 1 15 15 15 13 1 10 9 1 9 0 1 9 7 9 1 9 2 16 1 16 10 9 13 1 10 0 9 0 2 10 9 1 9 2 10 9 1 9 7 9 2 8
25 11 11 11 7 11 2 11 2 12 2 8 2 12 2 13 10 9 7 0 1 10 11 1 11 2
37 15 13 1 10 9 16 9 1 9 1 10 9 1 10 9 1 10 9 0 9 1 10 9 0 7 1 10 9 1 10 15 1 15 1 10 9 2
23 10 9 13 3 0 7 0 7 1 0 13 10 9 3 0 1 13 9 0 1 10 9 2
24 11 11 11 1 11 3 1 10 9 1 10 9 0 13 10 9 1 9 3 13 2 11 2 2
27 10 9 13 1 10 9 0 8 2 9 2 7 8 2 9 2 7 13 13 2 10 9 1 10 9 2 2
17 15 4 13 1 10 9 2 7 13 3 15 15 13 1 10 9 2
30 10 9 1 10 9 13 3 10 0 9 1 10 9 0 2 15 13 10 9 2 9 7 9 2 7 13 3 10 9 2
13 10 9 16 15 13 13 16 15 13 3 10 9 2
47 15 1 10 9 2 1 10 3 0 11 11 2 7 9 1 10 9 1 9 1 9 13 1 10 9 1 10 0 9 0 16 13 10 9 7 1 10 9 0 13 1 10 9 1 10 9 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
22 11 11 2 13 1 12 1 11 2 1 10 9 1 11 2 11 2 13 10 9 0 2
44 1 10 9 2 11 4 13 16 10 9 1 10 9 2 13 10 9 1 10 9 1 10 9 1 10 9 7 13 3 3 10 9 2 13 3 16 10 0 9 13 3 0 2 2
25 15 4 13 10 9 1 9 3 0 7 9 13 1 9 1 10 11 2 3 10 9 2 11 2 2
27 16 10 9 15 13 1 10 9 2 4 13 1 10 9 1 11 7 9 3 7 12 9 13 1 10 9 2
36 11 13 1 11 12 9 0 7 13 1 10 15 1 10 9 1 10 9 2 10 9 11 11 11 2 9 1 10 9 0 2 15 13 10 9 2
25 3 4 13 9 0 0 2 1 10 9 1 9 1 10 9 2 16 13 10 9 1 10 9 0 2
8 15 13 0 9 0 1 11 2
28 13 10 9 1 12 9 5 13 12 5 1 10 9 2 12 5 1 10 9 7 12 5 1 10 10 9 0 2
34 10 11 13 0 1 10 13 1 10 9 1 9 0 7 3 13 1 13 15 2 16 10 11 13 10 9 1 10 11 7 13 10 9 2
20 10 9 1 10 9 0 1 10 9 4 13 1 10 9 1 10 9 2 11 2
25 10 9 1 11 4 3 13 1 9 0 16 13 1 10 9 2 10 9 2 7 3 2 10 9 2
28 15 4 13 10 9 1 9 1 15 1 10 9 0 2 10 9 7 10 9 2 3 16 13 10 9 1 15 2
24 10 9 16 13 0 1 10 9 1 10 0 9 2 0 2 1 10 9 13 1 10 0 9 2
31 10 9 1 9 13 1 10 9 4 13 10 12 9 1 9 1 9 0 1 10 9 1 10 12 9 1 9 1 9 0 2
38 3 13 1 15 16 13 15 1 15 2 15 13 12 9 2 15 13 2 1 10 9 15 13 1 10 9 8 10 9 8 10 9 15 13 1 15 2 2
10 13 1 10 9 1 11 1 10 12 2
45 10 0 9 2 13 10 12 9 2 13 1 12 9 1 10 9 1 11 1 11 1 10 9 1 9 1 9 1 9 7 13 1 10 9 10 9 0 1 9 7 10 9 0 0 2
63 11 15 13 13 1 9 1 10 11 2 3 3 1 10 11 11 2 3 3 1 10 9 1 9 2 1 10 15 3 3 15 13 12 5 2 7 3 1 11 2 10 9 1 10 9 1 10 15 13 2 10 9 1 11 2 1 10 15 3 13 12 5 2
15 13 10 12 9 1 0 9 1 9 13 1 10 12 9 2
27 13 1 10 11 1 11 11 1 11 1 12 1 10 9 0 2 11 1 11 2 1 10 9 1 12 9 2
38 10 9 15 13 16 16 13 10 9 15 13 16 3 16 13 0 3 7 4 13 3 1 12 9 7 15 13 16 3 13 0 7 3 0 1 10 9 2
14 10 9 13 10 9 13 1 10 11 1 11 1 12 2
10 8 11 13 10 9 1 11 2 9 2
44 13 16 1 10 9 1 9 1 10 8 2 15 4 13 10 9 1 10 9 0 7 0 2 0 1 10 9 1 9 1 10 9 2 1 10 9 1 10 0 9 1 9 0 2
5 4 13 1 12 2
5 13 9 1 9 2
6 10 9 13 1 15 2
18 10 9 1 10 9 13 0 7 0 2 3 1 13 3 0 7 0 2
38 15 13 1 11 11 11 11 2 11 13 16 15 13 0 1 16 10 9 15 13 1 10 9 1 10 0 9 7 3 16 4 13 9 3 1 10 9 2
10 12 9 0 10 9 15 13 10 9 2
31 15 13 16 10 9 13 0 16 13 10 9 1 13 15 1 9 1 10 9 2 13 13 2 1 13 1 9 1 10 9 2
21 13 13 2 10 9 0 13 10 9 12 2 12 2 12 2 12 2 12 7 12 2
39 7 16 1 0 9 13 10 9 1 13 10 9 0 2 15 4 13 10 0 9 2 9 1 9 1 9 0 2 9 0 2 0 9 1 9 7 9 0 2
25 13 10 9 1 9 1 10 9 1 11 2 11 1 10 9 12 2 12 13 2 11 11 11 2 2
50 1 15 4 13 1 10 9 2 10 9 2 9 7 10 9 0 1 13 1 10 9 1 10 9 16 1 9 15 4 13 1 16 1 10 9 3 13 10 9 1 9 2 13 15 3 1 10 9 0 2
11 3 13 3 7 3 15 15 13 1 15 2
27 10 9 0 13 15 10 9 1 10 0 9 7 10 9 7 9 1 10 11 1 10 9 12 1 10 12 2
8 13 3 1 10 9 3 0 2
36 13 9 1 9 13 10 9 1 9 1 11 1 12 2 10 9 13 12 2 2 15 16 13 0 1 10 0 9 1 2 4 13 10 9 2 2
20 13 1 13 16 10 0 9 1 9 13 16 10 9 0 13 10 9 1 11 2
12 4 13 10 9 1 9 7 9 1 10 9 2
30 10 9 13 10 9 1 9 1 10 9 11 7 13 1 10 0 9 1 11 2 10 0 9 1 10 9 1 9 0 2
22 15 13 1 10 11 11 11 7 10 9 1 10 9 7 15 13 1 10 9 1 11 2
13 15 13 16 4 13 2 9 1 10 0 9 2 2
40 11 13 10 9 12 0 9 0 1 10 16 13 13 9 0 16 13 9 0 0 13 1 10 9 0 7 10 9 1 9 8 16 13 1 10 9 10 9 0 2
36 11 11 13 10 9 16 13 10 9 2 7 10 9 15 13 13 1 13 10 9 1 10 9 2 9 2 9 2 9 7 9 4 13 3 2 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 4 1 9 0 7 2 12 5 2 12 9 5 13 9 2
21 13 9 1 10 10 9 1 10 9 2 7 3 1 10 9 1 10 9 1 11 2
18 11 2 13 1 11 11 2 13 10 9 1 10 9 1 9 1 11 2
7 10 0 9 15 13 11 2
29 13 3 0 10 9 16 1 0 9 10 9 7 9 4 13 1 13 3 2 3 1 10 9 1 10 11 1 11 2
28 11 11 13 10 9 0 3 1 10 9 2 8 2 2 3 1 10 9 2 11 2 11 2 3 7 11 2 2
9 13 10 9 13 7 13 1 10 9
34 10 11 1 11 11 4 13 10 11 1 9 1 11 2 7 13 2 1 10 9 2 1 10 9 1 10 11 2 11 1 10 9 0 2
38 10 9 0 1 10 9 0 2 7 0 2 13 13 0 9 0 2 9 2 0 2 0 2 8 2 13 1 10 9 1 9 2 7 0 15 1 15 2
25 4 13 2 3 2 1 10 9 3 0 1 11 2 13 1 11 2 11 2 11 2 11 7 11 2
25 1 10 9 2 11 4 13 1 10 9 1 11 16 13 1 10 11 11 1 13 1 10 9 8 2
18 11 13 16 10 9 1 10 9 13 1 15 2 16 3 13 13 2 2
24 1 0 2 10 9 4 13 10 9 1 11 2 3 0 1 12 1 10 9 1 11 11 11 2
13 11 11 11 13 1 11 10 12 1 11 1 12 2
20 13 10 9 2 1 9 2 1 11 7 11 1 12 1 10 9 1 11 11 2
31 3 2 13 10 9 1 9 0 2 16 13 1 12 9 7 16 15 13 1 10 9 11 11 1 11 2 10 0 9 0 2
17 10 0 7 0 9 1 9 0 2 0 7 0 13 3 10 9 2
24 13 10 9 0 2 15 13 1 9 1 9 1 10 9 1 10 9 1 10 9 1 8 9 2
8 10 9 1 10 11 15 13 2
10 10 9 2 11 11 15 13 10 9 2
11 10 9 1 11 15 13 13 1 10 9 2
5 13 9 3 0 2
41 10 9 13 3 10 9 3 1 10 9 7 1 10 9 1 9 1 9 1 10 12 9 1 10 9 1 15 9 1 12 2 7 15 13 10 0 9 1 10 9 2
13 1 9 10 10 9 0 1 10 9 0 13 0 2
15 1 11 15 13 1 10 12 1 11 1 10 12 1 11 2
5 11 7 11 11 2
3 11 11 2
49 3 2 16 13 1 10 11 1 11 2 11 7 11 2 15 13 1 10 9 0 1 10 9 2 10 9 7 10 9 2 8 5 8 5 8 2 0 7 10 0 9 1 9 1 9 0 1 11 2
27 1 9 1 12 2 10 9 13 10 9 1 9 0 7 13 10 2 9 1 9 2 1 13 3 10 9 2
11 13 10 9 0 2 3 13 5 9 0 2
26 4 4 7 13 9 7 9 2 3 7 1 9 3 13 10 9 1 9 7 10 9 1 9 1 9 2
8 15 13 1 11 2 11 11 2
20 1 10 12 9 4 1 13 10 9 2 10 11 2 2 1 10 9 11 11 2
39 11 2 10 9 1 0 9 2 7 10 9 11 11 5 11 11 15 13 16 13 2 13 2 1 10 9 1 10 11 11 1 11 1 13 1 10 0 11 2
39 10 9 11 7 11 4 13 1 11 11 2 13 7 9 1 10 9 0 7 13 1 11 1 11 2 13 10 9 1 11 1 10 13 10 9 1 12 9 2
23 1 12 7 12 2 13 1 10 9 1 9 0 1 10 11 1 10 11 11 2 1 11 2
24 3 15 13 1 9 1 9 2 9 1 9 2 13 3 1 9 0 7 9 1 9 1 9 2
17 1 10 9 0 15 13 0 13 10 9 12 1 11 1 10 11 2
43 1 9 1 10 0 9 0 1 10 9 2 9 1 9 7 9 1 10 9 1 10 9 0 2 13 1 10 9 9 0 2 0 7 0 2 16 13 3 16 13 10 9 2
23 1 9 1 10 0 9 1 9 15 13 10 9 1 9 16 15 13 1 9 1 10 9 2
48 10 9 4 13 10 9 3 0 1 11 1 9 1 10 9 2 1 10 9 1 12 2 1 10 11 1 10 11 11 16 13 1 10 9 7 4 13 10 9 3 1 10 9 1 10 9 0 2
39 3 3 2 11 13 1 13 1 11 2 7 13 16 15 13 10 9 1 10 11 1 10 9 0 2 3 7 3 4 13 1 10 11 11 1 10 0 9 2
12 1 9 1 10 9 3 4 13 3 10 9 2
26 3 3 3 15 13 16 15 13 1 15 3 16 15 13 7 13 0 7 15 15 13 1 9 1 9 2
9 13 10 9 1 10 9 10 11 2
57 3 2 13 16 2 1 10 9 0 2 2 15 13 1 10 9 1 10 9 1 10 9 2 2 1 9 16 10 9 0 16 3 15 13 1 10 9 0 1 11 4 4 13 10 9 1 9 16 13 1 9 3 0 1 10 9 2
30 1 10 9 2 13 0 15 4 13 1 9 0 7 1 10 9 2 13 15 9 1 10 9 16 13 16 13 13 15 2
11 13 1 10 9 1 4 13 1 10 9 2
14 3 15 13 1 10 9 1 10 9 7 1 10 9 2
20 10 9 0 2 15 15 1 10 9 7 10 9 9 13 3 1 10 9 0 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
47 10 9 2 13 1 11 11 2 15 4 13 1 11 11 2 16 15 4 13 0 9 2 13 15 16 10 9 2 11 2 13 3 0 1 11 2 7 3 13 1 10 9 0 1 10 9 2
14 10 9 1 11 13 1 9 0 13 1 10 9 11 2
77 13 0 13 9 1 10 0 9 9 9 11 11 11 2 13 1 11 11 2 15 13 10 11 11 11 12 7 12 2 13 10 0 10 3 0 2 3 16 4 13 9 1 10 9 1 9 0 1 11 7 13 1 10 11 11 1 11 2 7 1 10 9 0 16 4 13 9 1 10 9 1 9 1 11 2 11 2
12 10 9 13 12 9 7 10 0 9 1 9 2
111 10 9 13 10 0 9 2 9 7 9 2 16 15 13 0 1 10 0 9 2 13 0 2 1 10 0 9 2 1 10 0 9 16 13 10 9 0 1 11 2 3 15 13 1 10 9 0 1 10 9 2 7 10 0 9 2 16 13 12 9 1 11 2 13 15 1 0 9 2 1 10 9 7 9 1 10 11 11 1 10 9 7 9 1 10 0 9 0 16 13 1 10 9 0 2 10 11 1 11 2 13 9 1 10 9 12 1 10 9 0 2
39 1 12 2 11 13 15 1 10 12 9 13 1 15 1 10 2 11 11 11 2 2 9 16 13 1 15 1 10 0 9 1 11 11 11 7 1 11 11 2
21 11 2 9 7 9 13 10 9 1 10 9 16 13 13 10 0 9 1 10 9 2
7 4 13 3 1 12 9 2
15 16 3 15 15 13 13 10 9 3 0 1 10 9 0 2
39 10 9 1 10 0 9 0 13 16 1 10 11 1 9 1 11 10 0 9 15 13 1 9 7 16 3 4 13 1 10 10 9 1 10 9 13 10 9 2
28 1 10 0 9 0 13 0 0 9 7 9 1 13 1 10 9 10 9 3 0 7 0 1 10 9 1 9 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
59 1 10 12 9 2 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
24 10 9 1 9 15 4 13 0 7 13 10 12 5 1 10 9 1 12 9 3 13 1 11 2
25 10 9 7 10 9 0 0 9 13 2 7 15 13 10 9 1 10 9 1 10 9 1 10 9 2
24 10 9 1 11 15 13 1 10 9 0 13 11 11 2 1 10 9 1 10 9 11 1 12 2
34 1 10 9 1 10 9 13 1 9 1 9 7 2 3 2 4 13 1 0 9 2 1 15 2 1 10 9 2 9 2 9 7 9 2
152 7 3 3 3 1 10 0 9 2 7 13 15 13 1 0 9 2 16 13 7 13 1 13 15 1 9 0 1 10 0 9 0 13 1 7 1 9 1 10 11 11 11 1 9 1 0 9 7 1 10 0 9 2 7 15 1 9 4 4 13 1 9 1 9 1 0 2 13 15 2 10 9 10 9 1 10 11 11 2 16 13 3 3 1 10 0 9 1 10 16 15 13 7 16 15 13 3 0 1 10 9 1 10 9 1 10 9 2 1 10 8 8 2 1 10 9 2 7 3 15 1 10 9 0 16 13 3 10 9 7 13 10 9 0 2 1 9 3 1 9 15 9 1 10 9 0 1 10 1 10 9 2
13 10 0 9 16 13 10 9 13 10 1 10 9 2
47 10 9 0 4 13 1 9 7 9 13 1 9 1 9 2 1 9 2 10 9 3 13 3 0 2 7 3 10 9 1 10 9 2 1 9 1 9 1 9 7 9 16 13 1 13 9 2
17 1 10 9 0 10 9 15 13 1 10 9 7 9 1 10 9 2
23 11 13 16 13 10 9 1 15 1 10 2 9 0 2 0 1 3 7 0 1 3 2 2
12 10 9 1 9 1 10 9 13 1 5 12 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
64 13 3 16 10 0 9 1 11 13 10 9 2 11 2 1 13 15 1 11 1 13 2 9 1 3 13 1 13 10 9 10 9 0 2 11 11 2 9 7 15 13 9 1 10 9 11 2 1 11 2 1 15 15 1 11 10 9 3 13 3 0 7 0 2
17 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 11 2
29 13 3 0 10 9 7 1 0 9 10 9 7 9 4 13 1 13 3 2 0 1 10 9 1 10 11 1 11 2
6 11 11 13 10 9 2
26 11 1 11 3 13 10 9 1 10 9 2 8 2 8 2 8 2 7 13 16 10 9 13 1 11 2
12 15 4 7 13 15 16 3 11 13 10 9 2
16 11 7 11 13 0 1 10 9 2 7 11 3 15 13 0 2
9 13 9 1 10 11 11 1 11 2
42 13 1 9 1 13 16 3 2 7 15 13 13 1 15 7 13 10 9 1 10 9 1 10 13 16 13 10 9 3 7 13 16 10 9 15 13 1 10 9 0 0 2
20 13 1 10 9 1 11 2 1 12 9 1 9 7 10 9 16 13 10 9 2
13 15 13 10 9 1 10 12 1 11 1 10 9 2
29 13 13 10 9 2 3 13 10 9 1 10 12 9 13 15 1 13 1 10 0 9 9 1 13 10 9 1 9 2
46 1 10 9 1 10 11 15 4 1 13 10 9 1 10 9 16 4 13 9 0 1 10 9 2 10 9 7 10 9 1 10 15 2 3 7 10 9 0 1 10 9 0 16 13 0 2
32 13 10 0 9 0 0 10 12 1 11 1 10 9 2 10 9 1 9 1 11 11 7 11 11 11 1 10 11 11 11 11 2
49 10 9 0 13 10 9 1 11 11 1 11 2 9 0 1 10 11 1 10 11 2 1 10 9 1 10 9 1 10 11 7 10 9 1 9 0 16 3 13 1 16 15 15 13 1 8 2 8 2
34 10 11 1 11 13 10 9 1 10 9 0 1 11 1 9 1 10 9 12 1 10 9 12 2 16 10 0 9 4 13 1 10 9 2
15 1 10 0 9 2 10 11 11 11 11 13 1 10 9 2
18 1 10 0 9 10 9 13 0 7 10 9 13 3 9 7 9 0 2
37 1 10 9 2 10 9 13 3 0 1 9 0 2 16 4 13 1 13 10 9 0 7 0 1 3 12 9 16 13 1 9 1 10 9 1 9 2
25 10 9 13 10 9 1 9 1 10 9 3 0 16 15 13 1 10 9 2 9 7 9 1 11 2
16 10 9 1 11 11 13 0 1 9 3 0 2 9 7 9 2
17 13 0 1 10 9 1 9 1 11 1 12 9 7 13 12 9 2
65 10 9 13 10 9 2 10 12 1 11 1 12 2 1 10 9 0 1 10 9 1 10 11 2 11 11 11 2 7 1 10 11 2 11 1 9 1 10 9 0 2 2 15 13 10 0 9 1 10 9 1 10 9 0 2 16 13 1 10 9 1 12 3 0 2
29 3 2 10 9 4 13 13 15 1 10 9 1 10 9 11 11 10 9 1 12 12 9 7 10 9 1 12 9 2
16 10 9 1 10 9 13 1 9 1 10 9 0 1 0 9 2
26 13 10 9 0 1 10 11 11 11 7 1 9 1 10 11 11 11 1 11 2 9 1 10 9 0 2
26 1 9 0 0 2 7 3 0 2 13 1 10 9 1 10 9 1 9 0 2 10 2 11 11 2 2
8 13 9 1 10 11 1 11 2
36 11 2 11 1 9 0 2 11 1 11 1 9 0 2 13 10 9 7 9 0 2 13 1 10 9 1 10 11 1 10 9 1 11 2 11 2
43 11 2 3 2 13 10 9 2 1 0 9 2 2 1 15 15 13 2 0 2 2 9 16 4 13 9 1 9 2 13 16 13 9 2 10 15 16 15 15 13 13 2 2
6 10 9 0 13 0 2
33 1 9 13 2 1 2 11 1 10 11 2 10 9 13 16 13 2 10 9 1 10 9 2 2 1 10 9 1 10 9 0 2 2
15 10 9 15 13 1 9 1 9 7 13 9 1 9 0 2
21 10 9 13 3 1 9 10 9 1 10 9 0 2 10 9 0 7 10 9 0 2
39 4 13 1 0 1 12 1 10 9 1 9 2 0 1 11 11 2 1 10 9 0 1 10 9 0 0 11 7 11 15 11 11 4 13 1 11 1 12 2
34 11 13 16 10 9 1 9 1 10 8 7 10 9 4 13 16 10 9 13 10 9 1 9 2 3 7 2 10 9 3 13 9 0 2
29 3 1 10 9 2 3 13 13 10 9 2 1 15 15 15 13 1 13 9 2 16 3 4 13 1 10 9 2 2
31 3 15 3 13 0 1 13 15 1 9 2 16 10 9 0 4 13 10 0 9 1 9 1 10 9 2 16 13 10 9 2
42 1 13 1 12 2 11 13 10 0 9 1 9 2 1 9 1 9 7 9 0 16 13 1 10 9 2 9 16 13 1 10 9 1 10 0 9 2 10 11 11 11 2
6 3 13 1 10 9 2
23 13 9 0 1 11 7 11 2 3 7 9 0 1 11 2 11 2 7 11 2 11 2 2
17 10 9 1 11 1 11 13 1 10 9 1 11 11 2 11 2 2
21 13 1 10 9 1 10 9 0 1 11 2 0 1 11 2 11 2 9 7 11 2
34 10 9 1 10 9 4 13 3 1 9 2 1 10 9 3 15 13 11 2 11 2 7 9 2 13 10 9 1 9 1 0 9 2 2
22 10 9 4 0 1 10 9 0 1 9 0 2 1 15 1 10 9 0 1 10 9 2
46 11 11 2 9 1 10 9 1 11 2 13 16 11 11 2 1 12 9 2 4 13 0 1 10 9 1 13 1 10 9 2 1 11 11 2 1 11 7 11 2 10 11 1 10 9 2
7 10 9 3 13 13 9 2
48 3 2 1 10 9 16 3 13 10 9 1 10 9 15 4 13 10 9 0 2 3 1 10 9 1 9 2 1 10 15 0 9 13 13 10 9 1 10 9 2 10 9 4 13 1 10 9 2
37 10 9 13 0 7 1 9 0 2 7 15 13 1 13 16 13 1 9 16 10 9 13 11 2 16 13 0 1 15 2 16 13 1 13 15 11 2
44 1 13 10 9 1 11 1 10 10 9 2 13 15 1 9 2 15 13 1 10 11 1 10 11 11 1 11 11 7 10 11 11 15 15 13 10 9 2 11 2 1 13 15 2
24 1 13 10 11 1 10 11 1 11 2 11 13 13 10 9 1 10 9 2 7 1 12 5 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
22 11 13 10 9 7 9 0 2 13 1 10 9 1 11 11 2 1 10 9 1 11 2
15 10 9 2 13 1 9 7 1 9 13 1 10 9 0 2
26 10 9 11 11 1 11 13 16 13 10 9 1 10 9 0 1 10 13 1 10 9 13 1 10 9 2
23 10 9 0 1 9 13 10 9 1 9 0 13 1 13 10 9 0 0 1 9 1 11 2
9 13 1 15 3 1 13 10 9 2
24 10 11 3 13 1 10 9 0 11 11 11 1 10 12 1 10 12 1 11 1 10 9 12 2
14 13 10 9 1 11 7 3 13 15 2 13 10 9 2
30 10 9 13 15 0 13 1 10 0 9 1 9 13 1 13 10 9 1 9 13 1 10 9 1 9 1 10 9 0 2
18 1 12 13 10 0 9 7 5 8 1 10 9 1 10 9 1 11 2
18 10 0 9 4 4 13 2 1 10 0 16 9 7 10 9 4 13 2
27 13 10 0 9 1 10 9 13 10 9 0 1 10 9 2 16 13 3 13 10 9 1 9 1 10 9 2
26 1 3 15 4 13 1 11 1 10 9 2 13 10 9 1 13 1 9 1 16 15 15 4 13 3 2
16 10 11 11 2 13 10 9 1 9 16 3 15 4 13 0 2
11 13 3 1 12 9 10 11 2 11 11 2
20 1 9 15 4 13 10 2 9 1 9 2 1 3 4 13 3 2 3 0 2
36 10 9 4 13 1 10 9 9 12 7 4 4 13 1 10 0 11 11 2 13 1 10 11 11 1 0 9 2 15 13 1 10 0 9 0 2
48 10 11 13 10 9 7 9 1 11 2 1 10 9 1 10 11 11 2 0 1 10 9 0 1 11 1 10 11 1 10 9 1 10 9 1 11 2 9 0 1 11 2 1 12 9 1 11 2
49 1 9 0 2 10 9 13 10 0 9 1 9 1 12 2 7 1 12 2 1 0 9 1 12 2 13 10 0 9 0 2 3 1 10 11 11 2 16 13 10 0 9 1 10 9 1 10 9 2
24 3 2 10 9 13 1 11 1 9 1 10 0 9 13 1 10 9 1 13 3 10 3 0 2
39 1 13 16 11 13 10 9 13 1 10 0 9 1 10 11 11 2 11 13 9 1 9 1 11 1 3 13 3 9 2 13 0 4 13 1 10 11 11 2
19 1 10 9 10 9 1 10 9 0 13 10 9 7 10 9 1 10 9 2
16 4 13 1 11 11 7 13 1 11 11 1 3 1 12 9 2
26 13 3 9 2 0 1 11 11 2 1 15 1 10 9 0 1 9 1 11 7 11 2 1 11 11 2
44 10 9 15 13 2 11 11 11 11 2 16 16 15 15 13 9 1 10 9 1 10 9 2 13 13 15 1 15 2 16 10 9 15 15 13 2 13 10 15 15 15 3 13 2
25 1 10 9 1 10 9 0 15 13 10 9 7 15 13 10 9 1 10 9 7 1 10 10 9 2
8 13 9 1 13 10 9 13 2
14 1 10 11 11 13 12 9 1 10 15 13 12 9 2
40 10 9 2 9 16 13 1 10 9 0 2 8 2 16 13 9 7 2 8 2 16 13 9 2 13 10 9 10 0 9 13 10 9 0 1 9 1 10 9 2
27 3 2 11 13 1 11 10 9 1 11 7 3 1 15 2 7 11 7 11 13 10 11 1 12 1 11 2
22 10 9 0 4 13 7 4 7 13 15 1 13 10 9 7 9 1 10 9 1 11 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
30 3 15 13 13 7 13 12 9 1 9 2 15 4 13 1 10 9 1 4 13 7 10 12 3 13 1 9 1 9 2
32 10 9 13 0 7 16 13 9 1 9 1 9 15 13 16 16 13 9 1 9 3 13 10 9 7 3 13 8 15 4 13 2
23 10 9 1 10 9 13 3 10 9 0 7 0 1 10 9 1 10 9 1 10 9 12 2
37 1 10 9 12 10 9 1 11 7 10 1 11 2 1 9 0 2 13 13 15 10 9 1 11 2 1 10 15 1 9 0 15 13 10 9 11 2
7 13 1 10 9 7 9 2
15 10 9 13 10 9 11 11 2 16 13 10 9 1 12 2
24 11 12 1 11 2 11 2 11 2 12 1 11 1 12 2 8 2 12 1 11 1 12 2 2
19 3 13 1 10 9 1 10 11 11 1 11 1 10 10 11 1 10 11 2
15 10 9 1 11 11 13 10 9 1 10 9 0 11 11 2
15 10 9 1 10 11 4 13 9 1 10 9 1 0 9 2
49 10 11 11 15 13 3 7 13 9 7 0 13 16 13 15 0 13 10 0 9 16 13 7 10 9 1 9 13 15 3 0 7 10 16 13 7 10 16 15 13 10 9 0 16 13 1 10 9 2
19 1 11 2 3 1 13 15 1 11 1 10 9 0 2 13 12 9 0 2
19 13 1 9 7 9 0 2 13 9 1 9 7 9 1 0 9 7 9 2
23 10 11 1 11 2 10 9 1 10 0 9 1 10 9 0 2 15 13 10 12 1 11 2
25 1 15 9 1 10 9 15 4 4 13 1 10 0 9 1 10 9 11 2 9 1 10 0 9 2
26 11 11 13 10 11 11 1 10 0 9 2 11 2 12 9 2 12 2 12 2 12 2 7 12 2 2
26 15 4 13 3 12 0 9 1 10 9 0 7 10 9 4 13 10 0 9 1 9 7 9 1 9 2
18 10 9 4 13 1 9 1 10 9 1 10 9 1 11 13 11 11 2
6 4 13 3 1 9 2
44 11 4 13 1 16 10 9 13 15 1 10 9 13 1 9 1 10 9 1 10 9 0 1 10 9 7 16 4 13 15 1 11 1 11 1 12 1 12 9 2 1 9 0 2
13 15 13 1 11 7 16 15 4 13 3 15 13 2
31 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 5 12 2 7 10 9 0 1 9 13 5 12 2
49 10 9 1 10 9 13 9 10 15 1 10 15 1 10 9 11 2 13 9 1 9 2 16 13 1 10 9 1 10 0 9 7 13 1 10 9 2 3 7 10 9 1 9 4 13 1 10 9 2
24 1 10 9 1 11 1 11 13 9 1 10 11 11 11 2 1 9 1 9 1 10 9 0 2
26 10 9 13 1 0 9 1 9 1 9 7 16 4 13 15 1 15 1 10 3 0 9 1 10 9 2
28 3 1 10 11 11 11 2 10 9 4 1 13 15 11 11 1 9 1 11 11 2 10 0 9 1 10 11 2
8 15 13 3 1 10 0 9 2
16 7 13 10 9 1 13 10 9 1 10 9 1 2 9 2 2
17 1 15 13 2 2 2 10 10 9 13 10 9 0 2 3 15 2
17 3 1 10 13 1 10 9 0 7 9 10 9 13 12 9 0 2
59 3 10 13 3 10 9 0 1 10 9 3 13 10 9 0 1 9 0 2 7 1 10 9 15 13 13 15 1 9 7 1 9 1 12 10 2 11 2 13 0 2 3 1 10 9 1 10 9 1 9 7 10 10 0 9 1 9 0 2
29 1 9 13 10 12 5 9 1 10 9 11 11 11 11 1 11 11 11 1 12 7 3 0 9 1 10 9 11 2
32 10 11 11 2 13 10 12 1 11 12 1 11 11 2 11 11 11 2 11 11 7 11 11 2 4 13 1 13 10 9 11 2
64 1 10 9 13 12 1 10 9 0 0 16 4 13 1 11 2 10 9 1 11 11 1 12 2 16 13 9 1 10 9 7 10 9 1 11 2 7 15 1 10 11 1 12 2 16 2 16 3 15 4 13 2 13 10 0 9 16 4 13 9 1 10 9 2
21 10 11 4 13 1 10 9 11 1 11 2 1 10 9 1 10 9 1 9 0 2
56 3 2 1 15 13 9 1 13 1 9 2 10 9 13 1 9 3 0 7 9 1 9 0 2 9 1 9 0 2 9 7 9 2 13 10 9 10 9 3 0 16 13 10 12 5 1 10 9 0 1 10 9 1 9 0 2
11 13 10 9 0 7 13 10 0 9 0 2
20 1 10 9 3 0 2 10 9 1 9 9 1 9 13 0 1 9 7 9 2
31 1 10 9 1 10 11 1 10 11 10 12 1 11 1 12 2 11 13 1 12 2 10 9 1 13 10 0 11 1 11 2
14 3 4 13 15 16 13 10 9 0 7 9 1 9 2
34 13 9 1 9 2 10 9 13 13 1 11 2 11 2 11 2 13 13 3 1 10 9 9 16 16 9 1 9 2 7 3 13 9 2
44 1 3 2 15 13 1 10 9 11 2 3 15 13 10 9 1 9 1 10 9 11 2 13 1 10 9 0 1 10 9 1 10 11 11 2 7 9 2 1 9 1 9 0 2
32 10 9 13 1 15 3 1 12 9 1 9 7 13 9 1 12 2 9 16 4 7 15 13 10 9 16 3 13 1 9 0 2
26 10 9 3 13 1 10 12 1 11 1 12 2 7 11 13 10 11 1 11 1 10 9 1 10 9 2
24 13 10 0 9 1 10 11 16 13 12 9 7 13 10 3 0 1 10 9 0 1 10 9 2
34 3 2 4 13 10 9 1 9 1 9 1 10 9 1 10 9 2 7 10 9 1 9 1 10 9 1 9 16 4 13 10 9 0 2
40 10 9 1 11 13 13 1 10 9 2 13 15 9 1 9 7 1 9 16 15 13 10 9 3 0 7 9 1 13 3 9 1 9 7 9 1 15 16 13 2
22 7 3 16 10 9 11 4 13 16 15 3 13 13 9 2 11 3 4 13 15 0 2
17 10 9 0 7 9 1 9 0 2 15 15 13 1 9 7 9 2
15 15 3 4 4 13 1 10 9 1 13 7 9 1 9 2
17 10 9 4 13 1 10 9 11 2 10 9 11 7 10 9 11 2
61 10 9 0 3 4 13 15 1 10 12 7 12 9 8 2 10 16 3 13 4 13 15 1 10 9 0 13 2 7 13 15 2 1 9 1 9 1 13 10 9 1 10 9 2 16 13 1 10 9 10 9 16 15 13 10 0 9 7 9 0 2
31 10 9 13 12 1 10 12 9 1 10 11 1 11 1 10 11 2 8 2 7 10 11 1 11 2 1 11 11 11 2 2
36 10 9 13 13 2 10 9 1 11 11 15 9 1 10 11 1 10 11 2 11 7 10 9 4 13 1 11 2 13 10 9 1 13 10 9 2
20 10 9 2 3 13 1 10 9 7 10 9 0 2 4 13 7 13 1 12 2
27 11 11 3 13 10 9 0 1 11 7 11 2 7 15 3 13 13 16 3 13 9 7 9 1 10 9 2
28 16 4 13 15 9 16 13 10 9 3 0 8 9 3 0 16 15 4 13 1 11 2 10 9 13 3 0 2
22 10 9 1 10 9 13 13 3 10 0 9 1 10 9 0 1 10 9 1 10 11 2
19 13 3 1 11 2 7 16 4 13 3 13 16 15 13 3 10 9 3 2
11 3 2 13 10 9 1 12 9 1 11 2
25 3 1 12 9 1 9 1 9 1 11 2 11 7 11 11 4 13 1 10 9 1 10 9 0 2
15 2 15 13 11 1 10 11 11 1 11 7 3 1 9 2
41 11 11 13 10 9 13 1 9 0 7 0 2 0 1 10 9 0 11 2 9 2 2 11 11 2 2 13 1 10 9 2 9 7 9 1 9 0 0 7 0 2
12 1 9 1 10 9 12 2 10 9 0 13 2
62 10 9 0 2 10 9 0 13 12 1 10 12 9 16 13 9 1 9 1 11 7 11 2 12 1 10 9 2 1 10 0 9 7 3 13 10 9 1 10 9 16 13 10 9 2 16 13 10 9 1 9 1 11 1 11 7 11 2 11 7 11 2
31 10 9 15 15 13 15 7 13 0 2 3 4 13 15 0 7 0 2 10 9 7 15 15 4 13 10 15 16 4 13 2
48 9 1 10 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2
13 1 10 9 9 0 13 1 12 9 1 12 8 2
6 13 0 1 10 9 2
31 10 11 11 2 8 11 13 10 9 1 9 0 1 10 9 1 11 2 13 1 12 1 10 9 0 1 10 11 11 11 2
39 13 10 9 0 1 10 2 9 1 9 2 1 10 15 10 9 15 13 16 13 1 10 9 10 9 16 3 13 1 10 9 1 10 9 7 1 10 9 2
62 10 9 1 10 9 13 10 9 1 10 9 0 16 13 10 9 1 9 1 10 9 1 10 9 2 16 3 4 13 10 9 7 10 9 0 1 10 9 2 1 10 10 9 16 15 13 1 10 9 1 9 7 16 13 1 10 9 1 10 9 13 2
25 11 11 7 11 3 4 3 13 7 10 9 1 10 9 13 1 10 9 7 9 0 1 10 9 2
15 10 9 13 10 9 7 9 1 10 9 1 10 0 9 2
14 4 13 0 1 10 9 1 9 1 11 9 2 12 2
15 10 12 1 11 1 12 2 15 4 13 1 10 9 0 2
39 10 9 13 10 0 9 1 12 9 1 9 2 7 1 15 15 13 10 9 0 1 9 0 16 15 13 1 10 0 9 0 0 1 0 9 0 7 0 2
40 1 11 15 13 2 0 1 11 11 2 10 12 9 9 7 0 1 9 0 2 1 10 12 11 2 10 9 0 9 16 13 1 11 2 3 4 13 9 0 2
30 4 13 3 1 12 9 1 10 9 2 7 13 3 10 11 1 10 9 1 9 1 11 11 11 12 2 10 11 11 2
17 13 10 9 1 9 1 12 2 13 15 1 9 0 7 9 0 2
40 1 10 9 13 1 9 11 11 11 2 15 13 10 9 1 9 1 10 9 8 7 10 9 1 9 1 10 8 2 16 7 10 11 13 10 0 9 1 8 2
21 1 10 0 9 15 13 3 9 1 9 8 7 0 1 11 1 11 2 8 2 2
22 1 12 9 13 12 1 11 2 9 1 10 9 1 3 1 10 0 11 11 2 12 2
18 1 0 2 11 3 4 13 1 9 1 10 9 3 1 10 0 9 2
49 10 11 13 4 15 13 1 10 11 11 7 10 9 15 13 1 10 9 1 11 16 13 10 9 16 13 7 13 16 10 9 1 1 11 15 13 10 9 16 15 13 13 15 1 10 9 3 0 2
25 10 9 3 13 1 9 1 0 8 0 2 7 3 13 10 9 1 15 3 7 15 3 7 11 2
26 1 12 2 10 9 12 1 10 9 1 9 1 10 11 11 15 13 1 10 9 0 1 10 9 0 2
30 3 1 10 9 2 0 7 13 1 10 10 9 2 10 9 1 10 9 2 1 10 9 0 2 0 2 13 3 0 2
23 10 9 1 10 9 11 11 11 4 13 1 13 1 10 9 0 1 16 13 1 10 9 2
42 1 9 1 10 9 1 10 9 7 1 10 10 9 1 11 0 1 10 9 2 10 9 3 13 13 7 13 2 7 3 13 10 9 0 1 10 9 0 7 3 0 2
23 10 9 0 13 10 9 3 3 2 10 9 11 15 13 1 11 9 13 3 1 12 9 2
56 10 11 1 11 7 11 2 11 2 4 13 16 10 9 13 1 10 9 1 13 10 9 13 3 9 2 10 12 5 2 7 10 3 9 2 12 5 2 2 1 10 9 13 1 3 1 12 9 1 12 9 1 10 10 9 2
17 11 13 13 10 9 1 9 0 2 1 10 2 9 2 1 15 2
20 11 11 2 1 10 9 11 11 2 13 1 10 9 1 10 9 1 10 9 2
7 9 2 9 7 9 0 2
11 3 15 3 13 9 1 9 16 13 15 2
11 13 16 15 13 10 11 11 1 10 11 2
19 13 1 10 9 2 13 2 7 13 3 1 12 9 2 13 1 0 9 2
20 10 9 13 1 9 0 7 2 1 9 2 3 0 1 10 9 1 9 0 2
9 4 13 9 16 15 4 13 15 2
35 1 10 9 10 9 13 10 9 0 2 1 9 2 15 13 0 0 9 1 10 0 9 2 13 1 10 9 1 9 7 1 10 9 0 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
12 11 11 13 10 9 1 9 1 10 9 11 2
26 10 9 15 4 13 1 10 0 2 8 8 2 16 13 1 10 9 1 10 9 1 9 1 10 9 2
20 13 10 9 1 10 9 0 13 1 10 9 2 10 3 9 11 11 1 11 2
9 15 13 1 13 1 9 1 11 2
22 4 13 0 1 10 11 11 2 12 1 11 2 13 12 9 7 13 10 9 1 11 2
42 15 13 1 15 0 1 9 1 9 3 7 1 9 2 13 10 9 1 9 1 12 9 1 9 2 13 1 10 9 0 7 13 1 11 11 2 3 9 0 1 9 2
15 1 10 9 11 2 10 9 13 1 10 9 10 1 11 2
39 10 11 2 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 1 11 7 11 2 1 10 9 1 9 7 9 1 10 11 2 1 2 11 2
28 15 13 3 0 16 10 9 2 13 8 2 3 1 10 9 1 12 1 12 3 1 10 11 7 10 9 11 2
29 1 13 10 9 11 1 10 0 9 7 13 10 11 11 1 10 9 4 13 10 9 16 4 13 13 1 10 9 2
15 13 16 13 3 10 9 1 10 9 0 1 9 1 9 2
67 1 0 9 2 9 0 2 11 7 1 9 0 2 13 1 10 9 0 2 11 2 11 2 11 11 1 11 2 11 2 11 8 2 1 10 13 9 1 11 1 12 1 10 9 1 11 11 2 5 5 11 1 11 7 1 11 9 1 10 9 1 11 2 9 1 11 2
16 10 9 13 3 0 1 9 9 1 10 9 5 7 11 11 2
17 1 9 1 10 9 13 10 9 9 16 13 10 9 7 13 9 2
37 10 2 11 1 10 11 2 13 1 15 2 4 13 3 1 10 9 0 2 1 15 11 2 7 3 1 10 9 1 10 9 2 1 15 11 11 2
10 11 13 16 15 13 1 10 9 12 2
30 10 9 4 13 3 10 9 1 10 9 1 10 9 0 2 16 10 9 4 13 1 12 9 1 12 9 0 10 15 2
35 10 9 7 10 9 4 13 1 9 1 10 9 16 13 1 10 9 0 1 10 9 1 10 9 2 16 13 2 2 16 13 10 9 0 2
25 11 13 15 1 10 9 1 0 9 1 10 9 0 1 10 9 0 2 0 1 10 9 1 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
54 16 1 15 15 13 13 15 2 13 10 9 3 1 15 9 2 15 13 10 9 0 7 0 7 3 13 10 9 7 9 16 3 15 13 2 0 2 1 10 9 13 15 1 4 13 1 2 9 0 2 7 4 13 2
40 10 11 2 7 11 2 13 10 9 13 1 10 9 0 13 1 10 9 1 10 9 0 7 0 1 10 9 0 1 11 2 1 10 9 1 10 11 11 11 2
42 1 10 9 3 0 13 10 2 9 2 7 2 11 2 2 10 9 2 9 1 9 0 2 10 9 0 7 13 1 9 2 3 10 9 2 7 10 9 1 9 0 2
17 16 10 9 13 1 10 9 2 15 3 15 13 2 3 3 2 2
33 10 9 1 10 9 15 13 8 2 3 1 13 1 11 1 10 9 1 10 9 1 11 1 12 2 16 4 13 1 10 11 11 2
32 13 9 1 10 9 11 11 2 9 1 10 11 1 10 11 2 13 1 10 9 7 16 4 13 9 0 1 13 10 9 0 2
24 10 9 1 10 9 1 9 0 1 11 11 1 11 13 9 0 1 10 0 9 1 10 9 2
31 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
14 10 9 2 11 2 4 13 1 11 11 7 11 11 2
50 15 13 1 10 9 4 13 1 10 9 11 12 2 1 10 9 15 15 4 13 16 13 1 10 9 1 11 1 11 7 1 11 9 1 10 9 13 1 15 16 13 10 9 1 9 13 1 10 9 2
20 1 3 10 10 9 0 2 1 10 9 2 13 0 10 9 1 10 9 0 2
22 1 10 9 15 13 10 9 13 1 10 9 1 9 2 9 2 9 2 9 7 9 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
71 1 13 15 10 9 1 11 12 7 10 9 1 10 9 1 11 12 1 11 2 10 9 0 13 10 9 1 11 1 10 9 1 10 0 9 2 10 9 11 12 1 11 2 16 13 1 10 9 2 1 10 9 0 7 0 1 10 11 9 1 10 9 1 10 9 11 1 10 9 0 2
17 11 4 3 13 1 15 1 10 12 9 0 3 0 1 10 9 2
35 13 0 2 3 7 4 1 13 15 3 9 1 10 9 1 9 2 4 7 13 1 12 9 10 9 2 7 10 16 13 1 16 4 13 2
8 13 10 9 1 10 9 0 2
35 10 9 0 13 10 9 1 11 11 2 11 7 10 9 1 10 11 1 11 7 13 1 11 1 10 9 0 1 11 1 10 9 1 12 2
19 3 13 9 1 10 9 1 2 11 0 2 2 12 2 2 1 11 11 2
10 10 0 9 13 10 9 11 11 11 2
18 4 13 7 15 4 13 10 9 0 1 9 1 9 0 1 10 9 2
58 15 1 10 9 7 1 10 9 13 1 10 9 2 13 13 3 1 10 9 2 3 16 13 1 15 2 7 16 10 9 15 13 1 9 1 10 9 2 1 4 13 1 9 2 1 10 0 9 1 10 9 0 2 1 10 9 0 2
50 10 9 11 1 9 12 2 16 4 13 1 11 1 12 9 2 13 10 2 0 9 2 9 7 9 2 16 13 1 10 9 0 7 13 16 2 1 10 9 7 10 9 2 15 13 1 10 9 2 2
51 3 1 16 13 10 9 8 2 11 13 10 9 1 12 9 2 11 11 2 16 15 13 1 10 11 1 11 2 2 11 11 2 16 15 13 1 10 11 2 7 11 11 2 15 15 13 1 10 11 2 2
18 15 13 0 1 10 9 1 9 1 10 9 1 11 2 11 7 11 2
37 1 10 9 2 11 11 12 2 11 13 9 1 9 1 11 2 1 15 1 11 1 10 12 5 2 11 1 10 12 5 7 11 1 10 12 5 2
12 10 9 1 11 11 15 13 0 1 10 9 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
18 1 10 9 15 15 13 1 9 2 10 9 13 3 12 12 1 9 2
10 13 3 1 10 9 10 9 11 11 2
35 10 9 0 0 13 9 1 9 2 11 2 2 1 10 9 0 9 2 9 2 16 4 13 15 1 9 1 9 1 9 1 10 9 0 2
14 10 9 13 15 0 2 16 15 13 3 1 0 9 2
15 13 10 9 1 10 9 2 7 10 9 0 13 3 0 2
10 4 7 13 3 15 13 3 10 9 2
47 13 12 9 2 1 10 15 12 13 1 10 9 1 11 2 7 1 10 15 12 2 10 3 9 2 11 11 2 13 1 11 0 2 7 10 3 9 7 3 0 2 11 11 2 1 11 2
16 10 9 13 10 9 1 10 0 9 0 7 0 1 10 9 2
31 10 9 13 10 9 0 1 10 9 3 0 1 10 9 0 2 2 3 13 2 3 1 13 7 1 15 15 13 2 9 2
28 2 13 10 9 2 4 13 10 9 0 7 3 3 13 10 9 2 4 1 4 13 15 2 2 13 10 9 2
8 11 15 13 13 1 10 9 2
23 13 10 9 1 9 1 10 0 9 2 1 11 11 11 15 13 10 9 16 3 4 13 2
25 10 11 2 10 11 2 13 10 9 0 1 10 9 1 9 0 9 13 1 11 1 12 7 12 2
39 10 9 13 10 9 3 0 2 10 9 3 0 7 10 9 3 0 2 3 15 9 13 1 10 9 2 16 13 10 9 15 13 10 9 1 10 9 0 2
18 11 13 10 9 1 10 9 1 11 1 10 11 1 11 2 1 11 2
15 10 9 4 4 13 7 0 9 4 4 13 1 10 9 2
31 10 0 9 1 10 9 2 2 8 8 2 2 13 13 1 11 2 11 2 11 7 11 11 2 7 13 3 1 9 0 2
20 3 13 10 9 1 10 9 1 10 9 11 2 11 2 16 13 15 1 15 2
34 10 9 4 13 13 1 11 11 2 1 9 1 10 9 16 15 4 13 1 10 9 1 10 9 2 7 16 4 13 10 9 1 11 2
31 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 9 12 2 7 10 9 0 1 9 13 9 12 2
35 10 9 13 1 10 9 0 16 10 9 0 13 10 11 1 10 9 0 16 12 9 13 10 9 0 1 10 9 2 16 13 9 7 9 2
25 1 10 0 9 15 13 1 10 9 10 11 11 1 11 2 1 15 13 1 12 1 10 0 9 2
12 13 10 10 9 7 11 7 11 1 10 9 2
12 15 4 13 1 12 9 7 3 15 13 13 2
15 2 1 9 10 10 9 4 13 1 10 9 0 2 13 2
31 10 0 9 1 9 13 16 2 10 9 0 4 13 10 9 2 7 13 1 16 2 10 9 13 0 1 10 12 5 2 2
22 15 13 3 1 11 11 2 11 11 11 2 11 11 2 11 11 7 11 11 1 9 2
4 13 1 11 2
14 13 3 1 16 10 9 13 1 10 11 12 1 12 2
6 1 12 13 10 9 2
31 10 9 0 13 1 10 11 16 13 1 10 10 9 0 1 10 9 16 13 0 16 13 11 2 1 9 7 1 10 9 2
18 1 10 9 10 9 1 10 9 13 0 13 10 0 9 1 9 0 2
42 10 9 0 4 1 4 13 1 9 1 2 9 12 2 2 13 10 9 0 1 10 9 12 5 7 12 5 7 10 9 1 10 9 1 0 9 0 1 10 0 9 2
21 10 11 1 10 11 2 11 2 15 13 1 11 1 11 10 10 9 3 1 11 2
38 12 9 1 10 16 11 1 10 11 11 2 11 2 3 4 4 1 13 16 13 7 13 10 9 1 9 16 10 9 13 1 10 9 1 9 1 9 2
21 1 9 15 13 10 9 1 10 9 1 10 9 13 1 11 1 12 2 13 3 2
11 15 13 3 11 7 3 10 9 11 11 2
14 10 9 13 3 0 7 15 13 3 15 10 9 0 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
16 13 10 9 1 11 7 1 10 11 11 1 10 11 1 11 2
19 11 11 13 10 9 1 9 0 1 10 9 11 1 10 9 1 10 11 2
37 1 10 9 1 2 11 11 11 11 11 11 11 2 2 10 9 13 1 11 11 11 1 10 9 12 1 9 1 12 9 3 15 13 1 12 9 2
23 11 11 2 11 11 2 2 13 1 11 2 13 1 10 9 1 11 11 2 2 15 13 2
18 11 13 15 1 10 9 3 0 1 10 9 12 3 1 10 9 0 2
51 16 13 1 10 9 1 10 9 0 11 15 13 2 1 9 2 1 10 0 9 1 11 1 11 7 11 11 1 11 1 10 9 16 13 10 9 3 0 1 10 9 2 1 10 9 1 9 1 10 9 2
30 1 9 4 13 15 7 1 0 9 1 9 1 9 2 0 9 2 7 15 13 0 3 16 15 13 9 1 9 0 2
11 11 11 13 10 9 0 1 10 9 11 2
27 2 13 16 0 1 10 11 1 10 11 2 9 4 13 11 1 10 9 0 2 2 13 11 11 1 11 2
45 11 11 3 15 13 1 9 0 2 3 10 9 15 13 10 11 11 2 16 13 9 1 10 9 11 2 3 1 9 1 9 2 1 10 16 10 9 4 13 0 1 10 0 9 2
8 10 9 2 13 7 3 13 2
21 3 1 10 9 1 9 2 10 8 2 9 13 13 9 7 13 15 1 9 0 2
24 10 9 1 10 9 13 10 9 1 10 9 16 13 1 10 9 7 10 9 1 10 9 0 2
21 16 13 2 13 1 10 9 1 9 1 9 1 10 9 15 10 9 11 15 13 2
41 3 13 9 1 10 0 9 13 10 9 2 1 15 16 13 1 3 7 9 1 9 2 16 15 9 16 13 13 16 15 13 10 9 3 7 13 15 1 10 9 2
48 13 10 12 1 11 1 12 1 11 2 3 10 12 11 15 13 1 10 11 11 2 1 11 10 12 1 11 1 12 2 1 11 11 1 11 12 7 16 13 1 11 10 12 1 11 1 12 2
35 1 12 1 9 1 10 9 2 8 4 13 2 11 11 2 1 12 5 11 2 13 1 15 11 7 11 1 11 1 10 11 11 11 11 2
33 10 9 13 1 13 10 9 1 10 9 2 13 15 10 9 2 13 15 10 9 7 13 15 1 13 10 9 1 10 9 1 9 2
12 1 13 10 9 13 1 9 1 10 9 0 2
59 11 13 1 10 0 9 0 13 1 9 0 2 16 13 1 13 10 9 0 1 10 9 16 13 3 10 12 9 1 9 2 4 13 10 9 15 0 1 9 2 9 1 0 9 7 10 9 16 1 10 9 15 7 3 10 9 4 13 8
27 10 9 13 10 9 3 0 1 10 9 2 10 9 0 13 1 12 11 11 2 15 1 12 7 1 12 2
53 10 11 13 0 10 9 2 10 9 1 11 2 10 9 16 3 13 1 10 9 1 10 11 7 13 15 1 10 9 1 11 2 3 1 11 2 15 15 4 13 0 1 15 1 10 9 16 3 13 1 11 11 2
9 10 9 0 15 13 1 12 9 2
11 10 9 13 0 7 10 9 13 3 0 2
46 1 9 1 13 1 10 3 8 1 10 9 2 15 13 1 10 9 10 9 4 13 10 9 1 3 12 9 1 10 9 16 15 13 0 1 10 9 1 10 9 1 9 1 9 0 2
26 11 11 11 11 2 2 12 1 11 1 12 2 11 1 11 2 9 1 11 2 2 13 10 9 0 2
3 11 11 2
19 11 13 9 1 10 9 1 11 12 2 3 1 9 1 10 9 0 11 2
52 1 10 9 10 9 1 11 11 3 13 10 9 1 9 0 1 10 9 0 9 2 13 1 10 9 15 11 11 13 1 15 1 10 0 9 1 10 9 1 15 16 3 3 13 11 1 10 11 1 10 11 2
56 1 10 9 11 3 13 10 0 9 0 16 13 1 10 9 0 1 13 12 5 2 10 15 15 13 1 9 1 10 9 1 10 9 2 10 15 13 10 9 1 10 9 2 15 15 13 10 9 1 9 1 11 1 10 9 2
9 13 1 10 9 1 11 7 11 2
8 10 9 13 10 9 1 9 2
18 10 0 9 13 1 9 13 11 11 2 11 11 7 11 11 2 11 2
19 3 1 10 9 0 2 10 9 1 11 7 9 13 0 9 1 10 9 2
50 2 13 0 13 15 15 1 10 9 2 7 13 3 0 13 15 16 10 9 2 7 11 7 11 13 2 16 3 13 10 0 9 7 3 15 4 1 13 2 2 13 11 11 11 2 9 1 10 9 2
51 10 9 1 9 1 10 11 11 13 3 1 9 0 1 9 1 10 9 13 1 9 13 1 10 9 7 3 13 1 10 9 1 10 11 1 10 11 1 10 11 11 2 11 11 1 11 1 11 7 11 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
22 1 13 10 9 2 11 2 9 1 11 2 4 13 1 9 1 11 2 9 1 11 2
25 10 9 0 13 10 9 1 10 9 1 11 11 1 11 15 4 4 13 1 10 9 0 9 3 2
50 1 12 2 10 9 13 10 0 9 2 1 0 9 1 10 9 1 10 9 2 12 9 13 1 12 13 2 9 1 11 1 11 2 9 1 11 1 11 11 2 7 3 4 13 1 10 9 1 9 2
8 1 10 9 4 13 12 9 2
14 10 9 15 13 1 12 1 10 9 1 11 11 11 2
30 15 4 13 1 10 9 1 10 9 1 11 11 1 12 2 1 9 1 11 2 11 7 11 2 11 11 7 1 12 2
10 7 9 13 9 7 1 9 9 0 2
9 4 13 1 10 11 11 1 11 2
12 10 0 9 13 1 10 9 3 0 1 11 2
31 16 13 11 11 2 1 11 10 9 3 4 13 1 10 9 0 0 2 7 1 10 9 1 9 1 10 2 9 0 2 2
36 1 12 2 13 1 10 11 11 1 3 3 15 13 0 13 10 9 1 9 1 9 2 7 13 13 7 15 4 1 13 1 10 9 0 0 2
69 11 13 10 9 0 1 10 9 1 10 9 1 9 1 10 9 7 1 10 9 1 9 16 4 1 4 13 1 3 1 12 9 1 10 12 9 16 13 10 9 2 12 1 11 1 12 1 11 2 2 13 1 10 9 10 9 1 0 16 4 13 10 9 1 10 9 1 9 2
28 1 10 9 13 1 13 1 11 7 1 11 2 3 13 1 10 9 1 10 11 11 2 9 1 10 11 11 12
19 10 9 13 1 10 9 1 10 9 1 11 11 11 13 1 10 12 5 2
27 10 9 4 13 0 9 1 9 1 10 9 1 9 1 11 11 11 3 1 10 9 0 1 10 9 1 9
55 11 2 11 11 2 2 11 2 11 11 2 7 11 2 11 11 2 13 10 9 1 10 9 1 11 11 1 10 9 13 10 11 11 2 15 2 3 1 9 2 13 10 9 1 9 1 16 10 9 4 13 1 10 9 2
13 13 10 9 1 10 9 1 11 2 11 11 2 2
36 7 3 1 4 15 13 2 13 10 9 1 13 1 10 9 7 0 9 1 11 11 2 11 2 13 1 13 1 10 9 7 1 9 0 0 2
38 13 15 1 10 9 3 0 2 13 10 9 1 9 1 3 1 10 12 5 8 2 3 1 12 5 8 2 2 16 13 9 3 0 1 10 0 9 2
10 13 9 1 11 10 12 1 11 1 12
8 11 15 13 13 1 10 9 2
29 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 2 1 10 15 13 1 9 0 7 13 9 2
32 1 10 12 13 1 10 9 11 1 10 9 11 7 1 10 9 1 9 11 11 11 1 11 11 2 3 13 0 1 11 11 2
23 10 0 9 0 2 13 0 2 16 13 10 9 2 0 1 10 9 1 9 1 9 0 2
24 11 11 11 15 13 10 9 1 10 9 1 9 1 10 8 2 9 13 1 2 11 2 2 2
13 11 4 4 3 3 13 1 10 9 1 10 9 2
34 1 10 9 4 13 13 4 13 1 10 11 11 2 1 9 1 0 9 1 10 9 11 11 11 2 1 10 9 1 11 11 1 11 2
49 10 9 1 10 9 13 3 0 2 7 10 9 3 13 10 9 0 13 1 16 13 1 10 9 1 11 11 2 1 15 7 15 13 10 9 1 10 9 13 15 1 13 11 11 12 1 11 11 2
8 12 9 0 13 1 10 9 2
14 15 13 1 10 9 11 11 10 12 1 11 1 12 2
40 1 11 1 10 0 9 4 13 1 0 9 1 10 9 0 1 9 1 9 1 10 9 2 9 15 4 1 13 1 11 7 1 11 1 12 1 10 0 9 2
9 11 11 7 11 13 10 9 0 2
23 10 9 0 11 11 2 16 13 1 9 1 11 2 15 13 13 10 9 1 11 7 11 2
15 3 13 1 10 11 11 7 3 1 10 9 1 11 11 2
59 10 0 9 1 10 9 1 9 0 16 13 1 12 9 1 11 13 9 1 10 3 1 12 9 7 9 16 13 1 10 9 2 10 11 11 11 7 11 7 10 11 11 2 9 0 2 13 1 10 11 1 11 7 1 11 1 10 9 2
11 15 9 0 4 13 7 13 1 10 9 2
33 10 9 16 13 16 11 13 0 1 10 9 0 0 13 10 9 0 7 10 12 9 0 2 16 13 12 0 9 7 9 1 9 2
6 10 9 13 0 9 2
24 1 10 9 9 12 1 10 9 0 1 0 9 13 1 10 11 1 11 2 3 1 8 9 2
21 13 9 1 10 9 0 1 9 1 10 9 1 1 10 9 12 1 10 9 12 2
31 1 9 1 10 11 11 11 2 11 11 13 10 9 1 10 9 1 12 9 1 9 0 1 13 10 9 1 10 11 11 2
26 1 10 9 1 11 2 11 7 11 2 10 9 12 4 13 10 9 1 13 15 0 1 10 9 11 2
28 2 11 11 11 2 11 11 11 2 10 11 11 11 11 11 2 11 2 11 11 11 11 2 12 2 11 2 12
38 1 10 12 11 2 11 11 2 12 4 13 1 10 11 11 11 2 10 11 2 11 12 7 11 2 11 12 13 10 9 11 2 12 7 11 2 12 2
17 1 10 9 15 15 13 8 8 8 2 2 2 16 13 9 2 2
21 10 9 15 13 1 10 12 8 2 7 13 3 1 12 5 5 1 9 0 0 2
21 10 9 11 11 11 13 3 0 7 13 9 1 9 1 3 1 12 9 1 11 2
38 15 13 9 1 10 9 1 10 9 0 2 1 10 9 2 1 10 9 0 1 10 9 2 1 10 9 2 2 3 13 8 13 0 1 13 10 9 2
43 10 11 0 2 1 3 12 9 2 15 13 1 10 9 0 1 10 9 0 7 0 0 11 2 1 10 9 1 10 16 10 9 0 2 0 13 15 1 10 9 3 0 2
29 1 11 11 2 4 13 1 12 10 0 9 1 9 0 7 13 3 1 12 9 1 9 2 16 13 10 9 0 2
33 13 9 1 10 9 2 1 10 9 1 10 9 2 7 3 1 10 9 4 13 1 9 1 10 11 1 11 2 16 15 3 13 2
49 1 10 9 2 13 13 1 10 9 1 10 9 1 10 9 0 1 10 13 16 16 3 2 13 3 10 9 0 1 9 2 1 10 9 15 13 1 10 9 1 12 7 12 9 1 13 9 2 2
66 15 13 10 9 1 9 2 1 15 13 16 10 9 0 2 0 2 7 0 0 1 10 9 1 9 3 13 9 7 1 10 9 7 1 10 9 2 1 13 2 1 9 2 9 16 13 10 9 1 10 9 2 1 10 9 2 10 9 2 10 9 1 9 2 8 2
29 11 2 10 9 1 11 3 4 13 0 9 7 15 15 13 1 10 9 2 7 15 3 13 9 0 1 10 9 2
35 1 11 2 15 1 10 0 9 0 13 1 13 1 10 9 1 10 11 1 11 2 3 15 13 9 1 10 9 13 1 2 11 0 2 2
24 11 11 11 13 10 9 0 1 10 9 1 10 9 1 10 9 1 11 11 1 10 9 0 2
38 13 9 1 0 9 1 9 0 7 0 1 10 15 15 13 2 11 7 11 1 11 2 2 3 13 1 10 9 0 7 13 10 9 1 10 9 0 2
17 11 13 12 9 1 10 9 0 0 0 2 3 1 10 9 0 2
6 9 0 2 11 11 2
31 11 11 13 16 13 1 10 0 9 0 1 10 0 9 2 15 15 4 13 16 10 9 1 9 1 11 4 13 10 9 2
13 1 10 9 13 13 1 10 9 1 10 0 9 2
28 10 9 3 13 2 1 10 9 2 1 10 10 0 9 0 7 0 1 10 9 2 16 13 1 9 9 0 2
40 1 9 2 10 9 0 15 13 1 10 9 13 1 10 9 1 0 9 1 10 9 1 9 2 9 7 9 2 0 1 10 7 9 9 2 9 1 9 2 2
56 2 11 15 1 10 9 2 15 13 9 1 9 7 9 1 10 9 2 16 2 1 9 1 10 9 13 2 13 7 13 10 9 0 2 10 9 0 2 10 9 0 2 0 2 0 7 0 16 13 10 9 2 2 15 13 2
16 10 11 11 15 13 1 10 9 7 4 13 1 9 1 9 2
21 10 9 13 10 9 1 11 2 10 9 0 16 13 1 10 0 9 7 10 9 2
63 1 10 9 4 13 9 1 10 9 1 10 11 1 9 1 9 0 1 10 9 13 10 9 3 0 2 1 9 1 10 9 1 11 2 1 10 9 1 9 1 10 9 2 1 10 9 1 11 11 2 7 13 10 9 0 1 11 2 10 11 7 11 2
30 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 7 9 2 1 10 9 1 11 7 9 1 11 2
27 10 9 15 13 7 2 0 1 10 9 11 2 16 13 10 9 1 9 2 13 10 9 1 10 9 0 2
16 1 12 10 11 11 13 10 11 11 8 11 11 1 10 9 2
33 1 10 9 2 10 9 1 11 13 10 9 1 11 1 11 2 1 15 15 10 9 2 1 9 13 1 9 2 15 13 1 11 2
41 1 9 1 9 3 2 11 13 3 1 10 9 0 1 10 9 7 15 13 16 13 10 9 16 15 13 13 10 0 9 1 10 9 16 3 13 1 13 1 9 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
52 10 9 1 11 11 11 13 4 13 10 9 2 0 1 15 3 16 13 1 10 9 2 1 10 0 9 2 15 13 4 13 9 1 15 10 9 1 10 0 8 1 11 11 2 3 13 1 10 9 1 11 2
33 10 12 11 11 11 1 11 2 13 15 1 10 12 11 11 11 1 15 15 13 0 11 7 15 1 10 12 1 10 9 1 11 2
26 1 10 9 1 10 2 9 0 1 9 2 2 1 10 9 12 10 9 1 10 9 13 10 12 9 2
56 16 10 9 0 11 11 13 13 10 9 1 10 9 1 11 2 1 10 9 11 12 2 10 9 13 1 10 9 0 13 10 9 1 10 9 0 1 1 10 9 11 12 13 1 11 12 1 13 9 0 1 13 1 10 9 2
13 10 9 0 2 11 2 13 10 9 1 10 9 2
25 10 9 0 15 13 10 11 1 10 11 11 13 0 1 13 1 10 9 0 7 0 2 13 1 2
55 1 4 13 1 10 9 2 1 10 9 13 1 10 9 2 10 9 1 10 11 2 1 10 3 16 10 1 10 9 2 9 7 9 13 0 1 10 9 2 13 10 9 0 2 9 7 9 1 10 9 0 1 10 9 2
12 13 16 16 13 1 10 9 10 9 13 0 2
12 13 1 13 1 11 3 1 4 1 13 9 2
55 10 9 1 10 9 1 11 11 2 11 2 9 7 11 7 1 10 0 9 0 3 0 1 11 1 10 9 1 10 9 1 9 1 10 9 7 9 0 4 13 1 10 9 7 9 10 9 0 3 0 7 1 0 9 2
31 11 11 11 4 13 10 9 1 10 9 11 7 13 10 9 9 1 13 1 10 11 0 1 10 9 1 10 11 11 11 2
72 3 2 16 15 13 10 9 1 9 7 3 15 13 10 9 16 3 13 1 10 9 2 3 15 13 10 9 2 7 10 9 13 16 2 13 10 9 2 10 9 13 1 13 1 10 9 2 1 9 16 10 0 9 3 3 4 13 15 2 16 2 1 9 2 4 13 1 13 10 9 2 2
56 1 9 2 1 10 12 2 11 4 13 1 10 0 9 2 13 1 9 12 1 12 2 13 10 9 0 7 13 3 9 0 7 9 2 1 10 9 1 13 9 1 0 9 0 0 7 13 0 10 9 1 10 9 1 15 2
19 10 9 13 10 9 1 15 13 3 2 1 9 0 2 1 10 9 0 2
14 4 13 1 9 16 13 10 9 1 10 9 0 11 2
10 10 9 13 3 10 9 16 10 9 2
20 13 1 9 7 10 0 9 13 10 11 11 11 11 1 10 0 11 1 11 2
8 15 13 1 10 9 1 9 2
37 13 0 1 11 1 10 9 1 12 9 2 13 3 10 9 13 1 9 7 13 10 0 9 1 15 15 15 13 10 9 1 10 11 1 11 0 2
11 10 12 9 4 13 1 10 9 1 9 2
30 13 1 13 1 9 2 9 2 9 7 9 1 10 9 1 13 9 0 2 3 1 10 9 1 10 9 7 10 9 2
19 15 2 3 2 13 1 15 15 15 13 13 1 10 9 7 1 10 9 2
14 15 13 16 13 10 9 1 10 12 16 3 4 13 2
17 10 11 13 12 5 12 8 9 9 7 12 5 12 8 9 9 2
53 1 10 9 1 10 9 2 13 0 9 0 2 1 15 2 1 10 9 1 9 7 9 1 10 9 16 15 13 13 2 11 1 10 11 11 2 2 15 13 13 10 9 16 3 15 4 13 1 9 1 10 9 2
17 10 9 2 3 0 2 15 13 0 1 10 9 1 10 9 0 2
41 1 13 15 1 10 15 4 13 10 11 11 16 2 1 13 15 2 13 9 0 2 7 1 9 7 1 9 2 16 13 16 15 15 13 1 10 9 7 15 13 2
27 10 9 2 1 10 9 11 2 13 9 2 9 0 16 13 10 9 0 1 10 9 2 3 10 9 0 2
27 1 9 2 4 13 10 9 0 1 10 11 11 1 10 11 1 10 11 2 11 1 10 9 1 9 2 2
11 10 9 4 13 15 3 0 7 10 9 2
21 11 3 13 10 9 1 13 10 9 1 9 1 10 11 2 11 1 11 1 11 2
10 10 9 1 9 13 0 1 12 9 2
26 11 11 13 15 1 10 9 3 0 1 11 2 1 9 1 11 13 1 10 9 1 3 1 12 9 2
33 2 15 15 15 13 3 7 1 15 15 13 1 10 9 2 10 9 16 15 13 10 9 2 10 9 15 13 0 2 2 13 11 2
15 15 13 1 10 9 1 10 9 0 0 7 10 9 0 2
35 10 12 1 11 4 1 13 10 9 1 11 1 10 12 1 10 9 1 10 9 12 16 13 10 9 1 10 9 1 11 7 10 9 11 2
12 10 9 4 13 13 10 12 9 1 9 0 2
21 4 13 1 10 9 1 13 10 9 1 9 0 1 10 8 2 3 10 9 0 2
9 1 10 9 3 15 13 1 9 2
15 10 9 4 13 1 10 9 1 9 1 9 1 11 11 2
29 10 9 1 4 13 11 3 4 13 9 2 1 15 15 13 1 10 9 1 9 7 9 1 13 0 1 10 9 2
45 10 9 0 1 10 9 1 11 2 1 9 0 1 9 2 0 9 2 0 7 0 9 2 0 9 0 2 0 9 7 0 9 2 4 13 1 9 0 3 3 0 1 10 9 2
19 10 9 13 10 9 12 1 10 9 1 9 0 2 13 12 9 1 9 2
25 10 12 1 11 1 12 2 10 11 13 13 15 1 10 11 2 13 10 11 11 11 2 11 2 2
19 0 9 16 13 9 7 10 9 7 10 9 3 0 1 10 9 1 11 2
38 1 10 9 2 10 9 1 10 9 13 13 10 9 1 10 9 2 10 9 7 10 9 2 13 10 9 1 0 9 0 1 10 9 0 1 10 9 2
18 2 11 2 13 10 0 9 13 1 10 9 1 10 0 9 9 0 2
36 10 9 0 1 9 1 10 9 0 7 1 10 9 1 10 11 11 1 10 9 13 1 9 1 10 9 1 9 1 9 11 7 9 1 9 2
25 1 10 9 2 11 11 13 10 0 9 1 9 7 9 0 1 10 9 16 13 13 15 1 15 2
11 13 0 1 10 12 9 7 3 3 13 2
20 1 12 11 13 10 0 9 1 10 11 1 10 9 2 13 10 9 1 11 2
16 3 3 1 10 9 4 13 1 10 9 1 10 11 1 11 2
3 13 15 2
5 11 0 7 0 2
16 10 9 13 16 13 10 9 1 11 11 2 9 7 9 0 2
49 2 11 2 10 9 1 9 8 13 1 10 12 5 1 11 7 11 2 4 13 13 10 9 1 10 9 0 1 10 9 1 12 9 0 1 11 7 12 9 9 1 10 9 1 9 1 10 9 2
46 3 0 2 16 13 15 13 1 10 9 1 11 2 1 16 1 12 10 9 4 0 1 10 9 3 1 15 1 10 9 11 12 1 11 7 10 0 9 1 15 2 9 11 1 11 2
40 1 2 11 1 9 1 11 2 15 15 13 3 2 11 1 10 9 0 2 16 11 11 11 11 13 1 10 9 16 13 3 1 13 1 10 9 0 2 0 2
18 10 9 1 9 2 13 1 10 9 1 13 10 9 0 1 10 9 2
42 15 16 3 4 13 0 13 16 10 9 0 13 16 13 10 9 0 1 9 1 10 9 7 9 0 2 15 15 4 13 1 10 9 1 9 7 9 1 10 9 12 2
25 1 3 2 13 0 1 15 1 10 9 7 1 9 2 15 13 3 2 3 2 16 13 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
38 15 4 13 9 1 9 0 1 10 9 1 10 9 0 2 7 1 10 2 11 10 9 2 2 1 2 11 2 7 1 2 10 11 1 10 11 2 2
14 10 9 4 13 1 0 9 1 12 1 11 11 11 2
22 10 9 4 13 1 13 15 1 11 1 10 11 2 16 13 3 10 9 15 3 0 2
34 10 0 9 2 4 13 1 10 9 11 2 10 9 0 2 7 10 9 15 13 1 10 9 0 1 10 9 1 11 7 1 10 9 2
59 15 13 10 9 16 13 1 10 9 0 2 7 3 15 13 10 0 9 1 10 9 13 1 10 9 15 13 2 15 13 16 15 13 16 13 15 1 10 9 3 1 9 2 1 10 15 16 1 10 9 13 10 9 7 15 13 10 9 2
54 13 1 10 9 1 11 3 11 2 15 13 9 1 12 1 12 2 13 10 9 2 1 9 15 13 16 3 4 13 1 10 9 1 11 1 10 9 1 11 2 13 15 10 9 10 9 2 16 10 12 9 13 0 2
11 3 10 0 9 7 9 0 1 10 9 2
47 10 9 1 10 9 0 1 10 11 1 10 11 1 11 2 11 11 11 2 4 13 10 9 1 9 7 9 1 10 9 1 10 9 0 1 10 9 1 10 9 10 9 1 10 10 11 2
6 13 1 11 7 11 2
38 0 13 10 9 1 10 9 1 11 11 3 11 15 13 15 3 0 7 13 13 10 9 1 9 1 9 0 1 10 9 2 11 2 11 11 7 11 2
15 13 10 9 0 2 10 9 0 3 0 7 10 9 0 2
37 10 9 13 2 2 2 10 9 7 10 9 7 10 9 1 9 15 13 10 7 15 13 1 11 7 15 13 1 9 1 10 9 1 10 9 2 2
27 10 9 13 10 9 1 10 9 7 13 13 16 10 9 1 9 3 13 1 10 9 1 13 9 7 9 2
63 1 10 9 2 10 9 1 11 13 1 10 9 1 10 9 1 9 0 1 9 0 2 16 13 10 9 1 10 9 2 10 9 7 3 10 9 2 15 13 2 15 10 9 7 10 9 1 10 9 2 1 9 16 13 0 10 9 1 11 1 10 9 2
8 2 13 1 10 9 7 3 2
12 13 10 0 9 0 2 13 1 11 12 9 2
46 10 9 1 10 9 13 1 11 1 10 9 1 10 9 2 1 9 1 10 0 9 1 9 1 10 11 1 10 9 1 9 16 1 12 7 12 13 10 9 1 9 13 1 10 9 2
28 10 9 15 13 1 10 9 0 1 4 13 10 9 0 1 4 13 1 13 15 2 1 10 9 1 10 9 2
13 11 13 1 11 1 11 10 12 1 11 1 12 2
9 1 15 2 11 15 13 1 9 2
7 3 2 9 13 13 9 2
28 11 11 2 11 2 12 2 13 9 1 11 11 1 10 11 1 11 10 2 11 7 9 1 10 9 1 9 2
7 3 13 10 9 1 9 2
8 10 9 13 1 10 9 12 2
70 7 16 13 15 13 16 13 0 1 13 7 13 1 9 1 12 1 10 0 16 3 15 13 7 1 10 9 7 13 1 0 9 7 1 10 9 1 10 16 15 13 15 9 2 3 4 13 1 13 3 1 10 9 16 13 16 3 13 1 15 7 3 3 13 10 0 9 1 15 2
20 3 13 1 10 9 1 11 2 13 1 11 11 2 10 11 2 2 1 12 2
36 3 13 10 0 9 16 13 9 1 10 9 0 7 3 13 16 1 11 16 15 13 10 9 2 3 15 13 10 9 1 10 9 1 13 15 2
41 3 3 2 3 4 13 1 10 9 1 10 9 0 13 1 9 1 10 9 7 1 15 2 1 10 9 1 10 9 2 16 1 3 3 15 4 13 1 0 9 2
53 10 9 4 13 1 10 9 1 11 2 3 10 9 1 10 16 13 11 7 10 9 2 10 11 11 2 3 9 1 10 9 0 11 2 2 4 13 1 10 9 10 9 15 4 13 10 9 7 3 4 4 13 2
25 3 2 15 15 13 12 9 1 9 1 13 1 10 9 2 15 13 13 16 13 0 1 10 9 2
43 10 9 1 11 13 1 3 9 1 10 9 1 11 2 1 10 9 1 10 9 2 1 15 15 10 9 1 10 11 2 9 1 10 9 1 11 2 13 10 9 1 11 2
47 1 9 2 3 7 16 13 10 0 11 11 2 13 15 15 16 13 16 4 1 13 15 10 0 9 1 10 9 1 10 9 2 13 15 1 15 10 9 7 13 13 1 10 9 16 13 2
14 10 12 1 11 1 12 4 13 9 0 1 10 11 2
24 10 9 13 0 1 10 9 0 2 1 10 0 9 7 1 10 9 0 0 1 11 2 11 2
16 10 13 10 9 0 8 2 9 1 9 1 10 9 0 2 2
32 10 9 15 13 1 10 9 1 9 7 2 1 15 2 1 10 0 9 1 10 9 2 15 16 15 13 3 3 0 1 13 2
30 10 9 13 1 10 9 7 2 0 1 10 9 0 2 15 13 1 13 16 10 9 1 10 9 13 1 10 9 0 2
24 10 9 2 10 9 7 1 9 10 9 13 16 15 13 9 16 13 1 10 9 0 2 0 2
31 1 10 9 10 9 13 1 9 10 9 1 16 10 9 2 1 9 2 9 7 9 0 2 13 7 13 9 1 9 0 2
17 10 9 0 13 10 9 0 1 10 9 0 7 0 0 7 0 2
29 15 3 2 1 11 11 3 4 3 13 3 7 13 1 10 12 5 1 11 2 1 10 9 1 11 1 10 9 2
38 3 3 1 16 13 10 9 2 10 9 0 13 1 11 11 13 10 9 0 1 10 1 11 2 7 3 1 10 2 9 2 0 2 16 13 10 9 2
17 10 9 13 9 1 9 1 10 15 13 10 9 0 2 13 15 2
21 13 12 9 1 9 7 13 1 10 9 1 9 2 16 3 15 13 3 1 9 2
22 13 16 10 9 13 9 0 0 1 10 9 1 16 13 2 7 13 3 9 1 9 2
12 11 4 3 13 1 10 0 9 1 11 11 2
18 10 9 1 9 15 13 11 11 7 13 10 9 3 0 16 4 13 2
15 11 13 10 9 0 1 9 1 9 0 1 10 9 11 2
28 10 0 9 1 10 9 13 10 0 9 2 7 3 10 9 3 0 13 15 7 15 13 1 9 1 10 9 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
32 1 11 13 3 10 9 1 11 3 0 2 7 13 9 2 9 7 9 2 13 1 10 9 1 10 9 11 11 1 11 11 2
11 1 10 9 12 13 10 9 1 12 9 2
34 10 9 15 13 13 1 10 3 9 11 11 11 1 12 1 9 1 10 9 1 9 1 11 2 10 9 15 13 10 0 9 1 12 2
49 10 9 0 1 10 9 13 10 9 1 10 9 1 9 7 9 1 9 2 16 13 13 16 10 0 9 2 1 9 10 0 9 2 13 0 7 3 7 10 3 0 7 7 3 13 2 9 2 2
33 4 1 13 2 3 13 1 10 11 1 11 11 2 1 11 1 12 1 10 9 1 11 11 11 2 13 1 10 9 1 0 9 2
16 1 12 4 1 13 10 9 1 9 11 2 16 13 1 12 2
51 10 9 0 1 10 9 1 10 0 9 13 1 8 2 8 1 9 1 11 1 11 7 12 1 9 1 11 1 11 2 2 1 15 15 13 1 9 1 9 2 10 9 16 15 13 0 1 10 9 0 2
35 1 10 9 2 10 9 1 11 2 1 3 3 1 9 1 10 9 1 10 11 11 2 4 1 13 1 10 9 1 11 1 11 2 11 2
30 13 11 10 11 7 10 9 2 1 10 9 0 15 13 11 2 10 0 11 11 2 13 1 9 0 2 9 7 9 2
34 1 12 15 13 10 0 9 1 10 9 2 3 1 10 9 1 2 11 2 11 7 11 2 7 1 10 9 9 1 12 8 12 5 2
19 10 11 13 1 10 10 9 1 10 11 2 12 9 1 10 9 1 11 2
73 10 9 1 11 1 11 2 11 2 7 11 1 10 9 0 2 13 10 9 0 0 2 16 13 10 9 0 1 10 9 1 9 0 1 9 7 9 0 2 0 13 1 12 1 9 1 10 11 1 10 9 7 9 0 1 10 9 1 9 0 2 4 10 0 9 13 10 9 1 11 1 12 2
7 1 15 15 3 13 9 2
37 1 12 13 1 10 9 9 2 9 1 11 11 1 11 7 3 3 13 10 0 9 1 2 8 8 1 10 9 2 1 10 11 11 11 11 11 2
34 13 3 0 1 1 10 10 9 15 0 10 12 1 11 1 10 15 1 12 9 13 10 9 1 10 9 1 10 9 0 1 10 9 2
27 10 9 4 13 15 1 15 1 10 9 2 1 9 0 1 10 0 9 2 10 0 9 7 10 9 0 2
32 10 9 1 15 13 16 10 9 13 3 9 1 10 9 1 13 1 10 11 11 16 13 10 9 1 10 9 13 1 10 9 2
15 1 15 13 0 2 3 7 15 4 13 13 1 0 9 2
38 2 15 13 1 11 2 13 10 9 1 10 9 0 2 3 0 2 13 9 1 10 9 2 4 7 13 15 3 0 1 16 13 10 9 2 2 13 2
23 10 9 13 1 10 9 4 4 13 1 10 9 0 1 12 2 12 2 12 7 12 9 2
8 11 13 10 9 1 9 9 2
40 3 10 9 4 13 1 10 9 0 13 15 1 3 0 7 3 3 15 4 13 1 10 8 2 8 1 9 13 1 10 9 2 7 1 9 0 1 10 9 2
31 10 0 9 1 9 13 10 12 1 11 1 12 2 1 11 2 1 10 9 11 1 11 2 10 9 0 1 10 9 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
43 12 9 1 9 1 10 9 0 1 10 9 12 11 11 7 11 11 15 13 3 1 13 10 9 1 12 9 2 16 13 15 1 10 9 9 1 10 9 0 0 1 11 2
59 1 10 12 9 2 11 13 13 1 10 12 5 0 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
30 10 9 13 3 1 12 9 7 1 15 13 10 9 2 9 7 9 2 9 1 9 2 9 2 9 7 9 1 11 2
26 1 9 0 2 13 0 16 13 10 9 1 11 12 2 9 1 10 9 12 2 7 9 1 11 12 2
21 10 9 13 1 9 1 9 0 2 7 13 13 1 10 9 0 0 2 11 2 2
14 10 9 0 4 13 10 0 9 2 10 12 1 11 2
35 7 1 10 9 1 10 9 1 9 0 2 15 4 13 10 9 0 1 9 0 3 1 10 9 2 1 15 1 10 0 9 1 10 9 2
42 1 10 11 1 11 2 12 2 7 10 9 1 10 9 16 13 10 9 10 9 11 13 13 1 11 1 12 7 10 9 13 1 10 9 11 1 11 7 1 10 9 2
37 10 9 1 10 9 2 1 10 9 0 2 3 13 10 9 0 13 1 10 9 1 9 1 10 9 0 1 9 7 9 1 10 9 1 10 9 2
24 1 10 9 0 13 10 9 0 2 3 16 3 13 10 9 13 3 1 10 9 1 10 9 2
28 1 9 1 11 1 12 10 11 11 11 15 13 1 9 1 10 9 11 1 11 1 10 9 7 3 15 13 2
38 3 13 10 10 9 3 0 1 10 11 11 2 1 10 9 11 2 11 7 10 11 11 2 1 10 9 1 10 9 16 13 1 10 9 10 10 9 2
11 10 9 1 10 9 13 0 1 15 9 2
17 10 12 13 10 0 9 1 13 10 9 0 15 3 1 10 15 2
7 15 15 13 1 10 9 2
35 1 9 13 1 9 2 7 15 13 3 1 10 9 1 9 1 10 9 7 15 13 1 10 9 1 10 0 9 2 9 13 1 11 11 2
22 1 10 9 1 9 0 2 11 11 2 10 9 1 10 9 1 10 8 13 9 0 2
18 1 12 15 13 10 9 2 1 0 9 1 9 2 1 10 12 9 2
34 10 9 13 1 10 13 10 9 1 10 9 2 13 1 10 9 11 0 2 1 10 9 11 1 10 9 0 2 13 10 9 1 11 2
94 1 10 9 1 10 11 1 11 1 11 1 11 11 1 11 2 7 13 9 11 11 1 11 2 11 11 1 10 9 1 12 2 15 4 13 10 0 9 0 1 9 1 0 9 1 11 2 3 1 11 2 11 7 11 2 1 9 1 10 9 13 1 9 0 9 3 1 10 3 9 1 10 9 2 11 11 11 1 15 2 7 1 10 9 1 10 9 0 1 10 9 1 15 2
20 10 9 1 11 13 10 0 9 1 11 2 1 3 1 10 9 0 0 11 2
18 11 1 11 13 10 12 1 11 1 12 1 11 1 11 2 11 2 2
22 11 1 10 11 13 10 9 0 2 0 1 10 9 1 11 2 9 0 1 11 2 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
19 15 1 10 9 1 11 11 13 11 2 11 11 2 11 11 2 11 11 2
66 10 9 0 0 15 13 1 10 9 0 1 3 3 15 13 1 10 9 7 10 9 2 13 0 9 1 10 9 7 1 3 9 16 15 13 1 9 1 9 1 10 9 2 13 1 0 9 1 10 9 2 0 9 1 9 2 3 0 9 1 10 9 7 10 9 2
23 11 13 10 9 2 1 9 2 2 9 2 2 1 10 9 1 11 2 11 2 1 11 2
4 13 10 12 2
61 11 13 1 9 0 1 4 13 10 9 1 10 4 1 13 10 9 1 10 9 10 15 4 1 4 13 1 10 9 2 15 4 13 1 10 11 11 11 7 3 4 13 1 10 9 3 16 13 10 9 0 2 3 10 9 4 13 1 10 9 2
27 3 13 1 16 10 11 4 13 1 10 9 7 10 9 15 13 1 9 0 2 1 13 9 1 10 9 2
45 1 9 12 1 11 1 10 12 2 4 13 1 10 12 5 2 1 12 9 1 9 1 9 2 3 12 9 1 9 2 1 12 9 1 9 1 9 2 3 12 9 1 9 2 2
21 3 15 4 13 1 9 1 13 10 9 1 11 2 3 13 1 9 0 9 0 2
23 10 0 11 4 13 10 9 1 10 9 1 10 9 1 9 13 1 10 12 1 10 9 2
24 10 0 9 1 10 9 2 2 11 2 2 4 13 10 9 12 1 11 1 12 1 9 0 2
11 10 9 4 13 1 10 9 1 10 9 2
15 10 12 1 11 1 12 13 13 10 9 1 10 9 0 2
28 10 9 1 11 15 13 1 9 0 1 10 11 11 1 11 1 10 9 1 10 9 0 2 1 12 7 12 2
42 16 13 2 13 13 15 1 11 11 2 3 3 16 13 15 3 1 10 9 13 11 11 2 7 16 11 13 3 0 2 1 9 1 10 9 1 11 1 13 15 2 2
49 10 2 11 2 0 2 13 10 9 13 1 11 11 1 10 9 1 10 15 10 9 0 1 10 9 13 16 10 9 13 10 9 13 3 7 3 13 1 10 0 9 1 10 9 1 15 4 13 2
12 10 10 9 15 13 3 1 11 7 10 9 2
17 3 13 0 9 1 9 1 10 9 1 9 7 10 9 3 0 2
69 1 10 9 2 9 1 11 13 10 9 0 1 10 11 2 15 13 10 10 9 1 11 3 13 2 1 11 12 2 16 13 10 9 1 11 11 12 1 2 11 2 7 9 2 2 11 2 9 1 11 1 12 7 12 2 7 11 12 1 11 12 10 11 7 11 12 10 11 2
25 2 11 2 2 13 10 9 0 7 0 16 4 13 1 9 1 10 16 10 9 13 10 0 9 2
23 11 11 11 2 13 1 11 2 11 2 13 10 9 2 9 2 9 1 9 7 9 0 2
12 15 13 1 10 9 0 2 0 7 0 0 2
20 10 9 13 1 10 9 1 1 10 0 9 1 9 2 3 0 1 12 2 2
19 15 4 13 1 10 9 0 1 13 15 1 13 10 9 0 1 10 9 2
23 0 1 9 0 2 1 15 2 7 9 1 9 2 13 10 9 13 1 10 3 9 2 2
40 10 11 13 3 1 10 0 9 2 15 1 13 10 9 1 10 9 0 7 15 1 13 1 10 9 0 10 9 15 4 4 13 1 10 9 0 1 10 9 2
15 13 9 0 1 11 11 1 10 11 11 1 11 1 12 2
24 1 13 10 9 4 1 13 10 12 5 9 1 10 9 2 12 2 7 13 1 9 1 12 2
26 1 12 4 1 13 10 9 2 11 11 2 1 10 9 1 2 11 2 11 2 11 2 11 7 11 2
21 10 9 1 9 13 1 10 9 1 10 9 1 10 9 0 13 0 10 9 0 2
11 11 11 13 15 1 10 9 1 10 11 2
13 1 9 13 10 9 1 9 0 7 3 9 15 2
15 10 9 11 13 16 11 13 12 9 1 3 12 1 11 2
40 1 10 9 1 9 2 11 13 16 11 13 10 12 5 1 10 9 1 9 1 8 5 8 10 2 9 1 9 2 16 15 13 13 12 9 1 9 1 9 2
58 1 10 9 15 13 9 1 10 0 9 0 1 10 9 1 9 1 10 9 3 15 13 16 10 9 1 11 4 1 13 1 10 0 9 2 9 16 13 3 0 1 10 9 13 1 10 9 1 10 9 2 11 11 1 11 1 12 2
13 10 9 1 9 13 1 12 9 2 2 5 5 2
22 11 11 13 10 0 9 1 10 9 3 1 13 1 10 0 9 12 9 1 10 11 2
16 1 10 9 1 10 9 2 10 9 1 11 1 11 15 13 2
40 1 10 9 1 11 13 0 13 3 0 9 1 9 10 1 10 9 0 7 0 1 10 11 7 10 9 0 2 3 1 9 1 9 1 10 9 7 10 9 2
7 13 1 9 1 9 0 2
3 11 11 2
16 10 9 13 3 3 7 15 13 10 9 2 13 1 10 9 2
7 10 0 9 13 11 11 2
30 1 10 0 9 1 10 11 11 11 11 2 11 13 1 9 1 10 0 9 1 10 11 1 11 10 9 1 10 9 2
19 13 10 9 1 9 0 2 10 9 0 1 9 2 9 0 2 0 9 2
34 13 1 9 1 10 9 0 1 10 9 1 10 9 1 11 12 1 12 7 4 13 1 9 0 3 11 12 13 1 10 9 1 12 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
39 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 13 10 0 9 1 9 7 9 2 13 3 1 10 9 13 1 10 9 1 8 8 8 11 2
39 1 9 2 1 10 0 16 13 10 9 11 12 7 10 9 11 11 2 4 1 13 1 10 9 1 11 16 13 10 9 1 9 1 10 9 1 10 9 2
33 3 2 10 9 13 0 1 13 1 9 7 9 2 7 3 3 1 13 7 13 0 9 2 3 7 3 0 7 13 13 10 9 2
30 1 10 9 1 12 9 15 4 13 10 9 1 10 11 7 13 9 10 9 1 9 7 9 1 15 15 3 13 11 2
37 10 9 13 1 10 9 1 10 9 2 3 15 13 10 9 1 10 15 15 13 10 11 1 10 11 7 10 10 9 1 10 9 11 1 10 9 2
22 15 13 3 1 10 9 2 11 2 7 4 13 1 11 2 12 1 11 1 12 2 2
19 1 10 0 9 3 15 13 1 10 11 1 11 2 13 10 9 1 12 2
40 1 10 9 1 9 0 2 16 10 9 13 1 9 2 15 13 11 2 7 1 10 9 11 2 1 15 16 13 10 9 0 7 11 2 1 16 13 10 9 2
13 10 9 1 10 9 1 0 15 13 3 1 3 2
28 11 13 10 9 0 3 0 1 11 1 9 16 13 1 9 10 9 1 10 9 1 9 1 10 9 0 0 2
17 10 9 13 1 10 9 1 13 10 0 9 0 1 10 9 0 2
23 10 9 3 0 13 13 10 1 11 2 1 10 15 3 15 13 16 13 10 9 3 0 2
19 11 11 13 10 9 1 9 0 9 1 10 9 1 10 9 2 11 2 2
37 3 13 10 9 0 1 9 0 1 10 9 1 9 13 1 9 7 12 9 1 0 9 2 13 1 0 9 0 1 9 0 16 13 10 9 0 2
13 3 13 1 10 9 12 1 10 9 0 10 11 2
40 10 9 1 9 1 11 1 10 11 2 1 15 13 16 15 13 1 10 9 1 11 8 13 3 9 1 10 9 7 10 9 1 11 2 12 9 0 1 3 2
36 10 9 0 2 9 0 1 9 2 10 11 11 2 13 10 9 1 9 9 1 11 11 11 13 3 1 10 9 1 11 1 12 1 11 11 2
21 15 13 1 7 13 16 13 12 9 7 16 13 10 9 4 7 13 3 1 12 2
65 13 0 9 7 9 1 11 2 1 10 15 13 12 9 2 10 11 11 1 10 11 2 10 11 11 1 11 11 2 11 11 7 10 11 11 2 2 3 1 10 11 2 11 1 11 2 11 1 11 2 7 2 11 7 11 2 2 15 1 11 1 10 9 2 2
5 2 9 7 9 2
20 4 13 1 12 2 13 1 12 2 7 13 1 10 11 11 11 11 1 11 2
13 1 9 10 0 9 1 11 13 1 10 0 9 2
15 13 1 11 13 1 10 11 2 12 1 10 11 7 11 2
7 3 13 1 10 10 11 2
26 11 11 13 10 9 1 11 0 13 7 13 15 2 2 11 2 2 3 13 16 10 9 15 4 13 2
23 10 9 3 4 13 2 15 16 13 10 9 1 0 9 7 9 0 0 1 10 9 0 2
40 13 0 1 10 9 11 11 1 10 12 1 11 1 12 2 1 10 15 13 10 9 2 11 2 13 1 11 1 12 7 10 9 11 2 13 1 11 1 12 2
6 11 11 2 12 2 2
5 2 3 4 13 2
27 7 16 10 11 11 1 10 9 3 13 9 1 9 0 3 15 1 10 9 13 1 10 11 1 10 11 2
22 3 0 11 4 13 7 13 3 1 10 9 13 16 10 9 0 13 10 9 1 9 2
20 11 11 2 9 2 8 8 2 13 1 12 2 13 10 9 7 9 0 0 2
9 2 13 10 9 3 0 7 0 2
98 10 9 1 11 13 1 9 0 9 1 10 9 2 13 11 7 11 11 2 3 7 10 9 1 11 13 16 13 2 0 1 9 2 2 16 15 3 13 0 1 16 10 9 13 16 10 0 1 9 1 10 11 4 13 16 11 13 1 9 0 7 16 2 1 10 9 1 12 9 2 4 13 1 10 0 9 1 10 9 1 10 12 1 11 1 12 2 1 10 9 3 13 1 10 9 1 9 2
42 11 11 2 10 9 4 13 1 11 2 3 11 2 11 2 11 2 7 13 1 9 1 10 9 11 11 1 4 13 1 10 9 1 11 11 7 11 11 1 11 11 2
23 15 13 10 9 2 10 9 1 10 9 2 10 9 2 3 7 10 9 16 15 13 0 2
37 4 13 1 0 9 0 13 1 10 9 0 1 11 3 12 9 3 1 10 9 1 11 11 7 13 10 12 1 11 1 12 1 10 9 11 11 2
19 11 13 10 9 0 1 9 0 16 13 1 10 11 1 11 1 10 11 2
5 3 4 13 15 2
16 10 9 0 15 13 1 11 3 12 9 7 3 13 10 12 2
16 13 10 9 0 16 4 1 13 15 1 9 1 9 1 9 2
68 10 9 15 13 1 10 9 1 10 16 13 10 0 9 1 10 9 1 10 9 2 10 9 13 1 10 0 9 0 13 1 10 9 1 9 1 9 9 7 10 9 1 10 9 1 9 0 7 1 10 9 2 7 1 10 9 0 13 1 10 9 1 10 9 16 13 0 2
45 2 11 2 2 2 11 11 2 7 2 11 2 2 1 10 9 2 13 9 1 9 2 7 16 2 11 2 15 13 1 0 9 1 10 9 2 1 10 15 13 10 9 1 11 2
14 1 13 15 13 10 9 16 13 10 9 1 10 9 2
35 11 2 10 0 9 0 1 11 2 13 10 3 13 1 10 0 9 2 1 15 3 12 9 4 13 2 10 9 13 10 12 7 12 9 2
49 1 3 1 11 11 2 13 10 2 8 8 8 2 2 10 9 3 1 10 9 0 3 10 9 4 13 10 9 1 9 7 13 10 9 2 13 15 15 7 13 1 10 9 3 13 1 10 9 2
34 10 9 0 1 9 1 10 9 1 11 1 11 1 12 15 13 1 16 2 1 15 9 1 10 9 2 15 15 4 1 4 13 3 2
21 7 1 12 13 9 1 10 9 0 1 9 2 12 9 4 13 1 12 5 2 2
37 2 1 10 9 2 11 11 13 3 1 10 9 0 13 1 13 10 9 1 11 2 2 13 10 11 10 9 1 10 9 0 1 10 9 11 11 2
10 1 12 2 10 9 13 1 12 9 2
33 1 10 9 1 10 11 0 13 10 9 11 2 0 9 11 13 11 7 10 11 2 9 1 10 0 9 13 11 2 11 7 11 2
28 11 3 3 13 10 9 1 10 9 3 7 13 1 9 1 11 11 1 13 15 1 11 11 1 12 9 0 2
23 3 1 13 2 11 13 16 11 1 11 13 1 9 2 0 7 13 0 9 1 10 9 2
72 10 9 2 16 15 13 1 9 1 10 11 12 1 10 11 12 1 11 7 13 10 9 0 1 10 9 1 11 2 13 12 9 1 9 1 9 7 9 1 9 1 10 8 1 10 9 2 1 10 15 11 13 15 1 10 9 0 2 1 9 0 1 12 9 2 16 13 1 10 9 0 2
52 1 9 1 13 3 10 9 13 1 10 9 2 16 13 1 10 9 0 0 2 13 13 9 2 9 2 9 2 8 2 10 9 1 10 9 1 11 15 13 1 9 2 9 2 9 2 9 2 9 7 9 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 9 2
17 10 9 15 13 1 10 12 9 3 2 7 3 1 10 0 9 2
32 7 10 9 2 11 2 10 9 16 13 1 4 13 1 10 0 9 7 9 7 11 2 13 10 9 2 7 4 1 13 15 2
11 10 12 1 11 1 12 4 13 1 9 2
11 11 13 10 9 1 9 1 10 9 11 2
24 11 1 10 11 15 13 1 9 0 1 10 11 11 2 16 3 13 16 10 9 13 10 9 2
34 1 10 12 7 10 12 1 11 2 13 9 15 13 1 11 1 10 11 2 1 10 9 11 1 11 2 10 9 0 1 9 7 9 2
16 11 11 11 2 7 10 9 13 10 9 11 11 1 10 11 2
7 13 9 0 7 9 0 2
21 9 11 2 16 3 13 10 0 9 2 3 4 13 10 0 9 7 10 10 9 2
40 11 13 10 9 7 9 0 2 1 10 9 1 9 2 9 2 9 1 11 2 1 10 9 1 11 2 15 2 11 7 9 1 11 2 15 2 11 2 11 2
14 10 9 1 10 9 13 13 10 10 9 1 10 9 2
13 1 12 13 1 10 11 11 11 2 3 13 9 2
9 10 9 13 10 9 1 10 9 2
25 0 9 2 10 9 13 1 10 9 0 1 9 1 10 9 2 3 13 15 0 1 10 9 13 2
12 10 9 1 9 1 10 9 13 1 5 12 2
53 1 10 9 15 13 10 9 2 11 2 2 1 10 9 11 11 2 13 1 10 9 12 2 16 15 13 1 10 9 1 10 9 1 10 11 11 1 11 2 7 3 15 13 1 10 9 1 11 11 1 10 11 2
18 11 13 1 10 9 1 10 11 1 10 11 7 15 13 1 10 9 2
37 10 9 0 1 9 1 10 9 1 10 9 0 13 10 9 10 9 1 12 9 2 10 12 5 1 9 1 9 1 10 0 9 1 10 0 9 2
10 13 0 1 11 1 10 9 1 11 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
6 3 15 13 10 9 2
22 10 0 9 1 10 9 13 1 10 9 12 2 1 10 9 1 10 9 11 1 11 2
21 13 10 0 9 1 11 11 11 2 7 13 1 13 10 11 11 1 10 10 9 2
28 10 9 1 11 2 1 10 9 1 2 11 13 16 15 13 10 9 9 0 0 2 13 15 3 10 9 0 2
49 10 9 1 10 9 13 0 2 10 9 1 9 0 2 10 9 0 2 10 9 0 2 10 9 0 3 15 13 10 9 2 9 7 9 2 3 1 13 9 7 9 1 3 13 1 9 1 9 2
43 1 10 9 1 10 0 9 2 15 13 1 10 9 11 10 9 1 10 9 0 3 0 2 1 10 15 15 13 1 9 1 11 13 1 10 9 1 10 9 1 10 9 2
22 10 0 11 13 1 9 10 9 1 11 2 13 16 13 10 9 16 13 1 10 9 2
34 11 2 11 1 11 2 13 10 9 7 9 0 2 13 1 10 9 1 11 11 1 10 9 1 11 7 1 10 9 0 9 1 11 2
31 16 4 13 1 10 9 1 13 10 11 1 10 16 13 11 2 3 13 2 3 1 10 9 1 11 11 2 9 0 3 2
22 3 2 11 15 13 1 11 2 10 9 1 11 2 7 11 13 1 10 9 1 9 2
22 13 12 9 2 0 9 10 9 2 16 13 10 0 9 1 10 9 1 10 9 0 2
13 10 9 13 0 7 0 2 15 13 13 1 9 2
16 10 12 0 9 1 9 4 13 1 12 9 0 1 10 9 2
54 10 12 1 11 2 10 9 15 13 2 10 9 1 11 13 3 1 10 9 1 11 2 15 4 13 1 9 10 12 1 11 7 3 15 13 10 9 1 10 9 1 10 9 16 3 4 13 1 10 9 0 1 11 2
12 11 13 10 9 0 2 13 1 11 2 11 2
60 1 10 15 15 15 13 0 13 1 10 9 1 10 9 0 2 16 3 13 10 9 1 10 9 13 2 7 10 2 9 2 1 15 1 2 9 1 10 11 2 2 1 9 1 10 2 9 1 10 9 0 2 15 13 2 3 3 2 0 2
15 2 7 3 4 1 13 1 15 2 16 15 13 1 15 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
31 11 13 10 9 1 9 1 10 11 1 11 7 15 13 1 11 11 11 2 10 9 1 11 16 13 1 10 9 1 11 2
37 10 9 4 13 15 1 10 9 0 1 13 1 10 9 1 10 9 0 1 10 9 2 3 1 16 13 10 9 0 1 10 9 3 1 13 15 2
26 13 10 9 0 2 10 9 1 10 9 12 7 10 0 9 0 1 10 11 7 10 11 1 9 0 2
32 10 9 1 10 11 13 0 8 10 9 1 10 9 1 9 0 16 10 9 4 13 2 3 3 15 13 1 10 9 1 9 2
26 7 15 16 10 9 13 10 9 16 13 10 9 1 10 9 13 10 9 1 10 9 0 7 10 9 2
7 13 10 9 1 12 9 2
16 1 15 9 2 10 9 4 13 1 16 10 9 13 9 0 2
34 1 10 9 1 9 7 9 13 1 11 2 10 9 13 10 9 1 9 0 9 1 9 2 9 1 10 9 2 9 2 9 7 9 2
25 10 9 4 13 15 1 10 9 1 10 9 2 8 2 8 8 8 8 2 5 2 8 2 8 2
21 13 10 9 1 10 11 1 10 11 7 13 10 0 9 1 10 9 1 10 9 2
17 13 1 11 11 2 10 9 0 4 13 10 12 1 11 1 12 2
10 1 15 15 13 9 1 9 7 9 2
42 10 9 1 11 1 10 1 15 13 1 10 9 7 3 11 4 4 13 16 3 15 13 1 13 16 4 4 13 11 11 11 1 10 9 1 9 3 4 13 10 9 2
28 11 11 11 1 10 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 2 9 2 9 7 9 0 2
48 10 9 13 3 1 10 9 1 9 1 9 2 10 11 2 1 10 9 11 2 7 12 9 0 2 11 1 10 9 11 2 11 11 1 11 1 10 9 11 2 7 11 1 10 9 11 2 2
20 11 11 13 1 9 1 10 2 9 2 7 1 10 12 9 13 11 11 11 2
29 1 10 9 13 13 15 1 10 9 0 7 1 12 13 10 9 2 3 16 10 12 1 11 1 12 13 10 9 2
33 13 10 9 1 10 9 7 10 9 1 10 9 4 1 13 7 10 9 15 13 1 10 10 9 1 16 13 1 10 9 1 11 2
5 15 13 1 11 2
10 10 9 4 13 1 3 1 12 9 2
34 10 11 1 11 1 10 11 7 3 1 10 11 1 11 2 1 9 2 11 11 11 11 11 2 13 10 9 9 1 10 9 1 11 2
37 9 11 11 7 11 2 11 1 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 13 10 9 7 9 1 10 11 11 13 1 11 2
27 10 9 13 0 2 0 7 15 13 3 1 10 9 1 10 9 11 11 2 11 11 7 10 9 1 9 2
11 9 2 9 1 9 0 1 10 9 1 11
17 1 12 2 10 9 13 10 9 1 2 11 11 11 11 11 2 2
32 1 12 2 1 10 9 1 11 1 10 9 0 7 10 9 1 11 2 11 11 13 1 11 2 13 1 10 9 1 10 11 2
41 10 11 2 11 2 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 1 11 11 2 1 10 9 1 11 7 9 1 11 2 11 2 11 2 11 2
24 12 9 3 3 2 11 13 1 11 2 3 13 10 9 1 10 9 1 11 2 3 1 11 2
51 10 9 1 11 13 0 9 1 10 9 12 2 10 15 4 13 2 1 15 2 1 10 9 0 1 10 9 1 10 9 12 2 7 10 9 1 0 9 0 2 3 13 1 10 9 0 7 1 10 9 2
29 1 9 2 13 10 9 12 2 10 9 0 13 1 11 2 9 3 10 9 0 13 10 9 7 10 9 1 9 2
18 10 9 13 16 3 4 13 3 1 12 7 12 9 1 13 1 9 2
46 13 7 13 1 10 9 0 11 11 11 2 9 1 11 2 7 1 10 9 1 10 9 0 1 11 2 15 1 10 9 1 11 2 13 10 9 1 11 1 10 9 1 13 10 9 2
47 11 13 9 1 9 11 2 11 2 8 2 11 2 1 9 1 11 7 1 10 0 11 2 7 11 2 11 2 8 2 11 2 2 1 10 9 1 11 7 10 11 1 10 9 1 9 2
31 13 0 3 10 9 13 0 1 13 9 0 1 11 1 0 7 0 2 10 9 16 13 3 0 1 10 9 0 1 11 2
27 10 9 2 9 1 10 9 0 7 9 0 13 1 10 0 11 1 12 9 1 10 9 1 10 9 0 2
14 15 13 11 11 2 9 2 11 2 1 11 1 12 2
31 3 2 10 9 4 13 1 10 9 2 9 7 9 1 10 9 7 9 1 9 0 7 0 2 0 1 13 15 3 2 2
18 10 9 0 2 13 1 11 11 2 4 13 1 10 11 11 1 11 2
41 1 10 9 0 1 11 11 11 15 13 10 9 1 11 11 1 11 11 11 2 7 1 10 9 0 4 13 10 9 0 1 10 9 1 11 11 2 11 10 11 2
39 1 9 0 11 13 10 9 13 1 11 7 11 2 9 2 7 3 13 10 9 2 13 3 10 9 1 9 0 1 10 2 9 1 11 2 1 10 9 2
11 10 9 1 10 9 4 13 1 10 9 8
43 13 15 1 10 9 0 16 13 1 10 9 1 10 16 13 0 11 7 3 13 1 3 13 1 10 9 16 13 10 9 0 16 13 3 15 13 10 0 9 1 10 9 2
22 10 9 13 16 10 9 1 10 9 2 4 7 13 15 1 10 9 16 13 10 9 2
24 1 10 0 9 1 10 11 2 13 1 0 9 13 3 12 9 7 3 13 7 12 3 9 2
24 13 1 10 9 1 10 11 11 2 2 11 7 10 11 1 10 11 11 2 2 11 12 2 2
43 10 9 13 15 1 10 3 0 9 1 10 0 9 1 12 9 2 10 9 1 9 1 11 7 10 9 1 10 9 2 11 2 2 1 10 9 1 3 12 12 9 13 2
15 1 0 9 13 1 9 10 9 0 1 9 1 10 9 2
15 11 11 13 10 9 1 9 1 9 0 1 10 9 11 2
60 11 4 13 1 12 1 10 9 1 7 13 1 10 9 3 0 2 3 13 2 1 1 10 9 13 1 10 9 1 10 15 2 4 13 1 9 1 14 15 16 13 2 7 3 4 13 10 9 1 10 9 2 16 13 1 11 11 1 12 2
26 3 13 2 16 2 10 9 1 9 16 13 1 0 1 15 2 7 7 10 9 15 13 1 9 0 2
15 2 10 9 1 10 12 9 7 10 0 9 1 10 9 2
20 10 9 13 13 10 10 9 0 1 10 9 7 10 9 13 1 10 10 9 2
22 3 4 13 16 8 8 13 10 11 11 1 11 2 12 13 1 10 9 1 10 9 2
35 3 10 9 13 1 9 1 10 0 9 1 10 9 0 7 15 13 1 12 9 3 0 16 13 10 9 3 2 11 11 7 11 11 11 2
22 15 13 16 4 13 10 9 0 1 10 9 2 7 10 9 13 13 15 10 9 0 2
4 13 1 11 2
21 3 10 9 7 10 9 15 4 13 7 13 15 1 10 0 9 1 10 9 0 2
5 1 12 13 12 2
21 13 13 15 10 9 1 10 0 9 16 15 4 13 10 0 9 1 9 1 11 2
69 13 10 9 0 1 10 11 11 3 1 10 9 1 11 2 11 1 10 11 2 10 11 2 11 2 11 2 11 7 11 1 10 11 1 10 9 1 11 2 7 11 1 10 11 2 11 2 11 2 11 2 11 1 11 2 11 1 10 11 2 11 7 11 1 10 9 1 11 2
4 2 13 0 2
56 10 9 1 10 9 7 10 9 1 10 11 11 1 11 11 11 15 13 1 10 9 1 10 9 7 10 9 1 10 9 1 9 1 9 1 10 9 1 10 9 1 10 9 7 10 9 1 10 9 7 10 9 1 10 9 2
20 7 15 1 15 15 13 1 10 9 0 7 1 10 9 13 3 1 10 9 2
10 15 13 10 9 1 13 15 15 3 2
35 1 9 7 9 2 10 9 13 10 9 0 13 1 10 9 16 1 9 1 10 9 1 11 13 1 9 0 10 0 9 1 9 3 0 2
40 3 13 1 10 9 1 10 9 0 1 9 7 9 0 2 7 13 16 1 3 1 12 9 4 4 13 10 9 2 3 1 9 0 1 10 12 9 1 9 2
43 16 4 13 3 10 11 11 10 9 1 11 3 13 1 9 16 4 13 15 10 9 1 10 9 1 15 3 2 15 13 1 10 9 2 9 7 1 15 3 16 15 13 2
14 10 9 13 10 9 1 9 2 9 0 7 9 0 2
23 10 12 9 13 10 9 1 9 2 13 10 9 1 9 2 1 10 9 1 10 0 9 2
36 10 9 0 4 4 1 13 1 10 9 1 15 2 13 1 15 16 4 13 15 10 9 7 13 1 10 9 0 1 10 9 1 10 9 2 2
14 13 10 9 1 9 0 7 1 9 0 1 9 0 2
33 11 0 11 2 11 2 11 2 12 1 11 1 12 8 11 2 12 1 11 1 12 2 2 9 0 0 7 9 1 10 9 0 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
28 10 9 4 13 1 11 7 11 2 10 9 13 10 9 1 9 1 10 9 2 11 2 11 7 11 11 2 2
12 3 15 13 16 13 15 1 10 2 9 2 2
38 10 9 13 1 0 9 2 3 0 1 10 0 9 2 7 13 9 1 10 9 2 9 2 9 0 2 9 1 10 9 0 2 7 9 1 9 0 2
33 10 9 13 10 9 1 10 9 1 10 11 2 10 9 1 10 9 3 10 9 13 0 2 1 10 9 3 0 1 10 9 0 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
48 10 3 0 9 1 9 0 1 10 9 1 11 2 13 1 12 1 10 9 1 11 2 10 0 9 13 1 9 1 10 9 1 10 11 1 11 2 1 15 15 10 9 13 2 11 11 2 2
9 11 13 10 0 9 1 10 9 2
20 3 1 10 9 1 10 9 1 11 7 11 2 7 1 11 1 10 0 9 2
12 13 9 1 9 1 10 9 1 9 3 0 2
23 10 9 13 0 1 10 9 1 10 9 0 1 11 2 13 9 1 10 0 9 1 11 2
12 13 10 9 1 12 2 8 11 1 12 2 2
13 3 13 10 9 0 7 13 10 9 1 10 9 2
15 1 10 12 1 11 1 12 13 1 10 11 11 11 11 2
23 10 9 13 10 9 7 3 3 9 10 9 1 10 9 13 10 9 0 1 10 11 0 2
15 13 10 9 1 0 9 2 16 13 10 9 0 1 9 2
37 10 11 4 13 3 10 12 1 11 1 12 2 13 3 1 10 9 13 9 1 10 11 7 11 11 2 3 7 13 15 1 10 2 11 11 2 2
15 10 11 1 10 11 13 10 9 0 13 1 11 2 11 2
27 10 0 9 13 10 11 11 7 10 9 0 7 0 2 3 7 10 9 13 1 10 9 1 10 9 0 2
39 3 1 10 9 0 2 1 10 0 9 1 9 2 2 10 9 16 13 10 9 0 1 10 9 13 1 10 9 1 10 10 9 7 3 2 13 15 3 2
29 3 11 13 16 11 11 13 10 9 1 11 2 15 4 13 3 3 1 16 10 9 16 15 4 1 13 4 13 2
42 13 1 10 9 2 10 11 11 3 3 13 1 10 9 1 10 11 11 1 11 2 3 1 10 9 0 1 11 2 2 7 4 7 4 13 1 10 9 1 10 9 2
23 15 13 1 10 12 7 10 12 1 11 1 12 1 10 11 11 1 10 11 1 11 11 2
22 1 10 9 0 2 10 9 13 0 1 15 1 10 10 9 0 2 13 1 12 9 2
45 11 15 4 13 1 10 9 1 9 0 1 7 15 15 13 1 10 9 0 2 7 15 4 13 1 10 0 9 2 1 10 15 4 13 15 3 9 1 10 9 7 1 10 9 2
49 1 10 9 1 9 1 10 9 2 11 4 13 10 9 1 10 9 1 10 9 0 0 2 1 10 0 9 16 2 13 1 15 2 15 13 0 7 0 2 13 1 10 0 9 1 10 9 0 2
24 15 13 13 1 10 9 3 0 2 1 10 9 1 10 11 11 2 11 11 2 1 11 11 2
20 1 0 9 13 1 10 9 15 4 13 1 9 1 9 1 9 7 9 0 2
58 13 10 9 0 1 10 9 16 13 13 9 1 9 0 1 9 1 9 0 7 9 1 10 0 9 10 9 0 16 13 10 9 13 10 9 0 1 10 9 1 10 9 7 9 0 1 10 9 1 10 9 1 10 9 1 9 0 2
52 1 10 9 2 12 10 9 0 1 11 11 11 3 4 13 1 10 9 2 4 13 1 10 9 0 2 11 0 2 1 10 12 2 1 10 9 1 11 11 7 1 10 9 1 9 1 10 9 1 11 11 2
17 10 0 9 3 0 13 10 9 2 1 9 15 13 10 0 9 2
10 4 13 10 12 1 11 1 10 12 2
32 13 10 9 0 2 13 9 1 9 1 11 7 1 11 3 13 1 10 9 1 10 9 7 13 0 9 1 9 1 11 12 2
10 10 9 13 16 13 1 9 1 12 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
20 10 9 11 3 15 13 1 10 9 1 10 9 11 2 15 4 13 1 12 2
20 13 9 0 1 10 9 1 9 1 10 11 11 2 11 2 2 11 2 11 2
60 10 9 13 9 0 1 9 12 1 10 11 2 13 13 2 9 1 10 9 1 9 1 10 9 1 10 9 7 9 1 9 2 7 1 10 9 1 10 9 1 12 9 2 13 1 9 2 9 2 9 0 7 0 2 9 0 7 9 0 2
23 11 11 11 13 10 9 0 0 1 10 9 11 2 9 1 10 11 11 1 10 9 12 2
33 1 12 2 10 9 0 13 10 9 1 10 9 0 2 1 0 9 2 9 1 9 0 7 8 2 9 2 10 0 9 7 9 2
65 3 1 13 13 10 9 0 1 10 9 1 10 9 0 1 10 9 2 10 9 3 13 13 10 9 0 1 10 9 2 3 7 10 9 13 1 9 1 9 7 1 9 1 10 9 0 2 3 7 3 1 9 0 7 1 9 2 9 0 2 9 7 9 0 2
5 0 9 2 12 2
29 10 11 11 1 11 2 11 2 2 13 10 9 10 15 13 10 9 7 9 1 11 1 11 0 2 9 7 9 2
4 13 15 13 2
23 1 10 11 11 15 13 10 0 9 1 10 9 1 10 9 11 7 10 9 1 10 9 2
17 16 15 4 13 16 10 9 2 3 9 2 13 9 1 10 9 2
24 1 10 9 2 10 9 15 13 1 9 7 9 7 13 1 9 1 10 9 0 1 10 9 2
22 11 11 13 10 12 9 1 10 9 2 16 4 13 1 12 9 13 1 3 1 15 2
22 10 9 13 10 9 1 10 9 0 2 7 10 9 1 10 9 1 11 11 1 11 2
40 10 9 15 4 13 12 9 3 1 10 9 2 16 10 9 2 0 1 10 9 2 13 1 10 9 1 16 1 10 0 4 13 1 10 9 0 1 9 0 2
13 11 2 1 11 11 2 13 0 3 1 10 9 2
41 3 2 1 15 16 3 13 10 9 1 9 1 10 0 9 1 9 2 9 7 0 9 2 10 11 11 13 1 10 9 10 9 11 11 1 10 3 0 9 0 2
34 10 0 7 0 9 15 13 10 9 1 16 1 10 0 9 13 10 9 3 15 13 10 0 9 1 9 7 9 0 16 13 1 15 2
29 7 7 1 0 9 1 10 11 11 1 10 9 1 10 11 11 11 12 7 1 11 1 10 9 11 11 11 12 2
16 13 10 9 1 10 0 9 1 11 1 10 0 9 1 12 2
37 10 9 1 9 11 15 13 1 12 9 2 13 1 9 2 9 7 15 2 1 9 0 11 2 1 10 9 1 9 2 8 2 8 2 8 2 2
27 10 9 1 10 9 13 10 9 1 10 10 9 1 9 1 10 9 2 11 2 7 10 9 2 11 2 2
17 13 9 2 9 2 9 2 9 2 7 15 13 1 10 9 0 2
31 13 16 10 9 1 10 9 13 0 7 15 13 13 1 10 9 3 3 7 10 9 13 0 2 10 9 4 13 1 11 2
37 1 9 2 16 13 10 9 2 13 3 1 12 9 1 13 15 16 3 15 13 10 9 2 5 12 2 16 15 13 3 10 2 9 1 9 2 2
17 10 0 9 1 10 9 11 13 10 9 11 1 0 9 1 9 2
55 11 4 13 16 10 9 0 13 1 10 9 0 1 10 9 1 11 1 10 0 9 1 9 2 13 1 10 12 13 1 10 9 1 10 11 2 2 3 13 9 0 2 0 2 16 15 4 13 7 13 1 10 9 2 2
38 13 13 16 10 9 7 9 15 13 1 9 0 2 13 16 1 10 3 10 9 13 10 9 3 0 2 1 15 15 15 13 9 2 0 2 7 0 2
63 3 11 15 13 1 10 9 1 11 13 1 10 9 15 13 1 10 9 2 7 15 13 1 10 9 1 10 9 11 2 2 10 11 1 10 9 2 8 1 15 0 1 10 9 1 9 3 1 11 2 3 15 13 12 9 13 9 7 13 1 10 9 2
24 11 3 13 13 1 3 9 10 0 9 16 13 1 13 12 9 2 15 13 7 13 10 9 2
68 15 13 0 1 10 9 1 10 9 3 0 1 9 1 11 11 2 10 11 11 2 7 10 11 2 7 13 13 0 1 10 9 2 9 16 15 13 1 10 9 1 12 10 11 11 1 11 11 1 11 11 2 10 9 0 1 11 11 1 9 1 10 9 1 11 11 2 2
11 9 1 11 1 10 11 11 2 11 1 11
16 10 9 1 10 9 3 13 15 16 13 0 1 10 0 9 2
21 3 10 9 1 10 9 15 13 1 10 9 7 15 1 15 13 9 1 10 9 2
35 10 9 13 1 13 10 9 0 3 16 13 10 9 1 9 1 10 9 1 11 2 1 3 15 13 9 7 9 0 2 1 9 7 9 2
34 11 4 13 10 9 1 9 7 9 1 11 2 13 1 10 9 1 11 1 10 11 2 11 2 11 11 2 1 15 13 1 12 9 2
24 15 13 1 9 1 10 9 1 9 0 7 9 0 16 15 13 1 9 13 1 9 0 0 2
13 10 9 16 15 13 15 13 3 11 1 10 11 2
23 11 11 2 11 2 12 1 11 1 12 2 13 10 0 2 9 0 16 15 13 1 9 2
27 3 2 3 2 4 13 15 1 10 9 16 4 4 13 1 10 0 2 9 2 1 9 1 9 1 9 2
49 10 9 11 11 15 4 13 1 10 11 11 10 12 9 1 9 2 10 9 0 13 13 1 13 15 15 2 10 9 13 15 1 10 9 1 11 7 13 9 16 10 9 13 1 3 1 10 9 2
27 10 9 1 10 9 13 10 9 0 1 10 9 1 11 1 11 1 12 2 7 13 11 1 10 11 11 2
28 1 12 14 1 10 11 11 7 12 9 3 3 13 13 10 9 1 11 1 15 15 13 1 10 11 11 11 2
26 11 12 13 1 13 15 11 11 2 9 1 10 9 2 1 4 1 13 11 11 2 9 1 11 2 2
7 13 10 9 1 11 11 2
43 1 10 9 1 11 2 11 13 1 10 9 2 11 11 2 2 13 10 9 1 11 1 10 15 0 2 1 9 1 10 9 1 16 4 13 1 10 9 0 1 10 11 2
25 10 9 13 13 10 9 0 1 11 2 1 10 15 15 13 10 9 0 0 1 10 11 11 11 2
29 9 2 10 9 0 2 10 9 1 10 9 13 10 9 10 12 1 11 1 12 7 13 10 9 0 1 10 9 2
30 1 10 9 2 13 13 1 3 16 1 10 9 0 1 11 3 15 13 9 0 1 2 13 1 13 2 1 10 9 2
56 10 9 1 10 9 13 1 1 12 9 1 9 13 1 9 1 10 11 2 11 2 11 2 9 0 2 11 2 11 11 2 9 0 7 1 13 10 9 1 9 0 2 16 13 1 3 1 10 12 1 12 1 10 9 0 2
41 1 10 9 1 10 12 9 2 15 13 1 15 3 0 2 13 1 10 9 1 10 9 2 10 0 9 13 1 10 9 11 11 2 1 10 0 9 1 10 11 2
65 13 2 1 15 2 1 10 9 0 1 9 0 2 10 9 4 3 13 2 13 10 9 1 10 9 1 10 9 2 9 2 9 7 9 15 13 3 13 2 16 13 1 9 10 9 1 10 9 2 10 9 2 10 9 7 10 9 1 10 9 1 10 9 0 2
26 3 13 9 1 9 7 10 9 0 16 4 13 10 9 1 2 9 16 13 10 9 7 9 0 2 2
17 10 9 13 16 15 13 0 9 7 15 1 10 9 3 13 9 2
34 10 10 9 13 9 2 15 16 13 10 9 3 0 16 13 1 9 3 7 10 9 3 13 2 13 3 7 13 10 9 1 15 0 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
21 1 12 13 1 11 2 7 3 12 13 1 10 9 2 16 3 13 3 10 9 2
60 11 11 2 11 1 10 11 2 11 1 10 11 2 12 2 11 11 2 11 2 12 1 11 1 12 2 2 9 0 16 13 10 9 3 0 1 10 9 1 10 11 1 10 9 1 10 9 1 10 11 2 13 10 9 1 11 7 10 9 2
22 10 11 1 10 11 13 10 9 0 16 13 9 1 10 9 1 11 11 2 11 11 2
49 11 2 16 4 4 13 10 9 1 10 9 0 2 13 10 9 1 9 1 12 2 3 15 13 16 13 10 9 0 0 1 10 9 1 9 0 1 9 0 7 9 0 1 9 1 13 10 9 2
26 11 0 2 9 1 9 2 9 7 9 1 9 2 13 9 1 0 9 1 15 16 15 13 9 0 2
35 13 10 9 1 10 9 15 13 11 12 1 10 9 1 12 1 16 15 13 10 0 9 1 10 9 1 10 11 11 1 10 11 1 11 2
38 11 2 10 2 11 13 10 9 7 9 0 2 1 10 9 1 11 2 11 2 9 1 11 2 1 10 9 1 11 2 1 2 11 7 9 1 11 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
13 1 9 1 15 2 10 9 13 10 9 1 11 2
9 10 9 0 13 9 13 1 9 2
18 3 1 9 2 13 1 11 11 7 11 11 1 11 1 12 2 12 2
60 7 3 15 13 1 10 9 1 2 9 2 3 1 12 9 2 1 15 11 11 2 11 11 11 2 11 11 11 7 11 11 2 2 11 11 7 11 11 11 13 10 9 3 3 0 2 13 15 1 10 9 0 2 0 7 1 10 9 0 2
46 1 10 9 1 10 9 2 10 9 0 13 1 10 9 3 0 1 11 2 15 1 9 1 1 9 1 10 9 1 10 9 11 11 2 10 11 11 13 1 10 0 9 1 10 9 2
32 15 13 16 10 9 1 11 13 1 10 9 0 8 2 2 9 2 2 7 8 2 13 2 1 15 15 13 2 9 0 2 2
14 10 9 1 10 11 15 13 1 10 9 0 1 11 2
15 13 10 9 1 11 11 2 10 9 0 3 1 10 11 2
47 0 2 9 0 16 13 3 9 2 3 13 9 7 1 15 13 0 7 3 13 9 2 15 9 10 9 16 13 0 16 1 13 15 1 9 1 12 9 13 9 7 15 9 10 15 15 2
22 4 13 1 10 11 9 0 2 10 9 0 1 9 2 1 10 9 11 1 10 11 2
17 11 11 13 10 9 7 9 0 2 13 10 12 1 11 1 12 2
17 10 9 3 4 13 7 10 9 1 10 9 15 13 1 10 9 2
28 10 8 4 3 13 1 7 3 1 10 9 1 9 1 13 7 13 10 9 0 7 3 10 9 0 1 9 2
26 7 3 2 1 10 9 13 1 2 11 11 15 11 2 15 4 13 10 9 16 15 13 1 10 9 2
44 10 11 11 11 11 12 13 3 10 9 1 10 0 9 1 9 1 9 3 7 13 12 9 15 16 13 10 12 2 12 9 1 10 9 7 10 12 2 12 9 1 10 9 2
14 3 13 3 1 12 9 1 10 10 12 9 1 9 2
16 3 3 3 15 13 10 9 7 10 9 1 10 9 7 9 2
61 2 10 9 4 13 1 9 10 0 9 1 10 9 1 13 16 10 9 7 10 9 2 4 13 3 2 13 10 9 11 11 1 11 1 10 13 2 13 1 10 9 2 10 9 11 11 1 11 2 1 13 10 11 1 10 11 11 1 10 9 2
17 11 11 13 1 10 11 11 2 11 2 10 12 1 11 1 12 2
20 10 9 2 13 3 0 7 0 2 10 9 13 1 10 9 7 13 3 0 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
11 10 9 15 13 13 1 10 9 1 11 2
21 15 13 0 13 15 1 10 9 1 9 16 10 9 11 13 1 10 9 1 9 2
21 10 8 11 11 11 13 10 9 1 10 0 9 7 10 9 3 0 7 3 9 2
51 10 11 3 15 13 0 1 10 11 11 2 16 10 9 1 10 0 9 13 10 9 1 12 9 13 1 10 11 7 15 13 10 9 1 10 9 7 13 1 13 1 10 9 1 10 9 1 10 11 11 2
24 1 15 9 3 13 10 9 2 3 1 2 13 2 2 2 9 2 2 7 2 3 0 2 2
35 1 10 9 1 10 9 2 13 9 1 9 1 10 9 1 11 1 11 1 10 9 1 10 9 1 10 12 7 10 12 1 11 1 12 2
20 2 2 16 10 9 3 13 10 9 2 2 3 1 15 15 4 13 2 2 2
36 3 13 16 13 1 10 9 2 10 9 2 10 9 7 10 9 1 10 9 2 7 10 9 1 15 2 7 3 3 15 4 13 10 9 3 2
25 10 9 4 0 1 15 9 1 10 9 0 1 12 9 1 9 16 13 10 9 1 2 9 2 2
24 1 9 1 11 13 9 0 3 1 12 9 7 1 10 9 1 11 11 7 11 1 12 9 2
40 10 9 1 10 9 1 9 7 9 1 11 1 12 13 1 10 9 11 2 12 2 12 2 1 10 12 2 12 2 9 13 1 9 1 9 1 10 9 11 2
24 15 3 0 13 10 9 1 9 1 11 10 9 4 13 1 11 11 3 12 9 13 1 11 2
13 11 11 13 10 9 0 1 10 9 1 11 11 2
32 11 11 13 10 9 0 1 10 9 1 11 1 10 8 11 2 1 15 13 10 9 1 10 11 11 2 10 9 1 9 0 2
27 3 3 10 9 1 9 3 0 1 9 0 7 3 13 3 13 10 9 1 9 7 10 9 1 10 9 2
110 10 9 2 4 13 1 10 9 1 10 10 9 0 2 11 2 11 11 2 10 11 16 13 1 10 9 16 10 9 1 9 4 13 10 9 1 9 1 10 11 11 2 1 10 15 15 13 10 9 1 13 15 2 15 1 10 9 8 9 1 10 9 13 10 9 1 10 9 1 11 11 1 11 2 9 11 11 11 11 7 3 16 10 9 0 0 2 4 13 1 11 2 3 16 10 9 13 9 1 10 9 7 9 0 13 1 9 7 9 2
30 10 0 9 1 10 9 1 9 1 10 9 13 15 15 4 13 10 9 1 10 9 9 1 9 7 1 9 0 9 2
36 2 13 9 1 10 9 1 9 16 10 9 4 13 2 2 13 10 9 2 16 13 9 1 10 11 11 2 15 1 10 9 13 10 9 0 2
20 10 12 1 11 1 12 4 13 10 11 1 11 7 15 13 10 12 1 11 2
37 10 9 0 13 10 9 1 10 9 1 13 9 13 1 10 9 1 10 9 11 11 2 16 13 10 9 1 10 9 0 0 1 10 11 11 11 2
45 3 1 13 10 9 0 1 10 9 2 11 15 13 1 10 9 0 7 0 2 10 9 0 1 15 15 13 10 9 7 10 9 16 13 9 1 9 1 9 1 10 11 7 11 2
24 11 13 10 9 0 2 16 13 10 0 9 10 12 1 11 1 12 7 15 13 1 9 0 2
55 13 1 10 9 0 16 15 13 2 11 4 13 16 1 10 2 9 2 1 10 9 2 13 0 16 10 9 13 1 10 11 2 1 10 9 3 0 3 1 13 0 16 13 15 16 4 13 10 9 1 10 12 9 2 2
28 7 13 1 9 1 10 9 7 1 10 9 1 0 9 16 13 1 15 10 9 13 13 13 7 13 10 9 2
22 10 11 11 13 10 0 9 1 9 0 16 4 13 1 12 5 2 12 9 1 9 2
40 10 9 0 2 16 4 13 10 0 9 1 9 1 10 9 1 10 9 2 13 10 9 0 12 9 2 16 7 10 9 1 9 7 9 13 12 9 1 9 2
41 16 11 13 10 0 9 1 9 2 10 0 9 13 10 9 7 9 1 10 9 16 13 1 10 9 0 2 7 3 13 1 13 1 11 7 1 10 9 1 9 2
36 11 13 15 1 10 9 1 9 3 0 1 10 9 2 16 1 10 12 13 1 12 5 2 7 13 3 3 12 9 10 12 9 1 10 9 2
12 11 11 13 0 9 1 10 9 0 1 10 11
33 1 9 1 10 9 1 11 0 2 1 12 7 12 9 2 1 9 0 16 15 13 1 10 11 2 13 10 9 1 9 0 9 2
29 10 9 1 10 9 1 10 9 0 7 9 0 11 11 11 1 10 11 7 1 11 11 1 11 2 1 9 0 2
21 1 10 9 2 10 9 13 13 1 0 9 1 10 9 2 1 9 7 9 0 2
31 3 2 1 10 9 16 13 10 9 1 10 9 7 10 9 15 13 9 0 2 15 15 4 13 10 9 0 1 10 9 2
28 10 11 1 10 11 13 10 9 2 1 9 7 11 15 13 1 10 9 1 9 13 1 9 7 13 1 13 2
30 15 1 10 9 1 10 9 13 10 9 1 10 9 0 1 9 1 10 9 0 7 1 10 9 2 3 0 7 0 2
17 11 13 10 9 1 10 9 1 11 2 1 10 9 0 1 11 2
20 9 0 2 9 2 9 7 9 2 2 7 15 1 9 1 9 0 2 0 2
26 1 9 1 16 10 9 7 10 9 0 13 10 9 1 11 2 1 10 0 9 15 4 4 13 3 2
55 1 9 2 15 13 10 9 1 9 3 1 10 9 0 2 7 10 9 1 13 1 9 0 10 9 1 10 9 1 10 9 1 10 9 2 15 16 13 10 9 7 9 1 10 9 3 1 13 10 9 1 10 0 9 2
3 10 9 2
44 10 9 2 11 11 11 11 11 15 2 13 10 9 2 11 1 11 11 2 16 3 13 1 10 9 2 7 16 3 15 4 1 13 2 16 13 15 1 10 9 1 15 0 2
17 16 13 1 11 13 1 9 1 10 11 11 7 13 9 1 9 2
32 13 9 1 9 2 9 1 10 9 0 1 10 0 9 0 2 9 1 10 11 9 0 1 10 9 0 9 1 9 7 9 2
23 10 9 13 16 15 13 10 15 13 15 16 3 13 10 9 2 7 1 9 13 10 9 2
14 4 13 11 11 2 13 1 16 3 4 4 3 0 2
11 15 13 10 9 5 12 1 10 11 11 2
17 11 7 11 11 2 10 9 9 1 11 2 15 13 1 10 11 2
62 1 15 2 1 10 9 2 10 9 7 10 9 1 11 2 3 13 10 0 9 1 10 9 15 13 10 9 0 2 13 7 13 2 16 3 4 13 10 9 1 11 16 15 13 9 1 10 9 2 10 9 7 10 9 0 7 0 3 13 1 11 2
32 3 2 1 15 15 13 10 9 0 2 7 16 1 15 3 2 9 1 9 2 2 13 10 9 1 10 9 1 10 9 0 2
8 15 13 1 10 11 1 11 2
30 1 13 10 9 1 9 2 15 15 4 13 1 11 10 9 1 10 9 7 13 0 1 10 9 15 10 9 13 13 2
27 13 9 1 10 9 1 13 15 7 13 1 10 9 2 7 3 13 1 9 1 11 13 1 11 1 12 2
27 10 9 13 1 3 1 12 9 1 9 7 13 10 9 1 13 9 1 10 9 1 9 0 1 9 0 2
28 10 9 1 10 9 1 10 16 11 4 13 15 10 9 16 4 13 0 1 10 0 9 2 10 9 1 9 2
15 13 10 9 3 7 4 13 1 10 9 10 9 1 9 2
7 10 9 13 1 10 11 2
21 1 15 15 13 9 1 10 10 9 7 9 2 3 9 2 9 2 9 7 9 2
22 4 7 13 10 9 3 1 10 9 7 15 13 16 10 9 1 9 3 13 1 9 2
17 3 7 10 9 1 9 1 10 9 1 9 15 13 1 10 9 2
46 1 10 9 1 10 9 3 1 11 7 1 10 0 9 0 10 9 13 10 9 0 2 13 3 1 13 10 9 1 10 9 2 11 2 16 13 1 10 9 1 2 11 11 11 2 2
70 10 9 0 1 15 10 9 4 13 10 9 0 1 10 2 9 1 9 2 2 13 10 9 1 9 2 10 0 9 7 10 9 0 0 1 10 9 7 2 7 9 2 16 15 4 13 3 2 0 1 10 3 0 9 1 11 11 11 7 1 9 0 7 2 7 9 0 2 3 2
32 10 11 13 9 1 9 1 10 9 2 15 16 15 13 13 10 12 9 2 3 1 10 12 9 0 1 10 9 8 2 8 2
16 1 12 2 10 9 4 13 1 11 7 4 13 11 2 12 2
29 10 9 13 15 13 1 9 1 10 11 1 11 1 11 1 11 7 1 10 11 1 11 1 10 11 1 10 11 2
53 1 10 9 12 2 2 2 11 11 11 11 2 7 10 9 1 9 1 10 0 9 2 13 1 11 11 1 10 0 9 0 16 13 13 2 3 2 10 9 11 11 12 7 11 12 2 10 3 0 1 11 11 2
9 10 9 4 13 1 10 9 0 2
22 0 2 11 13 1 10 9 1 11 1 13 1 11 2 15 15 4 13 1 10 9 2
11 3 1 0 10 1 12 13 10 0 9 2
78 3 2 16 3 15 13 16 10 9 13 9 2 10 0 11 2 1 10 9 16 1 0 9 1 10 9 2 1 10 9 3 0 2 1 11 2 10 11 11 2 4 13 2 15 13 10 9 7 9 1 10 9 1 10 8 9 1 11 2 7 15 13 0 2 1 3 13 10 9 3 7 1 10 0 9 1 11 2
20 10 9 13 3 0 1 16 13 10 9 1 9 1 9 16 15 13 3 3 2
20 13 10 12 9 2 1 10 9 1 11 2 7 15 13 10 9 16 13 9 2
20 13 10 12 1 11 1 12 2 11 11 4 1 13 15 1 10 9 1 12 2
34 11 11 13 10 9 1 12 9 2 12 9 2 1 10 9 12 9 13 1 9 0 2 13 1 10 12 11 11 11 2 11 2 11 2
22 1 11 1 10 11 13 12 9 2 12 0 2 7 12 9 0 1 9 0 7 0 2
10 10 0 9 1 10 11 1 11 13 2
14 13 10 9 1 13 1 10 9 7 1 10 10 9 2
26 10 12 1 11 1 10 9 2 10 9 11 11 13 10 9 1 10 9 1 10 11 1 10 11 11 2
44 1 15 2 10 9 4 7 13 10 9 1 13 10 9 2 3 1 10 9 1 11 3 1 0 15 13 10 0 9 2 16 15 13 1 11 1 10 9 1 10 11 1 11 2
26 13 0 9 2 9 2 9 2 9 2 3 1 9 0 0 1 10 9 1 10 11 1 11 1 11 2
20 14 2 15 4 13 10 9 1 11 2 10 11 11 8 8 2 7 3 0 2
51 15 13 10 9 1 9 7 10 9 3 13 3 0 1 0 2 7 1 0 13 15 3 0 2 13 16 0 2 16 15 13 1 10 9 1 3 1 13 15 9 0 13 15 16 15 13 0 7 10 9 2
22 16 11 13 9 1 10 9 0 2 13 10 9 1 11 13 10 15 16 13 1 9 2
10 13 10 9 1 9 2 3 1 9 2
7 10 9 11 11 11 11 2
70 10 9 13 1 15 10 9 1 13 1 13 15 9 1 10 9 1 11 7 1 9 16 10 9 13 1 9 1 10 9 13 1 10 9 0 2 4 13 1 10 9 0 2 3 13 13 15 1 0 2 3 16 10 16 13 3 7 16 3 13 15 16 13 3 1 15 2 15 13 2
24 10 9 13 1 10 13 15 10 9 3 13 10 9 1 9 1 10 9 7 9 1 10 9 2
13 1 9 2 15 15 13 3 1 10 9 1 9 2
56 13 10 0 9 1 10 9 1 10 9 11 2 1 10 15 4 13 1 9 1 10 12 2 16 10 9 0 2 11 10 11 7 10 9 10 11 11 1 11 2 4 13 1 10 9 0 2 11 2 1 10 15 3 13 9 2
23 3 2 16 13 10 9 0 1 15 1 11 13 10 9 3 0 1 10 9 1 10 9 2
38 13 16 2 1 9 0 2 16 10 9 13 3 13 16 3 13 7 3 13 10 9 0 2 2 15 9 13 16 10 9 15 13 1 10 9 0 2 2
61 10 12 9 7 9 0 1 12 9 13 1 10 9 2 9 2 13 1 10 12 1 10 12 1 11 1 11 2 11 2 1 10 9 2 10 9 1 9 2 2 1 10 15 11 12 15 13 1 2 13 10 0 9 1 10 9 1 9 0 2 2
29 10 9 1 9 0 13 1 10 12 9 1 10 11 11 15 13 3 1 10 9 2 7 13 1 9 10 9 0 2
15 13 9 7 9 2 1 11 11 7 13 10 9 1 11 2
19 1 9 0 1 10 11 2 16 13 1 12 9 2 10 9 13 12 9 2
17 3 2 10 9 1 9 1 10 11 11 4 13 1 12 7 12 2
22 10 9 0 7 10 0 9 15 13 1 10 9 0 1 9 1 10 9 1 10 9 2
31 11 7 11 2 10 9 0 0 1 10 11 11 7 3 0 2 4 13 1 12 1 10 9 1 10 9 1 9 1 11 2
10 4 13 10 9 1 12 9 2 5 2
17 10 9 1 9 11 11 13 9 1 9 1 11 10 9 1 3 2
20 1 10 15 15 4 13 7 13 1 11 2 15 13 10 9 7 1 9 0 2
40 10 0 9 1 13 15 10 9 3 0 7 1 13 15 10 9 2 13 15 16 13 1 2 9 2 0 2 1 0 10 9 2 16 10 15 16 13 13 0 2
34 1 9 1 11 10 9 13 13 10 9 1 10 9 0 1 10 9 0 13 1 10 9 7 10 15 4 13 1 10 9 11 1 11 2
30 10 9 0 1 10 9 4 13 1 10 9 1 10 11 11 1 11 7 1 9 1 9 1 11 7 1 10 10 9 2
25 1 11 11 2 10 9 16 15 13 13 12 9 1 10 9 7 10 12 9 1 9 1 10 9 2
43 10 9 13 3 16 9 3 1 10 9 15 13 1 10 9 1 10 9 10 9 1 10 9 2 10 9 1 9 1 10 9 7 10 9 1 10 9 0 1 10 9 0 2
37 11 12 2 1 10 9 2 16 3 4 13 13 1 11 1 10 9 0 1 10 9 1 10 9 12 2 4 13 9 1 9 1 10 9 1 11 2
43 3 2 4 13 16 10 9 1 10 9 1 10 0 9 1 12 4 13 1 13 9 1 10 9 2 2 10 11 4 13 1 10 9 1 10 0 9 2 7 3 13 9 2
54 10 11 8 13 10 9 1 9 13 1 11 1 10 11 11 1 10 11 2 11 11 1 11 11 2 3 11 2 11 7 11 2 2 13 15 1 10 9 8 1 10 11 11 7 11 1 9 1 10 9 1 10 9 2
36 1 10 9 0 1 15 13 10 9 1 10 9 1 10 9 1 9 2 0 1 0 9 11 1 12 9 2 7 13 1 10 9 7 1 9 2
42 10 9 1 10 9 0 1 11 13 1 13 1 10 9 12 2 16 10 11 11 1 11 13 10 9 1 10 9 1 9 1 10 9 1 10 9 0 1 10 9 0 2
25 10 0 9 13 9 1 11 2 1 10 15 10 9 1 10 9 16 13 10 11 11 15 4 13 2
41 1 12 2 10 0 9 0 1 11 15 13 1 15 15 1 2 11 2 1 2 11 2 2 10 9 1 9 16 13 1 10 9 1 12 2 12 2 12 7 12 2
31 10 11 11 7 11 11 2 0 11 2 2 3 13 1 10 11 11 2 13 10 9 0 1 10 10 9 1 10 9 9 2
38 10 0 9 1 9 2 9 7 9 1 10 9 1 9 2 1 10 9 2 1 10 9 1 9 1 13 15 1 9 7 1 10 9 1 10 13 9 2
18 10 9 4 13 11 11 2 9 1 9 1 9 9 1 10 9 11 2
21 1 12 11 16 4 10 9 7 15 13 10 0 9 3 15 13 13 10 0 11 2
31 1 9 2 10 9 13 10 9 1 9 3 0 2 1 0 2 10 9 0 1 10 9 1 11 2 11 4 13 3 0 2
32 10 9 13 1 9 0 1 0 9 1 10 9 7 15 13 1 10 9 1 10 9 16 13 10 9 7 13 13 1 10 11 2
8 10 12 9 0 2 12 2 2
52 10 9 11 13 1 10 9 1 10 11 11 7 4 13 10 9 1 10 0 9 2 3 1 10 12 4 13 10 9 1 11 2 9 1 11 15 13 10 9 1 10 9 7 13 3 1 10 9 1 10 9 2
16 10 9 13 2 10 15 1 15 4 13 1 10 9 7 13 2
38 3 1 10 9 2 15 13 10 9 3 1 9 13 1 11 11 2 10 9 1 11 2 2 13 10 9 1 10 9 0 2 7 15 13 12 1 13 2
43 1 9 1 10 9 2 10 9 13 10 9 3 0 1 15 15 13 1 10 9 0 2 3 16 10 9 13 0 3 7 13 10 0 9 0 1 10 9 1 10 9 0 2
11 3 13 1 9 7 9 2 13 10 9 2
31 10 9 16 15 13 1 10 9 1 10 9 11 7 11 13 2 3 2 10 9 0 1 3 9 1 10 9 1 10 11 2
30 10 9 10 9 15 13 9 1 10 11 1 10 11 1 10 13 1 10 9 1 10 11 1 11 1 12 9 1 12 2
24 15 13 1 10 9 0 13 1 10 9 13 2 1 10 15 15 13 10 9 1 10 9 0 2
27 1 15 13 10 9 2 13 1 10 9 0 12 9 1 9 2 16 15 7 10 9 1 9 13 10 9 2
29 16 15 15 13 1 10 9 2 15 13 3 0 7 15 13 3 1 10 9 7 3 13 1 15 1 10 0 9 2
44 1 11 2 15 13 12 9 2 1 9 7 9 2 10 15 15 13 1 10 12 9 1 10 9 0 1 11 2 7 12 9 13 1 10 9 1 10 9 1 13 9 1 9 2
24 10 9 4 4 13 1 0 9 1 10 9 1 10 15 4 13 2 11 1 11 7 11 12 2
21 3 13 3 10 10 9 0 2 3 10 9 13 1 9 7 9 7 1 9 0 2
35 3 2 10 9 0 13 9 0 1 10 0 9 0 2 16 15 4 13 1 15 3 0 2 16 15 13 3 0 7 15 13 1 10 9 2
29 11 4 13 1 9 1 11 2 11 15 13 16 13 10 11 2 7 10 9 15 13 3 3 1 10 9 1 9 2
53 3 13 10 9 16 13 10 9 7 13 1 10 9 1 10 9 16 1 11 2 11 11 1 11 2 11 2 11 2 11 1 10 0 1 10 9 0 7 10 0 2 7 13 3 1 10 9 1 10 11 1 11 2
49 13 9 1 10 9 11 11 2 15 3 13 0 9 1 10 9 0 2 7 1 10 9 11 11 11 2 8 2 2 9 1 10 9 1 11 11 2 12 2 2 9 0 7 0 7 0 9 0 2
15 10 0 9 1 9 1 10 9 11 13 1 10 0 9 2
56 10 9 1 10 9 13 1 10 9 1 10 9 1 15 1 10 9 2 10 9 11 2 15 13 10 9 1 10 9 2 9 0 1 9 1 13 0 9 1 9 1 9 0 1 10 9 1 11 1 10 9 1 10 9 0 2
27 1 9 2 10 9 11 11 2 11 11 7 11 2 1 12 1 10 12 9 0 2 13 10 0 9 0 2
26 10 9 7 10 9 1 10 10 9 15 1 10 9 0 1 11 1 13 10 0 9 1 10 10 9 2
24 3 1 10 11 11 0 2 10 9 0 1 11 15 13 1 10 9 9 7 9 1 10 9 2
20 11 11 13 10 9 0 2 1 13 2 3 10 9 7 9 13 1 10 9 2
10 3 13 3 10 9 1 10 11 11 2
47 10 11 4 13 10 9 1 9 1 11 1 10 9 1 10 9 2 7 4 13 3 3 1 10 11 11 7 10 9 4 13 1 0 1 9 1 15 1 10 11 11 7 1 10 11 11 2
62 11 13 3 13 1 11 1 13 15 1 10 9 1 9 1 13 10 9 1 10 15 15 9 4 13 2 7 11 15 13 1 13 15 2 1 9 11 2 16 3 13 15 0 16 13 10 9 15 13 16 13 10 9 0 1 13 10 9 1 10 9 2
14 10 0 9 4 13 3 1 10 9 1 10 9 0 2
19 11 13 10 0 9 1 9 1 10 9 1 11 7 1 0 1 10 11 2
26 1 10 9 1 9 1 10 9 0 1 12 2 13 9 1 10 9 1 10 11 1 10 9 1 11 2
17 10 9 0 13 9 3 9 1 4 13 0 2 13 2 1 9 2
13 10 9 13 9 1 10 9 1 16 10 9 13 2
15 1 10 9 0 13 10 9 1 12 9 1 12 9 0 2
21 1 4 13 1 9 2 15 15 13 9 7 9 7 4 13 7 13 1 9 0 2
29 1 11 1 12 13 10 11 1 11 7 13 3 1 11 11 7 13 3 3 1 11 11 16 13 10 9 1 11 11
6 15 9 3 13 0 2
8 2 10 10 9 13 1 9 2
61 10 9 0 7 0 13 10 9 3 0 1 11 2 3 1 10 9 1 13 9 1 9 0 1 10 9 0 2 1 15 10 9 2 2 9 15 16 13 10 0 9 1 11 2 13 7 15 13 1 9 1 9 0 1 10 9 2 2 13 11 2
37 1 10 0 9 1 10 11 11 2 1 11 7 10 9 1 10 11 1 11 2 3 3 15 13 1 11 11 2 10 9 16 13 1 10 9 0 2
18 10 9 1 11 13 1 9 1 10 9 1 11 11 1 11 1 9 2
50 10 12 1 11 1 12 2 1 10 12 5 9 1 10 9 1 9 1 10 12 9 0 1 11 11 1 12 2 10 9 11 11 4 1 13 10 9 1 11 11 1 10 9 1 11 2 11 7 11 2
7 11 11 13 10 0 9 2
22 4 13 9 1 10 11 11 11 1 10 9 11 11 11 1 11 2 1 10 9 13 2
57 13 10 9 0 1 9 16 13 9 0 1 9 2 0 1 12 1 12 9 0 1 9 0 16 13 1 9 1 10 9 0 1 12 1 12 5 1 0 2 7 1 12 1 12 9 0 1 9 9 0 16 13 12 5 1 9 2
15 3 2 13 1 9 1 10 15 15 4 13 9 1 9 2
21 13 1 10 9 1 10 9 7 10 9 1 10 11 11 1 11 7 10 11 0 2
14 3 13 10 9 2 9 16 3 3 13 10 9 0 2
22 0 9 13 1 10 13 9 16 15 4 13 3 1 10 13 1 10 9 3 3 13 2
17 15 9 13 16 2 10 9 2 11 11 4 13 11 1 10 9 2
56 11 1 10 11 13 10 15 1 10 9 1 10 0 9 1 10 9 0 2 9 2 9 0 1 13 9 7 9 2 1 10 15 13 1 9 3 0 1 9 1 9 0 1 9 2 16 13 15 1 10 15 1 10 0 9 2
36 10 9 3 13 10 9 1 10 9 0 1 13 9 0 2 0 1 9 2 9 1 9 2 9 0 2 9 1 10 9 7 9 2 1 15 2
26 1 10 0 9 2 0 9 13 15 1 10 9 1 0 9 1 9 2 15 15 0 1 10 9 0 2
15 13 10 9 0 2 11 11 2 11 11 7 11 11 2 2
8 15 13 1 10 9 1 9 2
28 10 9 1 11 13 1 10 9 10 12 1 11 1 12 7 10 9 1 11 15 13 10 12 1 11 1 12 2
24 1 10 9 2 13 1 13 10 9 0 2 0 7 3 7 2 1 10 9 2 15 13 0 2
17 1 10 9 15 13 10 9 1 10 9 16 13 10 9 1 9 2
37 1 10 9 13 10 9 2 7 4 1 13 1 10 9 0 2 2 10 9 2 2 2 1 10 9 1 13 10 9 16 15 4 13 1 9 0 2
23 1 10 9 1 8 8 13 15 9 2 1 10 9 8 3 1 9 2 7 10 9 3 2
22 1 13 1 10 9 4 10 12 0 1 13 0 9 13 1 10 10 9 1 10 9 2
25 1 12 15 13 10 9 13 1 12 9 0 13 1 9 1 10 9 1 10 9 1 11 1 12 2
36 1 10 9 1 10 9 2 10 9 1 11 13 1 10 9 0 7 15 13 1 10 9 1 10 9 0 1 10 9 1 10 9 1 10 9 2
16 1 12 13 10 0 9 1 10 9 1 10 9 1 10 9 2
22 1 10 12 9 13 10 0 9 1 9 7 3 13 8 5 1 9 2 11 11 2 2
44 10 9 1 9 0 1 11 13 9 0 1 10 11 11 2 7 13 10 9 1 9 0 16 13 13 9 1 11 2 11 2 11 2 11 11 2 8 1 10 0 9 1 9 2
20 10 9 1 9 9 1 9 13 1 12 7 10 9 9 1 9 13 1 12 2
24 9 0 2 13 9 1 10 9 1 9 2 9 7 9 2 9 1 10 11 11 1 10 9 2
14 15 13 3 10 9 1 9 1 9 7 9 1 9 2
23 10 9 0 11 11 4 13 1 10 9 1 10 9 0 0 1 10 9 1 9 7 9 2
20 0 9 1 11 13 10 0 9 1 9 2 9 7 9 0 0 1 10 9 2
35 1 10 11 4 13 10 9 1 3 13 2 10 9 1 10 9 2 7 4 13 1 16 10 9 1 9 0 2 3 4 1 4 13 2 2
25 10 8 1 11 1 10 11 2 11 4 13 10 9 8 16 4 4 13 1 10 9 16 15 13 2
67 10 11 13 10 9 1 10 9 13 1 9 16 10 9 13 10 9 1 10 9 1 10 16 4 13 9 0 0 16 4 13 1 9 2 9 2 9 2 9 2 9 2 2 3 1 16 10 9 15 13 7 13 10 0 9 1 9 2 1 10 13 3 0 10 9 0 2
32 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 9 2 1 10 9 1 11 2 11 7 9 1 11 2 11 2
35 1 12 2 10 9 0 13 1 10 11 1 13 10 0 9 2 13 10 9 1 10 9 1 10 0 9 1 13 10 9 0 1 10 9 2
16 13 1 11 1 10 11 2 9 2 1 10 11 11 1 11 2
27 1 9 1 10 9 12 2 11 15 13 1 10 9 1 9 1 0 9 1 10 9 0 1 10 11 11 2
40 1 15 15 4 13 1 10 9 0 1 10 9 2 13 1 9 2 9 9 2 9 2 9 2 9 0 1 9 7 9 1 12 9 1 10 9 1 10 9 2
7 13 9 1 10 11 11 2
36 1 10 9 16 13 10 9 1 10 9 0 11 11 11 11 1 12 2 11 13 16 4 13 13 1 10 9 16 13 10 9 1 2 0 2 2
27 1 12 13 10 9 1 10 13 15 10 9 1 11 2 11 11 11 2 10 9 15 13 10 11 1 11 2
21 4 4 13 12 9 2 10 11 11 11 2 7 10 11 11 7 11 2 3 0 2
11 11 13 10 9 1 11 2 11 2 11 2
16 1 10 9 1 10 8 8 2 15 13 1 10 11 2 11 2
30 1 10 0 9 1 10 9 10 13 3 1 10 9 1 10 9 13 1 10 0 7 0 9 4 4 13 10 9 0 2
46 1 12 11 11 13 1 10 9 11 12 2 3 1 10 9 11 11 11 11 11 2 3 13 10 9 1 10 0 9 7 1 10 9 1 10 9 13 9 1 10 9 11 1 11 11 2
39 1 10 9 2 15 13 1 10 9 1 10 9 1 16 10 9 1 10 9 1 11 13 16 13 10 9 1 10 9 16 13 10 9 1 10 9 1 9 2
10 1 10 9 2 10 9 4 13 9 2
17 10 9 15 13 0 1 10 9 0 8 12 2 8 2 11 11 2
13 10 9 4 13 1 12 9 1 11 11 11 11 2
4 13 12 9 2
20 10 9 0 15 13 1 15 2 16 11 13 1 9 1 11 2 10 0 9 2
17 11 13 10 9 1 10 9 11 16 13 1 10 0 9 1 11 11
25 13 1 10 0 9 2 3 15 4 13 15 15 13 1 9 1 12 9 1 9 2 9 7 9 2
36 10 9 1 11 11 11 3 13 1 11 1 2 10 11 2 13 10 9 7 9 1 10 9 1 10 9 1 9 0 1 10 11 11 2 11 2
31 16 2 1 10 9 1 10 9 0 2 10 9 4 13 4 13 10 9 1 10 9 2 15 4 4 13 15 1 9 0 2
17 11 11 13 9 1 9 1 0 9 16 15 13 1 10 9 0 2
54 1 10 9 16 13 1 10 8 10 0 9 1 10 9 13 2 10 9 8 1 12 9 1 0 9 2 9 8 2 8 1 8 2 8 1 8 7 10 9 0 0 1 11 7 10 9 13 15 9 2 3 12 9 2
26 15 13 1 10 9 0 7 9 1 11 2 10 11 2 7 11 7 13 10 9 0 1 10 9 0 2
38 11 2 11 2 1 2 11 2 11 2 11 2 1 10 2 11 1 9 2 13 10 9 0 2 13 1 10 9 1 10 11 7 11 7 10 9 11 2
38 3 10 9 1 10 12 8 3 15 13 1 10 9 1 10 9 2 16 3 15 4 0 2 7 7 15 4 13 13 1 9 7 9 2 9 2 8 2
46 2 1 10 9 2 13 15 15 1 10 9 1 11 2 1 15 3 15 15 4 13 15 2 2 4 13 1 10 4 13 1 10 9 1 10 9 1 9 0 1 10 9 1 10 9 2
5 10 9 13 0 2
13 10 9 1 9 13 1 12 8 2 2 9 8 2
25 10 9 1 11 2 13 1 10 9 1 10 11 10 9 1 11 2 7 15 13 1 10 11 11 2
17 1 9 15 13 1 13 1 13 10 9 2 10 9 7 10 9 2
30 1 9 2 9 3 0 2 13 1 10 9 2 13 9 3 0 2 1 9 1 12 1 12 7 3 1 12 1 12 2
22 1 9 2 10 9 1 11 13 10 9 0 1 10 9 0 2 3 1 10 9 12 2
31 10 2 0 9 2 16 13 10 9 0 1 10 9 1 9 2 4 4 3 13 1 10 9 0 13 1 10 9 11 11 2
9 11 11 13 10 9 0 1 9 2
14 10 9 13 3 10 9 1 11 11 11 11 11 11 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 9 2
28 13 1 10 9 13 10 9 7 13 15 1 10 9 2 10 15 4 13 15 1 9 1 10 9 1 10 9 2
20 10 0 9 1 11 13 1 10 9 1 10 11 0 1 10 9 11 2 11 2
7 13 10 9 7 10 9 2
23 10 9 4 13 1 16 10 9 0 1 9 0 13 13 15 1 10 9 0 16 15 13 2
43 10 9 1 9 1 10 9 0 13 3 0 1 10 9 2 9 1 10 9 2 9 1 9 7 3 3 2 1 10 9 0 2 10 9 3 13 1 10 9 1 10 9 2
10 15 13 10 9 0 7 3 15 0 2
23 13 10 9 1 9 7 9 2 10 9 13 1 13 7 4 13 10 9 1 10 9 0 2
21 4 13 1 5 10 0 9 1 10 9 1 10 9 1 9 1 3 1 10 9 2
14 13 3 10 9 7 3 1 10 9 0 1 10 9 2
44 10 9 1 9 1 11 2 11 11 2 13 3 1 16 10 9 0 1 10 9 13 9 0 1 10 9 1 10 0 9 0 1 10 9 1 10 9 1 10 11 11 7 11 2
20 1 15 9 1 10 9 13 1 12 9 7 13 12 9 7 12 9 1 9 2
24 1 1 10 9 1 10 9 2 11 3 13 9 1 10 9 0 16 13 13 1 11 11 2 2
28 3 13 10 9 13 11 11 2 11 11 11 2 1 10 9 0 1 11 2 13 3 10 9 1 10 9 0 2
25 1 0 9 2 13 1 10 9 11 11 2 11 11 2 7 1 10 9 3 13 0 11 11 11 2
35 10 9 13 1 10 9 10 11 1 10 9 1 11 1 10 9 16 13 2 13 10 9 7 10 9 2 13 1 11 7 1 10 9 2 2
38 10 9 1 9 13 1 9 1 11 7 10 9 0 7 10 9 0 1 10 9 4 13 1 9 1 11 1 10 11 1 11 1 10 9 1 12 9 2
48 1 11 10 9 1 10 9 4 7 13 15 10 9 0 2 1 15 2 13 10 9 1 16 16 13 1 10 9 7 15 9 1 10 9 2 15 15 13 1 10 9 16 13 15 10 9 0 2
15 11 11 11 2 15 13 1 10 9 1 9 16 15 13 2
54 1 10 9 1 10 9 11 2 10 9 1 16 10 9 13 1 10 9 1 10 9 2 10 11 2 1 11 11 2 1 10 9 1 10 9 0 7 10 11 2 15 13 0 13 1 10 9 1 10 9 0 11 11 2
67 10 9 13 10 9 1 10 11 1 11 11 1 10 11 2 1 10 9 3 0 1 10 9 1 11 2 9 1 10 15 13 1 13 10 9 13 3 1 10 9 1 10 9 11 1 10 9 2 16 13 13 13 1 10 9 1 10 9 1 13 15 1 10 11 1 11 2
16 10 9 13 12 9 1 11 2 9 0 2 7 1 12 9 2
45 1 12 2 11 11 2 10 3 9 1 9 0 7 9 0 1 10 9 2 13 10 9 1 11 1 10 11 1 10 11 7 10 9 1 10 9 1 9 7 9 1 9 7 0 2
21 11 11 2 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 1 11 2
13 3 3 7 1 11 2 3 1 12 9 4 13 2
42 3 10 10 9 16 3 13 3 1 10 9 2 7 13 10 9 1 9 7 1 9 2 13 9 1 10 9 2 3 13 1 4 13 7 13 9 1 9 1 10 9 2
14 15 13 3 7 13 13 15 3 7 16 15 13 15 2
15 13 16 1 9 1 9 3 13 15 13 16 13 10 9 2
12 1 12 13 10 9 1 11 11 1 10 11 2
31 13 1 10 12 9 10 9 1 9 1 9 0 0 0 7 10 12 9 1 10 0 9 2 16 13 10 9 1 10 9 2
31 13 10 9 0 1 11 1 11 2 1 15 13 10 9 13 11 11 11 2 16 13 1 10 12 9 1 9 1 10 9 2
44 10 9 0 1 10 11 11 13 0 1 10 15 7 0 1 10 10 9 0 2 16 3 1 10 9 0 7 0 10 9 1 10 9 0 13 2 7 13 3 3 7 3 0 2
61 3 15 13 10 11 1 11 7 11 1 12 2 13 3 9 0 2 7 1 9 2 10 11 1 11 11 1 9 1 9 1 10 11 11 15 13 1 12 1 11 2 13 3 10 9 1 10 9 1 10 9 0 2 9 0 2 0 7 1 9 2
22 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 11 2
25 10 9 1 9 13 0 7 2 16 13 10 15 3 0 7 10 9 1 10 9 2 13 10 9 2
30 3 0 15 13 1 9 1 9 2 10 9 1 10 9 0 2 1 9 0 2 1 10 0 16 10 9 1 10 9 2
28 1 10 9 2 3 11 13 10 9 1 13 9 0 1 10 9 7 10 9 7 13 10 9 1 9 1 12 2
26 1 9 1 10 0 9 2 10 11 11 13 10 9 0 7 0 2 7 0 1 10 9 7 10 9 2
38 10 9 1 9 13 10 9 1 10 9 2 16 15 13 1 13 9 1 9 0 1 10 9 2 1 9 3 1 13 9 1 9 1 13 1 3 0 2
10 11 13 1 10 9 1 10 9 0 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
39 1 10 9 0 2 10 9 13 16 10 9 1 11 3 13 0 1 10 9 2 7 11 13 10 9 1 13 1 10 9 11 13 16 11 13 1 10 9 2
8 1 15 13 9 1 10 9 2
17 13 3 1 10 9 2 11 11 1 10 11 1 13 1 10 11 2
12 1 10 9 1 10 11 3 13 9 1 9 2
31 1 15 2 10 9 13 1 11 13 1 10 9 11 1 13 10 9 1 10 9 13 3 2 7 13 10 9 1 9 9 2
29 3 15 13 1 10 9 1 9 11 7 11 1 10 11 2 7 10 9 0 1 10 9 11 1 10 9 11 11 2
18 13 9 0 1 10 11 1 11 11 7 11 2 11 11 2 1 12 2
25 13 10 9 2 11 2 12 1 11 2 11 11 11 2 11 11 2 11 11 2 11 2 11 11 2
28 1 10 9 2 11 13 2 2 10 10 9 15 13 1 9 1 10 9 1 10 9 7 3 16 3 4 13 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
21 1 13 10 9 13 1 11 11 16 13 9 1 10 9 1 10 9 1 10 9 2
16 15 13 2 11 2 7 2 11 2 7 1 15 2 11 2 2
15 0 9 1 10 9 1 10 9 3 4 13 1 10 9 2
10 13 10 9 1 12 12 9 1 12 2
54 10 9 1 10 9 1 10 9 1 11 4 13 1 10 9 1 10 9 0 8 10 9 0 0 2 7 4 13 10 9 1 9 1 10 9 2 1 16 10 9 1 9 1 11 13 10 9 1 10 9 1 10 11 2
33 10 9 13 0 1 10 9 1 10 9 1 9 1 12 9 2 12 9 2 7 1 10 10 9 1 10 9 0 2 12 9 2 2
7 13 1 10 9 1 9 2
11 13 10 9 0 16 13 10 9 1 9 2
35 10 9 1 11 1 12 13 10 9 13 10 12 1 11 1 10 12 1 10 12 9 9 0 2 12 9 2 16 13 10 9 1 12 8 2
32 1 9 8 13 10 8 2 9 2 2 13 13 2 13 9 1 10 9 2 2 7 1 10 9 0 1 8 13 10 9 8 2
27 3 1 12 2 10 9 11 4 1 13 10 9 13 3 1 10 9 7 13 1 9 1 12 8 12 9 2
28 3 0 2 13 16 2 13 16 1 10 9 10 9 13 0 7 3 15 13 13 1 10 9 1 9 0 2 2
25 3 3 2 1 10 13 10 9 0 15 13 0 16 13 1 10 9 0 7 15 13 1 9 2 2
69 2 16 13 1 10 9 11 11 2 4 13 16 1 12 10 9 13 1 10 9 0 1 12 9 2 7 3 3 15 13 10 9 1 9 2 10 9 7 15 13 10 0 9 0 2 10 9 0 13 10 9 1 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
6 10 9 0 13 0 2
38 3 2 15 13 1 10 9 1 10 9 1 13 10 9 1 10 9 2 3 16 3 4 13 10 9 1 10 9 7 13 10 9 0 1 1 10 9 2
44 10 9 1 9 1 10 12 1 11 1 12 2 13 9 0 1 10 9 0 1 9 1 10 9 9 9 5 12 2 1 10 12 1 11 1 12 2 10 15 13 10 9 0 2
43 3 2 1 10 13 1 11 2 15 13 1 10 9 0 2 15 13 1 10 9 1 11 11 13 10 9 1 10 9 0 1 10 9 1 9 1 11 1 9 1 10 9 2
11 3 13 16 3 15 13 9 1 10 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
23 1 9 1 9 1 10 9 2 10 9 13 3 0 1 13 8 8 15 13 10 9 0 2
17 3 13 16 13 10 10 9 1 11 1 9 0 16 4 13 15 2
33 10 9 3 13 16 10 9 13 1 10 9 10 9 2 15 16 9 10 9 1 9 7 9 15 10 9 1 11 13 1 10 9 2
21 10 9 13 9 1 9 1 10 9 0 0 2 8 2 7 0 0 2 11 2 2
4 11 13 9 2
38 1 9 2 10 0 9 1 10 9 0 11 11 13 1 10 9 1 11 2 15 3 4 13 1 9 1 10 9 11 2 7 1 10 9 1 10 9 2
50 1 10 0 9 1 10 11 11 7 10 0 9 1 9 1 10 15 11 11 2 10 9 1 13 9 13 10 0 11 2 10 9 16 13 13 1 9 1 13 15 1 11 7 10 10 9 1 13 11 2
7 10 9 15 13 15 0 2
35 1 12 1 12 13 9 1 10 2 11 11 1 11 2 2 7 1 12 1 12 13 9 1 10 9 1 9 2 9 0 7 9 1 9 2
19 13 9 1 11 11 2 9 2 9 1 11 2 15 13 0 1 11 11 2
37 16 10 0 9 1 10 11 11 1 11 13 10 9 0 0 2 1 11 1 12 2 11 4 13 9 1 10 9 1 9 2 13 1 13 10 9 2
25 1 12 10 9 15 13 1 0 9 2 1 10 9 1 10 11 11 11 11 11 16 13 10 9 2
10 15 4 13 1 11 11 12 1 9 2
12 11 11 13 10 9 0 13 7 13 1 11 2
20 10 9 1 10 9 15 13 1 10 9 1 3 15 13 10 9 7 15 13 2
35 1 13 10 9 13 1 11 13 3 13 10 9 0 0 2 1 10 9 1 11 1 9 1 10 9 0 7 11 1 9 1 10 9 0 2
9 9 0 7 0 13 1 9 0 2
40 10 9 0 3 13 9 1 10 9 1 9 1 13 15 1 10 9 3 0 1 9 1 3 13 10 9 7 1 10 9 13 10 0 9 1 10 9 3 0 2
19 13 0 1 10 9 1 10 11 2 12 2 16 13 1 10 9 1 11 2
33 10 9 0 7 0 13 10 0 9 1 9 1 10 9 1 10 11 0 1 10 9 1 9 1 10 9 0 1 10 11 11 11 2
20 13 1 12 1 11 16 13 1 10 9 1 11 2 4 13 1 10 9 0 2
20 1 12 13 1 11 16 13 1 10 9 16 15 13 13 10 9 2 10 11 2
24 1 10 9 0 13 10 0 9 1 11 2 15 16 13 10 9 1 10 10 9 1 10 9 2
27 10 9 4 13 10 9 1 10 9 7 15 4 13 0 9 1 13 15 1 10 9 7 9 1 10 9 2
38 3 4 13 9 1 10 9 1 13 10 9 0 1 10 0 9 2 15 15 13 1 10 9 1 10 9 0 1 13 7 13 1 10 9 16 13 0 2
17 11 13 10 9 1 9 1 9 1 12 9 0 1 10 9 11 2
12 11 11 13 10 9 1 9 1 10 9 11 2
21 11 13 10 9 0 0 1 9 7 9 0 2 13 1 12 1 11 11 2 11 2
41 3 0 13 11 11 1 10 9 7 4 7 13 12 9 1 16 13 16 10 9 0 4 13 2 10 9 1 10 9 7 10 9 2 16 13 10 9 0 11 11 2
12 13 3 16 10 9 1 9 13 1 10 9 2
75 4 13 16 11 2 3 15 4 13 10 9 1 13 2 10 9 7 4 13 1 16 15 13 1 9 1 13 10 9 7 13 15 1 15 16 13 1 11 11 7 1 15 16 15 13 1 10 9 2 1 9 1 9 13 1 9 7 16 15 4 1 13 2 1 9 0 7 3 13 9 0 7 0 2 2
44 10 9 1 9 13 1 10 0 9 2 16 16 15 4 13 1 9 1 10 9 12 2 3 15 15 3 2 2 4 13 1 10 0 12 9 16 4 4 1 13 3 1 9 2
19 4 4 13 10 9 1 9 0 1 9 0 1 9 7 9 1 10 15 2
18 7 13 10 0 9 1 10 9 0 1 11 11 16 13 10 9 13 2
33 10 12 1 11 2 13 1 10 9 1 11 1 11 2 10 9 7 12 9 3 1 9 2 13 10 9 1 10 9 16 15 13 2
18 11 13 10 9 0 1 10 9 1 11 2 13 1 10 9 1 11 2
79 16 10 9 13 1 10 9 2 7 10 9 13 1 11 2 15 1 10 9 2 2 16 15 13 16 10 9 1 11 0 9 3 13 10 9 1 11 2 16 3 10 9 1 13 10 15 1 10 15 2 16 1 15 10 9 13 1 9 2 7 15 13 16 13 10 0 9 1 13 0 2 1 15 15 13 13 1 15 2
106 1 10 9 2 11 8 11 2 2 11 4 7 13 1 11 1 10 11 11 11 2 7 2 16 11 13 13 1 10 9 7 15 13 1 13 15 1 9 1 11 11 2 10 11 1 11 3 15 13 1 9 7 15 13 2 3 13 16 11 15 13 1 11 2 2 15 13 10 9 4 7 4 1 13 1 10 11 2 3 16 1 15 0 15 4 13 7 3 13 1 16 11 13 3 1 4 13 10 9 16 4 13 1 10 9 2
23 10 10 9 0 0 1 10 9 4 13 1 11 2 3 2 11 2 2 13 1 11 11 2
16 10 0 9 0 2 10 11 11 10 11 2 13 0 1 9 2
44 10 9 1 11 11 3 13 1 9 0 7 9 0 13 10 9 13 1 10 9 16 13 1 10 11 11 7 1 10 11 11 2 3 11 11 2 2 9 1 11 2 11 2 2
19 10 9 13 16 3 13 10 9 13 11 2 15 1 10 9 0 1 11 2
53 1 10 0 9 1 10 9 1 10 8 2 10 9 13 1 0 0 2 16 16 13 9 1 9 2 13 3 9 2 1 10 13 10 9 1 9 1 10 9 8 1 10 11 1 10 11 1 10 9 1 10 9 2
44 12 9 0 2 10 9 13 1 12 7 12 2 4 4 13 1 12 9 0 1 9 0 2 11 1 11 7 11 1 10 9 1 10 11 2 11 1 10 9 1 10 11 11 2
25 1 9 1 13 0 2 15 3 13 1 13 10 9 1 9 7 10 9 1 10 9 1 0 9 2
44 13 10 9 0 7 1 10 9 1 10 12 9 13 10 16 3 15 13 2 1 10 9 1 11 7 11 15 13 10 9 3 7 4 13 10 9 1 9 8 1 10 0 8 2
30 10 11 4 13 1 9 1 10 9 0 10 9 1 11 11 16 4 13 16 13 10 9 0 1 10 9 2 11 2 2
20 10 10 9 13 1 11 11 2 11 11 7 8 11 3 16 15 13 15 9 2
44 10 9 2 16 15 13 1 10 12 1 10 12 5 1 10 11 1 10 11 2 15 13 1 13 10 0 9 1 9 2 16 13 9 1 10 9 3 0 1 10 9 1 11 2
48 1 12 15 13 16 3 1 10 9 1 10 9 16 13 10 9 2 13 10 0 9 1 10 9 2 8 2 1 10 9 12 2 7 15 13 3 10 9 1 10 9 7 10 1 11 2 11 2
37 1 10 9 2 11 11 2 15 1 10 12 9 7 10 9 1 10 9 1 11 1 10 9 1 11 2 13 10 0 9 13 1 10 9 1 11 2
12 15 13 1 7 10 9 15 13 13 1 9 2
21 13 1 13 15 16 3 13 10 11 11 1 10 11 11 1 11 7 10 11 11 2
27 15 9 10 9 16 13 1 9 2 3 0 1 9 7 1 0 9 2 9 16 15 13 1 10 9 2 2
25 10 9 1 11 13 10 9 1 10 0 9 1 9 0 1 10 9 1 11 2 11 11 2 11 2
21 13 3 1 10 9 16 3 13 3 3 1 9 1 10 9 2 1 0 2 0 2
15 10 9 3 13 7 13 1 10 9 1 10 9 2 9 2
25 10 9 13 9 0 2 13 1 9 0 1 10 9 7 10 9 1 10 9 3 1 10 9 0 2
18 10 9 15 13 10 9 4 13 1 10 9 15 13 11 11 1 12 2
6 15 13 9 1 9 2
6 13 1 11 2 11 2
12 11 11 13 10 9 1 9 1 10 9 11 2
27 11 13 1 12 1 11 11 1 10 9 1 11 0 7 11 11 2 7 1 12 4 13 1 10 11 11 2
14 10 9 3 13 1 9 2 13 2 8 8 8 8 2
12 15 13 1 10 9 0 1 10 9 1 9 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
64 16 13 10 9 1 9 2 1 10 9 1 9 7 10 9 2 7 13 1 10 9 10 9 7 1 10 10 9 2 7 13 1 10 9 1 10 9 16 13 10 0 9 1 9 2 13 10 9 9 1 10 9 1 10 9 7 10 9 16 13 10 0 9 2
38 1 10 9 1 8 2 9 1 10 9 1 10 9 11 2 10 11 13 10 9 1 10 9 1 10 9 11 7 10 9 0 1 9 2 11 2 0 2
15 10 9 1 9 13 1 3 1 12 12 9 0 1 12 2
45 1 15 15 3 15 13 7 1 9 1 10 9 1 10 0 9 2 10 9 0 1 11 15 13 10 0 9 1 9 1 12 2 10 9 1 12 7 10 0 9 1 10 9 0 2
11 10 9 1 11 15 13 13 1 10 9 2
12 10 9 13 8 0 7 10 9 0 1 9 2
13 13 9 3 1 15 13 10 9 16 15 13 3 2
23 13 1 10 9 9 0 11 11 2 11 11 2 1 10 9 1 10 9 7 9 3 0 2
24 10 9 1 10 9 0 1 11 13 1 10 9 0 1 10 9 1 9 1 10 9 1 12 2
35 1 16 13 1 16 15 13 4 3 3 13 1 10 9 1 10 9 2 13 15 10 9 3 0 13 15 10 9 16 15 13 1 10 9 2
21 13 13 10 9 2 16 1 9 15 13 9 0 16 13 10 0 9 1 10 9 2
9 1 9 13 15 16 3 9 13 2
39 13 10 0 9 1 10 9 1 10 9 0 13 10 11 1 11 2 9 1 12 1 11 1 12 2 2 10 11 11 1 12 2 10 11 2 1 10 9 2
23 16 10 9 16 13 13 3 2 9 0 2 10 9 13 0 7 10 9 13 3 7 13 2
23 10 0 9 13 13 1 10 9 1 9 1 9 1 9 0 1 10 12 9 1 10 9 2
39 10 9 11 13 10 9 1 9 1 10 9 1 11 11 13 1 10 9 1 10 11 11 7 10 9 1 10 11 11 2 13 1 10 9 1 11 2 11 2
39 1 10 9 1 10 9 12 11 2 12 7 12 11 2 10 9 12 2 10 9 9 12 7 10 9 12 2 12 11 2 12 7 12 2 13 1 12 9 2
38 4 13 16 10 0 9 13 1 13 9 7 13 10 9 1 16 12 9 0 2 13 1 9 0 2 1 13 1 0 9 1 9 2 4 13 1 9 2
12 13 12 9 13 10 9 7 13 10 0 9 2
47 10 9 1 10 12 1 11 1 11 1 10 11 11 4 4 13 1 12 1 11 11 2 11 11 1 10 9 11 11 2 11 2 7 1 12 13 1 11 10 9 1 9 0 1 10 9 2
41 13 1 10 0 9 1 9 7 9 15 13 10 9 2 10 9 1 10 9 7 1 10 0 9 1 10 9 15 4 13 1 10 0 9 2 11 7 9 1 11 2
21 10 9 7 10 9 4 13 1 10 9 1 10 9 7 13 1 9 11 2 11 2
43 1 10 9 1 10 9 1 10 11 11 2 11 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 4 1 9 0 7 2 12 5 2 12 9 5 13 9 2
17 7 16 10 9 0 13 10 9 0 2 10 0 9 13 3 0 2
42 1 13 10 9 15 13 1 11 11 2 15 1 10 4 13 10 9 1 10 9 11 1 15 16 13 9 1 10 9 1 10 9 2 11 11 2 2 15 13 1 9 2
14 11 13 1 10 9 7 13 1 9 3 13 1 9 2
38 15 13 1 10 9 16 13 12 9 1 9 1 11 12 1 10 9 7 9 11 11 13 1 10 9 1 11 1 10 9 1 9 1 10 11 1 11 2
25 1 10 9 10 9 1 10 9 2 11 2 11 1 10 11 7 11 11 11 13 16 13 12 9 2
38 13 10 9 0 2 10 9 1 9 13 1 10 9 10 9 3 3 2 8 2 1 10 9 2 13 16 16 10 9 4 13 2 10 9 3 15 9 2
14 10 9 1 9 7 9 15 13 3 0 1 9 0 2
21 4 13 1 12 7 1 3 4 13 13 10 9 16 13 1 12 9 1 12 9 2
32 0 1 10 9 1 10 9 1 11 11 2 10 9 11 13 10 12 9 1 10 9 3 0 1 11 1 13 1 10 9 0 2
23 10 9 1 10 9 1 9 1 11 1 10 9 3 0 1 11 1 13 11 11 10 11 2
22 1 9 2 13 1 11 3 13 1 13 10 9 0 2 10 9 0 2 15 13 11 2
15 10 9 2 16 3 13 9 2 3 4 13 15 1 15 2
39 3 10 9 15 4 13 1 10 9 1 11 11 7 11 11 2 15 4 13 10 9 7 10 3 1 10 9 1 10 2 9 1 10 9 2 2 9 2 2
29 13 10 9 11 12 10 11 2 15 13 10 9 0 1 9 0 7 10 9 16 13 3 10 0 9 1 10 9 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
18 10 11 11 2 11 2 11 11 2 13 10 0 9 1 10 9 11 2
24 15 1 15 3 15 13 0 1 10 9 1 11 11 2 9 0 16 13 9 1 10 9 11 2
40 10 9 2 13 1 9 7 13 1 12 9 2 4 13 10 9 0 1 10 9 1 11 10 12 1 11 2 1 9 1 10 9 1 10 9 11 12 1 11 2
36 3 1 10 9 2 10 9 13 10 9 1 9 0 2 1 10 15 11 11 13 1 10 9 3 0 1 10 9 1 10 9 1 12 7 12 2
30 1 10 11 1 10 11 1 12 10 9 0 1 9 1 10 9 13 1 5 12 7 10 9 0 1 9 13 5 12 2
22 16 15 4 1 13 2 13 7 10 9 1 11 13 1 10 1 10 9 13 1 11 2
28 3 2 1 11 1 12 10 9 13 1 11 10 9 2 13 15 1 10 9 0 7 13 1 15 9 1 9 2
28 12 9 0 2 10 9 8 13 10 9 11 10 11 2 13 1 11 1 11 11 2 1 10 9 0 11 11 2
20 13 1 10 11 11 11 7 13 1 10 9 1 11 12 7 11 12 1 11 2
32 15 13 15 10 9 0 16 15 13 11 1 10 9 7 15 13 2 3 2 1 7 10 9 15 13 1 10 9 1 10 9 2
86 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 15 13 0 10 8 8 13 10 9 7 9 0 16 13 10 9 1 10 9 1 11 2 0 1 13 10 0 0 9 1 9 1 15 9 1 10 11 1 11 2 11 11 2 2 13 1 15 13 10 9 0 7 3 4 13 1 9 1 9 1 10 9 0 2 1 10 9 1 10 9 2
30 10 9 13 1 10 9 1 11 2 1 10 1 11 2 1 10 11 1 11 2 2 16 13 9 1 10 9 1 11 2
29 10 9 1 10 11 13 10 9 0 16 15 13 3 1 10 11 1 10 11 1 11 2 1 10 9 0 1 11 2
53 11 11 1 11 13 16 13 10 9 1 10 15 13 0 1 4 15 13 2 13 16 13 10 9 1 9 16 15 13 3 1 10 9 7 10 9 1 11 11 2 7 15 1 9 15 13 1 10 9 1 10 9 2
46 13 3 2 7 3 1 13 10 11 2 15 13 1 10 9 2 13 10 9 2 11 11 1 10 11 2 11 2 11 11 1 10 11 2 11 2 10 11 1 10 11 2 7 3 11 2
31 3 13 1 11 11 11 1 10 11 11 11 2 7 13 1 13 10 9 1 10 9 2 13 12 1 12 9 7 12 9 2
26 10 10 9 1 10 9 13 3 0 7 10 9 13 15 9 1 10 11 11 11 1 1 10 9 0 2
43 3 2 2 10 11 11 11 2 13 10 9 11 1 4 13 10 9 1 0 9 0 2 7 16 10 9 0 13 10 9 1 0 9 1 10 12 1 10 9 11 11 11 2
30 15 13 9 1 10 11 11 1 10 11 7 10 11 1 12 7 9 1 10 11 11 1 10 9 7 10 11 1 12 2
18 10 9 13 10 9 0 1 9 12 9 1 10 9 12 1 10 9 2
7 13 8 4 1 13 9 2
22 10 9 13 10 9 1 10 9 0 2 13 10 9 1 13 10 0 9 1 10 11 2
40 15 3 13 10 9 0 1 10 0 9 1 9 16 13 9 0 2 13 16 15 3 13 10 0 9 1 9 1 9 2 7 16 13 9 0 0 1 9 0 2
22 10 9 1 10 9 3 15 13 0 2 15 16 13 16 10 9 15 13 1 10 9 2
8 11 13 10 9 1 11 11 2
33 11 11 2 2 11 2 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 15 1 10 9 0 1 9 3 0 1 11 2
37 1 10 9 1 11 12 1 11 2 13 1 13 1 11 11 2 7 13 13 16 15 13 1 11 1 10 9 1 12 2 7 10 9 13 1 9 2
17 13 1 15 2 1 10 9 12 10 9 13 10 9 1 10 9 2
31 10 9 13 10 9 0 1 10 9 0 2 3 7 13 9 1 9 0 2 1 10 9 1 10 9 1 10 9 1 9 2
47 11 11 11 2 13 1 11 7 11 1 11 11 2 11 2 13 10 9 0 1 11 11 16 15 13 10 12 1 11 1 12 1 11 11 2 1 10 9 1 12 9 1 9 1 10 9 2
52 1 9 1 10 9 0 15 4 13 10 0 9 1 10 9 0 1 10 9 2 15 15 13 0 1 10 9 11 11 2 1 10 15 15 13 0 9 1 9 0 2 9 3 7 3 1 10 9 2 9 2 8
38 11 13 3 1 10 9 2 0 1 15 1 10 10 9 1 11 11 2 10 0 9 1 9 2 3 10 0 9 1 10 9 16 13 1 10 10 9 2
48 10 9 13 1 13 10 12 11 1 11 11 1 10 11 11 2 11 11 11 2 13 10 9 1 9 7 9 2 0 1 10 9 11 11 2 1 10 9 2 11 2 2 1 11 2 11 2 2
32 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2 13 15 1 10 9 3 0 1 10 9 2
23 4 7 13 10 9 0 2 3 0 1 10 9 2 7 10 9 7 9 1 10 9 0 2
19 15 13 1 11 2 9 0 1 10 9 1 10 9 11 1 11 7 11 2
26 10 9 1 15 13 16 10 9 1 9 4 13 10 3 0 9 1 9 0 1 10 9 7 10 9 2
7 3 15 13 11 1 11 2
48 1 15 9 1 10 11 2 15 13 1 10 9 1 10 9 1 10 11 1 11 7 10 9 1 11 1 10 11 2 1 10 9 1 13 10 9 0 1 10 9 0 1 10 15 1 10 9 2
62 10 9 2 11 11 2 4 13 1 10 9 1 11 11 1 10 3 0 1 4 13 2 1 9 2 8 2 4 10 9 13 1 11 11 2 2 3 16 13 16 13 7 2 1 0 2 13 1 10 9 1 10 9 2 15 16 13 3 1 10 9 2
14 10 9 1 10 9 3 13 0 1 10 9 1 12 2
27 11 11 11 2 11 2 12 2 2 11 11 2 11 2 11 2 12 2 7 11 2 11 11 2 12 2 2
9 13 1 10 9 11 11 1 11 2
22 13 10 9 1 11 0 1 10 9 1 10 9 7 15 15 15 13 10 12 1 11 2
52 10 9 0 13 1 10 9 1 10 9 1 11 7 11 2 1 10 9 1 11 7 11 2 1 10 9 1 10 11 2 11 2 10 11 7 11 11 2 9 1 11 2 7 1 10 9 1 10 9 1 11 2
16 1 0 4 13 1 9 7 4 13 1 9 7 1 10 9 2
11 10 9 11 12 4 13 1 11 1 12 2
143 11 2 15 15 4 13 1 10 9 7 9 1 10 9 0 1 10 9 1 11 11 1 11 11 2 13 10 9 1 11 1 11 1 10 9 1 15 13 10 9 1 10 15 10 9 0 13 10 9 1 9 7 10 9 0 7 1 10 9 15 13 1 0 9 10 9 0 2 13 13 16 13 1 10 10 9 2 11 13 1 15 9 1 10 9 1 10 9 1 9 1 9 0 16 15 13 1 12 2 10 9 1 10 9 15 13 1 10 9 12 1 15 15 13 1 10 9 0 2 10 15 4 13 1 10 0 9 1 10 11 2 11 11 11 2 13 10 9 1 11 1 12 2
23 10 9 15 13 1 10 9 1 10 9 1 10 9 13 1 10 9 1 10 0 9 0 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
64 13 0 16 10 0 9 1 1 11 2 11 7 0 9 2 13 1 10 9 1 11 11 3 13 3 7 13 15 9 1 10 9 2 7 10 11 4 13 13 10 9 0 1 10 9 1 13 1 10 9 0 7 0 13 16 1 10 9 9 13 1 10 9 2
43 10 9 13 12 9 1 9 1 9 1 9 0 13 1 9 0 3 15 13 2 1 9 0 2 10 9 2 9 1 11 11 2 11 11 0 7 11 11 13 1 11 12 2
17 10 9 13 10 9 0 2 13 1 13 10 9 7 10 9 13 2
23 1 12 1 11 1 10 12 1 11 10 9 13 1 11 11 7 1 9 1 9 1 11 2
15 10 9 0 4 13 15 3 1 15 9 7 9 1 11 2
32 11 13 10 9 2 15 15 15 13 13 1 9 16 10 9 0 3 13 3 15 3 0 1 9 1 10 9 1 10 9 0 2
10 10 9 3 13 1 12 9 1 9 2
7 10 9 0 3 13 15 2
26 1 10 9 13 11 11 1 9 2 11 11 1 9 7 11 11 2 9 1 11 2 13 10 9 3 2
35 1 13 10 9 1 11 11 4 7 13 16 10 9 1 10 9 13 1 10 9 1 11 2 1 10 11 2 1 10 11 7 1 10 11 2
41 1 13 1 12 2 7 16 11 15 13 1 9 0 2 10 0 9 15 13 1 9 1 10 9 1 10 11 1 10 11 0 7 10 11 11 1 10 11 1 11 2
20 7 3 10 0 9 15 11 13 1 10 9 13 13 1 10 9 0 1 11 2
37 10 9 7 10 9 1 9 1 10 10 9 0 2 16 13 3 1 12 9 1 0 9 2 15 13 1 10 9 1 9 0 7 0 13 1 11 2
19 10 9 0 13 1 12 9 5 7 13 10 9 1 12 8 5 9 5 2
20 15 13 10 9 1 9 1 10 9 16 13 15 7 13 1 10 9 16 13 2
52 3 3 7 10 9 0 13 13 15 1 10 9 1 10 9 0 2 4 13 10 9 1 3 15 13 10 11 7 10 12 9 13 1 10 9 0 0 1 4 13 9 1 0 9 1 10 9 1 9 1 11 2
23 10 9 1 9 1 10 9 13 16 4 13 10 9 0 2 15 1 15 15 3 13 0 2
42 1 9 2 10 9 1 10 9 15 13 0 1 10 9 0 7 2 1 15 9 2 1 10 9 1 10 9 0 7 0 2 1 10 15 13 3 3 11 7 11 11 2
38 10 9 1 11 11 4 13 10 9 1 10 11 1 11 7 15 13 3 2 1 13 9 0 1 10 9 0 16 13 1 10 9 3 12 9 1 9 2
16 7 13 10 9 1 9 16 1 9 13 9 1 9 7 9 2
11 10 9 1 11 15 13 13 1 10 9 2
60 11 13 10 9 1 10 0 11 11 0 2 1 10 9 16 13 1 10 9 2 1 10 9 1 9 1 10 9 2 1 10 9 1 13 1 10 0 9 2 1 10 9 1 4 13 7 1 10 9 1 13 15 1 10 0 9 1 10 9 2
79 10 9 0 13 0 2 1 9 3 7 3 0 2 1 10 10 9 2 13 10 9 0 7 13 1 10 9 9 1 9 2 9 0 1 10 9 12 7 10 0 9 1 10 9 12 2 7 16 13 1 9 1 10 0 9 1 10 9 12 1 3 13 15 1 0 1 3 10 10 9 2 1 1 10 9 1 9 0 2
38 1 10 11 11 11 10 11 0 16 4 13 1 9 1 11 4 1 13 10 11 11 1 11 2 15 1 10 9 0 1 11 2 15 3 0 1 15 2
14 11 13 4 13 12 9 1 13 1 10 9 1 11 2
30 10 9 0 2 1 11 1 10 9 7 1 11 11 1 9 2 11 3 13 1 10 9 7 3 13 12 9 1 11 2
15 3 2 11 11 7 11 11 3 13 13 10 9 1 9 2
39 3 1 16 10 9 4 1 13 1 11 1 12 1 10 9 8 2 12 2 7 8 2 12 2 2 10 9 4 13 1 15 10 9 1 9 1 0 9 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
10 11 11 4 13 1 2 11 2 11 2
58 10 9 0 3 3 13 10 9 1 11 11 7 10 9 16 2 1 11 2 15 13 1 15 16 13 1 13 10 0 9 16 13 10 9 0 2 10 9 16 2 16 13 10 9 2 4 4 13 15 0 1 10 9 1 10 11 2 2
62 10 9 13 10 9 1 13 7 13 10 9 1 0 9 1 10 9 1 13 15 1 10 9 1 10 9 1 9 1 9 0 1 13 1 10 9 16 13 9 1 9 2 10 9 1 9 1 9 7 9 1 10 9 1 9 1 9 2 1 10 9 2
28 13 3 1 10 9 10 9 1 9 1 12 9 2 11 2 11 2 11 11 11 7 11 11 11 2 11 11 2
21 1 3 1 9 1 12 9 2 13 3 3 10 11 2 11 11 7 11 11 11 2
25 1 10 9 13 11 2 13 11 2 7 1 10 13 10 9 0 3 4 13 1 13 11 7 11 2
7 10 9 3 13 12 9 2
14 1 10 8 13 13 11 2 12 7 3 15 13 3 2
8 10 9 4 13 1 11 11 2
21 10 0 9 1 10 9 12 13 0 1 10 9 2 16 3 13 7 10 12 9 2
54 12 9 1 9 16 13 12 9 13 10 11 1 12 0 9 1 10 9 0 2 16 4 13 10 9 1 10 9 7 10 9 1 10 11 0 2 8 2 2 16 4 13 16 4 13 9 7 13 1 3 1 9 0 2
24 3 13 1 11 11 2 10 9 1 10 9 2 13 1 10 9 1 11 16 13 3 10 9 2
22 9 4 13 1 13 9 1 10 11 1 12 7 13 0 1 13 5 12 1 10 9 2
57 1 0 9 2 4 13 1 9 1 0 9 0 2 1 10 15 15 15 4 13 1 13 1 10 0 9 0 1 10 9 1 9 3 0 1 10 9 11 11 11 7 10 9 11 11 2 16 13 0 9 1 10 9 7 9 0 2
30 0 1 10 9 1 11 11 2 10 11 13 10 9 0 1 10 9 2 11 11 2 13 11 8 1 9 1 10 9 2
46 1 10 9 1 10 9 16 15 15 13 1 10 9 0 2 11 13 16 15 13 16 10 9 13 0 1 7 2 10 9 13 9 2 2 15 16 13 1 2 1 9 2 1 10 9 2
17 13 12 9 1 13 10 9 2 7 16 15 13 13 9 13 15 2
23 1 9 13 10 9 13 1 13 10 9 0 7 13 10 9 7 9 0 1 10 9 0 2
28 3 13 9 15 1 9 15 13 10 9 1 10 9 1 9 2 15 16 13 0 13 16 15 13 10 0 9 2
9 13 9 1 13 15 1 10 9 2
21 3 1 13 10 9 7 9 13 13 10 9 1 11 7 3 15 4 13 1 0 2
9 13 10 0 9 0 3 1 9 2
35 1 10 9 2 10 0 7 0 9 1 10 9 1 10 9 0 1 10 9 13 9 0 2 16 13 3 0 7 10 9 0 16 15 13 2
21 11 11 11 13 10 9 13 1 10 9 1 11 7 11 1 10 9 1 11 11 2
28 10 0 10 9 0 1 10 9 13 1 11 11 2 12 2 1 11 11 10 9 1 11 7 3 9 1 11 2
22 1 12 1 11 1 12 10 9 1 10 9 13 1 12 9 2 12 9 7 12 9 2
28 15 15 13 10 0 9 1 13 1 11 2 10 9 13 13 10 0 9 2 15 15 1 10 9 11 3 13 2
30 7 1 10 9 1 3 15 4 13 16 10 9 1 10 9 13 1 10 9 10 0 9 2 3 15 13 1 11 11 2
10 16 4 13 3 0 16 4 13 3 2
22 11 11 13 10 9 1 9 13 1 10 9 0 11 2 16 13 1 10 9 0 11 2
14 10 9 0 13 10 9 0 13 1 11 11 1 12 2
42 3 2 16 3 15 4 13 2 10 11 13 10 9 13 1 11 1 10 9 1 12 2 15 16 15 13 4 1 13 1 10 9 2 7 13 1 10 9 2 1 12 2
12 13 1 10 9 1 13 15 2 13 15 9 2
14 10 9 1 11 7 10 9 4 13 1 11 1 11 2
41 13 1 10 11 11 11 11 2 0 9 1 10 9 2 15 13 10 11 11 7 1 3 1 10 9 1 11 11 11 3 13 10 9 1 10 9 0 1 10 9 2
29 1 10 9 7 1 10 15 1 10 9 16 15 13 3 2 15 15 13 10 9 1 11 2 11 7 2 11 2 2
34 11 11 2 9 1 10 9 1 11 2 11 11 2 10 9 1 11 11 2 7 11 11 2 15 4 13 1 10 9 10 11 1 11 2
12 15 16 13 10 9 1 10 9 13 10 9 2
56 10 9 13 10 9 0 1 10 12 9 1 9 7 1 11 2 11 7 11 1 11 2 9 16 2 1 13 9 2 13 1 10 9 0 1 10 12 9 2 3 7 11 7 11 1 11 1 13 10 9 1 10 0 9 0 2
21 11 2 12 2 2 11 2 11 2 11 2 11 7 11 15 13 10 9 1 9 2
36 10 11 1 11 13 3 16 13 10 9 1 10 9 15 1 10 9 0 2 13 13 2 10 9 16 13 1 10 9 0 7 10 9 1 11 2
27 10 9 1 11 2 11 8 11 1 9 2 13 10 9 1 12 9 3 0 13 1 10 9 0 11 11 2
17 16 11 13 10 9 1 11 2 15 13 15 9 1 13 10 9 2
41 13 10 9 13 1 3 10 9 0 11 11 11 15 15 4 13 1 10 9 1 10 9 3 7 16 13 3 7 15 1 10 9 1 9 1 10 11 1 10 11 2
23 1 9 2 2 11 2 2 2 11 2 13 1 10 9 2 8 2 7 3 12 1 9 2
27 10 9 13 11 1 10 9 0 16 13 1 10 9 2 1 10 9 2 10 9 1 10 9 7 10 9 2
20 1 9 2 10 9 13 16 10 9 3 13 10 0 9 1 10 9 1 11 2
14 10 9 0 3 0 13 10 9 12 5 1 10 12 2
29 10 12 1 11 2 11 13 10 9 1 10 9 0 1 10 9 11 1 11 16 13 10 8 9 12 1 10 9 2
21 13 1 15 2 10 9 13 15 3 0 7 15 3 0 7 15 1 10 9 0 2
41 15 13 1 10 11 11 12 2 16 13 1 10 9 0 1 10 9 1 10 0 9 1 13 10 9 7 13 10 9 0 9 13 1 10 9 1 9 1 9 0 2
5 13 0 1 11 2
17 1 11 1 12 2 13 10 9 1 10 11 2 10 0 9 0 2
85 2 15 2 13 11 2 13 10 9 7 10 9 1 10 0 12 9 2 13 16 3 3 13 0 13 10 9 2 16 3 2 7 7 13 0 13 3 10 9 1 9 2 3 15 13 13 1 10 9 2 13 10 9 1 10 9 2 10 9 16 13 10 9 7 13 15 1 9 1 10 9 16 15 13 2 16 15 13 7 16 15 13 9 2 2
16 13 3 10 9 0 10 11 7 11 1 11 2 1 11 2 2
33 1 9 1 10 9 12 10 9 10 11 2 1 11 11 11 2 15 13 3 11 1 11 1 10 9 0 0 1 10 11 1 11 2
30 1 10 9 0 1 10 9 15 13 10 9 2 11 2 7 1 10 9 0 2 0 1 10 9 2 10 9 8 7 8
29 1 10 8 2 9 10 9 15 13 13 1 10 9 12 7 12 1 9 8 2 1 10 9 0 7 15 0 2 2
17 13 0 15 15 13 10 9 1 9 0 1 10 1 9 7 9 2
20 11 11 13 10 9 1 9 1 10 9 1 10 11 1 10 9 1 10 11 2
15 1 9 2 13 10 9 1 11 2 3 13 9 7 11 2
48 10 9 13 1 10 9 2 7 1 15 15 3 1 9 2 13 1 11 1 10 9 1 11 7 11 2 13 1 0 1 9 1 9 2 9 7 9 1 9 15 3 4 13 1 10 11 0 2
35 1 10 9 1 12 2 11 11 11 11 13 12 12 9 2 12 5 9 2 12 5 9 2 7 10 9 1 9 1 12 9 2 9 5 2
43 16 10 9 3 13 1 10 9 0 1 10 11 11 2 11 13 13 15 1 9 1 10 9 1 10 11 7 13 10 9 0 1 10 9 7 13 1 10 9 1 9 0 2
13 10 9 1 9 13 1 12 8 2 5 9 5 2
5 10 9 13 11 2
38 1 15 9 1 10 0 9 2 11 7 11 15 13 1 9 1 10 9 16 3 13 15 1 10 9 2 10 9 13 16 10 9 13 1 9 1 9 2
39 3 13 10 9 0 1 10 9 1 11 1 10 11 1 11 11 2 3 3 13 10 9 1 10 9 0 2 11 11 2 2 1 10 9 1 10 0 9 2
23 16 4 4 13 1 11 2 10 9 13 10 9 15 0 16 15 4 13 13 10 9 0 2
16 11 11 13 10 9 1 9 1 10 9 11 1 10 9 11 2
15 10 0 9 1 9 15 13 13 1 10 9 10 9 0 2
35 10 9 1 2 11 11 2 2 13 15 3 1 10 9 2 13 1 10 9 1 11 2 3 7 2 11 11 11 12 2 15 13 1 11 2
66 11 11 2 3 0 1 9 1 10 9 2 15 13 12 9 1 12 9 3 1 10 9 2 2 13 10 0 9 1 10 9 1 10 9 2 1 10 15 13 10 9 7 11 2 1 9 1 10 0 9 0 1 10 9 1 9 1 10 9 1 10 9 1 10 9 2
19 1 0 7 10 9 0 2 9 1 3 1 10 0 9 1 10 11 11 2
16 13 10 9 1 13 9 2 15 11 15 4 13 1 12 9 2
42 3 0 2 13 10 9 1 10 9 0 1 10 9 1 10 9 2 3 4 1 13 10 9 7 3 13 1 9 0 1 13 15 16 10 9 11 3 7 13 10 9 2
15 1 9 2 11 2 10 9 1 11 2 13 13 1 9 2
34 10 9 13 1 10 9 11 11 13 1 10 9 1 10 9 0 0 7 9 1 10 9 0 1 10 11 11 11 7 10 11 11 11 2
27 1 9 1 10 9 12 10 11 11 4 13 10 12 9 1 9 1 10 9 0 16 15 13 1 10 9 2
28 1 10 11 1 11 2 10 9 0 13 12 2 16 10 9 13 1 0 2 13 15 1 10 9 12 9 0 2
12 11 13 10 9 0 1 11 1 10 11 11 2
34 4 13 10 9 1 13 10 9 1 15 7 4 13 0 2 13 3 0 7 10 9 1 10 9 13 3 1 3 1 10 9 16 13 2
42 10 9 0 2 13 1 9 1 10 11 11 1 3 1 12 12 9 1 9 2 13 3 2 9 1 9 0 1 9 1 10 9 1 10 9 2 4 4 13 7 13 2
31 10 9 13 13 2 1 9 1 10 9 1 10 9 2 16 10 9 13 13 7 13 15 2 13 1 9 15 13 10 9 2
61 10 9 1 10 9 13 10 9 1 10 11 1 10 15 15 13 10 9 2 13 1 10 9 12 7 10 9 12 13 1 10 9 1 11 12 2 10 11 11 11 11 1 10 11 2 13 1 10 9 12 7 10 9 12 7 10 11 1 10 11 2
18 13 10 12 5 1 9 1 10 9 7 3 10 12 5 1 10 9 2
31 13 12 9 3 1 13 15 2 13 10 9 1 10 9 2 7 2 1 10 9 2 1 10 9 1 9 13 3 12 9 2
8 3 2 13 9 1 11 11 2
8 10 9 1 10 16 13 0 2
36 10 12 1 11 1 12 11 11 13 10 9 1 9 1 9 1 10 9 0 0 1 9 1 10 9 1 12 9 2 13 15 3 1 9 0 2
35 10 9 13 9 7 1 11 13 16 10 9 13 3 0 1 10 9 2 1 0 1 10 9 11 11 2 10 9 1 0 9 1 10 9 2
12 1 13 1 9 2 15 4 13 10 9 0 2
30 10 12 1 11 1 12 15 13 1 10 9 7 10 12 1 11 1 12 15 13 10 0 11 11 1 11 1 10 11 2
14 13 0 1 10 9 12 7 13 12 9 7 12 9 2
18 10 9 13 10 0 9 1 10 9 7 1 15 3 15 4 1 13 2
14 13 3 0 2 10 9 13 0 7 10 9 13 3 2
29 9 3 3 2 1 10 9 1 15 11 4 13 3 2 10 9 15 13 1 12 9 2 10 15 10 9 1 11 2
20 1 10 9 0 1 10 9 15 13 9 1 10 9 1 10 9 1 10 11 2
16 1 9 1 9 13 10 9 1 11 1 10 9 11 2 11 2
38 1 10 9 1 10 9 0 9 0 4 13 3 1 15 1 10 0 9 1 11 1 10 11 2 3 1 11 11 2 11 1 11 2 11 11 7 11 2
28 7 10 9 13 4 15 3 13 1 16 2 3 10 9 13 3 2 2 10 9 0 13 13 3 9 1 9 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
33 10 9 13 1 10 9 0 1 11 2 11 11 2 11 1 11 2 11 11 2 7 11 2 7 1 10 9 0 1 11 10 11 2
19 1 16 11 13 7 11 13 2 10 9 13 1 10 9 0 13 1 15 2
54 1 9 15 3 13 0 9 16 10 9 13 2 7 16 3 1 9 1 10 9 0 1 10 9 13 10 9 1 10 9 11 11 13 1 9 13 10 9 2 13 7 13 12 9 16 3 4 13 10 9 1 10 9 2
26 1 9 2 13 10 9 10 12 1 11 2 10 9 16 10 9 7 10 9 1 10 9 3 4 13 2
31 7 1 10 9 1 10 9 1 11 2 13 10 9 1 10 0 9 1 10 9 12 7 3 3 4 13 15 1 10 9 2
14 15 1 10 9 15 13 1 10 9 0 1 9 0 2
32 15 4 13 9 1 13 15 1 16 10 9 0 1 10 9 1 10 9 0 13 10 9 2 1 10 0 9 1 10 9 2 2
41 10 9 13 12 9 9 1 11 13 10 0 9 1 10 9 2 13 1 10 0 9 7 13 1 10 9 1 10 11 11 1 11 8 2 12 1 13 15 1 11 2
25 9 1 10 9 11 1 11 7 11 1 11 7 11 2 9 0 1 10 9 11 1 11 7 11 2
29 16 4 13 1 10 9 0 11 2 11 1 10 11 2 11 2 10 12 1 11 1 12 13 10 9 0 7 13 2
12 11 11 13 10 9 1 9 1 10 9 11 2
13 1 12 1 12 2 11 13 0 7 1 13 9 2
16 10 9 0 15 4 13 1 10 9 0 1 10 9 1 9 2
12 13 8 2 9 1 10 9 0 2 10 9 2
41 10 9 0 13 10 9 1 12 9 5 7 13 1 11 1 10 9 2 11 1 10 9 7 1 10 9 2 1 10 9 11 7 11 2 10 11 2 1 10 9 2
33 15 13 1 10 9 1 11 2 1 3 1 12 9 13 1 9 1 9 0 13 1 13 9 1 10 9 13 1 10 9 7 9 2
19 11 11 13 7 10 9 1 0 9 7 16 3 3 13 1 10 9 0 2
21 1 10 9 1 11 15 13 1 11 11 2 1 15 4 1 13 1 10 9 0 2
27 3 4 13 10 9 1 10 0 9 0 1 11 1 11 2 2 11 10 11 2 2 13 1 10 9 12 2
24 10 0 9 1 11 2 11 11 2 15 13 1 10 9 10 12 1 11 1 12 1 11 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
10 15 13 3 1 10 9 1 9 0 2
29 10 0 9 2 9 2 13 1 9 2 9 7 9 3 13 1 10 9 1 10 9 1 10 3 0 2 9 2 2
8 10 9 13 10 9 0 0 2
30 10 11 11 12 11 11 2 2 9 2 1 9 2 13 10 9 1 9 0 13 1 12 9 13 1 10 9 0 11 2
22 3 4 13 1 10 0 9 1 12 9 1 10 9 0 7 12 9 1 10 9 0 2
26 10 9 1 9 0 13 1 10 12 5 1 10 9 2 7 16 10 12 5 4 13 1 10 10 9 2
9 15 13 1 15 1 10 11 11 2
16 10 9 4 13 1 0 9 1 11 2 11 2 11 7 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
24 11 13 10 9 0 1 10 11 1 11 2 1 12 5 5 1 9 7 12 9 2 12 2 2
14 15 15 13 1 10 9 0 1 10 11 1 10 11 2
20 11 13 10 9 1 15 16 13 1 10 9 1 11 2 13 15 1 15 0 2
40 10 9 2 10 9 1 11 7 11 7 10 9 1 9 1 10 9 4 13 1 12 9 10 9 1 11 1 10 16 10 9 0 13 12 9 1 9 1 12 2
59 3 1 13 10 9 1 10 9 1 10 9 2 16 15 13 10 9 4 13 10 2 9 2 1 9 1 9 1 10 9 1 10 9 11 11 1 11 1 8 10 9 4 13 10 0 9 16 13 10 9 0 1 10 0 9 1 10 9 2
24 10 9 3 4 13 10 0 9 16 13 10 11 1 11 1 10 9 1 9 1 10 9 0 2
29 10 9 2 1 12 9 1 9 2 13 7 10 9 7 10 9 1 10 9 15 13 2 15 16 13 10 0 9 2
32 11 11 11 2 3 0 1 11 2 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 2 13 10 9 0 0 2
27 10 9 1 11 7 11 4 13 3 2 16 11 4 13 10 9 0 2 13 9 1 3 1 10 0 9 2
37 1 11 11 15 13 10 9 3 0 13 1 10 9 1 10 11 2 10 16 1 9 1 10 9 4 13 10 12 9 1 9 2 16 13 9 0 2
28 1 10 9 2 11 3 15 13 9 1 10 9 3 13 2 13 10 9 9 1 10 9 0 1 10 9 0 2
8 10 9 0 13 10 9 0 2
49 11 13 1 0 9 1 10 9 1 10 0 11 11 11 11 11 2 12 2 2 7 13 10 9 1 10 9 1 9 0 1 10 11 11 2 11 2 16 10 9 13 16 3 13 3 1 9 0 2
25 13 1 11 1 12 2 13 1 10 9 11 11 2 15 4 4 13 1 11 11 1 10 9 12 2
8 4 3 13 3 4 13 9 2
45 1 10 9 0 1 10 9 15 13 10 9 1 10 9 1 9 1 9 3 1 10 9 7 9 3 7 10 9 1 10 9 13 1 9 1 9 16 13 13 10 9 1 10 9 2
16 1 11 7 12 9 15 13 1 15 3 1 11 7 12 9 2
38 10 9 13 1 11 2 11 1 9 2 2 4 13 1 10 9 1 12 2 16 4 13 15 2 2 13 1 15 2 1 10 9 1 9 13 11 2 2
121 13 10 9 2 11 2 1 0 9 1 9 2 2 10 11 2 2 2 11 2 2 2 9 0 7 13 2 2 2 13 0 2 13 0 2 2 7 3 13 10 9 2 11 11 1 11 2 1 15 8 1 2 2 1 11 15 11 2 15 11 2 2 2 15 2 2 2 11 15 11 1 10 11 2 10 15 15 13 15 1 9 1 9 3 7 1 9 2 1 9 1 10 9 13 0 1 10 9 3 0 1 10 9 2 2 9 1 10 11 2 1 10 15 15 13 7 13 1 10 9 2
40 1 10 9 1 9 2 10 9 13 10 11 1 11 1 11 1 12 2 1 10 11 11 1 10 9 2 7 3 13 9 1 9 1 10 11 1 11 1 12 2
35 10 9 13 0 2 10 9 13 0 2 7 15 13 13 3 2 16 13 0 9 2 1 0 10 9 1 9 2 16 3 13 1 10 9 2
19 10 9 1 10 9 13 0 2 1 0 9 1 10 9 1 10 15 13 2
16 10 9 0 13 1 11 11 3 2 13 10 9 1 0 9 2
8 10 9 13 7 13 1 11 2
21 10 9 13 10 9 1 10 9 1 11 1 11 2 4 13 1 0 9 11 11 2
28 3 15 13 10 11 1 11 11 1 11 1 10 9 8 5 12 7 11 5 12 7 1 10 11 1 10 11 2
42 10 9 3 2 13 10 9 1 10 9 1 10 9 1 10 9 11 11 7 10 9 1 9 1 9 11 11 7 11 11 11 2 15 3 15 4 13 1 10 0 9 2
25 11 1 11 2 11 11 2 11 11 2 12 1 11 1 12 2 2 13 10 9 16 3 13 9 2
42 2 13 16 3 13 10 9 1 10 9 7 1 13 10 9 1 9 7 9 1 9 13 0 10 9 2 2 13 1 11 2 10 9 0 1 11 1 11 2 11 11 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
33 13 10 9 1 10 11 7 11 1 10 11 2 13 1 10 9 2 1 9 1 10 9 2 9 7 9 1 9 3 7 3 0 2
27 1 10 9 1 10 9 1 10 12 2 11 3 13 3 7 3 2 1 9 1 10 12 13 9 10 9 2
36 11 1 11 13 10 8 0 1 10 9 11 11 11 16 13 1 10 9 1 10 9 1 9 0 2 10 11 2 16 10 10 9 13 9 0 2
45 10 9 10 9 3 0 2 12 2 2 10 9 0 2 12 2 2 1 9 2 12 2 7 11 2 12 2 4 4 13 1 10 9 2 10 9 1 9 0 2 2 13 9 0 2
22 1 11 2 15 13 16 10 9 7 10 9 13 0 2 7 3 15 13 16 15 13 2
19 10 9 13 10 9 1 11 1 9 0 7 13 10 9 0 0 1 11 2
38 1 8 8 1 11 2 11 4 13 1 12 1 10 11 11 11 11 1 10 9 1 8 7 13 10 11 11 11 2 1 10 0 8 8 1 10 9 2
10 13 10 9 0 1 13 10 9 11 2
24 1 13 1 10 9 13 1 11 11 1 12 2 7 10 0 9 13 10 0 9 1 10 9 2
14 3 1 10 9 1 11 11 13 10 9 1 10 9 2
21 13 10 9 3 1 10 11 2 10 9 13 1 10 9 2 3 1 13 15 3 2
31 10 0 9 13 1 10 9 2 11 11 2 2 12 2 2 1 10 15 13 10 9 1 10 9 13 1 10 13 1 9 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
35 10 9 11 12 13 9 0 1 10 9 11 7 10 9 1 11 2 16 13 10 9 7 16 1 0 13 10 9 1 10 9 0 2 11 2
29 1 9 0 13 10 9 0 2 0 1 10 10 9 7 16 15 13 1 10 9 3 0 1 10 9 1 10 9 2
7 13 1 12 9 7 9 2
77 10 2 0 2 11 11 2 13 2 11 2 1 10 9 0 11 2 13 1 11 1 11 1 11 2 16 13 10 9 1 10 9 10 11 2 13 10 0 9 1 11 11 11 2 10 9 1 10 11 11 7 11 2 11 2 2 3 11 4 13 7 13 1 11 11 1 15 13 2 3 7 16 15 13 10 9 2
19 10 9 0 7 9 0 1 11 2 15 13 3 1 10 9 0 1 11 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
21 15 13 3 0 13 7 10 9 0 13 12 2 12 1 10 8 1 10 9 11 2
18 10 9 0 1 10 9 0 13 3 1 10 9 0 1 10 9 0 2
51 10 9 3 3 13 1 10 9 7 1 12 2 1 9 1 10 9 11 2 13 2 3 2 1 10 9 1 11 1 10 9 11 11 11 7 11 11 11 2 3 7 1 10 9 1 10 9 11 11 11 2
27 13 10 9 1 13 10 0 9 0 1 10 9 2 13 16 13 10 9 1 13 2 13 7 13 10 9 2
20 10 12 1 11 1 12 4 13 9 1 10 11 1 11 1 9 1 11 11 2
6 11 13 10 9 0 2
16 9 1 10 11 11 1 11 1 10 11 11 1 10 11 8 2
24 11 11 13 10 9 10 10 9 1 10 9 2 3 11 7 11 11 13 7 13 10 9 0 2
28 10 9 7 10 9 1 15 4 13 1 0 9 1 10 9 1 11 7 13 9 1 16 15 4 13 1 15 2
70 3 13 10 12 5 1 9 1 10 9 1 9 1 10 9 1 11 2 13 10 9 1 10 11 1 10 11 11 2 11 11 7 11 11 11 2 15 13 16 10 9 1 10 11 11 16 13 9 1 10 9 1 11 11 2 4 1 13 15 7 2 16 3 3 15 13 1 15 2 2
26 10 9 0 1 10 9 13 16 3 1 10 12 15 13 1 10 9 1 10 9 1 10 11 1 11 2
22 11 13 15 1 10 3 9 7 0 1 10 11 13 15 3 13 1 10 0 9 0 2
42 1 9 1 10 12 9 1 10 9 1 11 11 2 11 11 11 13 10 9 8 8 8 11 11 2 1 10 9 7 10 9 13 2 13 16 10 9 13 3 3 13 2
7 2 4 1 13 10 9 2
24 11 13 10 9 0 1 10 9 1 11 2 1 12 9 5 1 9 7 12 9 2 12 2 2
41 0 2 16 13 10 9 13 1 10 9 2 7 10 9 16 15 13 1 9 2 1 9 7 1 9 13 3 0 7 3 4 13 15 13 1 10 9 2 16 13 2
39 10 9 0 13 10 9 1 10 9 1 10 11 11 2 15 4 4 13 1 10 0 9 1 10 9 12 7 15 13 1 9 0 3 1 10 9 1 12 2
27 10 9 1 9 13 0 1 10 9 9 1 10 11 1 11 1 11 2 5 2 8 2 8 8 2 2 2
14 1 10 9 1 12 2 13 12 9 13 1 11 11 2
19 13 10 11 0 7 10 9 0 4 13 1 15 1 10 9 1 10 9 2
26 13 10 9 2 16 1 10 9 0 15 13 10 9 2 4 13 0 9 7 13 15 3 1 10 9 2
52 2 3 1 13 15 7 10 0 9 2 13 16 3 15 13 16 13 10 9 1 10 9 1 11 11 1 12 2 2 13 11 2 9 1 10 9 0 1 11 11 1 12 2 1 10 9 13 1 10 9 0 2
16 11 7 11 15 13 1 11 11 7 11 11 7 13 1 15 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
24 10 9 1 11 2 15 0 1 11 2 10 11 2 13 1 11 2 11 3 3 1 10 9 2
30 3 1 9 10 9 0 15 13 1 11 2 11 2 7 13 9 1 11 2 11 2 11 2 11 7 10 11 11 11 2
40 1 10 9 11 12 13 1 10 9 1 10 9 11 7 16 4 13 4 7 13 3 0 10 9 16 15 13 2 7 15 13 16 13 15 2 10 15 15 13 2
42 10 9 7 9 0 16 13 1 13 1 10 9 1 10 9 7 13 10 9 1 0 9 2 1 10 9 2 1 15 15 3 4 13 10 9 7 15 13 10 9 0 2
23 16 15 0 3 13 3 1 10 9 1 10 9 1 12 9 2 10 9 13 1 9 3 2
14 3 7 3 13 0 1 11 2 3 13 9 1 9 2
28 10 9 1 11 11 11 11 13 10 9 0 1 9 0 1 10 9 1 10 9 0 1 11 1 12 1 12 2
17 10 9 11 12 1 11 13 11 1 12 2 13 1 11 1 11 2
32 1 10 9 2 11 10 9 1 15 13 2 7 15 11 11 1 11 13 1 13 1 10 11 11 1 11 1 10 9 0 0 2
29 15 13 3 1 10 9 1 10 11 11 2 3 12 9 1 10 9 1 11 2 7 12 9 1 10 9 1 11 2
29 11 13 10 9 3 0 2 7 1 15 2 15 4 13 1 10 9 0 9 7 9 10 9 16 10 9 15 13 2
21 15 13 8 1 10 9 1 10 9 2 0 9 7 9 2 10 9 1 10 9 2
21 1 10 9 13 1 11 1 10 9 1 9 7 9 1 10 0 9 0 1 12 2
15 10 9 3 4 1 13 16 3 13 10 9 1 10 9 2
31 1 10 9 1 10 9 0 10 9 0 13 10 0 9 1 10 12 9 1 9 2 1 15 4 13 1 13 1 9 0 2
26 3 13 10 0 9 0 1 10 9 7 3 4 13 1 10 9 2 15 1 9 7 3 1 10 9 2
38 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 2 9 1 11 11 2 1 10 9 1 11 2 1 2 11 7 9 1 11 2 11 2
12 10 9 13 0 1 10 9 1 11 1 12 2
22 1 9 2 1 10 13 10 9 10 9 15 13 1 11 1 12 1 11 2 11 11 2
6 3 3 13 10 9 2
18 10 9 1 10 9 3 13 2 10 9 13 9 7 3 13 12 9 2
7 10 9 0 13 10 9 2
17 11 13 10 11 13 1 10 9 1 11 1 10 9 0 1 11 2
29 11 11 13 10 9 1 9 0 1 10 9 1 11 2 1 10 9 1 10 9 1 11 2 2 11 2 11 2 2
34 1 13 16 10 12 5 1 10 9 1 11 11 7 11 13 9 2 10 9 0 1 10 9 13 10 9 2 13 1 10 12 5 2 2
14 15 13 10 8 8 8 8 2 13 9 3 3 2 2
42 10 9 15 13 1 10 9 1 9 2 16 13 1 10 12 5 1 9 0 2 1 10 12 5 1 9 0 2 13 1 10 9 1 10 12 5 2 16 13 9 0 2
24 4 13 10 12 1 11 1 12 1 10 11 7 13 9 1 10 9 0 1 11 11 1 12 2
13 11 13 10 9 1 10 9 11 1 10 9 11 2
52 1 15 4 7 13 16 10 0 9 1 9 2 9 0 1 9 0 2 9 1 9 0 1 10 9 1 11 1 10 11 11 2 9 1 9 7 9 0 1 10 9 1 11 8 2 7 10 9 1 11 11 2
15 10 9 11 11 7 11 11 13 16 10 9 3 13 0 2
36 10 9 1 10 11 11 11 2 11 2 13 10 9 0 1 9 0 1 9 0 1 0 9 2 0 1 9 2 9 2 9 2 9 7 9 2
36 10 9 1 9 4 13 1 13 10 9 0 1 10 9 2 13 1 9 1 10 9 1 9 0 10 9 1 9 1 10 9 13 3 1 11 2
19 10 9 2 0 2 16 3 4 13 10 9 1 10 0 9 1 15 9 2
28 12 9 3 2 11 13 1 9 1 10 9 11 16 4 13 1 11 2 13 10 9 1 9 13 1 10 11 2
28 9 1 12 9 1 12 9 1 0 2 1 12 9 0 1 10 9 1 10 9 0 7 1 10 12 9 0 2
43 10 9 1 10 11 11 13 10 0 9 2 1 15 16 15 4 13 15 1 10 9 2 9 16 13 16 13 1 12 0 9 9 7 12 16 13 16 3 15 13 10 9 2
32 10 9 3 0 13 10 9 1 10 11 1 10 11 2 12 8 2 2 9 1 9 1 10 9 1 10 11 7 11 2 11 2
18 10 9 1 10 11 11 13 10 0 1 13 10 9 1 10 0 9 2
56 1 10 9 15 13 16 2 10 9 1 10 9 1 9 7 9 3 4 13 0 1 10 9 1 10 9 0 1 9 2 7 15 13 1 10 0 9 1 15 15 13 9 7 9 1 10 9 1 10 9 1 10 9 9 2 2
39 10 9 1 11 13 10 9 1 9 0 1 10 9 0 1 9 1 10 9 7 10 9 3 0 2 7 10 9 1 9 0 3 13 16 15 13 3 0 2
11 10 11 13 10 0 9 16 13 10 11 2
13 13 9 1 10 9 1 9 11 2 0 1 11 2
9 13 3 0 7 0 1 10 9 2
13 1 10 9 15 4 13 1 10 0 7 0 9 2
9 1 3 13 3 0 1 10 9 2
39 16 10 9 0 1 10 10 9 3 13 10 9 2 7 10 9 0 3 0 1 10 9 2 13 0 13 16 10 9 3 13 0 7 0 1 13 15 3 2
47 10 0 11 13 1 10 9 2 3 1 0 9 15 13 10 9 0 2 1 9 1 9 1 10 10 9 0 2 3 7 15 13 10 9 16 13 10 0 9 1 10 0 9 1 10 9 2
21 1 12 15 13 1 11 1 11 7 11 1 13 10 9 1 11 11 7 11 11 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 4 1 9 0 7 2 12 5 2 12 5 5 13 9 2
32 3 2 16 13 1 10 9 2 11 4 13 1 10 9 7 1 10 9 2 13 1 10 0 9 0 7 0 7 1 10 9 2
33 15 1 12 9 16 15 13 1 11 1 0 9 7 9 7 16 1 10 13 15 1 12 10 11 1 11 13 1 10 11 1 11 2
10 10 9 15 13 13 1 10 9 12 2
42 13 10 9 10 9 7 13 16 10 9 4 4 13 1 10 0 9 16 4 13 1 11 3 15 13 0 10 11 7 15 13 0 10 9 1 11 3 16 13 11 11 2
15 7 1 10 9 13 3 1 10 9 0 2 0 7 0 2
35 1 10 9 2 10 9 0 13 10 9 1 10 9 0 2 3 7 10 9 0 2 3 13 2 13 10 9 7 10 9 1 10 9 0 2
22 10 11 1 11 13 10 9 0 1 9 1 11 7 10 9 0 1 11 2 1 11 2
45 11 2 13 1 12 1 11 2 11 2 13 10 9 1 9 2 10 11 11 1 10 9 0 2 16 15 4 13 1 10 9 1 11 1 13 1 12 1 10 9 2 10 11 11 2
19 15 15 13 3 1 9 13 7 1 9 7 1 9 7 9 1 10 9 2
11 3 13 10 9 1 12 2 12 7 12 2
27 1 9 1 3 13 0 2 13 1 10 9 11 11 7 1 10 9 2 7 15 0 3 13 10 9 0 2
45 10 9 1 11 2 10 9 0 2 13 1 10 9 2 13 16 10 9 15 13 1 11 16 13 15 2 16 3 15 13 9 10 9 15 15 13 1 10 9 2 1 0 1 11 2
18 10 9 13 10 9 0 1 9 12 3 1 10 9 12 1 10 9 2
42 15 16 13 9 1 0 9 2 1 3 13 16 13 3 0 2 13 10 9 2 11 16 10 0 11 13 10 9 1 9 1 10 9 13 1 11 1 10 11 1 11 2
29 1 9 2 11 13 1 10 11 7 4 13 1 10 9 0 11 2 7 11 15 13 16 15 13 15 15 16 13 2
35 3 13 10 9 1 13 15 1 10 9 1 10 13 3 10 9 7 3 4 13 10 9 1 10 9 0 1 10 9 1 13 10 9 0 2
29 9 1 10 9 0 1 9 0 2 8 2 13 10 0 9 13 1 10 9 1 10 9 7 10 9 1 10 9 2
56 3 3 2 10 9 0 4 13 1 12 9 0 10 9 0 2 3 13 1 10 9 1 11 1 12 7 12 2 1 10 9 1 10 9 0 1 9 2 8 2 2 11 11 2 15 3 13 16 11 13 0 1 0 7 11 2
13 10 9 1 10 9 1 12 9 13 10 0 9 2
28 2 3 13 16 3 13 10 9 0 2 2 13 1 11 10 9 1 11 11 7 9 1 10 11 2 11 11 2
52 1 10 10 9 15 13 9 1 10 9 1 9 0 7 9 1 10 9 0 2 3 7 1 10 9 1 10 9 7 10 9 1 9 1 10 9 0 2 9 15 4 13 1 10 9 0 13 1 10 0 9 2
20 10 9 4 4 13 1 10 0 12 9 2 1 9 1 9 1 9 7 9 2
25 13 9 1 12 9 0 13 15 1 10 0 9 2 7 1 10 15 15 4 13 3 1 12 9 2
43 1 10 9 1 11 2 11 13 16 10 9 13 9 1 10 9 2 3 2 1 10 12 9 1 9 2 13 10 12 1 11 1 10 9 16 10 11 2 0 13 11 11 2
27 1 10 0 9 10 9 11 11 13 1 9 1 10 9 2 7 1 12 10 9 11 11 13 1 11 11 2
16 1 9 1 9 0 13 10 9 0 2 0 2 0 7 0 2
20 10 9 4 13 10 9 7 9 16 15 13 1 10 9 1 9 7 1 9 2
24 16 10 12 9 1 10 11 7 10 11 2 11 2 15 13 1 12 2 10 0 9 4 13 2
36 10 9 1 10 9 1 11 1 10 9 1 10 9 1 13 1 9 10 0 9 0 3 4 13 3 0 7 13 10 9 1 10 9 1 11 2
22 10 0 9 15 13 10 12 1 11 3 3 13 10 12 9 1 11 16 3 3 13 2
48 1 10 11 11 11 11 13 10 9 1 2 2 0 9 2 2 2 0 9 2 2 2 0 9 2 2 11 2 2 2 0 9 2 2 11 11 2 7 2 0 9 2 2 11 11 11 2 2
7 15 4 13 10 10 9 2
24 13 10 9 1 9 0 1 9 11 16 13 1 12 1 12 5 2 1 0 9 1 9 0 2
45 1 10 9 2 10 9 1 9 7 10 9 1 10 9 15 4 13 0 7 1 10 9 0 10 9 1 10 9 1 9 7 9 13 10 9 1 4 13 10 9 0 1 13 9 2
32 10 9 2 1 9 2 13 16 10 9 13 0 7 0 7 16 10 11 11 3 3 13 0 1 10 9 0 2 0 7 0 2
27 11 3 13 12 11 11 12 1 10 9 11 11 11 11 2 3 7 10 9 1 12 9 1 10 0 9 2
37 13 10 0 9 1 11 11 2 10 9 1 9 2 16 13 10 9 1 10 9 1 10 11 1 10 11 1 11 2 7 1 11 11 2 10 9 2
19 11 11 2 12 2 12 2 13 10 9 2 9 1 9 2 7 9 0 2
31 1 10 9 13 1 10 9 2 11 1 11 13 10 9 1 11 1 11 11 7 11 1 11 2 11 2 11 7 10 11 2
32 13 10 0 9 2 1 15 15 13 10 9 1 10 9 0 7 13 10 9 3 16 10 9 0 13 10 9 1 13 3 0 2
34 10 9 13 13 15 1 10 9 11 1 10 11 1 13 15 1 10 9 1 10 11 2 13 15 9 7 13 10 9 1 11 1 11 2
72 1 10 9 13 1 12 9 1 10 9 1 10 9 0 11 11 2 1 11 2 10 9 0 13 1 12 9 1 9 9 1 10 9 7 9 1 10 11 1 9 0 1 10 9 1 10 9 2 10 9 1 10 9 0 1 10 9 0 7 10 9 0 1 10 9 1 10 9 2 1 15 2
2 10 9
8 0 9 1 13 1 10 9 2
13 11 15 13 2 1 9 2 1 13 15 1 15 2
10 1 11 1 10 9 2 13 10 11 2
44 1 10 9 2 10 9 3 13 3 10 9 1 9 0 3 0 2 1 9 1 10 11 11 2 10 9 0 3 13 3 1 9 0 7 13 10 0 9 1 10 9 0 0 2
71 2 10 9 13 0 7 3 13 9 2 13 11 2 7 13 16 13 2 3 7 1 9 2 10 9 1 10 9 0 2 11 11 2 1 10 9 11 2 1 10 9 2 11 2 2 7 2 11 12 2 2 1 9 1 10 9 1 11 7 3 1 10 9 1 9 0 11 16 13 11 2
19 10 9 0 1 10 9 1 10 9 2 11 2 13 2 11 1 11 2 2
28 10 9 11 2 3 13 1 9 0 0 2 15 13 1 10 9 0 1 10 9 13 1 10 9 0 1 9 2
10 1 10 9 2 10 9 13 3 0 2
18 11 11 11 13 10 9 1 9 0 7 1 9 13 3 13 1 12 2
22 11 11 13 10 9 0 0 1 11 11 2 3 13 10 9 0 1 9 9 1 9 2
30 3 2 10 9 13 1 10 9 13 10 9 1 9 1 10 9 0 1 9 0 13 1 11 2 11 11 11 11 2 2
29 3 1 13 10 9 1 15 15 13 10 9 2 15 13 1 10 2 11 11 2 3 13 10 9 0 1 10 9 2
24 15 10 9 1 10 9 10 11 1 10 11 13 10 9 12 1 11 3 1 10 9 1 9 2
18 1 0 7 10 9 11 11 13 1 10 9 2 13 1 10 9 12 2
23 13 1 10 9 1 9 2 13 15 10 9 0 1 12 9 1 11 2 3 1 16 13 0
29 10 9 1 9 0 7 0 1 12 9 16 13 7 13 16 4 13 1 10 9 1 10 9 1 13 15 3 7 3
29 11 11 13 9 2 13 1 10 9 11 2 1 10 0 7 1 2 11 2 11 11 2 2 1 10 15 11 13 2
17 11 13 10 9 3 0 1 16 13 2 1 15 15 15 13 0 2
26 3 2 10 9 15 4 13 13 1 10 9 15 4 1 10 3 2 15 16 13 3 3 13 10 9 2
29 10 9 1 9 1 10 9 2 3 13 9 0 2 4 4 13 3 1 10 9 1 9 1 10 9 16 15 13 2
34 1 15 15 4 13 10 9 1 9 11 13 10 9 1 11 11 7 11 1 10 11 2 13 0 3 13 1 12 7 12 1 9 2 2
12 10 9 12 13 1 11 13 15 11 11 11 2
34 11 13 1 11 2 11 10 12 1 11 1 12 2 9 15 4 13 1 9 1 10 9 2 1 10 9 0 13 10 12 1 11 2 2
19 10 12 1 11 1 12 2 4 13 10 9 1 11 1 10 9 1 11 2
29 1 12 2 1 4 15 13 10 11 1 11 2 11 1 11 15 13 9 1 9 0 7 9 1 10 11 11 11 2
27 12 9 1 10 9 11 11 2 1 10 9 11 11 2 1 12 9 1 11 11 11 2 13 1 10 9 2
12 10 12 0 9 13 1 13 12 9 1 8 2
19 1 10 0 9 15 13 10 8 8 2 5 2 0 2 0 2 11 2 8
33 1 10 9 1 10 12 10 9 1 9 0 1 10 9 1 10 9 13 1 12 9 7 10 9 0 1 10 9 13 1 12 9 2
38 3 2 13 1 16 10 9 1 10 0 9 1 10 9 4 13 10 1 2 10 9 7 10 9 2 2 9 16 2 2 3 13 1 10 0 9 2 2
7 15 13 1 9 1 9 2
38 10 0 9 16 4 13 13 2 11 13 2 2 1 10 16 9 1 11 1 11 2 11 11 1 11 11 7 11 11 13 1 13 10 9 0 1 13 2
31 10 0 9 2 11 2 12 2 2 15 13 1 10 9 1 10 9 11 1 9 1 10 9 2 10 9 0 2 1 12 2
20 9 0 13 10 9 1 10 9 2 1 10 11 1 12 1 10 9 1 12 2
24 2 1 10 9 1 10 9 2 3 13 9 16 10 9 15 13 1 10 9 7 13 1 9 2
11 15 13 1 11 2 7 10 9 0 13 2
45 10 9 0 1 11 11 2 11 11 11 15 13 1 10 0 9 13 1 10 8 9 1 11 12 2 11 11 2 15 1 10 9 2 13 10 9 2 7 1 9 4 2 13 2 2
30 10 9 11 11 13 1 10 9 1 10 15 8 10 9 1 2 9 2 0 13 0 2 13 2 10 9 1 10 9 2
15 10 9 13 1 9 10 9 0 1 1 12 9 1 9 2
42 10 9 13 1 9 0 1 10 9 12 13 15 1 13 1 10 9 1 10 9 0 1 10 9 2 9 1 10 11 0 9 7 11 11 2 16 13 11 1 9 0 2
101 1 10 9 1 10 9 10 9 0 1 10 9 2 9 0 13 1 9 1 10 11 2 13 10 9 0 1 9 7 10 11 11 13 2 13 3 1 10 9 1 10 9 2 1 10 9 1 10 9 1 3 9 2 1 10 9 1 10 9 7 9 1 10 9 1 9 0 7 0 2 15 1 9 2 9 2 9 2 9 2 9 2 9 0 2 9 1 9 2 9 2 7 1 10 9 1 10 9 1 11 2
24 10 11 11 11 2 3 13 11 1 10 11 2 15 13 1 11 2 9 1 11 2 11 2 2
21 10 9 1 9 1 9 2 0 1 10 9 9 7 16 3 13 10 9 1 9 2
13 13 10 9 7 10 9 1 10 9 1 10 9 2
27 4 1 13 15 9 13 16 15 4 13 10 9 8 1 10 9 16 13 1 3 4 15 13 1 10 9 2
27 10 9 2 1 9 1 11 2 13 1 12 10 9 8 8 8 1 10 0 9 0 1 10 9 1 11 2
29 10 9 1 10 9 0 13 1 10 9 1 11 11 2 9 1 9 7 11 11 2 9 0 7 0 1 10 9 2
11 10 9 13 0 1 9 16 3 13 9 2
11 13 0 7 13 1 10 9 7 10 9 2
11 3 13 1 11 11 1 10 9 11 11 2
25 13 13 1 9 0 2 16 10 9 11 11 11 13 10 9 3 0 1 10 9 7 9 1 9 2
17 9 3 3 15 13 10 9 3 0 13 1 10 9 1 10 9 2
9 10 9 13 1 9 1 11 11 2
33 11 13 10 9 7 9 0 13 1 10 9 1 11 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2 11 2 11 2
19 11 11 13 1 12 1 10 9 1 10 9 13 1 10 9 1 10 9 2
30 10 16 13 1 10 9 10 9 7 13 10 9 1 10 9 2 2 3 13 16 15 13 10 9 16 3 13 12 9 2
49 11 11 11 2 11 2 11 2 12 1 11 1 12 2 10 11 2 11 2 12 1 11 1 12 2 13 10 9 9 2 9 0 16 15 13 0 1 10 9 12 1 10 9 9 7 9 2 9 2
16 15 13 12 1 11 11 1 10 15 13 10 0 9 1 9 2
25 10 9 13 16 10 9 3 13 1 10 9 16 13 0 1 9 7 13 1 10 10 9 1 9 2
67 1 10 9 7 2 10 9 1 9 15 13 1 9 1 9 2 10 9 0 1 13 9 1 9 0 2 3 13 3 1 9 0 2 7 9 1 9 7 1 13 0 7 0 2 9 0 1 13 9 7 13 9 1 9 7 9 1 0 2 13 3 1 9 1 13 2 2
7 12 1 10 11 2 11 2
13 10 0 9 12 13 1 10 12 5 1 0 9 2
16 10 15 3 1 10 9 4 13 9 1 10 9 0 1 9 2
47 1 10 10 9 4 13 16 11 11 13 13 1 10 11 11 2 1 9 3 15 13 10 9 1 10 9 10 3 9 11 11 1 10 9 1 9 15 1 10 9 1 9 7 3 1 15 2
41 15 9 13 16 15 13 1 10 9 15 0 13 1 9 10 9 2 7 3 15 13 13 3 9 3 13 4 13 1 10 9 1 9 2 0 2 1 10 9 0 2
33 11 2 16 4 13 10 9 0 1 11 15 13 1 15 2 16 3 4 7 13 15 9 16 4 4 7 13 10 9 0 0 3 2
22 3 1 12 9 13 2 2 13 1 3 10 9 1 16 15 13 3 1 13 1 9 2
31 11 2 11 7 11 2 1 10 9 1 10 9 1 11 2 13 10 9 1 10 9 2 10 9 0 7 10 9 13 13 2
26 3 2 11 13 10 9 1 9 7 9 1 13 1 11 2 7 10 9 1 15 7 10 9 13 0 2
21 11 11 11 12 13 10 9 1 0 9 1 10 9 1 9 1 10 11 1 11 2
7 11 11 13 9 1 11 2
32 13 3 0 2 3 13 9 1 10 9 2 16 13 9 4 7 13 12 9 3 2 1 10 9 3 13 9 7 1 10 9 2
33 4 13 1 10 9 1 12 9 2 10 9 1 10 9 0 1 10 9 7 10 9 1 10 9 1 11 1 10 9 0 1 11 2
34 1 12 2 15 13 1 10 9 1 10 9 11 11 2 9 2 2 13 1 11 2 11 2 11 2 10 9 2 9 0 1 10 9 2
12 3 13 12 9 1 9 1 3 1 12 9 2
17 11 13 16 10 9 13 10 9 0 1 10 9 0 1 10 9 2
46 13 1 15 2 10 0 9 1 9 1 9 0 2 11 11 2 11 11 7 11 2 2 9 16 4 13 10 9 1 9 0 3 0 2 13 11 11 2 11 1 11 11 1 11 11 2
5 2 9 7 9 2
25 1 10 9 11 2 0 2 13 16 10 9 1 11 15 13 1 15 3 7 1 9 1 10 9 2
6 13 9 7 9 0 2
32 3 10 9 15 4 13 1 10 9 2 13 13 10 9 0 7 0 1 10 9 0 2 13 15 3 10 0 9 1 10 9 2
18 13 1 9 1 11 11 2 1 10 15 13 3 1 9 1 10 9 2
24 13 3 16 10 9 1 11 11 1 11 11 2 4 13 1 10 9 1 10 9 1 9 2 2
12 1 10 9 15 13 10 9 0 1 10 9 2
11 2 1 9 1 12 9 13 1 9 2 2
43 2 15 15 13 10 9 1 10 9 7 3 13 15 16 4 13 2 7 13 13 10 9 16 15 13 10 9 3 2 1 10 9 1 10 9 2 1 10 9 1 9 2 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
30 13 10 9 1 8 9 7 4 13 3 1 9 1 9 7 9 1 9 2 9 1 9 1 12 7 1 0 1 12 2
26 3 13 3 1 13 15 10 9 7 9 11 11 2 11 13 11 11 10 12 1 11 1 10 9 12 2
23 13 10 9 16 10 9 13 11 11 4 13 10 9 1 15 1 10 9 1 10 9 11 2
16 13 1 9 10 9 12 1 11 1 12 1 10 11 9 11 2
68 1 10 9 0 10 11 4 13 1 10 11 11 2 11 11 11 2 11 11 7 11 4 13 9 2 7 10 9 2 1 10 11 11 16 10 9 1 10 11 11 13 1 10 9 11 11 13 10 9 1 13 10 9 1 13 1 3 4 15 13 1 10 9 1 12 7 12 2
18 10 11 3 13 10 9 0 1 11 11 2 15 16 3 13 1 11 2
26 1 10 0 12 9 2 10 9 4 13 0 9 13 1 10 9 1 13 1 10 9 1 9 7 9 2
55 10 9 8 11 11 11 2 11 11 11 1 10 9 2 4 13 1 12 7 13 9 1 10 9 1 12 2 3 4 13 1 10 9 2 3 13 1 11 11 11 2 9 1 11 11 2 1 10 10 9 1 10 11 11 2
36 10 9 11 11 13 10 9 0 1 9 1 11 2 11 2 11 11 2 11 2 2 13 1 12 2 7 16 3 13 1 10 9 1 11 11 2
63 1 10 9 0 13 10 9 1 10 9 1 10 9 7 10 9 1 10 9 1 10 9 0 1 10 0 9 16 10 0 9 0 13 3 10 9 2 10 9 0 4 13 1 10 9 1 10 9 7 10 9 1 10 9 3 0 1 10 9 13 9 0 2
19 10 9 1 9 7 12 1 9 13 1 10 9 1 11 1 10 9 0 2
16 10 9 4 13 10 9 7 10 9 16 15 4 13 12 9 2
33 13 1 9 1 10 9 10 9 0 1 10 9 7 9 0 2 2 9 2 1 10 9 0 0 1 11 2 16 13 10 0 11 2
26 15 13 1 10 0 9 1 9 1 10 10 9 9 1 11 2 7 1 11 2 11 2 11 7 11 2
9 1 10 9 0 3 15 13 0 2
23 10 9 0 4 13 1 12 1 10 9 0 1 10 11 11 11 2 13 1 11 11 11 2
10 3 2 12 2 10 9 13 2 11 11
22 7 13 9 1 9 2 7 11 7 11 2 1 10 9 2 13 10 9 1 10 9 2
10 11 7 11 13 9 1 10 10 9 2
26 10 9 4 13 10 9 0 3 13 16 15 4 13 16 13 1 10 9 0 1 10 9 1 11 11 2
28 10 9 0 1 10 9 1 11 13 10 9 1 9 3 0 1 10 9 3 13 1 10 9 1 11 7 0 2
18 10 9 1 9 13 10 9 13 1 9 0 16 13 1 10 4 13 2
23 3 15 13 1 10 9 0 9 1 10 9 1 11 7 13 10 9 3 1 10 9 0 2
12 1 10 9 9 4 13 15 1 11 1 11 2
47 10 9 0 1 10 11 13 13 10 9 2 3 10 9 2 3 7 13 10 9 1 11 16 15 13 1 10 11 1 10 9 1 12 9 1 9 7 3 13 13 7 10 9 1 10 9 2
9 13 13 0 2 7 3 15 13 2
14 13 15 3 9 1 10 11 1 11 7 10 9 0 2
55 1 10 9 1 12 15 13 1 10 9 0 2 4 13 2 1 10 9 11 11 11 2 11 1 11 2 11 7 11 1 10 11 1 11 1 11 2 11 11 2 2 1 10 15 13 3 10 9 1 11 2 11 7 11 2
64 2 10 9 13 12 9 1 9 7 3 15 4 13 15 7 15 4 13 1 9 10 0 9 2 0 9 2 10 9 16 4 13 10 9 10 9 2 2 13 11 2 16 13 1 10 9 1 13 10 9 7 13 15 1 10 0 9 16 4 4 13 1 11 2
47 10 9 1 10 9 13 0 7 15 13 1 10 9 10 9 0 7 1 9 0 16 15 13 1 15 1 10 9 0 1 10 9 2 7 15 13 2 3 2 1 13 15 16 11 13 0 2
43 10 9 2 9 7 9 0 2 11 11 2 13 10 9 1 9 0 1 10 9 1 10 9 2 15 1 10 12 16 15 13 3 1 10 9 7 15 4 13 3 1 11 2
7 15 13 10 9 1 9 2
33 13 15 3 2 13 10 0 9 2 10 9 7 10 9 1 9 2 13 1 10 9 0 7 13 1 10 0 9 1 9 1 9 2
28 1 10 9 2 1 9 1 10 9 2 15 13 13 16 4 4 1 13 1 10 9 7 13 3 9 1 15 2
19 11 13 10 9 0 1 10 11 1 11 11 2 9 1 11 11 2 11 2
26 13 1 10 9 0 13 1 10 9 1 11 2 9 1 11 2 1 10 9 1 10 9 1 11 11 2
18 10 0 9 1 11 15 13 1 9 1 10 9 12 1 10 9 12 2
21 9 7 9 1 11 1 11 2 13 1 11 10 0 11 11 1 10 11 11 11 2
22 10 9 0 1 9 4 13 1 10 9 3 0 13 1 10 9 1 10 9 1 9 2
26 13 10 0 9 1 9 13 1 10 15 13 1 10 9 2 13 9 2 9 2 9 0 7 9 0 2
23 10 9 0 1 10 9 13 16 10 9 1 9 3 4 4 13 1 10 9 1 10 9 2
48 10 9 11 11 2 11 11 2 15 13 10 9 1 10 9 1 11 1 11 2 13 1 15 9 1 11 11 2 11 11 2 15 4 13 1 10 0 9 0 1 9 2 11 2 11 11 2 2
19 4 7 13 1 10 9 16 13 10 0 9 2 9 16 15 13 9 3 2
11 3 13 10 9 0 1 13 15 1 9 2
27 1 15 15 13 10 9 1 11 11 2 1 10 9 1 10 11 11 2 7 1 9 1 15 10 9 0 2
27 1 12 2 10 11 13 10 9 0 1 10 9 2 3 3 1 9 13 10 9 0 7 0 2 11 2 2
78 11 15 13 1 10 9 1 11 12 9 1 8 11 15 13 1 10 9 1 11 2 1 10 13 9 0 16 13 1 10 9 1 11 2 1 10 9 1 11 8 2 1 10 13 10 0 9 1 10 11 11 1 11 2 9 8 9 2 13 1 10 9 12 1 10 11 1 11 11 7 11 1 11 1 10 11 11 2
12 15 13 3 2 10 9 13 0 2 3 0 2
38 13 10 9 1 10 9 1 13 1 10 9 2 13 15 7 13 3 10 9 1 10 15 16 3 15 13 9 1 2 3 2 13 1 15 1 10 11 2
35 1 9 1 10 9 0 13 15 1 10 9 1 10 9 1 16 10 9 1 10 11 15 13 1 9 2 13 13 2 16 13 10 9 0 2
20 10 9 13 3 0 2 7 13 3 0 2 1 9 0 1 9 0 2 0 2
20 10 9 13 9 7 1 10 12 1 10 9 1 15 15 4 13 7 3 13 2
9 11 15 13 0 1 10 9 11 2
28 10 11 9 12 3 13 9 2 7 13 0 9 0 7 13 10 9 0 1 10 9 0 1 9 2 11 2 2
15 10 9 13 0 1 11 2 13 15 1 12 1 11 11 2
25 11 11 7 11 2 11 2 11 2 12 2 11 2 11 12 2 13 10 9 7 0 0 1 11 2
23 13 1 10 11 2 1 11 11 7 3 1 10 11 11 11 11 2 3 13 10 9 0 2
7 2 10 9 15 13 3 2
30 10 9 1 9 13 12 9 2 10 9 0 7 10 9 0 7 0 2 16 13 10 9 0 7 0 1 10 9 3 2
33 13 1 16 10 9 3 13 16 15 13 1 12 9 2 3 1 12 9 15 13 16 13 10 9 7 3 3 1 16 15 13 0 2
25 10 9 0 1 10 9 15 13 1 13 3 10 9 2 16 13 16 10 9 0 13 0 7 0 2
19 10 9 0 4 13 1 12 1 10 9 1 10 2 11 1 15 11 2 2
22 13 0 16 1 12 13 10 9 1 10 9 1 11 7 10 9 1 10 9 1 11 2
19 10 9 1 9 7 9 1 10 9 13 10 9 0 1 13 10 0 9 2
31 11 11 13 10 9 0 1 9 13 10 12 1 11 1 12 1 11 2 11 16 13 1 10 11 11 1 10 9 11 11 2
13 4 13 9 2 15 15 1 15 15 13 10 9 2
14 11 11 4 13 16 1 15 2 13 10 9 0 2 2
13 10 13 10 9 1 11 16 13 10 9 1 11 2
12 3 4 13 15 0 1 10 11 7 10 11 2
9 3 10 0 9 2 11 7 11 2
11 3 2 10 0 11 11 15 13 1 9 2
44 13 10 9 1 10 9 0 1 9 13 1 10 9 1 10 2 9 2 2 7 10 9 13 1 0 9 16 1 10 9 13 1 15 15 15 4 13 1 2 0 9 0 2 2
38 0 9 2 1 10 11 11 11 11 2 11 11 2 11 11 7 15 2 13 16 10 2 9 2 4 1 13 1 10 9 13 1 10 9 1 10 9 2
29 10 9 11 2 11 13 10 9 1 10 11 11 2 11 11 2 11 11 7 11 11 2 0 1 9 1 10 9 2
36 1 9 2 16 13 9 0 1 9 2 13 0 1 13 10 9 1 10 9 0 1 9 2 16 4 1 4 13 1 10 2 9 1 11 2 2
20 13 10 9 1 10 9 1 9 1 11 16 13 9 1 10 9 7 15 13 2
16 10 8 2 12 15 13 1 11 2 11 2 11 7 1 9 2
13 10 9 13 1 10 9 7 10 9 15 4 13 2
17 1 10 9 1 10 9 0 1 10 11 1 11 13 3 10 9 2
5 1 12 13 12 2
41 7 3 13 0 1 10 12 9 11 2 11 2 16 13 12 9 16 13 10 9 1 9 1 10 9 7 1 12 9 1 9 0 7 13 3 1 10 9 1 9 2
15 15 13 16 10 9 1 11 4 13 1 10 9 16 13 2
46 10 9 1 9 11 13 3 10 12 1 12 1 10 9 1 9 1 11 2 1 10 12 9 2 1 10 0 9 1 9 3 1 16 10 11 13 10 9 1 9 13 10 9 1 9 2
31 10 0 9 1 9 7 9 13 10 9 1 2 10 11 8 11 10 11 2 2 1 10 15 10 9 1 11 13 9 0 2
33 1 10 0 9 15 13 10 11 11 1 10 11 11 1 10 11 11 1 10 11 11 2 16 13 9 1 11 1 9 7 9 0 2
17 7 13 10 9 2 10 9 15 13 2 7 3 13 12 1 12 2
20 10 9 13 1 10 9 1 10 9 0 1 13 10 9 0 13 1 10 9 2
31 1 0 9 1 10 9 0 0 3 13 1 9 1 10 9 0 1 11 2 13 0 13 9 0 1 10 9 1 10 9 2
20 1 10 0 9 2 10 11 13 10 0 9 1 10 11 7 10 11 11 11 2
28 15 9 3 15 13 1 13 9 0 16 13 9 1 10 9 0 2 7 13 13 9 16 13 3 7 3 0 2
20 10 9 13 2 0 2 4 7 13 15 1 9 1 9 16 13 15 3 0 2
63 1 10 9 2 13 10 9 10 16 13 1 2 10 9 1 9 2 9 1 9 2 9 2 9 2 9 2 1 10 9 2 13 8 2 9 1 9 0 2 2 13 9 0 2 2 7 2 16 10 9 13 10 9 15 15 4 7 13 15 13 9 2 2
41 1 10 0 9 10 11 13 13 10 9 1 15 3 9 16 13 13 10 10 9 7 13 10 9 1 8 8 2 16 3 15 13 1 10 9 2 10 9 1 12 2
34 16 11 13 1 10 11 2 3 13 1 10 9 0 8 8 8 2 11 2 1 9 1 10 9 8 8 1 10 9 11 7 11 11 2
17 11 4 13 1 10 9 1 10 11 2 1 10 0 9 1 12 2
20 3 1 9 15 13 1 9 2 15 3 7 3 1 10 9 7 13 9 0 2
32 10 9 1 10 9 13 1 11 2 1 10 0 9 1 10 9 1 11 1 10 11 2 3 15 13 1 12 7 13 1 12 2
31 1 10 9 2 10 9 13 9 1 10 9 11 7 13 1 9 1 10 9 1 11 7 1 10 9 1 10 9 0 0 2
32 15 13 16 10 9 0 13 10 9 16 13 10 9 0 1 10 11 11 1 10 9 1 11 2 13 10 12 1 11 1 12 2
12 10 9 1 9 0 7 9 0 15 4 13 2
16 1 10 9 1 9 1 9 0 2 10 9 13 13 9 0 2
38 10 9 0 1 10 11 12 13 3 1 10 9 1 9 0 2 11 11 11 11 2 1 9 1 9 1 9 16 3 15 13 1 9 1 4 13 15 2
19 10 9 13 10 9 1 10 9 0 2 16 13 13 3 1 10 9 0 2
10 10 0 9 13 12 9 7 12 9 2
29 1 12 2 3 1 0 9 7 9 0 2 13 10 11 11 1 9 1 10 12 9 1 10 9 1 9 7 9 2
18 10 9 13 10 9 0 1 5 12 9 1 10 5 12 1 10 9 2
20 3 3 4 4 13 0 7 3 4 4 13 1 10 9 1 0 9 1 11 2
20 1 10 9 13 10 12 1 11 2 11 13 16 4 13 13 15 1 0 9 2
32 1 12 13 10 9 1 10 9 1 11 1 3 13 1 13 10 9 1 9 1 10 9 2 10 11 2 2 5 2 5 2 2
18 4 13 9 2 9 2 9 0 7 0 2 7 9 1 9 7 9 2
19 10 9 13 9 3 0 16 13 1 10 9 0 1 9 1 9 7 9 2
25 3 1 10 9 0 1 11 2 9 2 10 9 15 13 1 10 9 1 10 9 0 1 10 9 2
27 15 7 10 9 4 13 1 11 11 2 10 0 9 16 13 15 3 16 10 9 1 10 9 1 10 9 2
7 1 10 9 15 15 13 9
26 13 3 0 9 1 10 9 1 13 10 9 2 10 13 10 9 3 0 7 1 10 9 15 13 9 2
59 10 15 13 9 2 7 1 9 3 13 1 10 9 1 10 9 2 1 9 1 13 10 9 1 10 9 3 0 7 4 13 9 7 13 1 9 2 9 16 3 13 15 1 1 1 15 2 7 1 9 13 1 9 7 3 1 9 0 2
39 11 15 13 10 9 1 9 7 9 2 7 3 2 15 13 10 9 9 13 1 9 1 11 2 11 11 2 2 9 7 9 1 10 11 1 16 13 11 2
37 16 13 1 10 9 1 11 11 11 11 11 11 2 11 13 16 10 9 1 10 9 13 10 0 9 2 13 10 9 7 2 10 11 1 11 2 2
10 10 9 13 0 1 10 9 1 12 2
20 10 9 1 10 9 8 7 8 15 13 10 9 1 9 9 1 15 3 9 2
24 13 15 1 10 9 1 10 9 1 9 7 9 13 13 3 9 2 9 7 9 1 9 0 2
21 13 10 9 1 12 9 16 13 10 11 1 11 12 2 16 3 13 9 1 9 2
43 1 10 12 9 1 10 9 2 1 12 13 2 2 11 11 13 9 1 12 9 2 11 1 12 2 11 1 12 2 7 11 1 10 11 2 11 7 11 2 15 10 15 2
43 12 1 10 9 1 11 2 8 7 8 2 2 13 1 12 9 1 9 1 10 11 2 4 13 0 7 1 15 13 9 1 9 1 13 10 9 0 1 9 1 10 11 2
19 13 3 1 9 0 2 9 11 2 9 1 9 1 9 7 9 1 11 2
31 1 10 9 2 13 3 3 7 12 9 1 9 0 2 13 9 2 9 2 9 1 9 2 9 2 9 7 0 9 0 2
31 11 15 4 13 1 10 9 1 13 15 1 9 7 3 4 13 3 10 9 1 10 9 1 9 0 7 3 0 7 0 2
20 15 13 1 11 2 11 11 2 11 7 11 1 10 9 1 10 9 3 0 2
44 10 9 1 10 15 10 9 13 10 9 1 10 9 13 0 7 10 9 3 0 1 10 15 15 13 10 9 1 10 9 7 10 9 1 10 9 13 0 2 16 13 1 9 2
25 10 9 13 1 10 9 1 10 9 1 10 9 0 2 7 13 10 9 1 10 9 1 10 9 2
50 13 9 1 10 9 0 11 2 11 13 1 11 1 9 1 10 9 1 12 2 16 13 0 1 11 1 4 13 1 9 7 9 1 11 11 2 0 9 0 7 3 9 1 10 9 1 9 0 11 2
56 11 16 11 13 2 1 10 9 2 10 9 1 10 9 9 7 2 1 9 2 1 10 9 2 3 16 13 10 9 1 10 9 16 13 0 1 13 10 9 1 10 9 1 13 1 10 9 0 2 7 1 9 1 13 3 2
23 1 9 2 10 9 13 10 9 1 10 9 7 10 10 9 1 10 15 15 13 10 9 2
15 10 9 1 9 0 13 11 11 7 1 11 2 11 11 2
11 11 13 10 9 1 10 11 11 2 11 2
12 4 13 3 1 9 1 10 9 0 11 11 2
11 10 9 11 13 10 9 1 9 1 9 2
16 13 10 9 0 7 10 9 1 10 9 0 1 10 0 9 2
30 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 1 10 11 2
7 10 9 13 1 9 0 2
29 15 13 10 9 0 2 15 13 1 9 0 2 13 1 10 9 11 11 7 15 13 1 9 13 1 10 9 0 2
30 10 11 13 10 9 0 1 10 9 2 13 1 10 9 1 10 15 13 9 1 10 9 1 0 9 1 10 11 11 2
18 10 9 0 4 13 1 10 9 0 1 10 9 0 7 9 11 11 2
39 13 16 10 9 0 13 3 10 9 1 9 7 10 0 9 1 10 9 7 16 10 9 13 3 13 3 1 10 9 7 13 1 9 1 9 1 10 9 2
4 13 3 0 2
34 3 13 10 0 9 1 9 0 1 10 0 9 2 11 2 1 10 16 15 4 13 10 9 2 1 10 10 9 2 1 10 9 0 2
31 1 12 13 10 9 1 9 1 9 1 10 9 1 11 7 1 10 9 8 13 1 10 9 1 10 9 1 11 7 11 2
38 10 9 15 13 16 13 1 10 9 11 11 7 15 1 10 9 2 9 1 10 9 1 10 9 0 2 13 1 10 9 1 10 9 2 11 11 11 2
59 1 10 12 9 2 11 13 0 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
12 1 3 1 12 9 15 15 13 10 9 0 2
31 10 9 3 13 0 1 10 9 2 3 16 13 9 1 0 9 1 9 7 9 0 13 1 10 9 0 7 1 15 0 2
32 3 1 16 10 9 4 13 1 10 9 12 7 10 12 2 10 9 13 1 9 1 10 9 7 13 10 9 1 9 1 9 2
46 11 11 11 2 9 0 1 11 2 13 16 10 9 13 9 1 10 9 1 10 9 1 9 1 9 1 9 0 7 9 1 9 7 3 16 10 9 15 13 1 9 1 9 7 9 2
37 11 11 1 11 13 16 10 9 2 13 0 1 9 1 10 9 1 10 9 2 7 13 10 9 2 1 10 9 1 9 3 0 1 0 9 2 2
38 2 13 10 9 1 15 1 11 2 13 1 10 9 2 16 13 10 9 1 10 9 2 1 10 9 0 7 9 1 11 2 2 13 10 8 9 0 2
33 13 10 9 10 16 13 1 10 9 1 12 9 2 15 1 11 2 16 13 10 0 11 2 7 15 1 11 2 16 13 1 11 2
25 1 10 9 1 10 9 2 0 2 13 3 10 9 1 10 9 7 10 9 1 10 9 1 9 2
23 1 15 3 15 13 15 0 7 3 4 1 13 16 15 13 3 7 13 9 3 1 13 2
5 4 13 1 12 2
12 10 9 13 10 9 2 1 15 9 1 11 2
34 10 9 4 13 1 10 9 11 11 15 4 13 1 9 1 10 9 16 2 1 9 3 13 9 2 7 1 9 3 4 13 9 2 2
6 1 12 13 1 11 2
52 10 9 1 10 9 0 15 13 1 10 12 1 12 1 10 9 7 10 9 2 1 10 16 3 13 12 9 0 1 9 1 9 7 9 2 3 7 10 9 0 7 2 9 2 16 15 13 1 10 9 13 2
25 13 1 10 9 1 16 10 9 13 9 0 7 2 1 1 15 2 13 1 10 9 1 0 9 2
7 10 9 13 1 10 9 2
39 1 9 1 10 9 1 10 9 2 1 10 9 13 1 11 2 15 4 13 1 10 9 1 10 9 1 10 9 2 9 16 13 15 3 1 12 9 13 2
45 11 11 11 11 11 2 13 1 0 10 11 1 11 7 10 11 11 11 1 11 2 13 10 9 0 13 10 12 1 11 1 12 1 11 11 7 10 12 1 11 1 12 1 11 2
32 1 0 9 2 13 10 9 0 3 4 13 9 0 1 10 9 13 1 10 0 9 16 15 4 1 13 1 10 9 1 11 2
11 10 9 1 10 8 1 10 9 13 0 2
29 10 9 1 11 13 15 1 10 9 1 9 1 10 9 1 11 2 13 1 10 9 9 0 1 10 11 10 11 2
9 15 13 16 1 12 13 10 12 2
33 11 2 0 2 15 13 16 3 13 13 15 3 3 2 7 11 2 13 15 2 13 1 11 16 13 15 16 13 9 1 10 9 2
20 10 9 0 13 1 11 1 12 9 1 9 1 11 7 1 10 12 9 13 2
43 2 10 9 13 16 3 13 0 10 12 9 1 9 16 13 16 13 13 10 9 0 7 16 2 3 2 13 16 13 10 9 7 0 1 13 2 2 13 10 9 1 11 2
14 11 2 9 2 11 10 11 13 10 9 0 1 12 2
42 10 9 0 13 10 9 1 9 0 1 12 1 12 9 1 12 5 8 13 1 10 9 0 7 9 1 9 2 9 2 9 2 1 7 1 10 9 1 9 0 2 2
42 10 12 1 11 1 12 2 10 9 13 10 9 1 10 9 12 1 10 11 11 11 3 13 10 3 0 9 0 1 10 9 2 7 1 10 9 12 1 10 9 0 2
19 13 1 10 8 13 1 10 9 7 11 13 1 10 9 10 9 1 3 2
20 10 9 13 3 16 13 0 2 16 3 1 10 9 1 10 9 13 10 15 2
34 1 10 9 0 4 13 1 10 11 1 11 1 11 2 7 1 10 9 0 15 13 1 11 2 7 3 4 1 11 2 3 1 3 2
7 10 9 0 13 10 9 2
63 10 0 9 0 13 11 11 2 11 11 2 2 16 13 3 9 1 10 9 7 1 10 9 1 12 9 2 11 11 2 11 11 2 2 13 10 9 1 9 7 10 9 4 1 13 1 9 7 13 10 9 1 10 10 9 1 10 9 0 1 10 9 2
35 10 9 0 2 16 15 4 13 1 13 10 9 2 13 1 9 0 1 10 9 13 3 10 9 1 9 7 10 9 1 9 16 11 13 2
21 15 16 15 13 4 13 1 10 2 9 0 3 0 1 10 9 1 10 9 2 2
20 10 0 9 13 1 15 1 10 9 1 10 9 3 1 10 0 9 1 9 2
35 7 2 1 9 2 13 10 0 9 13 7 13 9 1 10 9 1 11 7 11 2 9 1 10 9 0 7 9 1 10 9 1 10 11 2
42 3 0 13 9 1 10 9 1 10 9 2 7 9 1 11 11 13 1 9 1 10 9 1 10 9 13 1 16 4 1 13 1 10 9 1 10 9 0 1 10 9 2
25 10 9 3 15 13 1 10 0 9 1 11 11 2 13 10 9 12 1 10 11 11 12 1 12 2
23 10 9 15 13 1 9 7 10 9 0 13 3 2 15 7 4 13 15 1 10 0 9 2
12 10 9 1 9 1 10 9 13 1 9 12 2
29 1 10 9 1 12 10 9 1 9 1 11 13 1 12 13 1 12 7 1 12 4 1 13 13 1 12 1 12 2
38 13 10 9 0 7 1 9 0 2 10 9 0 2 3 1 9 2 10 9 1 9 1 13 10 10 9 7 10 9 0 1 9 7 9 1 10 9 2
26 10 2 9 0 1 12 9 2 15 13 1 10 9 7 15 13 1 15 1 10 9 0 1 10 9 2
39 10 11 15 4 13 1 11 1 10 9 2 7 13 10 9 1 13 15 1 10 11 11 2 1 0 9 0 2 16 10 9 4 13 1 10 0 11 11 2
24 1 9 0 2 15 13 1 10 9 11 2 10 11 2 11 11 2 11 7 1 10 9 11 2
30 10 12 1 11 1 12 2 10 9 1 10 0 9 0 13 11 1 10 9 1 9 16 13 1 10 0 9 11 11 2
25 3 13 1 10 11 11 2 10 9 13 3 0 2 7 1 3 13 1 10 9 16 13 1 15 2
68 1 11 1 12 13 0 3 10 9 11 2 11 11 11 2 9 1 0 9 16 16 13 10 9 1 12 9 1 9 1 12 2 8 7 8 2 7 15 1 10 12 1 11 1 10 12 2 4 13 1 10 9 1 3 1 12 9 1 10 9 7 10 0 9 1 10 9 2
16 15 13 1 10 0 9 1 10 9 1 10 9 11 7 11 2
56 11 11 11 2 11 11 11 13 10 9 1 10 9 11 11 11 7 13 12 9 0 2 12 9 0 7 12 9 0 3 0 2 3 1 0 9 7 9 1 10 9 0 2 10 9 13 1 10 0 9 3 0 2 10 9 2
27 11 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 11 11 2 2 13 10 9 7 9 0 2
21 2 10 9 13 16 10 9 13 10 9 1 10 9 4 13 10 9 1 10 9 2
23 1 10 9 15 13 1 9 11 11 1 10 9 7 11 11 2 11 11 2 1 10 9 2
37 4 13 1 10 9 0 1 10 9 11 2 16 13 1 10 11 11 2 12 9 1 10 9 1 10 9 1 11 7 12 9 1 10 9 1 11 2
63 15 13 1 0 9 13 1 10 9 3 13 2 1 10 9 1 10 9 2 1 10 9 1 10 9 1 10 11 2 2 15 1 10 11 2 1 11 11 2 1 10 9 1 11 2 10 9 7 9 2 1 10 9 0 2 7 10 9 2 1 11 2 2
28 15 13 16 13 3 12 9 2 9 0 2 9 9 0 2 12 9 1 9 2 9 0 0 13 1 10 9 2
29 10 9 13 1 9 1 10 9 11 2 1 13 10 9 1 10 9 1 9 4 13 3 9 1 9 1 10 9 2
9 1 10 9 11 11 13 12 9 2
26 1 9 1 16 10 9 1 9 11 13 3 0 2 10 9 1 9 11 13 10 9 1 9 3 0 2
14 3 13 0 2 3 13 9 7 15 13 3 1 13 2
56 11 2 11 7 11 2 11 2 9 1 11 11 2 11 1 11 1 11 11 2 11 7 11 2 13 10 0 9 3 0 1 11 7 11 2 16 1 10 9 0 1 0 9 2 16 13 10 0 9 1 9 0 1 10 9 2
43 13 1 10 9 1 10 9 1 11 2 1 2 11 2 1 10 9 1 9 2 1 10 9 7 1 10 9 1 9 2 1 10 9 1 10 11 11 7 1 11 1 11 2
32 10 0 9 1 11 11 1 10 11 4 13 16 12 9 0 13 10 9 1 10 9 3 0 7 16 13 1 10 9 1 9 2
43 10 9 12 2 3 1 10 9 0 2 15 13 3 1 10 12 0 9 1 11 2 15 15 13 1 10 0 9 1 9 16 15 13 1 11 2 1 10 11 11 1 11 2
21 11 12 4 13 10 12 1 11 1 10 12 1 10 11 11 1 10 11 2 11 2
48 10 9 2 10 9 0 11 11 2 13 10 9 1 12 2 1 10 15 13 1 12 2 1 10 15 13 1 10 0 9 1 9 0 3 1 10 9 0 1 10 9 2 16 3 1 10 9 2
12 15 15 13 1 0 1 10 9 1 10 9 2
24 10 0 9 2 1 11 2 11 11 2 13 10 9 2 10 11 2 2 1 10 9 11 11 2
19 1 12 2 11 11 4 13 9 1 10 9 1 10 9 1 13 10 9 2
11 11 11 1 10 11 7 10 11 2 11 2
12 3 16 13 10 9 4 13 9 0 1 9 2
10 10 0 9 1 10 9 13 10 9 2
35 13 10 0 9 1 11 1 13 1 10 11 12 0 2 13 1 10 9 9 12 2 7 10 9 13 1 10 9 12 1 10 9 1 9 2
27 10 9 3 15 15 13 10 9 0 7 0 2 1 10 15 13 13 10 10 9 7 10 0 9 1 11 2
34 10 9 0 13 10 9 1 9 7 9 2 7 13 10 9 7 9 16 15 13 1 10 9 1 10 9 0 1 10 9 1 10 9 2
41 9 1 10 9 0 1 11 2 9 1 10 9 1 10 9 2 13 16 13 3 10 9 2 1 0 10 9 1 9 1 9 2 16 13 1 10 9 1 10 9 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 9 2
50 10 0 9 1 10 8 0 15 13 10 9 0 2 1 10 16 15 4 13 1 0 9 0 2 7 16 1 10 9 13 15 1 10 3 0 1 11 13 1 10 0 9 1 10 9 9 1 10 9 2
14 9 1 9 1 10 1 9 1 12 9 0 1 9 2
26 13 10 12 1 11 1 12 2 15 3 1 13 12 9 2 1 9 1 9 13 1 10 9 1 11 2
25 10 9 13 13 10 9 1 9 16 13 1 10 9 13 15 3 1 10 9 1 9 1 10 9 2
9 11 11 11 13 1 10 9 0 2
58 10 9 1 10 11 13 10 11 1 11 11 1 11 10 9 1 9 0 2 10 11 1 9 12 2 1 10 9 2 11 10 11 3 2 3 15 13 15 2 7 16 13 1 9 13 3 1 12 9 1 10 9 2 13 10 9 0 2
24 4 13 10 9 1 9 2 7 10 9 13 16 13 15 3 2 13 3 0 9 1 10 9 2
31 10 9 1 10 15 10 9 15 13 1 9 7 15 15 13 1 10 9 1 9 7 1 10 0 9 1 11 10 0 9 2
10 3 3 4 13 1 10 9 1 11 2
15 13 0 1 10 9 7 1 10 9 7 15 9 13 9 2
63 10 9 1 9 0 13 1 10 12 5 1 10 9 2 7 16 10 12 5 4 13 1 11 2 10 12 5 1 11 2 10 12 5 1 11 1 10 11 2 10 12 5 1 11 1 10 11 2 10 12 5 1 11 2 7 10 12 5 1 10 10 9 2
76 10 9 3 13 1 10 9 2 15 1 10 9 4 13 2 10 11 2 1 10 9 16 13 1 10 9 1 10 9 16 15 13 2 13 1 16 13 10 9 13 10 9 1 10 9 1 0 9 2 16 3 13 10 15 13 10 9 11 7 11 2 15 15 4 13 10 9 0 1 10 0 9 1 0 9 2
13 11 4 13 10 9 1 10 9 1 9 8 8 2
26 3 2 10 9 13 1 9 1 7 13 10 9 1 10 9 1 10 9 1 16 15 4 13 1 11 2
32 9 2 10 9 13 0 7 15 13 0 2 7 2 16 8 13 0 2 8 13 10 9 0 2 10 15 13 16 8 13 0 2
12 16 13 13 1 9 13 1 10 9 1 9 2
16 1 9 10 9 15 13 13 1 10 9 1 12 1 12 9 2
17 11 11 4 13 1 2 8 2 11 11 11 7 13 1 11 11 2
10 4 13 9 0 1 11 7 1 11 2
13 16 15 13 15 13 1 13 15 16 3 4 13 2
47 15 13 1 10 9 2 15 13 10 0 9 2 15 13 1 13 15 15 16 4 1 13 7 10 9 16 13 1 10 9 2 10 9 16 13 3 1 10 9 1 15 13 15 1 10 9 2
23 10 9 4 13 1 10 3 12 9 3 1 10 0 9 2 10 0 13 10 1 11 2 2
35 16 15 13 1 10 9 2 13 10 0 9 1 11 2 10 9 11 11 2 10 9 16 15 13 1 13 1 10 9 11 1 10 9 0 2
20 10 9 1 11 13 3 10 9 16 1 10 9 1 10 15 13 0 10 9 2
34 10 9 1 9 4 13 2 10 9 4 13 15 2 10 9 1 9 1 10 9 15 13 2 7 10 9 4 13 1 10 0 11 11 2
21 10 9 15 13 1 9 2 10 9 13 10 9 1 10 9 2 16 4 13 0 2
29 3 16 13 0 1 13 12 8 2 8 2 7 13 15 1 13 10 9 0 1 10 9 1 10 9 1 10 11 2
30 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 1 10 11 2
25 13 9 1 10 11 11 1 11 7 11 11 1 15 1 12 7 12 7 3 1 10 12 7 12 2
13 10 9 4 13 1 11 11 2 11 7 11 11 2
10 4 13 1 10 9 1 9 1 9 2
7 10 9 4 13 7 13 2
30 10 9 15 4 13 10 9 1 13 10 0 9 1 11 10 9 12 1 11 1 12 3 2 1 10 11 10 11 11 2
25 15 1 10 9 1 10 9 1 10 11 11 2 1 10 9 16 13 1 10 9 7 1 10 9 2
100 3 13 0 1 10 9 12 9 2 11 2 11 2 11 11 2 11 2 11 7 11 11 2 16 13 1 10 9 13 10 0 9 1 10 9 0 0 2 7 11 11 2 16 13 1 10 9 0 2 16 13 9 1 10 10 9 1 10 9 2 10 9 11 2 10 9 0 11 2 10 9 0 11 2 10 9 1 9 1 9 11 7 11 2 1 10 9 0 0 1 11 11 2 2 7 10 9 9 11 2
46 10 9 0 2 1 10 9 2 13 1 10 9 1 12 9 1 13 2 1 12 9 0 1 9 7 3 3 0 1 10 9 1 10 11 1 11 2 16 13 10 9 13 1 10 9 2
67 11 11 2 1 10 9 2 4 13 16 2 1 10 0 9 1 9 0 2 15 4 13 10 9 1 9 7 9 1 10 9 1 9 2 7 2 16 4 13 2 2 15 4 13 1 10 9 1 10 9 0 1 10 9 2 3 1 10 9 1 10 9 1 10 9 2 2
14 1 10 9 1 12 2 13 12 9 13 1 11 11 2
14 1 9 13 10 9 0 1 10 16 15 13 3 3 2
42 10 9 3 13 13 11 2 9 2 9 2 9 7 9 2 2 11 2 9 7 9 2 2 11 2 9 2 9 7 9 2 2 11 2 9 2 7 11 2 9 2 2
32 1 10 9 0 12 2 10 9 0 11 11 13 1 11 11 12 2 10 9 16 13 13 10 9 0 1 0 7 8 9 0 2
61 10 9 3 0 13 10 9 15 10 9 15 13 13 3 1 10 9 2 13 1 9 2 15 4 13 1 15 1 10 11 11 1 10 11 11 1 10 9 1 16 10 9 15 13 3 1 9 1 13 15 1 0 9 2 7 10 0 9 1 11 2
23 13 10 0 9 1 10 9 1 10 9 2 7 10 9 3 0 1 10 9 1 10 11 2
34 4 13 15 1 9 16 10 9 1 9 2 10 9 0 2 10 9 7 10 9 0 4 13 1 10 9 7 15 15 13 1 10 9 2
11 1 10 0 9 13 11 9 1 11 11 2
41 3 2 10 9 0 13 10 9 16 4 13 10 9 0 7 10 9 1 16 1 3 3 12 9 15 4 13 13 3 1 12 9 2 16 10 9 13 13 1 12 2
22 3 15 13 1 12 1 10 9 1 10 9 13 1 10 9 1 10 0 9 1 11 2
8 11 15 13 0 1 10 9 2
88 1 10 9 10 10 9 13 2 13 0 10 9 2 9 2 9 1 9 2 9 0 7 9 2 0 7 0 2 1 10 9 1 10 9 2 1 10 9 7 9 2 1 0 2 0 7 0 9 2 13 2 1 9 2 10 0 9 7 2 7 9 1 9 1 9 2 9 7 9 1 9 1 9 0 7 3 7 3 9 2 1 10 16 15 13 9 0 2
11 13 8 0 7 13 10 0 9 7 9 2
3 11 11 2
27 1 12 10 9 1 9 15 13 1 12 1 12 1 9 1 10 9 1 11 7 11 1 9 1 10 11 2
43 10 12 1 11 1 12 13 1 11 11 2 13 10 0 9 1 10 11 11 1 3 2 13 12 9 2 12 9 2 12 9 2 12 9 1 9 7 12 9 1 12 9 2
47 10 9 2 10 9 13 10 9 2 13 1 10 9 1 9 12 9 2 3 10 9 1 10 9 13 1 10 9 1 9 1 10 9 2 1 9 2 12 9 2 12 9 2 12 9 2 2
43 10 9 2 1 9 2 13 10 9 1 9 0 2 16 13 2 2 12 9 2 2 16 13 10 9 0 16 15 13 3 1 9 0 7 0 1 10 9 1 10 9 0 2
37 10 9 1 9 0 0 4 13 2 1 10 9 1 9 2 1 12 2 10 9 1 12 9 13 1 10 9 0 2 12 1 15 9 1 9 0 2
44 16 4 1 13 10 9 2 13 16 13 13 10 9 2 7 1 10 9 7 10 9 1 10 9 2 1 10 13 10 9 2 11 13 10 11 11 7 13 15 13 15 16 13 2
31 9 1 10 9 2 15 13 1 9 1 10 11 11 11 1 10 11 1 11 7 3 1 10 11 11 1 10 11 1 11 2
65 1 0 2 1 10 9 13 1 11 11 1 10 11 11 1 11 2 11 2 2 1 11 9 10 9 13 0 1 10 11 2 12 1 10 9 12 7 12 1 10 9 1 9 1 11 2 3 1 10 11 2 12 10 9 15 4 13 0 1 10 9 12 7 12 2
11 10 9 4 4 13 1 9 1 9 0 2
11 10 9 0 1 10 9 0 3 15 13 2
29 1 10 9 0 4 13 11 11 2 10 9 1 11 7 11 7 10 9 7 9 2 1 9 1 10 0 9 0 2
13 3 1 15 4 13 9 0 1 10 9 1 9 2
20 15 13 1 10 9 0 1 11 1 10 12 9 1 10 9 2 13 3 0 2
25 13 0 7 4 1 13 1 10 9 3 7 13 10 9 1 9 2 7 3 15 13 1 10 9 2
29 10 9 13 10 9 1 9 2 1 13 1 10 9 0 15 13 12 9 0 10 9 0 13 10 9 7 10 9 2
12 1 9 4 13 10 10 9 16 13 3 0 2
34 3 11 15 13 16 10 9 1 11 11 1 11 15 13 1 11 2 10 11 2 11 11 1 11 2 7 13 1 10 9 1 10 9 2
26 11 11 13 1 11 3 1 9 1 13 1 10 9 16 13 1 10 9 0 16 13 1 11 7 11 2
15 0 9 1 10 9 0 2 0 1 9 0 7 1 9 2
61 3 1 10 9 2 11 4 7 13 1 10 9 1 0 13 11 11 2 9 1 10 15 4 13 1 10 11 11 2 3 1 13 15 10 15 1 10 15 15 13 1 0 9 3 16 11 13 10 9 1 9 1 10 9 11 11 2 9 1 11 2
23 3 3 13 1 10 9 7 15 9 16 13 13 13 1 10 9 1 10 9 1 10 9 2
32 3 3 13 1 9 1 10 9 2 1 10 9 1 9 2 9 7 11 2 12 2 7 10 9 1 10 0 9 1 10 9 2
36 10 9 0 1 11 2 13 9 1 9 0 1 10 11 1 11 2 15 13 13 1 12 9 2 13 1 10 9 11 2 10 11 7 10 11 2
10 1 10 9 2 15 13 16 13 0 2
30 15 13 10 9 1 10 15 15 13 1 10 9 1 10 9 1 10 9 3 10 9 8 10 9 1 16 13 0 9 2
24 11 11 11 2 11 1 10 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 0 2
23 10 9 2 11 2 3 0 7 0 1 10 9 1 9 7 9 13 0 7 0 7 0 2
18 10 9 0 0 2 10 9 1 9 7 9 2 2 2 10 0 9 2
32 13 1 10 9 1 11 2 11 13 1 10 9 0 1 11 2 11 2 11 2 11 7 11 1 11 2 3 7 11 1 11 2
24 10 9 13 3 1 11 11 12 2 3 1 11 2 1 9 1 11 11 11 0 1 11 11 2
30 9 3 10 9 1 10 11 13 9 0 1 9 2 9 1 9 0 7 10 10 9 16 10 9 1 9 0 4 13 2
43 3 1 16 10 9 13 10 11 11 1 12 9 1 11 2 10 0 9 4 13 2 10 9 15 13 10 9 11 1 13 12 9 11 1 11 1 10 11 1 9 0 11 2
28 10 9 13 10 11 1 10 9 11 2 1 10 9 11 4 13 10 9 1 11 0 2 13 15 3 1 11 2
7 4 13 1 12 12 8 2
79 1 13 10 9 2 11 13 10 9 1 11 11 2 11 2 10 9 1 9 13 1 11 11 2 1 10 9 1 13 9 0 7 9 1 9 2 13 9 1 9 0 2 13 9 0 1 0 9 1 10 9 2 13 9 1 9 2 7 13 1 9 0 1 9 1 11 11 11 2 11 2 11 2 11 11 2 7 11 2
36 10 9 13 10 0 9 0 7 1 15 2 10 9 1 9 8 2 11 10 11 2 2 13 3 13 1 10 9 0 1 10 9 1 10 9 2
16 11 7 11 13 1 9 10 9 2 11 11 11 11 11 2 2
17 9 1 10 9 0 2 3 3 10 9 0 7 10 9 0 0 2
32 10 12 1 11 1 12 13 10 9 1 11 11 2 3 13 1 10 9 1 10 9 2 15 15 13 3 3 16 13 10 9 2
15 1 12 4 13 1 10 11 1 11 1 0 9 1 9 2
12 3 15 13 10 9 13 1 10 9 1 11 2
66 10 9 3 13 1 10 9 1 2 11 7 11 11 1 10 11 2 2 0 2 8 8 2 2 3 4 13 15 1 10 2 0 9 1 10 9 2 2 9 2 8 8 2 2 10 9 1 10 9 11 1 10 9 0 1 10 11 11 2 3 1 11 2 1 11 2
24 13 9 2 7 13 9 2 13 10 9 0 16 13 1 13 9 1 9 16 13 10 9 0 2
31 4 13 1 10 9 11 1 11 8 11 2 15 2 11 1 12 1 13 1 10 9 13 1 10 9 13 1 9 1 9 2
12 10 9 1 9 13 1 12 9 2 9 5 2
17 13 1 9 7 10 0 9 13 10 11 11 11 1 10 11 11 2
32 10 11 13 10 9 1 9 0 1 9 0 2 1 10 15 15 8 9 1 10 9 13 9 0 2 15 1 9 0 1 9 2
23 13 1 11 1 12 7 15 13 1 11 1 11 2 13 0 9 0 1 10 9 1 9 2
35 1 15 16 15 13 13 1 13 9 1 10 9 2 15 16 15 13 1 10 9 1 15 15 15 13 13 7 10 9 13 1 13 10 9 2
37 3 10 9 7 10 9 4 4 13 1 10 0 9 1 9 0 7 1 9 13 1 9 0 1 9 1 10 9 0 8 9 1 10 3 9 0 2
13 13 1 10 9 1 10 9 7 15 13 3 3 2
33 11 11 2 11 2 12 2 12 2 13 1 11 2 7 3 4 13 10 12 5 1 10 11 1 11 2 7 13 3 12 9 3 2
19 10 9 1 9 15 13 10 9 1 11 1 10 12 9 1 10 0 9 2
15 3 1 13 2 11 15 13 1 11 16 3 13 13 15 2
15 10 9 7 10 9 4 13 2 10 9 4 13 10 9 2
20 13 3 0 16 1 15 3 15 13 15 1 13 7 4 13 9 7 9 13 2
15 3 3 13 0 10 9 2 10 9 13 1 10 9 13 2
20 13 0 2 13 1 10 9 1 11 7 15 4 13 10 9 1 7 1 9 2
8 10 9 1 10 9 13 11 2
80 13 1 10 9 1 0 9 2 15 1 10 3 0 13 15 13 11 1 11 10 9 11 11 4 13 1 13 9 0 1 10 9 7 1 10 9 0 2 9 15 10 9 11 13 3 2 13 16 10 9 4 4 13 1 10 8 2 9 2 13 3 13 1 9 0 0 2 3 3 2 10 9 1 10 9 1 10 9 13 2
13 11 13 10 9 1 10 11 11 1 11 2 11 2
41 11 13 10 9 0 1 9 7 9 1 9 0 1 12 9 0 2 11 11 2 13 10 12 1 11 1 12 2 7 11 11 2 13 10 12 1 11 1 12 2 2
34 9 13 10 9 0 1 13 10 9 0 2 15 13 10 9 10 9 7 10 9 7 10 9 16 13 0 2 7 16 13 15 15 0 2
30 10 9 0 1 10 9 1 8 2 9 13 12 7 12 9 2 10 9 2 10 9 7 9 2 10 9 7 10 9 2
28 15 13 1 10 9 2 9 16 10 11 1 11 11 4 13 1 10 0 9 16 3 13 10 9 1 12 9 2
24 11 11 7 11 2 0 9 1 10 9 2 13 0 7 3 0 2 12 1 11 1 12 2 2
7 13 12 9 1 10 9 2
39 13 16 13 13 8 1 11 2 13 1 13 9 5 9 1 11 7 10 9 13 10 9 13 4 13 10 9 3 0 1 10 9 1 9 1 10 16 13 2
74 3 13 0 10 9 1 13 3 7 10 9 16 13 10 9 3 13 9 1 9 1 9 0 7 9 7 9 1 9 16 15 13 13 2 13 10 9 1 10 9 7 3 15 13 16 10 9 1 9 16 15 4 1 13 15 4 13 1 10 9 1 9 0 1 9 0 7 15 15 4 13 1 0 2
29 1 11 4 13 1 10 11 1 11 7 10 11 2 10 0 13 10 9 4 4 13 1 10 9 1 10 9 11 2
9 10 9 1 10 9 3 15 13 2
36 10 9 13 0 1 9 0 16 15 13 13 1 10 9 7 13 1 10 9 1 10 9 1 9 1 10 9 1 10 9 0 1 11 7 11 2
29 11 11 11 2 12 1 11 1 12 2 13 10 9 1 9 7 0 9 2 3 13 1 4 13 1 10 9 11 2
21 11 13 10 9 1 9 1 9 0 0 0 1 11 2 3 13 1 10 9 11 2
28 16 13 11 2 11 2 11 7 3 11 2 10 9 15 4 13 1 0 1 11 11 2 10 9 13 10 9 2
43 1 13 16 10 9 0 3 0 16 13 0 2 10 9 4 13 1 10 9 1 9 1 9 2 16 1 10 11 11 2 12 13 10 0 9 16 13 10 9 1 0 9 2
23 10 12 9 7 12 9 3 13 1 10 9 1 11 2 11 8 2 1 10 9 1 11 2
6 10 12 9 13 0 2
40 1 10 9 4 13 1 10 9 11 1 11 16 13 10 9 0 1 11 11 1 11 2 13 16 15 13 13 15 7 13 1 9 13 10 9 1 10 0 9 2
19 9 1 9 7 11 11 7 15 1 11 11 11 11 7 11 3 13 9 2
15 9 1 10 9 2 10 9 4 13 15 1 10 9 0 2
13 1 10 9 15 13 10 9 1 10 9 1 9 2
29 10 9 1 10 9 1 11 2 10 12 5 2 13 1 3 1 12 9 7 3 10 12 5 13 1 3 1 12 2
62 10 9 13 1 9 2 11 11 2 11 11 1 11 2 11 11 2 11 1 11 2 11 11 2 11 1 11 2 11 11 7 11 2 11 11 2 11 11 1 11 2 11 11 11 2 11 11 7 11 2 11 11 11 2 11 11 11 2 7 11 11 2
33 10 9 9 13 1 10 9 13 1 11 2 1 10 9 1 13 10 10 9 13 1 10 0 9 1 10 9 13 1 9 1 11 2
50 10 13 10 9 1 10 9 1 10 16 13 9 11 11 2 13 10 9 0 1 9 2 13 10 9 0 2 13 1 10 10 9 0 7 13 16 15 13 10 9 0 13 1 10 9 0 2 2 13 2
38 1 10 9 0 10 9 4 13 1 15 1 10 9 0 7 11 2 1 9 2 2 15 9 1 10 0 9 2 7 2 15 9 1 10 9 2 2 2
28 3 2 10 9 1 9 0 0 2 13 1 11 11 2 4 13 10 2 11 11 2 2 13 10 9 1 9 2
45 11 11 13 10 9 0 1 9 1 11 2 11 2 11 11 13 9 0 1 11 7 10 11 1 11 1 10 11 11 2 10 11 1 10 11 7 11 2 1 10 9 1 12 9 2
16 11 11 13 10 9 1 9 1 10 9 11 1 10 9 11 2
46 11 13 16 10 9 13 1 10 2 9 0 7 0 2 1 10 9 0 2 7 16 3 15 13 1 10 2 9 0 1 9 13 1 10 9 0 2 13 1 10 9 1 10 9 0 2
37 4 13 1 12 2 13 15 1 10 0 9 1 4 13 1 10 9 3 1 2 11 11 10 11 2 2 2 11 2 7 2 11 11 10 11 2 2
36 10 9 1 10 9 2 1 10 9 8 10 9 3 13 0 2 1 15 15 13 0 13 0 9 16 13 1 13 1 10 9 10 9 3 0 2
12 10 9 9 0 1 10 9 13 1 12 9 2
46 15 16 1 9 13 7 13 13 9 0 1 13 1 9 1 0 9 3 7 3 15 13 1 10 9 1 9 1 9 16 13 11 7 1 10 9 1 13 9 0 1 9 1 13 9 2
35 11 11 1 11 11 13 1 10 9 12 9 1 12 7 13 2 2 1 10 0 9 0 2 11 3 13 10 9 0 2 7 15 13 0 2
13 10 9 1 9 13 1 12 8 2 2 9 8 2
41 1 9 2 1 9 1 13 15 15 1 10 9 0 3 0 1 10 11 1 11 2 3 4 4 13 1 9 0 2 0 2 16 1 10 9 15 4 13 1 15 2
20 10 0 9 13 11 1 10 11 11 1 11 7 11 2 12 9 1 10 11 2
17 1 9 2 10 9 15 13 10 0 9 7 15 13 9 1 11 2
15 13 10 12 1 11 7 13 1 10 9 1 12 1 11 2
16 1 10 9 1 10 9 2 15 13 10 9 7 10 9 0 2
26 15 13 1 10 0 9 0 13 1 13 10 9 16 13 10 9 1 13 10 9 0 1 11 7 11 2
20 1 10 9 15 13 3 0 10 9 1 10 9 3 1 10 9 1 10 9 2
8 3 3 13 10 9 1 11 2
22 3 11 3 13 15 1 0 9 2 7 1 10 11 7 10 11 2 1 12 11 11 2
44 7 13 12 1 12 1 11 1 10 9 16 13 1 10 9 1 10 11 2 7 3 1 11 11 3 1 12 1 12 2 13 1 10 0 9 1 10 0 9 1 9 1 11 2
41 11 11 2 1 11 2 13 10 9 9 1 11 1 10 1 10 9 11 11 2 13 15 1 10 9 1 10 9 0 1 10 9 2 7 15 13 12 1 12 9 2
32 10 9 13 0 7 0 10 0 9 1 10 9 7 10 9 1 10 9 1 10 9 13 0 2 13 9 3 1 9 1 9 2
19 11 2 1 9 2 11 2 13 10 9 1 11 2 1 10 9 1 11 2
21 10 9 0 4 13 13 12 9 1 10 9 0 1 11 2 11 2 1 9 0 2
20 1 10 11 0 15 13 3 0 9 2 9 2 9 2 9 0 1 10 9 2
34 11 2 11 2 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 2 11 7 9 1 11 2
25 10 9 13 10 0 7 0 9 1 10 15 15 13 10 9 1 10 9 1 9 1 13 10 9 2
18 15 4 13 9 1 10 11 1 10 11 16 13 9 1 10 11 11 2
30 11 11 13 9 1 9 1 11 1 10 13 10 0 9 1 11 11 11 1 13 12 9 1 10 9 9 1 10 9 2
48 1 9 1 10 11 1 11 2 11 2 11 13 1 9 10 9 1 10 9 0 7 10 9 1 10 9 0 2 16 9 7 9 1 10 0 9 2 2 1 10 15 3 13 1 9 1 9 2
16 10 9 0 1 11 13 16 10 0 9 15 13 1 11 0 2
16 1 10 9 1 11 2 9 1 11 2 13 10 9 1 15 2
25 10 9 0 13 10 9 1 10 9 1 15 13 1 10 9 1 10 9 1 9 7 9 1 12 2
21 1 10 9 1 11 1 11 1 12 2 10 11 11 12 15 13 1 11 1 11 2
19 1 9 1 0 9 15 4 13 9 7 9 16 13 9 3 1 10 11 2
12 10 0 9 1 10 16 4 13 1 10 9 2
35 10 9 0 2 0 7 0 16 1 10 9 4 13 11 7 11 7 3 13 13 15 1 11 2 1 10 9 1 9 16 13 1 10 9 2
16 3 13 1 11 7 10 11 1 16 13 1 11 2 11 2 2
16 4 13 1 10 0 11 1 11 2 1 10 9 1 10 11 2
18 15 13 3 1 9 2 9 9 2 15 10 9 13 9 1 10 15 2
36 1 10 9 0 1 10 9 11 15 13 10 9 1 10 9 11 11 2 9 1 10 9 11 1 11 11 2 15 13 10 9 2 9 10 9 2
23 1 10 11 11 11 2 15 13 1 9 9 7 9 0 2 13 10 9 0 1 0 9 2
33 15 13 1 15 1 10 9 2 13 9 2 9 2 7 9 2 9 2 2 16 15 13 1 15 9 1 10 9 7 1 10 9 2
38 3 4 1 13 15 0 16 13 16 13 1 10 9 13 15 16 4 7 13 2 16 3 15 13 3 4 1 13 2 16 13 10 10 9 1 10 9 2
27 3 11 1 11 13 1 10 11 11 1 11 7 10 11 1 11 11 1 10 9 1 10 9 11 11 11 2
18 10 9 13 10 0 9 0 1 10 9 0 7 13 1 10 9 0 2
23 10 0 9 1 9 4 13 9 1 10 9 2 10 15 4 3 13 1 10 9 0 0 2
17 10 9 13 1 0 9 7 1 10 9 16 13 3 13 10 9 2
29 15 1 10 9 3 0 1 10 9 13 10 9 1 10 9 1 9 2 9 16 3 13 10 0 9 9 2 9 2
16 11 15 13 7 4 1 13 11 1 11 2 13 15 2 11 2
25 13 0 10 9 1 10 0 9 1 10 9 1 11 2 11 11 7 10 11 2 10 15 13 0 2
26 10 9 11 12 1 9 7 11 4 13 1 9 1 11 1 11 2 11 1 10 9 11 12 1 11 2
29 10 9 1 9 1 11 7 10 9 0 7 10 0 9 1 10 10 9 13 11 3 7 10 10 9 1 11 11 2
17 10 9 0 13 10 11 10 0 9 1 10 11 1 10 9 11 2
15 10 9 1 10 9 13 3 13 3 1 12 9 1 9 2
14 15 13 1 15 1 16 10 9 0 13 15 16 13 2
25 13 9 1 10 9 2 12 9 2 13 10 9 1 10 9 0 7 10 9 0 2 1 9 2 2
20 11 13 1 10 9 15 15 13 1 9 2 1 10 9 0 1 11 11 11 2
30 3 3 2 10 9 1 11 1 11 2 11 11 2 13 1 10 11 1 3 4 13 0 9 1 10 9 1 10 9 2
23 3 10 15 13 1 9 1 9 7 9 2 9 1 9 7 9 1 10 11 11 7 9 2
41 1 10 9 1 11 2 11 13 9 9 1 10 11 2 13 1 10 9 1 11 7 13 9 1 10 9 11 11 2 11 2 2 9 1 10 11 2 8 12 2 2
18 12 9 3 3 13 1 11 2 3 13 12 9 2 7 1 13 9 0
47 8 13 1 12 5 9 1 12 2 10 9 11 11 11 2 15 13 13 2 7 10 9 1 10 9 13 0 1 15 16 15 4 13 9 1 10 9 1 12 9 7 12 9 1 10 9 2
57 9 15 3 4 13 2 7 8 8 1 10 9 3 0 2 1 13 10 9 2 1 9 1 9 1 11 11 11 2 11 11 2 11 2 11 11 2 11 2 11 8 15 16 1 10 0 12 9 4 13 0 1 10 9 10 9 2
24 10 9 13 10 9 0 13 1 10 9 13 16 4 13 3 1 10 9 1 9 7 13 3 2
20 12 2 10 11 0 1 9 1 9 1 11 3 2 10 12 1 11 1 12 2
26 3 10 12 9 15 13 1 13 16 10 9 13 1 10 9 16 10 0 9 13 16 13 0 1 13 2
18 13 1 10 9 11 7 10 9 11 1 10 9 1 9 0 1 11 2
13 15 13 9 1 13 7 1 8 0 7 0 0 2
16 13 1 10 9 1 11 2 15 13 1 10 9 1 10 11 2
19 1 11 13 1 11 2 3 11 9 0 13 13 1 11 16 13 10 9 2
11 1 10 9 2 9 1 9 7 10 9 2
10 15 15 13 7 13 13 15 1 15 2
16 15 15 13 13 12 9 7 15 13 1 10 9 1 10 11 2
32 3 13 9 1 10 9 0 2 7 3 10 0 9 1 10 9 2 10 15 4 4 13 3 1 10 9 0 1 10 9 0 2
34 1 9 2 11 12 13 10 9 1 10 9 1 10 9 1 11 11 1 10 9 1 9 2 1 9 10 9 3 0 1 10 9 0 2
11 13 10 0 9 1 10 9 1 9 0 2
50 10 0 9 1 12 9 2 11 2 11 2 12 2 2 13 1 9 1 11 11 2 11 4 4 13 1 10 9 1 11 11 11 2 11 2 11 2 12 2 1 10 0 9 1 10 0 9 1 12 2
20 9 1 9 0 15 4 13 1 10 9 1 9 11 2 3 1 10 9 11 2
13 11 13 1 9 0 2 15 13 1 10 9 1 13
29 1 10 9 2 13 1 10 9 0 1 10 9 16 10 0 9 0 13 13 9 0 1 10 9 3 0 7 0 2
11 10 9 13 16 10 9 13 15 16 13 2
23 13 10 9 1 9 0 16 15 4 13 1 13 1 10 9 16 15 13 1 10 9 0 2
20 3 10 9 1 13 1 10 11 1 11 13 9 3 0 7 15 13 0 9 2
9 10 9 0 13 9 1 9 0 2
9 1 9 2 11 13 10 9 13 2
30 1 3 1 10 9 2 13 10 9 2 1 8 9 2 7 13 0 2 10 9 1 9 1 9 7 9 3 0 3 2
10 1 10 9 13 10 9 1 10 9 2
21 16 13 9 7 13 10 9 0 2 9 2 9 2 9 2 2 2 13 10 9 2
82 15 15 13 3 1 12 9 2 10 9 1 10 9 13 1 10 9 1 10 9 0 2 11 11 1 11 11 2 11 11 2 8 2 13 1 16 13 13 10 9 1 10 9 1 11 7 10 9 1 10 9 0 2 16 13 13 10 9 16 15 13 3 0 1 10 9 2 1 10 9 0 2 0 7 0 2 13 7 13 1 11 2
27 11 11 11 13 10 9 0 16 13 10 0 9 1 9 0 2 12 9 2 12 9 2 1 10 9 0 2
42 10 9 2 16 4 13 12 9 1 9 1 9 1 9 2 9 7 9 2 3 4 13 3 4 13 11 2 16 1 11 7 1 11 2 10 8 16 13 9 2 13 2
12 11 0 13 10 9 1 9 1 10 9 11 2
13 13 3 10 9 0 3 1 10 9 1 10 9 2
31 1 10 9 2 10 0 9 13 10 9 1 0 9 0 2 7 13 2 1 9 2 10 9 1 10 9 7 1 10 9 2
28 3 1 10 9 7 1 10 9 0 2 13 0 9 11 7 11 16 15 13 3 7 15 13 3 1 10 9 2
27 1 10 9 2 10 9 0 15 4 3 13 1 9 7 9 2 16 13 1 11 7 1 11 2 10 11 2
18 1 9 2 1 9 1 10 9 13 3 0 1 9 1 10 11 0 2
31 1 10 9 2 10 9 1 10 9 2 1 10 9 2 1 10 1 9 2 2 10 9 7 10 9 13 3 1 10 9 2
13 1 12 10 9 1 10 11 15 13 1 12 5 2
9 15 13 15 16 3 15 13 8 2
61 1 10 9 13 1 10 11 1 10 11 1 10 11 11 1 10 12 1 10 9 1 9 1 11 2 15 13 16 2 1 9 1 9 7 3 1 15 3 3 15 13 1 1 11 2 10 9 1 9 7 10 9 1 10 15 13 0 10 9 0 2
9 10 9 2 11 13 1 10 11 2
16 3 2 13 1 11 16 13 15 16 13 13 15 1 10 9 2
40 10 9 13 10 10 9 1 9 7 10 9 0 1 13 9 1 9 0 7 0 1 12 7 12 9 1 10 9 2 13 10 9 1 9 1 10 9 10 9 2
31 10 9 13 0 2 10 9 3 0 7 10 9 0 13 10 9 1 9 1 9 1 10 9 16 13 10 9 1 10 9 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
10 3 15 13 1 10 9 11 11 11 2
35 10 11 1 11 2 1 11 2 11 11 2 9 2 11 11 11 2 4 13 1 10 9 11 1 12 2 1 10 9 1 11 2 3 11 2
21 15 4 13 15 9 3 1 10 9 1 10 9 2 9 7 10 9 13 9 2 2
38 10 9 1 9 7 9 0 1 10 11 1 11 1 11 2 10 11 2 11 11 2 4 13 3 8 10 9 0 13 10 9 16 13 10 9 1 9 2
15 10 9 3 4 13 15 1 9 1 15 16 13 1 9 2
14 11 13 13 7 3 13 1 13 15 1 10 9 0 2
20 3 4 13 0 2 7 9 0 2 1 10 9 10 9 13 10 9 3 0 2
21 13 10 9 10 9 1 11 11 2 13 1 10 9 16 13 10 9 7 12 9 2
36 10 9 11 2 13 15 16 13 2 10 0 9 1 10 9 2 1 15 1 13 3 1 10 9 3 1 10 9 1 13 1 10 9 1 11 2
29 10 9 13 10 9 0 7 10 9 3 0 13 10 9 1 10 12 9 2 12 9 2 1 10 9 1 10 9 2
19 10 9 4 13 1 10 0 9 1 10 9 3 1 10 9 1 10 9 2
13 10 9 8 11 11 16 1 12 13 1 12 9 2
11 9 1 10 9 7 9 1 11 11 11 2
46 13 10 9 2 15 13 1 10 9 13 1 11 1 11 7 3 15 4 13 1 10 13 10 9 1 11 1 11 2 10 9 13 1 10 0 9 7 16 15 13 10 0 12 1 11 2
19 10 9 13 10 9 2 8 11 2 8 2 8 2 2 0 9 1 9 2
36 3 10 9 2 0 7 3 15 2 1 10 9 4 13 9 7 13 2 16 13 9 7 3 9 16 3 15 4 13 12 5 10 9 1 9 2
76 2 1 10 9 2 11 13 13 1 15 2 9 1 9 2 10 9 0 1 10 9 2 3 3 13 1 11 11 1 10 9 2 10 9 2 10 9 7 9 2 7 2 1 15 2 13 13 15 13 10 9 1 9 2 1 9 7 1 9 1 10 9 1 10 9 2 2 13 11 11 2 9 1 10 9 2
66 10 9 0 2 0 1 10 11 11 4 13 1 12 1 10 9 1 10 9 11 2 9 7 9 1 10 9 1 10 9 0 0 1 10 9 2 9 1 10 9 0 1 11 11 7 9 1 9 1 10 11 1 10 11 2 13 1 13 9 1 10 9 0 1 11 2
8 11 15 13 0 1 10 9 2
23 16 3 4 13 10 12 9 15 13 3 0 13 15 9 1 0 9 1 10 9 1 12 2
18 10 0 9 1 10 0 9 1 10 9 1 9 1 9 13 10 9 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
17 3 13 9 2 3 13 10 9 2 13 1 10 9 1 9 0 2
71 1 13 1 10 15 2 10 0 9 3 0 15 13 1 13 1 10 9 12 2 1 10 9 1 10 9 0 2 1 9 1 10 11 1 11 1 11 2 1 11 11 2 11 2 12 2 2 10 11 11 2 11 2 11 11 2 12 2 2 7 10 11 2 11 2 11 11 2 12 2 2
7 15 13 9 1 10 9 2
37 1 10 9 0 1 10 9 1 10 9 2 10 9 11 11 13 10 9 1 10 11 2 1 9 1 10 9 0 1 11 11 11 7 9 11 11 2
14 3 13 1 9 1 12 16 11 15 13 9 1 11 2
71 15 3 13 1 9 7 1 9 1 13 2 16 13 10 9 1 10 9 11 11 2 4 13 10 9 0 1 10 0 9 16 13 10 9 2 7 3 13 10 9 1 10 11 2 16 10 9 16 13 1 10 9 3 4 13 2 1 10 9 0 1 10 9 16 15 13 1 13 9 0 2
43 10 0 9 1 10 9 13 0 10 9 1 10 9 16 13 10 0 9 1 10 9 0 1 9 1 3 13 9 0 3 12 9 3 1 10 9 1 10 0 9 1 9 2
34 11 11 2 11 2 11 1 10 11 2 11 11 2 12 1 11 1 12 2 13 10 9 1 9 7 9 0 0 1 10 11 1 11 2
24 10 9 0 1 10 15 15 13 10 9 1 10 11 1 11 2 11 15 13 13 1 11 12 2
36 1 9 0 2 13 12 9 1 9 2 10 9 1 10 9 1 10 9 1 15 2 13 9 0 2 7 10 9 1 10 0 9 2 13 9 2
29 11 2 13 16 4 13 10 0 9 1 9 2 1 10 15 4 13 0 2 15 10 9 2 10 9 7 10 9 2
17 13 0 7 10 9 4 13 13 1 10 9 2 0 2 3 0 2
59 4 13 1 9 0 2 1 10 9 0 1 13 15 3 0 1 10 9 0 7 3 0 1 4 0 2 1 10 0 9 2 0 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 7 3 1 10 9 0 2 2
13 10 9 13 2 3 2 10 9 1 9 7 9 2
17 11 13 10 9 2 7 13 10 9 0 1 9 1 13 10 9 2
25 10 11 5 12 9 1 10 11 1 10 11 2 9 1 10 9 2 3 13 1 9 1 9 0 2
94 1 10 9 10 9 4 1 13 9 0 1 10 9 1 11 2 3 2 11 13 7 10 9 1 15 16 15 13 10 9 1 11 1 10 0 9 1 10 9 12 1 11 11 11 2 2 1 4 13 10 9 13 13 9 1 10 9 1 13 1 9 10 9 1 10 9 1 10 9 2 10 9 13 10 9 1 10 9 3 15 13 1 10 9 1 9 1 10 9 1 10 9 0 2
11 10 11 13 1 10 9 1 10 0 9 2
19 1 10 9 2 10 9 13 9 2 9 2 9 7 9 1 10 9 0 2
14 9 0 1 10 9 11 1 11 2 10 9 1 11 2
25 1 3 1 10 9 0 13 0 1 10 9 2 3 16 10 9 15 15 13 11 13 0 7 3 2
20 15 13 10 9 1 10 15 1 11 11 3 15 13 9 1 10 9 0 0 2
22 10 9 1 11 1 10 0 9 7 10 0 9 1 10 9 2 13 16 3 4 13 2
18 3 13 7 13 10 9 2 11 11 2 1 9 1 11 1 10 9 2
33 2 2 10 9 0 1 9 15 13 1 10 0 12 9 0 1 3 12 1 10 9 12 2 2 1 10 9 3 13 12 9 0 2
36 9 0 1 9 1 10 0 9 0 2 13 10 9 1 10 9 1 10 9 13 1 10 9 13 10 15 15 13 11 2 10 9 1 10 9 2
29 10 9 11 15 13 1 10 9 9 1 10 9 1 11 2 15 1 10 12 9 0 1 10 9 1 11 2 11 2
12 10 9 13 10 9 1 10 11 7 10 9 2
13 15 3 2 13 3 0 7 10 9 13 3 0 2
32 10 9 0 2 10 9 0 1 9 2 10 9 7 10 9 0 1 13 2 13 3 13 1 10 9 7 9 1 10 9 0 2
20 1 9 2 10 9 2 3 1 10 9 0 2 13 15 1 10 9 1 9 2
23 10 0 13 9 1 9 1 9 2 7 10 9 13 10 9 1 9 0 1 10 9 0 2
20 11 13 15 1 10 9 0 1 10 9 0 1 10 0 9 1 10 9 12 2
29 1 11 2 10 9 1 10 9 15 13 1 10 0 9 2 7 3 13 10 9 0 1 10 0 9 1 10 9 2
13 3 13 13 10 0 9 1 10 9 1 10 9 2
19 1 9 1 10 11 2 10 9 13 1 0 9 13 0 9 1 10 9 2
17 10 9 16 15 4 13 1 15 2 9 2 9 2 9 2 9 2
42 10 9 1 10 11 11 13 1 15 7 1 9 1 10 9 1 11 7 10 9 1 10 11 2 1 11 15 13 10 9 3 0 7 10 16 13 1 13 10 11 11 2
21 3 13 0 13 3 1 12 9 7 13 10 9 1 13 1 10 9 1 10 9 2
12 2 3 10 9 11 3 13 15 1 10 9 2
33 11 2 15 1 10 12 9 13 1 10 9 1 11 1 10 9 1 11 2 13 10 9 0 7 0 2 1 10 9 0 2 0 2
22 10 9 4 13 16 10 9 13 10 0 9 1 10 9 1 9 15 3 4 4 13 2
28 1 9 2 10 0 9 1 9 1 9 1 9 1 10 9 1 10 9 7 10 9 1 10 9 11 4 13 2
9 13 1 11 2 1 10 9 12 2
7 10 9 13 13 9 0 2
21 1 12 13 1 10 9 12 9 0 2 1 10 15 13 1 9 12 9 1 9 2
29 1 9 2 1 10 9 7 9 1 10 10 9 1 10 9 13 10 9 1 10 9 0 11 11 2 15 2 11 2
11 2 3 13 0 16 10 9 3 13 9 2
19 13 1 9 12 9 0 13 10 9 7 3 13 9 7 4 13 1 15 2
13 10 9 11 11 3 13 10 9 2 3 15 13 2
30 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 7 11 2 1 10 9 1 11 7 9 1 11 2
27 10 9 1 10 9 15 13 3 1 10 11 1 11 2 7 13 1 10 9 11 2 1 10 9 1 11 2
11 9 2 15 2 0 1 9 1 10 9 2
12 10 0 9 13 1 9 2 9 7 9 13 2
15 1 13 10 9 1 10 11 2 4 1 13 10 9 0 2
18 10 9 13 4 13 3 1 11 1 10 9 1 9 1 11 1 11 2
53 10 9 1 10 9 13 16 10 9 1 9 1 10 9 7 10 9 4 13 1 10 9 1 10 9 16 13 9 1 10 9 1 9 2 13 13 2 1 10 9 2 7 3 1 10 9 1 10 9 1 9 0 2
14 1 3 1 9 2 3 4 13 1 15 16 15 13 2
37 11 2 1 10 9 9 7 2 9 2 2 1 9 2 13 10 9 15 13 1 11 7 2 1 0 2 1 11 10 9 1 9 13 1 9 0 2
34 11 13 10 9 1 12 9 1 9 2 12 9 2 2 3 1 3 4 13 10 9 1 9 2 7 13 15 1 0 9 1 10 9 2
28 10 9 2 16 3 13 9 0 2 13 3 1 0 1 10 9 0 1 10 9 1 15 9 9 12 1 11 2
10 15 13 10 9 1 11 11 1 9 2
38 13 16 13 13 15 1 9 1 9 0 7 1 3 9 10 9 1 9 1 2 9 2 2 1 15 9 15 13 16 15 13 9 1 10 9 3 13 2
57 10 9 1 9 4 13 1 0 9 16 15 13 13 10 9 1 10 9 1 9 1 8 2 0 1 12 9 1 0 9 7 13 10 0 9 1 10 9 1 10 9 11 11 2 16 13 1 10 9 1 10 9 0 0 1 15 2
25 13 1 11 11 2 13 10 9 1 10 9 0 16 13 10 9 2 9 7 9 2 13 10 9 2
7 10 9 7 10 9 13 2
30 13 1 10 9 2 9 7 9 1 9 2 15 13 1 3 7 3 9 1 13 1 10 9 13 10 9 1 10 9 2
22 10 9 13 0 3 1 10 9 16 13 1 10 9 0 1 13 16 10 9 13 3 2
11 15 13 3 1 11 10 11 13 1 11 2
30 10 9 1 10 9 4 1 13 1 10 9 2 4 1 13 1 10 9 9 1 10 9 1 10 9 16 13 13 11 2
44 11 11 1 11 2 13 11 11 2 2 11 11 2 2 2 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 2 13 10 9 0 0 0 1 10 11 1 11 2
25 15 13 16 11 13 10 9 10 9 14 2 0 1 9 0 0 1 10 0 11 0 1 11 11 2
21 1 9 2 10 9 4 1 13 0 9 0 2 1 10 0 9 16 10 9 0 2
32 1 10 2 9 1 10 9 7 9 1 10 9 1 10 9 1 11 2 2 11 13 13 10 9 1 10 9 1 11 1 11 2
19 3 10 9 4 13 10 9 0 7 2 1 15 2 0 7 1 0 9 2
18 10 9 0 1 13 10 9 1 10 9 2 0 7 1 10 9 0 2
22 10 9 4 13 3 1 10 11 0 2 7 10 9 1 10 9 0 13 10 9 0 2
38 10 9 1 4 13 13 10 9 0 1 11 2 13 1 12 2 1 10 9 1 10 9 4 13 3 10 9 2 13 15 1 10 9 16 13 1 12 2
38 1 12 13 10 0 9 0 1 9 1 11 2 13 3 1 9 1 11 2 7 16 13 11 2 1 10 9 2 1 11 2 11 11 2 1 10 9 2
26 1 10 9 1 9 1 10 9 1 10 9 1 11 2 11 11 13 1 11 11 12 7 13 10 9 2
26 13 1 9 7 15 13 1 10 12 1 13 1 10 11 16 13 2 16 3 4 13 10 0 9 3 2
20 13 10 9 7 9 0 2 9 1 10 11 11 11 2 13 9 7 9 0 2
18 13 3 10 12 16 15 13 13 10 9 2 13 1 9 10 0 9 2
103 7 16 1 10 9 15 4 13 10 9 1 15 7 15 2 9 1 11 1 10 11 11 2 11 2 11 11 7 1 10 11 1 10 9 2 7 10 9 2 1 11 2 10 9 1 10 9 1 9 13 16 10 11 4 1 13 9 1 10 9 0 2 15 16 15 13 10 9 0 0 1 10 9 1 11 2 7 3 4 1 13 10 9 1 10 9 1 9 2 0 1 10 9 1 9 1 10 9 7 9 1 9 2
20 13 9 1 0 9 2 3 0 9 2 13 3 3 10 9 7 13 3 0 2
30 10 9 4 13 1 9 1 10 11 11 11 2 7 3 10 9 15 4 13 1 10 9 13 16 15 13 1 15 0 2
69 15 13 2 10 9 0 1 10 9 1 10 9 2 16 7 3 13 1 9 10 9 0 1 10 11 2 11 7 11 2 9 3 10 9 0 13 3 0 1 9 1 10 9 0 1 10 9 2 2 7 10 9 0 1 10 9 1 10 9 0 16 4 13 10 9 1 10 9 2
85 15 13 1 10 9 0 1 1 12 7 12 9 1 10 11 1 10 9 2 15 15 0 1 10 9 1 10 9 13 16 13 3 1 10 9 0 11 11 2 10 9 1 10 15 13 1 9 10 11 1 10 11 2 7 10 9 1 9 1 0 9 4 4 13 1 12 7 12 9 15 1 10 11 2 15 16 15 13 1 10 9 3 0 9 2
68 1 9 1 13 9 3 3 0 1 10 0 9 1 10 9 15 13 3 3 1 10 9 0 1 10 9 7 13 1 10 10 9 10 9 9 0 7 9 16 15 13 2 1 10 9 16 15 3 13 2 3 4 13 15 10 0 9 1 9 7 2 7 9 16 15 4 13 2
12 10 9 16 13 9 1 9 15 13 9 0 2
41 1 10 9 1 11 2 1 12 2 12 12 12 9 2 12 5 2 13 1 10 9 1 9 1 9 2 1 12 12 12 2 12 5 16 15 13 1 10 9 2 2
21 1 10 0 9 0 1 10 9 0 2 15 13 10 9 1 9 0 1 10 9 2
38 11 2 11 2 12 1 11 1 12 2 2 1 9 11 11 2 13 10 9 2 9 7 9 1 9 1 9 0 7 13 9 2 11 1 11 7 11 2
16 1 9 2 1 10 9 15 13 13 10 9 1 10 9 0 2
35 16 11 4 13 1 10 0 9 2 3 13 0 1 10 9 0 2 1 15 15 3 13 9 1 13 15 1 10 9 10 9 1 13 15 2
35 13 3 9 0 1 10 9 1 10 9 2 9 1 10 11 1 11 1 10 11 11 2 9 11 1 10 9 7 9 0 1 10 11 11 2
9 3 13 9 2 9 2 7 9 2
25 10 12 1 11 1 12 13 10 9 2 16 10 9 3 15 13 3 1 10 12 1 11 1 12 2
8 11 15 13 0 1 10 9 2
29 11 2 1 10 0 16 9 9 1 11 11 7 11 11 2 13 10 0 9 0 3 1 13 15 1 10 9 0 2
20 10 9 13 16 10 9 1 2 15 1 10 9 4 13 15 1 10 15 2 2
26 1 13 10 9 2 1 10 9 12 2 11 7 10 9 1 10 9 13 3 1 9 1 10 9 0 2
14 4 13 1 10 11 11 2 11 2 1 10 9 0 2
27 10 9 1 0 9 15 13 1 11 2 9 1 11 2 1 11 2 9 1 11 2 7 11 2 11 2 2
26 1 13 10 0 9 2 11 15 13 1 13 1 10 9 7 13 3 1 11 7 1 15 1 10 9 2
20 4 13 1 10 9 13 1 9 1 10 9 2 1 10 15 15 13 11 11 2
22 1 9 1 9 15 4 13 9 1 8 9 7 15 13 9 1 10 9 7 10 9 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
25 1 13 15 10 9 2 10 9 13 13 1 10 9 2 7 13 16 13 16 11 13 4 13 9 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
42 1 10 0 9 2 9 1 11 11 4 13 10 9 0 2 7 1 9 3 0 2 1 10 9 13 1 10 9 0 2 12 9 1 10 10 9 1 10 9 8 2 2
11 13 10 9 13 1 12 9 2 12 2 2
18 13 13 9 1 10 9 1 10 9 1 10 9 16 13 1 11 11 2
16 10 9 13 1 9 1 10 9 7 11 13 1 10 9 0 2
26 1 12 2 13 1 11 11 11 2 10 9 0 1 11 11 11 16 13 10 0 9 1 10 9 0 2
17 13 1 0 9 1 11 1 10 9 7 3 4 13 9 1 11 2
38 11 11 2 11 2 13 10 9 0 13 1 11 11 2 11 11 7 11 11 7 13 1 10 9 0 11 2 11 11 1 10 9 0 2 11 2 11 2
52 10 9 1 10 15 15 13 1 10 11 11 10 9 1 9 13 10 9 13 11 2 11 2 9 13 10 9 1 10 9 0 16 13 0 2 2 1 10 9 1 10 9 1 11 2 1 10 9 0 1 11 2
11 10 9 2 11 11 2 13 15 15 13 2
30 10 12 1 11 1 12 11 11 4 13 1 10 11 7 13 1 12 9 1 2 2 11 2 11 2 10 9 1 11 2
12 10 9 1 9 13 1 12 8 2 9 8 2
41 10 9 1 10 9 13 13 1 10 9 10 9 1 10 9 1 9 1 13 9 1 9 7 9 1 9 2 3 1 13 3 0 10 9 1 10 9 1 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
44 3 1 13 15 1 9 0 2 11 15 13 1 10 9 1 10 9 16 15 13 1 11 2 13 11 2 7 13 10 9 1 9 1 10 9 1 11 2 3 13 13 10 9 2
23 10 0 11 11 3 15 13 0 1 12 9 0 7 10 9 1 12 9 1 10 10 9 2
21 10 9 1 9 7 9 0 2 13 1 10 9 10 9 1 10 9 1 9 0 2
81 15 1 10 9 3 0 2 1 15 1 10 9 1 10 9 2 13 10 0 9 1 10 9 1 9 16 13 10 9 2 1 15 10 9 1 12 9 1 10 9 7 12 1 10 9 1 10 9 1 9 13 1 4 13 10 9 1 2 9 2 1 13 1 10 9 1 9 1 10 16 2 1 10 9 2 13 12 9 1 9 2
48 10 12 1 11 2 13 1 13 9 1 10 9 12 11 11 11 11 2 13 1 11 11 5 11 11 12 1 10 0 9 2 7 13 10 12 1 11 1 11 9 2 11 11 8 11 11 2 2
23 10 9 0 13 13 10 9 1 10 0 9 0 1 10 9 1 10 1 11 11 1 11 2
10 3 2 13 10 0 9 2 13 11 2
49 11 11 13 10 9 2 8 2 8 2 0 16 4 1 13 10 0 9 16 2 13 1 10 9 2 4 1 13 15 3 1 2 10 9 1 10 0 9 2 3 10 9 15 13 1 10 9 2 2
18 10 11 13 1 9 1 9 1 9 1 13 10 9 1 10 9 0 2
40 10 9 0 13 10 9 1 9 0 2 13 1 0 9 16 2 1 10 9 3 0 2 15 4 13 1 10 2 9 0 2 1 10 9 1 4 2 13 2 2
26 10 12 5 9 13 1 10 9 1 9 1 15 9 1 10 9 11 1 11 2 3 10 9 1 11 2
21 1 9 1 10 9 1 11 2 10 9 11 11 15 13 1 13 10 9 1 9 2
11 10 9 1 11 15 13 13 1 10 9 2
69 10 9 13 1 13 15 2 15 2 9 1 10 9 2 13 10 9 16 15 15 13 1 13 9 1 9 7 3 7 3 2 10 3 9 13 13 9 7 13 1 9 1 10 9 16 13 1 10 0 9 2 9 0 1 10 0 9 0 1 15 1 10 0 9 0 1 10 11 2
26 10 9 13 1 12 1 10 0 9 1 9 1 11 2 16 1 12 4 13 1 11 2 11 7 11 2
28 11 11 13 10 9 3 0 1 10 9 2 13 10 12 1 11 1 12 1 10 11 11 2 0 11 11 2 2
25 10 9 1 10 11 1 11 7 11 11 15 13 13 1 10 9 0 1 10 11 1 11 2 11 2
19 1 9 15 15 13 10 9 1 9 7 9 7 1 9 1 10 0 9 2
18 13 9 1 9 7 9 7 9 1 10 11 11 1 10 11 1 11 2
17 4 13 0 1 10 9 1 10 9 1 10 9 0 1 11 11 2
30 11 11 11 11 2 11 2 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 13 10 9 7 9 0 2
17 11 13 10 9 1 10 11 13 1 9 7 9 2 13 1 11 2
26 10 9 2 1 10 15 15 13 10 9 0 2 4 1 4 13 16 13 1 10 9 0 1 10 9 2
18 4 13 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9
26 11 11 7 11 2 11 2 11 2 12 2 11 2 11 2 12 1 11 1 12 2 13 10 9 0 2
23 1 11 13 10 0 1 15 9 1 10 9 1 10 9 11 2 1 3 15 13 10 9 2
28 1 9 1 10 9 1 9 1 11 10 11 1 11 11 7 10 9 2 10 9 4 13 9 1 10 9 0 2
22 1 10 9 11 2 10 9 11 4 13 15 1 10 0 9 1 9 1 10 11 11 2
38 3 13 1 11 2 7 1 10 9 0 3 4 4 13 1 9 0 1 11 2 1 15 15 4 13 1 13 9 1 11 2 1 10 9 1 11 11 2
53 2 15 15 13 10 9 3 2 13 11 2 16 10 9 0 13 1 10 0 7 0 9 1 13 1 10 9 0 7 13 2 1 9 7 1 9 0 2 10 9 1 10 9 16 4 13 10 10 9 2 2 13 2
10 13 9 0 2 7 0 2 7 0 2
5 10 9 13 0 2
7 13 1 11 2 1 12 2
24 1 10 9 2 10 9 16 11 13 1 11 11 13 1 10 11 1 11 11 1 11 1 11 2
20 10 11 1 10 11 11 4 13 1 1 0 9 7 13 10 9 1 12 5 2
50 1 15 15 13 1 13 1 10 9 1 15 1 10 9 16 15 13 16 15 13 0 1 10 9 16 13 2 13 15 7 13 1 3 13 15 15 16 15 13 0 16 3 4 13 10 9 1 13 15 2
24 15 13 1 10 9 7 13 15 1 9 0 2 7 13 1 9 16 3 13 9 1 10 11 2
22 10 9 15 13 2 1 0 9 2 1 10 9 1 10 11 11 11 1 11 11 11 2
20 9 1 9 1 10 11 11 1 12 9 2 0 2 2 13 1 11 1 12 2
37 10 12 1 11 10 9 2 1 10 9 1 10 9 11 2 13 11 1 10 9 1 0 9 7 13 10 9 2 0 1 10 9 1 11 7 11 2
19 13 1 10 9 0 16 15 13 10 9 1 10 9 0 16 4 1 13 2
20 1 10 9 1 10 9 15 13 9 1 10 9 2 11 11 7 11 11 2 2
28 10 9 2 16 13 10 0 9 0 11 2 4 13 1 10 9 1 9 0 0 2 9 7 1 10 9 0 2
36 16 11 13 10 9 1 9 1 3 1 12 9 2 15 3 13 0 1 9 1 9 0 1 9 1 13 9 1 9 1 0 9 7 10 9 2
32 10 12 9 15 13 9 7 13 1 13 10 9 7 11 4 1 13 1 10 0 9 1 11 1 10 0 9 7 13 10 9 2
66 10 11 11 4 13 10 9 1 11 1 10 12 0 9 16 4 13 13 10 9 10 9 11 11 7 13 16 10 9 13 15 1 15 16 3 13 1 10 11 0 1 11 11 2 11 2 10 9 0 13 15 1 10 9 7 13 15 1 10 9 1 13 9 1 15 2
25 3 13 15 1 10 10 9 7 13 12 5 1 9 2 3 13 3 7 16 13 12 5 1 9 2
51 3 1 13 15 10 11 2 12 11 13 1 10 11 11 1 10 11 2 12 11 13 1 10 9 2 15 13 10 11 2 11 1 4 13 1 10 8 2 12 2 7 3 1 10 11 11 2 12 11 2 2
15 10 9 0 15 13 1 10 9 7 1 9 1 10 9 2
27 1 10 9 2 1 9 4 13 16 13 10 0 9 1 10 9 2 16 4 13 1 13 10 9 10 9 2
8 10 9 0 4 13 10 9 2
24 13 1 11 1 11 1 12 7 13 1 10 9 1 10 11 10 12 1 11 1 10 0 9 2
14 3 1 10 9 11 13 1 9 16 10 9 13 0 2
26 10 9 1 9 2 16 15 13 3 7 13 10 9 0 7 0 16 10 9 2 13 10 9 3 0 2
16 10 9 1 10 9 13 10 12 5 1 9 16 13 10 9 2
36 15 1 10 9 3 0 7 3 10 9 1 10 0 9 1 10 9 1 11 2 13 10 9 1 9 11 11 15 1 12 13 10 9 1 9 2
27 1 9 2 15 12 1 12 13 12 2 0 2 3 3 10 9 16 15 13 10 9 0 12 7 12 3 2
46 10 9 15 13 1 10 9 2 8 2 13 10 12 9 2 7 10 9 2 11 11 2 1 12 9 2 8 2 13 10 12 9 1 9 1 15 1 10 15 1 10 12 9 0 0 2
6 13 9 0 7 0 2
19 3 13 13 10 9 1 10 9 9 2 15 13 15 3 1 16 15 13 2
15 15 13 3 3 16 10 9 3 0 15 13 9 3 0 2
13 11 11 13 10 9 7 9 0 1 10 9 12 2
30 16 13 11 1 10 9 11 2 10 9 15 4 13 9 1 9 1 10 16 15 13 3 4 13 15 1 9 1 11 2
19 10 9 0 4 4 13 1 9 2 7 1 10 13 0 13 10 9 0 2
44 10 11 7 11 10 11 2 13 10 0 9 0 1 10 12 9 1 11 1 10 9 11 11 1 10 11 7 13 1 10 9 1 11 11 13 1 10 9 1 11 2 1 11 2
26 1 10 9 13 13 10 9 13 15 13 1 10 9 1 9 2 16 10 9 11 13 8 1 13 15 2
42 9 0 13 1 13 1 10 9 0 16 15 4 13 7 15 15 13 1 9 0 10 12 1 11 2 7 11 13 16 11 15 4 1 13 1 15 9 3 1 10 9 2
16 10 9 2 11 2 13 10 9 1 9 0 1 10 9 11 2
29 3 2 13 16 10 9 3 13 13 9 9 1 9 7 1 9 1 9 16 13 10 9 1 10 9 11 2 11 2
21 11 12 3 13 1 10 9 16 13 13 15 10 9 1 10 9 1 1 10 9 2
30 3 4 13 16 15 13 10 9 1 10 0 9 7 9 1 11 7 1 15 13 1 9 10 0 9 1 10 11 2 2
18 13 10 9 1 10 9 1 11 11 2 4 13 9 1 10 9 0 2
47 10 9 1 11 13 15 0 13 7 3 13 1 10 11 11 2 9 16 4 13 10 9 1 13 10 9 1 9 1 9 7 4 13 10 9 3 0 16 4 4 13 10 9 1 10 11 2
19 11 13 10 9 1 10 9 11 2 13 1 10 9 1 11 2 1 11 2
36 1 15 11 1 11 13 10 9 2 10 9 2 10 9 2 7 10 9 16 15 13 13 10 3 0 9 1 13 1 10 9 1 13 10 9 2
33 4 13 1 9 7 13 0 9 13 1 10 9 0 1 10 9 2 16 1 9 1 10 9 10 9 3 4 13 7 13 1 0 2
31 7 2 10 9 1 11 13 1 9 1 9 1 10 9 2 12 2 7 10 0 9 3 0 1 10 11 11 2 12 2 2
14 10 9 4 4 13 1 10 9 0 10 12 1 11 2
47 10 9 15 13 1 10 9 0 2 9 0 2 9 1 9 1 10 9 1 9 2 1 10 9 0 2 9 7 9 1 9 2 1 10 9 0 1 10 9 2 3 7 9 1 10 9 2
26 11 13 10 0 9 3 0 1 11 2 7 10 9 0 7 0 1 10 9 1 10 9 0 1 11 2
34 10 9 1 10 11 13 15 1 10 12 9 0 16 13 10 9 1 11 1 10 9 1 11 2 1 10 9 1 10 9 0 1 11 2
24 1 9 1 13 15 1 10 9 1 10 9 2 13 10 9 10 16 4 7 13 0 1 15 2
11 10 9 4 13 3 0 1 10 0 9 2
19 10 11 1 11 13 10 9 1 10 15 13 10 0 9 1 10 9 0 2
9 10 9 15 13 0 7 3 0 2
21 1 9 15 13 10 9 1 10 9 1 10 9 13 1 11 1 12 2 13 3 2
5 13 11 1 11 2
27 11 2 1 9 11 11 7 11 11 11 2 13 15 1 10 9 0 1 10 9 1 9 1 11 1 11 2
30 10 9 1 11 11 2 1 9 2 11 11 11 2 2 13 1 12 2 13 15 1 12 9 1 10 9 0 1 11 2
13 11 13 10 0 9 1 11 1 13 10 9 13 2
20 11 11 13 10 9 0 2 16 13 1 9 9 1 10 9 1 9 1 11 2
40 1 12 2 1 10 0 9 0 2 13 10 9 1 11 2 9 1 9 2 9 1 10 15 13 10 9 1 10 9 0 16 3 3 13 1 10 9 1 11 2
104 1 0 9 2 13 13 10 9 1 10 9 0 2 9 7 9 2 9 2 1 15 0 0 2 9 0 7 9 0 2 2 13 3 9 1 10 9 1 10 9 7 10 9 1 9 1 9 0 1 10 9 2 13 1 10 9 1 10 9 1 2 9 0 16 4 13 10 9 1 9 1 10 9 1 9 1 9 2 9 7 9 0 2 2 13 16 10 9 0 7 10 9 0 0 13 9 1 10 9 0 7 0 0 2
9 2 16 16 15 13 13 1 11 2
14 10 9 1 9 13 1 10 12 9 1 10 9 0 2
8 10 9 4 13 1 11 11 2
39 3 10 9 3 0 15 4 7 13 13 10 9 7 0 9 1 11 2 1 11 2 13 1 10 9 11 11 1 11 1 12 2 13 10 9 1 10 9 2
16 10 9 0 2 13 1 9 2 13 10 9 2 0 1 9 2
14 3 13 9 1 10 9 2 1 9 13 1 11 11 2
22 1 10 9 10 9 1 10 9 4 13 10 0 2 10 9 2 0 2 1 10 11 2
25 15 13 7 3 2 10 9 1 9 1 11 13 1 11 3 13 10 15 9 16 4 13 1 11 2
6 11 11 2 12 2 2
43 1 10 11 1 10 11 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
24 11 13 9 1 9 1 9 2 9 1 9 7 9 1 11 11 11 11 1 11 11 2 11 2
18 1 10 0 9 2 10 9 13 1 12 9 1 12 12 2 12 9 2
20 13 10 9 1 10 9 0 1 11 7 9 1 9 1 10 11 11 1 11 2
65 3 13 4 1 13 9 1 9 1 9 7 15 13 13 10 9 1 9 1 9 2 15 16 15 13 10 9 1 10 9 1 11 11 2 10 9 1 10 11 2 1 10 11 12 2 16 13 1 11 1 9 1 10 12 7 13 1 11 2 11 11 7 10 11 2
19 1 15 3 2 13 1 9 1 10 0 9 2 1 10 15 13 1 11 2
29 1 10 0 9 2 13 10 9 0 1 13 9 7 9 16 13 16 10 9 0 13 2 1 16 10 9 15 13 2
16 10 15 3 3 13 10 0 11 15 13 10 9 1 10 9 2
16 11 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2
14 3 13 1 10 9 2 7 3 1 15 15 13 2 2
38 3 13 9 1 11 11 2 11 7 11 1 10 12 5 1 9 13 1 15 16 4 13 1 10 0 9 13 1 10 9 2 3 7 4 7 13 15 2
26 3 2 4 13 9 1 11 1 10 10 9 1 11 2 9 1 11 2 3 15 4 13 11 11 11 2
11 10 9 13 10 11 12 1 11 1 12 2
75 11 13 16 10 9 16 4 13 11 7 10 9 1 11 1 10 11 1 13 9 1 10 9 1 10 9 7 3 13 15 15 1 10 9 16 15 13 16 13 0 10 9 0 1 11 2 13 10 9 7 13 16 10 8 9 1 10 9 0 13 10 9 2 13 7 13 1 13 13 2 1 0 9 2 2
27 1 10 9 0 9 15 13 10 11 1 11 2 2 10 11 1 11 2 7 10 9 1 2 10 11 2 2
20 1 10 0 9 2 10 9 13 12 9 1 10 11 11 1 9 1 11 11 2
34 11 2 1 9 11 2 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
41 3 13 10 9 1 13 9 0 3 3 1 9 7 0 9 1 9 16 4 13 9 1 10 9 1 9 16 15 4 13 1 10 0 9 1 10 9 1 10 9 2
22 10 0 9 11 13 10 9 1 10 11 11 9 16 13 10 0 9 1 12 7 12 2
55 3 2 3 13 0 1 1 10 3 12 9 0 7 9 1 9 2 16 13 9 1 10 9 2 7 1 10 9 1 11 7 11 2 15 1 11 11 2 16 15 13 1 9 1 9 1 9 2 16 10 9 13 3 0 2
20 9 0 2 1 10 9 15 13 11 1 10 13 10 9 2 10 9 4 13 2
43 10 9 13 1 10 9 16 10 9 1 10 11 11 1 11 1 11 2 1 10 9 1 12 9 2 13 0 9 1 12 9 0 7 13 1 12 3 15 4 13 1 9 2
6 13 10 11 1 11 2
7 11 13 1 11 2 11 2
29 0 15 1 13 15 10 9 1 10 9 7 3 13 1 10 9 2 7 1 13 10 9 3 1 10 9 1 9 2
28 1 10 9 8 13 3 12 9 16 13 1 5 8 2 7 12 9 16 13 1 10 0 9 1 10 8 8 2
46 10 9 0 1 10 9 1 12 4 13 10 9 13 9 0 7 11 13 1 10 9 1 11 7 11 11 2 3 10 9 15 4 13 7 13 1 13 15 1 9 2 13 10 9 0 2
48 10 11 4 1 10 9 13 10 9 0 10 15 13 1 9 7 15 13 11 2 9 16 13 1 10 11 11 2 15 1 10 9 16 13 16 15 13 1 10 9 0 16 4 1 13 10 9 2
21 1 10 9 0 1 9 0 2 10 15 11 13 3 0 1 10 9 11 2 11 2
4 3 15 13 2
16 11 2 9 0 2 13 10 0 9 1 10 9 0 11 11 2
21 10 9 13 0 2 13 1 9 2 0 2 0 1 12 5 1 0 2 3 13 2
27 15 4 13 10 0 9 1 10 9 0 2 7 3 13 9 0 3 7 3 13 0 1 3 16 10 11 2
14 8 2 9 9 8 2 13 10 9 0 1 10 9 8
26 13 13 16 10 9 2 3 15 13 1 10 9 1 11 2 10 9 0 1 10 9 7 10 0 9 2
26 10 9 1 10 9 1 10 9 13 16 4 13 1 10 9 1 11 2 10 15 13 10 9 1 15 2
55 10 9 13 0 1 13 15 1 10 9 7 13 15 1 10 9 1 13 1 11 16 2 10 9 16 13 10 9 1 10 9 15 13 15 9 1 10 9 2 2 15 15 13 1 10 9 0 1 10 9 15 13 11 11 2
16 3 15 13 10 9 0 2 15 13 10 9 7 15 13 0 2
18 15 13 16 1 3 1 11 1 10 9 3 13 10 12 9 1 11 2
33 10 9 1 10 9 2 3 10 9 13 0 9 1 10 9 2 7 3 10 9 0 13 0 9 1 9 7 9 2 11 12 2 2
20 10 9 13 10 9 3 0 2 13 10 9 12 1 10 9 1 11 1 12 2
9 10 9 13 1 11 7 10 11 2
20 1 10 9 1 9 16 13 3 1 10 9 2 10 9 4 13 9 3 0 2
23 10 9 3 13 10 9 1 13 9 2 16 1 11 2 13 9 1 10 9 1 10 9 2
23 15 4 13 9 1 10 0 9 2 2 1 15 10 9 0 13 1 10 9 1 12 9 2
42 1 10 11 1 11 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
49 10 9 13 1 10 9 0 8 2 2 3 13 1 8 2 2 16 13 10 9 2 2 13 1 10 9 8 2 9 2 9 2 2 8 2 9 2 9 2 7 8 2 9 2 9 2 9 2 2
21 3 15 13 1 10 9 13 1 10 9 1 10 9 1 16 10 13 1 10 9 2
11 3 10 9 13 1 10 0 9 1 9 2
36 10 9 1 11 2 15 13 13 1 10 9 1 10 9 1 11 1 11 2 11 2 13 15 1 10 12 9 1 10 9 0 2 9 1 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
71 10 9 15 13 16 13 9 16 1 13 0 1 10 9 7 13 10 0 9 0 0 1 0 3 13 10 9 0 2 1 3 4 13 10 9 1 9 1 10 9 0 2 7 1 9 3 13 10 9 0 2 1 13 9 1 10 9 16 15 4 13 7 13 9 1 9 1 10 9 2 2
19 9 3 0 2 1 8 7 8 1 10 12 7 12 13 1 3 0 9 2
59 10 9 1 10 9 0 13 10 0 9 1 13 9 1 13 15 1 9 1 9 0 2 9 2 2 15 13 3 16 1 0 13 10 9 0 9 1 9 1 10 9 1 10 9 2 15 16 13 16 0 9 1 9 15 13 1 10 9 2
12 10 9 13 1 9 7 13 13 15 12 9 2
45 9 13 10 9 0 16 15 13 1 9 1 13 9 1 10 9 3 0 16 13 1 10 9 2 13 13 1 10 9 1 9 0 1 10 9 16 15 13 1 10 9 1 10 9 2
19 11 13 1 11 13 15 13 1 10 11 2 13 16 4 13 1 10 9 2
30 1 9 10 9 3 13 10 9 16 15 13 1 10 9 13 10 9 0 1 11 7 11 1 11 7 10 9 0 3 2
6 13 2 7 4 13 2
38 3 10 9 13 1 10 9 1 11 11 1 10 9 11 11 1 10 9 2 11 2 11 9 2 13 1 13 1 11 3 1 16 15 13 9 7 9 2
54 1 10 9 2 11 13 1 10 0 9 1 10 9 0 2 10 0 9 10 11 2 12 15 13 1 10 0 9 0 2 1 9 1 16 1 10 8 2 9 3 13 2 10 9 1 10 9 1 10 0 7 0 9 2
13 11 13 10 9 9 1 11 11 1 11 1 12 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
13 15 13 1 10 9 13 1 10 9 1 10 9 2
39 15 13 1 10 9 11 1 11 2 11 10 12 1 11 1 12 2 10 0 9 1 11 12 1 11 2 11 2 11 11 1 11 2 7 1 11 1 11 2
43 11 11 1 11 13 16 2 10 9 3 0 1 11 11 13 13 16 10 9 1 0 9 2 9 1 10 0 7 0 9 4 13 3 13 1 10 9 1 10 0 9 2 2
20 11 8 11 2 11 11 13 10 9 0 15 4 1 4 13 1 10 11 11 2
19 15 16 3 13 0 13 16 10 9 13 1 9 1 13 7 15 13 15 2
43 1 10 9 1 10 9 1 10 11 11 2 10 11 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 13 1 9 0 7 2 12 5 2 12 5 5 13 9 2
17 1 10 0 9 1 9 2 10 0 9 1 11 2 11 13 11 2
21 11 13 9 1 10 9 0 1 10 9 1 10 11 7 1 9 0 1 11 11 2
29 13 9 1 11 7 11 1 10 11 1 11 2 16 15 13 1 10 9 12 10 2 11 1 11 1 10 9 2 2
25 3 1 13 12 9 1 10 11 1 11 11 2 3 13 11 2 11 1 12 15 13 1 10 9 2
32 15 13 10 9 1 10 11 11 1 10 11 1 11 2 10 9 1 8 15 3 4 13 1 11 7 10 11 1 10 11 11 2
27 10 11 0 4 13 1 11 11 12 9 7 3 13 1 10 0 9 1 10 9 1 12 9 1 9 3 2
26 10 9 13 0 1 11 2 10 0 9 1 10 9 13 1 11 2 7 13 10 9 1 9 1 11 2
10 1 9 3 13 7 10 9 4 13 2
53 10 9 0 1 11 13 10 9 13 7 13 1 10 9 0 2 13 10 9 1 10 9 0 2 1 10 0 9 0 1 3 1 10 9 1 9 2 9 7 9 2 4 15 13 15 1 15 1 3 1 10 9 2
22 11 2 11 13 10 9 0 0 1 9 2 0 1 10 9 1 9 11 11 7 11 2
20 10 9 0 1 10 9 0 4 13 1 10 9 0 0 11 11 5 11 11 2
61 10 9 0 13 1 9 2 3 7 1 9 0 7 0 0 1 10 9 1 10 9 7 1 10 9 0 16 15 13 1 10 9 0 16 15 13 1 10 9 1 10 9 2 4 13 1 10 9 1 11 16 13 9 1 10 9 0 13 1 11 2
32 11 11 13 10 9 1 9 0 9 1 10 9 1 10 9 2 0 1 8 0 2 1 10 9 1 11 1 10 11 1 11 2
45 10 9 1 10 9 12 13 10 9 1 11 2 13 11 7 13 10 11 11 1 10 9 1 10 0 9 1 11 2 7 10 0 9 15 4 7 13 13 10 1 10 9 1 9 2
49 1 9 0 2 15 13 10 9 1 13 10 9 1 10 9 1 9 16 4 13 9 1 10 9 2 8 2 8 2 1 10 9 0 2 7 16 3 13 0 1 13 15 16 13 10 9 1 11 2
34 10 9 4 3 13 1 13 1 10 9 0 2 11 11 2 2 7 3 3 13 15 16 15 13 3 2 16 10 15 13 1 11 11 2
25 10 9 0 13 16 10 9 1 10 9 0 15 13 13 3 1 13 1 10 9 1 10 9 11 2
39 10 0 9 1 10 9 7 10 9 1 10 9 1 11 11 2 10 9 16 13 2 10 11 11 2 7 2 11 11 2 2 3 13 10 9 1 9 0 2
18 10 9 13 0 1 11 2 11 2 11 7 1 3 9 1 11 11 2
30 10 11 11 1 11 13 10 9 0 13 1 10 9 1 11 2 1 10 9 0 1 10 11 11 1 11 2 11 2 2
32 10 11 11 11 13 10 9 1 9 1 11 7 10 9 13 1 10 11 11 1 11 2 10 9 1 9 3 0 1 10 9 2
34 15 13 10 9 1 0 9 0 2 9 7 9 16 13 10 9 7 10 9 1 10 9 15 10 9 13 1 15 9 1 9 7 0 2
14 10 9 4 1 13 15 2 1 0 1 10 9 0 2
23 11 11 2 1 10 9 2 4 13 16 1 9 1 10 1 3 2 15 13 9 0 2 2
15 15 13 1 9 0 1 10 9 1 9 2 9 7 9 2
25 13 10 9 1 10 9 11 9 3 7 13 3 10 0 9 1 11 2 11 2 2 12 9 2 2
36 1 9 2 10 9 1 9 0 1 12 13 1 12 1 12 2 15 15 15 13 16 10 9 15 4 13 15 3 1 10 12 1 12 1 12 2
29 3 15 13 12 12 9 2 7 11 13 1 10 9 7 13 12 12 7 13 1 13 10 9 2 1 15 15 13 2
37 10 9 0 2 12 2 15 4 13 7 13 10 9 1 11 2 11 7 11 2 10 9 16 15 4 13 1 10 9 11 12 7 9 11 2 11 2
28 10 9 13 13 3 15 13 10 9 2 10 9 1 10 9 2 10 9 2 10 9 1 9 7 9 2 8 2
31 16 10 9 16 13 1 10 9 13 9 7 9 2 13 10 9 7 15 13 1 9 3 3 2 11 2 12 2 12 2 2
35 10 9 3 0 7 0 13 2 10 9 0 16 10 9 15 4 13 2 7 16 10 0 9 4 13 1 10 9 1 10 0 9 1 9 2
27 13 10 9 1 10 9 3 0 2 13 15 1 13 1 10 9 2 7 13 16 3 13 3 1 10 9 2
30 3 1 10 9 1 12 7 12 2 9 1 9 0 1 15 11 7 9 1 11 2 4 13 1 13 10 9 0 0 2
9 10 9 13 10 9 0 7 0 2
35 10 9 1 9 4 13 3 1 10 9 16 13 1 9 0 0 2 7 10 9 1 9 4 13 3 1 9 1 9 16 13 3 1 9 2
53 1 12 15 13 1 15 10 9 0 16 15 13 1 13 10 9 1 13 15 1 0 1 10 9 0 2 13 1 9 8 0 1 10 9 0 11 2 16 13 4 13 1 9 1 10 9 1 16 15 15 4 13 2
23 11 11 2 8 12 1 11 1 12 1 11 2 9 2 11 2 13 10 8 9 0 0 2
31 11 11 11 2 11 2 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 13 10 9 2 9 7 9 0 2
38 11 13 16 1 11 13 10 9 0 2 16 13 1 9 0 2 16 2 4 13 1 10 9 1 11 16 13 10 9 1 9 7 4 13 10 9 2 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
21 10 12 1 11 13 1 9 1 10 0 9 1 10 9 2 11 11 1 10 11 2
30 9 0 7 0 16 13 3 1 10 9 0 7 9 1 15 13 10 9 1 9 16 10 9 13 1 10 9 1 9 2
43 10 9 1 12 9 15 13 1 1 10 9 1 12 7 12 9 2 9 1 0 9 1 9 7 9 2 16 13 1 10 9 1 10 9 16 1 0 9 15 13 1 11 2
22 11 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
9 4 3 13 3 10 9 1 9 2
40 1 11 1 12 2 1 10 9 1 10 0 11 11 0 16 13 1 9 16 13 1 10 9 1 11 1 0 9 1 11 8 1 11 2 15 4 13 7 13 2
61 13 12 12 9 1 9 2 1 10 15 10 12 5 4 13 1 10 0 9 2 10 12 5 1 9 0 1 7 1 9 0 2 10 12 5 1 9 2 12 5 0 2 12 5 1 13 2 1 7 1 9 0 2 7 10 12 5 1 0 9 2
17 15 4 13 3 1 10 9 0 2 13 10 0 9 7 0 9 2
10 1 10 9 3 15 4 13 1 9 2
47 1 10 9 10 9 4 13 10 9 7 9 2 13 1 9 1 10 9 2 13 9 3 7 1 9 7 13 1 0 9 1 10 9 1 9 2 9 0 2 9 1 9 7 9 2 8 2
21 10 9 1 10 9 1 9 15 4 13 3 1 9 7 3 15 13 10 9 0 2
21 15 13 1 11 11 2 11 1 11 2 11 2 11 2 7 2 3 2 11 11 2
49 10 9 0 1 10 12 9 7 10 0 9 1 11 7 11 13 1 10 11 1 11 1 12 13 1 10 9 0 1 13 10 9 1 4 1 13 10 9 1 11 13 10 9 1 10 11 1 11 2
39 3 13 1 10 9 1 10 11 11 11 11 11 11 2 10 9 1 11 11 11 11 5 11 11 2 13 0 3 1 13 10 9 1 11 11 7 11 11 2
9 10 9 15 13 9 1 12 8 2
31 10 9 16 13 0 9 13 11 11 2 11 11 2 8 13 1 12 16 13 13 1 13 1 10 9 0 10 9 3 0 2
18 10 9 15 2 8 2 8 15 13 16 13 10 9 1 10 12 5 2
14 1 10 9 1 12 2 13 12 9 13 1 11 11 2
22 10 11 13 1 10 9 3 13 1 9 2 1 12 9 1 9 7 12 9 1 9 2
43 13 1 0 9 2 1 10 9 0 1 11 2 10 9 0 1 11 7 15 9 2 3 7 10 9 1 10 9 1 10 9 2 3 13 16 15 9 13 9 1 10 9 2
46 11 4 4 13 3 1 10 2 9 1 9 2 1 10 10 0 9 2 7 10 9 1 10 9 12 7 12 13 16 3 1 10 9 2 10 9 13 3 0 9 2 13 15 1 9 2
27 11 2 3 0 2 0 7 16 13 0 1 10 9 0 2 13 9 1 10 9 1 15 1 13 10 9 2
41 10 9 9 0 13 10 9 1 10 9 1 10 9 0 1 15 15 13 2 1 10 9 0 10 9 0 2 16 13 9 16 13 1 10 9 3 0 1 10 9 2
18 10 12 9 4 13 1 10 9 0 7 3 4 13 1 10 0 9 2
20 13 1 12 9 1 9 1 12 9 2 9 2 9 2 9 7 9 1 9 2
19 11 11 13 10 9 0 2 1 10 9 1 11 2 9 1 10 9 0 2
20 11 11 11 7 11 11 11 13 10 0 9 1 10 9 1 10 9 0 11 2
8 13 10 0 9 1 10 9 2
24 3 0 2 3 13 1 10 11 11 1 10 9 2 11 7 10 9 13 1 11 7 15 13 2
7 13 1 11 11 1 12 2
42 10 9 0 11 11 15 13 3 1 0 9 0 1 10 9 1 10 11 12 1 11 2 1 13 1 10 9 11 11 2 7 13 3 1 10 9 1 10 9 11 11 2
20 9 0 15 13 1 9 1 2 9 1 10 15 1 9 0 13 10 0 9 2
13 12 9 1 10 9 0 7 10 10 12 1 9 2
23 10 11 11 13 10 9 10 9 1 9 1 11 11 16 13 10 12 9 1 9 1 9 2
14 1 0 10 9 0 1 10 9 0 13 0 7 0 2
13 11 11 13 10 9 1 9 11 1 10 9 11 2
24 3 4 13 1 10 9 0 13 1 10 9 2 3 1 9 2 9 0 2 7 9 1 9 2
14 10 9 2 9 2 9 7 9 13 10 9 2 9 2
44 13 10 9 1 9 1 11 2 7 3 1 13 10 0 9 1 10 2 11 11 11 2 9 13 1 10 11 1 12 2 13 10 9 1 10 9 1 11 1 10 11 1 11 2
28 10 11 1 11 11 2 11 2 13 10 9 3 0 13 1 10 9 0 16 13 1 9 1 9 7 1 9 2
25 13 1 10 9 1 10 9 11 2 11 15 13 2 0 2 12 2 7 11 10 9 2 12 2 2
24 10 0 9 0 0 2 1 11 1 12 1 11 1 12 2 13 1 9 7 9 1 10 9 2
7 15 13 9 1 10 9 2
46 10 9 1 9 3 13 3 3 13 9 2 3 15 13 1 9 0 1 3 9 1 9 2 1 9 1 10 9 0 2 2 7 3 9 0 1 9 7 9 7 10 9 1 10 9 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
37 15 13 0 9 1 9 1 9 0 1 10 9 2 13 1 9 0 1 10 11 7 10 9 2 7 13 10 0 9 1 9 0 1 10 9 0 2
45 13 1 10 9 1 11 11 2 11 11 2 1 10 9 2 16 13 10 11 11 2 9 1 10 0 2 1 10 9 11 11 2 3 16 11 11 2 10 9 0 2 13 13 9 2
64 13 9 1 10 0 9 1 9 0 1 10 9 11 2 1 15 2 11 11 2 11 11 2 11 11 2 11 11 11 2 12 2 2 11 11 2 11 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11
33 1 10 9 2 1 10 11 15 13 16 10 9 1 11 1 10 9 13 10 9 1 11 2 16 4 13 3 3 1 10 9 0 2
9 13 1 10 9 1 11 1 12 2
47 1 10 15 4 7 13 10 9 0 2 16 13 10 9 1 10 9 1 9 2 9 7 2 1 15 2 9 2 13 1 9 10 0 9 0 1 10 9 3 7 10 0 9 1 0 9 2
25 10 9 13 13 1 9 0 2 15 4 13 1 9 0 1 9 13 1 9 2 9 7 10 9 2
41 13 10 9 1 10 9 1 9 0 2 7 9 13 1 9 2 15 4 13 1 10 9 0 1 10 9 0 1 10 9 1 9 7 9 1 10 9 1 10 9 2
12 10 9 1 9 13 15 16 3 9 0 13 2
21 10 9 0 1 10 0 9 13 11 11 2 11 11 2 11 11 2 7 11 11 2
36 10 12 9 0 1 10 11 1 11 2 1 15 2 13 1 9 2 3 10 11 2 1 10 0 9 1 10 16 13 10 9 0 1 10 9 2
33 1 12 4 13 1 10 9 0 10 11 12 2 13 1 11 2 7 1 10 9 11 1 12 9 1 9 15 13 10 11 12 11 2
24 11 13 16 1 10 9 3 13 13 10 9 2 7 13 16 3 2 3 15 13 1 15 2 2
11 3 15 13 10 9 0 2 10 9 0 2
43 1 13 10 9 2 11 7 11 2 11 2 7 11 11 2 11 2 13 1 10 11 2 11 2 11 2 4 13 1 11 11 7 11 11 1 10 9 9 12 2 9 12 2
32 10 9 0 1 10 9 1 10 9 1 11 13 1 12 9 2 1 9 2 0 9 0 7 9 0 2 1 10 9 1 11 2
14 7 10 9 1 10 9 4 13 3 9 1 10 9 2
18 13 10 9 1 12 9 0 2 3 0 2 13 1 10 9 7 9 2
24 3 11 13 1 11 16 13 1 10 11 11 1 10 9 2 9 2 2 13 1 11 1 12 2
14 10 9 13 10 9 2 1 10 9 1 11 11 11 2
27 10 9 13 10 9 3 0 2 16 7 15 13 1 13 1 10 9 0 0 2 0 7 0 2 10 9 2
14 13 1 12 2 11 13 1 10 9 0 3 1 11 2
23 10 9 13 2 7 2 10 9 0 1 16 10 12 13 13 1 16 4 1 13 15 9 2
15 10 9 1 9 15 13 1 10 12 8 8 12 8 3 2
38 3 1 10 9 1 13 2 11 13 13 1 11 1 10 9 7 15 13 1 10 9 1 13 13 1 15 2 13 1 10 9 13 1 10 9 1 11 2
33 2 3 13 10 9 2 13 10 0 9 15 16 13 3 2 7 10 9 4 13 15 7 13 15 2 2 13 11 1 9 1 11 2
22 10 9 13 0 9 7 1 9 3 13 12 9 7 11 13 10 9 7 13 10 9 2
30 15 15 13 9 1 10 9 13 1 10 9 0 2 7 1 10 9 13 1 12 1 12 9 1 13 10 10 9 0 2
44 10 12 1 11 1 12 13 1 10 0 9 1 9 1 2 11 1 11 2 2 10 9 0 1 10 9 11 2 11 1 10 15 15 13 10 9 0 16 13 1 10 10 9 2
15 10 0 11 11 2 15 4 13 1 13 1 11 1 12 2
13 10 9 1 9 13 1 12 8 2 5 5 5 2
39 11 13 10 9 1 12 9 1 9 0 0 13 1 10 9 11 2 0 1 10 9 1 11 2 12 9 2 7 9 1 11 2 10 9 2 11 11 2 2
18 10 9 4 13 1 10 9 1 9 1 9 1 9 13 1 11 11 2
43 11 11 11 2 12 2 12 2 2 13 10 9 0 2 9 1 10 11 11 2 12 2 2 9 0 1 12 9 2 16 13 9 0 0 16 4 13 1 11 1 10 8 2
28 1 9 10 9 13 13 10 0 7 15 9 1 10 9 1 10 9 0 16 13 10 9 1 10 15 16 13 2
62 11 11 11 11 2 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 13 10 9 2 13 7 0 0 16 13 1 10 9 0 2 1 0 1 10 11 7 13 10 9 0 1 0 9 1 9 1 9 0 1 10 9 1 9 1 11 2
27 13 10 9 16 15 13 3 1 10 9 1 9 2 3 15 13 1 10 9 7 1 0 9 1 9 0 2
21 4 13 1 10 9 1 12 1 12 2 7 13 1 9 1 10 11 2 11 11 2
17 15 13 1 10 0 9 2 13 15 16 13 7 15 13 1 13 2
10 3 3 2 13 3 7 13 1 11 2
31 10 9 1 9 4 13 1 9 1 10 9 2 3 9 2 1 10 9 16 15 9 1 9 15 13 10 9 0 1 11 2
5 9 1 10 0 2
17 2 15 13 0 9 1 9 2 9 2 9 7 9 2 2 13 2
32 10 9 16 13 10 9 1 9 13 11 2 10 0 9 0 1 10 9 0 1 9 1 9 7 10 9 1 10 9 1 9 2
27 1 10 9 13 1 15 9 1 10 9 0 13 10 9 1 9 1 9 1 10 9 7 10 9 1 9 2
18 1 11 1 12 2 13 10 0 9 1 10 0 9 13 1 10 9 2
26 11 11 11 1 11 13 10 8 2 0 9 2 9 2 9 7 9 0 13 10 12 1 11 1 12 2
38 15 9 16 13 11 4 13 16 1 9 10 9 16 13 4 4 13 3 13 10 9 16 15 13 3 7 16 3 15 13 1 15 1 9 1 10 9 2
33 1 13 15 1 10 9 7 13 15 10 9 1 13 2 13 10 9 1 13 15 1 9 2 9 16 3 13 15 0 2 16 13 2
23 1 10 9 0 1 10 9 2 3 9 1 11 15 4 13 1 9 7 1 10 9 0 2
13 2 11 2 13 15 1 10 9 3 0 1 11 2
17 1 15 13 10 9 1 11 11 2 16 4 13 10 0 9 0 2
20 1 11 13 3 1 10 0 9 0 1 10 9 11 2 1 10 9 1 11 2
77 3 15 4 7 15 4 13 10 9 0 16 1 10 9 13 10 9 2 10 9 1 10 9 2 15 16 13 0 1 13 9 2 13 2 13 2 13 2 13 13 1 10 10 9 7 1 15 15 16 2 1 9 0 2 13 0 1 13 10 9 1 9 2 13 10 3 0 9 1 9 1 10 9 1 10 9 2
32 15 13 1 10 0 12 2 1 15 15 11 10 11 13 10 9 1 10 9 11 1 11 1 10 9 3 0 1 13 10 9 2
57 1 10 12 9 1 10 11 7 1 10 12 1 10 9 1 3 11 2 15 13 1 9 1 9 7 9 1 10 9 0 1 13 10 9 1 10 9 2 3 1 13 15 9 0 1 10 9 1 10 9 1 10 9 7 9 0 2
12 10 9 15 13 1 10 10 9 1 10 9 2
48 3 2 1 0 13 10 9 1 10 9 0 15 16 13 10 9 16 15 13 1 13 2 7 16 1 10 9 10 9 13 13 3 1 10 9 1 9 0 2 3 3 1 10 0 9 0 2 2
76 13 1 10 11 2 9 11 2 15 13 1 11 1 10 11 11 11 2 3 15 13 1 11 11 16 13 9 1 9 1 10 11 11 1 10 11 2 3 13 10 9 1 9 1 10 9 2 3 3 13 1 10 9 1 11 16 13 9 1 9 1 10 11 11 1 11 2 13 10 9 1 9 1 9 0 2
13 16 13 0 2 3 4 13 1 9 0 10 9 2
30 10 11 11 2 11 11 1 9 2 13 10 9 13 1 10 9 0 11 11 2 1 10 9 1 11 2 11 11 2 2
25 13 10 9 3 0 2 3 0 2 16 10 9 3 13 3 3 2 7 3 13 16 13 1 9 2
34 10 9 13 0 9 2 7 1 15 13 9 1 2 7 15 13 3 2 2 2 3 15 13 2 7 2 13 1 11 2 2 1 15 2
22 1 9 2 10 12 1 11 1 12 2 4 13 1 0 9 0 1 10 9 11 11 2
23 11 13 0 1 11 11 2 11 1 10 9 1 9 1 9 7 0 1 11 11 1 9 2
7 10 9 13 0 2 0 2
41 1 10 12 9 4 13 1 10 9 1 10 11 3 13 12 9 1 12 9 2 1 10 12 9 4 13 1 10 11 11 11 2 13 9 1 10 0 9 11 11 2
10 10 10 9 4 3 13 1 9 0 2
44 10 9 15 13 1 9 1 10 0 9 2 1 10 9 1 2 9 2 7 3 1 9 1 10 12 1 11 1 12 2 10 2 9 2 4 13 1 10 9 1 2 9 2 2
28 11 15 13 10 0 11 1 11 16 13 1 10 9 1 11 7 15 13 16 10 11 1 11 13 10 9 0 2
35 10 9 0 13 1 12 1 15 15 13 10 9 1 0 9 1 9 2 1 10 15 10 9 1 10 9 13 0 3 1 10 9 1 11 2
15 13 1 4 15 13 1 10 9 7 13 0 1 10 9 2
21 1 10 15 2 15 13 10 12 9 16 3 2 11 1 11 2 13 1 10 9 2
15 10 9 13 3 2 1 10 9 0 2 2 1 10 9 2
28 1 3 2 4 13 10 9 0 2 1 10 12 5 0 1 12 7 12 2 7 13 1 12 5 2 1 9 2
19 1 0 16 10 9 1 10 9 2 11 4 13 0 9 1 11 15 13 2
25 1 10 9 15 13 0 9 1 9 2 1 10 15 13 10 9 2 3 7 11 2 10 9 0 2
5 1 15 15 13 2
36 7 13 16 15 13 16 13 1 9 10 0 9 16 13 1 10 9 1 10 9 1 10 9 10 10 9 13 16 10 9 13 0 9 1 9 2
18 15 13 2 1 9 2 16 16 10 9 15 13 2 1 0 15 13 2
22 10 9 13 10 11 1 11 1 10 9 2 13 10 9 1 15 16 3 13 10 9 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
15 15 13 15 10 9 16 13 8 0 7 15 13 8 0 2
32 3 15 13 10 9 1 10 9 1 10 9 2 7 10 9 1 10 9 0 2 13 1 15 16 13 7 15 1 15 15 13 2
45 1 10 9 10 9 1 10 9 0 1 10 11 2 1 10 9 1 9 2 13 9 2 13 1 10 9 0 2 10 9 1 9 7 10 0 9 13 1 9 1 9 1 10 9 2
29 13 3 10 9 0 1 9 1 3 9 7 11 7 10 0 9 1 10 11 11 2 10 9 1 11 3 13 9 2
18 15 13 13 1 10 9 0 1 9 1 10 0 9 1 9 7 9 2
12 11 11 2 9 2 13 1 10 9 1 12 2
16 13 10 9 2 9 1 10 9 1 11 2 11 11 1 11 2
49 1 10 9 1 10 9 1 10 15 10 9 15 13 1 13 1 10 9 2 11 11 13 1 10 9 16 13 1 10 9 15 9 1 10 9 1 9 2 15 16 13 9 1 10 0 9 1 11 2
25 13 16 11 4 4 13 10 9 2 1 15 15 13 1 11 7 15 13 16 10 9 13 3 0 2
40 10 9 15 13 1 10 9 12 2 9 1 10 15 15 13 1 10 9 1 10 2 9 0 2 2 1 10 13 1 10 0 12 9 16 13 10 9 3 0 2
74 13 1 10 9 1 2 11 11 2 2 11 13 15 1 10 9 1 10 9 1 9 16 13 10 9 1 9 1 12 3 13 9 1 10 11 11 7 1 10 11 11 1 10 11 11 11 1 10 11 11 2 11 2 2 10 9 1 9 16 1 10 9 15 13 1 10 0 1 10 9 1 10 11 2
41 10 0 9 2 13 1 10 0 9 0 2 13 10 9 1 11 2 10 9 16 13 1 11 1 10 9 1 13 1 10 9 13 1 10 9 1 10 0 11 11 2
29 1 10 9 1 3 13 10 9 1 13 1 10 9 2 3 4 13 1 10 9 16 15 4 13 1 9 3 0 2
10 13 10 9 3 0 7 13 10 9 2
26 10 9 3 13 9 1 7 4 13 1 10 9 0 1 10 9 2 13 1 9 2 7 9 1 9 2
36 13 1 11 11 7 11 11 2 11 2 13 1 11 11 11 2 11 2 2 11 11 2 11 2 2 11 11 2 11 2 7 11 2 11 2 2
29 3 1 12 9 1 9 3 15 13 9 1 10 9 13 10 9 1 10 0 9 1 12 2 1 10 9 11 11 2
11 2 2 3 13 10 9 1 11 1 11 2
13 2 11 11 11 2 4 13 1 13 10 9 0 2
18 10 9 3 13 3 0 2 7 3 13 10 0 9 1 13 1 9 2
26 10 9 1 9 7 1 9 1 10 9 2 9 0 7 0 2 13 10 9 1 10 9 16 15 13 2
7 13 10 9 1 1 13 2
36 1 10 12 9 1 10 9 4 1 13 10 9 1 10 9 2 1 12 9 2 3 1 10 9 11 11 7 1 10 9 11 11 7 11 11 2
12 15 13 16 13 7 10 9 13 1 0 9 2
14 1 11 13 10 0 9 15 16 13 1 10 10 9 2
19 15 13 1 10 9 0 1 10 1 10 9 0 2 0 1 10 9 12 2
28 10 9 13 0 2 13 13 2 13 9 7 9 2 7 1 10 9 13 0 1 10 9 1 9 7 1 9 2
12 1 10 9 0 2 15 13 3 1 10 9 2
5 13 1 9 0 2
22 1 12 1 11 1 12 10 9 1 10 9 13 1 12 9 2 12 9 7 12 9 2
20 10 9 2 11 2 9 0 11 11 2 2 13 1 11 7 3 4 1 13 2
56 10 9 13 16 3 4 13 0 1 13 2 16 15 4 13 10 9 2 10 9 1 16 10 9 1 10 12 5 1 10 9 4 1 13 10 9 1 10 9 2 7 3 13 3 13 15 2 13 10 12 5 0 10 10 9 2
30 9 12 10 9 1 10 9 15 13 1 11 12 2 1 10 15 13 1 11 1 12 2 16 15 13 1 11 11 11 2
21 10 9 3 9 2 13 1 0 1 10 9 2 4 4 13 3 1 10 9 3 2
8 10 9 13 1 10 0 9 2
17 1 11 11 11 15 9 13 10 12 1 11 1 12 1 11 11 2
10 1 10 9 0 13 3 1 12 9 2
20 9 1 15 2 15 13 9 15 3 4 13 1 10 9 1 9 1 0 9 2
62 1 9 1 15 2 10 9 13 10 9 2 13 15 1 10 2 9 1 9 1 10 11 11 13 1 10 9 0 0 1 10 9 1 10 9 0 2 2 7 3 1 10 2 9 1 9 1 10 11 11 1 10 9 13 1 10 11 1 10 11 2 2
33 10 9 1 10 9 13 9 0 2 13 16 12 1 10 0 9 1 9 1 10 9 15 13 1 10 9 2 11 11 7 11 11 2
30 11 13 1 2 13 10 9 0 2 0 16 13 10 9 2 10 15 2 13 2 3 15 4 1 13 1 9 0 2 2
38 13 9 16 13 1 9 10 9 1 10 9 2 1 10 9 1 10 9 1 11 1 12 7 10 9 1 10 9 1 10 11 11 1 10 9 1 12 2
8 13 10 9 1 9 1 12 2
9 10 9 13 9 1 10 9 11 2
28 10 9 1 10 9 15 13 1 12 1 10 9 0 11 11 2 13 1 10 9 0 1 10 3 9 11 11 2
26 10 9 11 13 1 12 1 10 9 0 1 10 11 1 11 11 1 10 11 11 11 1 11 1 11 2
70 10 9 4 13 1 11 11 2 7 13 1 10 0 9 13 1 15 1 10 9 1 11 1 9 7 0 9 1 10 9 1 10 15 13 2 1 10 9 1 13 9 1 10 9 2 1 10 13 1 9 1 9 7 9 2 13 10 3 0 1 10 9 0 10 9 0 1 11 11 2
37 10 9 11 12 2 1 9 8 2 13 10 9 1 9 1 10 11 1 11 2 10 9 4 13 1 10 9 13 1 10 9 1 10 9 11 11 2
38 10 9 1 10 9 1 10 9 13 3 0 2 3 0 10 0 9 1 0 9 2 1 0 9 2 1 0 9 16 13 1 10 9 1 9 1 9 2
11 10 9 1 11 15 13 13 1 10 9 2
27 1 12 7 12 13 10 9 1 9 0 1 11 2 13 15 1 15 1 10 0 1 13 9 1 10 9 2
25 1 9 2 10 9 1 9 13 16 3 15 4 13 9 0 7 16 3 4 13 15 9 1 15 2
21 10 9 16 10 9 13 10 9 2 15 13 10 9 7 15 13 0 10 9 0 2
25 10 9 0 1 10 11 11 13 1 10 9 1 9 1 10 11 11 11 7 9 1 10 11 11 2
70 3 10 9 3 0 1 10 9 13 10 15 15 4 13 10 9 1 10 9 0 1 11 7 1 11 2 1 10 9 1 11 11 2 1 10 9 1 10 9 10 11 11 1 11 11 2 7 1 10 9 0 2 11 11 2 1 9 1 10 9 1 9 1 10 11 11 1 11 11 2
36 10 0 9 1 9 13 1 10 9 1 0 9 1 10 9 1 11 11 2 16 15 13 0 1 13 10 9 1 9 1 10 11 1 11 11 2
26 13 10 9 16 3 4 13 15 2 3 16 3 13 3 0 13 16 13 1 10 9 0 7 10 9 2
31 1 13 1 11 1 12 2 11 13 16 13 1 13 1 10 9 1 10 0 12 9 1 10 9 1 1 10 9 1 11 2
40 10 11 11 1 10 9 2 8 2 8 2 2 8 2 12 2 2 15 13 1 9 2 15 16 13 1 10 9 1 11 13 15 1 10 9 0 1 10 11 2
35 10 12 1 11 1 10 12 13 10 9 13 1 10 11 11 2 1 10 15 13 12 2 9 1 10 9 1 2 11 11 2 7 0 9 2
15 1 9 2 10 9 1 10 9 0 13 1 10 9 0 2
28 10 9 15 13 1 10 9 0 2 0 1 11 2 1 10 9 1 11 7 13 10 9 1 10 9 1 11 2
15 1 11 7 0 1 9 2 9 7 9 2 9 7 9 2
33 10 9 0 1 10 9 13 3 2 3 1 12 9 0 1 9 2 1 10 16 11 13 1 10 12 7 10 12 5 2 2 13 2
36 10 0 9 10 11 11 1 11 13 3 13 15 10 9 0 1 10 9 7 13 3 1 10 9 0 2 13 1 15 10 9 0 10 0 9 2
20 13 9 0 1 10 9 1 9 1 10 11 11 2 11 2 2 11 2 11 2
56 1 9 7 13 1 0 1 11 3 3 9 15 13 1 10 9 2 10 9 0 15 13 1 10 9 1 10 9 1 11 2 9 3 13 10 9 1 12 9 13 1 12 2 1 10 9 0 1 10 9 1 10 9 1 11 2
30 10 12 1 11 1 12 2 4 13 1 10 11 11 1 10 9 12 2 12 2 3 13 1 12 9 7 13 12 9 2
15 10 9 0 13 1 10 11 11 2 3 13 1 12 9 2
27 10 9 13 3 0 2 13 1 9 0 10 9 7 10 9 1 9 1 9 2 9 2 11 11 2 2 2
34 10 9 1 9 15 13 1 10 9 0 1 13 1 9 1 15 2 1 10 9 13 10 9 1 10 9 1 10 9 0 7 10 9 2
17 16 11 13 2 13 1 11 13 1 10 11 0 3 1 10 9 2
22 10 9 4 13 10 9 1 16 15 13 1 10 9 0 13 9 0 1 10 9 0 2
48 2 3 13 0 9 1 9 16 13 0 9 1 9 1 9 1 10 9 1 11 2 11 7 10 9 1 10 9 1 11 11 1 9 0 1 10 9 1 9 0 2 2 13 11 11 1 11 2
18 15 13 1 10 0 9 1 10 9 2 15 1 10 9 1 10 9 2
62 10 9 13 16 1 13 9 0 1 10 9 4 7 13 10 9 0 2 1 10 15 3 13 2 2 16 13 10 9 1 3 0 9 4 7 13 10 9 0 2 7 1 13 9 0 1 10 9 4 7 13 10 9 0 2 1 10 15 3 13 2 2
16 1 12 10 9 11 1 10 11 7 10 11 13 10 0 9 2
66 1 11 15 15 13 10 9 16 3 13 10 9 2 10 9 1 9 1 10 9 2 10 9 1 10 9 7 10 9 0 2 3 13 11 1 11 1 11 7 3 11 2 7 10 9 2 11 11 2 2 10 0 9 1 10 9 7 10 9 1 10 9 7 10 9 2
17 3 14 1 10 9 1 11 3 15 13 1 10 9 7 10 9 2
39 1 10 9 2 10 9 1 9 4 13 1 9 0 2 16 4 13 1 10 9 0 2 10 9 2 7 9 7 9 1 9 7 9 1 9 0 7 0 2
32 10 0 9 13 1 3 1 7 10 9 4 13 15 13 13 1 10 9 8 11 2 3 10 9 2 16 13 1 10 9 0 2
48 10 0 9 2 1 11 11 11 1 10 9 15 4 13 1 13 15 1 9 1 10 9 1 10 9 1 11 2 4 1 13 10 9 2 3 10 9 1 9 7 10 9 0 1 10 9 12 2
11 15 13 3 3 7 10 9 13 3 0 2
27 10 11 1 3 1 12 9 13 0 2 0 7 0 2 10 9 13 1 10 9 2 9 1 10 10 9 2
27 1 10 9 3 0 2 10 9 0 1 11 15 13 1 9 0 2 1 9 10 9 7 10 9 13 0 2
61 7 3 3 13 1 9 10 9 0 3 2 7 3 10 9 1 9 1 10 0 9 2 13 1 9 16 3 13 1 10 9 1 10 11 10 9 1 11 11 11 2 10 9 9 1 10 11 11 11 11 2 3 7 9 1 9 0 7 9 0 2
22 3 2 10 9 15 13 3 1 9 0 16 13 1 10 9 10 0 9 1 10 9 2
26 9 1 11 11 2 9 1 10 11 11 1 10 9 4 13 1 10 9 0 16 4 13 1 10 9 2
10 11 2 10 9 2 13 1 10 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
36 10 9 1 11 15 13 1 13 10 9 1 9 1 11 11 1 15 15 11 15 13 7 13 16 10 11 13 1 1 15 16 3 13 1 15 2
21 1 11 11 15 13 10 0 9 1 10 9 2 10 9 0 3 0 1 10 11 2
49 4 13 1 10 9 0 1 9 1 12 1 10 9 1 11 11 1 11 11 1 10 9 0 1 10 9 0 2 11 13 10 9 1 9 1 10 9 1 0 9 0 1 15 9 1 10 9 12 2
26 1 9 2 15 13 10 9 1 10 0 8 9 2 15 16 13 1 10 9 13 10 9 1 10 9 2
20 11 13 1 10 9 2 2 13 0 13 1 11 7 13 1 10 11 11 11 2
25 11 2 3 0 13 15 1 9 1 10 9 1 11 2 15 13 1 13 9 1 10 9 1 9 2
14 4 13 1 9 1 8 2 0 2 0 7 0 2 2
34 1 11 11 15 13 10 9 1 9 1 10 9 7 10 9 1 10 9 1 10 9 1 9 1 10 9 1 10 9 7 10 0 9 2
29 1 15 15 13 3 7 15 13 2 7 3 15 13 1 10 9 2 16 0 16 1 10 16 15 13 3 13 0 2
48 10 9 1 10 9 13 1 10 9 0 2 1 10 9 0 1 10 9 1 10 11 2 9 0 7 10 9 11 2 1 10 11 11 2 16 4 13 10 9 1 13 10 0 9 1 9 0 2
83 11 11 7 11 11 2 9 1 10 9 2 13 10 9 1 10 0 9 2 7 13 9 0 1 10 9 7 9 1 10 9 7 9 13 1 10 9 2 15 16 13 10 2 9 2 9 1 10 9 7 9 2 7 1 10 9 0 2 7 15 13 3 1 10 9 2 1 9 2 13 3 10 9 7 9 7 3 13 3 1 15 2 2
42 10 9 1 11 11 4 13 10 2 9 2 16 15 4 13 1 16 3 13 1 10 9 12 9 7 9 1 9 7 16 1 9 3 13 3 1 13 1 11 1 11 2
16 12 9 13 10 0 9 7 11 11 11 13 1 10 11 11 2
28 1 3 2 4 13 10 9 0 2 1 10 12 5 0 1 12 7 12 2 7 13 1 12 5 2 1 9 2
14 4 13 9 1 10 11 11 11 11 11 11 1 12 2
21 10 9 1 9 1 10 9 4 13 1 12 9 1 9 0 1 10 9 1 9 2
18 1 12 2 11 4 13 1 10 11 8 1 12 9 1 9 3 9 2
25 15 4 13 3 3 1 10 9 7 4 13 16 10 9 1 10 9 13 0 1 10 9 16 13 2
18 1 9 1 10 9 0 2 11 13 10 9 1 9 2 3 1 11 2
15 4 1 13 15 1 10 9 1 9 1 10 0 9 0 2
17 10 9 15 13 1 15 0 2 13 11 1 10 0 9 1 9 2
36 13 1 9 10 12 1 11 1 12 1 10 12 9 7 4 13 1 10 9 11 2 11 2 11 1 11 2 1 2 11 2 11 1 10 9 2
43 10 9 1 11 13 1 10 9 1 15 2 1 0 9 7 13 1 10 9 2 2 4 7 13 0 3 7 3 13 10 0 9 1 9 7 10 9 1 10 9 2 13 2
40 11 11 2 2 11 11 2 2 2 13 10 12 1 11 2 13 10 9 3 0 1 11 7 11 11 7 13 3 10 9 3 0 1 10 9 1 10 12 9 2
14 4 1 13 1 10 9 7 13 1 12 5 1 11 2
19 13 3 0 1 16 10 9 15 13 1 16 10 9 4 13 1 15 9 2
35 10 9 1 10 9 13 9 16 4 1 13 3 1 10 12 1 11 1 12 2 7 9 16 15 13 1 10 9 1 13 10 9 1 9 2
13 11 11 11 1 11 2 9 1 11 2 2 11 2
23 10 9 7 10 0 9 4 13 1 10 9 11 11 1 10 11 2 11 1 11 1 12 2
28 13 13 2 10 9 13 9 1 11 11 1 10 9 7 13 10 9 11 1 10 9 11 2 8 7 11 0 2
16 3 1 9 13 10 9 1 12 2 13 1 11 2 8 2 2
8 10 10 9 15 13 1 9 2
11 11 3 13 10 9 1 10 11 11 11 2
32 10 9 1 10 11 13 10 9 0 16 15 13 1 10 9 1 10 9 2 1 10 9 1 11 2 11 7 11 2 11 2 2
20 11 13 10 9 16 15 13 1 10 9 0 1 11 1 10 9 1 10 11 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
19 10 9 0 13 16 12 11 13 16 10 9 1 9 0 13 3 1 10 9
19 10 9 1 10 9 1 9 1 10 15 11 13 13 0 1 13 10 9 2
14 10 12 5 1 10 9 13 9 7 9 1 10 9 2
19 11 11 11 11 2 8 11 2 12 1 11 1 12 2 13 10 9 0 2
16 10 9 13 0 2 0 7 3 0 2 4 13 1 10 9 2
46 10 11 11 13 10 9 1 9 1 12 9 16 13 1 10 11 11 1 10 9 0 2 0 1 12 7 1 4 13 13 1 10 11 1 10 11 11 1 11 11 1 10 11 11 11 2
16 11 11 13 10 9 1 9 1 10 9 11 1 10 9 11 2
11 15 4 4 7 13 10 9 7 13 9 2
39 7 10 9 2 10 9 0 2 13 2 1 10 9 1 11 2 11 7 3 0 2 1 9 1 10 0 9 1 10 9 2 13 3 1 13 1 10 9 2
22 10 13 13 15 1 10 11 11 11 2 9 3 10 9 1 10 9 13 1 12 9 2
16 1 10 9 13 13 10 9 7 13 1 13 10 9 1 9 2
48 10 9 2 1 10 12 16 15 13 2 4 13 1 10 9 1 10 0 9 7 13 10 9 1 9 0 1 10 9 0 15 0 2 1 10 9 2 1 10 9 1 9 7 1 10 9 0 2
16 13 1 11 11 1 11 2 3 1 10 9 1 0 9 0 2
23 8 11 15 13 13 10 9 0 0 1 10 9 2 1 10 0 9 1 9 1 10 9 2
25 1 10 9 2 10 13 9 16 15 13 9 2 3 13 10 9 0 16 8 13 1 10 9 0 8
64 1 10 9 2 12 2 2 1 10 0 9 1 10 2 9 2 2 10 9 0 4 13 16 3 13 0 16 10 9 13 10 9 1 9 2 1 10 9 2 1 13 1 10 9 1 9 2 1 13 10 9 7 1 10 9 1 13 1 9 2 9 7 9 2
24 15 15 13 1 10 2 9 2 1 10 9 1 10 9 2 2 1 10 12 1 11 1 11 2
34 10 9 13 7 15 13 2 16 3 11 13 10 12 5 1 10 11 1 10 9 11 11 11 11 2 0 9 1 11 11 1 10 11 2
51 1 4 1 13 10 9 1 10 9 2 15 1 10 9 16 3 4 13 1 10 9 7 1 10 9 0 13 10 1 10 9 2 10 0 9 1 12 9 1 9 0 16 13 0 0 1 10 9 2 13 2
29 1 11 1 12 2 11 13 10 9 1 9 1 10 11 2 12 9 11 1 9 1 10 11 11 1 10 9 0 2
24 15 2 1 11 11 13 9 1 10 9 1 10 9 2 10 11 2 11 2 1 10 9 9 2
17 1 11 13 10 0 9 1 10 9 11 2 3 1 11 11 11 2
15 10 9 2 8 4 4 13 1 9 1 10 9 1 9 2
42 10 9 4 4 13 1 10 11 1 11 1 13 16 13 0 16 10 9 13 16 13 10 9 0 7 3 13 10 9 0 2 13 13 2 10 9 13 1 5 9 2 2
72 2 3 1 12 9 1 10 0 9 1 10 11 1 11 11 11 2 11 2 1 10 10 9 15 13 10 11 1 10 9 1 10 11 11 1 11 2 11 2 1 11 2 1 10 9 1 13 1 9 1 10 9 0 10 9 1 10 9 1 10 9 7 13 10 9 1 9 1 9 7 9 2
45 10 9 13 16 10 0 9 1 9 13 1 10 9 7 16 13 15 1 0 9 16 3 13 1 13 10 15 3 7 13 10 9 1 9 7 9 1 15 13 15 10 9 1 9 2
15 1 10 9 0 1 10 11 11 12 15 13 1 12 9 2
37 10 9 1 10 9 13 1 16 13 10 9 0 2 1 9 16 13 0 9 1 15 2 13 10 9 0 7 9 2 16 13 10 9 1 9 0 2
24 1 10 9 1 10 9 2 10 9 13 10 9 0 1 2 1 10 15 13 9 7 13 9 2
14 10 9 4 13 0 7 10 9 3 0 1 9 0 2
34 10 9 4 13 1 0 9 1 10 0 9 1 9 1 11 11 1 12 2 3 11 13 9 1 9 7 1 10 15 11 13 10 9 2
19 15 13 1 12 9 1 12 9 10 15 2 13 1 10 9 1 12 9 2
30 15 13 1 13 3 13 1 10 9 1 10 9 1 10 9 2 13 9 0 7 0 1 13 10 0 9 1 10 9 2
20 1 12 13 1 10 9 1 10 9 0 2 1 10 9 1 11 7 11 11 2
11 12 1 10 12 9 13 9 1 10 11 2
11 10 9 15 13 1 10 9 1 10 11 2
50 10 9 1 9 9 1 10 15 4 13 1 10 9 11 2 7 1 10 9 13 1 12 1 12 9 8 1 12 9 2 13 10 9 1 9 1 10 9 1 9 1 10 9 1 10 9 7 10 9 2
64 4 13 10 12 1 11 1 12 7 4 13 1 11 11 2 1 9 15 3 13 10 0 9 2 3 7 1 15 15 15 13 1 11 11 2 16 15 13 16 13 15 1 10 9 1 9 2 7 3 3 11 11 2 15 13 15 3 10 9 1 11 11 2 2
19 10 9 13 15 7 16 13 13 1 10 9 13 9 0 13 1 10 9 2
46 13 10 9 1 11 1 10 11 2 0 9 1 11 7 10 11 2 7 3 10 11 2 1 9 1 10 9 9 1 10 9 2 3 15 13 9 0 2 3 7 3 1 10 9 0 2
34 10 9 13 1 10 9 1 11 1 12 9 13 1 10 9 11 7 1 9 1 10 9 1 9 0 9 2 12 5 8 2 10 11 2
25 0 1 15 0 2 13 3 0 10 9 1 9 0 2 13 13 2 16 15 13 1 9 0 0 2
31 3 1 10 0 9 1 11 11 2 10 9 2 1 10 7 10 9 2 15 4 13 1 10 11 11 7 10 0 11 11 2
13 4 1 13 10 0 9 1 10 11 7 13 0 2
17 10 11 11 13 10 9 0 1 9 1 10 9 7 1 10 9 2
45 13 10 9 1 13 15 1 15 3 0 13 1 10 9 1 9 7 15 1 10 9 0 9 1 10 15 3 9 15 4 13 2 4 13 3 1 10 11 2 11 11 7 10 11 2
50 10 9 0 0 2 11 2 13 3 10 9 1 13 10 9 1 9 1 10 9 0 1 10 9 12 1 11 2 13 10 0 9 16 13 10 9 1 10 9 1 10 9 0 2 16 13 1 10 9 2
25 10 9 3 13 3 3 2 11 11 8 2 7 15 13 1 16 15 13 13 9 3 1 15 13 2
49 1 9 0 2 0 7 0 2 13 12 9 1 10 9 1 10 9 1 9 2 11 2 10 9 11 11 7 11 11 2 16 13 1 10 9 0 13 1 15 1 10 9 1 10 9 1 11 11 2
28 1 10 9 11 7 11 13 13 10 9 1 10 9 1 10 9 11 7 13 1 13 10 9 0 1 10 9 2
28 10 9 1 10 11 13 11 11 1 11 2 7 1 10 9 10 9 15 13 1 10 9 0 1 11 7 11 2
16 10 11 11 13 10 0 9 1 10 9 1 9 0 11 11 2
62 1 10 12 9 2 10 9 1 11 13 0 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 9 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
22 3 2 11 15 13 1 13 10 9 1 12 9 0 1 10 9 0 2 1 10 12 2
37 10 9 4 13 1 0 9 1 10 9 11 11 1 11 11 11 1 10 11 2 11 2 11 1 10 11 2 11 11 2 11 7 11 7 11 11 2
7 13 1 9 0 7 0 2
35 11 7 11 2 13 16 10 9 1 10 9 2 11 2 4 13 1 11 11 11 11 2 10 9 1 9 1 10 0 9 1 9 2 11 2
50 1 9 1 10 0 9 16 13 1 11 1 10 0 9 1 10 9 11 11 7 0 9 1 10 9 1 10 9 2 10 9 0 2 11 11 2 13 16 3 13 10 9 1 10 9 0 1 10 9 2
24 3 1 11 11 13 1 4 13 2 3 1 10 9 0 1 13 10 9 0 0 7 10 9 2
7 1 10 0 9 15 13 2
26 10 12 5 1 10 10 9 4 13 1 10 0 9 7 12 5 13 1 10 9 1 3 1 12 9 2
22 7 16 10 9 13 0 1 16 10 9 4 13 1 9 10 9 0 13 1 10 9 2
55 10 9 1 15 13 1 10 9 1 16 15 13 13 10 9 1 11 7 3 10 1 10 9 0 1 9 1 9 7 10 9 13 3 0 2 13 0 16 10 0 9 3 4 13 1 12 9 13 1 15 1 12 9 0 2
17 10 9 0 2 13 11 7 11 4 13 10 11 2 12 2 12 2
27 15 1 10 0 9 13 1 10 9 1 10 9 3 0 1 10 9 1 13 1 10 9 1 10 0 9 2
10 10 9 0 1 10 9 15 13 0 2
22 13 1 10 9 0 2 9 7 9 1 10 9 2 0 2 9 7 9 2 1 11 2
27 11 11 2 9 0 1 0 9 1 11 11 2 4 13 13 10 9 1 9 7 13 15 1 10 0 9 2
9 2 15 13 10 9 7 10 9 2
11 15 13 10 11 10 11 7 10 11 11 2
20 11 11 13 10 9 1 9 1 10 9 1 10 11 1 10 9 1 10 11 2
54 10 11 13 10 9 0 1 11 1 10 13 3 1 12 9 1 10 9 8 12 9 1 10 9 2 1 10 9 1 16 13 1 10 9 0 16 13 10 9 7 10 9 2 0 2 1 10 9 0 16 13 10 9 2
18 3 13 10 9 1 10 9 1 11 1 11 11 7 10 9 1 11 2
18 3 4 13 9 1 10 9 1 9 3 1 10 9 0 7 13 9 2
32 10 9 1 11 15 13 0 1 10 9 1 10 9 0 1 11 1 10 9 0 1 10 11 1 11 1 10 9 1 12 9 2
33 11 2 3 1 11 2 12 2 12 2 11 2 13 10 9 0 2 9 7 9 1 10 11 11 1 11 2 3 13 1 12 9 2
6 13 0 1 10 9 2
30 11 11 13 10 9 1 9 0 2 1 10 9 0 2 3 1 3 1 10 9 1 0 2 7 10 9 0 7 9 2
34 10 9 1 9 13 10 9 0 7 9 1 9 1 10 9 0 0 7 0 1 10 9 0 7 0 2 13 10 9 1 9 1 9 2
21 1 11 10 9 0 15 13 0 1 10 9 3 0 1 11 2 1 10 9 0 2
23 10 9 0 2 11 11 2 15 13 0 1 10 9 0 3 15 9 10 9 1 9 0 2
16 10 11 13 10 9 0 0 16 13 10 12 1 11 1 12 2
24 0 9 10 9 3 0 2 1 10 9 2 13 10 13 1 10 9 0 11 1 10 9 0 2
86 10 0 9 3 13 1 10 9 1 3 15 13 1 10 9 1 10 9 1 16 10 9 0 13 1 10 9 2 10 9 13 13 1 15 16 15 4 4 1 13 2 10 9 1 10 9 0 2 2 9 7 9 1 10 9 0 13 1 10 9 10 4 13 10 0 9 1 9 2 13 15 1 3 1 10 9 0 2 9 13 3 1 10 11 11 2
36 10 9 13 10 9 2 16 13 1 10 12 1 10 12 2 15 13 16 10 9 13 1 11 10 9 1 10 11 1 10 11 2 9 1 11 2
12 11 11 2 1 9 0 11 11 7 11 2 2
10 10 9 4 13 1 0 9 1 12 2
6 3 15 13 10 9 2
39 11 11 15 13 1 11 16 10 9 1 2 11 11 2 13 10 9 16 15 13 1 10 9 2 16 2 3 15 16 13 1 11 4 13 15 1 11 2 2
22 1 10 9 2 10 9 0 1 10 12 1 11 1 12 13 10 0 9 1 10 9 2
58 1 10 9 2 15 13 1 10 9 1 10 0 9 2 13 1 10 9 0 1 0 9 2 9 1 15 15 13 1 16 11 13 16 10 9 15 13 1 10 9 3 10 9 13 1 10 9 0 1 10 9 1 9 2 9 7 9 2
19 1 3 13 10 9 2 10 9 1 11 13 13 1 10 9 1 10 9 2
6 13 9 1 10 9 11
25 15 13 1 10 0 9 13 2 2 8 8 8 8 8 8 8 8 2 8 8 8 8 8 8 2
28 2 13 16 10 9 13 10 9 1 10 9 7 15 13 10 9 1 9 3 0 2 2 13 10 9 0 13 2
43 10 9 1 10 9 4 13 1 13 1 15 7 1 15 13 10 9 0 2 1 10 9 1 10 9 2 1 11 7 11 2 7 15 4 13 10 11 1 11 1 10 9 2
10 10 9 2 11 11 15 13 10 9 2
8 10 9 4 13 0 7 0 2
25 9 1 10 9 1 10 9 3 15 13 0 1 9 1 10 9 7 10 11 9 1 10 9 0 2
10 1 10 11 1 11 13 0 10 9 2
32 1 10 9 13 0 2 10 9 2 10 11 1 11 1 11 11 1 10 11 11 2 11 2 7 11 1 11 8 2 11 2 2
19 13 10 9 1 15 3 15 4 13 2 1 10 9 7 1 10 9 3 2
119 15 13 1 11 1 12 2 7 15 15 13 10 9 1 10 9 1 10 11 2 7 1 0 1 10 9 0 11 1 11 2 12 2 2 13 1 9 11 11 2 12 2 2 9 0 7 9 0 2 1 10 15 13 16 11 1 11 13 0 1 10 9 0 1 10 9 2 16 13 2 13 0 7 0 1 15 2 7 13 1 10 9 1 0 2 2 3 7 2 1 4 13 9 1 9 0 7 0 1 10 10 9 2 1 9 1 9 2 9 7 9 2 2 9 16 13 3 0 2
23 13 10 9 7 9 7 10 9 13 1 10 9 1 10 9 7 1 10 9 1 10 9 2
18 1 0 16 10 10 9 2 11 11 11 13 0 9 13 1 10 9 2
11 10 9 1 10 9 0 13 1 12 5 2
20 13 1 9 7 10 0 9 13 8 8 8 8 1 10 8 8 8 8 8 2
11 15 3 13 10 9 3 0 1 10 9 2
51 10 9 4 13 1 10 9 1 11 2 16 13 10 9 1 10 9 0 1 0 2 13 10 9 1 12 9 13 1 12 9 1 9 2 1 10 9 12 9 13 10 9 3 3 1 10 9 1 10 9 2
56 13 10 10 9 3 1 10 9 1 11 2 1 12 9 2 3 16 10 9 4 13 1 9 1 9 7 1 10 9 3 0 2 0 2 0 2 9 2 10 11 1 11 13 10 9 1 12 7 13 1 0 9 11 1 11 2
26 16 1 10 11 3 13 9 10 2 11 13 12 7 12 9 1 9 2 9 2 9 2 9 7 9 2
19 13 10 9 1 10 8 0 13 10 9 1 13 1 10 9 1 0 9 2
21 10 9 4 1 13 7 16 4 13 0 13 2 1 10 9 0 1 11 7 11 2
33 16 10 9 4 13 10 9 1 10 11 11 4 13 15 1 10 9 3 0 7 0 1 11 9 0 7 0 1 10 11 11 11 2
46 11 12 1 9 9 1 10 9 2 13 13 1 15 1 10 0 2 2 13 1 9 1 9 2 7 13 1 9 0 7 9 2 15 16 13 9 7 10 9 1 10 9 1 10 9 2
12 3 13 16 13 0 16 3 4 13 3 8 8
21 10 9 13 0 1 13 16 3 11 15 13 1 9 2 7 3 7 1 9 0 2
8 11 15 13 13 1 10 9 2
14 1 10 9 13 11 11 2 13 11 11 2 9 2 2
13 10 9 13 3 1 9 0 1 9 7 9 0 2
5 10 9 13 0 2
29 12 9 3 11 13 10 9 1 10 9 1 10 15 15 13 10 2 9 7 10 9 1 9 2 1 10 9 0 2
18 10 9 13 10 9 0 1 5 12 9 1 10 5 12 1 10 9 2
11 13 1 12 3 13 10 0 9 1 9 2
40 10 9 2 13 1 10 9 11 11 11 2 13 16 10 9 13 10 0 9 1 10 9 3 1 3 12 9 1 9 1 9 0 7 15 13 1 10 9 0 2
36 13 10 10 9 2 0 1 10 7 10 9 2 7 16 3 13 1 10 9 13 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2
23 10 9 1 10 9 3 13 9 1 9 1 10 0 9 1 9 1 10 9 1 10 9 2
29 11 7 11 9 1 11 1 12 2 12 1 9 1 10 9 11 1 11 2 12 12 1 11 1 11 2 1 12 2
4 13 9 0 2
30 10 12 1 11 9 1 9 15 13 1 10 12 8 16 13 9 1 10 9 2 3 1 9 10 9 7 0 1 12 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
28 10 9 4 13 1 9 0 2 1 9 16 10 9 1 15 13 3 10 0 9 1 10 9 0 1 10 9 2
22 3 1 10 9 1 10 9 2 3 15 4 13 10 0 9 1 10 9 1 10 9 2
25 15 13 1 10 9 1 10 9 2 16 4 1 13 1 10 9 1 10 9 13 0 9 1 9 2
10 3 13 10 11 11 1 11 1 12 2
31 3 13 10 9 1 10 11 2 11 3 0 1 10 9 1 9 0 2 16 13 12 9 1 11 1 12 9 7 12 9 2
22 10 9 1 10 0 9 0 13 10 9 2 11 2 11 11 11 11 11 2 1 11 2
39 10 9 1 9 3 2 1 10 0 9 1 10 9 2 11 13 1 10 9 1 10 9 1 7 2 11 2 13 1 10 9 1 10 9 0 2 12 2 2
37 7 16 4 13 15 4 13 1 9 1 13 9 2 13 1 9 3 0 7 13 9 1 9 1 10 9 1 9 1 0 9 16 15 13 3 3 2
19 10 9 13 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
20 3 2 15 16 4 13 10 9 1 10 9 4 13 10 9 1 10 9 2 2
9 1 9 1 9 13 10 0 9 2
30 10 0 9 13 10 9 0 10 11 0 2 1 11 11 7 11 11 1 10 9 1 10 9 1 9 3 13 11 11 2
37 10 9 1 9 2 9 4 3 13 1 10 0 9 0 2 7 3 15 13 1 10 12 9 1 10 12 9 1 10 9 0 2 16 13 1 11 2
14 10 15 13 3 13 9 1 15 3 13 2 7 9 0
24 15 13 10 9 1 9 7 15 4 13 3 3 2 1 3 0 9 2 13 1 10 9 2 2
16 10 9 15 4 13 1 10 11 1 13 10 0 9 1 11 2
34 15 1 10 0 9 0 1 11 7 11 4 4 13 1 11 2 13 10 9 0 1 11 11 11 2 11 11 2 11 11 7 11 11 2
30 1 12 2 13 1 10 9 0 1 11 2 11 15 13 10 9 1 10 9 1 9 3 16 4 13 10 9 1 9 2
13 11 13 3 13 15 1 10 9 16 15 4 13 2
27 13 3 13 10 9 1 10 9 11 11 1 10 0 9 2 7 3 1 15 1 10 9 1 10 9 12 2
19 11 13 10 11 7 15 13 1 13 1 11 11 11 11 1 10 9 12 2
28 10 9 2 1 9 0 11 2 13 1 12 1 12 9 1 10 9 16 13 1 10 9 1 10 9 7 3 2
24 9 3 11 13 10 9 7 13 11 11 11 11 2 8 2 10 11 1 11 2 1 10 9 2
20 4 13 1 12 9 1 12 9 2 13 15 1 10 9 0 10 9 1 9 2
21 1 12 2 13 1 11 1 10 9 0 2 7 1 11 2 1 11 1 12 9 2
21 13 1 11 2 4 13 1 10 9 11 7 13 10 9 10 12 1 11 1 12 2
68 1 12 15 13 10 11 0 1 10 9 1 10 9 1 10 9 1 11 7 0 9 13 1 10 9 2 11 2 2 16 1 10 9 12 13 1 10 13 1 10 9 2 1 9 1 10 13 1 10 9 1 11 2 3 1 9 2 13 10 11 1 11 3 1 9 1 9 2
14 10 9 4 13 1 11 1 10 9 0 11 11 11 2
10 7 16 15 1 10 9 0 15 13 2
23 10 9 0 11 13 10 9 1 2 9 1 10 9 2 7 2 10 9 1 10 9 2 2
25 10 8 9 0 11 8 11 13 16 13 1 10 9 11 11 1 13 15 1 10 9 1 11 11 2
23 1 10 9 2 10 9 15 13 2 7 11 13 16 4 1 4 13 2 10 0 9 2 2
13 3 15 13 9 1 9 0 7 9 1 9 0 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
17 11 11 11 11 13 10 9 0 1 10 9 1 11 11 11 11 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
11 10 9 1 9 0 7 1 10 9 0 2
15 13 10 9 13 1 0 9 7 1 15 3 4 13 15 2
25 15 13 1 10 9 1 10 9 16 15 13 1 10 9 0 11 2 11 2 12 16 13 1 11 2
23 1 12 13 10 11 1 10 11 2 10 9 1 0 9 1 9 1 9 1 9 7 9 2
44 10 9 0 2 1 9 0 7 9 0 2 15 13 1 9 1 9 2 13 1 9 2 1 9 0 3 0 2 13 1 10 9 7 1 10 9 1 10 15 1 10 12 9 2
14 10 9 13 0 9 1 15 16 3 13 11 7 11 2
22 3 2 1 7 10 9 13 0 2 10 9 13 1 9 10 9 1 2 11 11 2 2
33 11 11 11 2 11 2 11 2 12 1 11 1 12 2 2 13 1 11 11 2 13 10 9 0 16 13 1 10 9 1 9 0 2
21 13 1 0 10 9 9 2 1 15 10 9 1 9 7 1 9 16 13 1 11 2
25 10 9 0 1 10 9 0 7 0 7 1 9 1 13 9 0 1 10 9 1 11 7 1 0 2
18 13 1 16 15 13 10 9 16 13 10 9 7 13 13 15 1 15 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
21 16 13 0 2 13 0 1 15 8 1 10 9 16 9 1 10 9 1 9 0 2
41 10 12 9 0 13 2 10 0 9 1 9 1 11 2 10 0 9 1 10 0 7 0 9 0 2 13 12 9 3 0 1 9 2 9 2 10 11 1 11 2 2
18 10 9 13 10 0 9 1 10 9 2 7 15 13 3 3 15 13 2
28 1 10 0 9 2 10 9 15 13 1 10 9 1 10 9 1 10 9 0 7 0 2 7 3 3 1 15 2
23 13 1 11 2 13 13 15 2 7 4 13 1 10 9 1 9 11 1 13 1 0 9 2
31 9 1 10 9 2 11 4 13 1 9 1 9 0 7 0 1 10 9 1 10 8 9 1 10 11 1 11 11 11 11 2
14 10 9 13 3 10 9 1 10 9 1 11 7 11 2
26 3 13 9 2 13 9 1 9 1 9 0 7 9 1 10 9 1 9 7 9 1 10 9 1 11 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 5 12 2 1 10 15 12 5 12 4 1 9 0 7 2 12 5 2 12 5 12 13 9 2
32 15 3 13 1 2 11 2 2 10 9 1 10 11 1 10 11 2 16 11 15 13 1 13 16 11 4 4 13 1 10 9 2
14 2 11 13 15 1 15 0 7 13 1 10 9 0 2
38 10 9 13 1 10 9 10 9 0 7 10 13 2 3 1 10 9 0 1 10 9 1 10 9 1 10 9 1 10 0 11 11 11 1 11 1 11 2
23 11 15 13 3 2 10 9 0 7 0 7 10 9 1 10 9 13 1 15 10 9 0 2
35 11 11 11 2 9 1 9 2 13 16 3 10 0 9 15 13 1 13 10 9 1 9 1 10 9 2 9 1 10 9 7 9 1 10 9
22 10 9 4 13 1 11 11 12 2 10 11 11 9 0 9 1 11 11 7 11 11 2
14 10 9 1 10 9 13 0 7 10 9 3 13 3 2
80 3 2 1 9 1 10 9 1 9 1 10 11 11 2 11 7 10 9 1 10 9 1 10 16 13 10 9 1 0 9 2 11 11 13 10 0 9 1 10 9 11 11 1 11 7 13 10 9 1 11 1 10 9 1 9 1 10 0 9 11 7 10 9 1 10 9 1 11 1 11 1 10 0 8 1 9 1 10 11 2
24 10 9 1 9 13 10 9 1 9 1 16 13 10 9 1 13 9 7 13 9 0 2 0 2
32 9 1 10 9 13 10 9 1 10 9 2 10 9 2 10 9 0 2 9 0 2 1 10 9 1 10 9 13 1 10 9 2
10 4 13 9 1 11 11 7 11 11 2
19 13 12 9 7 15 13 1 10 9 0 2 1 10 9 7 9 1 9 2
19 9 9 1 10 9 12 13 0 10 9 7 10 11 1 10 12 9 0 2
48 10 9 1 10 15 4 13 10 9 13 1 13 2 9 2 13 0 1 9 1 10 9 7 9 1 10 9 2 7 4 13 1 10 9 1 9 1 9 2 1 13 10 9 1 10 9 0 2
21 1 12 9 15 13 7 15 13 1 10 9 1 8 1 7 15 13 1 13 15 2
17 10 0 9 2 10 9 11 13 1 11 10 12 1 11 1 12 2
49 1 9 1 10 9 7 9 1 9 0 1 10 16 15 13 9 0 1 10 9 0 7 0 1 10 9 0 2 11 4 13 10 9 1 10 9 0 1 9 11 2 16 13 10 9 0 7 0 2
31 10 9 0 13 10 9 1 10 9 13 1 10 9 2 15 10 9 13 1 9 1 11 1 11 2 9 1 11 7 11 2
23 1 10 9 1 10 9 11 13 13 15 3 2 3 3 10 9 1 10 9 13 13 15 2
38 11 11 2 11 2 11 2 13 10 1 11 11 2 11 11 7 13 10 1 11 11 2 11 2 13 10 9 1 9 0 16 13 10 9 1 10 11 2
13 10 9 1 9 13 1 12 8 2 5 9 5 2
41 3 13 9 7 9 1 3 10 10 9 2 13 1 10 11 11 11 1 11 2 16 13 10 0 9 1 10 9 0 7 0 9 1 10 9 1 13 10 9 0 2
31 10 12 9 13 1 0 9 1 10 9 1 9 0 1 10 9 11 2 15 1 10 0 9 1 10 11 1 10 9 11 2
21 10 9 11 13 1 10 9 13 10 12 9 1 9 7 11 13 1 10 0 9 2
5 10 11 2 12 2
25 1 9 2 16 10 9 11 11 15 13 1 10 9 2 13 16 10 12 9 4 1 13 1 12 2
18 10 9 13 10 9 0 1 12 5 9 1 10 12 5 1 10 9 2
42 3 15 13 10 9 1 10 9 1 12 12 9 2 3 0 2 10 0 9 1 10 9 13 2 1 9 1 10 0 9 1 10 9 2 13 10 9 1 10 9 0 2
16 13 9 1 11 11 11 1 11 1 10 11 7 11 1 11 2
32 4 1 13 2 1 9 7 3 13 1 13 15 7 7 13 10 9 3 2 3 7 2 13 1 15 3 1 12 9 1 11 2
12 1 9 12 13 1 10 9 1 12 12 9 2
24 3 15 13 10 9 1 13 15 3 1 9 7 4 13 10 9 1 10 9 0 16 13 3 2
11 11 15 13 3 7 13 10 9 1 11 2
57 2 1 9 4 7 13 16 13 3 0 13 1 11 1 10 9 2 7 1 10 9 1 10 9 2 2 4 13 1 9 1 10 9 11 2 11 2 1 13 10 9 1 9 1 10 11 1 10 11 11 1 10 11 2 11 2 2
17 10 9 13 0 9 1 9 7 1 0 13 10 9 1 9 0 2
15 10 11 1 11 13 10 9 0 16 13 9 0 1 9 2
34 10 9 1 10 9 11 15 13 1 10 9 11 1 10 0 9 1 11 16 13 0 1 10 9 1 10 9 1 10 9 1 10 11 2
34 2 10 11 1 10 11 11 2 13 10 0 0 9 1 10 9 0 1 9 11 2 10 9 1 11 7 10 0 9 1 10 0 9 2
26 1 10 0 9 3 13 1 10 9 2 11 2 1 9 1 10 9 0 2 8 2 8 2 11 2 2
14 10 9 4 13 1 10 9 3 0 10 9 13 0 2
52 10 9 1 10 9 7 1 9 1 10 15 1 9 7 1 9 16 15 13 1 10 9 1 9 1 13 10 9 16 13 7 3 13 15 1 10 9 3 1 10 9 1 10 9 2 3 1 10 9 1 9 2
76 1 10 9 0 0 2 16 13 10 0 9 0 2 10 9 0 13 10 9 0 7 10 9 3 1 9 7 11 2 1 10 9 0 7 0 0 2 16 13 1 10 11 11 11 7 1 10 11 11 2 3 1 10 9 0 1 9 2 15 4 13 10 9 1 10 11 7 1 10 9 0 2 11 11 2 2
30 3 1 10 9 1 9 2 13 1 10 9 10 9 7 1 10 9 0 2 7 1 10 9 3 13 10 11 11 11 2
3 13 0 2
37 11 11 11 2 11 11 2 2 10 0 9 9 1 11 2 11 2 2 13 10 9 1 13 15 1 10 11 1 10 12 9 1 13 10 9 0 2
30 12 9 1 10 11 4 13 9 1 10 9 2 7 1 10 9 0 1 12 2 10 11 13 9 1 9 1 10 11 2
11 15 13 1 11 2 11 2 11 7 11 2
10 10 9 13 15 16 15 13 1 13 2
16 13 10 11 11 1 11 11 2 9 1 9 0 1 10 9 2
16 9 0 3 13 2 0 9 1 9 2 7 3 13 1 9 2
14 10 9 13 10 8 1 10 9 1 10 12 1 11 2
11 1 10 9 12 13 10 9 1 12 9 2
8 11 11 2 2 9 7 9 2
18 10 9 13 9 0 1 10 10 9 7 9 1 9 3 1 10 9 2
10 9 2 10 9 0 2 15 0 2 2
22 1 11 13 10 9 9 1 10 9 2 11 11 11 2 1 10 9 1 10 9 11 2
44 2 9 1 9 1 11 11 13 11 1 9 16 13 15 7 13 1 10 9 7 9 2 10 15 13 10 9 0 1 10 9 1 11 11 2 2 13 11 1 10 9 1 9 2
59 10 9 1 11 13 1 10 9 10 9 13 15 16 13 10 9 1 11 1 10 9 1 15 13 3 10 9 1 10 9 7 3 2 1 0 9 2 15 13 1 10 9 0 1 11 1 9 1 16 13 10 9 0 2 9 16 13 0 2
32 1 10 9 0 10 9 0 1 12 9 1 9 13 3 1 12 9 1 11 10 15 2 7 3 10 9 0 9 3 1 9 2
80 10 9 13 1 10 9 0 3 1 10 12 2 3 1 10 9 0 2 13 1 10 9 1 3 13 8 2 13 10 9 11 11 2 15 1 10 9 1 10 5 0 2 7 10 9 11 11 2 9 1 11 11 16 1 12 9 13 3 10 9 2 1 10 9 0 16 2 9 13 2 13 1 9 16 10 9 13 1 11 2
25 10 9 13 1 10 9 2 9 2 9 7 9 2 7 3 1 10 9 1 10 9 1 10 9 2
34 10 9 0 2 3 10 0 2 13 10 0 9 7 10 9 15 13 1 10 9 0 2 1 10 15 13 9 1 10 10 9 1 11 2
20 10 9 1 11 11 11 15 13 1 10 11 11 2 1 3 1 11 7 11 2
6 10 9 13 1 11 2
36 10 12 9 0 1 10 9 2 3 13 10 11 11 11 2 4 13 1 9 1 10 9 0 1 10 9 0 2 16 13 10 9 1 10 9 2
19 1 10 9 2 11 15 13 9 1 9 1 10 15 7 13 15 3 0 2
33 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 13 10 9 1 9 0 16 13 1 10 9 1 11 11 1 10 11 2
43 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 2 0 9 15 4 1 10 9 13 1 10 9 1 10 9 2 9 13 1 10 9 1 10 9 7 10 9 2
38 10 9 13 10 9 0 1 11 2 9 1 9 11 1 10 11 7 1 13 1 9 9 13 15 1 10 12 2 12 2 12 2 12 2 12 7 12 2
30 10 12 9 1 11 1 10 11 11 2 12 11 2 11 2 11 2 13 10 9 0 1 10 11 1 10 11 11 11 2
29 1 10 9 0 1 10 9 0 2 0 2 12 2 7 1 10 9 0 2 0 2 12 2 13 10 9 1 9 2
19 1 10 9 15 16 13 3 1 10 9 1 10 9 7 1 10 9 0 2
32 10 11 11 11 11 13 10 9 0 1 10 12 9 1 9 16 13 9 0 1 10 9 1 11 2 11 2 1 0 9 0 2
34 10 9 1 10 9 2 2 11 11 2 2 2 10 9 13 2 2 4 13 1 10 9 1 10 0 9 2 1 12 2 1 11 11 2
24 11 2 9 1 10 9 1 9 0 10 9 2 13 10 0 9 1 10 0 9 1 10 9 2
14 10 9 11 11 4 13 10 12 1 11 1 10 12 2
9 13 10 9 1 10 9 1 15 2
39 13 1 9 13 1 10 9 2 15 13 16 1 10 9 10 9 4 13 15 16 13 9 2 13 10 0 9 16 15 13 10 9 0 1 10 9 16 13 2
40 13 1 9 0 2 1 10 0 9 16 10 9 2 7 1 10 9 0 15 13 10 9 1 11 11 2 9 0 2 3 1 9 0 1 9 1 10 9 12 2
62 3 10 9 1 10 9 13 0 2 16 13 0 1 13 7 15 13 9 0 2 7 15 1 10 9 3 2 16 13 10 9 3 0 1 10 9 2 16 13 9 1 10 9 2 7 1 10 9 7 10 9 2 13 15 10 9 1 10 9 0 0 2
13 11 12 13 10 9 0 0 1 10 9 1 11 2
52 11 7 11 2 1 9 8 2 1 8 2 9 2 9 7 1 8 2 0 2 9 2 2 9 15 13 10 9 3 0 1 9 13 1 10 9 7 9 1 10 11 11 2 15 1 10 0 9 13 10 9 2
10 10 9 15 13 3 3 1 10 9 2
8 9 2 11 11 12 11 11 2
47 13 1 11 12 7 1 10 9 11 11 11 12 9 7 10 9 0 0 2 10 0 9 1 10 9 13 1 12 9 2 10 9 11 7 10 11 2 1 10 9 1 12 7 12 9 3 2
43 10 9 1 9 0 2 1 0 1 9 1 10 9 1 0 9 2 3 15 4 13 1 10 9 1 9 1 10 9 2 16 13 0 16 15 3 13 10 9 0 1 9 2
21 10 0 9 0 13 10 9 1 10 9 0 7 1 10 9 0 1 9 1 9 2
26 10 9 1 10 9 15 13 3 7 10 9 13 15 16 4 13 15 1 10 9 1 9 7 9 0 2
26 11 11 11 2 11 11 2 7 10 9 2 10 11 4 13 1 13 11 10 9 3 1 10 0 9 2
28 10 11 2 10 9 13 10 9 1 10 9 16 3 15 13 7 13 10 9 1 11 2 1 10 9 1 11 2
10 10 9 0 3 0 7 13 1 11 2
60 1 10 9 8 1 10 9 2 15 13 16 15 13 9 1 9 2 7 16 13 10 9 1 10 9 1 10 15 11 13 10 9 2 10 9 7 9 16 13 10 9 13 7 13 1 0 9 2 15 13 13 1 10 9 1 16 15 13 3 2
33 10 9 4 13 9 1 9 9 1 9 1 11 1 10 9 7 9 1 11 2 3 16 15 13 10 9 1 10 9 3 0 2 2
22 1 11 2 11 2 10 9 0 3 4 13 3 9 0 13 1 10 9 7 9 0 2
25 13 10 9 1 10 9 2 10 9 7 10 9 2 13 9 7 0 9 13 1 9 7 9 0 2
42 15 13 10 0 9 1 9 16 15 13 1 10 9 3 9 1 12 9 1 9 2 1 9 1 12 9 7 1 10 9 1 10 9 1 11 2 11 2 7 1 11 2
44 1 10 9 1 10 11 12 1 11 1 12 2 10 0 9 1 10 9 0 1 11 11 1 11 13 1 9 10 9 7 10 9 1 10 9 1 10 11 1 11 2 11 2 2
19 4 13 1 10 0 9 1 9 1 11 11 11 11 1 10 9 0 11 2
34 1 10 0 9 2 15 13 16 10 9 4 13 1 10 9 1 11 11 11 2 13 16 3 11 13 10 9 3 0 1 10 9 0 2
67 3 2 13 9 1 10 9 11 11 2 9 1 10 9 1 10 9 11 2 9 1 10 2 11 11 11 11 11 2 2 9 1 10 2 11 11 11 11 2 2 9 0 1 10 2 11 11 11 11 2 11 2 2 7 9 1 10 9 0 1 10 11 1 11 7 11 2
46 10 11 11 13 10 9 1 11 1 12 1 11 1 12 1 10 9 2 15 13 1 9 0 3 1 10 9 2 7 13 1 10 9 3 0 1 10 9 7 10 9 1 11 1 12 2
41 13 10 9 4 13 1 0 2 1 10 9 1 10 11 11 2 1 11 2 13 3 10 0 9 2 11 2 9 9 16 4 13 15 1 2 11 1 10 11 2 2
24 10 9 0 1 11 13 16 10 9 0 4 13 10 9 1 11 1 10 9 1 10 9 0 2
25 13 9 1 10 0 9 7 9 2 15 15 13 3 3 1 11 2 3 16 13 10 0 9 2 2
25 1 15 9 2 3 13 0 9 1 10 9 1 10 9 2 1 15 1 3 1 10 9 1 9 2
23 1 10 9 3 13 2 0 13 13 10 9 1 10 0 9 11 2 7 10 9 3 13 2
20 15 13 1 11 2 10 9 1 9 0 7 13 0 16 13 1 10 11 11 2
24 10 9 1 10 9 13 3 0 2 15 13 1 10 9 1 10 9 10 0 9 1 10 9 2
76 3 1 12 15 13 1 0 9 10 9 1 9 2 10 9 11 11 13 1 10 9 13 10 0 9 1 10 9 15 13 2 10 9 11 2 0 9 1 10 11 2 4 4 13 1 9 2 2 7 1 11 1 11 2 10 0 9 2 0 2 10 9 16 4 1 13 1 15 2 1 13 9 2 13 9 2
14 1 10 9 0 13 10 9 0 1 10 11 1 12 2
93 10 9 1 10 11 13 13 1 10 0 9 1 10 9 0 7 1 9 2 15 1 10 9 0 7 0 2 3 1 10 9 3 0 2 1 10 9 1 13 1 10 9 1 10 9 2 9 1 10 9 7 9 1 0 2 16 4 13 7 13 10 3 0 7 0 9 7 9 2 13 7 13 3 1 10 8 2 3 7 13 10 0 9 1 9 1 0 9 15 0 7 0 2
39 2 1 13 10 0 9 16 13 1 10 9 2 10 9 1 11 4 4 13 3 1 9 1 13 1 10 11 1 10 9 1 10 9 2 2 13 10 11 2
11 13 1 10 11 1 10 11 11 1 11 2
22 13 1 10 9 1 3 13 10 9 2 11 13 7 13 1 11 7 1 10 9 11 2
19 10 9 0 1 10 9 4 13 1 9 2 1 9 1 10 9 12 2 2
14 1 9 1 10 12 1 10 12 13 10 12 7 3 2
38 3 13 10 9 2 13 16 1 12 10 9 1 11 2 1 10 9 1 11 7 11 2 1 10 9 1 10 12 1 11 2 13 3 10 9 10 9 2
8 15 1 15 13 10 9 0 2
18 15 15 13 13 10 9 1 10 11 1 10 9 1 11 2 7 13 2
5 15 13 1 11 2
47 10 9 13 16 10 12 5 1 10 9 0 4 1 4 13 1 9 0 2 2 1 9 7 9 0 1 10 0 9 2 2 1 16 1 10 9 15 4 13 1 10 9 13 1 10 9 2
55 10 11 1 11 11 13 10 9 0 2 13 1 12 1 10 11 2 8 1 8 8 2 1 10 11 1 11 11 11 2 11 11 11 2 16 13 9 1 10 9 16 13 1 11 7 11 2 7 1 11 7 11 2 11 2
24 11 13 10 9 1 11 16 15 13 1 10 9 1 11 2 1 10 0 9 1 10 9 0 2
17 10 9 13 3 0 2 13 1 13 0 9 2 7 4 13 0 2
41 10 9 13 1 9 0 2 7 1 10 9 1 9 0 1 9 0 2 13 10 9 1 13 9 2 10 9 12 1 11 2 1 12 9 5 5 2 12 8 2 2
28 10 9 13 10 9 0 1 9 1 9 2 0 1 10 9 7 16 9 1 10 9 1 10 9 0 1 9 2
30 10 9 0 13 10 9 0 7 15 13 1 13 1 10 0 9 0 7 10 0 9 1 9 0 16 13 1 0 9 2
66 13 11 11 11 8 2 8 9 1 10 9 1 9 2 9 2 9 2 9 7 9 1 10 9 1 9 1 10 9 0 1 11 2 2 11 11 11 13 10 0 9 0 16 13 1 10 0 9 10 9 0 2 16 15 13 3 1 13 1 10 0 9 1 10 9 2
21 10 9 15 13 1 10 9 1 10 8 2 1 10 9 1 9 0 7 9 0 2
56 10 9 1 10 11 1 10 9 2 11 11 11 11 2 7 10 9 0 1 10 9 2 11 11 11 2 15 13 1 10 9 1 11 11 2 16 13 15 16 10 9 4 13 1 10 9 1 11 2 11 2 13 1 9 0 2
49 1 12 10 8 8 13 10 9 1 9 0 1 3 13 10 0 9 1 11 16 13 10 9 1 10 9 1 12 2 1 12 15 4 13 10 0 9 0 1 3 3 15 13 10 9 1 11 2 2
8 10 9 13 10 9 8 0 2
22 1 9 2 1 10 9 12 2 13 1 10 0 9 1 10 15 3 3 15 4 13 2
18 10 9 0 1 10 11 1 10 11 13 3 0 9 1 10 9 0 2
48 15 13 9 0 1 10 9 0 9 2 3 1 9 1 9 0 7 1 9 3 0 2 1 9 2 10 9 0 3 13 2 10 9 0 0 7 10 9 1 10 9 13 1 10 9 0 2 2
28 1 10 9 1 9 1 11 2 10 9 1 11 11 2 15 13 10 0 9 1 9 1 10 9 0 1 12 2
19 3 1 15 16 4 7 13 10 9 1 10 9 15 13 10 9 1 8 2
22 10 9 13 10 0 9 2 13 9 7 9 1 10 9 1 9 1 13 15 1 9 2
61 11 11 11 2 12 1 11 1 12 2 13 10 0 9 0 7 9 2 0 9 1 11 11 11 2 11 2 16 13 10 9 1 10 9 11 2 11 11 11 2 2 1 3 3 13 1 10 9 1 9 1 9 2 1 3 13 10 9 1 11 2
26 1 9 1 10 9 1 10 9 0 2 10 9 4 1 13 9 0 1 10 9 1 10 9 1 12 2
26 13 10 9 13 1 10 9 0 0 16 2 13 1 10 0 9 2 13 10 0 2 0 7 0 9 2
26 10 9 13 1 3 1 10 9 1 10 9 2 7 15 13 16 13 1 12 9 7 15 7 1 12 2
36 3 3 2 1 10 9 1 9 2 7 1 9 10 9 1 9 2 13 0 7 10 9 1 10 9 2 13 3 10 12 5 1 10 11 0 2
14 3 10 9 12 13 11 11 7 10 9 12 11 11 2
17 13 1 10 9 1 10 9 1 12 2 1 10 9 1 12 9 2
16 11 13 10 12 1 11 1 12 1 10 9 1 10 9 11 2
22 10 9 13 10 9 1 11 2 11 11 2 2 2 11 2 7 2 11 11 12 2 2
31 2 11 2 2 10 11 1 10 11 2 2 13 1 10 9 1 9 2 13 10 9 1 9 7 9 0 1 10 0 9 2
4 15 13 11 2
23 1 15 13 0 9 10 0 9 1 10 9 11 11 1 10 11 1 11 1 11 1 12 2
64 10 9 16 13 1 13 10 9 1 10 9 11 13 16 10 9 1 9 1 10 9 12 1 10 9 1 12 1 12 9 13 1 12 9 2 7 15 1 10 9 13 12 9 2 1 9 16 10 11 11 1 11 2 11 2 4 13 1 10 11 1 10 11 2
15 10 11 13 10 0 9 1 11 11 11 3 1 10 9 2
47 11 4 13 1 11 1 12 1 10 9 0 1 11 2 3 13 0 12 9 7 15 4 13 10 9 0 7 10 9 1 10 9 0 2 3 1 4 13 1 10 9 0 16 13 9 0 2
12 16 13 13 9 2 9 0 16 13 3 0 2
31 1 7 10 9 3 15 13 2 10 9 13 10 9 1 10 9 1 11 3 1 10 9 1 10 9 2 10 13 11 11 2
26 1 10 9 2 1 10 0 9 2 12 2 11 13 3 10 9 9 12 2 10 10 8 1 10 9 2
14 10 9 0 1 9 1 11 4 3 13 1 9 0 2
59 3 2 1 9 15 15 13 15 1 15 2 11 2 11 7 11 15 13 10 9 1 10 9 1 10 9 3 1 4 13 1 10 9 3 0 2 1 10 9 1 9 1 10 9 1 10 9 7 1 9 10 9 1 10 9 7 10 9 2
42 11 13 10 9 1 9 2 1 10 15 10 9 13 3 1 11 11 2 10 9 1 9 16 4 2 1 9 2 13 10 9 1 9 0 2 9 7 10 9 1 9 2
33 1 10 9 2 13 1 12 7 1 12 10 9 1 9 2 1 9 1 10 9 1 10 9 7 1 10 9 1 10 0 11 11 2
33 10 0 9 2 1 9 3 0 7 9 3 0 2 13 0 2 1 10 9 0 2 1 10 0 9 1 10 9 12 2 1 12 2
7 15 4 13 10 9 0 2
6 15 13 11 7 11 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
23 10 9 15 13 10 12 1 11 1 12 1 10 9 1 10 11 11 7 10 11 1 11 2
21 1 10 9 15 4 13 1 11 11 2 7 1 10 9 12 1 11 11 2 11 2
43 10 9 1 11 2 13 1 16 10 9 7 9 0 7 9 1 11 11 2 11 11 2 13 10 9 1 9 13 2 12 1 11 1 12 2 2 9 1 10 0 9 2 2
43 10 11 1 10 9 13 1 9 0 2 15 1 10 9 1 10 9 0 7 1 10 9 1 10 9 2 13 3 10 9 0 1 10 0 9 1 10 9 0 1 11 11 2
61 1 10 9 12 10 9 0 13 10 9 0 1 10 9 1 9 0 1 9 0 1 10 0 9 1 10 9 2 10 9 16 15 13 1 9 2 13 15 1 10 9 0 7 0 1 12 9 2 1 9 0 1 9 7 1 9 1 0 9 0 2
31 11 11 11 11 2 1 9 2 2 11 10 11 2 2 13 10 9 0 1 10 9 0 11 13 1 10 9 11 1 12 2
18 1 9 1 10 9 1 9 11 2 15 13 1 11 7 13 10 9 2
50 10 9 8 3 4 4 13 1 9 0 1 9 1 11 11 3 16 15 13 10 0 9 1 9 1 9 1 10 9 0 1 10 9 0 9 7 9 1 10 9 0 1 10 9 2 13 1 10 9 2
142 10 9 1 9 1 9 7 10 9 1 10 9 16 10 11 11 1 11 13 1 10 12 0 9 1 10 9 0 1 11 11 1 11 1 10 11 13 1 9 1 10 9 1 10 9 16 13 1 3 7 1 10 0 11 1 10 0 9 1 10 9 1 9 7 13 16 16 10 9 3 13 10 9 2 10 9 13 0 3 7 1 10 0 9 1 9 1 9 13 3 10 9 15 13 1 13 1 10 9 16 13 1 10 9 2 2 13 10 9 7 9 1 10 9 1 9 1 10 9 2 11 11 2 15 13 16 2 1 12 7 12 9 1 9 2 10 9 13 10 9 2 2
20 10 9 13 11 11 7 11 11 2 13 1 0 9 1 9 7 1 9 0 2
18 10 10 9 15 13 1 10 11 7 10 9 3 13 10 0 9 0 2
17 10 9 13 16 10 9 1 10 9 13 0 1 0 9 1 9 2
23 3 1 9 1 9 2 9 1 9 0 2 9 2 1 9 0 1 10 9 9 1 11 2
16 13 2 13 2 13 3 13 7 13 2 7 3 13 1 9 2
33 2 15 15 13 13 1 11 3 7 1 10 11 7 13 11 7 11 11 11 11 11 16 15 13 10 9 1 13 1 10 11 2 2
20 13 10 9 1 3 1 11 2 3 16 3 13 7 15 13 10 9 1 11 2
19 4 7 13 10 9 1 10 9 1 10 12 12 5 7 3 1 10 9 2
19 1 10 9 10 9 0 7 10 9 13 9 0 1 10 9 1 10 9 2
61 10 9 11 3 15 13 3 1 10 9 13 1 10 9 1 11 11 9 1 10 9 1 10 9 0 1 10 9 1 10 9 2 15 1 10 0 9 13 2 2 13 9 1 15 16 13 2 16 16 3 2 4 1 13 1 9 16 13 15 2 2
32 1 13 1 3 10 10 9 0 1 11 2 1 10 9 15 13 9 0 2 1 9 2 2 15 13 10 9 1 10 9 0 2
27 13 9 0 1 10 11 1 10 11 1 12 1 12 2 7 9 1 10 11 11 1 11 1 12 7 12 2
17 1 3 2 10 9 0 4 13 10 9 1 0 9 1 0 9 2
24 1 10 9 2 10 9 13 9 3 1 9 0 7 4 13 10 9 1 10 9 1 10 9 2
23 10 9 1 10 9 15 13 1 10 9 1 3 4 13 1 10 9 1 9 1 10 9 2
34 10 9 11 1 11 13 10 9 0 0 0 7 15 0 2 1 12 9 1 0 2 12 9 1 9 7 1 12 1 12 9 1 9 2
10 4 13 3 10 12 1 11 1 12 2
32 13 10 9 0 2 9 1 10 11 11 1 11 1 12 9 2 8 2 8 2 2 13 2 10 0 9 1 10 9 0 2 2
12 1 10 15 13 10 9 1 9 7 0 9 2
65 11 13 1 10 9 10 9 0 1 10 11 2 9 15 13 1 10 9 0 1 9 1 10 9 0 2 13 1 10 9 1 16 13 1 10 9 1 9 0 2 7 1 10 9 1 11 2 13 7 13 10 9 1 9 15 13 10 9 1 10 9 1 10 9 2
28 10 9 13 0 7 15 13 13 1 10 9 1 10 9 1 9 1 9 0 7 9 0 1 9 1 10 9 2
18 10 9 1 10 9 7 3 10 9 3 0 2 4 13 1 10 9 2
7 10 9 3 0 4 13 2
14 13 1 10 9 2 2 11 1 10 11 1 11 2 2
20 1 10 9 1 12 2 4 1 13 10 9 0 1 10 9 1 10 11 0 2
43 10 9 13 10 9 1 10 9 16 13 1 10 9 1 10 9 0 2 13 1 9 0 2 9 9 2 9 1 9 7 10 9 16 13 10 9 1 10 9 0 1 15 2
18 13 10 9 1 10 9 1 10 9 15 4 13 3 1 11 11 11 2
19 16 10 9 13 3 13 10 0 2 1 10 3 2 3 13 10 9 0 2
23 10 0 9 13 10 9 1 13 10 9 1 9 1 15 1 10 9 0 1 11 2 11 2
24 16 10 12 9 13 10 9 0 1 10 9 2 10 12 1 11 1 12 11 13 1 10 9 2
27 3 15 4 13 10 9 1 10 9 2 16 4 13 1 9 7 13 3 0 1 15 16 13 1 10 9 2
83 10 9 13 10 11 9 0 2 13 1 10 9 1 12 2 13 1 12 1 10 9 0 0 16 15 13 1 12 2 1 10 9 1 9 0 0 2 0 2 1 10 9 0 0 2 8 8 2 2 13 1 12 2 1 12 1 10 9 11 0 7 0 2 7 1 12 1 10 9 0 0 2 1 3 13 0 9 0 1 9 3 0 2
32 3 13 9 3 4 1 13 10 9 1 10 9 0 7 4 13 1 12 1 10 9 1 11 11 2 1 10 15 13 12 9 2
30 3 1 13 1 10 9 2 11 4 1 13 1 10 9 7 0 9 1 10 9 9 2 9 0 1 10 9 1 11 2
15 10 9 4 13 7 13 1 1 10 9 10 9 1 9 2
79 9 1 10 9 0 2 9 1 10 11 1 11 2 12 2 2 9 1 10 9 1 10 9 1 9 2 12 2 2 9 0 1 10 11 1 11 2 12 2 7 10 9 1 10 9 1 12 2 3 1 12 2 9 1 9 1 12 9 1 9 2 1 12 9 1 9 2 13 1 10 11 11 11 7 11 1 11 2 2
21 1 10 9 2 7 13 1 10 9 2 4 13 10 9 2 13 1 7 10 9 2
30 10 9 13 1 10 9 1 10 9 7 1 9 1 15 10 9 0 13 13 10 9 0 2 7 10 9 3 13 0 2
47 10 10 11 1 10 11 0 13 1 12 7 12 11 2 12 7 12 11 2 2 3 2 7 1 12 7 12 11 2 2 12 7 12 11 2 2 13 1 10 9 10 9 1 10 9 0 2
24 15 15 13 9 0 7 9 1 10 9 2 15 2 10 9 9 2 0 3 2 0 7 9 2
30 1 0 9 13 3 1 10 9 11 11 2 10 9 16 13 1 12 9 2 9 7 10 10 9 16 13 10 9 0 2
9 2 3 13 9 1 10 0 9 2
37 1 10 9 0 1 2 11 2 2 11 13 10 0 9 0 1 10 9 2 1 10 15 13 10 9 1 10 2 11 11 11 11 2 1 12 2 2
7 13 10 9 1 9 0 2
44 1 10 0 9 1 10 9 12 15 13 10 9 1 10 11 16 13 0 9 1 10 9 2 10 9 15 13 9 1 10 9 2 10 9 2 9 1 9 2 9 0 7 9 2
16 10 11 13 1 15 2 1 15 1 10 9 16 13 1 9 2
29 10 9 13 15 1 10 9 1 10 11 1 11 2 12 2 2 16 13 9 1 10 9 1 9 0 1 10 11 2
20 1 10 0 9 13 10 9 0 7 1 10 9 10 9 0 12 1 11 11 2
17 15 13 10 9 1 10 0 9 1 10 11 1 10 11 11 11 2
13 15 13 9 1 9 7 9 1 9 1 10 9 2
71 15 2 16 13 2 1 15 2 2 10 11 2 7 2 10 11 2 2 13 10 0 9 0 0 16 10 9 1 10 9 0 2 9 1 12 2 12 7 12 2 12 7 9 0 1 2 9 0 2 2 13 13 2 9 1 12 7 3 9 0 2 13 1 9 1 12 7 3 9 2 2
35 3 1 13 15 1 10 9 1 10 9 1 9 0 2 10 9 7 0 11 2 11 11 2 13 0 9 1 11 1 13 15 1 10 9 2
19 10 9 3 4 13 1 10 9 13 3 10 9 1 9 3 0 1 11 2
30 1 10 0 9 2 1 9 1 10 9 11 2 15 13 10 9 3 0 1 9 0 2 9 0 0 7 9 1 9 2
13 10 9 11 13 10 0 9 0 1 10 9 11 2
18 10 11 11 13 10 9 0 13 1 10 11 11 1 10 11 11 11 2
6 13 1 9 11 12 2
65 1 10 9 1 12 15 13 1 10 0 9 1 10 9 0 16 13 10 9 1 10 0 9 1 10 9 9 1 11 2 13 10 9 1 10 13 15 10 9 1 11 1 12 2 7 13 15 11 1 10 0 9 2 12 2 2 1 9 1 10 9 11 11 11 2
11 3 15 13 1 10 9 16 13 9 0 2
17 13 0 1 10 9 1 9 1 11 1 12 9 7 13 12 9 2
17 10 9 0 2 1 10 9 1 11 2 13 9 3 0 1 9 2
45 1 12 9 1 13 10 9 2 1 10 11 11 1 11 1 9 1 9 1 12 5 8 2 13 1 11 1 13 1 10 11 11 2 7 10 9 0 13 10 9 1 10 9 0 2
24 10 9 0 7 9 1 10 9 1 10 9 13 11 11 11 2 7 3 13 10 9 1 15 2
35 10 12 1 11 2 10 12 9 1 9 0 2 12 9 2 13 1 11 11 2 4 13 10 9 0 2 3 16 15 4 4 13 1 11 2
27 11 11 11 2 11 2 11 1 12 2 8 2 12 1 11 1 12 2 13 10 9 2 9 7 9 0 2
21 10 8 16 4 13 13 3 10 9 8 5 8 5 8 13 15 10 8 1 9 2
40 1 10 0 9 7 3 1 12 2 2 11 2 13 10 9 0 0 1 11 11 2 1 10 15 13 2 11 1 11 2 2 16 4 1 13 1 10 9 0 2
26 10 9 15 13 1 10 12 9 2 16 10 9 1 9 1 10 9 12 13 10 9 13 1 10 9 2
42 13 9 1 10 11 11 3 13 1 10 9 11 2 16 15 13 3 1 9 0 9 16 13 16 10 9 1 10 9 1 10 11 11 7 10 11 11 3 13 3 0 2
22 10 9 1 10 9 1 10 0 9 13 10 9 1 12 9 13 2 7 10 9 13 2
40 3 1 9 2 7 1 15 1 10 9 1 10 9 2 4 13 10 12 9 16 13 1 9 1 10 9 16 13 16 10 9 4 13 1 10 9 7 10 9 2
20 10 9 2 9 13 10 9 0 0 1 10 9 0 7 9 1 10 11 11 2
35 1 9 2 10 9 13 16 13 0 13 10 9 1 10 9 7 3 1 9 10 9 15 13 1 9 16 15 4 13 1 15 1 10 9 2
47 1 12 2 3 13 9 7 9 1 10 11 1 10 11 11 1 10 11 2 15 4 4 13 1 9 1 10 9 12 1 10 9 1 13 7 13 10 9 1 10 9 1 10 11 1 11 2
25 1 9 10 9 1 11 2 11 2 7 1 11 2 1 11 2 3 13 0 13 3 10 9 0 2
12 10 12 9 4 13 1 10 9 0 1 12 2
32 3 2 11 0 16 10 9 2 2 1 9 7 1 9 2 2 16 13 13 10 9 13 1 10 2 9 1 10 9 0 2 2
75 13 1 11 1 10 11 2 0 9 0 1 11 1 10 15 13 10 9 2 13 9 1 11 11 1 12 7 12 2 7 10 9 1 10 11 13 9 1 11 2 1 3 15 13 1 12 2 1 10 9 1 10 1 10 11 2 1 15 13 1 12 1 10 9 1 10 9 1 11 11 1 10 11 11 2
45 1 13 1 12 10 9 15 13 1 12 2 11 15 13 1 10 9 1 11 11 2 1 10 9 1 10 11 11 1 11 11 7 11 16 13 1 10 9 1 10 11 11 1 11 2
22 13 15 10 9 1 13 15 2 13 3 9 1 10 9 1 10 9 7 10 9 0 2
37 10 9 2 11 2 13 10 9 1 11 11 11 2 16 13 1 10 11 11 1 15 15 13 3 11 7 10 11 11 2 1 10 11 7 10 11 2
15 1 3 10 0 9 15 13 1 10 9 1 10 0 9 2
27 1 11 3 13 10 0 9 16 13 1 11 2 11 13 10 9 7 13 1 10 9 0 10 9 1 9 2
31 10 8 8 4 13 1 12 9 16 13 1 10 9 11 3 1 10 12 1 11 1 12 2 3 15 13 10 9 1 9 2
35 3 4 13 16 16 3 4 13 11 10 9 2 10 9 1 16 10 9 13 10 9 1 10 9 15 13 15 0 7 16 13 0 1 15 2
25 10 9 1 10 9 13 10 1 13 15 1 10 10 9 3 16 15 4 13 10 9 1 10 9 2
20 1 10 9 2 1 10 9 3 4 13 3 2 1 15 15 4 13 10 9 2
46 10 9 7 10 9 0 3 13 10 0 9 1 10 9 7 9 0 13 1 10 11 7 10 11 1 10 10 9 1 10 9 1 10 9 1 9 1 10 9 2 10 9 7 1 9 2
25 15 13 10 12 9 2 12 9 7 12 9 1 12 2 7 3 1 12 13 12 8 7 9 12 2
17 13 10 0 9 2 10 0 9 16 13 1 10 9 0 10 9 2
15 1 9 1 10 9 15 13 1 10 9 10 9 11 11 2
35 1 9 1 10 9 7 9 0 0 2 10 9 0 13 3 1 15 1 10 9 2 13 10 9 2 1 9 2 1 10 12 9 1 9 2
16 10 0 9 13 10 9 1 11 11 7 11 11 1 10 9 2
15 4 7 13 3 16 4 13 3 16 3 13 0 13 9 2
30 15 4 13 10 9 1 10 9 1 10 9 0 2 3 3 1 10 9 0 7 3 1 10 9 0 2 0 15 13 2
22 10 9 13 10 9 1 10 15 4 13 15 9 1 13 10 9 0 1 10 9 9 2
37 11 2 3 13 1 11 1 11 2 13 10 0 9 1 9 1 10 11 1 13 15 16 10 9 15 16 13 13 13 7 1 10 11 3 13 9 2
62 1 10 12 9 2 10 9 1 9 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
17 15 13 12 9 1 10 11 11 12 7 12 1 10 11 11 12 2
9 15 3 13 9 7 9 1 9 2
25 10 9 13 1 9 1 10 9 0 16 15 13 7 16 13 0 9 1 13 9 1 10 9 0 2
53 3 3 2 10 11 15 4 13 1 11 11 2 11 2 11 2 1 13 3 1 11 2 3 11 11 2 1 10 12 9 2 15 13 1 11 11 2 10 12 1 11 1 12 2 16 11 13 1 12 9 1 9 2
42 1 15 2 10 9 13 10 9 0 7 0 7 2 1 15 2 13 10 9 13 3 1 9 1 0 9 16 3 13 10 9 1 0 9 1 11 11 11 7 11 11 2
62 1 10 12 9 2 10 9 1 11 13 0 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
13 1 10 0 9 13 12 9 16 13 3 1 11 2
34 11 13 16 3 7 13 10 9 13 1 9 16 13 9 2 7 1 15 13 15 1 10 9 16 4 13 1 10 9 9 1 10 9 2
14 3 15 2 1 11 11 2 15 4 13 10 9 0 2
12 10 9 1 9 13 1 12 8 5 5 5 2
32 10 9 13 9 8 1 10 11 8 11 7 11 8 11 11 2 1 3 12 9 1 10 9 11 11 2 10 9 1 9 2 2
37 1 13 15 2 15 13 1 11 11 16 13 1 10 11 2 16 15 13 3 1 13 15 1 13 9 1 10 11 2 11 2 11 2 11 11 11 2
38 10 9 0 13 10 9 1 9 0 16 13 10 9 1 10 9 1 9 3 0 7 0 16 15 13 0 9 1 10 9 0 13 1 9 7 9 9 2
22 10 9 0 0 15 13 1 13 9 0 2 13 10 9 0 1 10 9 1 10 9 2
34 13 10 9 0 0 3 0 2 10 9 0 13 1 12 5 8 2 0 9 0 2 0 1 10 12 5 2 7 0 9 1 9 0 2
61 1 9 1 10 9 2 11 3 4 13 16 3 1 10 9 3 15 4 13 2 1 9 1 10 9 2 2 10 9 1 9 1 10 9 1 9 0 2 2 1 10 9 3 3 1 13 10 9 1 10 9 7 10 9 1 2 10 9 0 2 2
46 10 9 13 11 11 11 2 0 1 11 2 11 2 7 0 1 11 16 15 13 1 11 1 9 1 10 9 12 1 9 0 1 9 1 10 9 0 3 1 13 12 9 1 0 9 2
35 13 10 9 0 3 1 10 9 1 10 11 11 2 7 13 0 1 10 11 11 11 3 7 1 10 15 13 3 10 9 2 9 7 9 2
21 16 13 10 0 9 0 2 13 3 1 10 11 11 7 1 10 9 13 1 11 2
6 13 1 11 1 11 2
23 11 15 13 1 13 10 9 1 10 9 2 10 9 13 1 3 1 12 9 1 10 11 2
35 10 9 13 12 8 1 0 1 10 9 1 9 1 9 1 12 5 1 0 7 4 13 3 1 16 10 9 15 13 1 10 9 1 11 2
31 10 9 1 11 11 7 13 15 1 9 15 13 1 10 9 1 10 9 0 2 1 10 15 13 3 1 10 9 11 11 2
13 1 11 11 2 10 9 3 4 13 16 13 13 2
51 4 13 2 1 15 2 10 9 0 1 11 11 2 12 2 2 1 9 11 11 2 12 2 2 1 9 1 11 11 11 2 12 2 2 1 9 11 11 2 12 2 7 1 9 11 11 11 2 12 2 2
24 1 10 12 8 15 13 9 0 1 9 1 11 1 10 9 1 0 9 1 11 7 11 11 2
25 11 11 13 1 10 9 0 2 9 1 10 9 2 16 13 10 0 9 1 10 9 1 9 0 2
33 1 9 1 10 9 1 12 2 11 7 10 9 13 16 10 9 1 11 1 10 0 9 4 13 15 1 3 2 13 15 13 3 2
38 10 9 1 11 11 15 13 1 10 12 9 1 10 0 9 1 10 9 7 13 12 0 9 13 1 9 1 9 7 1 10 0 9 1 10 9 11 2
39 10 9 2 16 13 10 9 0 1 10 9 11 7 11 11 11 7 10 9 11 7 11 2 4 13 1 10 0 11 1 12 7 13 13 15 3 1 12 2
16 10 9 0 13 10 9 1 11 11 1 11 13 1 9 0 2
34 15 11 13 10 9 7 9 0 2 13 1 10 9 1 9 1 10 11 2 9 1 11 11 2 1 10 9 1 11 7 9 1 11 2
24 1 12 2 10 11 15 13 10 9 11 11 11 11 2 1 9 2 11 11 1 11 11 2 2
40 1 10 9 12 2 1 10 9 1 11 1 10 11 2 13 10 0 9 1 13 10 11 1 11 11 7 11 11 1 10 11 1 11 7 11 11 1 10 11 2
34 1 9 0 2 10 9 15 13 1 10 9 1 10 15 13 10 9 0 1 10 9 7 9 7 1 10 15 10 9 13 10 9 0 2
12 13 9 1 9 1 12 9 1 10 9 0 2
23 10 9 0 1 10 9 1 9 13 1 10 11 1 11 2 1 12 2 13 13 10 11 2
28 1 10 9 13 9 16 15 4 13 1 13 9 2 13 1 9 0 7 4 13 2 1 9 2 9 11 11 2
18 10 9 13 1 12 9 1 10 9 10 11 7 13 1 10 9 3 2
23 10 11 2 9 13 0 1 9 7 13 10 9 0 2 16 13 10 9 1 10 9 0 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
28 4 13 3 9 1 10 9 1 9 15 13 1 12 9 1 10 9 1 12 9 2 10 0 9 1 10 9 2
31 10 9 13 10 9 16 13 10 9 0 7 9 0 1 4 13 1 0 2 7 1 15 3 13 1 10 9 1 9 2 2
12 1 12 13 3 10 9 1 10 11 11 11 2
22 16 10 9 0 4 13 10 9 1 3 9 2 3 15 13 10 9 1 10 9 0 2
11 10 9 1 9 13 1 11 1 10 9 2
42 4 13 10 9 1 11 11 7 10 9 1 9 1 10 9 3 3 15 4 13 12 9 2 15 15 4 13 1 12 9 7 4 13 10 12 9 1 13 15 10 9 2
38 10 9 13 9 1 13 10 9 1 10 9 7 1 10 9 1 10 9 1 13 10 9 2 7 4 13 1 10 9 0 1 10 9 1 10 9 0 2
54 10 9 0 13 10 9 1 11 1 10 12 0 9 1 10 9 2 1 9 1 10 11 2 3 2 4 13 10 10 9 0 16 15 4 13 1 12 1 9 1 10 1 12 1 10 15 3 15 13 7 15 13 11 2
20 1 9 10 0 9 16 4 13 11 13 1 10 9 1 9 2 1 11 11 2
41 11 11 7 11 2 11 2 11 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 13 10 9 0 1 9 0 2 1 9 1 10 9 7 10 9 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
22 10 9 4 13 1 10 9 1 10 9 2 1 15 15 10 9 4 13 1 9 0 2
19 10 9 1 10 9 0 2 12 9 13 13 1 10 9 1 9 1 11 2
10 15 13 9 0 1 10 9 1 11 2
14 1 10 9 1 13 1 10 9 15 13 7 13 0 2
6 7 10 8 13 0 2
32 11 13 15 1 15 16 4 13 2 3 7 4 13 16 13 16 13 11 11 2 7 10 9 11 3 13 16 10 9 15 13 2
38 1 9 2 16 13 1 10 9 1 10 9 11 1 10 11 10 11 1 11 13 16 13 10 0 9 7 11 11 2 10 9 16 3 15 4 13 0 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
17 4 13 1 11 1 10 9 1 10 9 10 12 1 11 1 12 2
25 10 9 0 13 10 0 9 16 13 10 9 1 0 9 15 4 4 3 3 13 1 10 9 0 2
30 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 1 10 11 2
12 11 4 13 1 10 9 1 10 12 9 0 2
27 9 1 10 11 11 11 11 11 7 9 1 11 11 11 7 11 11 11 2 9 0 1 10 9 12 5 2
28 15 4 13 9 1 10 9 0 3 1 10 9 1 10 9 1 10 9 11 7 1 10 9 0 1 10 11 2
10 1 10 9 13 10 9 1 9 0 2
20 15 13 1 10 9 1 9 1 10 9 2 8 2 7 10 9 2 8 2 2
14 3 15 13 1 10 9 1 11 7 15 13 10 9 2
19 10 9 13 10 9 1 9 13 13 15 1 10 9 2 1 9 3 0 2
10 10 9 1 11 2 15 13 1 11 2
28 13 10 9 1 13 10 9 1 10 9 0 2 0 2 7 10 9 0 2 2 9 2 9 2 9 2 9 2
71 1 10 9 2 13 13 16 1 0 9 1 10 9 0 1 10 9 1 11 11 2 15 13 1 10 9 1 12 9 3 2 9 2 9 16 13 3 3 2 16 1 11 1 11 3 13 10 3 2 9 2 7 16 1 10 9 10 9 4 13 2 12 1 11 7 12 1 11 11 2 2
22 1 10 9 1 10 0 9 15 13 12 9 1 9 13 1 9 0 2 16 13 9 2
31 10 9 13 0 2 10 9 13 10 0 9 0 0 7 10 9 2 10 9 2 1 15 9 16 4 13 3 1 10 11 2
9 11 11 15 13 13 1 10 9 2
24 1 11 1 12 2 13 11 2 10 9 11 16 13 10 9 1 9 13 1 11 1 9 11 2
20 1 10 11 1 9 2 9 1 10 11 11 2 15 13 10 9 1 10 9 2
37 11 11 13 1 10 9 1 9 2 7 15 13 3 1 12 1 10 13 10 11 1 10 9 1 11 2 16 4 13 1 10 11 7 1 10 11 2
14 1 13 11 2 13 3 7 0 16 4 1 13 0 2
6 11 11 2 9 2 2
20 3 2 10 9 13 10 9 0 1 10 15 15 13 13 10 9 1 9 0 2
30 11 13 0 9 1 9 16 13 1 10 9 7 10 9 2 16 15 13 3 3 1 10 9 1 11 11 11 1 12 2
12 1 10 9 1 10 9 13 10 9 1 11 2
20 10 0 9 13 2 10 9 0 2 10 9 3 9 7 10 9 1 11 2 2
36 1 0 16 3 13 13 15 10 9 1 9 1 10 9 2 13 16 11 13 10 9 3 13 9 1 0 9 7 1 3 15 8 13 10 9 2
8 13 10 9 0 2 1 9 2
17 15 2 1 10 9 2 13 1 10 9 1 10 15 13 10 9 2
14 11 2 13 10 9 1 9 0 0 1 10 9 11 2
17 10 12 1 11 1 12 10 11 7 11 13 10 9 9 1 11 2
51 10 9 15 13 1 10 9 1 10 9 1 10 9 1 10 9 1 11 2 10 9 1 10 9 7 10 9 1 9 1 10 9 1 13 10 9 1 9 16 13 3 10 9 1 10 9 7 1 10 9 2
30 1 10 9 15 13 10 11 11 12 2 10 11 11 2 10 11 11 2 10 11 11 2 10 11 11 7 10 11 12 2
21 4 13 10 9 0 7 15 4 13 10 10 9 1 13 10 9 1 10 9 9 2
22 1 9 2 1 10 9 13 9 1 13 1 13 10 9 2 8 16 13 10 9 0 2
50 13 13 10 9 0 2 11 7 11 11 2 11 11 2 11 11 7 11 11 2 1 15 2 13 10 9 1 12 1 10 12 9 0 1 10 11 2 7 13 1 16 11 4 13 9 0 1 3 0 2
20 1 10 9 2 9 7 9 13 10 9 16 13 16 10 9 13 0 1 9 2
22 10 9 4 13 1 9 2 7 10 9 9 4 13 1 13 9 1 3 1 12 9 2
26 10 9 1 12 9 4 13 1 10 9 1 10 9 1 10 9 0 1 11 11 2 1 10 0 9 2
28 10 9 1 9 7 9 13 4 13 3 1 10 9 0 2 16 3 10 9 13 13 3 1 10 9 1 15 2
27 11 13 15 1 10 9 16 13 1 15 8 15 2 1 10 16 13 10 9 3 0 7 1 15 13 9 2
12 3 15 13 0 9 7 1 9 7 1 9 2
53 13 1 10 9 1 10 11 7 13 1 10 9 0 1 11 11 1 11 7 11 11 1 11 1 10 9 2 11 1 11 7 11 1 10 15 2 11 1 10 9 7 10 11 1 10 9 7 9 2 15 1 11 2
15 10 9 4 3 13 2 11 2 8 8 8 8 2 2 2
38 10 9 15 4 13 1 9 0 1 10 9 1 11 11 1 11 11 2 8 11 11 1 10 11 7 10 9 11 11 2 9 1 10 11 11 1 11 2
9 9 0 2 3 0 9 7 9 2
68 1 10 9 12 11 13 10 9 1 13 1 11 11 11 1 9 1 10 11 11 1 10 9 1 10 11 11 2 16 15 13 1 12 1 10 11 11 11 11 11 2 11 2 2 10 9 1 10 11 11 1 11 2 11 2 2 1 10 15 3 1 10 9 11 11 13 9 2
13 1 10 9 1 10 9 7 2 3 2 13 9 2
22 10 9 0 1 9 13 1 12 9 2 1 10 15 10 9 13 1 9 12 1 12 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
31 3 13 9 0 0 2 3 13 9 0 2 3 13 9 0 0 2 4 4 13 1 9 0 7 3 13 9 1 10 9 2
19 16 13 11 2 15 4 13 15 1 10 0 9 16 13 3 7 1 9 2
19 13 0 13 16 15 13 10 0 9 1 10 9 1 10 9 11 11 11 2
40 10 8 11 13 10 9 1 9 1 10 11 11 1 12 2 10 9 1 9 1 10 11 1 11 1 12 2 13 10 9 1 9 1 10 11 1 11 1 12 2
12 13 10 9 1 13 10 9 0 1 11 11 2
13 3 10 9 4 13 1 10 9 1 10 9 0 2
30 11 11 13 10 9 1 9 1 9 0 13 1 11 12 10 12 1 11 1 12 1 10 15 13 3 10 11 11 12 2
39 1 10 9 12 10 9 15 13 3 1 9 0 2 1 10 9 0 2 10 9 13 1 9 0 7 10 9 2 13 1 10 0 9 0 7 1 10 9 2
12 10 9 1 10 10 9 13 10 9 1 9 2
15 3 2 3 15 13 10 9 1 10 9 1 11 7 11 2
49 1 10 9 13 9 1 12 9 16 13 9 0 1 10 9 0 7 3 10 9 1 9 1 9 0 13 1 10 2 11 11 1 11 1 11 11 2 2 16 4 1 13 10 9 0 2 11 2 2
40 15 13 15 1 10 9 16 13 1 10 9 10 9 11 1 10 13 10 9 1 10 9 11 11 2 15 4 13 1 10 9 1 9 1 10 9 1 9 0 2
78 3 13 16 11 13 1 2 11 2 2 9 0 2 11 11 2 2 10 9 1 0 9 0 2 16 1 10 9 15 13 1 11 2 11 11 2 2 10 9 3 13 1 10 9 2 16 13 13 1 10 0 9 1 16 13 10 9 1 15 2 16 15 15 13 1 10 9 1 11 1 10 9 11 2 11 11 2 2
24 10 9 2 9 0 7 11 1 9 0 2 11 11 2 13 10 9 1 9 1 10 9 11 2
27 11 13 10 9 1 11 1 10 9 1 10 9 1 9 7 9 1 9 1 10 12 1 13 10 9 0 2
14 1 9 1 15 2 15 4 13 1 10 11 11 0 2
15 2 10 9 7 10 9 13 2 1 9 2 9 0 2 2
31 1 0 9 2 13 1 12 9 1 11 2 16 15 13 10 9 0 1 10 9 11 2 9 13 1 10 9 1 10 11 2
31 16 13 10 9 13 0 4 1 13 10 9 7 13 3 2 7 1 0 13 10 9 16 4 7 13 1 10 13 1 11 2
53 13 1 11 2 11 7 11 13 13 15 10 9 2 7 4 13 1 11 15 13 1 10 9 2 1 16 13 1 10 9 1 13 3 10 9 15 13 0 1 10 14 9 2 7 1 10 9 13 10 9 7 13 2
29 15 13 2 3 3 2 9 1 9 7 9 0 2 7 1 10 9 15 13 9 7 9 1 9 1 9 1 9 2
39 1 7 3 15 13 1 15 2 11 13 10 9 0 1 0 9 15 0 2 1 9 10 0 11 8 13 10 8 7 13 9 1 13 9 1 8 1 9 2
19 1 12 4 13 11 1 11 2 7 4 13 1 10 12 9 1 0 9 2
63 13 1 11 1 12 2 4 13 1 11 1 10 9 0 0 2 7 13 1 9 0 1 10 9 1 12 9 2 12 1 15 9 2 13 1 10 9 1 11 16 4 13 1 9 1 12 9 13 1 9 0 13 12 9 2 16 13 12 9 7 12 9 2
18 15 13 10 9 16 3 13 10 9 0 7 3 10 9 1 10 9 2
31 10 9 1 10 9 0 13 0 2 7 15 13 1 0 0 2 4 4 13 15 1 10 0 9 1 10 9 7 10 9 2
31 15 15 13 1 15 13 15 1 0 9 2 7 3 1 10 13 15 10 9 4 13 15 1 9 1 10 9 1 9 0 2
28 1 9 0 2 11 11 13 1 0 9 0 1 9 1 10 9 11 2 1 0 9 1 11 11 7 11 11 2
22 1 9 1 10 0 9 10 9 13 3 0 1 9 0 7 10 9 0 13 1 12 2
20 1 11 7 11 2 10 11 11 13 1 10 10 9 7 9 10 12 1 11 2
20 1 10 9 1 11 13 16 10 9 0 13 1 9 1 9 1 9 7 9 2
12 1 10 9 3 4 1 13 10 12 9 0 2
17 3 13 10 9 1 9 7 13 9 1 11 2 11 7 11 11 2
34 1 10 0 9 2 11 11 4 4 13 1 10 0 9 1 9 1 0 9 1 9 16 13 9 1 9 7 1 9 1 9 1 9 2
16 13 9 1 9 0 1 9 0 0 9 16 13 13 9 0 2
35 9 3 3 13 1 10 9 2 13 1 0 9 13 1 0 9 1 9 3 0 2 16 15 13 10 9 1 11 7 10 9 1 11 11 2
11 1 10 9 12 13 10 9 1 12 9 2
52 10 9 0 2 16 13 11 2 13 0 1 13 1 10 9 16 13 10 9 1 10 9 0 1 10 9 0 2 9 16 15 13 13 1 10 9 1 13 16 13 10 9 0 1 10 9 1 11 11 1 12 2
18 11 11 13 10 9 1 9 1 10 9 11 1 10 9 1 10 11 2
13 13 10 0 9 3 0 2 0 2 0 7 0 2
59 1 10 12 9 2 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
17 10 9 0 7 0 7 1 10 9 0 1 10 9 1 9 0 2
61 10 9 3 4 13 9 1 10 10 11 2 12 2 3 13 16 10 11 13 2 15 13 11 7 13 10 0 9 1 10 11 11 2 13 1 13 9 0 1 9 0 2 1 10 9 1 13 10 9 0 16 13 1 10 11 9 1 10 9 0 2
35 10 12 5 9 13 9 1 11 1 12 2 10 12 5 9 15 13 1 11 1 12 2 7 10 12 5 1 11 11 1 12 2 5 2 2
13 13 3 16 10 9 13 1 10 9 1 9 0 2
79 1 13 15 11 11 13 10 9 16 13 16 10 9 1 10 11 16 13 1 10 11 2 11 7 9 0 13 3 1 10 9 1 10 11 10 9 0 2 3 16 10 9 1 10 11 2 9 2 7 1 10 9 16 3 13 1 10 11 15 13 1 10 9 1 9 1 10 11 2 7 10 13 10 9 3 13 3 9 2
16 1 9 1 15 13 10 9 0 1 10 15 3 15 4 13 2
25 10 9 1 10 9 0 4 3 13 2 16 13 10 11 15 13 2 1 10 9 2 0 9 0 2
51 10 9 1 11 7 11 13 10 9 1 10 9 1 10 9 2 13 1 10 9 11 11 2 10 9 11 1 11 7 11 11 11 2 7 10 9 11 11 7 11 11 2 11 2 13 3 11 1 10 9 2
47 2 15 13 1 10 0 9 3 1 10 9 1 9 1 9 1 0 9 1 10 9 0 1 0 9 1 13 10 9 2 2 13 1 10 9 10 9 0 7 9 0 1 11 2 11 11 2
32 13 10 9 1 10 9 11 1 10 9 0 2 10 9 3 0 1 10 9 11 11 16 4 2 1 10 9 2 13 7 13 2
52 1 11 1 12 2 1 10 9 1 10 11 11 2 4 13 9 0 1 10 11 11 11 11 11 2 11 1 11 1 10 11 7 10 11 11 7 11 1 10 11 1 9 0 7 11 1 10 11 11 1 11 2
49 9 0 1 9 1 9 0 2 9 2 9 2 9 1 9 0 2 7 15 13 1 9 0 2 9 0 2 9 2 9 0 2 9 0 2 9 1 3 1 12 9 1 10 9 1 10 9 12 2
24 8 10 9 1 10 9 13 10 9 0 15 13 10 9 1 10 9 7 10 9 1 10 9 2
30 11 11 11 2 10 9 13 2 2 11 2 9 1 11 2 13 1 0 9 10 9 15 4 13 2 1 11 11 2 2
12 0 9 1 9 13 3 1 10 9 1 11 2
14 15 13 1 16 10 9 0 1 10 9 13 10 9 2
33 13 1 10 9 12 1 11 2 11 2 16 10 9 1 11 4 13 1 9 0 1 10 9 1 10 12 11 11 1 10 11 12 2
19 3 2 10 9 13 1 10 9 7 10 9 2 1 9 15 13 10 9 2
21 10 9 3 2 10 9 1 10 9 1 11 11 11 15 13 1 9 1 11 11 2
8 9 0 1 10 11 1 12 2
48 13 1 10 9 1 10 9 0 1 11 7 10 9 1 11 2 1 10 9 1 11 1 10 11 2 1 10 15 1 11 7 10 11 2 1 10 9 1 11 2 7 1 10 11 11 7 11 2
51 16 4 13 10 9 1 10 9 2 10 9 0 11 11 4 13 10 9 1 13 9 16 13 1 10 9 1 9 1 9 0 16 13 9 1 1 10 11 1 11 1 10 9 1 2 13 1 10 9 2 2
16 10 9 7 15 15 4 13 3 0 1 10 9 1 10 9 2
18 10 11 11 4 13 1 9 1 10 9 12 1 10 9 0 11 11 2
30 1 10 12 9 1 9 0 16 13 1 11 2 10 12 13 1 10 9 0 2 13 13 2 9 1 3 1 12 9 2
27 10 9 1 11 13 3 2 1 10 9 1 10 9 16 13 1 10 9 11 11 7 1 10 9 11 11 2
69 3 2 10 9 0 3 13 10 9 1 10 11 1 11 1 10 9 10 9 1 9 1 10 9 2 9 0 7 9 0 0 16 15 13 1 10 9 2 16 15 4 13 10 9 2 7 9 0 7 0 0 1 10 9 1 10 9 0 0 1 9 16 15 13 1 10 9 0 2
10 13 0 1 10 9 1 9 1 11 2
29 15 4 13 10 9 1 9 2 7 4 13 16 3 15 13 10 9 3 0 7 1 10 9 16 13 10 9 13 2
42 1 11 1 12 2 10 9 2 1 15 10 8 0 9 11 11 7 8 9 1 10 11 2 13 1 10 9 12 9 1 10 9 2 15 4 13 1 10 9 11 11 2
29 15 13 1 10 9 8 1 12 9 2 7 10 9 1 10 8 1 11 8 2 8 8 8 8 2 1 12 9 2
61 1 10 0 9 1 10 9 2 15 13 1 10 9 0 2 7 13 1 10 9 1 10 9 1 10 12 9 2 13 1 11 2 11 2 1 12 2 1 9 2 13 1 9 0 1 9 0 2 13 10 9 11 2 1 10 9 1 11 7 11 2
23 1 9 1 16 10 9 13 0 4 7 13 15 10 9 2 7 13 3 13 7 3 13 2
35 13 1 10 9 1 10 9 1 12 7 13 1 9 7 9 1 10 9 1 9 7 1 9 2 12 2 7 9 1 10 9 2 12 2 2
18 11 13 1 10 9 1 9 1 11 1 11 2 10 9 1 10 9 2
20 3 13 9 0 16 15 13 3 1 11 7 13 0 1 10 9 1 10 9 2
32 13 10 9 0 0 16 13 1 9 1 10 11 11 12 1 11 1 10 9 1 11 11 2 1 10 11 2 0 9 1 11 2
18 3 1 11 7 11 2 13 15 1 10 12 9 3 0 1 10 9 2
19 3 15 13 10 0 9 1 8 2 8 10 15 3 13 3 1 10 9 2
25 10 11 13 3 10 9 2 11 11 11 11 2 2 1 10 15 4 4 13 1 12 10 0 9 2
52 11 2 9 1 8 8 8 8 8 8 11 8 8 8 2 1 9 9 0 13 0 9 0 0 0 7 9 1 9 2 13 10 9 0 1 10 11 0 1 10 9 1 10 9 11 2 8 8 8 8 2 2
27 3 4 13 15 16 10 9 0 1 10 9 13 10 2 9 0 2 3 15 13 10 10 9 1 10 9 2
17 3 10 9 13 10 9 1 10 16 9 1 9 15 13 10 9 2
6 9 0 7 9 0 2
42 10 9 1 10 9 2 1 0 13 1 9 7 9 0 1 10 9 2 16 13 10 0 9 2 13 10 0 9 1 9 0 3 1 10 9 0 2 0 1 10 9 2
21 3 3 0 13 10 9 1 10 9 1 10 9 2 3 0 13 1 9 10 9 2
46 11 13 9 1 10 11 1 11 1 10 11 7 1 10 9 1 12 13 10 9 1 10 11 1 10 11 11 1 10 9 1 11 2 13 15 1 10 0 9 1 9 0 1 10 9 2
23 1 16 10 9 4 13 3 1 15 1 10 15 2 4 7 13 3 10 9 1 10 9 2
21 10 9 13 10 9 2 15 1 10 9 0 7 1 10 9 7 9 1 10 9 2
13 11 13 1 10 9 1 13 15 1 10 0 9 2
41 10 0 9 1 11 2 13 10 0 9 7 13 3 0 2 13 9 1 15 13 15 7 11 15 13 3 3 2 10 9 13 3 0 7 10 9 1 9 13 0 2
33 10 9 0 11 11 13 16 2 1 10 13 15 2 2 1 10 0 9 2 11 13 1 3 0 7 10 10 9 3 16 15 2 2
11 2 15 13 9 1 11 11 7 11 11 2
32 1 11 11 2 10 9 1 10 9 2 10 9 11 4 13 1 9 0 13 9 0 1 10 9 0 7 0 16 3 13 13 2
12 10 9 15 13 1 3 1 10 9 1 9 2
43 15 16 13 4 13 1 10 9 1 10 9 1 11 1 12 2 15 1 10 9 13 12 9 13 1 9 7 9 1 11 15 16 15 4 13 1 10 9 13 1 10 9 2
44 10 9 1 13 9 13 10 16 1 11 13 13 15 1 10 9 7 13 10 16 2 3 2 13 10 9 16 3 13 1 3 0 7 16 13 1 15 0 1 10 9 1 9 2
27 10 9 13 3 9 1 10 11 2 10 9 1 9 1 9 16 13 13 1 9 0 9 2 9 7 9 2
16 10 9 13 0 2 10 9 10 9 7 10 9 10 0 9 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
24 3 11 13 10 9 1 10 9 1 10 9 3 7 10 11 15 13 10 9 1 10 0 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
23 10 9 4 13 1 12 7 10 9 3 15 13 7 12 9 0 2 13 13 2 1 12 2
28 1 10 9 16 13 9 1 11 2 12 2 2 11 13 1 10 9 0 2 10 9 0 0 1 10 9 12 2
35 1 9 0 2 11 11 13 10 12 1 11 1 10 9 1 10 9 0 2 16 3 13 10 9 1 9 1 10 9 16 13 1 10 9 2
26 3 1 10 9 1 10 9 11 2 10 9 13 10 9 1 10 9 7 10 9 13 1 13 10 9 2
20 2 11 11 2 13 10 9 0 1 9 7 9 16 13 1 9 1 10 9 2
28 11 2 1 12 5 5 2 13 10 0 9 3 0 1 10 9 7 10 0 0 1 3 1 9 1 10 9 2
62 10 9 1 9 0 9 1 9 0 13 1 13 2 3 2 10 12 0 9 2 10 3 0 2 3 1 12 7 12 9 2 1 10 9 1 12 16 13 10 9 1 9 7 16 2 3 2 13 10 9 9 0 0 2 9 1 9 7 10 9 0 2
17 13 1 10 11 1 10 11 1 11 2 13 1 10 11 1 11 2
30 1 10 9 13 11 11 2 11 2 11 2 10 11 2 11 7 11 1 9 1 9 7 3 16 13 1 10 9 0 2
21 10 9 4 13 7 1 10 11 7 3 1 10 11 1 11 16 15 13 1 0 2
56 11 11 1 10 9 1 11 1 10 2 9 1 10 9 1 11 2 13 10 9 0 1 10 9 0 2 2 0 9 3 1 12 13 0 16 2 3 3 2 13 10 9 1 10 9 1 10 9 7 16 15 15 13 1 3 2
22 11 11 11 2 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 0 0 2
41 10 9 1 9 4 13 1 10 9 11 1 11 11 2 1 10 9 1 10 9 1 10 9 11 1 10 0 9 1 10 9 11 11 11 1 3 13 9 1 9 2
19 10 9 13 1 9 10 9 1 9 1 10 9 1 10 9 1 9 0 2
16 10 9 4 3 13 1 10 9 11 11 11 9 1 10 9 2
28 10 9 4 13 1 11 11 7 4 13 3 1 11 7 3 1 16 15 13 2 11 7 11 13 13 10 9 2
8 13 1 11 1 11 1 12 2
34 1 9 1 10 9 7 9 1 10 9 0 0 1 10 9 11 8 9 2 7 13 1 10 9 11 11 2 10 9 3 13 0 9 2
16 1 11 15 13 1 11 1 12 1 10 9 0 0 11 11 2
8 13 3 10 9 1 11 13 2
7 10 9 13 3 3 0 2
34 11 15 13 1 9 1 12 7 3 3 4 1 13 1 11 2 3 13 1 11 11 2 13 1 10 9 1 10 9 1 10 9 9 2
34 11 11 2 12 1 11 1 12 2 9 1 10 11 2 11 2 11 2 13 10 9 2 9 7 9 0 13 3 1 11 2 11 2 2
32 4 13 15 1 9 2 2 13 9 1 10 9 11 11 2 1 10 9 1 9 1 11 11 1 10 9 1 11 2 9 2 2
5 13 1 12 9 2
17 10 0 9 13 1 11 11 8 7 13 1 9 1 10 0 9 2
25 1 9 1 10 9 2 13 10 9 0 2 7 4 13 9 1 10 9 1 13 13 10 9 0 2
35 11 13 1 15 1 10 9 3 0 1 11 11 1 0 9 2 10 11 11 11 2 13 1 12 1 10 11 11 11 11 7 11 11 11 2
31 13 10 9 0 2 0 9 0 1 11 11 7 9 1 10 9 11 2 10 9 7 10 11 13 1 11 11 7 11 11 2
20 10 9 3 0 1 10 9 13 3 9 1 10 9 1 10 9 2 10 11 2
20 11 11 2 9 1 10 9 11 2 13 1 9 13 1 10 9 2 11 2 2
16 1 9 3 0 2 4 13 0 9 7 9 13 1 10 9 2
37 10 9 1 10 9 3 13 9 2 1 9 0 2 7 10 9 13 1 9 0 2 3 0 0 2 0 7 0 2 3 1 10 0 9 0 2 2
20 10 9 4 13 10 0 11 11 1 12 7 13 12 9 1 11 0 1 12 2
16 10 9 15 13 1 10 9 1 10 9 0 1 10 9 0 2
25 1 12 2 10 0 9 8 2 11 1 10 11 13 10 11 11 1 10 9 1 10 9 2 9 2
15 1 10 9 0 0 2 10 9 15 13 1 12 9 0 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 4 1 9 0 7 2 12 5 2 12 9 5 13 9 2
20 11 13 1 16 3 13 15 15 13 1 10 9 2 15 10 9 13 10 9 2
76 9 0 0 13 10 9 15 13 1 10 9 0 1 11 2 11 2 11 7 11 2 11 2 11 7 11 11 2 15 15 10 9 0 13 1 9 1 9 0 0 1 10 9 2 7 15 1 10 9 0 15 13 1 10 9 1 9 0 2 11 2 2 9 0 9 2 11 2 7 9 0 0 2 11 2 2
27 1 12 10 9 11 11 1 10 11 15 13 1 9 1 15 2 13 3 10 0 9 1 11 7 10 11 2
14 13 0 7 15 13 0 2 7 3 13 15 16 13 2
43 4 13 1 15 1 10 9 11 11 11 2 11 11 2 11 2 11 2 10 9 1 12 9 2 13 3 1 10 9 1 11 11 7 11 10 11 2 2 7 11 11 11 2
15 4 13 3 10 0 9 1 11 2 1 11 1 10 9 2
38 13 3 3 1 10 9 0 7 15 13 9 1 10 9 2 13 3 0 13 3 1 13 1 10 12 1 10 9 7 13 0 1 10 12 1 10 9 2
26 10 9 13 10 9 1 11 11 2 11 1 11 2 2 13 10 9 1 10 10 9 13 1 10 9 2
60 15 13 1 12 9 2 15 3 13 1 10 9 1 9 1 9 1 9 1 9 1 10 9 0 0 1 9 1 10 9 1 10 9 0 7 0 1 10 9 1 9 2 1 10 9 13 1 10 9 2 1 10 9 1 10 9 1 0 9 2
14 13 12 9 1 10 9 0 1 12 9 2 9 5 2
14 3 2 10 9 4 13 10 9 0 13 11 11 11 2
24 10 9 1 9 0 4 13 1 12 2 1 10 9 1 10 9 1 11 11 2 11 7 11 2
31 15 16 4 13 10 9 1 10 11 13 10 9 0 13 9 1 10 9 7 13 13 12 9 1 10 9 16 4 13 3 2
34 1 10 9 13 0 2 15 13 1 9 2 15 13 1 10 9 9 2 11 2 7 15 15 13 10 9 1 9 2 9 0 7 9 2
25 11 11 13 10 9 1 11 2 13 1 10 9 1 11 11 2 16 13 10 9 0 1 10 9 2
34 10 9 13 1 10 9 3 3 7 0 2 3 7 1 3 1 13 11 11 3 4 1 13 16 13 0 7 0 1 13 1 10 9 2
18 10 9 13 10 9 1 10 9 1 10 9 1 16 15 13 1 15 2
46 1 10 9 1 12 2 10 11 11 1 11 4 1 13 1 13 10 0 9 1 10 9 1 9 2 1 0 9 1 13 13 1 10 9 1 9 13 3 9 1 10 9 7 10 9 2
29 10 9 1 11 11 2 1 9 2 11 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
56 10 9 13 9 1 10 9 11 11 16 15 13 3 0 13 2 1 10 9 1 10 9 1 11 2 1 10 9 1 11 10 9 1 9 0 2 10 0 9 0 2 2 13 1 9 1 11 11 11 7 10 9 1 10 11 2
31 10 9 15 13 1 10 9 0 1 11 11 7 13 9 1 10 9 2 8 5 11 11 11 2 9 1 8 11 11 11 2
25 1 9 1 10 9 1 10 9 7 9 2 10 9 1 8 2 9 7 10 9 15 13 3 0 2
18 1 9 0 10 9 13 10 9 0 2 0 2 0 1 10 0 9 2
14 3 13 1 11 11 2 1 10 15 4 13 15 3 2
16 3 13 12 10 9 0 13 7 13 1 11 1 11 7 11 2
22 13 10 9 1 11 11 2 9 1 11 11 2 1 10 9 1 11 2 2 11 2 2
23 11 2 11 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 13 10 9 0 2
14 10 9 1 10 9 15 13 3 1 10 9 1 9 2
8 3 13 1 10 0 8 11 2
42 10 9 13 1 9 16 10 9 16 13 10 9 1 10 11 11 2 15 13 1 10 9 1 13 1 9 1 10 9 0 7 3 13 13 10 9 1 9 0 7 0 2
16 1 10 9 12 13 10 9 1 13 13 10 9 1 10 9 2
41 3 3 13 9 16 10 9 1 11 1 11 13 1 10 0 9 1 11 2 7 1 9 2 10 9 1 10 15 10 9 13 10 9 1 10 11 15 13 1 11 2
17 10 11 1 11 11 13 10 9 13 1 11 11 2 11 2 11 2
23 4 13 9 1 10 9 1 9 1 10 9 1 10 9 1 9 1 10 11 2 11 11 2
25 11 11 7 11 11 13 10 9 1 10 9 16 13 2 1 0 9 2 10 9 0 1 0 9 2
16 10 9 13 1 11 11 2 11 11 2 11 11 7 11 11 2
14 10 9 1 10 9 13 13 10 10 9 7 13 9 2
28 10 9 1 10 11 13 10 9 0 7 9 0 1 10 11 11 7 10 9 1 11 1 10 11 11 1 12 2
26 1 9 10 0 9 1 11 13 1 9 10 9 1 10 0 9 2 0 9 7 0 9 1 10 9 2
31 1 12 13 10 9 0 0 2 1 10 15 3 13 11 11 2 1 10 15 13 8 2 11 2 9 1 10 9 1 12 2
13 10 9 4 4 13 1 9 7 13 10 9 0 2
17 10 11 11 11 13 10 9 1 9 1 11 1 10 9 1 11 2
15 10 9 13 0 7 0 9 2 0 1 10 9 1 9 2
35 1 12 9 1 9 10 9 0 2 10 9 11 11 2 13 10 9 1 10 9 0 1 15 9 1 10 9 2 1 13 3 1 12 9 2
14 13 13 0 1 10 15 3 3 13 10 11 2 11 2
38 1 9 1 10 9 15 4 13 1 9 1 10 11 1 10 11 2 15 13 13 10 9 15 13 10 9 1 10 9 1 11 1 10 9 1 9 0 2
39 10 11 13 10 9 0 7 0 0 13 1 10 9 1 11 2 1 10 9 1 9 11 2 3 7 4 13 1 11 11 1 10 11 1 11 11 1 12 2
60 10 9 11 1 11 2 12 5 2 7 11 1 11 11 2 12 5 2 13 13 1 10 9 16 3 13 3 1 12 9 1 9 2 7 1 15 13 9 0 1 10 9 1 9 1 10 12 1 10 12 7 1 10 12 1 10 12 1 11 2
42 3 1 10 12 7 12 9 1 11 2 10 9 13 10 0 9 1 10 9 2 11 2 10 9 1 11 2 2 7 10 0 9 2 11 2 11 2 2 10 9 0 2
48 10 9 2 10 9 2 9 7 10 9 2 13 9 1 10 9 0 1 10 9 1 10 9 12 2 10 15 1 10 0 9 2 7 10 9 15 13 1 13 0 9 1 9 2 16 13 11 2
20 13 10 9 11 1 10 9 0 1 9 1 12 1 10 9 1 10 9 0 2
14 3 13 15 0 15 13 10 9 1 10 9 1 11 2
13 13 12 9 1 10 9 1 10 9 1 12 9 2
18 15 13 1 10 9 1 16 11 13 2 7 13 2 2 10 9 2 2
12 15 13 1 10 9 1 0 9 13 11 12 2
25 13 15 1 10 9 2 10 9 10 11 11 13 1 10 9 1 10 9 1 13 1 10 12 13 2
22 1 10 0 9 12 15 15 13 3 0 9 15 16 13 9 1 10 9 1 12 9 2
43 10 9 1 10 11 3 4 13 3 10 9 1 10 9 0 1 10 9 2 1 10 15 10 9 13 3 0 2 1 9 1 10 9 1 10 9 7 1 10 9 1 9 2
9 10 9 1 10 9 13 10 9 2
33 10 9 3 13 2 10 0 9 1 13 15 13 10 9 1 9 2 7 13 16 1 10 13 3 0 13 9 16 1 0 15 13 2
64 3 13 1 3 3 2 10 12 1 11 1 12 2 16 15 13 3 10 9 0 1 10 9 1 10 9 2 11 2 1 10 9 0 1 10 9 1 11 2 3 15 13 0 9 7 15 13 10 10 9 0 0 1 13 1 10 9 1 10 9 0 1 9 2
13 11 2 13 10 9 1 9 0 1 10 9 11 2
50 11 4 13 1 11 2 7 3 1 10 9 2 13 1 10 10 9 11 1 16 13 1 11 7 15 13 13 15 13 10 9 7 1 15 15 13 1 11 11 7 4 0 13 1 10 9 1 15 3 2
20 1 10 9 2 3 15 13 15 13 10 9 2 13 1 9 2 2 9 2 2
28 1 10 9 11 11 13 10 9 1 10 9 0 16 4 1 4 13 10 9 1 10 9 0 1 10 9 0 2
34 13 10 9 1 10 12 5 1 10 9 7 10 12 5 1 9 1 10 9 2 9 2 9 1 10 9 0 7 9 1 9 1 9 2
22 10 9 0 13 0 9 1 10 9 0 2 15 4 4 13 1 7 10 9 13 0 2
39 10 9 11 1 10 11 11 11 2 16 13 11 11 2 4 4 1 4 13 1 10 9 11 15 3 15 4 13 10 9 0 1 10 9 1 10 9 12 2
26 10 9 1 11 2 9 1 2 13 1 0 9 1 11 11 2 10 9 0 1 10 9 1 10 9 2
14 4 13 0 1 10 9 1 9 1 11 1 12 9 2
11 2 11 2 4 13 7 13 1 11 11 2
25 4 13 1 9 7 9 1 9 2 1 10 9 13 1 10 9 2 1 9 0 7 9 1 9 2
79 10 9 1 9 1 9 2 11 11 11 2 4 13 10 9 1 16 10 9 2 4 1 13 15 2 1 13 1 2 11 7 11 2 2 3 15 13 10 9 0 1 10 9 1 10 8 1 13 12 9 2 7 4 13 3 16 10 9 1 11 13 16 11 4 13 1 9 2 16 10 8 13 9 2 16 3 0 2 2
19 1 13 10 9 1 9 10 0 9 13 13 7 13 9 13 1 10 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
32 2 3 15 13 10 9 2 1 10 9 2 1 16 13 1 10 9 1 10 9 12 9 3 16 3 15 13 10 9 16 13 2
16 10 0 9 1 9 2 12 1 12 2 15 13 1 9 0 2
18 10 9 3 4 4 13 1 11 1 12 2 7 3 4 13 1 3 2
20 1 10 9 15 13 10 9 1 9 1 11 16 13 1 11 1 10 9 0 2
26 13 12 9 0 1 10 11 0 1 10 9 2 13 10 9 1 12 15 11 11 13 1 12 7 12 2
17 10 9 0 4 13 9 7 13 2 13 7 13 2 1 9 0 2
49 13 3 9 0 1 10 11 11 2 11 2 12 2 2 1 10 9 1 10 9 11 2 0 9 1 10 9 0 9 1 10 9 2 10 3 0 11 11 11 2 7 10 11 2 11 2 12 2 2
21 10 9 13 10 0 9 1 10 9 0 3 0 1 10 9 1 9 0 3 0 2
12 15 4 13 10 9 16 15 4 13 10 9 2
12 1 10 15 15 13 10 0 9 1 10 9 2
42 10 9 3 0 15 15 13 11 11 1 10 12 2 12 3 16 10 9 3 0 15 15 13 10 9 11 11 1 10 12 2 12 2 3 3 10 10 9 13 10 9 2
30 10 9 1 11 11 13 1 10 9 7 10 9 1 11 2 9 15 13 10 9 7 3 13 9 1 9 0 7 0 2
20 10 11 4 4 13 1 9 1 9 7 13 10 7 15 9 1 10 9 0 2
17 10 9 1 10 9 1 10 9 13 0 7 13 1 10 9 0 2
17 10 9 13 1 0 9 7 1 10 9 16 13 3 13 10 9 2
26 10 0 9 13 7 13 10 9 1 9 0 13 4 13 1 10 0 9 1 9 1 9 7 9 0 2
31 13 10 9 1 9 1 9 1 12 1 10 9 1 9 1 11 11 11 3 11 13 1 11 11 7 11 2 13 0 9 2
19 11 11 13 10 9 0 1 10 11 1 11 2 9 1 11 11 2 11 2
28 13 16 10 9 3 4 4 13 7 13 3 13 1 10 10 9 15 13 1 10 9 7 10 9 1 10 9 2
29 10 9 1 11 11 2 1 9 2 11 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
26 3 4 1 13 9 1 10 9 1 11 1 12 1 12 2 1 10 0 9 1 11 11 11 7 11 2
17 1 10 9 0 1 10 9 2 10 9 0 1 10 9 13 0 2
16 10 0 9 13 16 10 11 13 1 10 9 3 1 12 9 2
29 13 10 9 0 1 10 0 9 1 10 9 2 10 9 1 10 11 2 3 15 4 13 3 10 9 16 10 9 2
47 13 10 9 1 16 10 9 15 13 1 3 0 2 11 11 13 1 9 0 2 2 1 10 9 0 10 9 1 13 10 9 4 4 13 1 9 2 3 1 10 9 0 1 10 9 2 2
35 1 10 9 11 11 2 16 4 13 9 1 9 1 10 9 1 9 7 16 13 1 10 9 1 10 9 1 10 9 2 10 9 13 0 2
15 10 9 15 13 1 10 9 0 1 10 15 13 12 9 2
34 10 9 0 15 13 10 9 1 10 9 4 13 2 13 10 9 13 1 10 9 1 9 0 2 1 11 11 2 1 10 9 1 11 2
42 10 11 11 0 2 11 11 2 13 10 9 1 9 1 10 9 11 2 9 1 10 9 0 1 10 9 0 1 10 9 1 11 1 10 9 2 1 10 9 1 11 2
12 15 13 10 9 1 9 2 7 13 1 15 2
28 10 9 1 9 13 1 9 10 9 1 9 9 2 10 9 1 9 13 1 3 10 12 5 2 16 13 11 2
16 3 2 11 13 1 10 9 1 11 2 13 1 10 9 11 12
21 1 10 0 9 2 1 12 15 13 10 0 9 16 13 1 11 1 9 1 11 2
42 13 9 1 11 1 11 7 11 2 8 2 2 9 1 11 1 11 7 9 1 11 1 11 11 7 1 11 2 9 1 11 11 1 11 7 11 2 12 9 1 11 2
27 10 9 1 10 9 1 11 11 15 13 3 3 0 2 3 10 9 1 11 15 13 13 1 10 0 9 2
25 10 9 1 9 13 1 12 9 7 3 1 10 12 5 1 10 9 13 1 10 9 1 9 0 2
19 1 10 9 1 9 13 10 9 0 10 9 11 7 10 9 2 10 11 2
10 10 9 0 13 13 10 9 1 9 2
18 1 15 13 0 1 13 10 9 0 1 13 15 7 13 1 10 9 2
18 1 10 9 0 11 1 11 2 10 9 1 11 13 9 1 9 0 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
38 16 11 3 13 13 9 1 10 9 2 10 9 1 10 9 13 1 16 11 13 1 10 0 9 1 10 9 7 13 10 0 9 1 10 9 1 11 2
15 10 9 13 3 2 15 3 0 7 13 1 10 9 0 2
17 1 12 13 10 9 11 11 1 9 0 13 1 10 9 1 11 2
23 10 0 9 13 1 10 9 1 11 7 11 13 1 3 1 12 9 1 10 9 1 11 2
18 10 9 1 3 12 5 1 0 2 9 1 12 5 1 0 2 9 2
16 1 10 0 9 15 13 1 10 9 1 11 10 9 1 9 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
13 4 13 3 1 15 1 10 9 7 3 1 3 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
31 4 13 1 13 10 9 1 10 9 0 1 10 9 0 1 11 11 1 12 2 3 1 9 0 1 10 9 0 11 11 2
41 1 10 9 0 1 11 11 11 15 13 10 9 1 11 11 1 11 11 11 2 7 1 10 9 0 4 13 10 9 0 1 10 9 1 11 11 2 11 10 11 2
22 1 10 9 0 3 13 10 9 1 9 7 1 0 2 7 1 9 7 1 0 9 2
22 11 4 13 10 9 0 1 10 9 1 10 9 1 10 0 9 1 10 9 1 11 2
45 10 9 15 13 1 10 9 1 9 2 1 10 15 13 10 9 0 2 10 9 1 9 2 7 9 2 7 16 1 10 9 10 9 0 13 10 9 1 9 7 10 9 1 9 2
21 1 10 9 15 13 2 3 10 9 1 10 0 9 1 10 11 1 11 7 13 2
46 10 9 1 13 15 13 1 4 13 10 9 0 3 7 4 13 10 0 9 16 13 10 9 11 2 1 10 9 7 15 13 10 0 9 7 9 16 15 13 3 1 10 9 1 9 2
38 10 9 15 13 1 10 11 2 12 7 10 11 2 12 7 15 4 13 1 10 9 13 11 11 11 11 2 7 3 10 11 2 12 13 1 13 15 2
21 1 10 9 12 10 9 13 10 0 9 2 1 10 9 1 10 9 1 10 9 2
33 1 10 9 0 13 1 12 13 7 15 13 10 15 1 10 9 2 7 15 1 15 3 2 16 10 9 13 3 13 1 10 9 2
26 1 10 0 9 2 1 10 9 3 0 1 10 11 11 13 0 10 9 7 2 1 9 2 10 9 2
46 1 9 2 9 11 11 15 13 10 9 1 9 1 11 11 1 10 11 7 4 13 1 11 1 12 2 1 8 12 1 10 9 2 10 9 1 10 9 1 10 9 0 11 11 11 2
53 4 13 1 11 11 11 11 2 11 11 7 11 11 7 13 1 11 11 2 16 3 13 10 9 0 7 13 9 1 10 9 0 1 10 9 2 0 1 11 11 2 11 11 11 2 11 11 7 10 0 11 11 2
43 10 0 9 4 13 16 10 9 4 4 13 1 10 9 0 1 11 1 11 16 13 1 13 1 11 10 9 0 13 1 10 9 1 10 9 0 3 1 10 9 1 11 2
14 1 10 9 1 11 3 3 15 4 13 10 9 0 2
16 13 0 1 10 9 1 10 9 2 10 12 1 10 0 9 2
27 1 13 15 10 0 9 1 8 15 13 1 10 9 2 1 11 15 4 13 10 9 11 1 10 8 3 2
27 1 9 1 9 10 9 1 9 0 15 13 3 1 9 1 9 3 0 2 15 1 9 1 9 7 9 2
34 13 1 11 11 2 11 7 11 11 2 10 9 13 10 9 1 9 1 10 9 11 0 7 10 9 1 9 1 10 9 11 1 11 2
44 11 2 9 1 10 11 11 13 1 10 9 0 10 12 9 1 9 2 10 9 16 13 1 13 1 10 9 16 4 13 15 1 13 1 0 10 9 10 9 0 1 10 11 2
11 3 13 1 10 11 11 1 0 9 0 2
10 1 12 13 10 0 9 13 1 11 2
20 13 1 10 9 1 9 3 15 13 10 9 1 9 1 10 9 1 10 9 2
12 11 7 9 1 11 2 11 2 11 7 11 2
28 10 9 2 9 2 8 8 8 2 7 2 8 2 2 13 10 9 0 13 3 1 11 2 3 13 9 0 2
51 3 1 10 9 1 9 2 11 11 11 13 3 10 9 1 9 2 13 10 9 1 9 1 9 0 7 4 13 1 10 9 1 9 1 9 1 11 11 1 10 11 7 1 9 1 9 1 10 11 11 2
21 10 12 1 11 2 13 15 1 10 9 13 1 2 10 9 2 2 11 11 2 2
15 10 11 11 1 11 1 12 4 13 1 10 11 1 11 2
10 13 1 10 11 1 12 9 13 0 2
17 10 9 13 1 3 1 12 9 1 0 9 7 1 10 10 9 2
59 1 10 0 9 1 10 9 2 10 9 1 11 1 11 2 11 11 13 10 9 11 11 1 10 9 11 11 2 15 4 4 13 1 9 1 0 2 7 13 16 15 13 13 3 1 3 1 11 11 16 13 10 9 1 9 1 10 9 2
45 1 9 1 11 2 11 2 13 15 3 0 7 0 1 4 13 10 0 9 1 11 2 13 10 9 7 15 13 1 11 13 1 10 9 1 10 9 1 13 1 9 10 9 0 2
48 10 9 2 11 11 11 11 11 2 15 4 13 1 10 9 1 10 9 2 11 11 2 11 2 2 7 3 13 9 1 11 11 2 10 9 16 13 1 10 9 1 2 11 11 2 11 2 2
29 16 10 0 9 13 10 1 11 2 1 10 9 13 3 10 9 0 2 9 2 1 11 2 11 7 11 2 11 2
15 10 9 0 13 1 12 9 1 9 0 2 8 5 2 2
20 10 9 16 13 10 9 1 11 1 10 9 1 10 9 1 10 9 4 13 2
38 10 0 12 9 1 9 2 10 9 1 10 9 16 13 1 10 9 10 11 1 11 7 11 2 15 4 13 1 10 3 9 1 10 2 12 9 2 2
37 13 9 1 10 9 7 13 1 13 1 10 9 1 10 9 1 9 2 15 13 14 11 1 10 9 7 9 0 15 13 1 10 9 1 10 9 2
11 1 12 13 1 10 11 1 9 7 9 2
48 10 9 2 11 2 2 10 9 1 9 1 13 9 0 2 4 4 13 1 2 0 2 1 10 9 11 11 2 10 15 15 4 13 1 10 9 1 10 2 0 9 1 10 9 1 11 2 2
24 4 13 7 13 10 9 15 16 13 13 9 0 2 3 0 2 13 1 0 9 7 0 9 2
52 10 9 13 16 10 11 3 4 13 9 16 13 10 9 1 9 0 7 10 9 1 10 9 0 2 3 7 16 13 10 0 9 1 10 9 0 7 13 3 10 9 1 10 9 0 1 9 1 13 1 12 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 12 2
36 15 4 13 9 0 9 1 10 9 1 11 2 9 11 2 11 2 9 2 11 2 11 2 7 3 1 10 9 0 1 11 11 1 10 11 2
58 10 9 2 15 13 1 10 9 1 13 1 10 9 2 7 1 10 9 15 13 1 13 15 1 10 9 1 10 9 2 3 16 11 2 13 1 10 10 9 0 1 10 11 1 10 9 2 7 13 0 1 13 1 11 7 10 9 2
75 1 9 1 10 9 4 13 1 10 9 1 10 15 13 3 0 2 15 13 1 11 7 13 13 15 2 15 3 13 2 10 9 4 13 3 0 2 15 13 0 1 10 9 1 0 9 2 4 13 1 9 2 1 10 9 1 13 10 9 13 3 0 16 10 9 13 9 2 7 1 11 15 4 13 2
37 1 12 7 12 15 13 1 10 9 1 10 9 10 9 11 2 16 13 2 11 2 2 9 16 13 16 1 12 10 9 4 13 1 10 9 0 2
31 13 10 9 1 9 1 10 9 1 10 9 1 10 9 16 13 13 15 1 10 0 9 16 15 13 10 11 1 10 11 2
31 1 9 12 7 1 3 4 13 15 2 15 10 9 7 9 16 13 7 15 13 16 3 15 4 13 2 16 15 13 3 2
59 10 0 9 7 0 9 2 11 2 13 10 9 0 1 11 2 13 1 10 0 9 1 11 11 2 1 11 11 11 2 2 3 9 1 10 11 1 11 2 1 9 1 10 9 11 2 11 2 2 11 2 11 2 7 11 2 11 2 2
13 3 2 15 15 13 1 10 11 1 11 1 12 2
5 3 7 15 13 2
10 13 12 9 0 1 11 7 13 0 2
6 4 13 1 11 11 2
18 10 9 13 9 1 10 0 9 0 1 10 9 1 10 0 12 9 2
19 11 11 13 16 3 4 13 9 1 10 9 0 2 16 13 10 9 0 2
14 1 3 1 3 2 10 9 13 1 13 10 0 9 2
33 1 10 9 1 11 2 11 11 2 2 10 9 1 11 1 9 1 10 9 1 10 9 0 13 3 3 3 1 10 9 0 2 2
37 10 9 1 9 13 3 1 9 2 7 13 13 15 1 10 9 0 2 7 15 13 1 7 2 2 2 10 9 13 0 7 3 1 9 0 2 2
20 1 11 2 10 9 0 13 1 13 10 9 1 9 1 10 9 1 10 15 2
44 10 9 3 4 13 10 9 0 1 10 9 1 10 9 2 7 10 9 13 10 9 1 9 0 1 10 9 1 10 11 2 7 10 9 0 1 10 9 0 7 1 10 9 2
33 1 9 1 10 0 9 0 2 10 9 0 1 10 9 15 13 2 1 11 13 2 11 11 11 11 2 16 15 13 3 10 9 2
11 10 9 1 11 15 13 10 12 2 12 2
32 10 9 15 13 1 10 0 5 12 1 10 11 11 2 7 13 15 1 10 0 9 1 9 2 13 9 1 9 1 10 9 2
19 1 10 9 13 1 10 9 1 15 7 11 11 1 10 9 11 15 11 2
26 13 1 10 9 0 13 16 10 9 3 0 13 10 1 13 10 9 2 13 1 9 7 3 13 15 2
34 1 10 9 1 11 2 12 2 10 5 2 12 11 2 13 3 1 10 9 7 10 9 1 10 11 11 2 3 13 13 1 9 0 2
18 1 12 2 1 10 0 9 0 2 10 9 13 7 10 9 13 3 2
20 10 9 13 9 1 9 0 1 9 7 9 1 10 0 11 1 10 9 0 2
48 1 10 9 1 9 13 2 11 11 11 2 2 2 11 11 11 11 2 11 11 11 2 2 2 11 11 2 2 2 11 2 7 3 2 11 11 2 1 10 9 12 2 3 15 13 10 9 2
40 10 9 1 9 1 10 11 1 11 15 13 1 9 1 10 9 13 1 10 9 1 10 9 7 13 10 9 1 9 9 1 9 13 1 9 0 1 9 0 2
5 1 12 13 12 2
45 13 1 10 9 1 11 2 10 9 13 10 9 1 10 9 7 10 9 1 10 9 2 10 9 2 10 9 1 10 9 1 9 1 9 7 10 9 0 1 10 9 7 10 9 2
15 1 10 9 1 10 11 13 3 10 9 1 9 13 0 2
31 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 5 12 2 7 10 9 0 1 9 13 5 12 2
12 1 10 9 12 11 11 13 10 9 1 11 2
7 3 4 1 13 3 3 2
22 15 13 9 16 16 15 13 10 9 2 10 9 13 1 10 9 13 3 0 10 9 2
26 11 11 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 13 10 0 2 9 0 13 0 2
13 1 10 9 1 12 2 11 11 4 13 10 9 2
18 1 10 9 2 11 7 11 11 13 10 12 5 1 10 9 1 11 2
26 10 9 13 10 9 1 9 11 11 2 12 1 9 0 2 11 11 12 7 10 11 11 1 9 0 2
16 10 0 9 13 10 0 9 1 9 1 10 11 7 10 9 2
42 16 4 13 3 1 11 11 11 2 16 15 13 1 12 2 10 11 4 13 1 0 9 1 10 2 11 11 2 10 12 1 11 1 12 2 3 3 1 10 9 0 2
24 13 9 13 1 10 9 1 11 7 4 13 16 4 13 15 1 10 9 16 3 4 13 3 2
48 10 12 1 11 1 12 15 13 10 9 1 10 9 11 1 10 9 1 10 3 9 0 1 10 0 7 0 11 7 11 1 9 1 10 9 11 1 10 9 7 11 0 1 10 9 1 11 2
26 10 9 1 10 9 13 1 13 10 9 1 9 1 10 9 0 1 10 9 0 1 15 13 10 9 2
9 13 10 9 7 4 13 1 11 2
16 1 15 16 13 9 0 2 15 13 1 10 9 1 10 9 2
21 10 9 15 13 13 1 9 2 10 11 3 0 7 10 9 1 10 9 3 0 2
23 1 10 0 9 13 10 9 12 9 2 13 3 10 9 0 2 1 12 2 7 12 9 2
36 10 9 13 3 1 11 2 3 7 10 11 4 7 13 3 10 11 15 13 2 7 1 9 0 2 10 9 2 9 1 11 2 10 0 11 2
40 3 1 10 12 7 12 1 10 9 1 10 11 2 10 9 13 1 16 15 4 13 10 9 1 10 9 1 11 7 16 10 9 13 1 9 1 10 11 11 2
18 15 13 1 10 9 1 12 9 1 12 9 1 10 9 0 2 11 2
15 1 11 15 13 2 16 3 4 13 10 9 2 10 9 2
28 1 9 0 10 9 0 7 9 4 1 13 15 2 10 9 1 13 1 10 9 0 7 10 9 1 9 0 2
41 10 9 1 10 9 1 15 9 13 3 0 16 10 9 0 1 15 1 11 1 11 7 10 11 11 1 11 13 1 10 9 7 10 9 1 9 13 1 10 11 2
21 1 10 9 2 10 9 1 10 9 7 9 0 3 15 13 9 1 10 9 0 2
40 1 10 9 1 9 13 3 16 10 9 13 16 10 11 2 1 10 12 2 4 13 1 10 11 10 9 13 1 13 1 11 11 2 1 9 1 10 11 0 2
8 11 15 13 13 1 10 9 2
25 11 13 1 11 1 16 15 13 2 7 15 3 13 1 10 9 13 15 3 1 10 9 1 9 2
66 1 15 2 11 11 1 0 13 13 13 1 15 15 11 2 11 13 1 11 11 2 11 2 7 13 3 2 1 10 9 11 11 15 13 10 9 1 10 12 9 2 11 7 11 2 2 1 3 13 15 1 11 10 9 1 11 2 0 9 1 10 9 9 1 11 2
43 1 9 2 13 10 9 1 10 2 11 11 2 2 3 10 9 1 10 13 10 9 1 10 11 2 13 16 10 0 9 13 13 1 10 9 1 11 11 1 10 11 11 2
30 1 9 2 10 9 0 1 9 2 10 9 1 9 0 2 13 16 15 1 15 10 9 0 13 1 9 1 10 9 2
70 4 13 1 10 3 0 9 1 9 0 1 10 9 7 13 10 11 2 10 11 7 10 11 2 11 10 15 13 10 0 9 7 3 13 10 9 0 7 7 10 9 3 0 1 10 11 11 11 10 15 4 13 1 11 11 11 11 10 9 3 13 9 1 10 1 10 11 7 11 2
30 1 9 1 10 9 13 0 13 1 9 10 9 1 10 9 1 10 9 7 1 15 13 3 0 13 1 9 10 9 2
15 10 9 15 13 1 10 9 1 9 13 1 11 7 11 2
18 11 13 10 9 1 9 0 1 12 9 0 1 10 9 1 10 9 2
23 1 10 9 13 3 1 12 9 7 9 0 1 10 11 11 2 11 7 9 1 10 9 2
4 2 1 15 2
9 13 13 15 1 10 9 1 9 2
32 10 9 1 9 13 13 15 1 10 12 2 16 4 13 15 1 9 1 10 11 11 2 11 11 11 2 11 11 2 12 2 2
60 0 9 2 1 11 11 2 11 11 7 11 11 4 13 16 15 13 1 10 0 11 2 16 10 9 1 10 9 0 13 10 9 1 9 1 11 2 0 1 10 9 7 16 10 9 0 1 10 0 7 0 9 2 4 13 10 0 9 0 2
16 10 9 13 1 0 9 1 10 9 1 10 0 7 10 9 2
40 1 10 9 2 10 12 1 11 15 13 9 1 9 1 10 11 1 11 0 1 11 16 13 10 9 1 10 11 11 2 10 11 1 9 7 10 11 1 11 2
11 15 13 1 9 1 11 1 11 1 12 2
36 1 10 0 9 1 10 9 1 9 13 1 10 9 1 9 7 10 0 9 0 2 13 10 9 1 9 1 11 1 10 0 9 1 10 9 2
21 10 9 13 10 9 0 1 10 9 0 10 9 13 11 7 10 9 0 13 12 2
22 10 9 13 3 3 3 1 10 9 1 11 11 10 11 1 12 2 10 9 3 13 2
11 1 10 9 13 9 13 1 10 9 13 2
40 1 10 0 9 0 1 10 9 0 1 11 15 13 10 9 0 2 9 2 13 1 15 1 10 9 15 4 13 1 9 1 11 2 1 9 0 0 7 0 2
20 13 1 9 1 2 11 2 7 0 9 1 10 9 0 1 10 9 1 11 2
11 10 9 1 9 9 7 11 13 10 9 2
49 10 0 11 11 13 10 9 3 13 10 9 0 1 10 9 1 10 11 11 11 2 11 11 2 1 15 15 15 13 13 1 10 9 15 4 4 13 1 10 9 1 9 2 16 15 13 15 9 2
7 11 1 10 9 0 0 2
14 1 12 4 13 1 10 9 1 11 2 1 9 11 2
24 10 9 13 1 10 0 2 9 2 7 0 2 11 2 13 9 13 1 9 2 3 10 9 2
24 11 2 1 9 2 8 8 2 13 15 1 10 12 9 0 1 10 9 1 11 1 10 11 2
18 11 13 10 9 0 0 1 9 0 13 1 10 9 1 10 3 9 2
24 11 13 10 9 1 10 9 1 8 9 2 10 9 1 10 9 1 9 7 0 1 9 0 2
15 10 9 1 10 9 13 10 9 1 9 1 9 7 9 2
40 10 9 0 13 3 3 0 7 10 9 2 1 15 15 10 9 15 13 2 13 15 10 0 9 0 1 10 9 1 10 9 1 9 0 13 9 1 10 9 2
13 16 10 11 13 2 2 1 3 13 1 10 9 2
14 7 4 13 15 1 2 9 2 7 2 9 0 2 2
51 10 9 2 13 9 0 7 0 1 10 9 2 4 13 13 1 11 16 13 10 9 1 9 2 9 7 9 7 13 1 15 1 13 15 10 9 7 13 15 1 10 9 2 15 15 13 13 15 15 13 2
34 10 9 1 10 11 11 1 11 13 3 0 1 10 9 1 13 10 9 2 7 16 13 13 10 9 0 4 13 9 7 13 10 9 2
11 10 9 2 11 11 2 13 0 10 9 2
7 15 13 1 10 11 0 2
14 3 13 10 9 3 0 1 10 9 1 9 7 9 2
79 10 11 1 10 11 11 2 11 2 2 13 1 11 2 13 10 9 0 13 1 10 9 1 10 9 1 11 16 2 3 1 13 1 10 9 0 1 10 9 0 7 0 2 13 0 1 9 7 9 0 0 2 16 13 10 9 1 10 9 1 9 0 2 10 9 0 2 10 9 1 10 9 7 10 9 1 10 9 2
23 1 10 9 13 10 9 1 12 1 11 2 9 2 1 10 13 1 11 1 10 9 0 2
25 10 9 16 13 1 10 9 13 1 10 9 3 0 7 0 2 10 0 1 10 11 1 10 11 2
13 10 12 5 1 10 3 1 12 9 13 1 11 2
36 0 9 2 9 7 9 1 9 2 3 7 0 9 1 9 1 9 8 2 7 3 9 7 9 1 10 9 1 9 13 15 1 10 9 0 2
31 11 13 10 9 1 10 9 0 1 10 11 11 1 10 11 7 4 13 1 10 9 1 9 0 1 10 9 1 10 11 2
28 1 10 9 10 9 4 13 1 10 9 1 9 0 11 2 7 13 10 9 4 13 15 3 1 10 9 11 2
36 1 9 1 16 10 9 13 15 1 10 9 3 0 1 11 11 2 13 1 9 1 9 1 9 1 9 2 3 4 13 1 10 0 9 9 2
12 3 13 1 12 9 9 2 7 12 1 9 2
23 1 10 0 9 1 0 9 13 1 12 15 15 13 10 9 1 11 1 11 1 10 9 2
41 1 10 9 1 10 9 0 1 10 12 9 2 10 9 1 11 1 11 7 1 10 0 9 11 11 2 11 2 15 13 9 3 3 1 10 9 1 10 9 11 2
12 10 9 1 9 1 10 9 13 1 9 12 2
33 15 13 10 9 16 13 1 10 9 7 15 13 16 7 15 7 10 15 13 10 9 2 1 15 15 4 13 1 10 15 16 13 2
33 11 11 13 10 9 1 10 9 0 2 1 15 9 0 2 7 1 9 1 3 1 10 9 7 16 13 10 9 1 1 12 9 2
48 1 10 11 11 2 10 9 13 9 0 0 2 9 7 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 2 11 11 2 11 2 11 2 11 7 11 2 1 15 2
23 11 13 10 9 1 10 9 0 1 10 9 1 11 2 13 1 10 9 1 11 2 11 2
131 1 11 1 12 13 1 13 10 9 1 10 9 0 1 11 7 1 3 15 13 1 11 16 13 10 9 1 9 1 9 1 10 11 11 1 10 9 11 1 11 7 3 13 10 9 1 10 9 2 1 10 13 10 0 9 0 4 13 1 10 9 1 9 1 11 2 3 1 11 2 16 3 4 13 1 11 7 1 3 1 10 9 0 2 11 2 11 7 9 1 4 13 1 11 1 12 15 4 13 15 1 11 3 13 9 1 9 0 1 10 11 11 11 16 13 0 9 7 1 12 13 10 9 0 1 13 15 1 10 9 2
15 10 0 9 13 16 10 9 7 10 9 13 1 10 9 2
21 10 9 13 1 9 10 9 1 10 9 1 10 9 2 7 13 10 9 1 9 2
6 11 11 11 2 11 2
30 11 1 9 1 11 15 13 10 9 1 11 2 7 15 13 9 13 15 9 1 9 1 11 7 13 15 1 10 9 2
11 9 3 0 1 4 13 9 7 10 9 2
11 15 1 10 9 15 4 13 1 11 11 2
25 1 10 9 4 13 10 9 2 7 1 10 9 10 9 1 10 9 3 15 13 3 1 10 9 2
25 10 9 13 13 16 10 9 0 3 4 13 1 9 1 9 16 13 10 9 1 13 10 9 0 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
11 13 3 9 2 10 9 13 3 3 0 2
29 1 10 9 16 4 13 3 2 10 9 0 1 10 9 13 13 10 9 1 11 11 1 10 9 1 11 11 11 2
7 11 13 1 10 10 9 2
49 11 13 10 9 1 3 13 9 1 10 9 0 1 11 2 15 13 1 10 9 1 9 2 1 3 13 2 7 13 16 13 3 1 10 9 7 10 9 1 13 9 2 13 1 15 1 9 2 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
21 15 13 1 10 10 9 7 10 9 13 0 2 3 7 15 4 13 10 9 0 2
19 3 2 13 1 10 9 0 10 0 9 7 9 16 10 9 13 10 9 2
31 3 1 10 9 1 10 9 1 10 9 11 2 11 11 4 13 7 13 1 11 11 3 4 13 10 12 1 11 1 12 2
26 10 9 0 0 9 4 13 10 9 0 2 10 9 11 13 0 3 3 1 10 9 1 10 9 11 2
21 10 9 13 16 10 9 13 3 2 11 11 2 16 10 9 4 13 1 10 9 2
19 1 10 0 13 10 9 0 11 11 2 13 1 10 9 1 11 1 12 2
18 10 9 1 9 3 13 0 1 13 3 10 9 7 15 13 1 8 2
19 1 12 10 9 4 13 1 10 11 11 11 2 11 1 10 11 11 2 2
14 1 10 9 15 4 13 9 13 1 10 9 1 9 2
21 10 12 5 1 10 9 1 11 11 13 2 1 10 0 9 2 12 9 1 9 2
15 1 10 9 2 1 12 9 2 13 12 0 9 1 11 2
14 13 13 10 15 3 7 3 4 7 4 13 10 9 2
29 10 0 9 12 1 11 1 12 13 1 10 9 16 15 13 13 2 11 1 11 2 11 2 7 11 2 11 11 2
22 13 10 9 1 12 9 2 1 9 1 12 2 7 10 9 1 12 5 2 9 5 2
4 11 11 12 2
23 3 15 4 13 1 9 1 10 9 2 1 10 16 15 4 13 10 0 2 8 8 2 2
12 1 15 2 1 9 13 10 9 9 2 9 2
15 13 1 12 9 1 9 1 9 0 7 12 1 9 0 2
43 3 1 10 9 0 1 11 2 11 13 3 1 11 2 11 2 12 2 2 10 9 16 13 1 10 9 16 13 10 9 1 9 7 13 10 9 2 4 3 13 1 9 2
22 1 10 9 10 9 1 9 7 9 4 13 3 1 9 1 10 9 1 10 11 11 2
25 11 13 9 1 10 11 11 2 7 9 1 0 2 2 13 12 9 7 4 13 1 10 0 9 2
30 10 9 2 3 7 15 13 1 10 9 1 10 0 9 7 1 15 16 13 2 4 13 1 10 11 1 11 1 12 2
18 10 9 13 1 9 1 11 11 2 15 13 10 9 1 11 1 12 2
31 15 13 16 10 12 13 1 11 11 12 16 13 10 0 9 11 7 15 13 1 10 9 11 1 10 9 0 0 1 11 2
13 1 10 9 15 13 9 13 15 1 10 9 0 2
47 10 9 0 4 13 16 1 10 9 15 13 10 0 9 2 16 10 9 3 15 13 2 2 1 15 15 4 13 16 10 11 13 0 1 10 9 1 10 0 9 7 13 1 9 1 9 2
26 4 1 13 7 2 3 1 13 10 9 1 13 10 9 1 9 1 10 9 2 13 10 9 1 9 2
20 3 15 13 1 10 0 9 1 11 2 11 7 11 1 13 15 3 1 15 2
25 10 9 13 13 1 10 9 7 13 10 9 1 9 2 7 1 10 9 13 10 9 1 4 13 2
39 10 11 11 1 10 9 4 7 13 3 12 9 1 9 1 10 9 1 11 11 16 3 13 0 7 16 15 13 3 1 10 9 1 10 9 1 10 11 2
23 10 0 9 1 10 9 7 10 9 13 1 10 9 1 10 9 7 10 9 1 10 9 2
5 10 9 13 0 2
36 13 1 15 10 9 0 7 1 10 9 4 13 15 10 9 0 16 13 16 4 13 1 3 1 10 3 9 16 13 9 3 0 7 3 0 2
26 10 0 9 1 9 15 13 1 10 9 1 0 9 2 1 10 9 1 2 10 11 11 1 10 11 2
58 10 9 2 11 11 2 11 4 13 3 10 0 9 16 13 2 10 9 1 10 10 9 0 1 10 9 0 1 9 1 9 2 1 2 10 10 0 8 1 9 1 9 2 2 13 10 9 0 1 10 9 1 9 0 2 8 2 2
6 13 1 11 2 11 2
20 3 1 15 4 13 1 9 1 12 1 11 2 1 10 15 13 1 12 9 2
5 15 13 1 11 2
41 1 10 9 2 10 0 11 1 11 7 11 1 11 13 10 9 1 15 13 1 13 15 2 1 9 1 13 1 10 9 3 0 7 10 11 16 13 10 9 0 2
53 10 9 0 2 3 13 1 9 0 2 13 3 1 13 10 9 13 15 7 13 9 3 2 13 10 9 0 7 13 10 0 9 1 9 1 10 9 2 10 9 2 10 9 2 10 9 7 10 9 2 1 15 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
25 1 13 1 10 9 4 13 9 0 1 10 9 2 7 10 0 9 13 13 1 10 9 1 9 2
9 13 10 9 1 10 9 1 3 2
21 3 13 10 9 1 10 11 11 2 1 15 15 15 13 1 10 9 1 10 9 2
42 1 10 11 1 10 11 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
96 1 10 9 0 7 9 0 1 11 11 11 2 11 11 2 2 10 9 1 10 9 1 9 16 11 11 11 15 4 13 1 12 13 16 13 1 10 0 9 1 13 10 9 1 9 13 1 10 9 1 9 2 15 16 13 10 9 1 10 9 2 13 1 10 9 0 7 0 2 1 10 9 1 10 16 13 2 1 10 9 0 1 10 9 0 1 9 1 13 10 9 1 10 9 2 2
44 13 3 10 9 1 9 1 0 9 2 1 10 16 13 1 10 9 12 1 4 4 13 1 10 11 1 11 1 10 11 1 12 9 1 9 2 10 12 5 1 10 9 2 2
13 3 13 1 9 7 1 9 1 9 13 10 9 2
8 1 9 3 13 10 0 9 2
48 10 9 8 15 13 1 11 1 10 9 0 1 11 7 15 13 1 10 0 9 1 10 9 12 13 1 10 0 9 0 8 10 9 16 13 1 13 15 1 10 9 0 7 1 9 1 13 2
41 1 1 10 9 1 12 10 9 16 15 13 0 1 13 10 9 13 1 10 9 1 11 2 15 16 13 1 10 11 10 9 15 0 1 10 9 1 9 1 9 2
60 1 10 9 1 10 9 1 10 9 15 13 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 7 11 11 2
20 11 11 13 10 9 1 9 1 10 9 1 10 11 1 10 9 1 10 11 2
12 10 9 1 9 1 10 9 13 1 5 12 2
21 1 11 1 12 13 9 1 10 11 11 16 13 10 9 1 10 9 0 1 11 2
20 3 13 10 9 2 2 1 10 9 16 13 9 15 4 13 16 13 0 2 2
20 1 9 16 13 15 13 10 9 1 10 9 2 9 7 0 9 1 10 9 2
23 9 1 11 11 2 11 2 11 11 2 11 11 8 4 13 10 9 1 10 9 1 11 2
10 10 9 0 1 9 13 10 12 8 2
17 11 11 8 11 11 2 8 12 2 13 10 9 2 7 9 0 2
52 11 11 13 1 10 9 11 11 1 11 1 10 11 3 15 13 10 9 1 10 16 13 10 9 1 9 1 11 11 2 15 1 10 0 9 2 10 15 13 3 10 12 1 11 1 12 1 10 9 1 9 2
23 10 11 13 1 10 11 11 2 1 9 1 11 11 2 10 15 13 9 1 10 9 11 2
28 3 4 13 9 0 2 7 15 16 13 1 11 11 1 2 10 3 0 9 1 9 0 1 10 0 9 2 2
12 11 11 13 10 9 1 9 1 10 9 11 2
23 10 9 13 1 10 9 1 9 16 15 13 2 7 13 1 11 2 16 15 13 3 0 2
42 10 9 16 13 10 9 12 1 10 9 11 1 12 9 7 12 1 10 9 11 9 1 11 11 2 11 11 7 11 11 11 16 3 13 10 0 9 1 10 9 0 2
24 15 13 1 10 9 13 1 9 1 10 9 7 15 13 1 10 9 16 15 15 13 1 0 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
14 13 10 9 16 13 10 0 9 1 11 2 11 11 2
18 16 13 10 9 13 10 9 2 3 4 13 10 9 0 1 10 9 2
12 2 15 13 1 9 15 16 13 1 10 9 2
26 10 9 0 13 10 9 1 9 0 13 1 10 9 1 10 9 1 10 11 11 1 10 9 12 8 2
16 10 9 1 10 9 12 13 12 9 1 9 7 10 3 9 2
34 11 11 15 13 16 3 13 0 1 13 15 2 7 13 9 1 9 1 10 9 13 1 10 9 1 9 2 15 13 13 13 10 9 2
24 10 9 13 1 10 9 0 7 1 10 9 1 9 1 10 9 0 10 9 0 1 10 9 2
83 10 11 1 11 15 13 10 12 1 11 1 12 2 3 1 10 2 11 1 11 2 12 2 1 12 9 1 9 1 10 9 13 1 11 11 7 10 9 0 1 11 12 1 10 11 11 11 11 2 1 3 1 12 9 1 10 9 1 0 9 1 11 11 2 11 11 7 11 11 10 15 1 10 9 1 11 1 11 2 11 1 11 2
45 3 2 16 10 9 13 10 9 2 13 1 13 1 9 1 0 9 2 4 10 9 1 10 9 1 11 11 1 13 10 9 3 15 4 13 10 9 1 9 16 4 1 13 15 2
18 13 1 9 1 10 9 1 10 8 1 10 9 1 12 1 11 11 2
39 13 1 13 1 12 9 3 1 10 9 2 7 13 10 12 9 1 9 1 9 2 7 3 13 9 1 16 10 9 4 13 1 10 11 11 11 1 12 2
26 1 10 9 4 13 1 10 11 11 2 1 3 13 1 8 3 15 13 13 1 11 11 1 11 11 2
9 13 1 11 1 11 2 11 2 2
31 10 9 13 1 9 1 10 9 11 11 7 13 13 10 9 1 10 9 1 10 8 9 2 13 10 12 1 11 1 12 2
24 13 10 12 1 11 1 12 2 10 15 3 13 10 9 1 10 11 1 10 11 1 11 11 2
17 3 1 13 2 10 9 13 10 9 2 7 13 1 13 1 11 2
20 13 1 10 9 11 11 2 1 10 9 2 13 1 10 9 12 7 3 13 2
43 13 1 10 9 16 15 13 3 3 2 13 15 1 10 9 3 0 7 4 13 1 11 1 12 16 13 10 0 9 2 16 4 13 1 10 11 11 7 1 10 11 11 2
7 4 13 1 10 9 11 2
25 1 10 9 0 15 13 10 9 1 10 9 1 10 9 1 10 9 0 1 9 7 1 0 9 2
16 1 10 9 13 12 9 7 15 13 9 1 10 11 11 0 2
27 1 9 1 15 16 13 1 10 9 1 9 2 10 9 1 10 9 1 9 13 1 10 9 1 10 9 2
45 3 1 10 9 1 10 11 10 11 2 3 13 1 10 11 2 13 10 9 8 1 10 9 2 7 4 13 3 12 9 2 10 10 11 13 3 1 10 11 11 1 10 11 11 2
16 15 13 13 1 10 9 1 10 9 1 10 9 10 10 9 2
30 10 9 13 0 2 1 10 9 7 10 9 13 7 13 3 0 1 10 9 7 1 10 9 1 12 7 12 9 2 2
16 10 11 13 9 1 11 2 11 1 11 2 7 1 11 11 2
20 11 13 10 9 0 1 10 9 16 13 11 7 11 1 10 9 1 11 11 2
30 10 9 1 11 15 13 0 1 10 9 1 10 9 1 11 2 3 1 12 9 1 10 9 1 10 9 1 10 9 2
34 1 3 10 9 0 13 10 12 9 0 2 10 9 15 0 13 1 9 3 10 0 9 16 4 13 16 13 10 9 1 10 0 9 2
34 1 10 9 0 1 11 11 15 1 10 0 9 1 10 11 11 2 10 9 1 10 11 11 13 15 3 0 7 15 1 10 10 9 2
12 3 10 9 12 7 12 13 1 10 0 9 2
33 1 15 10 9 15 13 1 10 9 0 1 10 9 11 2 1 11 2 11 7 11 1 10 9 12 2 13 1 12 9 1 0 2
30 10 9 15 4 13 1 10 3 13 2 3 16 13 10 0 11 11 2 9 0 1 10 9 2 2 13 1 9 0 2
34 10 9 3 15 13 1 3 0 9 1 10 9 2 3 1 9 3 13 3 7 9 1 10 9 2 3 13 1 9 1 10 9 12 2
14 3 13 10 9 0 1 10 15 10 9 13 3 0 2
16 9 11 11 11 11 13 10 9 0 16 13 1 10 11 11 2
22 10 9 7 10 9 1 10 9 1 9 15 13 1 10 11 7 11 1 11 1 11 2
12 1 10 9 7 9 0 1 11 15 4 13 2
20 9 0 1 10 9 0 2 12 11 2 2 13 1 10 0 11 11 1 12 2
52 1 10 9 1 0 9 2 11 13 1 11 11 2 15 3 13 9 1 10 9 1 10 11 11 2 2 1 13 1 10 9 16 13 1 10 9 2 15 15 13 1 10 9 1 13 1 10 9 1 10 9 2
24 10 9 0 1 11 13 10 13 10 9 0 2 13 1 9 2 9 1 9 7 9 1 9 2
55 10 9 1 10 9 1 9 1 10 9 7 10 4 13 13 10 9 0 1 10 9 2 10 0 9 0 13 2 3 1 10 9 2 0 1 10 9 1 10 9 16 15 13 2 13 10 9 2 12 2 2 3 3 2 2
34 16 13 3 3 10 9 0 2 10 9 0 1 10 9 9 7 1 10 9 0 1 9 13 0 2 1 9 0 3 1 9 1 9 2
54 10 9 11 11 2 1 9 2 2 9 1 9 1 10 9 2 7 1 9 2 9 9 2 2 13 10 9 0 3 0 15 4 4 13 1 11 7 11 1 10 9 1 10 11 1 11 2 1 10 9 9 1 11 2
33 10 9 1 10 9 1 9 1 10 9 13 10 11 1 10 11 1 10 11 11 11 2 16 13 10 0 9 1 10 9 1 11 2
38 10 9 0 4 13 3 16 15 4 13 9 1 9 1 9 0 2 7 15 4 4 13 1 9 1 9 2 3 16 15 3 13 0 1 13 10 9 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
9 3 3 13 15 16 3 13 15 2
13 15 1 10 9 15 13 3 3 1 10 0 9 2
46 13 1 11 11 1 12 1 9 1 10 9 11 1 10 11 1 12 9 1 9 0 7 10 0 9 1 9 0 2 9 1 10 15 13 4 13 13 16 10 9 13 0 1 10 9 2
35 10 9 1 10 9 1 9 0 2 11 11 4 13 1 10 9 1 13 10 0 9 13 10 9 16 13 7 10 9 15 13 1 12 9 2
39 11 13 16 10 9 0 13 2 1 10 9 1 10 9 1 9 2 2 15 16 2 3 13 3 10 9 0 1 10 9 1 10 16 15 13 10 9 2 2
17 1 10 9 0 13 11 11 2 9 2 7 11 11 2 9 2 2
32 1 10 9 2 13 1 10 9 1 10 9 1 16 13 1 10 9 1 13 9 16 13 1 13 10 9 0 2 0 7 0 2
25 13 1 15 16 2 3 16 10 9 4 13 11 11 2 10 15 1 10 12 9 13 10 9 0 2
33 1 9 1 9 13 1 9 1 11 2 8 8 2 11 2 16 13 10 11 1 11 2 13 1 10 0 9 1 10 9 1 9 2
29 3 2 13 10 9 1 9 7 9 11 2 10 9 13 10 3 9 2 11 11 2 2 1 3 3 1 10 9 2
29 1 15 2 1 9 0 7 3 2 10 9 4 13 10 0 9 1 10 9 1 16 15 13 10 9 1 10 15 2
32 3 3 1 13 10 9 1 10 9 1 11 2 15 15 13 1 10 9 7 3 15 13 3 16 15 13 10 9 1 10 9 2
28 1 3 13 9 1 10 9 1 10 11 11 7 15 13 1 9 1 10 9 7 1 10 9 0 1 9 0 2
39 1 10 9 11 10 11 4 7 13 10 9 7 10 9 16 13 0 2 10 9 1 9 13 13 16 10 9 13 3 0 1 9 7 10 9 3 13 0 2
65 10 9 1 10 11 11 13 0 2 15 1 15 1 9 13 15 1 10 9 1 11 1 9 1 10 9 1 10 9 1 12 9 1 9 16 13 15 16 13 1 10 9 3 2 10 9 16 3 13 1 10 9 2 3 1 11 2 9 1 10 11 1 11 3 2
13 11 11 11 13 10 0 9 1 11 2 11 11 2
22 10 9 13 15 13 10 9 16 15 13 1 12 9 1 16 3 13 10 12 5 0 2
37 11 11 2 0 2 11 2 13 10 9 1 10 9 1 9 1 9 0 13 1 11 11 11 2 1 9 0 1 11 11 2 7 13 1 11 11 2
32 9 4 13 16 1 10 9 7 9 1 9 1 10 9 4 9 1 10 9 1 3 12 9 1 10 15 12 13 0 1 9 2
24 10 9 2 10 9 1 10 9 11 2 11 2 0 2 11 7 11 2 13 13 1 10 9 2
22 10 0 9 15 13 1 15 9 1 10 12 9 1 9 2 1 10 9 1 0 9 2
21 15 13 16 15 13 10 9 7 2 3 15 13 1 11 16 3 13 16 13 0 2
27 10 11 11 4 13 1 10 9 1 11 10 11 2 9 0 16 13 1 11 11 7 16 13 1 10 11 2
12 1 13 12 9 13 10 9 1 10 9 11 2
19 10 9 15 4 13 1 10 9 0 2 13 1 10 0 9 1 10 9 2
42 1 10 9 0 2 10 9 1 12 9 4 4 13 1 9 0 2 7 7 2 10 9 3 0 2 2 7 3 10 9 0 7 0 15 4 13 1 9 1 9 0 2
8 9 13 10 12 1 11 1 12
28 3 3 13 0 15 13 10 9 1 9 1 13 0 9 0 2 0 1 10 0 9 1 10 11 1 10 11 2
52 10 9 0 1 9 1 10 8 13 10 9 0 1 10 9 1 9 1 10 9 2 1 10 9 2 1 10 0 9 15 13 10 9 2 3 15 2 13 2 10 9 2 15 13 2 7 3 15 13 1 9 2
30 1 9 2 16 13 12 2 4 1 13 2 16 13 12 10 9 13 12 2 12 1 10 0 7 12 1 10 9 2 2
26 10 9 1 9 1 10 0 9 1 10 9 1 11 11 3 15 13 1 10 9 0 0 1 10 9 2
30 11 11 2 11 2 12 1 11 1 12 2 13 10 9 1 9 1 11 16 13 1 10 11 1 11 11 11 1 11 2
30 3 1 10 9 16 13 10 9 7 12 2 11 1 11 13 1 10 11 11 1 10 0 9 7 15 13 1 10 9 2
15 15 15 13 0 9 2 3 9 1 10 9 7 0 9 2
42 10 9 0 2 15 13 10 9 1 9 0 16 13 1 13 1 10 9 1 11 7 11 2 15 13 10 11 1 11 1 10 9 0 11 11 7 13 10 9 1 11 2
16 15 13 1 10 9 0 16 13 10 9 7 10 9 1 9 2
26 10 9 4 13 10 9 3 13 10 0 9 1 10 9 1 3 1 12 9 7 13 13 15 13 3 2
24 11 11 2 11 11 2 11 0 2 12 1 11 1 12 2 13 10 9 2 9 7 9 0 2
13 3 0 13 1 10 9 16 1 15 15 13 11 2
57 16 10 9 3 3 13 1 0 9 2 10 9 15 13 1 9 0 7 3 2 10 9 1 10 12 9 4 13 1 13 1 10 15 1 10 9 1 10 9 0 2 9 2 9 2 9 2 2 8 2 8 2 8 1 11 2 2
29 13 0 10 9 0 15 13 11 7 3 16 10 9 15 13 1 10 9 16 13 15 9 1 9 15 11 4 13 2
12 2 4 13 15 3 10 9 1 10 9 0 2
16 3 4 13 1 12 9 0 13 1 12 7 12 9 1 15 2
36 13 10 9 0 9 16 13 3 1 12 9 2 13 3 1 10 11 11 11 11 1 11 2 1 9 1 10 15 13 10 10 9 0 7 0 2
26 11 13 0 1 10 9 16 10 9 4 13 1 10 9 2 7 11 15 13 16 10 9 13 10 9 2
16 16 4 7 13 12 9 1 16 13 10 9 1 11 1 12 2
23 1 9 2 12 9 16 15 13 1 10 9 15 13 1 10 9 16 13 15 2 3 13 2
19 10 9 11 11 13 10 0 8 1 10 9 1 10 9 0 16 3 13 2
15 3 15 13 3 1 10 9 0 7 3 0 7 1 9 2
33 1 9 1 10 9 0 16 13 10 9 2 13 13 15 1 10 9 7 1 10 9 13 2 7 13 13 15 1 10 9 1 9 2
21 10 9 13 13 1 10 9 11 2 11 2 13 1 10 9 11 11 11 2 11 2
32 15 13 10 9 9 12 1 10 9 2 15 4 13 10 12 1 11 1 12 2 1 11 7 11 3 3 4 4 13 10 9 2
20 3 15 13 10 9 3 0 16 13 1 10 9 2 1 10 12 5 1 9 2
21 11 11 2 8 12 1 11 1 12 2 11 2 11 2 11 2 13 10 9 0 2
42 10 11 1 11 1 15 11 2 10 11 0 1 10 11 11 2 10 0 11 11 2 10 9 1 9 11 2 9 13 1 13 10 9 1 9 2 7 10 9 1 9 2
18 11 11 13 10 9 16 13 1 11 11 2 11 11 2 7 11 11 2
44 13 16 10 9 0 2 13 10 0 9 2 13 3 1 10 0 9 2 13 1 10 9 0 7 13 3 10 9 1 10 15 15 13 2 3 16 15 13 1 15 10 9 0 2
19 13 10 0 9 16 15 13 1 10 9 1 9 7 10 9 0 1 13 2
11 1 11 1 12 11 13 10 9 1 11 2
27 11 11 2 11 13 10 11 12 1 11 1 10 12 9 16 13 1 10 9 0 2 1 10 9 0 0 2
24 16 3 13 10 9 2 11 13 15 16 13 2 7 3 15 13 2 2 10 9 0 13 0 2
38 11 13 1 13 15 1 10 0 9 1 11 11 11 1 11 1 12 2 3 7 11 11 15 13 1 13 1 9 1 10 9 1 8 8 8 8 8 2
22 1 9 13 10 9 2 1 11 11 2 13 2 11 2 2 16 13 9 1 10 11 2
16 13 10 9 1 10 11 11 2 16 13 1 10 0 11 0 2
46 10 9 1 10 11 11 11 1 11 15 4 13 1 9 2 9 1 10 9 0 2 9 2 9 2 9 1 10 0 8 7 9 1 10 9 16 13 1 10 9 1 9 2 11 11 2
35 10 11 15 13 10 9 7 1 9 1 9 2 1 10 9 2 15 13 9 1 10 9 1 10 9 7 10 9 1 16 13 1 10 9 2
22 10 9 13 1 10 9 13 1 10 9 1 11 1 10 12 9 1 10 9 1 3 2
11 3 7 13 10 9 7 15 13 3 3 2
22 4 7 13 10 10 9 1 9 4 13 2 15 15 13 2 15 13 10 9 0 2 2
16 13 1 10 9 1 9 1 12 2 1 10 9 1 12 9 2
58 9 2 3 13 1 13 10 9 7 3 13 2 4 7 13 9 2 3 13 13 1 10 9 2 16 13 13 10 9 0 2 13 15 15 1 10 9 2 13 15 10 9 2 16 13 15 16 13 2 7 16 13 10 9 10 16 13 2
73 11 15 13 2 1 9 2 16 11 7 11 15 13 2 13 16 10 9 1 11 13 10 0 9 1 9 3 13 10 9 0 13 1 10 9 2 16 11 7 11 2 8 2 7 11 7 11 2 8 2 13 10 9 0 1 15 2 15 15 15 13 15 7 13 10 9 1 11 1 13 1 11 2
24 10 0 9 1 10 9 13 1 10 9 1 11 11 1 10 9 1 11 2 13 1 10 11 2
35 11 11 15 13 10 0 9 1 9 0 1 10 0 9 1 10 9 2 3 4 13 10 9 0 7 10 9 1 10 9 1 9 1 11 2
16 1 9 4 1 13 16 3 15 13 16 10 9 3 13 0 2
32 10 9 0 1 10 0 9 2 11 11 2 15 13 1 11 11 2 13 1 10 9 0 2 1 10 9 13 1 10 9 11 2
38 16 13 10 9 1 9 1 15 7 10 9 2 1 10 9 1 10 9 2 10 9 1 9 1 10 9 15 13 1 10 9 1 9 3 1 10 12 2
21 3 15 13 2 13 15 16 4 7 13 7 13 3 2 1 10 9 13 10 9 2
14 10 0 9 13 1 11 11 11 12 1 10 9 12 2
16 11 11 13 10 9 0 2 13 3 1 11 2 11 0 2 2
15 1 10 9 1 10 9 2 11 13 12 9 0 1 9 2
10 1 12 13 10 9 1 12 12 9 2
34 13 0 9 2 10 9 7 10 15 13 0 2 15 7 15 16 4 13 1 11 1 10 3 0 8 15 0 16 4 13 1 10 9 2
16 11 11 13 10 9 1 9 1 10 9 11 1 10 9 11 2
43 10 11 2 10 9 1 10 9 11 7 11 2 4 13 1 12 2 1 9 1 10 9 1 9 7 1 9 1 13 10 9 1 9 1 11 11 1 11 8 1 10 9 2
32 11 11 11 2 8 12 1 11 1 12 2 13 10 9 0 2 13 3 1 10 9 1 11 11 1 11 7 11 11 1 11 2
13 11 13 1 11 11 1 10 9 1 12 0 9 2
21 1 10 0 9 13 10 9 0 2 10 9 1 10 9 7 10 1 10 9 0 2
16 1 13 10 9 0 1 10 9 13 1 9 1 9 7 9 2
22 3 13 16 13 9 2 7 1 10 9 2 3 13 16 13 1 10 9 1 10 9 2
13 10 9 13 1 9 3 16 10 9 4 13 0 2
13 13 9 1 11 11 1 12 9 1 12 7 12 2
27 3 4 7 13 10 0 9 1 10 9 1 10 0 9 2 10 9 1 11 7 10 9 1 11 2 11 2
24 10 9 13 1 10 9 0 1 10 9 1 10 11 2 16 13 10 9 1 10 9 1 11 2
62 10 9 4 13 1 10 9 2 3 3 4 13 10 9 13 1 11 16 13 10 9 1 10 9 1 10 9 1 10 9 1 12 9 7 10 9 13 1 9 1 10 9 1 11 11 2 9 0 2 7 11 11 2 15 4 13 10 9 1 0 9 2
14 1 10 11 0 10 9 15 13 1 9 1 9 0 2
58 10 9 1 11 13 10 9 0 2 13 13 1 9 0 2 16 4 13 10 9 1 10 9 1 10 9 1 11 2 10 9 1 12 9 1 9 7 10 9 0 1 12 8 2 10 15 15 4 13 3 1 10 0 12 9 1 9 2
16 10 0 9 2 11 11 11 2 13 10 9 0 9 1 11 2
13 13 9 1 9 0 9 16 13 1 10 0 9 2
35 3 1 13 15 7 1 0 9 2 10 12 1 11 15 13 10 9 0 1 11 2 15 1 15 15 3 15 13 9 2 13 10 9 0 2
8 15 4 13 1 13 1 13 2
28 11 1 11 2 10 0 9 0 1 10 9 2 7 1 10 9 2 13 9 1 10 0 9 0 1 10 9 2
32 11 11 1 11 11 2 12 2 9 2 9 0 0 9 1 10 9 7 9 0 2 13 0 1 11 11 12 1 10 9 12 2
15 10 0 9 15 13 10 9 12 2 13 1 9 1 9 2
22 10 9 4 13 3 1 11 1 11 16 15 13 1 10 9 0 16 13 3 1 9 2
19 10 9 11 13 9 1 10 9 1 10 9 16 15 13 1 9 1 9 2
19 15 13 1 10 9 0 7 1 9 16 15 13 1 10 9 1 10 9 2
11 4 13 9 7 13 0 9 1 9 0 2
19 15 13 1 1 10 9 13 11 2 7 10 9 13 0 1 13 10 9 2
47 10 9 13 1 10 9 2 13 9 7 9 0 2 10 9 15 13 11 2 11 13 9 1 10 9 0 8 2 0 2 2 13 0 1 9 2 7 13 10 9 1 10 0 9 1 9 2
30 1 10 0 9 1 10 9 10 9 3 1 10 9 1 10 9 13 1 10 0 7 0 9 4 4 13 10 9 0 2
12 10 9 1 9 13 1 12 8 2 5 12 2
8 3 4 13 11 11 7 11 2
12 10 9 13 0 1 10 9 2 1 3 0 2
15 10 9 13 10 9 1 9 1 10 9 1 11 11 11 2
12 1 10 9 15 13 0 9 1 10 10 9 2
29 10 1 11 13 13 1 11 1 11 7 1 10 3 13 4 1 13 15 1 11 2 13 10 9 3 1 10 9 2
13 2 9 1 9 1 10 9 16 13 3 9 1 9
46 1 11 1 10 0 9 2 10 9 1 11 11 7 11 11 11 15 13 1 10 11 11 2 10 9 0 13 1 10 9 0 11 7 11 11 2 2 16 13 10 12 5 1 10 9 2
33 10 9 0 13 0 0 3 1 10 0 9 2 1 15 15 3 13 9 1 16 13 1 15 1 10 9 3 0 13 1 10 9 2
29 7 2 1 9 1 15 2 1 10 9 1 12 1 12 1 9 1 11 12 2 10 9 13 13 15 1 10 9 2
30 3 2 10 9 0 2 0 2 3 4 3 13 1 9 2 1 15 15 3 15 13 9 0 7 15 13 3 11 11 2
33 16 3 13 12 9 7 13 1 10 11 11 1 11 4 13 1 10 9 1 10 11 11 1 11 2 13 1 10 9 1 9 0 2
38 1 11 1 12 7 1 0 9 0 1 11 11 11 13 10 9 7 4 13 11 1 10 11 11 7 2 7 0 2 9 1 10 11 1 11 1 11 2
23 11 13 1 10 9 1 11 1 12 1 10 11 11 11 11 11 11 2 1 10 9 11 2
32 15 1 10 9 0 1 10 9 13 10 1 11 11 1 10 9 1 10 9 1 9 1 10 11 2 9 2 10 9 1 11 2
17 15 13 1 10 9 1 11 13 10 9 2 7 13 3 1 9 2
36 3 3 13 10 9 0 1 10 9 0 2 0 2 3 13 1 9 1 11 16 13 1 10 11 11 2 3 10 9 13 10 11 1 10 11 2
26 10 9 9 1 10 11 11 15 13 13 10 9 1 12 9 3 2 12 13 2 12 13 1 9 12 2
12 10 9 13 10 9 1 13 15 1 10 9 2
31 10 9 13 0 1 10 12 1 11 1 12 2 1 9 1 10 0 9 2 1 10 9 2 1 10 12 1 11 1 12 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
28 1 11 1 12 2 10 0 11 11 4 13 10 9 1 9 0 1 10 9 1 11 7 11 13 9 1 9 2
15 11 11 2 12 2 12 2 2 9 2 9 7 9 0 2
14 4 13 0 1 10 9 1 9 1 11 1 12 9 2
30 10 9 8 13 9 16 13 10 9 0 1 10 9 0 1 10 9 0 2 13 15 1 10 0 9 13 9 1 9 2
25 10 9 1 11 13 1 10 9 1 10 9 10 9 0 2 7 3 10 9 0 1 10 9 0 2
31 10 9 1 11 11 11 2 1 11 2 3 4 4 13 1 10 9 1 9 3 1 10 9 16 15 13 10 12 1 11 2
21 13 15 15 15 13 2 13 3 2 13 15 1 9 1 10 9 15 15 4 13 2
44 10 9 13 10 5 9 0 13 12 9 7 13 0 1 10 9 2 15 15 13 16 15 3 13 10 9 3 7 10 9 1 9 16 15 13 16 13 1 10 9 1 10 9 2
27 10 9 7 9 1 11 11 0 15 13 0 7 15 13 1 10 9 1 11 1 10 9 1 11 1 9 2
50 0 1 10 9 2 10 9 13 10 9 1 9 7 9 1 12 9 2 1 15 2 11 15 13 1 10 0 9 1 10 9 1 10 9 1 10 9 1 13 9 2 7 10 8 8 1 10 12 9 2
28 1 13 9 11 1 11 2 9 1 10 9 2 10 9 1 11 11 7 10 9 2 3 15 13 1 10 9 2
27 10 9 0 1 11 13 10 9 1 9 0 2 0 2 9 7 9 7 9 2 2 0 0 7 9 0 2
9 13 9 1 13 1 13 10 9 2
17 11 13 1 11 1 12 9 2 7 3 13 10 9 1 10 9 2
43 1 10 9 12 2 10 9 15 13 1 9 1 10 9 2 7 12 9 3 2 1 12 2 10 9 0 11 15 13 9 1 10 9 2 16 13 10 9 0 1 11 11 8
27 1 12 2 10 0 9 13 10 9 1 9 0 2 15 16 13 1 10 9 1 10 9 1 10 11 11 2
22 10 9 1 10 9 0 2 7 10 9 0 1 10 9 2 13 9 1 10 9 0 2
18 10 0 9 1 10 2 9 2 13 1 10 9 1 11 7 1 11 2
42 1 13 2 13 1 10 9 11 11 13 15 10 12 9 1 10 9 3 13 16 10 9 13 3 0 2 3 16 3 13 3 16 0 1 13 10 9 1 10 9 2 2
25 10 9 1 11 11 2 0 9 1 9 1 11 2 13 15 1 10 9 0 3 0 1 10 9 2
37 11 10 9 0 2 2 13 1 11 1 10 12 9 1 13 10 11 1 10 11 7 13 1 10 0 11 1 11 2 9 1 10 9 1 10 9 2
46 1 10 9 1 10 9 1 10 9 1 9 1 10 9 2 10 15 16 4 13 1 10 11 13 1 0 9 2 1 9 1 16 13 1 9 7 13 10 9 1 13 10 9 1 9 2
38 15 1 10 9 3 0 13 15 1 11 11 2 16 13 10 9 0 2 3 7 10 0 9 2 11 0 2 2 1 10 9 11 11 2 1 12 9 2
20 10 9 0 15 4 13 1 15 9 1 10 9 1 9 1 10 12 0 9 0
15 3 4 13 3 10 9 7 10 9 0 7 3 4 13 2
36 11 2 7 2 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2 1 2 11 2
23 13 0 1 10 12 1 11 1 12 2 16 4 13 1 10 0 11 11 1 11 1 12 2
37 2 10 9 13 1 10 9 1 11 13 2 10 9 0 2 13 15 1 10 9 0 0 2 3 9 13 1 9 0 13 1 9 1 9 7 9 2
110 1 10 9 15 13 10 9 1 10 9 2 1 10 9 0 2 15 9 1 10 13 10 9 0 1 12 1 10 9 1 9 1 9 2 3 7 10 9 9 0 2 10 9 0 2 7 10 9 1 10 9 0 2 0 7 13 10 9 0 1 10 0 9 0 2 10 9 13 1 10 9 1 10 9 1 10 9 1 9 0 2 0 7 13 10 9 1 11 11 2 10 9 1 10 9 13 13 1 10 9 2 7 10 9 4 13 1 10 9 2
43 3 1 10 9 1 10 11 11 2 10 9 1 11 13 10 9 1 11 1 7 10 9 13 10 9 0 16 3 4 1 13 15 2 7 1 10 16 11 15 13 12 9 2
27 11 11 13 10 9 0 0 2 13 1 12 2 16 13 10 9 7 13 9 1 9 0 7 1 9 0 2
28 10 0 9 2 11 11 11 11 2 15 13 1 10 0 9 7 13 9 1 10 9 9 0 2 13 1 12 2
53 10 9 0 4 13 10 9 13 10 9 1 9 7 1 9 0 1 10 9 7 13 1 9 2 10 9 0 13 1 10 9 1 10 9 1 10 9 7 10 9 13 16 4 13 13 15 10 9 1 10 9 2 2
40 1 10 9 13 3 16 13 1 10 9 11 11 2 1 10 9 11 2 11 2 11 7 11 2 1 10 0 9 16 15 4 13 1 10 9 1 10 9 0 2
41 1 15 9 2 13 0 13 16 10 9 4 13 10 9 0 7 4 13 1 9 1 13 1 15 3 9 1 10 9 1 10 9 7 13 15 1 9 1 10 9 2
8 13 1 10 9 1 12 9 2
18 4 13 1 11 1 12 2 7 3 4 1 13 9 1 10 0 9 2
13 10 0 9 16 13 10 9 0 13 1 10 9 2
22 11 12 13 3 1 9 10 9 1 10 9 11 7 11 2 3 1 10 9 11 5 2
21 15 15 15 13 1 10 9 0 2 3 15 13 7 9 1 9 7 9 7 15 2
11 13 3 1 11 2 9 0 1 10 9 2
29 1 10 9 12 10 9 2 11 11 2 13 10 9 1 2 11 11 2 11 2 2 13 1 10 9 1 11 11 2
34 13 3 0 13 1 10 9 16 4 13 10 9 0 1 10 0 9 2 13 10 9 1 11 7 1 1 11 1 11 7 11 2 3 2
12 11 11 13 10 9 1 9 1 10 9 11 2
33 1 10 9 1 12 2 12 5 1 11 13 0 2 3 16 10 9 0 2 12 5 2 7 3 16 10 9 0 2 12 5 2 2
10 15 13 10 2 8 2 1 10 9 2
72 10 9 4 13 1 10 9 2 13 9 15 10 9 0 2 16 15 15 4 13 1 9 1 9 0 1 10 9 1 11 2 1 9 1 10 9 13 1 10 9 1 12 1 10 9 0 7 0 2 10 15 13 9 1 9 1 0 9 16 13 16 1 10 0 9 1 11 15 13 9 0 2
20 15 13 1 0 9 10 9 7 13 10 9 1 10 9 1 9 1 10 9 2
17 1 15 10 9 1 9 13 1 2 9 0 2 16 3 15 13 2
19 4 13 1 10 11 1 10 11 11 7 13 0 1 10 11 11 1 11 2
14 15 13 7 15 13 8 9 1 13 10 9 1 9 2
42 1 0 2 10 0 9 13 10 9 3 8 1 11 2 9 1 9 7 9 2 9 1 9 2 9 1 10 9 2 9 1 9 2 10 9 1 10 9 1 4 13 2
48 10 9 13 16 11 2 16 3 13 10 9 3 0 1 10 9 2 13 12 9 1 9 1 13 1 11 11 1 10 0 12 9 1 10 9 2 12 9 1 10 15 2 2 13 1 11 11 2
24 11 13 10 9 1 9 1 10 9 7 9 0 11 11 13 1 11 1 12 1 9 1 11 2
31 10 9 1 11 11 11 2 8 11 11 2 10 12 5 11 1 10 9 2 4 13 1 10 11 11 1 11 2 1 11 2
45 3 0 2 10 9 3 2 1 12 10 9 1 9 0 1 10 9 8 1 10 9 11 11 2 9 1 10 9 11 11 7 11 11 2 4 13 1 10 11 11 1 11 11 11 2
15 1 10 9 15 13 10 9 0 1 10 9 1 12 9 2
35 13 13 15 1 10 9 0 16 15 13 3 3 1 10 9 1 10 9 2 3 1 9 0 2 1 10 9 1 10 15 10 9 13 0 2
13 10 9 1 9 1 11 13 0 7 1 0 9 2
22 10 9 4 13 13 1 10 9 1 10 9 0 0 1 9 1 13 9 0 1 11 2
21 10 9 1 9 11 4 13 3 1 11 2 12 2 1 10 0 9 1 11 11 2
39 1 9 4 13 16 13 10 9 2 7 3 15 1 10 9 3 0 2 2 16 4 13 1 10 9 1 9 2 4 13 1 10 9 1 10 10 9 2 2
28 10 9 4 13 1 10 9 12 1 11 11 2 1 10 9 11 11 1 2 11 2 9 1 11 11 1 11 2
21 1 15 2 10 9 1 9 0 15 13 1 9 7 4 13 3 16 15 13 0 2
9 9 1 10 11 11 1 11 1 12
23 13 2 3 2 9 13 10 0 9 0 2 1 9 1 10 9 1 10 9 11 1 11 2
20 1 10 9 2 13 1 11 11 1 12 9 2 13 12 9 7 12 13 0 2
21 13 15 9 7 9 0 2 1 10 10 9 4 13 15 9 1 10 9 1 9 2
48 1 10 9 1 11 13 10 9 0 1 9 0 1 10 9 1 10 9 0 2 13 10 11 1 11 11 1 12 2 1 9 1 11 11 13 1 11 11 2 11 11 7 11 11 2 1 15 2
29 10 11 7 9 3 13 1 10 0 9 0 2 16 1 15 1 15 10 9 1 9 0 4 13 10 9 0 0 2
15 10 9 11 12 1 11 3 15 4 13 1 11 1 12 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
81 10 9 13 2 1 9 3 13 1 10 9 1 9 2 9 2 9 1 11 11 2 2 13 10 9 13 1 9 7 9 1 10 9 1 9 13 16 13 3 0 7 2 12 2 13 9 1 9 0 16 13 13 3 1 10 9 1 10 0 9 1 10 9 7 2 12 2 13 10 9 1 9 1 9 2 1 9 0 7 0 2
59 1 10 12 9 2 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
46 11 13 10 0 9 1 10 9 1 10 11 11 1 10 9 9 10 12 2 15 13 13 1 10 9 1 10 9 2 1 10 15 10 9 13 13 15 1 9 1 10 9 1 11 11 2
20 1 4 13 1 11 1 15 2 11 13 16 13 1 9 1 10 9 1 9 2
26 11 11 11 2 11 2 12 1 11 1 12 2 13 10 9 2 9 2 9 2 9 0 7 9 0 2
36 1 9 2 1 0 9 2 11 4 1 13 10 0 9 13 10 10 9 0 1 10 10 8 8 7 9 1 10 9 3 7 10 9 0 0 2
44 10 9 1 11 2 11 11 7 11 13 0 7 13 3 3 1 10 9 1 10 9 7 3 1 10 9 1 13 1 10 9 0 7 13 10 0 9 1 10 9 1 10 11 2
34 11 13 16 10 9 0 1 11 13 1 10 9 1 10 11 13 3 0 9 1 10 13 1 10 9 1 11 10 12 1 11 1 12 2
18 1 12 4 13 1 10 9 0 11 7 11 11 1 10 9 1 9 2
12 10 9 1 9 13 10 9 0 1 11 11 2
47 1 10 9 0 2 13 3 1 9 1 10 9 0 7 13 1 15 2 15 13 12 9 1 9 2 13 1 9 2 3 13 2 13 1 10 9 0 2 1 10 9 1 9 1 10 9 2
25 13 0 1 10 9 0 2 10 9 0 2 10 9 2 7 10 9 7 10 9 1 9 1 9 2
20 15 13 1 10 9 1 11 11 7 11 11 2 1 12 7 12 9 2 3 2
26 11 11 11 2 12 1 11 12 1 12 1 11 12 2 13 10 9 0 0 13 3 1 11 2 11 2
30 1 15 2 13 10 3 0 9 13 1 10 9 2 2 11 11 2 2 2 10 9 1 11 11 2 2 2 11 2 2
53 3 1 11 11 2 10 9 0 4 1 13 1 10 9 1 13 10 9 0 1 10 1 10 9 0 1 10 9 2 7 13 13 1 10 9 0 1 11 2 16 15 13 1 10 9 10 0 9 1 10 9 11 2
25 15 13 1 15 1 13 10 9 1 11 1 8 2 11 2 9 1 11 2 15 4 4 13 3 2
59 16 15 13 9 1 10 9 2 15 13 1 11 13 7 13 1 9 1 9 1 10 9 2 16 15 13 0 2 10 9 15 13 1 15 1 10 9 1 16 1 3 13 11 7 11 13 4 13 1 11 2 13 2 10 9 7 1 11 2
33 10 9 0 11 11 13 9 0 1 10 9 0 1 11 2 9 1 10 16 13 10 0 11 16 13 10 0 9 1 11 7 11 2
16 1 12 15 13 9 1 9 7 10 9 1 10 9 1 9 2
41 1 13 1 0 9 2 13 10 9 1 9 1 9 9 1 10 9 13 1 10 9 1 10 9 11 11 11 2 15 16 13 13 10 9 0 1 13 15 1 9 2
47 4 13 15 1 10 0 9 0 7 10 9 1 9 2 10 9 1 11 2 10 9 0 2 9 0 2 10 9 1 11 2 10 9 9 0 2 10 9 0 0 7 10 9 1 9 0 2
30 3 11 15 13 1 11 3 13 10 11 11 11 2 2 11 0 0 2 2 2 1 10 15 13 13 0 9 1 9 2
9 9 1 9 15 13 1 11 11 2
9 3 13 7 3 10 9 16 13 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
4 9 1 10 11
48 1 10 9 1 10 9 1 10 0 9 15 13 10 9 1 10 9 0 1 10 9 7 3 1 10 9 13 1 10 9 1 10 11 2 11 2 11 11 7 11 2 3 7 10 9 1 11 2
35 1 11 2 15 1 10 0 9 0 13 1 13 1 10 9 1 10 11 1 11 2 3 15 13 9 1 10 9 13 1 2 9 0 2 2
24 10 9 2 13 1 9 2 13 1 9 2 11 2 3 13 2 1 9 16 15 13 1 9 2
43 10 9 11 11 2 15 13 1 9 2 13 1 11 1 13 10 0 9 1 10 0 9 3 7 10 9 1 11 11 1 10 11 13 10 0 9 1 11 1 10 0 9 2
52 11 13 10 9 0 1 10 9 2 11 11 11 2 2 1 9 2 11 11 1 9 7 11 1 9 1 9 2 2 16 13 10 15 0 1 10 9 1 9 13 1 10 9 1 13 15 1 10 11 1 9 2
21 1 10 9 4 13 15 1 12 9 2 1 13 0 7 3 2 1 10 9 9 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
27 1 9 2 7 16 11 1 10 9 13 0 1 11 2 15 13 9 1 16 10 9 0 3 13 10 0 2
46 10 9 9 13 9 1 10 9 1 9 16 2 1 10 9 2 13 1 10 9 1 10 9 7 1 10 15 1 10 9 0 1 9 2 9 2 9 7 10 9 1 9 7 9 0 2
9 3 2 10 9 13 1 11 11 2
29 10 9 16 15 4 13 13 16 3 13 0 16 10 9 13 12 9 1 10 9 2 3 7 10 9 3 15 13 2
22 11 11 11 11 13 10 9 0 1 9 1 9 7 13 3 1 12 9 1 9 0 2
49 13 0 1 9 0 1 10 9 0 1 11 2 13 9 1 2 8 11 11 2 1 11 2 13 8 8 8 1 10 9 0 1 11 2 11 2 2 3 1 12 13 10 9 1 9 7 9 0 2
48 1 10 11 11 11 2 13 1 10 9 1 11 11 7 11 11 11 2 1 10 15 13 1 10 9 1 10 9 2 12 2 7 1 15 1 11 11 2 1 15 13 1 2 11 11 15 2 2
25 1 15 10 9 1 9 13 10 9 10 0 9 13 10 11 2 10 11 2 10 11 7 10 11 2
27 1 10 9 15 15 13 2 3 7 3 3 2 10 11 11 0 7 0 7 2 1 9 2 10 12 0 2
17 12 2 13 10 9 7 9 0 1 9 13 3 1 11 10 11 2
37 10 9 13 1 2 3 3 10 9 7 9 2 7 1 10 9 1 9 0 1 10 15 16 15 13 1 9 0 16 13 10 9 1 9 7 9 2
35 10 0 9 1 10 11 1 10 0 9 1 11 11 7 10 0 9 1 10 9 1 10 9 2 10 9 1 12 1 9 2 13 10 9 2
28 3 16 10 9 1 9 4 13 2 11 3 13 10 9 7 9 1 15 2 1 9 1 10 0 9 1 9 2
15 10 9 2 9 1 11 15 13 1 12 9 7 12 9 2
8 1 10 9 15 13 13 3 2
16 10 9 1 9 16 13 9 1 9 7 9 13 1 9 0 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
26 10 9 15 13 1 9 1 10 9 1 10 9 0 1 10 9 0 1 7 3 1 10 12 9 0 2
15 10 9 12 15 13 16 10 9 1 13 4 1 10 12 8
26 3 3 13 1 10 12 8 2 7 2 3 2 1 11 2 7 13 10 9 1 16 4 13 15 3 2
19 16 7 10 9 0 11 11 2 11 2 13 1 10 9 1 2 11 2 2
31 10 9 13 1 12 9 1 10 9 0 2 10 0 9 3 0 13 1 10 9 1 10 9 3 1 2 11 1 15 2 2
22 1 13 1 12 13 9 1 10 11 11 2 11 1 11 7 1 12 7 12 9 0 2
18 11 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
39 13 0 13 16 10 9 3 0 1 10 15 15 4 13 3 4 13 0 7 16 3 15 1 15 13 2 10 4 13 10 9 1 9 1 10 15 13 0 2
14 13 1 9 1 10 0 9 1 10 9 1 11 11 2
33 3 3 13 15 13 1 11 1 10 9 1 9 1 13 10 9 1 10 9 2 13 10 9 7 13 10 9 1 0 9 1 11 2
36 1 12 10 11 1 11 11 13 1 10 9 2 10 0 9 1 12 9 0 0 16 13 10 9 1 15 16 1 10 9 13 10 11 11 11 2
24 13 1 15 2 13 15 13 16 11 13 10 9 7 15 13 16 15 15 13 1 10 9 0 2
14 10 11 11 4 13 1 12 7 10 11 11 1 12 2
21 10 9 11 11 15 13 1 2 10 9 1 9 2 1 0 13 7 15 0 2 2
27 3 13 0 2 7 13 15 0 2 1 0 9 2 0 9 2 9 0 2 9 1 9 2 8 7 8 2
18 10 9 13 1 9 7 13 1 16 15 1 10 9 13 7 4 13 2
12 11 7 11 15 13 1 10 9 1 10 9 8
46 10 9 1 10 9 8 15 4 13 1 9 2 9 7 9 0 1 11 11 11 9 1 10 9 2 16 13 1 10 9 1 11 11 11 11 1 10 10 9 0 1 10 11 11 2 2
49 10 9 0 1 10 11 15 13 3 1 16 10 9 0 1 10 9 2 16 13 10 0 11 1 10 11 2 13 10 9 7 10 9 1 10 9 1 10 9 0 16 13 10 9 11 11 1 11 2
34 13 1 9 16 10 9 13 10 9 3 1 10 10 9 0 2 10 9 13 16 10 9 16 15 4 13 3 4 13 0 1 10 9 2
23 1 11 2 11 13 1 10 0 9 1 10 9 11 1 12 12 9 0 1 10 0 9 2
28 10 9 13 13 10 9 1 10 9 1 12 9 1 9 2 12 9 1 9 2 7 13 12 0 9 1 9 2
20 10 9 13 16 10 9 1 9 0 9 1 11 15 13 1 10 9 12 8 2
39 10 9 2 9 1 10 9 1 10 9 2 4 13 1 0 9 1 15 9 1 10 9 7 0 9 4 13 10 9 1 13 10 0 9 1 4 13 15 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
11 1 12 2 10 9 1 9 0 13 12 2
21 11 11 11 1 11 11 2 12 2 2 13 10 9 2 9 2 9 2 9 0 2
23 13 9 10 9 0 3 15 13 10 9 16 13 10 9 1 10 9 1 10 12 9 2 2
38 10 9 1 10 9 15 13 1 12 9 13 1 9 0 2 7 10 1 10 9 13 10 9 0 1 10 9 13 10 9 1 9 7 10 9 1 9 2
17 16 15 13 1 9 11 13 1 10 9 1 9 10 9 1 9 2
29 1 9 1 9 2 10 9 0 4 13 15 10 3 0 1 10 9 2 1 10 4 13 1 1 10 3 12 9 2
37 13 1 10 9 1 10 9 1 11 2 1 10 9 1 10 9 1 11 2 1 10 9 1 10 9 1 11 7 1 10 9 1 10 9 1 11 2
33 9 1 10 11 11 11 1 10 11 11 11 13 9 0 1 10 9 1 10 9 11 1 11 2 11 2 7 1 10 9 1 11 2
14 1 10 9 1 9 13 7 15 13 3 1 10 9 2
34 1 9 1 10 9 12 13 9 1 10 9 0 2 1 13 1 10 9 1 13 1 13 1 10 9 0 0 1 10 9 1 10 9 2
42 1 11 11 2 9 0 1 10 11 2 2 10 9 7 9 0 13 10 9 7 9 1 10 9 2 16 13 10 0 9 7 10 0 9 1 9 1 10 9 1 11 2
13 13 0 16 10 9 1 0 9 0 13 15 3 2
31 10 9 13 10 0 9 0 16 13 3 3 10 10 9 1 9 1 9 2 1 15 9 10 9 1 9 7 9 2 9 2
18 15 4 13 10 9 3 10 9 13 7 3 9 7 9 1 10 9 2
24 15 1 10 9 1 10 9 2 3 13 1 10 9 1 10 9 2 13 1 10 9 1 11 2
24 0 1 10 9 0 13 10 9 9 1 11 2 3 7 10 9 0 0 1 10 9 1 9 2
15 11 2 3 4 13 2 13 10 9 1 10 9 1 9 2
22 1 10 9 2 10 0 9 13 10 0 9 1 10 11 1 11 2 0 1 10 9 2
28 1 13 1 10 9 3 15 15 13 1 9 7 0 9 16 13 1 10 9 2 13 10 9 1 13 10 9 2
11 15 13 16 15 13 10 9 16 3 13 2
40 16 1 9 3 13 15 0 2 10 9 13 1 10 9 13 16 10 8 13 1 9 0 11 2 1 9 1 10 11 2 16 13 10 0 9 1 10 9 2 2
15 7 1 12 13 10 0 9 13 1 10 9 1 9 0 2
42 10 0 2 10 11 2 15 13 1 10 0 9 1 11 7 11 1 9 1 10 9 1 2 10 11 2 2 10 9 4 13 9 1 10 9 0 2 1 11 1 12 2
61 1 9 2 10 9 13 0 9 1 9 1 10 9 0 1 10 9 7 1 0 9 7 9 2 1 3 10 9 9 2 16 15 13 10 9 7 10 9 13 1 9 1 13 10 9 1 10 9 2 7 2 1 15 2 10 9 1 10 9 2 2
14 3 15 4 13 9 1 9 1 9 1 10 0 9 2
20 15 4 13 1 10 11 13 10 9 3 1 10 9 0 2 3 9 0 2 2
31 11 11 13 10 12 1 11 1 12 1 11 7 13 10 12 1 11 1 12 1 11 2 13 10 9 7 9 1 9 0 2
13 12 9 3 1 13 10 9 4 13 10 0 9 2
15 11 11 2 13 10 9 0 9 1 10 9 1 10 9 2
17 0 7 0 2 11 13 10 9 0 13 1 10 9 0 7 0 2
19 3 1 11 13 1 11 2 11 4 1 13 7 13 1 10 9 1 9 2
10 1 10 9 13 10 9 1 12 9 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
31 3 1 10 9 3 15 4 13 9 4 13 10 9 1 10 9 2 7 10 9 13 10 9 7 9 1 13 10 9 0 2
7 3 3 15 13 10 9 2
16 15 13 1 10 9 1 10 9 0 2 13 1 10 9 0 2
28 11 11 13 10 9 1 9 1 9 1 10 9 1 10 15 15 13 10 8 11 11 11 2 9 1 10 9 2
27 13 3 1 10 15 1 10 9 0 7 0 2 7 11 13 1 11 1 10 9 1 10 9 9 1 9 2
45 10 9 1 9 3 3 15 13 1 10 9 7 1 10 9 0 1 10 9 2 1 9 11 13 1 10 9 1 10 9 0 1 10 11 2 10 11 7 10 9 1 10 10 9 2
19 10 12 1 11 1 12 10 9 13 13 10 9 1 12 9 1 10 9 2
29 10 9 13 0 1 10 9 0 1 9 1 9 2 7 9 0 13 3 3 1 10 9 0 2 16 13 10 9 2
31 10 9 1 9 13 16 13 10 9 1 10 11 1 10 9 1 9 11 7 10 9 13 0 2 3 0 9 1 10 9 2
13 3 13 9 1 9 0 1 10 12 1 10 12 2
50 10 9 1 9 1 10 9 0 1 10 9 1 9 0 1 9 1 10 9 0 2 13 11 2 13 15 1 10 9 1 10 16 13 1 13 15 1 10 9 0 2 10 9 16 3 13 1 13 2 2
21 1 11 1 10 12 15 13 10 9 16 13 1 10 9 13 9 1 9 0 10 2
19 1 12 5 1 11 11 1 10 11 1 11 7 1 12 5 1 11 11 2
55 1 10 9 1 13 10 9 1 10 9 1 11 7 13 10 9 0 0 1 9 1 10 9 2 10 9 11 7 10 9 0 11 11 11 13 1 10 0 9 11 1 11 1 9 0 2 10 9 13 2 10 9 1 11 2
9 10 9 4 13 15 1 9 0 2
33 10 9 1 9 15 13 1 9 0 1 10 9 1 10 9 0 11 7 9 2 1 10 15 11 11 2 13 1 13 10 9 11 2
15 10 11 1 11 11 4 13 1 10 11 1 11 1 12 2
34 11 11 13 1 11 2 11 2 1 9 13 1 11 11 2 11 1 10 11 2 3 13 1 10 9 11 11 11 11 2 11 11 2 2
20 10 9 2 11 11 11 4 13 1 11 1 12 2 16 15 3 13 12 9 2
37 13 3 0 3 7 13 10 9 1 9 1 10 9 1 10 9 1 13 9 1 15 13 7 15 8 3 7 15 13 1 10 9 0 1 0 9 2
31 15 13 10 9 1 16 10 9 0 4 13 3 2 16 2 1 0 2 15 13 16 10 9 0 13 10 9 1 9 0 2
8 13 9 0 16 3 15 13 2
11 12 9 1 11 13 10 9 1 13 15 2
8 15 13 11 7 15 13 11 2
34 11 13 3 10 0 11 1 11 1 11 11 2 12 2 1 10 11 2 10 15 13 1 10 9 1 10 9 1 9 1 9 1 12 2
23 10 9 4 13 16 10 9 13 9 1 9 0 2 16 1 9 15 13 1 9 0 9 2
31 13 12 9 2 10 9 0 13 10 9 1 10 10 9 7 13 3 10 9 1 10 9 1 10 9 16 13 0 1 3 2
10 1 11 2 8 11 2 13 10 9 2
21 13 3 13 10 9 0 16 1 10 9 13 10 9 1 10 9 0 1 9 0 2
30 10 9 0 13 1 13 9 10 10 9 1 10 9 1 10 9 8 1 11 2 11 2 7 10 11 2 11 11 2 2
31 1 10 9 16 4 13 1 10 9 2 13 15 16 15 13 1 10 9 13 2 10 9 1 10 9 2 13 1 10 9 2
14 3 13 1 10 9 11 7 1 10 9 1 9 11 2
38 13 0 1 15 1 10 9 0 1 9 7 9 1 9 2 3 7 1 10 9 1 9 1 9 1 10 9 1 11 2 11 11 7 10 9 11 11 2
22 11 11 13 10 9 0 2 9 0 0 1 0 2 0 2 16 13 1 10 9 11 2
26 15 13 16 11 4 13 2 2 15 3 13 15 2 7 15 16 13 15 2 3 15 9 1 15 2 2
28 11 11 13 10 9 1 9 1 9 13 1 11 11 16 13 9 1 9 2 9 2 9 7 9 1 11 11 2
35 3 1 0 2 10 9 0 4 13 10 0 9 1 10 9 2 1 10 9 16 13 10 9 1 9 1 10 9 11 11 11 2 11 2 2
23 10 9 3 0 1 10 9 16 4 13 1 10 9 11 11 2 4 13 1 9 0 0 2
17 15 13 1 10 0 9 1 10 9 11 2 13 1 9 1 9 2
14 3 3 15 4 4 1 13 10 9 2 1 9 0 2
28 1 10 9 12 13 13 15 10 9 1 11 2 15 16 13 16 11 15 13 13 1 10 0 9 1 10 9 2
20 3 15 13 10 9 1 10 2 9 2 7 3 15 13 10 9 0 1 11 2
24 3 10 9 9 1 10 9 0 2 16 13 1 10 9 1 10 9 7 13 10 9 0 0 2
10 13 3 0 7 13 10 9 1 9 2
9 10 9 7 10 9 13 15 0 2
9 10 9 0 3 0 13 11 11 2
8 11 15 13 13 1 10 9 2
30 1 9 15 15 13 1 10 9 2 9 0 2 9 7 9 0 2 16 13 13 1 10 9 2 10 9 7 10 9 2
15 13 1 10 9 0 1 10 11 2 13 1 13 9 0 2
40 10 9 15 13 10 11 0 13 10 9 2 10 9 0 1 10 9 13 9 1 10 9 0 1 10 9 1 10 9 1 10 9 2 13 15 1 10 11 11 2
35 10 9 11 0 1 10 0 2 12 9 2 2 11 11 2 2 11 2 11 11 2 11 2 7 11 2 13 1 10 0 9 1 10 9 2
11 1 12 2 13 13 9 1 10 9 0 2
18 10 9 1 10 9 1 11 2 13 1 10 9 2 4 13 1 9 2
59 1 10 12 9 2 11 13 0 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
38 11 11 7 10 9 1 10 11 1 11 13 1 10 9 13 1 10 9 0 1 10 9 3 7 11 2 11 7 11 13 1 9 0 1 13 10 9 2
23 3 1 13 7 13 0 9 2 10 12 13 13 1 10 9 1 13 10 9 1 10 9 2
10 10 9 13 1 12 13 1 12 9 2
32 10 9 0 4 13 10 9 1 10 9 16 13 10 9 0 1 11 10 0 9 1 11 1 11 16 13 10 0 8 1 11 2
19 10 0 9 4 13 1 13 1 15 11 13 3 1 11 1 10 9 0 2
20 4 13 1 10 9 16 15 13 1 9 9 2 9 2 0 1 10 9 11 2
57 10 9 1 9 9 2 11 11 2 1 10 9 1 9 0 7 3 0 1 10 9 7 1 9 1 10 16 15 13 0 2 13 16 2 10 9 1 10 9 1 11 13 10 9 16 4 13 1 10 9 16 4 13 10 9 2 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 8 2
35 10 9 13 10 9 1 11 7 10 9 0 2 13 9 0 1 10 9 1 11 11 2 16 13 9 1 10 9 0 1 11 1 10 9 2
19 10 9 13 1 10 12 9 2 10 11 2 7 15 13 10 9 11 11 2
41 1 9 2 16 10 9 0 1 10 9 4 13 2 3 13 10 9 1 13 2 1 15 15 10 9 0 1 10 9 2 13 1 10 9 1 12 2 4 13 15 2
19 10 9 12 7 12 1 11 13 10 9 1 10 11 1 10 11 2 11 2
22 10 9 0 15 13 2 10 9 1 9 2 15 1 9 2 15 0 7 15 1 9 2
12 10 0 9 1 13 9 1 9 1 9 0 2
34 10 11 1 10 11 1 11 13 10 9 10 9 13 1 10 11 1 11 11 7 10 9 4 13 1 10 11 1 11 1 10 9 12 2
29 3 13 9 2 1 10 9 0 2 10 9 1 10 15 3 13 3 3 7 10 9 2 1 10 9 1 10 9 2
63 1 10 12 9 2 10 9 1 11 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
36 11 13 4 13 7 4 13 10 9 1 11 1 11 2 9 16 13 10 9 1 10 11 16 13 16 13 1 10 9 1 10 11 11 1 11 2
43 11 11 2 15 13 10 9 2 15 13 3 1 10 9 1 11 11 2 10 9 1 10 9 13 1 10 9 11 2 2 3 1 10 0 9 0 1 10 9 1 10 9 2
19 1 10 9 1 12 2 10 9 4 13 1 10 9 1 11 11 7 11 2
45 10 9 16 10 0 9 16 13 1 10 9 12 13 1 9 13 1 11 11 13 10 9 1 13 10 9 0 1 10 9 2 1 15 11 11 2 10 9 1 9 1 10 11 11 2
22 3 10 9 13 2 1 11 1 11 2 11 1 11 2 11 11 11 7 10 9 11 2
29 1 9 0 2 10 9 0 13 9 3 3 15 13 2 9 3 3 13 9 7 9 3 15 16 13 13 10 9 2
12 10 9 15 13 1 12 7 11 13 1 12 2
16 4 13 1 10 9 2 9 2 9 7 10 9 1 9 0 2
20 11 11 4 13 10 9 3 0 10 10 9 7 11 15 4 13 3 7 11 2
35 10 9 1 9 0 4 13 1 10 9 12 7 12 2 13 10 9 0 2 10 9 1 9 1 10 9 2 10 9 0 2 7 10 9 2
19 4 13 1 12 3 1 16 10 9 0 15 13 1 4 13 1 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
41 10 9 3 0 16 15 13 13 15 1 10 9 0 11 11 11 2 15 13 16 1 12 11 13 1 10 9 1 11 7 16 1 12 15 13 10 9 1 11 11 2
14 3 4 13 10 9 7 9 1 3 13 1 10 9 2
15 10 12 1 11 1 10 12 2 11 13 10 0 9 0 2
31 10 9 15 13 1 3 1 2 10 10 11 2 2 7 1 15 15 4 13 2 13 2 13 10 9 2 13 10 9 2 2
5 3 13 9 0 2
24 13 1 10 11 11 2 11 2 11 2 11 2 7 15 13 1 10 11 11 1 11 1 12 2
12 10 9 16 13 10 9 0 4 13 1 11 2
35 13 1 11 11 2 10 9 13 1 10 9 16 13 1 10 9 1 10 9 0 9 15 4 13 7 13 1 10 9 1 10 9 1 11 2
75 2 1 10 9 1 16 10 9 1 10 9 13 0 2 3 13 9 1 9 7 9 1 10 9 2 2 13 10 9 2 15 13 16 2 1 10 9 2 10 9 13 10 9 0 7 13 0 1 10 9 7 3 10 0 9 1 11 2 15 3 13 1 9 1 10 16 13 10 9 1 10 9 1 11 8
9 13 10 9 1 11 1 11 11 2
47 10 9 13 10 9 1 9 1 10 9 2 7 1 10 9 1 10 9 1 10 9 4 13 10 9 0 16 3 13 0 1 11 12 2 13 3 1 10 9 1 10 9 1 9 1 9 2
19 10 11 12 15 13 1 9 1 9 2 13 12 9 1 10 9 1 9 2
27 10 0 9 1 10 9 15 13 1 11 10 8 0 7 13 10 9 1 9 0 0 7 9 1 9 0 2
35 15 4 13 7 13 10 9 1 11 2 13 10 0 9 1 10 9 7 13 13 16 10 9 1 11 13 10 9 7 13 9 1 10 9 2
28 10 9 4 13 1 12 9 13 3 1 10 9 2 16 13 1 10 9 0 13 1 9 7 13 1 10 9 2
25 1 10 0 9 1 11 11 2 1 12 7 12 2 10 9 2 11 11 2 13 1 10 9 12 2
26 15 4 13 15 10 9 1 13 1 3 1 10 9 2 10 9 7 10 9 13 1 11 7 10 9 2
5 13 10 9 11 2
24 10 9 4 7 13 16 13 13 1 10 9 16 4 7 13 15 3 1 3 1 9 1 9 2
24 13 10 9 1 12 9 2 7 13 10 9 10 12 2 16 4 13 1 10 9 1 10 11 2
20 13 16 10 9 13 1 16 15 3 4 1 13 1 10 9 13 1 10 9 2
22 10 11 11 13 10 9 1 9 0 7 10 9 1 9 1 10 9 0 1 10 9 2
17 9 12 10 0 9 13 3 2 7 3 3 15 13 1 10 9 2
26 13 1 10 9 2 11 4 13 3 1 10 9 1 10 9 1 9 1 11 16 15 13 1 9 0 2
48 10 12 5 1 11 1 12 2 10 9 1 10 11 2 11 11 11 2 13 16 10 11 13 3 1 10 11 7 15 13 16 4 13 12 9 2 12 1 3 1 15 13 1 10 0 9 0 2
8 11 15 13 13 1 10 9 2
26 16 10 0 9 1 11 11 13 3 1 9 0 2 11 11 13 1 9 0 10 0 9 1 10 9 2
20 13 9 7 1 10 9 1 9 13 9 1 10 9 1 13 10 9 3 3 2
22 15 13 1 12 9 1 9 7 1 12 9 1 10 9 1 11 2 10 9 1 9 2
36 1 10 9 2 10 9 0 3 0 4 4 13 16 13 1 10 0 9 3 15 13 10 0 9 10 0 9 1 10 9 1 10 0 9 11 2
18 10 9 13 0 7 10 9 4 13 0 1 9 12 1 10 9 0 2
38 1 10 9 2 10 9 13 1 10 10 9 0 2 1 10 0 7 1 10 10 9 0 2 1 9 1 11 2 3 15 13 10 9 1 10 12 5 2
24 15 13 10 8 1 10 9 1 11 11 2 11 7 11 2 15 4 13 3 1 10 9 12 2
63 10 9 0 1 2 11 2 4 13 1 9 1 11 1 12 1 10 11 2 11 7 13 10 0 9 15 11 13 1 10 9 11 11 2 15 3 3 13 9 1 2 11 1 11 2 2 2 11 11 2 2 2 10 11 11 2 7 2 11 1 11 2 2
22 11 2 11 2 2 11 2 11 11 2 11 11 2 11 2 11 2 11 11 7 11 2
33 10 9 11 3 13 10 9 1 10 9 1 10 0 9 2 7 16 10 9 4 13 1 10 9 0 2 15 13 1 13 10 9 2
24 10 9 4 13 0 2 4 13 15 2 15 4 13 15 3 2 2 13 1 10 9 1 11 2
54 3 1 13 10 9 1 9 1 10 9 1 9 2 10 9 1 9 1 10 9 7 2 3 2 10 9 1 10 9 1 0 9 1 10 9 1 12 9 2 7 13 10 9 1 10 9 1 10 9 15 13 3 0 2
34 15 2 9 1 10 9 7 1 10 9 0 1 10 11 0 2 13 1 10 0 9 1 16 13 9 1 10 9 7 1 16 15 13 2
23 1 10 0 9 10 9 13 1 0 9 1 3 1 10 9 16 13 0 1 10 9 0 2
13 10 9 13 1 13 3 10 9 0 1 10 11 2
30 10 9 0 13 10 9 0 1 11 1 11 11 2 10 9 1 10 9 1 11 2 11 2 2 13 1 10 9 12 2
35 10 9 11 11 3 13 1 9 0 2 11 11 2 1 10 9 12 1 10 15 15 13 1 10 9 13 1 10 9 1 11 11 1 11 2
21 9 1 9 11 11 11 10 11 7 11 7 1 11 11 11 11 1 11 7 11 2
4 9 0 0 2
42 10 11 11 1 10 11 11 4 13 1 10 9 13 12 8 2 12 2 7 3 15 13 12 9 2 1 9 1 10 0 9 1 9 0 16 13 10 12 9 1 9 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
34 3 13 9 1 9 1 10 11 1 11 2 1 11 11 2 2 12 7 12 2 7 1 15 1 11 2 1 11 11 2 2 12 2 2
29 1 12 10 9 13 1 10 11 11 11 1 10 9 1 11 11 11 11 1 10 9 11 11 7 10 9 11 11 2
11 1 4 13 2 11 13 13 1 10 9 2
21 1 10 9 1 11 1 11 2 9 15 13 1 9 1 9 0 1 9 1 9 2
17 11 13 10 9 1 12 9 1 9 1 9 0 1 10 9 11 2
9 9 2 10 9 12 3 13 9 2
41 10 9 13 16 10 9 4 13 10 12 1 11 1 12 2 7 16 10 9 16 15 10 9 15 4 13 1 10 0 9 2 11 2 3 4 4 13 1 10 9 2
19 1 9 13 10 9 1 10 9 7 10 9 4 7 13 1 10 9 13 2
34 15 13 12 9 3 3 2 7 10 9 15 13 3 1 9 1 10 9 7 10 10 9 16 15 13 1 13 1 10 9 1 10 9 2
29 10 9 0 2 3 7 3 10 9 1 9 1 9 13 1 11 1 2 13 9 1 10 9 1 9 3 0 2 2
13 10 9 1 9 4 13 3 1 10 9 11 11 2
16 10 9 1 10 9 13 0 1 10 9 7 0 11 1 11 2
17 1 10 11 1 10 11 1 11 2 13 10 9 1 9 7 9 2
39 10 9 15 13 16 4 13 1 10 9 1 2 10 9 2 10 9 7 10 9 2 1 10 9 2 1 9 1 10 9 13 1 10 9 0 1 10 9 2
17 13 0 1 9 2 1 15 10 9 0 2 7 3 13 10 9 2
22 11 11 11 2 2 10 9 2 2 1 11 2 13 10 9 1 9 1 11 2 11 2
24 11 13 13 10 9 1 9 2 7 13 9 1 11 11 2 10 9 2 16 13 1 10 11 2
30 4 4 13 10 11 2 1 11 2 7 1 9 1 16 3 13 1 10 9 13 16 15 4 1 13 1 13 9 2 2
17 9 1 10 0 9 0 0 2 1 9 13 10 0 9 0 0 2
53 7 10 9 16 10 9 13 10 9 16 13 0 13 0 13 10 9 0 1 11 1 10 9 0 2 1 9 0 2 9 2 9 2 1 9 0 1 9 0 2 9 1 9 9 7 9 0 7 9 0 1 9 2
20 11 13 13 15 1 10 9 1 15 3 1 11 2 16 13 13 15 1 15 2
28 13 1 10 9 0 1 0 9 2 11 13 3 13 10 9 16 15 13 1 10 9 10 12 1 11 1 12 2
32 3 16 3 13 3 2 3 13 1 15 13 16 15 13 7 3 13 1 10 9 16 10 15 11 4 13 16 13 0 1 15 2
28 11 13 10 9 13 1 10 9 13 1 10 9 1 11 7 10 9 1 11 11 2 1 10 9 0 1 11 2
28 10 9 15 13 1 10 9 1 10 9 0 2 7 1 10 9 4 13 1 10 9 16 15 13 1 10 9 2
20 13 9 1 9 1 9 1 10 9 3 2 1 15 15 10 9 0 13 0 2
13 1 12 11 13 1 11 7 11 13 1 11 11 2
18 1 12 2 13 1 10 9 0 7 0 1 10 9 11 16 15 13 2
17 10 9 13 0 7 0 2 1 10 9 13 10 9 7 10 9 2
25 1 9 1 10 12 5 1 10 9 7 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
15 11 15 13 1 11 2 0 9 2 3 9 1 11 11 2
36 1 13 10 9 2 11 13 10 9 13 1 10 11 1 10 11 11 2 11 8 11 2 7 11 11 1 10 9 0 2 11 2 1 8 12 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
30 1 10 12 10 9 1 9 0 1 10 9 1 10 9 13 1 12 9 7 10 9 0 1 10 9 13 1 12 9 2
19 10 9 1 10 9 13 1 16 13 10 9 1 10 15 10 9 15 13 2
26 11 11 2 11 2 11 1 11 2 11 2 12 1 11 1 12 2 13 10 9 7 9 1 9 0 2
24 1 11 2 10 9 13 1 10 9 10 11 12 1 11 1 10 12 1 10 12 8 1 11 2
32 11 2 13 1 11 2 9 0 1 11 2 7 16 10 9 0 9 13 1 10 9 1 10 11 11 0 2 7 1 9 0 2
12 11 15 13 1 9 0 1 9 1 10 9 2
50 15 4 13 10 0 9 1 10 9 1 9 2 7 3 15 13 0 9 1 10 9 1 10 9 0 1 10 0 9 2 15 16 13 10 0 9 1 10 9 1 10 9 1 9 13 1 10 9 0 2
16 1 13 1 3 10 9 15 13 1 9 1 10 9 1 11 2
15 11 11 13 10 0 9 0 16 13 1 10 9 1 11 2
11 13 3 10 12 2 12 2 12 7 12 2
5 15 13 1 11 2
12 10 9 1 9 1 10 9 13 1 5 12 2
15 13 11 2 0 1 9 10 9 16 13 9 1 10 9 2
37 10 9 1 10 9 13 10 12 2 10 9 13 1 10 9 1 1 11 7 10 12 9 1 10 12 9 2 10 9 15 13 1 9 1 11 2 2
10 10 9 1 9 3 13 10 9 0 2
25 10 9 13 1 10 9 1 10 11 1 13 1 10 0 9 13 3 13 11 11 2 11 11 2 2
22 10 8 2 11 1 11 11 2 11 13 1 10 9 1 13 1 16 15 13 10 9 2
50 1 10 9 13 10 9 1 10 9 11 11 11 1 10 9 1 10 11 2 3 15 13 13 10 9 1 11 11 2 16 10 9 4 13 1 9 1 9 1 10 9 2 3 13 3 1 10 11 11 2
19 10 9 4 13 3 1 10 9 9 13 11 16 15 13 3 1 9 0 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
26 10 9 1 11 2 1 9 2 11 11 2 2 13 1 12 2 13 10 9 1 10 9 0 1 11 2
10 3 13 10 9 1 10 11 1 11 2
9 15 13 16 3 13 2 16 13 2
9 4 13 1 0 9 0 7 0 2
5 2 3 13 15 2
59 3 13 1 10 9 1 10 11 2 15 13 1 10 9 1 10 9 12 1 10 11 11 2 13 9 0 3 1 10 9 2 13 1 10 9 12 1 10 9 0 2 3 13 1 9 1 10 9 1 10 9 0 1 11 2 11 7 11 2
16 13 3 0 1 10 0 9 2 13 1 10 9 1 10 11 2
49 13 13 1 11 7 11 2 16 15 13 16 2 10 10 9 2 4 13 1 10 9 7 10 9 16 13 10 9 0 7 15 13 1 10 9 0 10 9 1 10 9 2 7 10 9 1 15 9 2
40 3 1 10 9 11 11 7 11 2 3 9 2 13 10 9 1 10 9 0 1 10 9 10 9 0 1 11 2 13 7 13 1 10 11 11 1 11 1 12 2
26 10 9 0 2 10 9 3 0 2 10 9 3 13 2 10 9 1 9 0 7 15 1 10 9 0 2
22 1 9 2 3 13 10 9 0 1 10 9 1 9 0 1 10 9 1 15 16 13 2
29 10 0 9 0 2 11 11 11 2 16 15 13 1 11 2 4 13 10 9 1 11 7 13 9 1 10 0 9 2
17 1 10 9 10 9 13 0 3 1 15 15 13 7 13 10 9 2
9 9 0 0 1 10 11 7 9 2
30 10 9 13 1 10 9 2 13 10 1 10 9 1 10 9 0 2 11 11 2 2 10 15 13 1 10 9 10 9 2
15 11 11 1 10 9 1 12 13 16 13 1 12 7 12 2
37 13 1 10 9 1 10 9 1 11 7 11 2 1 10 9 1 11 2 1 10 9 1 11 7 11 2 7 1 10 9 1 9 2 11 7 11 2
38 16 1 10 9 2 9 8 0 0 15 13 1 10 9 2 1 7 3 1 10 9 2 3 7 3 1 10 9 10 9 2 3 7 3 1 10 9 2
17 10 9 1 10 9 0 7 15 13 10 0 9 15 13 11 11 2
18 10 9 1 2 11 1 11 2 4 13 1 10 9 1 9 0 11 12
8 10 9 15 13 1 10 9 2
16 10 12 9 13 10 12 9 1 11 2 10 9 7 10 9 2
27 10 9 1 10 9 13 3 3 2 10 9 4 13 1 10 0 9 7 9 0 2 13 10 9 11 11 2
28 10 9 4 13 3 1 10 10 9 0 1 10 9 0 2 13 10 9 1 10 9 0 1 10 9 11 11 2
29 14 2 13 9 1 9 7 3 1 13 1 10 9 1 9 13 1 10 9 1 11 1 9 1 15 1 10 9 2
67 10 9 10 11 11 13 10 9 1 13 1 13 1 10 9 2 1 10 9 7 1 10 9 3 7 13 10 9 16 13 9 0 7 0 2 13 16 1 9 1 16 13 3 3 13 10 9 1 11 7 11 2 3 1 16 10 9 13 10 9 1 9 7 9 1 9 2
25 1 10 0 9 1 9 0 2 10 0 9 9 13 1 10 9 1 9 1 10 9 1 9 0 2
16 10 9 0 0 1 11 13 13 2 10 9 2 1 9 0 2
17 3 2 10 9 4 13 16 13 1 10 9 9 16 13 10 9 2
38 1 11 11 2 11 7 11 1 11 2 11 13 10 0 9 1 9 1 11 2 13 1 10 9 10 9 1 10 9 2 3 11 11 11 7 11 11 2
35 10 9 13 0 0 7 0 2 0 1 9 1 10 11 1 10 0 9 1 9 0 10 15 15 13 1 10 9 7 16 13 1 10 9 2
26 13 9 0 1 12 9 2 13 1 9 0 16 13 9 1 0 9 7 13 10 9 1 10 0 9 2
24 11 13 10 0 9 1 9 1 10 9 1 11 11 0 11 2 13 10 12 1 11 1 12 2
32 15 13 13 1 11 1 10 11 1 13 10 9 1 10 9 7 1 11 1 11 1 13 1 10 9 10 9 1 10 9 0 2
19 10 11 13 13 1 10 9 0 1 0 2 16 13 1 11 1 9 2 2
17 10 9 1 11 13 9 13 10 9 1 10 9 13 9 1 9 2
13 10 9 1 10 9 0 4 3 13 1 10 9 2
40 3 2 15 13 16 10 9 4 13 13 10 9 16 13 1 10 9 1 10 9 1 9 1 9 1 10 9 0 7 1 10 9 1 10 9 1 10 9 1 11
58 10 9 0 3 15 13 1 15 7 1 10 9 11 11 1 9 0 0 10 15 7 13 15 1 9 0 1 10 9 1 13 1 15 1 9 1 13 10 9 1 10 11 7 3 13 15 1 16 13 0 1 9 1 16 10 11 13 2
26 9 1 15 2 13 0 13 9 0 1 10 9 1 9 2 9 1 9 8 7 8 2 7 10 9 2
28 2 13 9 16 3 15 13 1 10 11 7 15 13 15 0 2 16 4 13 15 1 10 10 9 2 2 13 2
14 10 9 1 9 13 1 10 9 1 9 13 1 9 2
30 10 9 1 11 1 10 0 9 7 13 1 9 13 1 9 0 2 15 4 13 1 9 7 15 13 1 10 9 0 2
65 13 13 1 10 9 12 7 13 1 10 9 1 10 11 2 11 2 1 12 1 10 0 9 0 0 1 11 7 11 11 2 1 10 9 1 10 9 7 9 2 10 9 11 11 11 2 1 10 9 1 9 7 10 9 1 9 0 1 10 9 7 10 15 13 2
21 11 11 4 3 13 1 10 9 3 0 1 10 9 1 10 9 0 1 10 11 2
16 11 13 10 9 0 1 9 0 0 1 10 9 1 10 9 2
88 2 11 13 3 0 1 13 7 3 13 16 15 13 15 0 16 15 13 1 10 0 9 0 2 7 15 11 2 7 11 7 15 2 16 3 13 10 11 0 2 13 16 4 1 13 10 9 1 9 3 0 7 10 12 9 1 11 11 2 2 13 15 1 0 9 1 10 0 9 2 13 10 0 9 1 12 7 1 13 13 16 10 9 13 1 10 9 2
22 10 9 2 8 2 2 3 13 1 9 2 13 10 9 13 1 10 9 1 10 9 2
78 3 13 9 1 16 4 13 15 9 1 10 9 1 10 9 7 1 10 9 1 9 13 9 1 13 15 7 13 15 2 1 15 15 2 3 4 13 10 9 1 10 9 16 2 1 10 9 2 1 10 9 7 10 9 16 13 2 4 13 2 7 1 15 0 9 2 3 3 1 10 9 0 7 1 10 9 0 2
10 3 13 9 1 10 9 1 10 9 2
35 15 13 10 9 16 13 9 1 10 9 0 2 1 9 0 2 7 16 13 10 9 1 10 9 7 10 9 0 1 9 1 10 9 0 2
22 11 7 11 2 10 9 0 13 10 0 9 0 1 9 15 4 4 13 1 11 11 2
18 10 9 13 10 9 0 1 5 12 9 1 10 5 12 1 10 9 2
56 1 10 9 2 1 0 9 7 9 0 2 10 9 13 1 10 9 0 2 1 15 10 12 9 13 1 9 7 2 1 10 3 13 3 1 15 2 10 9 1 9 3 13 0 1 10 9 0 1 10 9 7 1 10 9 2
9 4 13 10 12 1 11 1 12 2
45 10 11 1 11 13 10 9 0 0 13 10 12 1 11 1 12 1 10 9 11 12 2 13 3 9 1 10 11 11 1 9 1 11 1 11 7 11 2 9 0 1 10 11 11 2
42 1 10 9 1 9 4 13 3 0 10 9 1 9 7 9 2 16 15 1 15 15 4 13 10 9 1 9 2 16 13 13 15 1 10 9 1 11 3 1 10 9 2
25 1 10 3 9 1 11 1 10 9 0 15 13 16 10 9 0 13 1 15 7 13 15 3 0 2
14 13 3 0 3 15 4 8 10 9 0 1 10 9 2
26 10 9 13 16 1 15 15 13 16 10 9 1 11 11 13 0 2 1 11 13 3 9 1 10 9 2
41 13 1 10 9 1 9 2 10 9 1 9 4 13 13 1 10 0 9 0 2 13 13 2 10 9 1 10 9 4 4 13 3 7 13 13 10 9 1 9 2 2
13 10 9 1 9 13 1 12 8 2 2 9 8 2
11 10 9 1 10 9 13 11 7 11 11 2
10 10 9 4 13 1 11 11 1 12 2
19 9 3 0 2 1 3 0 7 0 0 2 3 0 2 9 0 2 9 2
57 15 13 16 10 9 7 9 0 1 10 9 1 9 3 13 10 9 1 11 2 7 10 9 1 10 9 7 16 10 9 1 9 7 9 4 13 15 1 9 1 10 9 1 11 2 1 10 9 1 9 7 10 9 1 10 9 2
39 10 9 0 1 11 13 1 10 9 1 10 9 3 13 10 9 2 8 8 2 12 2 0 10 9 1 10 9 0 7 15 1 10 9 1 10 9 0 2
7 10 9 1 9 13 0 2
25 15 13 10 0 9 1 9 1 15 9 1 10 9 11 0 1 11 2 11 13 3 1 10 9 2
15 11 11 2 13 10 9 1 9 0 0 1 10 9 11 2
3 9 0 2
11 11 3 13 16 13 13 9 0 7 9 2
33 15 13 16 10 9 0 13 10 9 0 2 1 9 11 11 2 1 10 9 16 10 9 3 4 13 10 9 16 13 0 9 0 2
31 3 13 10 9 2 2 4 13 1 11 10 0 9 2 9 1 11 2 16 1 10 9 13 1 10 9 1 10 9 2 2
28 10 9 0 13 10 9 1 10 9 1 12 8 12 8 12 8 3 7 10 9 15 13 1 10 12 9 0 2
33 11 11 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 13 10 8 9 1 9 0 16 13 1 12 9 1 10 11 2
15 13 10 11 0 2 15 1 10 0 9 1 9 0 9 2
22 11 13 3 1 10 9 7 15 13 2 13 15 1 11 16 15 13 10 9 1 15 2
21 10 11 11 13 10 9 0 1 9 0 16 15 13 3 1 10 0 9 1 11 2
12 10 9 1 10 9 13 9 1 8 2 8 2
32 10 9 1 11 12 1 9 1 12 9 1 9 4 13 10 9 1 9 1 10 9 12 7 10 15 1 9 1 10 9 12 2
28 15 0 2 13 1 10 9 7 9 1 10 9 13 1 10 9 7 9 15 1 10 9 3 0 1 10 9 2
8 10 9 13 3 1 10 9 2
32 11 2 9 1 11 11 2 11 2 13 10 9 0 2 0 1 10 9 11 1 9 1 10 11 11 1 11 11 11 1 11 2
45 10 9 4 13 15 13 10 9 2 1 10 9 1 13 10 9 11 2 15 16 13 1 10 9 13 9 1 9 7 1 9 1 10 13 10 11 1 10 0 7 10 9 1 9 2
16 1 10 9 0 7 10 0 9 1 11 2 11 14 10 9 2
22 13 10 9 0 2 1 9 0 2 7 0 9 1 11 9 2 11 2 1 11 11 2
20 1 9 1 9 15 13 10 9 0 2 13 1 13 10 9 0 1 10 9 2
13 10 9 13 1 10 0 9 1 11 1 10 12 2
28 10 9 13 9 7 9 1 11 11 2 16 1 13 9 1 10 9 1 10 9 1 11 11 13 1 9 0 2
33 1 4 13 0 10 9 11 13 10 9 1 10 9 2 13 13 10 9 1 11 11 1 11 1 11 2 13 10 9 0 1 11 2
10 4 13 11 2 11 2 11 7 11 2
53 3 3 2 1 10 9 2 10 9 13 1 11 2 11 2 11 2 11 2 3 10 9 13 1 9 1 10 9 11 12 1 11 10 12 1 11 2 7 10 9 0 13 10 12 5 1 11 4 13 1 10 9 2
55 4 4 13 1 10 9 2 1 10 0 9 2 7 1 10 11 11 2 2 13 9 1 10 9 0 2 7 1 10 11 11 2 12 2 2 7 4 13 10 9 3 0 2 13 1 9 2 15 15 13 0 1 10 9 2
15 13 1 10 9 0 11 7 1 10 9 12 1 10 9 2
23 16 13 13 16 4 1 13 3 0 1 10 9 16 13 2 7 15 3 3 1 10 9 2
19 15 13 3 11 15 13 7 16 4 13 10 11 1 13 10 9 1 9 2
40 13 13 16 11 11 13 12 9 1 10 9 1 10 11 1 10 9 8 12 2 16 10 9 1 10 9 0 13 1 13 1 10 9 1 9 0 1 10 9 2
44 10 9 13 10 12 1 11 1 10 9 11 1 10 11 13 1 11 1 0 9 13 1 10 9 11 11 2 15 13 12 5 2 7 11 11 2 16 13 12 5 2 3 0 2
6 15 13 1 9 0 2
26 10 11 4 13 1 10 3 0 9 0 1 11 2 9 13 13 9 1 9 0 1 0 9 1 9 2
23 13 9 1 10 9 10 12 1 11 1 12 7 1 10 9 15 13 0 9 1 10 9 2
16 10 9 13 15 1 10 9 3 0 1 10 15 15 13 9 2
12 15 13 10 0 7 0 9 1 10 9 0 2
33 1 9 2 15 15 13 1 13 1 11 2 11 12 2 2 9 1 10 9 2 1 15 13 13 2 13 15 3 10 9 11 2 2
36 13 10 12 1 11 1 12 2 16 13 1 12 9 13 10 9 2 11 11 11 11 11 2 13 1 10 9 1 10 9 0 2 11 11 11 2
40 10 9 4 13 1 9 1 10 9 0 1 11 12 1 11 2 16 13 15 10 9 1 10 11 1 11 2 11 12 7 11 11 1 9 2 0 9 1 12 2
25 10 0 9 1 9 2 15 13 1 10 9 1 10 9 1 10 9 2 10 9 7 10 11 2 2
28 1 9 2 10 9 0 13 1 11 13 10 9 1 10 9 1 10 9 11 2 10 9 1 10 9 11 2 2
11 13 12 9 2 1 10 12 3 1 11 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
6 13 0 1 10 0 2
32 13 10 9 2 1 10 9 13 9 2 3 13 10 9 16 13 15 1 9 2 3 9 2 3 13 10 0 9 16 15 13 2
14 9 0 11 11 2 9 1 11 2 11 2 12 2 2
40 3 2 1 10 13 15 1 10 9 1 10 0 9 2 16 3 15 13 9 1 13 10 9 2 11 15 13 0 1 10 9 7 13 16 2 10 9 13 2 2
35 13 3 2 16 15 13 1 13 1 10 9 1 10 9 7 10 9 1 10 9 2 1 10 9 7 1 10 9 2 15 13 1 10 9 2
34 1 0 13 16 13 16 10 9 4 13 1 7 1 15 2 1 10 0 9 1 13 15 7 13 15 1 10 15 9 1 10 9 0 2
21 15 13 1 10 9 2 11 2 1 11 2 0 1 10 9 2 11 2 1 11 2
58 1 15 1 10 9 1 10 9 2 10 9 9 1 10 0 9 16 13 16 3 13 10 9 0 1 10 9 1 10 11 11 2 1 9 1 10 9 1 10 11 1 13 15 12 9 1 10 0 9 2 1 15 15 3 13 1 9 2
9 13 1 9 1 13 1 10 9 2
36 3 13 10 9 1 9 13 1 10 9 1 9 8 2 15 15 13 1 10 9 16 13 1 10 9 1 10 11 11 2 12 9 1 12 13 2
25 13 10 9 1 10 11 11 11 2 15 4 13 1 10 0 11 1 11 2 1 10 9 1 13 2
13 3 15 15 13 13 10 9 1 13 1 10 9 2
10 13 1 10 9 0 2 13 13 9 2
10 3 2 10 9 0 0 13 10 9 2
9 0 16 3 4 1 13 10 9 2
23 1 10 0 9 15 13 10 9 1 0 9 1 11 1 11 1 10 9 0 1 0 9 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
47 11 11 13 15 1 10 9 16 0 9 4 13 10 9 1 10 9 0 7 13 16 10 9 13 1 10 1 10 9 2 7 13 1 9 7 11 15 15 4 13 1 15 3 13 3 0 2
21 11 11 4 13 1 11 11 7 13 1 11 11 12 2 12 2 1 10 9 12 2
31 10 9 13 1 15 1 10 9 1 10 9 3 0 1 10 15 13 2 3 10 9 1 9 1 10 9 1 11 7 11 2
11 3 13 16 15 13 10 9 1 10 9 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
43 15 1 10 0 9 2 7 3 10 3 0 2 16 13 10 9 0 13 10 9 0 1 10 9 2 16 13 1 10 9 1 10 9 15 1 10 9 3 0 1 10 9 2
15 13 10 9 0 7 0 1 9 2 9 7 10 0 9 2
10 10 9 1 9 0 13 10 0 9 2
16 10 9 13 12 5 2 15 1 10 9 1 9 7 1 9 2
20 10 9 15 13 1 15 2 15 13 10 9 1 10 9 2 7 3 15 13 2
11 15 13 10 0 9 14 2 0 7 0 2
29 1 9 2 10 9 0 13 10 9 1 11 1 11 2 13 1 10 9 0 15 1 10 9 3 0 1 10 9 2
22 1 10 9 1 10 11 11 1 12 2 11 13 10 9 1 9 1 13 10 11 11 2
13 11 11 11 11 2 13 16 15 13 10 9 0 2
32 10 11 1 11 4 13 1 11 11 2 9 1 10 9 2 3 1 4 13 10 9 1 9 0 15 13 10 9 1 9 0 2
47 10 9 1 10 9 1 11 2 11 11 2 13 3 10 2 9 2 1 10 9 2 16 13 10 9 16 15 4 13 10 0 9 16 4 13 1 10 9 1 11 7 10 2 9 0 2 2
23 9 3 13 0 1 11 1 10 0 9 0 1 11 2 12 2 13 1 0 9 1 11 2
19 11 11 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 0 2
30 10 9 13 10 9 1 10 0 9 7 9 1 10 9 13 1 10 9 1 9 3 0 13 1 10 15 13 10 11 2
26 10 9 11 11 13 1 10 9 12 2 13 1 9 1 9 1 11 1 11 7 13 1 10 9 0 2
32 10 9 13 10 9 1 10 11 2 11 13 1 10 11 11 11 1 11 1 12 13 1 10 11 11 10 9 12 1 10 9 2
16 3 2 1 10 9 12 2 12 2 13 1 0 9 1 11 2
10 11 11 11 13 1 11 11 2 11 2
31 3 15 13 2 7 15 9 13 16 15 15 13 15 0 2 3 15 13 10 9 1 9 2 16 3 13 7 9 13 0 2
12 15 13 1 10 9 1 10 11 1 10 11 2
35 10 9 11 11 4 13 1 10 9 0 13 10 9 1 10 9 1 10 9 11 11 11 1 0 7 0 9 0 1 10 9 0 1 11 2
11 10 9 13 10 9 0 1 12 9 0 2
28 10 9 15 13 1 3 9 1 9 0 1 9 0 7 0 2 1 10 9 2 9 2 9 2 9 7 9 2
15 13 12 9 1 9 7 13 9 1 10 9 0 1 11 2
31 11 11 2 1 11 2 8 8 2 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 13 10 8 9 1 11 2
29 15 15 13 2 1 11 11 2 9 1 10 9 7 9 1 10 11 11 2 2 1 8 8 16 8 5 8 2 2
15 11 13 10 9 0 1 9 0 2 13 1 10 9 11 2
41 10 9 16 3 4 1 13 1 10 9 3 4 13 9 1 10 0 9 8 2 8 2 1 10 16 4 7 13 10 9 13 1 10 9 1 10 11 2 12 0 2
15 10 9 4 13 3 13 0 10 2 9 2 7 10 9 2
47 10 9 0 13 16 10 9 3 0 1 10 9 13 10 11 11 7 11 0 2 7 13 16 1 10 9 2 3 13 9 1 10 9 0 2 7 1 9 7 1 10 9 16 13 1 13 2
40 1 9 2 13 10 9 1 10 9 13 0 1 10 9 13 1 10 9 2 1 15 15 10 9 15 13 1 13 9 1 10 9 1 10 9 7 1 10 9 2
11 3 13 10 12 9 2 13 11 7 11 2
48 3 2 15 13 10 9 1 10 9 1 11 1 9 0 1 10 9 1 10 9 1 0 9 7 10 9 1 9 13 1 9 1 10 9 2 10 9 2 10 9 2 10 9 7 10 9 0 2
7 11 11 13 10 9 0 2
20 15 1 10 0 9 1 13 9 1 10 9 3 0 13 10 9 1 9 0 2
47 10 11 2 12 4 13 1 10 9 12 1 10 9 1 9 7 9 0 11 1 10 9 1 9 0 0 13 1 13 10 9 1 9 0 7 1 9 1 9 0 13 1 10 9 3 0 2
17 15 13 1 13 1 10 9 16 13 1 10 9 0 1 10 9 2
21 1 3 1 10 9 2 1 10 9 2 13 3 10 9 16 4 13 1 10 9 2
9 15 13 10 9 7 13 10 9 2
12 10 9 1 9 1 10 9 13 1 9 12 2
29 10 9 15 13 1 11 1 12 7 1 10 9 1 10 9 1 10 9 1 11 2 10 9 15 13 1 12 9 2
38 1 10 9 13 1 10 11 1 11 2 11 11 13 16 2 16 10 9 13 10 9 1 10 9 13 1 11 13 10 12 5 1 10 12 0 9 2 2
41 2 1 10 9 1 9 15 4 13 10 9 1 10 9 7 15 4 13 10 9 0 3 15 13 9 0 1 10 9 0 2 3 13 0 10 9 0 2 2 13 2
18 11 13 10 9 1 10 9 1 11 2 9 1 10 11 1 10 11 2
24 3 2 15 13 1 10 9 11 1 11 2 11 2 7 1 10 11 10 9 1 13 15 13 2
34 3 13 16 16 13 1 9 10 9 15 13 1 10 9 1 10 9 2 13 10 9 16 13 10 9 3 1 13 15 1 13 10 9 2
38 1 11 13 13 1 10 0 9 1 9 7 9 2 13 0 9 1 9 1 10 9 1 9 1 10 9 0 2 13 10 9 1 9 7 1 10 9 2
34 16 15 13 9 1 15 1 10 9 1 9 0 7 9 0 13 3 2 1 3 13 8 4 13 10 9 1 10 9 7 1 10 9 2
53 10 11 11 1 11 2 1 9 13 1 9 2 1 9 14 2 11 11 11 2 13 1 11 2 11 2 13 10 9 13 1 9 0 1 9 13 1 13 10 9 1 9 7 9 1 15 9 1 10 10 11 11 2
30 16 15 13 1 15 11 13 1 9 3 0 1 10 9 11 7 10 9 11 13 15 9 1 11 1 3 3 12 9 2
43 13 9 1 10 9 1 11 16 13 10 9 1 10 9 2 2 11 11 11 2 2 7 16 13 3 10 9 0 1 10 9 2 16 3 13 10 9 0 0 1 10 9 2
50 1 10 9 2 10 9 4 1 13 7 13 10 9 2 15 16 13 10 9 1 10 9 2 16 15 13 16 15 15 4 13 10 9 2 1 10 9 2 1 10 9 2 7 3 2 1 10 9 2 2
16 10 0 9 1 9 2 9 7 9 0 15 13 0 1 9 2
42 10 9 1 11 2 1 9 1 11 2 13 10 9 0 0 13 1 10 9 11 12 10 12 1 11 1 12 1 11 11 7 11 2 11 1 11 2 11 7 11 11 2
23 10 9 1 9 1 9 15 13 3 2 13 1 9 1 12 9 1 9 1 10 0 9 2
12 1 10 9 1 12 13 10 9 1 12 9 2
29 10 9 13 1 10 2 12 1 10 9 1 9 1 10 11 11 7 12 2 1 11 2 11 12 2 9 1 9 2
31 10 9 0 13 3 1 10 9 11 2 11 11 11 11 11 11 2 2 16 13 13 9 1 9 0 0 1 10 9 11 2
27 1 9 1 10 9 0 2 10 9 1 10 9 15 13 0 9 1 9 2 15 15 15 13 1 10 9 2
57 11 13 10 9 1 9 1 10 9 1 10 11 11 2 15 9 0 2 1 13 10 9 1 10 9 13 1 10 9 0 1 10 11 11 2 1 11 1 10 11 2 10 12 1 11 2 9 0 1 10 9 2 13 1 10 11 2
64 10 12 1 11 1 12 2 11 12 13 1 11 2 13 10 12 1 11 1 10 0 9 2 7 16 10 9 10 9 11 15 13 1 11 1 9 2 1 10 9 0 2 13 1 10 11 1 11 2 1 10 15 13 1 10 9 1 9 1 16 11 15 13 2
19 3 15 13 1 15 1 10 9 7 4 1 13 15 10 12 9 15 13 2
28 1 10 9 2 1 10 9 1 11 2 13 16 15 4 13 2 1 10 9 7 10 9 16 13 3 10 9 2
24 15 13 1 15 15 13 3 10 9 1 11 2 13 10 9 11 1 9 10 11 2 11 2 2
14 13 0 2 7 10 9 3 0 7 15 1 11 11 2
43 15 1 10 0 9 1 9 0 2 13 1 10 11 2 16 13 10 16 15 13 9 1 9 1 0 9 1 3 13 10 9 1 10 9 1 9 0 1 10 9 1 9 2
16 13 16 13 1 10 9 16 13 16 15 13 3 1 15 13 2
21 3 10 0 9 1 11 2 3 10 9 13 9 3 1 1 10 9 1 9 0 2
26 10 9 1 10 9 0 1 11 4 13 7 13 1 9 7 10 9 15 13 1 9 0 1 10 9 2
14 13 0 10 9 1 10 11 11 12 11 11 1 11 2
22 10 9 1 10 9 13 3 0 1 10 9 1 9 2 1 9 0 1 3 3 0 2
23 13 1 10 9 1 16 10 9 0 4 4 13 2 16 1 10 9 4 13 1 10 11 2
18 10 9 4 13 10 10 9 7 10 9 0 4 13 12 9 1 9 2
19 10 9 15 13 1 9 0 2 7 10 9 13 10 9 1 10 9 12 2
17 13 1 9 13 3 10 9 7 4 13 16 13 1 10 0 9 2
12 1 9 0 12 2 3 13 0 1 0 9 2
32 10 9 15 13 1 12 9 2 10 0 9 1 10 9 0 10 11 2 7 10 9 3 13 9 0 1 10 9 7 10 9 2
27 2 3 13 10 9 16 13 10 9 1 10 9 7 10 9 7 10 9 15 13 1 9 2 2 13 11 2
48 10 9 1 10 9 1 11 1 10 9 0 0 1 10 11 13 13 10 9 0 2 1 10 9 16 15 13 10 12 9 1 10 9 1 10 12 1 11 2 1 10 9 0 7 1 9 0 2
37 10 9 0 1 10 11 1 11 1 10 11 1 10 11 11 2 11 2 2 11 11 2 13 3 16 10 9 13 1 10 9 1 11 11 1 11 2
40 11 11 13 9 1 11 11 2 10 0 9 0 2 1 9 1 10 15 15 15 13 10 9 1 10 9 1 11 7 1 10 9 1 9 0 1 10 0 9 2
18 1 12 13 10 11 11 1 11 1 10 11 2 16 13 10 0 9 2
86 7 10 9 1 11 15 13 0 9 1 10 9 1 9 7 13 1 0 10 9 2 15 16 13 1 10 9 1 10 9 1 9 2 10 2 9 2 2 9 2 7 10 9 1 9 1 9 1 9 0 7 0 2 16 1 10 3 4 13 3 1 10 9 0 3 13 1 10 9 0 1 10 9 2 7 1 10 9 1 10 9 2 1 4 13 2
37 10 9 7 10 9 13 1 11 7 11 1 9 2 7 15 15 13 16 15 13 2 7 15 2 1 13 10 9 2 15 13 9 13 7 15 13 2
24 3 1 13 10 9 15 13 1 11 2 13 15 1 9 1 12 1 10 9 2 10 9 2 2
18 13 10 9 0 7 0 2 9 16 15 13 0 8 10 9 1 9 2
19 1 10 9 2 1 9 2 15 13 1 10 9 11 16 13 9 1 11 2
20 13 3 0 1 10 9 1 11 11 2 16 10 9 13 1 9 10 9 0 2
46 10 11 1 11 13 10 13 0 10 12 1 11 1 12 2 1 11 12 1 11 7 11 12 1 11 2 3 1 16 13 9 1 10 11 1 10 11 1 11 10 12 1 11 1 12 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
23 1 12 2 1 10 9 1 10 9 1 11 1 10 9 0 2 4 13 9 1 10 9 2
21 10 9 0 1 10 9 0 4 1 13 1 7 15 13 1 10 9 1 10 9 2
15 10 12 4 13 1 9 1 10 9 11 11 12 1 12 2
55 10 9 11 13 3 0 13 10 9 1 10 9 7 1 10 9 1 9 1 10 9 2 13 10 9 1 13 10 10 9 1 10 11 11 2 13 10 9 3 0 7 13 9 0 1 10 0 9 0 15 15 0 4 13 2
31 1 11 2 10 0 9 0 13 1 9 12 9 13 10 9 1 10 9 1 10 9 7 2 3 2 1 10 9 3 0 2
23 11 13 10 0 9 1 10 9 15 3 4 8 2 13 1 10 9 7 9 11 11 11 2
32 1 10 11 11 11 2 10 9 1 10 11 15 13 1 9 1 10 9 11 11 2 13 1 10 9 10 12 1 11 1 12 2
15 4 13 12 9 1 9 2 15 1 15 13 1 10 9 2
25 1 10 12 2 12 13 12 9 1 12 9 2 7 1 10 12 2 12 13 12 9 1 12 9 2
11 11 13 10 9 1 9 0 13 1 12 2
24 10 9 13 10 9 1 15 15 13 3 3 1 10 9 2 7 3 1 10 9 7 10 9 2
37 10 9 1 9 1 10 9 0 7 10 9 0 13 10 9 1 10 10 11 11 1 11 2 11 1 10 9 1 9 2 11 11 11 2 1 12 2
13 10 9 1 9 13 1 12 9 2 2 5 5 2
14 10 0 9 1 10 9 13 1 11 11 11 1 12 2
35 10 11 1 11 11 13 10 9 0 13 1 10 9 1 11 11 2 11 2 3 1 10 9 1 11 11 2 13 10 9 1 10 9 11 2
53 1 9 2 1 9 1 0 9 1 13 9 1 0 9 2 11 2 2 9 0 2 2 1 9 0 2 15 13 16 10 9 1 9 0 1 11 2 9 0 2 13 1 10 9 1 11 11 1 3 13 12 9 2
27 3 0 2 10 2 0 2 9 1 10 9 2 10 11 7 10 11 15 13 1 9 1 10 9 1 12 2
27 1 9 10 0 9 1 9 2 15 11 13 3 2 4 3 4 13 10 9 16 4 4 13 1 10 11 2
20 13 12 9 3 3 7 13 10 9 10 9 1 9 2 1 0 11 1 9 2
20 10 9 4 13 1 12 2 7 1 10 9 3 4 13 1 9 0 1 11 2
16 4 13 9 2 16 10 10 9 13 10 9 1 10 9 2 2
34 10 9 1 9 0 7 10 9 13 1 9 13 4 13 1 10 9 1 10 9 2 13 9 1 9 2 9 1 11 7 9 1 9 2
5 10 9 13 0 2
28 11 11 2 10 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 2 9 7 9 1 9 0 0 2
30 13 1 10 9 1 12 9 1 9 1 11 2 10 9 1 9 2 7 1 12 9 1 11 2 9 1 10 11 11 2
17 11 15 13 2 13 16 4 13 0 2 1 3 13 15 13 2 2
33 10 9 11 2 11 1 10 9 1 9 1 10 9 9 13 10 9 0 16 13 1 10 9 11 7 15 13 10 9 1 12 5 2
33 10 9 1 0 9 13 10 9 1 10 9 1 10 0 9 2 0 2 16 10 9 1 10 9 13 10 9 1 9 1 10 9 2
6 13 10 11 1 11 2
27 13 2 1 9 1 9 2 10 9 0 1 2 11 11 2 2 1 10 0 9 1 10 11 7 10 9 2
28 3 2 11 3 13 16 3 15 13 10 9 0 2 13 13 2 15 13 1 9 1 10 9 1 10 9 2 2
20 10 9 1 9 3 13 0 2 7 13 0 13 10 9 1 3 1 12 9 2
28 1 9 2 10 9 3 7 3 13 1 13 2 16 10 9 13 1 3 0 9 7 3 13 10 9 1 13 2
27 1 10 9 0 2 1 9 2 15 13 1 10 9 1 11 1 10 9 1 10 9 1 10 9 1 9 2
16 10 9 1 9 15 13 3 3 16 15 4 13 10 9 0 2
22 1 10 11 1 10 11 11 10 9 13 10 9 1 9 1 10 12 7 10 12 9 2
21 1 9 2 11 15 13 1 10 9 7 13 13 1 9 3 1 10 9 1 9 2
35 10 9 2 1 9 1 10 11 11 1 10 11 11 2 11 2 2 13 1 10 9 2 1 9 16 15 13 13 1 10 0 9 1 9 2
15 10 9 11 13 1 10 9 8 8 2 9 1 9 2 2
13 13 3 0 16 15 13 1 10 9 1 10 9 2
60 13 13 16 1 10 9 1 9 2 15 13 10 9 1 10 9 2 11 2 2 1 10 9 0 11 11 11 11 2 15 13 10 9 1 10 9 0 2 13 3 1 10 9 1 10 9 3 0 1 9 1 10 9 0 1 10 9 1 12 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
32 10 9 1 10 9 8 1 10 2 9 2 10 11 2 10 11 7 11 13 10 0 9 2 10 9 1 10 11 2 1 11 2
29 10 0 9 0 1 10 11 1 10 11 1 10 9 13 10 9 0 1 11 11 11 2 2 11 11 11 11 2 2
23 10 9 13 3 10 9 1 10 9 11 11 11 2 7 10 9 1 10 9 11 11 11 2
20 16 15 13 16 13 9 16 13 9 2 11 1 9 13 10 9 1 10 9 2
28 2 10 11 2 13 1 10 11 11 2 1 10 16 13 1 11 2 1 10 9 16 13 10 12 9 1 9 2
18 4 13 1 10 9 0 11 11 1 12 2 1 10 9 1 11 11 2
28 10 9 2 11 13 1 11 7 1 9 1 10 9 2 13 10 0 9 16 15 13 1 15 1 10 9 0 2
40 13 2 0 1 10 9 1 11 1 11 11 7 10 9 1 11 11 2 1 15 1 10 0 9 0 1 10 10 9 2 7 10 9 0 1 10 9 1 9 2
12 9 10 11 2 1 11 11 2 9 1 11 2
20 3 13 15 3 1 10 9 1 11 0 2 7 9 16 4 1 13 0 9 2
34 10 0 9 1 10 11 2 12 13 10 12 1 11 1 12 2 7 10 0 9 1 10 9 0 13 10 12 1 11 1 10 0 9 2
8 3 15 13 1 9 1 9 2
13 15 13 0 1 10 9 10 9 16 13 1 11 2
24 10 9 11 13 10 9 1 10 9 1 9 1 11 2 7 13 9 1 10 9 12 7 12 2
43 11 11 2 12 1 11 1 12 2 2 13 10 9 0 2 15 13 1 9 7 3 13 1 10 11 12 2 1 10 0 9 1 11 11 2 11 13 10 9 1 9 0 2
28 10 9 1 16 10 9 1 10 9 13 10 9 0 11 11 15 13 10 9 1 1 3 13 13 10 9 2 2
30 10 9 4 4 13 1 10 9 1 10 9 3 0 2 15 16 13 10 9 1 9 1 10 9 1 9 1 10 9 2
40 10 9 13 3 0 1 9 1 16 1 9 1 12 15 13 10 9 1 9 2 15 16 13 1 10 9 13 9 0 1 10 9 1 9 1 9 1 10 9 2
42 10 9 0 4 13 1 10 9 1 9 1 9 1 10 9 16 15 13 1 9 1 11 1 12 1 11 1 12 7 13 10 9 3 13 10 9 3 15 13 10 9 2
24 1 10 9 1 9 10 9 0 13 10 9 0 1 10 9 0 1 10 9 0 1 10 9 2
47 1 10 9 2 10 9 1 11 11 1 10 9 2 11 11 11 13 10 9 1 10 9 16 10 9 15 13 1 13 10 11 1 11 1 12 7 10 12 9 1 10 9 1 10 9 0 2
19 13 10 9 1 10 11 11 11 11 11 11 11 2 1 9 1 12 9 2
11 10 9 1 11 15 13 13 1 10 9 2
18 2 3 15 13 16 15 13 1 10 9 1 10 9 0 2 2 13 2
17 1 9 2 10 9 16 13 10 9 3 15 13 10 9 15 13 2
83 10 0 9 1 10 9 1 10 9 13 1 10 9 0 16 3 15 13 1 10 9 0 1 10 9 7 3 1 10 9 2 10 9 7 9 1 10 9 0 3 13 9 1 10 9 8 1 10 9 7 13 10 9 0 1 9 2 1 10 9 3 0 13 9 16 13 0 9 0 1 10 9 0 1 9 16 13 13 10 9 1 9 2
24 10 9 13 0 1 10 9 1 11 7 15 13 1 9 0 3 1 9 3 13 10 0 9 2
22 13 9 0 13 1 9 1 10 15 15 4 13 9 0 2 1 9 7 1 9 0 2
11 11 11 13 13 2 7 13 10 0 9 2
8 13 3 1 12 9 1 13 2
36 1 10 9 2 11 13 13 10 9 1 10 9 2 16 4 1 13 1 10 9 1 10 3 13 9 1 10 9 11 11 2 1 9 1 9 2
17 1 12 2 1 10 9 0 1 11 2 13 1 10 9 1 9 2
14 3 15 13 9 0 1 3 10 10 9 1 10 9 2
16 15 13 1 10 9 1 11 2 11 2 11 2 11 7 11 2
57 1 10 9 1 10 11 10 9 16 15 13 1 3 9 13 15 1 2 11 2 11 2 1 12 9 7 13 10 9 15 10 9 12 9 13 1 10 0 9 2 15 13 15 1 2 11 2 11 7 11 2 11 2 1 12 9 2
46 3 3 2 12 1 11 1 12 2 4 13 9 0 1 10 11 11 1 11 2 0 9 1 10 15 13 12 7 12 9 2 1 10 9 3 12 13 9 1 10 9 1 11 7 11 2
30 10 9 16 10 9 3 13 9 13 9 1 9 1 9 1 0 9 2 15 3 13 9 1 10 9 0 1 10 9 2
25 10 9 13 1 10 12 9 2 9 1 10 16 10 9 1 10 9 0 13 10 9 1 10 9 2
45 1 10 0 9 0 2 12 2 2 10 9 0 1 0 9 0 1 11 2 13 10 9 1 1 12 7 12 9 2 13 10 9 1 11 11 10 16 13 10 9 3 0 1 9 0
15 13 10 9 1 10 9 1 10 9 7 11 4 13 9 2
13 10 11 11 15 13 0 3 1 10 9 0 0 2
11 11 13 10 9 1 3 9 13 1 9 2
72 9 0 11 11 13 2 1 3 1 10 9 2 10 11 11 11 2 10 11 11 1 11 11 1 9 2 1 10 11 2 8 2 2 9 1 9 2 10 11 1 10 11 9 2 10 11 11 11 9 1 9 2 10 11 1 11 2 10 11 11 2 7 1 10 9 7 10 11 1 11 9 2
39 10 9 13 1 10 11 11 0 2 13 3 2 1 9 7 13 10 9 0 1 9 0 7 10 9 0 1 10 9 2 15 16 3 13 1 11 7 11 2
15 10 9 0 2 0 7 0 13 1 10 9 1 0 9 2
48 15 3 4 13 2 1 9 2 1 12 9 10 9 1 11 9 7 13 3 0 7 0 1 15 7 10 9 16 15 13 2 15 9 7 9 2 10 0 9 3 3 15 4 1 13 1 15 2
11 1 10 9 1 9 1 11 13 12 9 2
30 15 13 10 9 1 10 9 1 11 11 2 16 13 1 10 0 11 11 11 13 10 9 1 13 10 9 1 11 11 2
17 11 11 11 2 11 2 12 2 12 2 13 10 9 7 9 0 2
18 3 13 10 9 12 1 10 11 11 1 11 10 12 1 11 1 12 2
22 16 3 13 10 9 0 1 10 9 2 10 11 4 13 9 0 1 9 0 7 0 2
23 10 9 9 11 11 11 11 7 10 9 11 11 1 11 11 11 2 12 9 1 11 11 2
15 10 9 3 13 3 0 7 1 0 10 9 3 13 0 2
22 11 2 10 9 0 11 11 13 10 11 16 10 9 11 11 13 0 1 10 0 9 2
34 1 13 2 10 9 1 10 9 13 3 0 2 1 10 0 9 0 10 9 1 10 9 0 15 13 1 10 12 5 7 10 12 5 2
11 10 9 16 13 15 13 9 1 13 15 2
38 0 7 3 2 13 0 16 10 9 4 13 3 0 7 0 7 3 15 13 1 9 2 7 15 16 3 4 1 13 13 16 3 13 2 7 15 2 2
8 13 3 1 10 9 1 11 2
32 7 13 10 9 1 9 2 13 1 13 1 9 1 9 7 9 1 10 11 11 2 15 16 13 3 10 9 4 13 10 9 2
13 10 9 1 10 9 13 0 7 10 9 13 0 2
13 3 13 12 9 2 1 10 15 12 13 3 0 2
14 13 9 1 10 9 0 2 7 3 13 10 9 0 2
10 13 10 9 9 13 10 9 1 9 2
19 1 10 9 13 10 11 11 1 4 13 15 1 9 7 1 9 1 11 2
36 11 2 11 2 11 13 10 9 7 9 0 2 1 10 9 1 11 2 11 2 9 1 9 2 1 10 9 1 11 7 9 1 11 2 11 2
11 15 4 13 10 3 0 9 1 10 9 2
10 15 13 10 0 9 1 9 7 9 2
45 1 12 2 12 13 10 9 1 11 13 1 10 9 7 1 10 9 12 2 12 2 12 2 12 7 12 2 12 13 9 1 10 11 11 1 11 1 9 1 10 9 11 1 11 2
24 10 9 13 13 10 9 0 1 10 9 1 9 1 10 11 9 7 9 2 8 7 8 2 2
14 10 9 7 10 9 1 10 9 9 4 13 1 12 2
49 10 9 0 2 1 9 13 16 10 9 13 10 9 3 15 4 13 10 9 2 13 10 9 3 0 2 1 10 9 16 4 7 13 8 10 15 15 13 15 2 10 9 13 16 4 13 10 9 2
14 10 9 13 3 10 0 9 7 10 9 1 10 9 2
29 11 3 4 13 1 13 1 11 7 3 16 13 9 2 16 15 13 1 11 7 3 1 10 9 1 1 10 11 2
26 11 11 11 11 2 11 2 13 3 12 8 8 2 11 12 7 11 12 2 1 9 1 9 7 9 2
12 1 12 15 13 16 13 0 1 10 9 0 2
14 10 9 0 15 4 13 1 10 9 2 9 7 9 2
25 11 13 0 1 13 10 9 1 10 12 1 11 1 12 2 1 10 9 10 9 4 13 1 11 2
30 1 10 0 9 13 1 9 1 10 9 7 9 11 1 11 2 16 13 1 10 0 9 13 10 12 1 11 1 12 2
35 10 9 13 10 9 1 11 2 1 10 15 2 1 10 9 2 10 9 11 1 9 1 10 9 0 13 1 10 9 0 1 10 9 0 2
13 10 12 1 11 1 12 13 10 9 1 8 9 2
43 1 9 1 16 10 11 1 11 13 10 9 7 10 9 2 10 9 0 9 3 15 13 2 2 1 15 15 3 3 15 4 13 10 9 1 10 9 2 2 13 10 9 2
19 10 12 1 11 1 12 15 13 1 11 10 12 9 1 10 9 1 9 2
11 13 1 11 1 9 7 13 0 1 15 2
21 10 11 15 13 1 10 12 9 3 0 1 10 9 2 11 11 2 11 7 11 2
21 4 13 9 1 10 11 1 10 11 1 11 1 10 11 11 1 11 2 11 2 2
40 11 11 2 11 3 15 13 1 10 9 1 10 9 0 11 11 2 11 11 2 11 11 11 11 2 2 12 2 2 16 15 13 1 10 9 3 0 7 9 2
25 10 9 13 10 15 3 0 1 15 2 9 2 1 13 1 11 2 7 1 10 9 15 13 0 2
29 3 4 13 1 0 9 1 9 0 7 9 16 13 1 10 9 12 7 16 13 10 9 1 0 9 1 10 9 2
42 2 10 9 3 0 13 10 9 1 10 9 1 10 9 0 16 4 13 1 10 9 2 2 13 11 11 2 9 0 1 10 9 1 11 11 2 1 10 16 13 11 2
8 3 13 10 9 1 9 9 2
25 13 10 9 1 12 9 7 1 9 10 9 3 15 4 13 16 15 13 13 10 9 1 10 9 2
52 1 11 13 1 10 9 15 11 2 12 2 1 10 0 11 11 7 1 15 11 11 2 12 2 2 1 11 11 7 11 11 2 3 13 10 9 1 10 9 0 7 1 10 9 2 1 10 9 1 10 9 2
17 1 0 9 2 1 12 10 9 0 13 12 5 1 10 9 0 2
4 13 1 11 2
20 15 13 1 0 9 2 7 13 10 9 7 0 9 1 10 9 1 9 0 2
22 10 0 9 1 10 9 1 9 15 13 1 11 1 10 12 1 10 9 0 0 11 2
49 8 8 8 8 8 8 8 2 8 2 2 2 2 1 9 2 2 1 10 9 1 10 9 13 3 2 2 2 13 10 0 9 1 9 1 10 9 0 11 11 2 13 10 12 1 11 1 12 2
13 13 9 0 2 10 9 1 11 3 15 13 15 2
15 1 10 9 1 11 13 1 10 9 1 11 7 11 11 2
17 10 9 2 3 13 1 10 9 1 11 2 13 10 0 9 0 2
28 3 13 9 1 10 11 11 11 2 1 10 9 1 10 9 1 11 2 11 7 9 1 11 1 10 11 11 2
61 13 10 9 1 10 9 1 9 1 10 9 2 9 1 10 15 4 13 10 9 0 2 11 2 9 1 11 11 2 9 1 11 11 2 2 3 1 13 10 9 1 9 0 2 0 1 15 16 15 13 1 10 0 9 0 2 13 1 10 9 2
5 15 13 1 11 2
54 15 4 13 16 11 11 2 11 2 13 10 9 1 10 3 0 12 9 1 9 2 16 11 11 2 11 2 7 11 11 2 11 2 15 13 10 12 0 9 7 16 11 11 2 10 11 2 15 13 10 0 12 9 2
46 7 13 16 10 9 4 13 1 10 9 2 11 2 9 0 2 9 0 2 13 10 9 15 13 3 9 2 9 7 10 0 9 1 9 0 1 9 1 15 15 13 10 9 1 8 2
10 11 11 4 13 10 9 1 10 9 2
28 10 9 13 0 1 10 9 1 9 16 13 10 11 2 0 9 3 10 11 11 11 4 7 13 10 9 8 2
67 3 16 11 13 1 15 16 2 15 13 13 9 1 10 10 9 1 10 9 2 2 13 10 0 9 1 10 9 2 15 13 3 16 1 10 9 1 10 11 1 11 2 13 16 15 1 10 9 3 15 13 2 2 2 13 16 11 4 1 13 15 1 9 7 3 2 2
25 1 12 13 1 9 1 10 9 1 10 9 1 11 2 7 1 12 1 12 2 1 15 1 11 2
38 10 9 2 10 11 11 12 2 3 3 13 1 10 9 1 11 11 2 13 13 10 9 1 11 1 10 9 1 10 9 0 7 13 10 0 9 0 2
40 10 12 1 11 1 12 2 1 10 9 1 9 2 11 13 1 10 9 10 9 1 11 11 1 10 11 2 16 13 1 10 0 9 10 9 1 10 9 0 2
17 13 10 9 1 11 10 9 1 9 1 10 15 13 9 1 11 2
41 11 4 0 7 13 13 1 10 9 1 9 1 10 11 11 11 1 11 2 11 2 3 9 1 11 2 11 2 2 7 10 11 11 11 1 11 11 2 11 2 2
17 13 1 9 1 9 7 9 0 16 13 10 9 1 10 9 0 2
50 10 9 1 11 13 9 0 2 15 16 15 13 1 10 9 0 1 10 9 0 1 9 16 15 13 1 10 9 7 15 16 13 1 15 10 9 15 13 1 10 9 0 1 10 9 1 9 1 11 2
33 1 0 2 10 9 1 10 10 9 0 13 10 12 9 1 9 2 13 1 3 1 12 9 1 9 7 3 1 12 9 1 9 2
20 15 13 1 10 9 1 10 11 11 1 10 9 2 3 13 10 9 1 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
34 1 10 9 1 12 13 1 10 9 1 11 2 15 13 1 2 7 1 12 7 12 13 3 1 9 1 10 9 1 11 2 11 2 2
27 13 10 9 13 15 16 13 15 2 3 7 13 1 3 2 10 0 9 1 15 16 4 13 1 10 9 8
37 10 9 8 2 0 11 11 4 13 3 10 9 1 9 1 10 11 11 2 1 10 16 13 9 1 10 9 1 10 0 9 2 13 10 9 0 2
35 15 13 1 10 9 7 9 0 7 13 10 9 2 1 16 4 1 13 0 9 1 9 2 1 10 3 0 7 3 0 2 15 4 13 2
21 1 11 2 10 9 13 1 10 0 9 0 7 15 13 10 9 13 1 10 11 2
17 1 10 9 4 13 10 0 9 0 2 10 0 11 1 10 11 2
33 11 7 11 13 1 9 16 13 10 11 1 10 8 1 11 2 11 2 13 10 9 3 13 16 13 10 9 1 9 1 10 9 2
11 10 9 13 10 0 9 15 13 10 9 2
34 11 2 1 10 16 10 9 13 1 9 0 1 10 9 2 13 12 9 1 9 1 10 9 1 9 1 10 12 9 13 1 10 9 2
33 1 9 1 9 2 12 9 3 0 2 1 10 9 2 13 10 9 1 10 10 9 7 13 1 10 9 2 1 9 2 9 2 2
16 3 15 13 10 9 11 11 2 3 15 13 0 9 7 9 2
6 2 3 13 10 9 2
11 15 15 13 10 9 1 10 9 1 11 2
16 10 9 4 13 1 10 9 1 9 0 0 15 4 13 3 2
42 1 12 2 15 13 16 10 9 1 10 9 1 10 9 1 9 16 13 10 9 13 1 10 9 0 10 9 1 10 9 2 10 9 7 9 7 9 0 1 10 9 2
31 11 13 1 11 12 9 1 9 2 1 9 1 15 15 11 13 3 10 9 0 1 11 2 16 3 13 1 13 3 9 2
20 10 9 3 13 16 10 9 4 4 13 1 10 9 1 10 9 1 9 0 2
37 1 10 9 1 10 9 2 11 7 10 9 2 11 2 11 7 11 2 13 10 9 1 11 13 15 15 1 11 2 15 4 13 10 9 1 11 2
40 13 10 0 7 0 9 0 1 10 9 2 13 1 9 2 9 0 2 8 9 2 9 0 7 0 9 16 13 1 10 9 3 0 1 10 11 11 7 11 2
21 10 9 1 10 0 9 13 1 9 1 10 9 2 10 9 7 10 9 1 9 2
19 15 13 1 9 2 16 13 1 10 9 0 2 10 9 7 1 10 9 2
14 10 9 0 1 10 9 13 10 9 0 7 10 9 2
13 3 2 10 0 9 13 1 10 12 9 10 9 2
28 15 3 1 12 9 1 9 7 10 9 1 9 15 4 4 7 13 10 9 2 3 7 15 13 10 9 0 2
13 10 9 13 1 10 9 1 10 9 3 3 0 2
17 10 9 13 12 9 7 10 9 0 1 10 9 13 1 11 11 2
16 3 1 10 9 1 11 2 10 9 13 3 10 9 1 11 2
4 14 9 0 2
44 10 9 15 13 10 9 11 7 11 1 10 9 1 12 9 2 13 13 15 12 9 1 10 13 15 10 9 2 12 1 10 13 1 10 9 1 10 9 2 12 1 13 15 2
33 1 9 2 1 10 11 1 10 11 10 9 1 9 4 13 1 9 1 9 16 13 1 9 0 7 9 1 9 1 9 13 9 2
27 13 3 0 1 9 1 10 9 12 2 11 4 1 13 1 10 9 1 10 9 1 11 2 3 1 11 11
45 16 15 13 10 0 9 1 9 7 9 2 13 1 10 9 1 11 11 11 2 13 1 10 9 1 13 10 9 0 1 11 2 13 9 1 10 9 1 10 9 0 1 10 9 2
34 3 13 0 1 10 9 1 9 0 10 9 1 9 0 1 13 10 9 0 2 7 13 3 9 0 1 10 9 1 9 1 9 0 2
8 9 1 10 9 2 11 11 2
33 1 10 9 1 10 9 15 13 15 1 10 0 11 7 15 1 10 9 16 13 0 1 10 9 1 10 10 9 1 10 9 0 2
40 11 11 11 13 11 1 11 7 1 11 1 10 11 1 11 2 9 1 11 7 11 1 10 11 1 11 7 1 10 11 11 1 11 2 1 10 15 3 13 9
12 4 13 1 10 9 11 11 2 1 11 11 2
34 10 13 1 10 9 0 8 2 8 2 2 9 2 2 7 8 2 8 2 2 9 2 2 2 13 9 1 10 9 16 13 10 9 2
24 1 10 12 9 16 13 3 2 3 13 9 0 3 16 15 13 9 1 10 9 1 10 9 2
7 4 13 1 10 9 12 2
13 2 1 11 11 4 13 3 7 13 1 13 9 2
37 10 9 1 9 0 1 11 13 10 12 1 12 1 11 9 1 10 0 9 1 12 2 3 7 10 9 0 1 10 9 13 1 10 12 1 12 2
18 10 9 13 10 9 0 1 9 12 9 1 10 9 12 1 10 9 2
11 10 10 9 13 1 9 0 2 11 12 2
23 1 10 9 2 10 9 13 1 9 1 11 11 2 8 2 2 9 1 10 9 11 12 2
17 3 2 15 13 1 10 9 16 15 15 13 1 11 1 10 9 2
39 10 9 1 10 12 13 10 9 1 10 0 9 1 9 16 13 1 13 1 10 9 12 1 10 9 1 10 11 1 15 1 10 9 1 10 9 0 0 2
24 13 9 0 1 10 11 1 11 7 9 0 1 10 0 9 1 9 7 1 10 11 11 11 2
20 15 13 1 12 7 12 7 13 10 10 9 1 10 9 0 1 10 9 0 2
21 13 10 0 7 0 9 1 10 0 9 13 11 11 16 15 13 9 7 3 9 2
46 1 11 1 12 13 9 1 11 1 11 11 1 13 1 10 9 1 10 15 13 2 11 11 2 16 13 1 10 9 1 13 1 10 0 9 2 3 1 13 1 0 9 1 10 9 2
32 13 0 10 9 1 9 7 9 1 10 11 12 9 1 10 0 9 0 2 10 11 12 2 16 13 12 8 7 13 9 0 2
19 11 11 4 13 1 11 11 7 13 1 11 11 12 2 1 10 9 12 2
19 10 9 1 10 10 9 1 0 9 1 10 9 0 13 10 0 9 0 2
20 10 9 13 0 2 1 12 5 1 0 2 7 0 7 13 10 0 9 0 2
35 13 10 9 0 1 11 16 13 9 0 1 11 2 11 7 9 0 0 1 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
11 10 9 1 10 9 13 1 11 2 11 2
26 10 9 1 3 3 1 12 9 1 10 0 9 3 3 1 0 9 1 9 1 10 0 9 1 9 2
22 11 11 8 12 2 13 10 9 1 9 0 7 0 0 1 10 9 7 9 1 11 2
66 1 10 9 0 2 7 1 3 1 15 2 15 13 1 10 9 1 10 9 16 2 13 1 10 9 0 2 13 10 9 1 10 9 1 10 9 0 1 16 10 9 1 9 1 10 9 13 1 13 10 9 1 9 2 13 1 10 9 0 2 7 4 13 1 15 2
17 10 9 0 3 13 16 3 13 3 9 7 13 15 1 10 9 2
9 0 9 1 13 10 9 1 9 2
42 1 13 10 9 1 10 11 1 10 11 7 10 11 1 10 9 13 1 13 10 9 1 10 9 0 3 1 10 9 7 15 13 1 9 16 13 10 9 1 10 11 2
17 11 11 13 10 9 1 10 9 1 11 2 1 10 9 1 11 2
56 1 10 9 1 12 2 11 13 10 9 1 10 15 10 12 5 13 0 2 12 5 9 2 12 5 0 2 12 5 0 2 12 5 9 1 10 11 2 10 12 5 1 10 9 2 7 10 12 5 13 1 12 7 3 9 2
25 10 9 0 1 12 2 1 12 1 11 2 13 10 9 0 1 10 12 9 2 0 1 10 9 2
13 2 10 9 4 13 13 10 12 9 1 9 0 2
9 3 15 13 1 10 9 1 9 2
21 1 10 9 13 1 10 9 15 13 16 15 2 13 7 13 2 10 0 9 0 2
49 13 10 0 9 1 9 0 7 0 2 9 7 9 2 15 3 0 2 15 9 16 13 15 0 2 15 13 10 8 1 10 0 9 7 13 0 2 9 0 7 10 9 8 0 2 0 12 8 2
35 16 3 10 9 10 9 1 11 11 13 10 0 8 0 1 10 0 9 2 4 13 13 10 9 10 9 1 11 1 9 1 10 0 9 2
14 2 13 16 3 4 1 13 16 13 1 10 9 0 2
17 7 1 10 9 12 13 1 9 1 10 11 11 1 10 9 0 2
34 11 1 11 2 11 2 11 11 2 13 10 12 1 11 1 12 2 11 2 13 10 12 1 11 1 12 2 2 9 1 10 9 0 2
11 1 13 1 9 7 1 9 15 13 15 2
54 1 12 15 13 1 11 11 7 1 10 9 8 2 0 2 3 1 10 9 1 11 2 13 1 11 7 3 1 11 2 3 13 1 13 9 13 1 10 9 0 2 10 9 1 10 9 15 13 10 9 1 9 0 2
20 13 1 9 10 9 3 0 1 11 2 13 1 10 9 0 1 10 9 0 2
29 1 3 4 13 1 0 9 3 13 1 9 13 1 16 10 9 13 0 2 16 13 0 16 11 11 13 10 9 2
22 15 13 13 10 9 3 1 13 10 9 1 10 9 7 13 15 1 16 4 4 13 2
20 1 10 9 2 11 13 10 9 1 10 9 1 10 9 1 10 9 1 11 2
29 13 1 10 9 2 1 10 9 16 10 9 1 10 9 1 11 2 1 3 13 10 9 2 1 9 1 12 9 2
26 10 9 1 0 13 15 0 2 1 9 1 16 10 9 1 10 9 2 10 9 1 9 2 13 0 2
35 10 9 11 11 13 10 0 9 1 10 15 13 16 10 9 13 2 10 9 0 2 7 1 10 15 10 9 13 1 3 9 7 10 9 2
47 10 9 12 1 11 1 12 10 9 1 11 11 2 1 10 3 1 10 12 1 10 9 1 11 2 13 1 10 9 2 7 4 1 13 15 9 16 13 2 11 11 13 3 1 9 2 2
41 3 2 10 9 13 1 9 1 10 11 1 11 2 1 12 1 12 2 13 15 1 9 0 1 0 9 2 1 10 9 1 10 2 11 1 10 11 11 11 2 2
17 10 9 1 9 1 12 9 1 9 4 4 13 3 3 7 3 2
38 2 10 9 1 10 9 16 4 13 10 9 3 13 3 0 7 13 2 13 11 2 16 13 10 9 0 16 13 10 0 9 1 10 9 1 10 9 2
18 10 9 13 10 9 0 1 9 12 9 1 10 9 12 1 10 9 2
28 1 10 9 2 10 9 3 0 7 0 2 11 2 4 13 10 0 9 2 7 10 9 3 15 4 13 13 2
23 10 11 13 1 12 9 0 1 10 9 2 10 11 11 7 11 7 10 9 1 10 11 2
26 10 9 1 10 9 2 11 2 13 10 9 1 9 1 11 7 13 9 1 10 9 2 10 9 11 2
39 11 13 16 10 9 0 4 13 0 9 1 11 10 12 1 11 1 10 16 13 9 1 13 0 9 16 13 15 1 9 7 9 1 10 9 7 10 9 2
28 10 9 0 0 13 10 9 0 1 10 9 0 1 10 9 2 10 9 1 9 7 10 9 0 1 9 0 2
31 10 12 0 1 10 9 13 1 10 9 0 7 10 12 9 1 10 11 13 1 10 9 1 10 9 7 15 10 9 0 2
39 13 2 1 9 2 16 10 9 13 9 7 9 0 16 13 16 2 13 1 16 10 9 1 10 9 0 1 9 1 10 9 0 4 13 1 10 9 2 2
17 10 9 13 10 9 0 13 1 12 9 13 1 9 1 0 9 2
16 13 10 9 0 1 11 1 10 12 1 10 9 1 12 9 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
41 11 11 2 13 1 9 1 10 9 1 12 1 11 1 12 2 13 1 11 1 12 13 10 9 1 10 9 1 12 9 2 13 10 9 1 10 9 1 10 9 2
38 11 11 4 13 1 12 1 10 11 11 11 1 2 0 11 1 10 9 1 9 0 1 10 0 9 2 1 10 9 1 11 11 1 11 2 12 2 2
40 10 9 0 13 1 10 12 5 1 11 7 11 2 7 10 12 5 1 10 9 1 12 2 16 11 11 13 10 0 9 1 9 1 9 1 10 11 11 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
28 1 10 9 1 10 9 0 2 1 10 9 1 9 13 3 1 12 10 9 16 10 9 13 1 10 9 0 2
36 1 10 9 2 13 1 15 11 11 1 10 11 11 11 11 11 2 11 2 1 12 9 2 13 1 10 9 1 12 9 0 1 12 7 12 2
16 13 1 10 9 0 1 10 9 2 13 10 9 1 9 0 2
20 9 1 10 0 9 7 3 3 9 0 1 11 1 10 9 1 11 1 12 2
26 10 11 2 12 11 13 10 0 9 1 11 11 11 2 11 2 13 1 10 11 11 1 10 11 11 2
10 15 13 10 9 2 9 2 9 2 8
22 7 1 10 9 2 10 9 13 3 0 7 1 9 1 10 9 0 2 3 13 9 2
29 10 9 7 9 1 10 11 1 11 12 13 1 10 9 1 9 1 5 1 10 12 9 1 10 11 12 1 11 2
37 11 13 16 13 13 10 9 0 1 10 9 1 10 9 7 1 15 13 0 9 1 9 1 10 9 16 15 4 13 1 10 9 1 10 9 0 2
20 15 13 16 4 13 1 9 1 10 9 11 1 15 0 15 13 10 9 0 2
61 1 10 9 2 1 9 1 10 9 0 16 13 11 2 7 10 9 16 13 9 1 11 2 11 13 9 1 10 9 1 10 9 0 2 7 10 9 7 10 9 0 4 9 1 10 0 9 1 10 9 2 7 10 9 13 1 9 1 13 15 2
10 11 11 15 13 1 0 2 7 0 2
15 10 9 0 3 13 13 1 10 9 1 10 9 1 11 2
22 11 13 10 9 1 9 0 0 13 1 10 12 16 15 13 0 1 10 11 11 11 2
44 1 9 1 10 9 2 3 13 1 10 0 9 1 9 9 2 16 13 10 9 1 10 9 16 11 4 13 1 9 1 11 2 15 15 13 10 9 1 16 15 15 13 9 2
23 1 12 2 11 11 7 11 11 13 16 10 9 0 1 10 9 1 10 9 4 13 9 2
40 1 10 9 1 9 8 2 10 9 1 10 9 1 10 9 4 13 10 9 1 10 11 2 11 2 7 2 1 10 9 2 13 9 1 9 7 1 9 0 2
27 10 11 11 4 13 1 10 9 2 11 11 11 11 2 1 10 12 5 11 8 11 11 7 13 1 11 2
10 13 0 9 1 10 9 1 9 0 2
25 1 9 2 10 9 1 9 4 4 13 1 10 9 1 9 2 7 15 13 9 0 1 9 0 2
31 1 12 2 1 10 9 2 11 11 2 10 9 1 11 2 13 15 1 11 2 13 1 10 9 1 9 1 9 1 9 2
16 10 9 1 9 13 0 2 3 16 4 1 13 15 1 9 2
41 10 9 0 3 15 4 13 1 10 9 3 1 11 2 3 7 13 1 10 9 0 1 13 9 1 10 9 0 10 0 4 13 1 11 2 10 9 11 15 13 2
40 10 9 1 10 9 0 1 10 9 1 11 13 16 10 9 0 1 10 9 11 4 13 10 0 9 1 13 15 1 13 1 10 9 1 9 0 1 10 9 2
37 11 12 13 10 0 9 1 10 0 9 2 1 10 15 13 2 9 0 2 7 1 15 13 1 11 11 2 1 10 9 1 10 11 11 1 11 2
22 10 9 15 13 1 16 10 9 1 10 9 4 13 15 1 9 1 13 10 10 9 2
23 1 15 9 1 10 9 11 2 10 9 1 11 13 15 1 10 9 0 13 1 10 9 2
63 11 11 2 11 2 7 11 11 13 10 9 0 13 1 10 9 12 9 12 9 1 9 9 7 12 9 12 9 1 9 9 1 12 9 1 9 2 1 10 9 1 10 11 0 1 10 9 1 10 11 2 9 1 11 2 1 10 9 1 10 9 0 2
16 13 1 11 1 10 9 3 13 10 9 1 9 1 9 0 2
31 16 10 9 3 15 13 1 10 9 1 9 1 12 9 1 11 2 10 9 15 13 1 10 9 1 10 0 9 1 9 2
23 13 10 9 16 4 13 3 1 9 10 9 0 1 10 9 0 1 10 9 1 10 9 2
66 10 9 4 4 13 1 10 9 11 11 7 11 11 2 16 3 4 13 1 10 9 0 7 0 13 1 10 9 0 16 15 13 1 11 1 10 9 2 7 16 13 1 13 1 13 15 1 10 0 9 1 10 9 9 0 7 15 1 10 0 9 0 1 11 11 2
57 1 10 9 13 10 9 11 11 7 11 11 2 7 7 10 9 1 10 9 2 10 9 11 11 2 10 9 11 11 11 2 10 9 11 11 7 11 11 2 10 9 11 11 7 10 9 1 9 11 11 2 13 9 1 0 9 2
13 0 1 11 11 2 13 8 2 9 1 10 9 2
15 2 13 10 9 0 1 9 7 9 1 10 9 1 11 2
8 15 9 10 9 0 7 0 2
13 10 9 1 9 13 1 12 8 2 5 5 5 2
8 13 3 7 3 4 13 9 2
51 1 10 9 4 13 1 10 9 1 10 9 2 7 3 2 7 1 9 0 2 1 15 1 10 9 0 1 0 2 13 1 10 9 1 10 9 2 13 1 13 10 9 7 13 1 10 9 1 10 9 2
24 1 10 9 0 1 11 13 0 10 13 9 0 2 13 1 9 0 1 9 13 1 9 0 2
24 1 12 13 1 11 7 13 1 10 11 1 11 11 1 11 11 3 13 9 11 7 11 11 2
45 10 9 1 10 11 11 11 2 16 13 9 10 11 1 10 9 1 3 1 12 9 1 13 2 4 13 16 13 1 9 0 16 13 10 9 1 11 1 13 10 8 1 10 11 2
70 1 16 10 9 1 11 2 13 11 2 1 10 15 3 15 13 10 9 2 4 13 1 15 16 13 9 7 1 10 9 1 11 2 9 1 16 15 4 13 10 9 2 16 3 13 0 1 10 9 2 11 3 13 9 1 10 0 9 1 4 13 15 1 10 9 3 0 16 15 2
29 1 10 9 1 15 1 12 2 11 15 13 1 10 9 1 13 1 13 1 11 2 13 16 10 9 13 10 9 2
11 11 4 13 12 5 7 11 2 12 5 2
28 11 11 13 10 9 0 2 16 3 13 0 2 11 15 4 13 10 9 3 0 16 15 13 3 0 16 13 2
20 16 13 13 15 2 11 13 3 10 9 16 13 1 10 9 2 7 13 9 2
37 11 13 10 9 1 9 2 13 1 12 9 1 11 1 10 9 12 2 12 9 0 1 10 9 1 0 7 15 13 1 10 9 11 11 1 13 2
12 11 13 8 1 10 0 9 1 10 11 11 2
26 1 11 11 13 16 10 9 13 13 1 10 9 0 3 3 2 16 10 9 13 3 1 11 1 12 2
55 3 13 10 9 16 16 15 13 10 11 11 13 16 1 10 9 11 15 16 13 13 13 15 15 13 3 9 2 13 9 16 3 15 13 2 1 11 11 12 7 13 10 9 16 10 9 2 3 13 15 1 10 10 9 2
43 1 10 9 1 12 10 0 9 13 1 10 9 2 3 15 13 9 1 10 9 7 15 15 13 1 9 13 1 10 15 1 10 9 2 1 10 9 1 11 1 10 11 2
29 16 15 15 13 2 11 7 10 9 1 9 0 7 8 0 15 13 1 10 9 2 15 3 4 13 1 10 9 2
36 1 10 9 0 2 10 0 9 13 10 9 13 10 0 12 1 11 1 10 9 11 11 2 16 13 10 9 1 9 7 9 13 1 10 9 2
40 15 16 3 15 13 1 13 13 10 9 1 10 9 16 8 13 1 9 7 1 10 9 1 10 9 0 16 13 13 1 10 15 10 0 9 0 16 15 13 2
26 13 11 7 11 1 10 11 11 1 11 3 1 13 1 10 9 2 3 1 10 11 1 11 1 11 2
24 1 3 16 11 11 2 11 13 10 9 0 1 9 1 11 1 12 2 13 10 0 9 0 2
19 11 13 1 11 13 1 10 9 1 9 2 7 1 11 1 10 9 0 2
26 15 13 11 11 1 11 2 1 9 1 10 3 9 1 11 11 11 1 11 2 1 10 9 1 12 2
13 10 9 1 9 13 1 12 8 2 2 9 8 2
31 11 13 16 2 13 1 10 0 9 1 9 1 11 2 9 2 10 9 1 9 1 9 2 11 2 15 4 13 1 9 2
42 3 3 1 10 9 2 10 12 1 11 1 12 10 11 13 10 9 9 13 1 12 9 2 12 9 3 2 1 9 0 1 10 9 1 11 2 1 10 9 1 11 2
15 1 10 9 2 13 10 9 1 10 9 1 10 9 0 2
46 1 12 13 1 10 11 11 2 7 13 3 0 1 10 9 1 10 9 7 9 1 9 11 11 7 1 10 9 11 11 11 2 15 15 13 1 10 9 2 10 9 7 9 11 11 2
21 1 12 9 2 11 11 15 13 1 10 9 1 9 1 9 16 15 13 10 9 2
11 13 1 10 9 1 9 1 11 1 12 2
55 10 10 9 3 13 13 11 10 11 2 12 2 12 7 12 2 12 2 2 11 11 2 12 2 12 2 2 11 2 12 2 12 2 2 11 2 12 2 12 2 2 11 2 12 2 12 2 7 11 2 12 2 12 2 2
11 13 0 9 1 10 9 1 11 11 11 2
13 1 10 9 10 9 1 10 9 4 13 15 9 2
35 10 9 2 1 11 1 10 9 2 4 13 1 10 9 1 9 1 9 2 7 16 11 11 3 13 1 9 1 9 1 15 13 1 11 2
13 4 13 1 9 1 10 9 1 9 1 11 11 2
33 10 9 3 0 2 0 1 15 2 1 10 9 1 9 7 1 11 2 7 1 15 9 2 2 7 1 10 9 0 1 10 9 2
26 10 9 9 1 9 4 4 13 3 1 10 0 9 1 9 7 1 9 1 12 7 3 9 1 9 2
34 7 15 13 3 16 8 2 13 10 9 2 9 16 3 3 13 1 2 8 2 8 2 2 3 8 13 9 1 10 9 1 10 9 2
19 13 3 0 1 13 1 10 9 2 3 16 10 9 13 3 0 7 0 2
29 1 9 2 12 9 0 2 11 11 7 11 11 2 13 10 9 1 10 11 12 15 13 10 12 1 11 1 12 2
41 3 15 15 13 1 10 0 11 11 10 15 4 13 1 10 11 7 13 10 9 0 1 9 2 10 9 15 4 13 1 12 2 13 1 4 13 3 1 10 11 2
53 10 9 1 11 11 11 1 11 7 10 9 0 1 10 9 0 1 10 9 7 9 1 10 11 11 2 11 11 2 15 4 13 1 10 0 7 0 9 1 9 0 16 13 3 10 9 1 9 9 2 8 2 2
13 13 10 12 5 1 10 9 1 9 0 1 9 2
17 3 2 10 9 1 10 11 11 11 4 4 13 1 10 9 0 2
11 2 3 15 13 15 16 13 2 2 13 2
21 1 9 1 10 9 2 11 11 13 10 2 9 1 11 2 9 1 10 9 11 2
23 1 12 2 10 9 15 13 1 10 9 0 1 4 13 1 10 9 1 9 13 1 3 2
36 3 12 9 2 10 9 1 9 15 4 13 1 10 9 0 16 15 13 1 10 9 2 1 15 1 10 9 1 9 3 3 13 10 9 0 2
32 10 9 1 10 9 13 1 13 1 2 11 11 11 2 10 9 3 13 1 11 11 2 10 16 3 13 10 2 11 11 2 2
11 10 9 1 10 9 13 12 9 3 0 2
19 15 3 13 9 1 10 9 2 13 1 10 10 9 1 10 16 15 13 2
27 3 1 10 9 2 10 9 13 10 0 9 10 12 1 11 2 4 10 0 9 13 1 10 9 1 11 2
21 10 11 13 15 1 10 9 3 0 1 10 9 0 1 11 7 1 10 9 0 2
40 11 11 11 2 9 1 10 11 2 2 11 11 11 2 9 1 10 11 7 11 2 9 2 2 11 11 2 11 2 0 9 1 10 11 11 11 1 11 2 2
33 1 10 9 2 15 13 16 10 9 4 13 1 12 9 1 9 1 9 2 4 15 13 1 10 9 0 3 1 12 9 1 8 2
25 7 10 9 15 13 1 10 9 1 9 1 11 2 3 16 10 9 3 13 10 9 1 10 11 2
19 11 11 1 10 11 2 10 11 2 11 2 12 2 13 10 9 0 0 2
55 0 1 10 9 16 15 13 10 9 1 10 2 11 0 2 7 1 13 15 0 1 2 10 9 1 9 7 9 2 16 3 13 1 13 2 1 12 10 0 9 11 1 10 11 15 13 10 9 1 13 15 1 11 11 2
23 11 10 11 13 10 9 1 10 9 1 11 11 1 11 2 3 1 10 9 11 1 11 2
25 11 11 11 11 13 10 9 1 9 9 0 13 1 11 2 1 10 9 1 10 11 2 11 2 2
39 11 11 2 1 10 12 9 1 9 2 4 13 1 7 1 10 11 2 13 1 9 10 9 2 10 9 2 10 9 2 10 9 7 1 9 1 10 9 2
27 10 9 4 13 1 10 9 1 11 7 11 11 2 16 16 10 9 11 2 11 2 11 13 8 2 9 2
19 10 9 13 9 0 13 1 9 1 10 9 10 9 0 4 13 10 9 2
14 1 10 9 2 15 13 9 0 1 10 9 1 11 2
32 2 10 9 13 3 3 1 10 9 1 11 2 3 7 15 3 13 13 1 10 0 9 16 15 13 10 9 2 2 13 11 2
15 10 9 1 10 9 4 13 1 10 9 1 9 1 9 2
10 11 15 13 1 12 1 10 9 0 2
58 10 12 13 10 9 7 13 16 13 2 10 0 7 0 9 2 1 10 11 2 1 0 9 1 10 9 0 1 10 9 1 9 7 1 10 9 1 10 15 4 3 13 1 4 13 7 13 2 13 0 13 1 10 9 1 9 2 2
31 13 0 3 1 13 1 10 9 15 11 11 1 9 7 1 11 2 11 7 11 11 1 10 11 1 11 1 11 11 11 2
46 16 1 10 9 1 10 9 8 2 10 9 1 10 9 2 3 3 1 10 9 0 2 15 13 1 10 0 9 2 16 13 1 10 9 1 0 9 1 9 15 13 7 3 3 0 2
36 10 9 13 1 10 9 1 9 1 9 7 9 2 15 16 13 1 0 1 10 9 1 9 1 11 2 9 13 1 9 3 0 16 10 9 2
76 15 13 2 3 3 2 1 10 9 7 9 1 10 15 10 9 4 3 13 3 0 1 16 10 9 13 3 0 1 10 9 1 10 11 2 1 9 1 11 2 11 1 11 2 10 9 0 2 1 11 11 7 2 1 9 2 10 9 1 10 11 1 11 11 11 2 9 1 9 1 10 9 2 1 12 2
40 10 9 0 13 11 11 11 1 11 2 11 2 13 1 12 2 2 16 13 1 9 1 10 9 1 11 2 7 11 11 2 13 10 12 1 11 1 12 2 2
32 9 1 10 9 2 13 1 9 10 9 0 1 10 9 1 9 0 7 3 3 11 1 11 2 9 16 13 1 12 1 12 2
21 13 16 13 1 10 9 1 10 9 16 13 7 1 15 3 15 13 10 12 9 2
40 3 1 10 9 0 10 9 0 15 13 1 0 9 1 10 9 0 3 3 1 10 9 0 1 10 9 2 7 3 1 10 9 1 0 9 13 1 10 9 2
41 10 9 2 16 3 4 13 1 13 10 0 9 3 1 10 9 1 9 13 1 10 9 11 2 13 13 1 9 10 9 2 16 13 10 9 1 10 9 13 3 2
22 10 9 13 0 9 0 7 9 13 13 1 10 9 15 1 10 3 0 1 10 12 2
13 4 13 1 0 9 1 10 9 1 10 9 12 2
13 13 9 1 9 2 16 4 13 1 13 3 0 2
28 11 11 2 1 10 9 0 2 11 1 11 2 7 13 15 1 10 0 9 2 13 10 9 2 11 11 2 2
15 10 9 13 13 10 12 9 13 10 9 1 10 9 0 2
28 1 9 1 15 2 4 13 16 10 9 2 0 2 15 4 13 1 2 10 9 1 10 9 1 10 9 2 2
39 10 9 1 10 11 11 16 13 10 9 1 10 9 1 10 9 0 2 4 13 1 10 2 11 11 2 2 2 11 1 11 2 7 2 11 7 11 2 2
26 10 9 1 13 10 9 4 4 13 16 10 9 13 3 0 3 1 10 9 7 16 4 13 10 9 2
87 13 12 9 1 9 16 13 10 9 1 11 2 10 9 1 10 9 16 13 10 9 1 10 11 11 2 11 10 9 2 9 2 9 2 9 16 13 10 9 0 1 10 0 11 11 2 0 9 1 11 2 9 13 1 13 10 9 0 1 10 11 2 3 7 0 9 16 13 10 9 1 10 9 16 13 9 1 10 9 0 1 11 1 10 9 12 2
30 15 13 1 9 1 9 2 7 15 13 16 15 1 10 9 0 13 10 9 1 10 9 0 13 1 10 9 1 9 2
20 4 13 10 0 9 1 11 7 10 10 9 1 10 9 2 10 9 13 2 2
43 10 9 0 13 3 1 10 9 0 1 10 9 1 10 9 1 10 11 11 2 3 4 13 10 9 1 10 9 1 10 9 7 0 9 16 4 13 10 9 1 10 9 2
18 10 0 9 13 13 2 16 13 16 13 2 13 1 10 9 1 11 2
28 1 12 9 15 13 16 4 4 13 1 9 1 10 9 1 12 1 11 2 7 9 0 13 16 13 1 12 2
17 3 10 10 9 13 10 9 10 9 7 10 9 1 10 9 0 2
16 10 9 3 0 2 3 7 3 13 10 9 7 3 10 9 2
6 3 4 13 1 9 2
17 4 13 1 0 9 1 10 9 11 11 2 10 9 2 12 2 2
17 11 13 10 9 11 11 2 10 9 1 10 9 1 10 11 11 2
49 11 11 13 10 9 0 0 13 1 12 16 3 13 12 9 0 1 10 9 7 9 0 2 10 11 11 11 1 11 7 10 11 11 1 11 2 13 1 12 7 16 13 10 0 1 10 9 0 2
19 10 9 0 13 3 15 4 13 1 10 9 7 15 4 13 1 0 9 2
42 13 1 15 7 1 10 9 13 1 10 9 2 9 1 9 7 9 1 10 9 2 10 15 15 13 0 2 2 10 9 15 13 13 1 10 9 10 9 7 10 9 2
11 15 13 10 9 1 10 9 2 11 2 2
29 3 2 10 9 0 1 11 1 10 9 13 13 7 13 1 9 0 2 16 13 15 1 10 9 0 1 10 9 2
13 13 1 10 0 9 2 15 13 1 10 0 9 2
23 13 10 9 1 9 16 13 0 1 13 9 2 13 12 9 0 7 0 1 10 9 0 2
77 11 7 11 2 13 1 10 9 1 9 2 2 8 8 2 2 2 8 8 2 2 2 8 2 2 2 8 2 2 2 8 8 2 2 7 2 8 8 8 8 2 2 13 10 9 1 9 1 10 9 2 11 11 11 2 16 1 10 9 2 1 12 2 13 1 10 9 11 2 13 3 9 1 10 9 12 2
11 15 13 1 9 7 10 9 7 0 9 2
18 10 9 0 1 10 9 13 11 2 16 15 13 1 10 9 1 11 2
20 1 10 11 2 13 11 11 1 11 2 9 1 10 9 1 11 13 10 9 2
38 10 9 0 1 11 2 1 9 2 11 11 11 2 13 10 9 0 1 12 9 2 12 9 2 1 9 2 13 1 11 2 11 2 1 10 11 11 2
9 10 9 2 3 2 13 3 0 2
13 10 9 0 15 13 1 3 1 12 9 1 9 2
14 2 10 0 9 2 1 10 0 9 1 9 15 13 2
48 1 9 1 13 10 9 1 10 9 2 10 9 1 10 9 2 9 2 1 13 10 9 1 10 11 4 4 13 1 10 9 2 11 11 2 2 16 1 9 0 4 4 9 1 2 9 2 2
38 1 9 13 1 10 9 11 2 11 1 10 9 1 10 9 11 11 11 7 10 9 1 11 7 1 10 9 1 10 9 11 2 11 1 10 9 11 2
22 10 11 1 10 11 13 10 9 13 1 10 9 9 1 10 11 11 1 11 2 11 2
45 10 0 9 13 12 7 12 9 13 3 3 1 10 9 7 10 9 1 9 1 9 7 10 1 10 9 13 9 2 13 13 10 9 1 9 1 9 2 15 1 9 7 15 3 2
3 9 1 9
19 13 3 16 13 10 9 1 10 9 4 1 13 10 9 1 9 1 9 2
14 10 9 13 10 9 1 0 9 2 13 1 10 9 2
40 13 10 9 1 12 9 2 12 9 0 2 2 7 15 13 1 12 8 2 12 5 2 1 10 9 1 10 9 11 2 9 1 11 2 2 13 1 10 11 2
19 7 10 9 4 13 3 0 2 16 13 9 1 13 9 0 1 10 9 2
20 10 9 4 13 12 9 1 9 10 9 11 7 11 1 9 1 11 11 11 2
42 16 10 9 1 10 9 13 1 10 9 1 1 10 11 2 10 9 13 3 10 9 0 10 9 1 10 11 1 10 11 2 1 10 15 3 13 10 9 1 10 9 2
18 10 9 4 3 13 3 10 9 1 10 9 7 10 9 16 15 13 2
40 10 9 1 11 11 2 11 4 13 9 0 7 11 11 1 12 2 1 10 9 1 10 9 12 2 12 1 10 12 1 11 2 1 9 1 10 11 1 11 2
13 10 9 13 10 9 0 1 11 1 10 9 0 2
136 1 9 1 10 11 1 10 11 13 7 13 10 9 1 11 11 2 7 9 1 10 0 9 13 10 9 0 1 10 0 9 1 10 9 1 11 2 15 13 1 10 9 7 15 13 1 9 1 10 11 11 11 2 1 9 1 9 13 1 9 0 3 13 3 7 10 9 1 10 9 1 9 13 11 2 11 2 11 2 11 10 1 11 2 13 1 10 9 1 11 2 1 11 2 1 16 10 9 1 11 7 11 13 16 13 1 10 9 10 9 1 9 0 1 9 13 1 15 0 1 11 11 1 11 1 10 9 3 1 10 9 1 10 11 0 2
33 10 0 9 1 10 9 1 10 9 1 11 2 16 13 1 10 9 1 10 11 2 15 13 1 9 1 10 9 0 11 2 11 2
14 3 2 1 11 13 10 9 3 15 13 0 7 0 2
35 10 9 13 16 10 9 1 13 13 1 10 9 7 15 13 1 15 0 1 9 1 10 9 2 10 0 9 13 1 10 9 1 10 9 2
37 10 9 0 1 10 9 4 13 1 10 9 0 2 5 2 7 10 9 11 2 8 2 2 15 1 9 2 1 1 10 12 9 0 16 13 8 2
8 13 10 9 0 1 10 9 2
3 11 11 2
37 15 1 10 9 0 1 9 13 10 9 1 11 7 10 9 2 7 10 9 4 13 10 0 9 9 1 10 9 13 1 10 9 3 1 10 9 2
14 10 9 1 9 4 13 1 13 1 10 9 1 11 2
22 12 9 1 10 9 1 9 16 13 1 10 9 11 7 16 13 1 10 11 1 11 2
17 13 9 3 0 7 4 9 1 9 1 9 1 9 0 7 9 2
14 13 0 3 1 10 9 7 1 10 9 1 10 15 2
31 10 9 7 10 9 13 0 2 10 9 13 0 0 0 2 15 9 16 10 9 2 7 10 0 13 9 0 1 10 9 2
24 1 10 0 11 2 15 4 13 12 9 7 12 9 2 16 3 3 15 4 13 10 9 0 2
20 10 9 7 9 13 11 0 2 10 9 2 2 10 9 1 9 7 9 0 2
24 10 11 1 11 7 10 11 0 1 11 13 10 11 1 10 11 10 11 12 1 11 1 12 2
15 13 1 10 9 0 1 10 9 1 10 9 1 10 11 2
15 13 1 10 9 1 13 7 3 15 13 3 0 2 3 2
33 1 4 1 13 15 2 13 15 9 15 13 11 1 11 2 11 15 13 7 11 15 13 13 1 10 9 2 1 10 9 1 11 2
36 3 2 1 10 12 5 9 9 1 11 11 13 10 0 9 1 10 0 9 1 10 9 0 1 9 1 0 9 0 16 13 1 10 9 0 2
18 10 10 9 13 1 0 9 2 13 10 0 9 1 9 1 10 9 2
73 10 0 9 1 10 9 2 16 4 13 1 9 3 1 9 1 10 9 1 9 0 7 3 1 10 4 13 1 10 11 1 11 1 10 11 2 10 9 1 10 9 13 16 10 11 13 1 10 9 1 10 9 1 10 9 1 16 10 9 1 9 3 13 1 10 9 1 10 9 11 10 11 2
30 10 9 13 9 3 9 7 9 2 16 13 3 1 10 9 7 13 10 9 0 16 15 13 1 10 9 1 10 9 2
13 10 9 13 0 7 3 4 13 3 1 12 9 2
29 1 10 9 1 12 2 15 13 1 0 1 9 10 9 0 1 11 7 11 2 10 0 9 1 12 9 1 0 2
12 10 9 1 9 1 10 9 13 1 9 12 2
12 10 9 0 15 13 2 1 9 2 1 9 2
9 3 4 4 13 1 10 9 1 9
15 13 10 9 1 9 1 9 7 13 2 13 10 11 11 2
38 11 5 11 15 13 1 12 2 9 1 10 9 1 10 9 1 9 1 0 9 0 7 11 11 2 1 9 0 1 9 2 9 7 9 1 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
7 10 9 13 3 15 13 2
15 15 1 10 9 3 0 1 9 0 13 10 11 11 11 2
11 10 9 1 11 15 13 13 1 10 9 2
18 13 1 11 11 1 9 16 15 13 10 9 2 9 7 9 11 11 8
34 10 9 0 1 10 9 2 1 11 11 2 13 2 11 8 11 11 2 11 11 2 2 2 3 4 13 2 7 13 1 0 9 0 2
14 15 13 16 13 10 0 9 3 7 13 10 0 9 2
24 3 15 13 0 9 1 9 7 9 2 16 3 15 13 1 10 9 0 1 10 11 11 11 2
16 11 11 11 2 12 2 12 2 13 10 9 2 7 9 0 2
26 1 16 13 1 10 11 1 10 11 2 11 11 2 13 1 10 9 2 13 10 10 9 1 10 9 2
20 11 13 13 15 2 7 13 1 11 13 10 9 16 15 15 13 1 4 13 2
34 11 11 11 2 11 2 11 2 12 1 11 1 12 2 11 1 11 2 12 1 11 1 12 2 2 9 0 7 9 1 11 1 11 2
30 10 9 1 9 7 9 13 10 9 11 2 10 9 11 11 2 11 1 11 7 10 9 11 1 11 7 11 1 11 2
19 10 12 1 11 1 11 13 9 1 10 9 11 11 1 11 2 8 2 2
56 15 13 10 9 2 10 9 1 3 12 9 2 4 13 1 10 9 7 10 15 2 3 0 2 13 10 9 1 12 9 7 9 2 1 10 9 2 13 1 13 15 15 3 0 13 1 9 10 9 3 0 1 10 9 0 2
19 15 13 10 0 9 1 13 1 10 1 11 7 1 10 9 13 1 11 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
57 13 3 9 1 9 1 10 9 1 11 11 11 2 7 3 3 1 10 1 10 9 0 11 11 11 2 16 15 13 2 15 3 13 3 10 0 9 2 7 10 3 0 2 2 16 15 13 1 10 9 7 15 13 15 1 11 2
40 10 9 0 13 10 9 1 9 13 2 16 11 11 13 10 2 11 1 11 2 2 7 16 13 1 10 9 1 9 0 2 7 1 9 1 9 7 13 9 2
55 11 11 2 11 2 12 1 11 1 12 2 11 11 2 12 1 11 1 12 2 13 10 9 0 1 9 0 2 13 1 9 7 9 1 10 9 1 10 11 1 11 2 1 10 9 1 10 9 0 1 10 11 11 11 2
12 11 13 10 9 1 9 0 1 10 9 11 2
25 1 10 12 9 9 1 10 9 1 9 0 2 10 9 13 16 13 10 0 9 15 13 10 9 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
32 10 8 1 11 13 10 0 9 1 16 15 13 1 10 0 9 1 10 9 1 10 16 15 13 9 2 9 7 9 1 9 2
29 13 10 9 11 11 13 16 3 4 13 10 16 13 10 0 9 2 9 1 10 0 2 10 11 1 10 11 2 2
28 15 13 10 9 0 1 10 12 5 2 15 16 13 1 15 16 13 1 10 9 9 1 9 1 9 3 0 2
21 3 2 4 13 1 10 9 1 11 7 10 9 2 3 1 13 10 9 7 9 2
23 10 9 15 15 13 1 15 3 0 2 10 9 13 0 7 10 9 13 0 7 3 0 2
29 11 2 11 2 13 10 9 1 10 9 0 2 13 1 10 11 2 1 10 9 0 3 0 1 15 1 10 9 2
29 15 13 10 9 0 1 10 9 2 15 0 2 10 9 0 15 9 2 9 1 9 7 1 9 2 9 1 9 2
51 1 10 9 2 16 13 1 10 11 10 0 9 1 10 0 9 1 10 11 1 11 1 10 11 11 2 11 2 2 10 11 1 11 13 10 9 0 1 10 9 1 10 10 9 2 1 9 1 10 15 2
24 15 1 10 0 9 1 10 9 0 13 10 9 0 1 9 7 9 1 10 9 1 10 9 2
56 11 11 11 13 1 11 11 2 11 2 11 11 2 10 12 1 11 1 12 2 16 1 10 9 0 13 1 10 9 12 1 11 1 12 2 11 13 10 0 9 1 10 9 1 10 9 1 10 9 1 10 9 1 10 9 2
14 11 13 10 0 9 16 4 13 15 1 10 0 9 2
49 15 1 10 9 1 11 2 8 2 13 10 9 10 12 1 11 1 12 2 13 10 9 1 10 9 1 10 9 2 15 13 7 13 1 10 9 7 13 1 10 9 12 2 12 1 10 9 12 2
54 10 9 1 10 9 2 11 11 11 11 13 1 13 10 9 16 10 9 9 13 10 9 1 10 9 1 10 0 9 16 15 13 1 13 9 2 10 9 7 1 15 3 4 13 15 10 9 0 1 9 7 10 9 2
6 3 13 1 9 0 2
17 10 0 9 13 16 10 9 1 11 13 10 9 2 9 1 9 2
23 10 9 0 3 7 13 15 2 7 10 9 2 10 9 2 9 2 7 15 1 9 2 2
15 3 15 13 13 10 9 1 11 2 13 1 11 3 0 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
33 15 13 16 10 9 0 4 7 13 15 1 11 1 4 13 1 9 1 9 0 7 3 13 16 10 9 0 4 13 1 10 9 2
40 10 9 0 11 11 13 1 10 11 11 1 11 11 2 11 2 1 10 9 16 15 13 1 9 1 9 1 10 8 9 1 11 11 11 2 13 3 10 9 2
35 11 11 13 16 2 4 13 15 10 9 1 10 0 1 1 10 0 1 10 9 2 2 10 9 3 0 1 10 16 13 3 1 10 11 2
26 10 9 4 13 1 9 9 5 12 1 10 12 1 11 1 12 1 10 0 9 1 9 1 11 11 2
20 15 13 9 1 15 1 10 9 1 11 2 3 10 9 13 1 10 0 9 2
10 4 13 1 11 2 11 7 11 11 2
11 15 0 13 10 9 0 1 9 2 9 2
26 1 10 9 13 10 9 0 1 0 9 1 10 9 12 2 12 7 10 11 1 11 1 10 0 9 2
36 10 9 2 13 1 10 11 8 8 11 11 11 2 4 13 9 1 12 9 16 2 1 10 9 1 9 16 15 13 3 2 3 13 9 0 2
25 1 13 10 9 1 9 2 13 10 9 1 13 1 10 9 0 2 3 1 9 1 13 1 12 2
16 4 13 1 0 9 1 10 0 9 1 10 11 12 1 12 2
18 10 9 13 10 9 0 1 5 12 9 1 10 5 12 1 10 9 2
6 10 9 3 13 0 2
18 15 13 0 1 10 9 1 11 11 7 10 3 3 0 9 1 11 2
28 1 10 0 8 13 13 10 0 9 12 2 12 1 0 9 1 10 9 0 2 9 1 11 7 9 1 9 2
21 10 9 1 10 9 0 13 10 9 1 9 7 9 2 1 10 9 11 7 11 2
64 10 11 1 11 1 10 11 7 10 11 1 10 11 1 11 2 13 1 10 9 11 11 2 13 13 2 10 9 0 1 10 15 13 1 9 10 9 0 3 1 10 9 0 2 10 9 0 2 7 10 9 1 10 9 2 10 9 2 7 10 9 0 2 2
10 1 10 9 13 9 7 10 9 0 2
13 15 13 3 3 15 1 10 9 7 1 10 9 2
34 10 11 13 10 9 7 9 0 2 13 1 10 9 1 10 11 1 10 9 1 11 2 11 2 1 10 9 0 1 10 11 1 11 2
15 1 10 9 13 10 9 16 13 10 12 9 1 10 9 2
17 10 9 1 9 4 13 3 1 9 0 7 0 1 10 9 0 2
9 13 10 10 9 0 1 10 9 2
30 13 13 1 11 7 3 11 1 10 9 1 10 9 2 13 10 9 1 10 9 0 2 2 16 10 0 9 13 11 2
30 1 15 15 13 9 0 7 0 2 10 9 3 1 10 11 1 10 11 2 9 1 0 9 3 1 10 9 1 11 2
29 10 9 13 1 11 13 3 7 0 1 13 1 11 2 16 10 9 3 13 1 10 15 13 1 10 9 1 11 2
20 14 2 16 16 13 1 10 11 2 2 3 13 1 9 1 15 1 10 9 2
18 3 1 10 9 2 11 13 10 9 1 9 0 1 13 15 1 9 2
20 13 3 3 10 9 2 1 10 9 3 13 1 15 2 7 15 13 3 0 2
8 10 9 11 13 9 1 11 2
35 1 10 9 2 10 9 15 13 1 9 0 1 9 1 10 9 0 2 3 13 10 9 0 1 10 9 0 2 10 9 0 7 10 9 2
37 1 12 15 15 13 10 9 1 11 2 11 2 11 7 9 2 7 15 3 13 1 13 10 11 1 11 2 1 9 1 10 9 11 11 7 11 2
39 1 9 2 10 9 1 10 9 1 11 13 0 2 3 16 1 9 1 10 9 7 10 9 1 9 1 9 4 7 13 10 9 10 12 1 11 1 12 2
40 1 9 1 10 0 9 0 2 4 13 10 9 0 1 11 7 11 2 10 9 0 13 2 13 10 9 1 10 9 7 13 9 1 10 9 0 1 10 9 2
38 15 1 10 9 3 0 1 10 9 3 7 13 12 9 7 15 13 13 12 2 3 7 13 16 4 13 1 13 15 1 10 10 0 9 1 10 9 2
41 1 10 8 1 9 1 9 11 11 4 13 1 10 9 0 1 10 9 1 9 0 2 10 9 1 9 1 11 2 13 1 10 9 0 7 3 3 0 1 9 2
41 3 1 10 9 13 2 16 13 1 10 9 1 9 7 9 0 1 10 9 1 10 9 2 4 7 13 3 10 9 1 11 11 2 0 9 1 10 9 1 9 2
45 15 13 1 9 3 1 10 9 1 10 9 1 10 9 15 4 13 1 12 1 0 9 2 11 11 11 2 11 11 2 11 1 11 2 11 1 11 2 11 11 7 11 11 2 2
28 11 7 10 0 11 11 1 10 11 11 11 11 13 9 1 9 10 12 1 11 2 16 13 10 9 1 9 2
14 10 9 2 0 2 1 10 9 2 7 10 9 0 2
15 11 13 1 10 9 1 3 1 12 9 3 1 10 9 2
22 10 9 13 1 10 9 15 13 0 7 4 1 13 15 10 9 1 9 1 0 9 2
32 15 16 3 13 0 13 16 10 0 2 9 2 1 9 13 2 1 9 2 10 9 1 9 3 0 1 10 9 1 10 9 2
53 10 9 11 13 13 1 10 9 1 8 8 16 13 2 9 1 9 2 2 2 9 2 1 8 2 8 1 2 13 2 2 2 16 13 10 9 1 10 9 1 10 9 13 1 9 1 9 1 11 1 10 9 2
38 4 13 1 9 2 7 10 9 4 13 1 10 9 2 10 9 0 1 9 0 2 1 12 9 2 13 1 10 9 0 1 10 0 9 0 1 11 11
24 10 11 13 10 9 7 10 9 1 10 9 0 2 10 9 1 10 9 7 9 1 10 9 2
5 13 9 7 9 2
18 2 15 13 1 10 12 9 7 3 15 13 7 15 13 1 10 9 2
32 3 2 10 9 8 13 12 9 2 10 9 2 16 3 15 13 1 10 9 1 9 11 7 15 0 2 13 1 10 9 11 2
17 10 9 0 7 0 1 9 1 9 5 4 4 13 1 10 9 2
31 10 11 11 1 11 1 11 2 11 11 7 11 2 13 7 13 10 9 1 10 9 0 1 11 1 10 9 0 7 0 2
27 1 10 11 2 11 2 13 10 9 2 12 2 7 13 1 10 9 1 10 11 1 10 12 1 10 12 2
36 3 15 10 9 7 15 2 3 15 13 1 15 0 16 13 2 16 13 16 3 13 10 9 16 15 13 8 8 16 15 16 13 9 15 13 2
10 10 9 11 11 13 16 13 12 9 2
11 11 11 3 13 1 11 11 1 10 9 2
42 2 10 0 9 13 10 9 0 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 11 11 2 11 11 7 11 11 2
14 13 10 9 1 16 3 15 13 16 15 13 10 9 2
9 15 15 4 13 7 15 4 13 2
22 3 13 9 1 9 2 9 0 2 9 7 16 15 13 9 7 3 1 9 0 0 2
15 15 13 11 11 7 11 11 1 10 9 1 10 9 0 2
29 16 4 13 1 10 9 2 10 9 1 11 7 11 2 15 13 1 10 9 0 1 10 9 0 1 9 1 11 2
5 15 13 1 11 2
26 10 9 0 13 10 9 1 10 9 7 1 10 9 1 10 9 7 10 9 13 10 9 1 9 0 2
14 13 12 9 1 10 9 0 1 12 9 2 9 5 2
37 15 13 1 13 10 12 9 11 11 11 11 2 1 10 9 0 1 12 8 12 8 2 1 12 11 2 1 10 9 0 1 12 8 12 8 2 2
14 15 1 10 9 0 1 10 9 4 13 1 10 9 2
12 13 10 0 9 1 11 2 13 1 11 11 2
26 10 9 15 13 1 9 0 2 12 9 2 7 10 9 1 10 0 9 13 13 15 1 10 9 0 2
21 11 2 12 16 15 13 1 10 2 9 1 9 2 1 10 9 0 1 10 9 2
17 13 10 9 1 9 1 9 13 9 1 9 1 13 1 10 9 2
12 10 9 13 0 1 13 10 9 1 9 0 2
16 1 10 9 1 10 9 1 11 2 15 13 1 12 1 11 2
55 1 10 9 16 10 9 13 1 10 9 2 10 11 11 7 10 9 16 1 15 7 15 13 2 11 11 2 13 10 9 3 0 1 10 16 3 15 13 1 10 9 10 9 9 1 10 9 13 1 11 7 11 1 11 2
58 10 12 1 11 1 12 13 10 0 9 2 11 2 2 13 1 10 9 1 0 9 1 13 15 1 10 9 1 10 9 7 1 10 9 1 10 9 2 2 13 10 9 1 9 7 13 1 10 9 1 10 9 1 10 9 1 9 2
25 10 9 13 0 9 2 13 10 9 11 11 2 16 13 1 10 9 2 10 11 11 1 11 2 2
53 10 9 1 9 2 13 10 9 0 2 4 7 13 10 9 0 2 7 1 0 9 13 1 13 1 10 10 9 0 16 3 13 1 10 13 1 15 7 13 0 2 3 7 15 13 1 10 9 1 10 0 9 2
6 0 9 1 10 11 2
29 10 9 1 10 9 15 13 9 2 7 3 0 2 16 10 11 13 0 15 12 2 3 2 1 10 9 0 2 2
29 3 1 10 11 11 10 11 13 10 9 13 1 9 1 9 13 1 10 11 11 16 13 10 9 1 0 1 9 2
24 10 9 16 13 10 11 13 3 0 7 13 10 9 1 10 9 0 1 13 15 10 0 9 2
16 11 13 10 9 1 9 7 10 9 1 9 1 10 11 11 2
13 16 10 9 15 13 1 10 9 13 1 10 9 2
53 1 10 9 1 11 11 2 11 13 9 1 9 2 1 15 10 11 11 2 13 3 1 13 1 11 1 10 11 11 11 2 11 2 16 13 1 10 9 1 11 2 7 11 11 2 10 9 1 10 9 11 11 2
11 10 9 11 13 10 9 1 10 9 0 2
5 15 13 1 11 2
17 10 0 9 2 11 11 13 10 11 2 10 9 1 9 1 9 2
49 7 10 9 13 3 16 3 1 4 13 1 10 11 1 10 11 2 11 11 11 2 2 1 11 2 4 13 15 1 11 2 1 10 13 1 10 9 2 1 10 15 13 10 9 1 3 12 9 2
25 1 9 0 2 12 2 2 4 13 1 11 2 7 11 13 1 9 1 11 2 3 13 13 15 2
32 10 9 2 13 1 11 1 10 0 9 1 10 11 1 11 2 4 13 7 13 10 9 1 9 0 1 9 1 10 0 11 2
27 10 9 0 4 13 1 13 10 9 1 10 9 16 15 13 2 7 1 15 9 4 13 1 9 1 9 2
25 3 2 3 13 9 7 9 1 9 2 7 3 13 1 9 10 9 1 10 9 1 10 9 0 2
18 11 13 10 9 0 1 10 9 1 11 2 13 1 10 9 1 11 2
23 1 12 2 13 1 10 9 1 10 9 1 9 2 15 4 13 1 11 2 11 7 11 2
16 11 15 13 1 13 2 7 13 16 10 9 4 4 1 13 2
30 1 9 2 16 10 9 15 13 1 11 11 1 9 1 12 1 11 2 15 13 3 1 12 9 1 10 2 11 2 2
12 13 3 1 10 9 13 1 11 2 11 11 2
13 11 13 10 9 0 1 9 0 1 10 9 11 2
11 11 11 11 3 13 1 9 1 10 9 2
15 15 13 1 9 2 9 2 9 0 2 9 7 10 9 2
19 13 10 9 1 9 8 7 13 1 9 13 10 9 7 10 9 13 0 2
23 1 12 10 9 4 13 9 1 11 7 11 15 13 3 3 13 1 11 1 11 7 11 2
16 1 10 9 13 10 9 1 0 9 1 10 0 9 1 9 2
24 11 2 11 2 11 2 11 2 11 7 11 13 9 2 7 10 9 13 3 10 9 1 11 2
17 1 10 9 0 1 12 13 12 9 2 13 1 12 9 1 9 2
20 1 15 2 1 10 9 0 1 9 15 13 16 10 9 15 13 1 10 9 2
32 8 8 9 8 0 9 12 2 12 2 1 12 1 11 2 1 10 15 15 13 10 9 1 10 11 7 11 11 1 11 11 2
20 10 12 1 11 1 12 4 13 1 11 1 3 4 13 1 9 0 9 3 2
30 15 13 10 9 1 11 11 3 1 11 16 13 10 9 0 1 9 1 2 9 2 2 1 10 0 9 1 10 9 2
16 13 10 9 1 10 9 1 11 11 2 11 11 2 1 12 2
31 16 10 9 4 13 9 1 9 1 10 9 1 11 2 11 7 10 9 2 10 11 2 13 0 7 13 9 1 10 9 2
36 10 9 0 0 1 12 2 3 13 1 9 0 13 1 10 9 1 9 1 9 1 10 12 1 11 1 12 2 16 13 1 10 9 0 0 2
26 15 13 0 1 15 9 1 10 2 11 11 2 10 9 1 10 11 11 1 10 9 9 1 11 11 2
23 15 4 13 1 9 1 9 2 9 3 0 2 3 1 10 9 2 7 13 1 10 9 2
8 11 15 13 13 1 10 9 2
20 11 3 13 3 13 10 9 1 11 11 2 11 2 7 13 1 10 9 0 2
43 10 9 0 1 9 2 11 2 13 10 11 10 9 0 7 13 16 10 9 0 15 13 1 9 1 12 9 1 9 7 9 0 13 1 10 9 1 10 9 1 0 9 2
17 11 15 13 13 10 9 3 7 10 9 2 7 10 9 3 13 2
37 13 9 1 10 12 1 10 11 1 11 2 11 1 11 2 11 2 11 11 2 11 11 2 11 7 10 11 11 1 11 11 11 11 11 2 11 2
18 13 9 1 11 11 2 15 1 10 9 1 10 9 1 9 1 11 2
14 3 1 10 9 3 13 10 9 1 9 1 10 9 2
8 15 13 10 9 1 10 9 2
25 1 10 9 2 3 13 0 3 1 10 9 11 7 13 10 9 1 10 9 2 9 1 10 11 2
33 10 9 4 13 2 7 15 13 10 9 1 4 15 13 1 10 9 0 2 10 9 0 13 0 7 10 9 3 4 13 3 0 2
11 13 9 1 10 9 1 9 1 10 9 2
24 1 10 0 9 1 11 2 1 10 9 1 10 9 11 4 13 10 2 9 2 1 13 9 2
9 15 13 1 11 1 11 7 11 2
44 1 9 1 2 11 2 10 11 11 2 10 9 1 11 11 2 15 13 16 11 4 1 4 11 9 3 1 10 9 1 11 11 5 12 2 3 10 0 9 1 11 4 13 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 8 2
24 1 3 1 10 9 16 15 13 1 10 9 2 7 10 15 13 1 10 9 15 16 13 0 2
10 9 1 11 10 12 1 11 1 12 2
35 1 9 2 10 9 1 11 3 15 13 13 1 10 9 1 10 9 3 13 2 7 10 9 0 4 13 3 1 4 13 1 9 3 0 2
11 13 10 9 1 10 9 8 1 10 9 2
29 1 12 11 13 3 7 13 1 11 12 2 13 10 9 1 10 9 1 11 2 1 10 15 10 9 13 12 9 2
24 15 13 16 10 9 15 13 10 9 2 7 13 12 9 1 9 2 13 10 15 15 15 13 2
4 11 2 12 2
6 4 13 1 11 11 2
19 13 1 11 2 1 10 0 9 7 9 1 9 1 10 0 0 9 11 2
20 10 9 13 0 2 13 3 1 12 9 0 7 9 1 9 0 7 1 9 2
8 10 9 13 1 9 1 9 2
70 10 9 1 9 1 10 0 9 15 1 10 9 0 2 0 7 0 2 15 13 1 9 1 10 9 1 10 0 9 0 16 13 10 9 1 10 9 7 16 13 3 1 10 9 1 8 2 7 1 15 1 10 9 2 9 1 10 10 9 16 13 9 0 1 10 9 1 10 9 2
23 10 9 16 13 1 9 2 1 10 9 1 10 9 1 10 9 2 4 13 1 10 9 2
33 1 3 1 10 9 2 13 15 3 0 7 9 9 3 13 7 10 16 15 13 1 9 2 16 3 13 15 7 13 1 10 9 2
7 13 1 10 11 11 1 11
27 1 11 7 11 4 13 10 12 1 11 1 12 2 7 1 11 13 10 12 1 11 1 12 2 1 11 2
26 1 12 13 12 9 1 11 11 1 11 7 1 11 2 7 12 9 1 11 2 11 7 11 1 11 2
24 1 10 0 9 2 11 13 16 11 2 1 10 9 2 3 13 1 10 9 0 1 10 9 2
21 4 13 10 9 1 10 10 9 1 9 1 10 9 7 15 15 4 13 1 9 2
36 1 10 9 1 10 9 2 11 15 13 1 9 0 7 1 9 1 10 9 2 11 13 10 9 1 10 0 9 1 0 9 2 11 11 11 2
14 15 1 10 0 9 1 9 16 4 13 1 10 9 2
19 13 13 9 2 9 1 13 1 10 9 9 1 9 1 10 9 11 11 2
82 10 9 13 10 9 1 3 9 0 1 10 9 1 13 10 9 13 10 2 0 9 2 16 13 15 1 10 0 9 0 7 1 15 2 15 13 13 1 10 9 0 16 15 13 1 10 0 9 9 1 0 9 1 9 13 1 10 9 16 15 13 1 10 9 16 13 15 9 7 13 15 16 15 13 1 10 8 0 1 10 9 2
29 1 10 9 13 1 10 9 15 4 13 1 9 10 9 1 10 9 1 9 1 9 1 10 9 1 10 9 0 2
12 13 10 0 9 0 7 9 1 0 9 0 2
19 3 4 4 13 1 10 9 1 10 9 1 9 3 7 1 9 1 9 2
20 1 12 10 9 13 10 9 1 9 1 5 12 9 1 5 12 1 10 9 2
16 9 1 10 9 1 11 1 11 2 11 11 7 11 11 11 2
11 13 10 9 1 9 0 7 1 9 0 2
15 10 9 1 10 9 8 13 9 1 10 0 9 1 11 2
12 10 9 1 9 1 10 9 13 1 5 12 2
15 11 11 11 2 11 2 12 2 13 10 9 7 9 0 2
57 1 10 9 2 10 9 1 16 3 15 13 1 10 9 13 10 9 0 1 10 9 1 9 1 10 9 2 2 3 2 10 11 3 13 1 10 9 1 9 7 1 13 15 15 13 1 9 1 9 2 0 7 1 9 2 2 2
23 15 13 1 13 10 9 1 10 9 2 13 1 10 9 1 10 9 1 13 10 0 9 2
10 4 13 0 12 9 7 3 13 9 2
30 16 15 13 1 15 15 4 13 1 10 3 12 9 1 10 9 2 13 3 12 9 2 13 1 11 11 7 11 11 2
39 13 10 9 0 2 10 9 11 11 11 2 10 16 13 10 9 1 11 16 11 11 13 13 1 10 9 11 1 11 1 10 9 1 13 10 9 1 9 2
6 9 1 10 9 1 11
23 1 9 2 1 10 9 12 2 10 9 1 11 11 2 11 2 15 4 13 1 10 9 2
16 10 9 3 15 4 4 1 13 3 1 10 9 1 10 9 2
68 3 13 9 7 9 1 10 9 1 10 9 1 16 15 13 10 9 1 9 1 10 9 7 3 4 13 10 2 9 2 13 1 9 1 11 7 10 9 1 9 2 1 10 9 1 10 9 0 1 10 9 1 10 9 2 3 10 9 13 1 13 1 10 9 3 15 13 2
31 10 9 16 15 13 1 10 9 4 13 1 10 9 1 9 1 9 7 1 13 10 9 0 1 10 9 7 10 9 0 2
19 13 10 9 1 12 9 16 13 10 9 0 2 3 10 9 7 10 11 2
17 3 15 13 10 9 1 11 1 9 1 11 2 3 1 9 2 2
78 10 9 1 11 7 11 10 11 13 10 0 9 0 1 10 9 1 11 2 7 1 0 9 0 3 16 1 15 15 13 15 1 10 0 9 0 16 13 3 1 9 1 10 9 13 1 11 1 11 2 3 1 10 9 1 9 1 9 1 9 2 1 0 1 10 9 1 10 9 0 2 1 10 15 13 10 9 2
15 3 1 10 9 11 1 11 13 10 9 1 10 9 0 2
23 10 9 1 10 9 4 13 3 0 1 13 1 10 9 1 10 9 1 10 15 4 13 2
45 10 9 13 0 7 13 2 3 13 7 13 2 7 9 0 1 9 1 9 7 1 9 2 7 1 10 9 10 9 1 10 9 4 13 1 0 9 0 7 9 13 1 9 0 2
41 10 11 11 11 11 2 11 2 2 1 9 11 1 11 11 2 13 10 9 16 13 7 15 13 1 10 9 1 10 11 11 11 2 10 11 1 10 11 1 11 2
12 1 9 12 13 1 10 9 1 12 12 9 2
13 15 13 3 3 2 0 9 7 13 1 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
28 15 13 1 11 11 7 13 1 11 11 2 9 0 3 0 1 10 9 2 16 13 10 0 9 1 9 0 2
15 3 2 1 10 0 9 2 11 13 0 9 1 10 9 2
28 10 9 13 10 9 1 0 9 13 15 3 1 12 9 2 7 16 10 9 13 1 9 0 1 10 10 9 2
15 10 9 13 15 1 10 9 0 2 1 1 13 1 9 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
22 11 13 10 9 7 9 0 2 13 1 10 9 1 11 11 2 1 10 9 1 11 2
30 10 9 0 1 11 11 2 1 9 11 11 11 11 2 13 10 9 0 1 10 9 0 1 9 1 11 11 2 11 2
36 11 11 11 11 11 12 13 10 9 1 9 0 13 1 10 9 2 16 13 10 12 1 11 1 12 7 13 10 12 1 11 1 10 0 8 2
20 10 12 1 11 1 12 2 13 13 10 9 1 9 1 10 9 1 10 9 2
44 1 10 9 1 11 2 11 13 10 9 1 9 7 9 2 10 0 1 15 2 7 10 16 15 13 1 10 9 13 10 1 11 11 1 10 2 11 1 11 11 1 11 2 2
8 13 10 0 9 7 9 0 2
6 13 0 1 10 11 2
28 9 1 15 13 10 11 1 10 11 2 1 11 2 10 11 1 11 2 1 11 1 10 11 7 10 9 0 2
32 10 0 9 1 9 1 10 9 0 13 10 9 0 16 13 10 9 0 3 0 2 15 0 1 10 9 1 9 1 10 9 2
22 3 2 15 13 1 10 9 1 9 1 10 9 2 1 15 1 10 9 9 1 11 2
38 11 13 13 1 9 7 9 2 1 9 1 13 10 9 1 10 0 9 1 10 9 7 1 9 1 13 15 3 0 2 7 3 13 3 0 9 0 2
16 1 10 9 15 13 1 9 1 10 9 11 11 2 1 11 2
26 11 4 13 1 10 0 9 7 13 0 13 10 9 0 1 11 12 13 11 11 11 1 10 9 11 2
9 10 9 13 10 9 11 11 11 2
18 10 9 13 3 10 9 1 10 9 2 13 1 15 10 9 1 11 2
5 15 13 1 11 2
12 0 3 13 15 9 1 15 15 13 1 15 2
19 1 9 16 15 4 4 13 10 9 15 4 13 10 9 0 1 10 9 2
25 13 1 10 0 9 2 11 2 11 2 11 2 11 7 11 2 10 12 9 1 10 9 1 11 2
31 1 10 9 10 9 0 1 11 13 7 10 9 13 1 10 9 2 3 3 1 10 9 0 15 13 1 10 9 3 13 2
51 16 10 9 1 11 13 11 2 15 13 1 13 1 10 9 13 0 9 1 9 2 1 16 10 9 13 1 10 9 0 1 10 9 1 10 11 11 1 10 11 2 15 4 13 1 10 11 1 10 11 2
23 1 10 0 9 2 10 9 13 1 10 9 0 1 9 16 15 13 1 11 7 1 11 2
21 2 7 11 7 11 11 4 4 13 1 10 11 7 10 11 2 10 9 0 2 2
26 10 9 11 4 13 1 10 9 16 15 13 10 9 2 11 11 11 7 11 11 2 1 10 9 12 2
26 11 15 13 9 1 10 11 11 1 10 11 13 1 12 2 1 10 15 1 12 13 10 11 11 11 2
30 10 9 13 1 10 9 1 10 16 10 9 0 4 13 15 1 9 7 9 16 13 13 1 10 9 7 9 15 13 2
11 1 10 0 9 1 12 1 12 13 9 2
27 15 13 1 0 9 1 10 9 16 3 13 12 9 7 16 15 4 13 2 16 3 13 9 13 15 3 2
24 11 11 1 11 13 16 2 11 1 11 2 4 13 1 10 9 9 7 10 9 9 1 9 2
51 9 1 10 12 13 0 1 10 11 11 2 16 13 11 2 9 0 1 10 9 11 2 2 10 11 11 2 9 1 10 9 1 10 11 11 2 7 10 11 11 2 9 1 10 9 1 10 11 11 2 2
9 11 11 2 9 1 10 9 2 2
7 3 15 13 1 10 9 2
27 13 1 11 2 11 0 2 7 13 1 11 11 2 11 11 2 7 1 10 9 1 10 9 11 11 11 2
32 13 13 3 1 10 9 1 11 11 16 13 10 9 0 1 10 16 3 3 13 9 1 13 1 10 9 10 15 13 10 9 2
13 10 9 0 2 1 9 2 15 13 1 10 9 2
20 10 0 9 13 1 10 9 1 10 9 2 0 2 0 7 0 1 0 9 2
36 1 10 9 10 9 4 1 13 15 11 11 11 2 9 16 1 9 15 13 1 10 11 7 1 10 9 1 10 11 1 10 9 1 10 9 2
12 11 13 10 9 1 13 1 10 9 1 9 2
20 3 1 12 10 9 15 13 1 10 11 11 1 10 9 1 10 9 1 0 2
43 1 12 2 11 13 1 0 1 10 11 1 11 2 10 9 13 1 11 2 11 2 3 15 13 1 10 0 9 1 9 7 9 1 10 9 1 10 8 11 2 11 11 2
35 10 9 13 16 13 0 15 13 16 1 10 9 1 9 3 4 13 15 3 9 7 3 13 15 16 13 13 15 0 1 1 9 10 9 2
26 3 11 2 11 7 11 15 13 1 10 9 1 9 1 9 1 11 2 3 1 16 10 9 13 3 2
10 4 13 10 12 1 11 1 10 12 2
52 10 11 13 10 9 0 2 16 13 3 1 9 13 1 9 10 9 2 13 10 9 1 9 1 10 9 2 13 9 7 9 1 11 3 16 1 10 13 10 9 1 11 8 15 13 1 10 9 1 10 9 2
12 11 11 13 10 9 1 9 1 10 9 11 2
20 11 13 1 0 9 0 1 11 7 13 10 9 0 1 10 9 13 1 9 2
52 1 10 9 15 4 13 1 10 9 1 10 9 0 1 0 1 9 1 10 9 7 9 1 10 9 2 7 15 13 1 10 9 15 13 10 9 0 1 10 9 10 9 2 16 10 9 3 13 1 10 9 2
36 10 9 0 4 3 13 1 10 9 0 1 10 0 9 1 10 9 2 13 10 9 1 10 2 9 1 10 11 2 1 10 9 8 2 0 2
35 1 10 9 2 11 13 16 10 9 13 10 9 3 0 1 9 1 0 9 2 10 15 2 1 10 9 0 2 3 4 4 13 7 13 2
20 1 15 16 13 9 0 7 3 13 10 9 1 10 9 2 11 13 1 15 2
59 1 10 12 9 2 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
59 7 3 10 9 4 13 1 10 9 0 2 10 9 13 16 15 13 1 9 1 10 9 16 15 4 13 1 10 9 2 13 13 2 10 9 3 13 3 10 9 1 10 9 1 10 9 1 9 1 9 2 3 15 4 13 1 10 9 2
4 13 1 11 2
7 4 13 9 0 1 11 2
29 10 9 13 9 1 10 15 2 13 1 10 9 16 13 2 1 9 1 9 1 11 2 9 1 11 7 9 11 2
7 13 10 0 9 1 9 2
16 13 0 9 1 9 2 7 10 9 13 0 1 10 9 0 2
36 10 9 1 11 2 10 9 13 1 3 10 0 9 1 10 9 0 2 4 13 1 10 9 0 1 10 9 0 1 10 9 1 10 9 0 2
19 11 11 10 9 13 2 2 11 7 15 13 10 0 9 1 10 9 2 2
23 10 9 13 10 9 1 12 9 1 9 0 1 3 1 0 9 1 10 9 1 10 9 2
17 16 3 10 9 0 13 0 15 13 1 10 9 1 10 9 0 2
47 10 9 13 10 9 1 12 5 5 2 10 15 12 5 5 13 13 1 9 2 2 10 9 1 12 9 2 7 10 9 1 9 13 1 12 8 2 5 5 2 1 9 0 1 12 2 2
16 1 9 1 10 9 10 12 5 13 0 7 0 1 10 9 2
10 10 9 16 13 1 9 0 13 0 2
20 1 13 10 9 2 10 9 7 10 9 16 13 1 11 4 13 1 10 9 2
14 1 9 7 9 9 13 13 1 10 9 1 10 9 2
50 1 15 2 11 4 13 1 12 9 16 2 1 11 11 1 10 9 0 2 13 1 10 9 7 10 9 1 0 9 1 11 16 13 10 10 9 1 10 9 7 10 9 7 13 10 9 1 10 9 2
10 11 11 4 13 11 11 1 10 9 2
45 1 9 2 16 10 9 1 9 13 1 10 9 1 13 10 9 1 10 9 0 1 11 11 10 11 11 2 12 2 2 3 13 1 11 2 0 9 4 1 13 1 10 9 0 2
14 13 10 9 16 15 13 9 16 3 13 15 10 9 2
42 3 1 13 10 9 1 12 9 1 9 1 10 11 2 1 11 11 11 7 3 1 11 11 11 2 2 11 11 13 10 9 1 12 7 13 10 9 1 10 11 0 2
21 1 10 12 10 9 15 13 1 0 9 1 10 9 11 11 7 1 11 1 11 2
18 0 9 13 10 0 9 1 13 13 10 9 1 9 0 7 0 9 2
10 10 9 0 13 1 12 9 1 9 2
59 1 9 2 1 12 13 10 0 9 1 10 9 1 9 0 0 1 10 11 7 2 1 12 2 10 0 9 1 1 10 9 1 9 1 9 2 1 10 0 9 0 9 11 11 1 10 11 2 0 1 10 9 1 10 9 1 9 11 2
29 13 0 10 9 16 13 10 9 11 1 10 9 2 1 15 13 2 10 11 1 11 2 11 1 11 7 11 11 2
17 10 11 13 1 9 2 7 10 9 4 13 1 9 0 1 9 2
21 16 16 15 13 9 7 13 1 9 13 3 10 9 13 2 3 13 10 0 9 2
79 1 11 3 4 13 13 15 1 10 9 1 10 12 9 0 1 11 1 13 11 7 11 10 9 4 13 1 10 11 2 1 10 11 11 2 15 1 10 0 9 1 10 9 16 3 13 10 11 11 12 2 12 1 10 9 0 1 12 1 10 9 1 11 2 11 7 10 11 16 13 15 1 10 9 3 0 16 13 2
15 10 9 10 11 11 11 11 11 7 10 11 2 11 11 2
32 1 9 2 13 9 1 11 2 7 9 1 9 2 1 10 15 13 9 1 11 2 11 7 11 2 15 1 9 7 1 9 2
68 1 10 9 1 10 9 1 12 7 1 12 10 9 0 1 10 9 13 9 2 1 9 2 1 11 7 10 9 0 1 9 2 1 10 9 1 9 11 11 2 10 9 11 7 11 11 2 15 13 1 9 1 10 9 1 9 13 10 0 9 1 10 11 7 3 9 0 2
2 13 3
10 13 1 10 9 1 13 10 9 1 8
17 8 3 0 2 0 7 0 2 15 13 13 1 9 7 13 9 2
20 1 9 1 15 2 2 10 11 11 2 13 10 0 9 13 2 7 13 2 2
36 11 13 10 8 0 1 10 11 1 11 2 2 11 2 11 2 13 1 9 0 1 10 9 1 10 11 11 1 11 2 9 0 1 11 2 2
40 10 0 9 1 11 1 10 9 1 11 15 13 1 10 9 1 11 2 11 2 11 2 7 13 10 11 2 11 2 11 7 11 1 9 1 12 9 7 9 2
129 10 9 0 13 16 10 9 4 13 10 9 16 13 1 10 10 9 1 10 9 1 13 10 9 1 9 0 1 9 2 3 15 1 10 9 15 13 0 3 2 1 15 10 9 1 9 15 13 1 10 9 1 10 9 2 13 3 10 9 2 15 16 13 10 0 9 0 16 13 10 9 1 10 9 1 9 1 10 13 10 9 2 13 13 2 10 9 9 1 9 1 10 9 7 10 9 2 16 13 10 9 16 13 10 9 1 10 13 1 9 1 10 9 0 10 9 0 1 13 15 9 7 9 16 10 9 0 13 2
22 1 9 2 10 9 0 13 10 9 2 13 10 9 0 1 10 9 1 1 10 9 2
59 1 10 12 9 2 11 13 0 1 10 12 5 0 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
3 13 11 2
37 11 7 11 13 10 9 10 0 11 1 10 0 9 0 1 10 9 1 11 7 11 1 10 9 0 1 10 16 10 9 4 13 9 1 0 9 2
37 2 11 11 11 11 2 2 1 9 2 2 13 1 10 9 2 2 13 10 9 2 0 9 1 10 9 11 11 11 11 1 10 9 0 11 11 2
29 4 10 9 13 9 1 10 9 2 7 13 3 3 1 10 9 2 13 15 16 13 10 9 3 7 10 10 9 2
39 10 9 0 1 10 9 7 10 9 1 9 0 1 9 7 1 9 15 13 1 9 1 10 9 1 12 9 1 9 1 9 0 1 12 9 1 10 9 2
26 7 2 13 1 10 9 16 13 16 3 13 10 9 1 10 9 1 10 9 7 15 16 13 10 9 2
26 10 9 13 9 2 10 9 13 2 13 1 10 9 10 9 2 7 10 9 1 10 9 1 10 9 2
59 1 10 12 9 2 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 0 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
47 10 9 4 13 10 9 0 2 13 15 1 10 0 9 1 10 9 0 1 10 9 7 10 9 0 1 15 16 13 13 1 10 9 2 10 9 2 10 9 7 10 9 1 10 9 0 2
42 10 9 13 10 9 1 10 9 0 15 1 10 11 1 1 10 11 2 10 9 4 13 10 9 1 10 0 9 1 10 9 1 11 11 13 1 10 11 1 10 11 2
17 4 13 1 10 9 7 13 0 1 10 9 13 16 13 3 0 2
28 13 1 10 9 1 10 9 1 11 2 10 9 1 10 0 9 1 10 11 2 13 10 9 0 1 12 5 2
27 10 9 11 12 13 15 1 10 12 9 13 1 10 9 1 9 0 9 11 2 13 1 10 11 11 11 2
28 1 10 9 1 10 9 2 10 9 13 10 9 0 1 2 1 10 15 13 9 7 2 12 5 2 13 9 2
37 1 15 9 1 10 9 10 9 4 13 3 1 9 2 9 7 9 7 15 4 13 1 3 0 9 2 13 15 15 1 9 0 2 0 7 0 2
51 10 0 9 0 15 13 10 11 13 12 9 2 11 11 2 0 1 10 9 11 11 2 7 11 11 2 10 9 0 1 10 11 1 11 10 11 2 16 13 10 9 1 9 1 10 11 11 1 11 12 2
40 3 15 13 9 1 10 9 3 3 7 15 1 9 0 2 1 1 11 1 12 7 12 2 3 13 1 9 10 9 1 9 0 7 9 1 9 1 10 9 2
35 1 10 9 2 13 10 9 13 1 10 11 2 1 0 15 3 13 1 15 7 13 16 4 1 13 8 2 7 3 13 0 1 3 0 2
11 13 15 1 10 9 0 3 0 1 11 2
28 10 9 4 13 10 12 9 1 9 16 15 13 4 1 13 1 11 7 3 13 0 13 1 10 9 3 13 2
9 13 1 2 11 1 10 9 2 2
20 3 13 1 12 8 1 9 1 9 1 9 2 1 9 13 10 9 3 0 2
24 10 10 9 4 13 9 0 1 9 1 10 9 7 1 4 13 1 11 1 10 7 10 9 2
51 1 10 9 1 10 9 12 2 9 8 1 10 9 0 2 2 10 9 15 13 1 10 0 9 1 9 7 1 9 2 15 16 4 13 9 1 15 1 10 9 3 0 1 10 9 2 10 9 0 2 2
14 10 9 3 3 2 10 9 15 13 1 11 1 9 2
55 10 9 1 10 9 1 11 13 10 9 1 9 13 1 12 9 1 0 9 2 16 13 1 9 1 9 1 10 9 13 3 2 9 2 9 2 9 2 9 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 2
19 3 2 11 7 11 13 13 15 2 7 10 12 0 13 1 10 9 0 2
21 1 10 9 1 10 9 2 10 9 13 1 8 2 1 15 15 10 9 13 0 2
25 10 9 13 16 1 10 9 1 10 9 15 13 9 0 2 1 1 9 11 2 11 1 11 11 2
12 11 4 7 13 3 10 0 9 1 9 0 2
14 4 13 10 9 2 10 9 7 10 9 1 10 9 2
27 3 2 10 11 8 11 13 1 10 9 0 1 11 11 0 2 10 9 0 1 0 9 1 9 7 9 2
36 2 3 13 1 1 10 9 1 16 10 9 0 13 1 10 9 7 15 13 1 10 9 2 13 12 9 16 4 1 13 0 2 2 13 11 2
22 13 1 10 9 13 1 10 0 9 0 2 10 9 4 13 1 9 1 10 10 9 2
22 13 10 0 9 1 9 1 9 1 9 2 9 2 8 2 2 3 4 13 10 9 2
20 11 11 13 10 9 1 9 1 10 9 1 10 11 1 10 9 1 10 11 2
30 15 13 1 10 0 9 1 10 0 9 1 2 4 13 15 15 4 13 2 2 7 15 16 3 15 13 3 4 13 2
51 11 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 1 10 9 0 1 9 0 2 0 1 10 9 11 1 12 0 1 11 11 7 11 11 11 2 1 10 9 1 10 9 13 1 8 8 2
12 10 9 16 13 15 13 1 15 7 3 0 2
13 10 9 13 0 1 9 7 9 1 10 11 11 2
28 13 9 1 9 0 1 12 9 2 7 13 1 10 9 0 13 8 2 9 2 1 9 0 13 1 10 9 2
17 10 9 13 9 3 7 15 2 7 15 13 1 13 15 1 15 2
48 1 10 14 2 9 2 11 13 1 10 8 2 8 2 7 1 10 9 15 13 16 15 13 10 9 1 10 9 1 10 9 0 2 7 10 9 0 13 11 11 2 8 10 9 11 2 11 2
10 13 10 9 3 0 1 10 9 0 2
29 1 9 11 13 16 10 9 3 4 13 10 9 15 15 13 2 7 16 4 13 10 9 9 1 9 1 10 9 2
11 10 0 9 4 13 1 9 1 10 9 2
25 13 1 10 9 9 1 9 2 13 10 9 0 2 15 13 9 1 10 9 7 9 1 10 9 2
23 1 9 2 10 9 11 4 13 9 7 13 1 11 1 10 9 1 10 9 1 12 9 2
13 1 13 10 9 13 9 3 1 10 9 1 11 2
12 13 1 11 2 11 4 13 1 9 1 9 2
7 15 4 13 3 1 11 2
59 1 10 12 9 2 11 13 0 1 10 12 5 0 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
23 3 1 10 9 1 9 0 2 7 0 2 2 11 13 9 1 10 9 2 10 0 11 2
6 9 2 9 7 9 2
41 13 3 9 1 10 11 1 10 11 7 1 10 11 1 10 11 2 9 0 1 10 15 13 1 10 9 1 11 11 11 7 11 11 2 1 10 9 1 10 9 2
6 3 13 1 12 9 2
19 13 9 1 11 1 11 11 11 2 11 11 2 11 11 11 7 11 11 2
45 10 12 1 11 1 12 2 11 1 11 13 1 10 9 1 10 9 0 0 7 1 10 9 0 1 9 1 10 9 10 9 11 11 12 2 9 1 10 12 1 11 1 12 2 2
30 3 3 13 9 1 10 9 1 10 9 0 11 11 1 11 2 7 15 13 3 1 10 9 1 10 9 0 1 12 2
46 1 10 9 2 16 13 10 0 9 1 10 9 1 10 9 1 15 15 13 10 11 1 11 2 3 13 9 1 10 11 1 11 2 2 10 9 13 3 1 13 15 1 10 9 0 2
44 11 11 11 11 2 11 2 12 1 11 1 12 2 11 2 12 1 11 1 12 2 2 13 9 2 9 7 9 1 9 2 9 1 9 2 9 2 9 7 9 0 7 0 2
47 10 9 13 10 0 9 1 10 9 16 13 3 1 10 9 16 13 12 9 2 11 1 10 11 2 11 7 11 2 2 11 1 10 11 2 11 7 11 2 7 11 2 11 7 11 2 2
20 10 9 16 15 13 1 10 9 13 3 10 9 3 1 9 16 3 15 13 2
15 11 13 3 10 9 1 9 3 0 16 4 13 1 11 2
11 15 13 9 1 9 2 10 9 1 9 2
21 10 9 0 7 9 0 2 1 9 2 8 2 13 10 9 0 3 1 10 9 2
26 1 9 1 10 9 1 10 9 2 3 15 13 15 13 10 9 3 7 15 15 13 3 1 10 11 2
31 10 11 11 13 10 9 0 3 0 1 9 0 1 11 2 1 10 8 11 12 13 1 10 9 0 11 7 10 9 11 2
35 1 9 2 10 9 13 1 13 16 10 9 1 10 9 2 9 2 1 9 13 15 3 16 10 9 7 2 7 9 1 10 9 1 0 2
26 10 9 1 11 11 13 9 2 9 2 9 2 9 7 9 0 2 13 1 10 9 1 11 2 11 2
15 10 11 4 13 9 1 10 11 10 12 1 11 1 12 2
41 10 9 3 0 7 3 0 1 10 9 4 13 15 1 16 15 13 1 10 9 16 13 9 1 10 9 1 9 13 7 10 9 1 9 2 13 10 9 7 9 2
22 7 3 2 13 16 13 9 13 2 15 15 13 7 15 4 13 15 16 15 15 13 2
18 11 13 10 9 7 9 1 10 11 11 1 10 9 1 11 2 11 2
37 13 1 10 9 0 0 1 10 15 2 10 9 4 4 13 1 10 9 0 1 4 13 1 10 9 7 4 13 10 9 0 7 15 3 0 2 2
40 1 10 9 15 4 13 12 9 2 1 10 9 0 1 12 9 2 7 1 10 0 9 13 0 16 15 13 10 12 9 2 1 10 9 16 13 10 12 9 2
31 11 13 3 10 9 0 1 10 11 1 10 9 2 1 10 13 16 10 9 1 16 11 13 1 15 10 9 0 13 0 2
67 3 15 13 1 10 9 1 10 10 9 2 7 10 9 4 13 1 10 9 1 11 2 13 1 10 9 1 9 1 9 2 10 9 1 11 11 13 1 10 9 1 3 2 9 7 9 2 3 15 4 13 1 9 7 9 2 10 9 0 16 10 9 13 1 10 9 2
34 1 9 1 10 9 15 13 10 9 13 10 9 1 10 9 1 9 10 15 15 13 1 9 2 16 15 4 13 15 1 10 9 0 2
19 11 11 13 12 9 1 10 9 1 10 11 11 2 13 1 10 9 12 2
32 15 15 4 13 16 3 13 9 7 13 10 9 7 1 10 9 3 13 16 13 15 7 16 13 16 10 9 1 9 13 0 2
18 10 9 13 3 11 13 1 10 9 2 7 13 0 1 10 9 11 2
31 10 9 0 13 0 2 12 5 1 0 2 7 0 0 2 7 16 10 9 0 13 0 7 0 0 2 1 12 5 2 2
7 4 1 13 1 10 9 2
33 10 12 1 11 1 12 2 10 0 9 0 0 4 1 13 1 11 2 1 12 9 12 9 7 12 13 9 1 10 9 1 11 2
40 10 12 9 4 13 9 16 13 10 9 7 9 1 10 9 0 2 13 10 9 1 9 16 4 13 1 10 9 1 10 9 0 9 1 10 9 1 10 11 2
6 13 12 9 1 12 2
20 3 1 13 13 1 10 9 16 10 9 15 13 1 10 9 7 9 1 9 2
8 13 9 0 1 9 7 9 2
31 3 3 13 15 9 7 13 1 9 2 7 16 15 4 13 1 9 1 10 9 2 1 9 15 13 10 9 16 4 13 2
10 11 8 12 15 13 13 1 10 9 2
22 3 1 13 10 9 0 2 13 1 10 11 1 11 2 3 13 3 0 9 1 9 2
41 16 13 10 0 9 1 10 9 2 15 15 13 10 9 1 11 2 16 15 13 1 10 9 1 13 1 10 11 1 11 2 3 4 7 13 15 1 10 9 0 2
16 13 10 9 0 1 10 9 1 13 1 10 9 1 9 0 2
37 1 10 9 1 10 11 11 11 2 1 10 9 3 1 16 11 15 4 13 7 13 1 12 2 11 13 1 11 1 3 13 1 10 9 1 11 2
54 1 10 11 15 13 1 10 9 1 9 0 1 10 11 11 2 10 9 11 11 11 1 10 11 2 10 9 11 11 11 2 10 9 11 11 2 10 9 11 11 11 2 10 9 11 11 2 7 10 9 11 1 11 2
34 16 13 1 11 2 10 9 13 16 1 10 9 13 10 0 9 7 15 13 0 1 13 1 10 0 9 2 16 13 1 9 1 9 2
23 13 3 2 10 9 1 10 9 0 1 9 0 7 10 9 1 10 9 1 9 1 9 2
21 10 9 1 10 9 0 15 13 1 9 1 10 9 1 9 1 9 0 13 11 2
23 11 13 10 9 0 1 12 5 2 5 2 7 16 10 11 13 1 10 12 5 2 5 2
58 4 13 15 12 9 1 9 0 9 13 1 10 9 7 3 1 9 2 10 9 0 13 15 10 9 13 3 1 10 9 1 10 13 0 1 13 9 0 2 10 9 13 10 0 9 1 10 9 16 1 10 9 3 4 13 1 15 2
18 16 11 13 13 15 13 1 11 2 13 3 1 11 2 1 15 13 2
43 3 2 13 16 10 16 15 13 10 9 0 2 1 13 12 9 1 12 9 2 13 15 3 0 7 13 12 9 1 12 2 3 16 1 10 0 9 10 9 13 3 0 2
35 1 10 9 1 11 10 9 0 2 10 9 1 9 13 1 10 11 11 7 11 2 13 10 9 3 3 1 10 9 1 12 9 1 9 2
33 10 9 1 11 13 13 15 1 10 9 1 11 1 9 0 3 3 13 9 1 16 11 4 13 1 9 1 11 1 10 0 9 2
19 9 1 11 11 11 11 1 11 7 11 1 11 7 11 11 11 7 11 2
18 10 9 0 2 16 13 1 10 9 2 4 13 10 9 1 10 9 2
31 10 9 1 11 2 11 11 2 13 10 9 1 1 12 9 1 9 2 3 12 9 2 7 1 12 9 1 9 1 9 2
9 3 2 13 3 1 10 11 11 2
24 10 9 1 9 4 13 2 3 13 2 3 7 9 1 9 1 10 9 9 4 13 7 13 2
14 3 10 9 1 10 9 15 13 0 1 10 9 0 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
31 11 2 1 9 2 13 1 11 11 1 11 2 7 1 11 2 13 1 10 9 2 10 11 11 11 11 11 2 1 11 2
36 10 9 1 9 2 11 11 11 2 13 16 1 10 9 10 9 0 15 13 1 10 9 0 2 13 10 9 1 13 0 1 9 1 10 9 2
19 1 10 9 10 9 13 10 9 0 1 12 9 7 10 9 1 12 9 2
12 11 3 15 13 16 11 3 13 9 1 9 2
29 1 9 2 8 11 4 13 0 1 9 0 1 9 15 13 10 9 2 13 0 1 9 1 9 2 9 7 9 2
12 7 10 9 1 10 11 2 3 13 10 9 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
31 1 10 9 11 15 13 1 10 9 1 10 9 1 11 1 10 9 2 9 16 3 13 13 1 10 9 1 11 11 11 2
11 10 9 1 11 15 13 13 1 10 9 2
15 10 9 13 9 7 15 4 13 9 13 9 1 10 9 2
20 11 13 10 9 9 1 10 9 11 11 11 2 13 10 12 1 11 1 12 2
13 3 3 15 13 2 13 15 13 7 13 1 9 2
32 3 2 1 10 9 13 1 9 4 13 15 10 10 9 1 13 10 0 9 2 9 1 10 9 2 9 7 9 1 9 8 2
16 3 13 10 2 11 2 2 10 9 1 9 0 0 7 0 2
17 11 13 10 9 1 10 11 13 1 9 7 9 2 13 1 11 2
22 1 13 15 13 0 10 9 0 2 13 1 10 9 1 9 7 9 1 9 7 9 2
35 1 12 13 1 9 0 1 10 9 11 11 11 1 10 9 1 11 2 1 10 9 1 13 15 1 10 9 16 4 13 15 1 10 9 2
40 10 9 1 11 1 11 15 13 13 1 10 9 1 10 9 1 11 2 1 12 9 1 10 9 2 7 1 9 1 10 9 11 2 13 1 10 11 1 11 2
28 1 10 0 9 2 10 9 13 1 10 9 0 2 3 0 1 10 9 2 2 16 15 13 1 10 9 0 2
75 10 12 1 11 1 12 2 11 11 11 9 1 11 11 13 16 4 13 11 1 10 9 1 12 9 1 10 11 11 2 1 10 9 9 1 10 9 2 3 16 10 9 9 0 2 1 5 12 9 2 13 10 9 1 11 1 11 1 10 11 1 11 11 10 12 1 11 7 13 12 9 1 10 9 2
41 3 10 9 13 0 2 13 0 2 0 2 1 3 1 10 9 13 3 3 2 10 9 13 0 2 13 3 3 0 2 10 9 13 0 7 10 9 13 3 0 2
28 10 0 9 13 10 9 0 0 1 10 9 7 9 0 2 15 13 9 1 9 1 10 9 1 10 0 9 2
45 13 1 10 11 11 7 11 11 2 10 9 1 9 13 1 10 9 4 13 1 10 9 1 10 11 11 1 11 11 2 11 11 2 7 13 1 10 9 1 10 11 2 11 11 2
7 3 10 9 0 13 0 2
32 10 9 3 4 13 10 9 7 10 9 16 13 1 10 0 9 1 10 9 1 9 7 1 9 1 10 9 7 1 10 9 2
17 1 12 15 13 10 9 1 10 9 0 1 10 11 1 10 11 2
41 1 11 1 10 9 12 2 11 11 11 11 2 0 1 10 9 11 2 13 10 12 8 1 11 2 3 1 10 9 13 11 11 2 2 9 1 3 13 10 9 2
15 4 13 1 10 11 11 11 11 11 11 1 11 2 11 2
18 10 9 13 3 1 9 0 2 7 16 10 9 13 3 1 10 9 2
10 12 9 2 12 5 2 15 13 9 2
14 10 9 15 13 15 16 13 0 2 0 7 3 0 2
16 11 4 13 15 1 10 9 7 15 9 4 13 16 13 15 2
8 10 9 13 0 7 10 9 2
31 11 11 11 2 11 2 11 2 12 1 11 1 12 2 2 13 10 9 0 2 15 13 1 9 0 1 10 11 1 11 2
43 13 10 0 9 2 1 10 9 1 10 9 1 10 11 11 1 3 1 11 2 9 2 7 9 2 13 3 1 13 15 1 3 1 9 7 9 2 15 3 0 7 0 2
16 10 9 2 1 12 9 2 15 13 1 10 9 1 9 9 2
23 10 12 9 13 13 10 9 2 7 10 9 1 10 9 4 13 9 1 9 0 7 0 2
77 13 10 0 9 1 9 0 2 7 10 3 0 13 10 9 1 9 0 2 16 3 15 13 9 1 10 9 2 10 0 9 1 10 9 2 2 7 10 9 1 9 0 2 0 7 0 9 1 10 9 2 2 16 3 16 13 0 9 2 13 15 1 10 9 1 10 0 9 1 9 1 15 9 1 10 9 2
14 10 9 13 9 0 7 15 13 1 9 1 10 9 2
7 10 9 15 13 1 12 2
39 1 10 9 2 11 13 16 2 10 9 16 13 9 1 10 9 1 9 4 13 9 1 10 9 1 10 9 2 3 1 10 9 13 1 0 9 0 2 2
33 11 13 13 1 11 13 16 15 1 10 9 13 1 13 10 9 1 15 0 2 7 15 13 1 15 0 1 10 9 1 10 9 2
43 10 9 11 7 11 13 1 10 9 1 10 9 2 13 1 10 9 16 4 13 10 9 1 11 2 1 9 10 12 4 13 2 16 10 9 15 13 0 7 13 10 9 2
25 3 13 13 15 10 9 13 2 12 9 3 2 16 3 4 13 10 9 1 13 9 1 10 9 2
18 15 13 1 10 11 1 11 7 15 4 13 1 10 11 11 1 11 2
19 7 3 15 13 2 16 10 9 7 10 9 1 9 0 15 13 3 0 2
28 10 9 15 13 0 1 10 9 1 10 11 2 13 15 1 10 9 10 0 11 2 11 11 2 11 7 11 2
24 10 12 1 11 1 12 2 10 9 1 9 13 1 11 11 1 10 12 5 9 1 10 9 2
10 10 9 15 13 1 9 1 10 9 2
8 13 10 0 9 1 10 9 2
22 1 9 2 10 7 10 9 10 1 9 1 9 13 3 0 2 1 10 9 7 9 2
19 10 9 4 13 1 12 1 10 11 1 12 9 7 13 0 1 12 9 2
28 7 10 9 1 10 9 13 10 9 0 16 13 1 10 0 9 1 9 1 10 15 15 15 13 1 9 0 2
13 10 9 12 13 10 12 5 9 0 1 10 9 2
19 15 13 10 12 1 11 1 12 7 15 15 13 9 0 1 9 1 11 2
14 10 9 2 9 7 3 9 15 13 1 10 9 0 2
24 10 9 0 13 0 1 10 9 2 12 12 2 7 12 9 1 11 11 1 9 1 10 9 2
5 13 10 0 9 2
19 10 12 9 13 9 7 13 1 9 1 10 11 1 11 1 9 1 11 2
25 15 15 13 10 9 1 10 11 7 15 13 10 9 3 0 1 11 10 3 0 9 0 1 11 2
65 10 9 13 0 1 13 7 1 10 9 1 10 9 1 10 9 7 1 10 9 15 13 1 10 9 12 7 10 9 15 13 1 10 9 12 2 10 9 13 0 1 10 9 1 10 9 1 11 2 1 9 1 10 9 12 2 16 15 13 1 9 1 0 9 2
25 9 13 10 9 13 1 11 11 1 13 15 1 10 9 0 1 9 0 1 11 7 0 1 11 2
35 10 9 16 13 1 11 7 13 15 1 10 9 1 10 9 0 2 13 0 9 1 10 9 1 10 9 7 3 1 10 9 0 11 11 2
13 10 9 13 1 11 2 10 12 1 11 1 12 2
16 13 10 9 0 16 15 13 1 10 9 1 10 9 1 11 2
22 1 9 2 10 9 4 13 1 10 9 1 10 13 15 2 0 2 1 10 0 9 2
45 10 9 2 15 3 15 13 1 9 7 9 0 2 15 15 13 0 9 7 9 1 10 9 2 2 13 1 13 15 1 9 3 0 2 7 2 1 15 2 3 0 1 10 9 2
38 11 11 4 1 13 1 10 9 0 13 16 9 1 11 1 11 13 16 10 9 1 9 13 9 1 9 16 1 10 9 1 10 9 15 13 1 9 2
52 10 9 10 9 15 4 13 3 7 3 3 2 10 9 15 15 4 13 3 7 10 9 1 10 9 13 10 9 7 2 3 7 13 10 0 9 1 10 9 2 15 13 10 9 1 10 9 2 2 0 9 2
46 15 13 9 1 10 9 0 7 1 0 9 7 0 2 1 9 7 1 9 2 1 10 9 0 1 10 11 2 1 13 15 1 10 9 1 10 9 1 10 15 15 4 1 9 2 2
26 16 10 9 0 13 10 9 2 1 9 10 9 13 9 1 10 11 11 7 10 9 1 10 11 11 2
39 3 15 13 13 1 12 9 10 11 11 1 11 1 10 9 11 11 7 10 11 11 1 10 9 11 11 1 15 13 10 9 1 12 1 10 9 1 11 2
17 10 0 9 13 10 12 5 9 1 10 11 11 1 11 1 12 2
17 10 9 3 13 0 1 9 1 4 13 1 10 9 11 11 11 2
39 1 10 9 9 13 10 9 1 15 2 7 15 9 13 16 15 13 1 10 9 2 3 7 13 0 10 9 16 13 10 9 2 1 10 9 1 10 9 2
31 10 9 15 13 1 9 1 1 9 1 10 11 2 3 10 9 4 13 1 10 11 2 13 10 9 16 13 9 7 9 2
33 10 11 11 3 15 13 11 2 11 7 11 2 10 0 9 1 9 13 1 10 9 7 13 1 9 1 9 0 1 11 7 11 2
15 11 11 13 10 12 1 11 1 12 1 10 11 1 11 2
53 10 9 2 9 2 13 9 0 1 10 9 7 1 10 9 16 3 13 1 13 15 2 7 16 10 9 13 3 1 10 0 9 1 10 11 11 1 11 2 10 9 0 2 9 1 11 7 1 11 1 10 9 2
26 10 0 9 0 7 0 2 15 13 13 10 9 1 11 7 13 16 13 9 1 0 9 0 1 11 2
14 7 10 9 15 13 1 15 15 3 13 2 10 11 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
40 3 10 9 1 9 4 4 13 7 13 1 3 10 10 9 0 2 1 11 2 2 7 10 9 1 10 9 1 11 2 1 11 2 11 11 7 11 11 2 2
14 10 9 2 13 1 8 7 9 0 13 10 0 9 2
17 1 10 9 1 11 2 11 3 13 10 9 0 1 10 9 0 2
54 7 10 8 9 7 8 9 13 3 3 2 15 13 10 0 9 1 11 11 1 9 1 10 9 7 9 1 9 1 9 9 0 7 0 1 10 9 1 9 2 15 1 10 9 1 13 10 9 13 10 9 1 9 2
11 13 10 9 16 13 10 12 9 1 9 2
36 10 0 9 1 10 9 2 10 12 5 0 1 15 1 10 9 1 9 0 2 13 13 1 12 8 1 10 9 16 15 13 1 10 0 9 2
15 10 9 1 9 7 9 4 13 0 1 9 0 7 0 2
21 3 2 15 13 10 9 1 11 11 16 8 12 9 1 9 1 9 1 10 9 2
42 10 9 2 1 12 9 2 13 0 2 1 10 9 2 1 10 11 11 7 13 1 13 2 1 10 9 7 10 9 2 1 10 9 1 10 9 0 1 10 0 9 2
45 13 0 16 10 9 13 0 2 7 4 13 15 1 9 2 0 2 2 1 10 9 1 9 2 0 2 2 1 9 2 7 1 10 9 7 10 9 1 9 2 0 1 9 2 2
134 13 10 9 1 13 15 1 9 1 10 9 1 10 9 11 7 10 9 1 9 7 13 15 16 10 12 1 11 1 10 9 1 9 2 1 10 9 1 10 9 1 10 12 9 1 11 11 2 10 9 1 10 9 11 2 1 9 1 10 9 1 9 4 13 10 0 9 1 9 1 9 1 10 9 0 1 10 9 11 2 16 13 1 10 9 1 9 1 10 9 0 0 2 0 7 0 2 3 7 0 9 2 9 2 9 1 9 1 10 0 9 16 13 10 9 1 9 1 10 9 2 9 0 2 9 0 7 9 0 1 10 11 11 2
47 10 9 1 10 9 1 9 2 7 3 10 10 9 2 1 10 11 0 1 11 2 13 1 10 9 11 11 2 7 11 1 10 11 2 2 13 1 10 11 11 2 2 4 13 1 11 2
11 15 13 7 15 13 1 10 9 7 9 2
22 10 9 4 13 1 9 1 10 9 0 7 4 4 13 1 10 9 2 9 7 9 2
41 1 10 9 2 13 10 9 0 16 13 13 10 9 0 1 10 0 9 1 10 9 11 2 9 16 15 13 3 1 10 9 0 7 9 0 16 13 10 0 9 2
33 13 3 0 1 10 9 2 13 10 0 9 1 9 7 9 0 2 9 2 9 2 9 7 9 1 10 9 1 9 7 10 9 2
18 10 9 13 16 10 9 13 15 1 15 13 2 15 15 13 10 9 2
49 9 0 7 1 9 0 2 9 7 11 2 1 0 9 16 9 1 9 1 12 9 0 2 11 11 1 11 2 1 10 15 3 13 3 7 10 9 1 10 9 2 7 10 1 11 11 1 11 2
17 11 11 8 2 11 2 12 1 11 1 12 2 13 10 9 0 2
12 10 9 13 1 0 7 0 1 9 7 0 2
22 11 11 2 11 11 2 2 0 9 1 11 11 2 11 11 2 2 3 13 13 9 2
23 1 10 9 13 11 10 9 0 2 1 12 10 9 13 3 10 9 0 1 2 11 2 2
35 10 9 1 11 2 11 11 11 2 15 13 1 16 1 10 9 1 10 9 2 13 10 9 1 10 9 1 12 9 1 10 3 9 9 2
26 1 10 9 1 10 9 4 13 1 9 9 7 11 11 13 10 9 1 10 0 9 1 11 11 12 2
6 3 13 9 1 9 2
46 3 2 1 10 9 13 1 10 9 2 15 4 1 13 10 9 1 12 9 16 4 1 13 13 10 12 5 1 10 9 13 1 10 9 2 1 9 1 9 1 10 9 1 10 9 2
28 7 10 9 3 10 12 9 0 2 15 4 13 1 9 7 1 9 2 2 0 1 13 0 9 1 10 9 2
33 16 13 1 10 9 2 10 9 13 10 9 0 1 10 0 9 7 15 13 13 1 15 9 1 10 9 2 1 13 1 10 9 2
26 1 9 1 4 13 1 9 1 10 9 0 2 11 13 10 0 9 0 1 13 15 3 1 10 9 2
16 10 9 13 10 0 9 1 10 9 7 10 9 1 10 9 2
28 10 12 5 1 10 12 9 1 9 0 13 1 10 9 2 10 9 1 9 1 10 12 5 1 13 12 9 2
14 3 4 13 9 1 0 9 0 1 9 1 10 9 2
16 3 1 10 12 5 1 10 9 13 1 10 9 1 9 0 2
18 11 12 13 1 13 3 3 12 9 7 1 12 13 9 1 10 9 2
31 15 13 16 2 1 10 9 1 10 9 1 12 2 10 12 5 1 10 9 0 13 0 2 16 7 10 12 5 13 0 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
29 4 13 11 2 11 11 2 11 11 7 11 11 2 3 16 10 9 0 13 1 9 1 11 2 11 7 8 11 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
34 13 10 9 1 12 9 2 10 9 0 1 12 9 5 7 10 9 0 1 12 8 2 8 1 12 9 1 10 9 1 10 9 11 2
18 10 0 9 13 10 9 11 1 11 1 9 1 11 11 7 11 11 2
23 10 9 4 13 1 0 9 1 11 11 2 11 11 2 11 11 2 11 11 2 1 15 2
26 1 10 9 1 9 7 9 1 10 9 1 12 2 10 9 16 13 1 10 9 12 13 10 0 9 2
16 10 9 4 8 2 13 1 10 9 0 11 7 10 0 11 2
69 3 2 10 9 0 1 10 9 2 16 10 9 4 13 16 10 9 1 10 9 1 10 9 13 12 9 1 9 2 16 10 9 16 15 13 1 10 9 13 0 2 1 12 9 1 9 1 10 9 2 7 16 10 9 13 10 9 3 0 1 10 9 0 1 3 1 12 9 2
23 15 13 15 7 3 13 10 9 1 9 16 13 2 13 3 0 7 3 15 4 7 13 2
57 15 13 1 9 0 2 13 15 12 9 0 0 1 9 7 9 7 13 1 9 10 9 0 2 2 16 1 11 13 3 9 2 7 13 3 1 9 0 2 13 10 9 0 1 10 9 7 13 15 1 13 1 2 10 9 2 2
33 10 9 13 0 1 9 1 10 9 7 15 15 13 1 10 9 1 10 9 1 10 9 1 9 16 13 1 10 9 1 10 11 2
27 10 9 13 16 9 1 9 1 10 8 4 13 7 13 2 16 10 15 4 13 1 9 13 10 9 0 2
18 1 11 15 4 13 3 1 10 9 0 7 3 3 1 10 9 0 2
31 10 9 1 10 9 0 2 11 11 11 11 2 15 13 0 1 13 9 1 13 10 9 1 10 8 16 2 4 13 2 2
24 10 9 15 13 1 10 9 2 7 10 9 0 13 10 9 9 1 10 9 3 1 10 9 2
13 10 9 15 13 3 3 1 10 9 16 13 13 2
12 1 0 2 3 15 13 1 13 1 9 0 2
50 2 10 9 13 10 9 1 9 16 13 1 9 1 10 11 11 1 11 2 7 13 3 1 10 9 1 10 9 7 13 9 1 10 9 1 10 9 1 10 9 2 2 13 11 11 2 9 1 9 2
44 10 9 1 10 9 1 11 2 12 2 13 10 9 1 10 9 1 10 9 2 7 1 10 9 0 1 10 9 0 2 13 1 10 9 1 11 2 13 1 10 0 9 2 2
31 3 2 13 10 9 13 11 11 2 9 1 10 9 16 13 1 11 2 7 1 9 2 11 11 2 9 0 1 10 9 2
59 1 10 12 9 2 11 4 0 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
11 10 9 1 9 15 13 10 12 1 11 2
17 1 10 9 13 10 9 0 7 15 13 1 10 9 1 9 0 2
32 10 9 0 3 15 13 1 13 1 10 9 13 15 1 13 1 10 9 7 13 3 10 9 1 10 9 13 15 1 10 9 2
34 11 13 3 10 0 9 0 1 9 0 2 1 3 1 12 9 1 9 1 9 2 9 0 1 15 1 9 1 11 2 11 7 11 2
24 1 10 9 10 9 0 1 11 13 1 10 9 1 10 9 7 3 3 1 10 9 1 9 2
31 3 15 13 3 9 0 2 7 9 3 0 7 15 16 3 13 9 4 13 10 9 1 13 15 3 9 1 10 9 0 2
14 11 1 11 2 11 2 11 7 11 1 9 2 11 2
27 15 15 13 1 11 15 15 4 13 1 10 9 16 13 15 1 10 9 0 7 13 10 9 2 11 2 2
5 4 13 12 9 2
26 10 0 9 2 3 15 13 1 11 2 1 9 1 10 3 9 2 11 11 13 7 13 13 10 9 2
15 11 13 10 9 8 16 1 10 9 15 4 13 11 11 2
26 13 2 13 7 13 11 2 13 1 10 9 1 11 7 1 12 9 4 13 2 1 9 1 9 0 2
53 1 9 1 10 0 9 2 10 9 1 11 10 11 13 10 9 1 0 9 0 1 10 9 1 10 13 10 0 9 1 10 12 9 0 1 11 2 11 7 11 2 10 9 1 10 9 15 13 3 9 1 9 2
38 11 11 13 13 15 1 10 9 1 11 2 13 1 10 9 1 9 1 10 11 11 1 10 11 1 11 13 0 9 1 10 15 15 13 1 10 9 2
35 1 10 9 13 10 9 1 9 1 0 9 13 1 10 0 12 1 11 1 12 2 9 1 10 16 15 13 1 9 1 9 1 0 9 2
38 1 9 0 2 1 10 0 9 2 15 13 10 0 9 0 3 13 10 11 1 10 11 1 11 2 11 11 7 11 2 0 9 1 10 11 1 11 2
15 3 13 16 3 15 13 3 9 16 13 9 1 10 9 2
60 11 2 9 0 1 10 11 1 11 2 13 8 9 1 9 7 3 13 9 1 10 9 1 9 2 9 7 9 7 9 1 10 9 1 9 7 9 2 1 9 7 9 0 2 1 9 2 9 7 9 2 1 9 7 9 7 1 9 9 2
47 1 15 2 1 9 1 10 9 0 2 10 9 2 15 13 1 10 9 1 10 9 0 2 13 2 3 0 2 0 1 10 0 9 2 1 10 3 1 10 9 16 13 1 10 9 0 2
37 1 10 9 13 10 9 1 10 0 9 1 9 0 2 10 9 1 11 11 2 11 11 11 11 2 2 13 1 10 9 11 12 1 11 1 12 2
25 7 13 1 10 9 0 9 0 9 12 2 10 12 9 0 12 7 12 7 15 0 12 7 12 2
14 15 1 10 9 3 0 13 10 9 0 11 11 11 2
11 10 9 1 11 15 13 0 1 10 9 2
30 1 9 2 13 10 0 9 2 16 5 13 3 1 10 9 0 7 16 4 13 10 0 9 0 1 10 10 11 11 2
25 11 11 2 10 9 0 2 13 10 9 1 9 1 10 9 2 13 1 9 7 9 10 0 9 2
7 13 10 9 1 10 9 2
18 10 12 9 2 11 7 11 2 13 1 13 10 9 1 10 9 11 2
43 1 10 11 1 10 11 1 10 11 11 2 10 9 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 4 1 9 0 7 2 12 5 2 12 5 5 13 9 2
38 10 9 3 0 13 1 12 9 1 9 7 10 9 1 1 12 9 2 7 15 3 0 13 16 13 15 3 1 12 9 1 9 7 13 10 12 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
21 11 13 15 1 10 3 10 9 15 10 9 0 13 1 10 9 0 1 10 9 2
21 3 13 1 10 0 9 1 8 2 8 1 11 2 1 0 9 1 9 7 9 2
17 10 9 13 3 3 10 9 3 1 10 0 9 1 1 10 9 2
41 10 11 13 1 9 10 11 1 10 9 10 9 1 11 2 13 1 0 1 10 9 3 13 0 10 9 1 10 9 0 11 11 2 3 1 10 9 1 10 9 2
36 9 2 1 10 9 11 2 13 2 2 2 9 1 10 15 10 9 2 1 10 9 1 10 9 7 3 3 2 15 13 10 9 1 10 9 2
14 10 12 5 1 10 9 13 9 7 9 1 10 9 2
30 11 3 4 13 9 1 10 9 11 2 1 12 15 13 10 9 1 9 1 10 9 1 9 1 10 9 7 9 0 2
16 1 12 9 15 13 16 1 11 13 10 0 9 1 10 9 2
32 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 13 10 9 0 1 9 16 3 15 13 1 10 9 1 9 0 2
23 10 9 13 1 10 9 1 10 11 2 13 1 10 9 1 9 2 7 13 1 10 9 2
23 13 1 11 11 1 10 9 16 15 13 16 13 10 9 2 13 10 9 1 10 12 11 2
7 10 0 9 13 11 11 2
40 10 11 11 15 13 1 12 9 15 1 10 9 0 7 1 11 11 2 1 12 9 10 11 0 2 1 13 1 3 7 1 9 1 13 1 10 12 1 11 2
28 10 9 0 4 13 1 9 13 1 11 1 11 2 1 11 16 13 10 11 1 11 1 10 9 0 1 11 2
22 1 9 1 10 9 2 10 9 13 10 9 1 10 9 0 10 12 1 11 1 12 2
34 1 11 1 10 9 0 15 13 16 11 13 10 9 0 13 11 1 15 10 11 15 13 10 9 7 13 10 9 1 11 1 1 9 2
16 9 13 1 10 9 1 10 9 0 2 3 13 9 3 3 2
19 1 12 10 9 13 10 9 1 9 1 5 12 1 5 12 1 10 9 2
52 10 9 15 4 1 10 9 1 0 9 7 9 0 1 10 9 1 9 0 2 13 1 10 9 1 10 9 1 9 0 16 13 9 1 9 2 1 9 16 13 10 9 1 9 0 13 1 10 9 1 9 2
41 11 2 1 9 11 2 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 1 11 11 2 1 10 9 1 11 7 9 1 11 2 11 2 1 2 11 2
4 13 12 9 2
21 1 9 15 13 10 9 1 10 9 1 10 9 13 1 11 1 12 2 13 3 2
20 13 10 9 0 2 11 2 7 15 13 1 10 12 1 11 1 10 0 9 2
31 1 9 2 1 10 9 2 3 1 11 2 1 13 15 13 1 11 2 9 0 11 11 2 2 10 9 1 11 7 11 2
23 10 9 11 13 13 15 0 1 10 9 0 16 3 3 13 1 10 9 1 10 10 9 2
16 15 13 10 9 0 13 1 11 11 1 10 9 7 10 9 2
29 10 9 13 9 1 11 2 7 3 1 10 9 4 13 1 10 9 1 11 2 3 13 9 1 9 0 7 9 2
39 1 11 11 2 10 9 1 9 13 15 16 13 10 9 0 7 1 9 1 10 9 2 1 10 9 0 1 9 2 2 1 10 16 11 13 3 3 2 2
14 10 9 8 0 16 13 1 10 9 13 15 7 0 2
13 10 9 0 13 0 2 13 15 7 13 15 0 2
76 10 0 9 1 10 9 2 13 1 10 9 1 11 2 13 1 10 9 7 1 10 9 2 3 2 13 11 1 13 10 9 0 1 9 7 13 10 9 1 10 9 1 9 1 13 9 1 10 9 1 10 9 2 15 3 13 0 1 10 9 7 9 1 9 2 13 16 15 13 1 10 9 1 15 2 2
54 10 9 1 11 2 16 4 13 13 12 9 1 13 1 10 9 1 10 9 2 13 16 1 15 15 15 13 2 10 9 16 4 13 1 10 9 1 11 10 9 0 1 13 10 9 12 1 10 9 3 13 1 9 2
19 11 11 13 16 16 11 11 13 9 1 11 2 4 13 16 3 4 13 2
13 13 0 13 16 15 3 13 12 9 1 10 9 2
48 10 0 9 1 0 9 11 11 2 10 9 7 0 9 1 11 13 10 9 0 1 9 0 13 3 1 10 9 1 11 11 1 10 11 1 10 9 1 11 1 11 2 1 10 9 1 11 2
46 10 0 12 9 1 10 9 13 3 0 7 15 13 13 3 1 10 9 8 0 1 10 9 0 2 1 10 0 11 13 1 10 9 1 10 9 7 10 9 3 1 10 9 8 0 2
18 11 11 10 11 13 10 9 0 1 10 11 11 8 11 2 12 2 2
53 1 9 13 9 1 0 9 0 13 1 10 9 16 13 16 10 0 9 13 1 10 11 2 7 3 13 9 1 10 9 0 1 15 2 7 16 10 9 1 9 1 10 9 13 3 9 1 13 10 9 7 9 2
30 10 9 0 11 2 11 11 5 11 11 2 11 2 13 10 9 2 1 10 15 13 12 5 7 10 9 0 12 5 2
21 1 10 9 1 10 9 2 15 15 4 13 9 2 10 9 16 4 13 10 9 2
23 11 13 10 9 0 7 13 10 9 1 10 0 9 1 7 10 9 11 13 1 12 9 2
75 10 9 11 11 2 13 1 10 9 2 9 7 9 7 15 13 1 12 0 1 10 11 1 11 11 2 3 13 10 9 1 9 11 1 10 11 2 10 9 11 11 13 10 9 2 7 10 9 11 11 11 15 13 1 10 9 0 11 11 11 1 11 11 2 12 9 1 11 2 1 9 1 10 9 2
34 10 9 3 0 1 10 9 13 10 9 0 13 1 11 11 2 3 13 1 11 2 11 2 7 10 11 2 13 3 11 2 11 2 2
48 11 11 1 11 4 13 15 1 10 9 1 11 11 2 3 3 1 4 13 15 1 10 0 9 1 10 11 11 1 11 2 7 16 4 15 13 1 10 9 2 13 10 9 1 10 9 0 2
23 10 11 13 1 15 10 9 11 2 11 2 16 3 13 9 11 2 11 7 11 2 11 2
42 10 12 1 11 1 12 2 1 10 9 0 1 10 9 0 2 11 13 1 10 9 11 1 10 9 1 9 7 13 10 9 1 9 1 10 9 7 9 1 10 9 2
29 10 9 13 1 10 9 0 3 0 2 1 10 9 1 11 11 1 9 2 11 11 1 9 7 11 11 1 9 2
13 10 9 13 9 1 10 11 12 8 8 1 12 2
12 10 11 1 11 9 13 1 11 11 1 12 2
30 1 9 2 10 9 15 13 0 16 15 13 16 4 13 3 12 9 1 10 9 7 10 9 15 4 13 1 10 9 2
15 10 9 15 13 10 9 1 9 0 1 10 9 11 11 2
21 15 13 15 1 11 15 3 4 13 10 9 2 7 15 13 2 8 8 8 8 2
25 3 2 15 13 0 1 10 9 13 1 10 9 1 10 9 0 2 7 16 13 9 1 10 9 2
23 10 9 0 4 13 1 10 9 7 9 16 13 10 9 11 11 7 11 2 11 2 11 2
35 1 12 11 13 10 9 1 10 9 11 1 11 3 13 1 11 1 11 11 7 13 1 11 11 7 11 11 1 10 9 0 1 11 11 2
25 15 15 13 1 9 1 9 1 13 10 9 1 10 9 1 10 9 13 10 8 1 10 9 0 2
22 11 13 10 9 13 1 10 9 1 11 1 10 9 1 10 9 11 2 11 7 11 2
81 1 10 9 2 10 9 0 3 3 15 13 0 1 10 0 9 0 2 13 1 10 9 2 3 1 9 2 3 7 0 2 1 0 9 1 9 7 9 2 3 7 1 10 9 1 0 9 7 9 0 2 7 16 3 10 9 0 2 0 15 13 1 10 0 9 2 10 9 1 0 2 13 1 9 1 10 9 1 10 9 2
9 4 13 15 0 3 1 12 9 2
40 1 9 2 10 9 4 13 1 9 0 2 1 9 16 2 1 10 9 11 8 11 13 2 2 11 13 10 9 0 1 10 9 0 1 13 15 13 10 9 2
36 15 1 10 0 9 16 13 1 10 9 1 11 13 13 10 9 1 13 9 1 0 9 13 9 1 0 9 2 1 0 8 7 8 2 9 2
7 1 12 13 10 9 0 2
16 11 11 13 10 9 1 10 9 1 10 9 1 11 2 11 2
27 13 9 7 2 13 1 10 9 2 13 1 9 0 1 10 9 13 1 10 9 1 11 7 11 11 11 2
15 15 13 3 1 0 9 2 9 1 9 7 3 9 0 2
37 11 4 13 1 10 9 0 11 2 16 10 9 0 9 0 1 13 10 9 1 12 2 1 10 9 1 13 13 1 10 9 1 10 9 1 11 2
36 16 1 10 9 2 10 9 1 11 7 11 13 1 13 10 9 0 1 10 9 2 3 4 13 16 4 13 9 0 1 11 1 10 12 9 2
20 10 9 1 11 2 11 2 13 15 1 10 12 9 1 10 9 0 1 11 2
57 11 11 13 10 9 1 9 1 10 9 1 9 0 11 11 2 13 1 12 7 16 13 10 9 1 10 9 1 11 2 12 2 2 11 2 12 2 2 10 11 11 2 11 2 12 2 7 10 11 11 2 11 11 2 12 2 2
81 10 9 9 1 10 0 11 11 2 13 1 10 9 1 11 2 13 10 9 11 2 10 9 15 13 1 10 0 9 1 9 1 2 12 7 2 12 5 8 1 10 9 13 3 1 13 15 1 10 9 1 9 1 12 5 8 1 10 0 9 15 13 10 9 1 9 9 1 10 9 1 9 0 7 10 9 1 9 7 9 2
9 13 15 13 1 10 9 2 11 2
33 11 11 2 11 2 12 1 11 1 12 2 11 1 11 2 12 1 11 1 12 2 2 13 10 9 0 2 9 1 10 11 11 2
28 11 3 13 16 15 4 13 3 16 13 16 15 13 1 11 2 15 13 16 10 9 13 0 7 11 4 13 2
25 10 9 1 10 15 15 13 1 11 13 1 9 1 10 9 2 13 3 7 3 12 9 1 9 2
50 10 9 1 9 12 13 1 11 1 10 9 1 10 11 2 13 10 9 0 1 11 11 2 11 2 1 10 9 1 9 2 2 13 1 10 3 12 9 2 9 1 9 7 9 1 9 7 9 0 2
56 9 1 9 13 10 11 1 10 9 0 1 11 1 10 9 1 12 9 1 10 11 8 11 2 1 10 9 1 10 9 1 10 11 1 10 11 2 11 11 7 11 11 2 9 0 1 10 9 1 12 2 4 13 10 9 2
29 1 10 11 11 2 10 12 0 9 0 2 11 2 11 7 11 2 13 10 2 11 1 11 2 10 12 1 11 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
16 13 10 0 9 1 13 10 9 1 9 2 1 11 1 12 2
19 3 4 13 1 11 1 10 9 8 1 10 11 11 2 3 13 12 9 2
23 13 9 1 10 9 0 1 11 1 10 9 2 3 9 1 10 11 1 9 0 1 11 2
48 1 12 7 12 9 1 9 2 10 9 13 1 9 1 10 9 0 2 1 9 1 16 10 9 4 13 9 1 9 1 0 9 0 1 10 9 1 10 0 9 1 9 0 1 11 1 12 2
68 10 9 9 1 10 11 11 1 10 9 12 2 12 4 13 9 7 3 4 13 3 10 9 16 4 13 15 1 10 9 7 1 10 11 11 13 10 9 16 3 13 9 1 10 0 9 1 13 10 9 1 10 9 2 1 15 10 11 2 11 7 15 3 1 10 0 9 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
36 11 11 13 13 2 3 7 3 13 13 3 9 3 13 1 10 9 7 1 10 9 0 2 1 15 13 1 13 15 1 10 9 1 10 9 2
38 10 0 9 0 13 1 10 9 13 10 9 1 10 9 7 9 1 10 9 2 3 9 1 10 9 13 1 10 9 1 10 9 7 1 10 9 0 2
43 3 0 2 13 10 9 1 10 9 11 1 10 9 1 10 9 1 10 9 7 1 10 9 1 10 9 2 16 1 10 9 0 13 9 0 1 10 0 9 1 11 11 2
19 13 1 10 0 9 2 3 0 1 9 7 3 15 13 7 13 10 9 2
34 15 1 15 4 13 1 13 7 10 12 1 11 10 11 1 11 11 11 15 13 1 11 7 13 2 2 2 15 4 1 13 7 13 2
9 13 9 1 10 9 0 11 11 2
17 1 4 13 9 10 12 1 11 1 12 2 13 1 10 9 0 2
13 1 10 9 13 10 10 9 1 11 13 1 11 2
13 11 13 1 11 2 11 10 12 1 11 1 12 2
20 11 11 4 13 1 11 11 11 7 13 1 11 11 11 11 11 12 2 12 2
45 10 9 0 4 13 16 10 9 13 3 0 1 10 9 0 7 13 15 3 9 1 10 9 1 9 0 1 13 10 9 1 9 7 9 7 10 16 15 13 1 13 7 13 9 2
32 10 9 7 10 9 1 9 2 9 2 9 2 9 3 2 13 10 9 1 9 7 1 9 2 16 15 13 13 1 10 9 2
18 11 13 1 10 11 7 3 13 16 15 13 10 9 0 1 10 11 2
19 10 10 9 2 10 0 2 13 10 9 3 0 1 10 9 2 10 11 2
11 1 12 4 13 9 0 1 10 12 11 2
33 3 10 11 11 11 4 13 1 13 0 9 2 1 9 1 9 9 2 9 2 16 13 16 15 13 0 0 1 15 7 10 9 2
28 3 10 13 3 1 10 9 7 3 1 10 9 3 13 10 9 1 10 9 1 13 15 2 1 9 3 0 2
36 10 9 1 10 9 13 0 7 13 1 0 7 0 9 7 15 13 1 12 9 1 10 15 10 15 13 9 13 1 15 9 1 10 9 0 2
48 11 13 1 10 9 1 10 11 11 12 10 15 15 13 1 9 10 12 1 11 1 10 11 2 11 11 2 3 13 1 9 1 0 9 1 13 1 13 10 9 1 11 11 2 0 11 11 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
40 10 9 2 16 13 9 1 10 9 13 15 1 13 1 15 2 15 13 3 0 1 10 9 1 9 1 10 9 1 11 7 1 10 2 9 0 1 9 2 2
30 1 15 2 13 2 13 7 13 1 16 10 9 13 10 9 1 10 9 2 9 1 10 9 1 9 0 1 10 9 2
26 3 2 13 9 0 0 1 10 11 11 2 4 13 1 10 11 11 1 10 11 1 10 11 1 12 2
11 13 10 9 0 1 10 9 1 10 9 2
39 2 13 16 4 1 13 3 16 10 0 9 1 11 3 15 13 2 2 13 11 11 2 9 1 10 11 11 1 11 11 7 15 1 10 9 1 10 9 2
25 10 9 0 2 1 9 13 10 9 1 10 9 2 15 13 10 9 16 1 15 3 4 1 13 2
14 13 12 9 16 15 13 10 11 1 10 9 1 11 2
20 10 9 2 1 15 13 1 10 0 9 2 4 4 13 1 10 9 1 10 8
14 11 13 10 12 1 11 1 12 1 11 11 2 11 2
16 13 10 0 9 1 13 15 1 12 9 7 1 12 9 0 2
35 1 9 0 1 10 11 1 11 2 13 10 9 0 1 10 9 2 1 10 13 1 10 12 9 1 9 1 10 9 1 10 11 11 11 2
24 16 11 11 13 10 9 0 2 11 15 13 1 9 1 10 11 1 11 7 10 11 1 11 2
11 1 10 9 2 10 9 15 13 1 9 2
38 3 2 13 10 9 13 1 11 12 1 12 1 10 15 15 13 10 9 1 10 9 11 11 12 1 11 7 11 2 9 1 10 9 11 11 1 11 2
42 15 1 10 9 4 4 13 2 1 11 11 2 11 2 4 3 13 10 9 0 2 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 3 1 11 11 2
31 13 12 9 1 10 11 2 13 10 9 1 15 10 9 2 10 9 8 2 1 10 15 13 12 9 7 12 9 1 9 2
28 11 11 11 13 10 9 13 1 10 9 0 2 1 10 11 11 11 1 11 1 12 2 7 13 3 1 11 2
10 12 9 0 13 1 10 9 10 11 2
12 15 13 7 1 10 9 0 2 11 15 13 2
20 1 9 1 10 9 2 10 9 15 13 1 10 9 0 7 13 1 10 9 2
22 10 9 0 13 1 10 0 9 1 10 0 9 1 10 9 7 3 1 9 1 12 2
22 15 13 16 10 9 13 1 15 3 1 10 12 9 16 15 13 1 9 1 0 9 2
24 11 4 13 1 10 9 1 11 2 11 11 2 7 11 4 13 9 1 10 9 1 10 11 2
41 1 10 9 2 10 9 1 10 9 13 2 0 3 1 10 9 2 2 1 15 15 13 0 16 10 9 13 1 10 9 0 1 10 9 2 9 2 9 7 9 2
30 1 9 2 10 9 13 10 3 13 1 10 15 16 13 1 10 9 1 10 9 2 1 15 1 11 2 11 7 11 2
35 1 0 9 2 10 9 1 13 3 4 13 15 0 1 10 9 3 0 2 13 1 10 11 11 2 7 13 1 10 0 9 9 1 11 2
29 2 13 10 9 16 4 1 13 0 1 10 9 1 9 1 10 9 7 3 4 13 15 1 10 9 0 16 13 2
20 10 9 2 11 11 2 13 1 10 9 1 10 9 1 11 1 11 11 11 2
15 10 9 13 3 10 9 1 10 9 0 1 10 10 9 2
57 15 1 10 9 3 0 7 3 0 13 10 9 1 10 9 11 16 1 7 13 1 10 9 3 4 4 1 13 12 9 0 7 16 15 13 10 0 9 1 9 1 10 9 0 2 7 16 13 10 9 1 13 1 10 11 0 2
36 3 11 4 13 16 10 9 1 10 11 13 2 0 2 7 15 4 13 2 1 9 2 1 10 0 9 1 9 1 9 1 10 9 13 3 2
34 7 0 2 10 15 13 13 15 9 1 15 0 2 7 7 3 15 4 13 15 1 10 9 0 1 10 9 2 1 10 15 15 13 2
13 10 9 1 11 2 11 13 9 1 9 1 12 2
13 10 9 1 11 13 13 1 11 7 2 1 11 2
12 11 11 11 11 13 10 9 1 10 9 12 2
47 10 9 0 11 11 11 11 13 0 1 10 12 9 13 1 10 9 16 13 10 9 1 10 11 12 1 11 1 10 0 9 1 10 9 1 10 9 1 8 2 9 7 9 0 2 11 2
28 1 11 7 11 1 12 2 13 1 11 11 3 1 13 1 10 9 1 11 8 8 1 9 1 11 1 12 2
23 3 3 1 10 0 9 15 13 13 10 9 1 9 1 10 9 7 1 9 0 1 11 2
60 1 3 12 9 1 10 9 15 4 13 10 11 12 1 11 1 12 1 10 9 1 10 9 11 11 1 11 1 12 9 1 9 1 0 9 16 15 13 1 10 9 1 11 7 15 13 12 9 2 10 9 13 10 9 1 13 1 10 11 2
34 10 12 1 11 2 15 13 10 9 0 1 10 9 1 11 11 11 2 11 12 2 1 10 9 7 9 1 10 9 0 1 10 9 2
12 10 9 13 10 9 7 13 0 1 10 9 2
28 0 1 0 10 9 16 15 13 9 7 9 2 1 9 2 16 13 2 0 2 2 3 13 10 9 7 9 2
17 15 2 1 11 11 2 1 10 9 1 9 13 15 16 3 13 2
8 13 10 9 1 11 7 11 2
32 10 9 4 13 1 10 12 1 11 1 12 1 11 2 10 12 1 11 1 12 1 11 7 10 12 1 11 1 12 1 11 2
81 13 1 15 1 10 0 9 0 2 2 11 11 2 2 13 1 12 2 13 1 11 10 0 9 1 9 0 13 1 10 9 0 9 10 0 9 1 9 2 10 9 13 1 0 9 2 13 15 13 1 10 9 1 9 1 9 2 15 16 15 4 13 1 13 15 3 1 9 1 10 0 9 1 0 9 1 9 0 1 11 2
31 11 11 2 10 9 0 15 13 2 3 1 15 2 1 9 1 11 11 2 15 4 13 1 13 1 10 8 9 11 11 2
32 1 9 1 10 9 1 11 1 12 2 13 9 16 13 3 1 15 2 1 10 9 16 4 13 10 9 1 10 9 1 11 2
9 11 11 15 13 13 1 10 9 2
23 10 9 13 1 10 9 1 9 15 10 9 0 13 1 3 2 13 1 9 1 9 13 2
16 10 9 2 13 10 9 2 1 11 7 1 9 4 13 0 2
10 15 13 16 13 3 9 1 10 9 2
77 3 13 1 13 3 16 10 11 1 11 2 9 0 0 2 4 13 0 9 1 9 1 10 9 1 9 2 7 16 10 16 13 3 3 13 9 1 10 9 0 2 11 11 8 11 7 11 11 11 2 4 13 1 15 10 9 1 0 9 2 16 2 15 13 2 1 9 0 2 1 10 9 11 7 11 2 2
38 13 10 0 9 1 9 13 10 9 1 9 3 15 13 10 9 1 9 1 10 0 9 10 9 4 13 1 0 9 1 13 9 7 3 13 10 9 2
20 13 9 0 2 1 9 7 4 13 3 3 1 10 9 9 1 10 1 11 2
10 3 3 15 13 10 9 1 10 9 2
33 11 15 13 10 12 1 11 7 13 10 12 1 11 1 12 10 9 1 11 16 13 2 1 9 2 13 10 9 0 13 1 11 8
40 8 3 2 10 9 7 9 13 3 16 11 13 1 10 9 1 10 9 1 10 9 1 11 2 10 15 15 4 13 1 11 1 12 2 2 13 15 1 11 2
17 13 1 11 2 11 2 7 3 13 1 11 2 11 1 10 11 2
17 10 9 0 13 12 9 0 2 15 1 9 7 15 1 9 0 2
17 10 9 13 10 9 0 7 0 2 9 1 10 15 11 3 13 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
14 11 11 11 13 15 1 10 9 16 13 1 10 11 2
44 13 3 1 11 2 3 15 13 1 10 9 15 10 9 11 1 11 13 1 13 1 11 2 7 1 10 13 15 1 10 9 1 11 11 2 13 1 11 2 7 3 1 11 2
24 10 9 13 1 11 2 12 9 7 12 9 13 10 9 16 15 13 1 9 0 7 9 0 2
52 10 11 11 11 11 2 13 10 9 13 1 9 1 9 7 9 1 0 9 0 9 1 10 9 1 11 2 1 10 9 1 9 11 2 10 11 11 11 2 9 1 9 9 11 7 1 10 0 9 11 11 2
21 3 1 12 11 13 10 9 7 4 13 1 11 11 2 3 1 9 1 11 2 2
13 13 3 10 9 1 9 1 11 11 2 12 2 2
13 11 11 11 2 13 1 12 2 13 10 9 0 2
57 10 0 9 4 13 1 12 9 0 1 10 9 11 11 1 9 1 9 0 2 10 9 0 4 13 1 12 9 2 12 9 7 12 9 13 10 9 8 1 9 1 12 9 0 0 9 9 0 9 0 13 1 9 0 7 0 2
8 4 15 13 1 10 0 9 2
31 10 9 16 13 10 9 9 1 16 13 3 0 1 13 15 0 1 10 9 1 9 2 13 15 1 13 15 1 10 9 2
21 11 13 10 9 1 10 9 1 11 2 11 2 1 10 9 1 3 1 12 9 2
28 10 9 13 10 9 0 1 10 11 2 11 11 11 11 2 7 10 9 1 9 0 11 1 10 0 9 0 2
78 10 9 15 10 9 13 13 10 9 1 9 2 1 15 1 15 10 9 0 13 1 10 9 2 13 1 10 9 2 9 3 7 13 15 1 10 9 7 9 12 9 10 15 1 15 2 16 13 1 10 12 9 13 10 9 1 12 2 3 7 10 9 13 10 9 1 10 9 1 12 9 1 10 9 0 7 11 2
17 10 9 4 13 13 10 12 9 1 9 0 7 12 9 1 9 2
25 10 9 0 7 9 0 15 13 1 10 9 1 9 0 13 1 9 0 2 9 7 9 2 9 2
17 15 13 10 9 1 9 3 0 1 9 1 13 3 1 10 9 2
6 2 15 13 1 11 2
21 3 1 10 12 15 13 7 13 10 9 2 11 1 9 1 11 2 11 11 2 2
20 10 9 13 1 11 7 13 13 7 10 9 4 13 1 3 1 11 1 9 2
15 1 10 9 0 1 10 9 15 13 10 11 1 10 11 2
63 10 9 1 9 13 1 10 9 12 2 16 13 1 10 9 11 11 1 10 0 9 1 10 9 0 2 9 1 10 15 13 10 9 1 10 9 7 13 1 11 11 2 7 10 15 1 10 15 13 3 1 10 0 9 1 10 9 0 1 10 0 9 2
16 10 9 1 10 9 13 2 7 13 1 10 9 2 1 9 2
34 16 11 11 13 10 0 9 4 13 2 13 2 10 9 16 10 9 13 16 13 1 10 9 2 1 3 0 7 3 0 16 15 13 2
31 1 0 13 12 9 3 1 10 9 2 3 10 9 1 9 13 0 9 1 9 1 13 10 9 0 0 1 10 9 0 2
10 3 13 9 1 9 1 10 9 0 2
20 1 9 7 1 10 9 10 9 15 13 1 10 9 1 9 1 10 9 0 2
64 13 0 9 1 11 7 10 9 3 15 13 13 2 1 10 9 11 15 13 1 10 9 3 11 15 13 0 1 15 15 4 13 1 0 7 15 13 10 9 13 1 16 15 15 13 10 9 1 15 2 1 10 9 13 1 10 9 1 11 1 13 1 11 2
28 13 13 15 1 10 0 9 1 10 9 1 11 2 3 1 10 0 9 1 11 11 2 11 11 7 11 11 2
24 10 9 13 10 0 9 1 10 11 2 12 9 12 7 0 1 10 9 2 11 1 11 2 2
12 1 9 12 13 1 10 9 1 12 12 9 2
36 10 9 1 10 9 13 1 10 9 2 16 13 9 0 2 9 0 7 1 9 2 13 1 9 13 1 10 9 2 7 10 9 1 9 0 2
35 1 12 2 10 9 4 13 1 9 1 11 2 11 1 9 0 2 2 7 4 13 2 13 1 10 9 0 1 11 1 10 9 1 11 2
32 1 10 9 15 13 10 9 1 10 9 1 9 7 1 10 9 2 1 9 2 1 3 3 13 9 1 13 10 9 1 9 2
14 10 9 0 13 10 9 1 10 9 0 1 11 11 2
28 10 9 1 11 11 1 10 9 1 9 2 0 7 9 2 13 3 3 1 10 9 1 10 9 0 2 11 2
39 13 3 12 9 16 11 13 13 10 9 0 16 13 1 10 9 1 10 9 7 2 9 1 15 2 10 9 1 9 2 13 1 10 9 0 1 15 0 2
22 9 13 1 9 0 16 10 9 1 10 9 13 1 10 9 1 10 9 0 11 11 2
26 15 13 10 9 10 11 11 11 8 8 2 16 13 15 1 10 9 1 9 1 10 9 1 10 11 2
14 3 10 9 13 0 2 10 9 3 0 13 1 9 2
46 1 0 2 11 15 13 16 13 10 10 9 1 2 10 9 7 9 1 10 9 0 15 4 4 13 1 10 0 9 1 10 9 2 1 10 9 1 9 7 9 1 10 9 1 9 2
19 10 12 1 11 1 12 15 13 10 0 9 2 13 10 9 1 9 1 8
9 10 9 12 13 10 9 12 9 2
30 13 2 5 2 8 2 7 2 8 2 5 2 12 9 1 11 2 7 13 10 9 1 9 1 2 5 2 8 2 2
14 13 0 1 11 2 3 15 13 1 10 9 1 11 2
12 11 11 13 10 9 1 9 1 10 9 11 2
25 7 1 12 9 1 9 1 11 7 10 9 0 2 3 7 1 10 9 1 11 11 2 11 2 2
10 15 13 1 13 1 10 9 3 13 2
19 10 11 11 13 10 9 1 10 9 11 13 1 10 9 0 11 1 12 2
30 10 9 1 10 0 11 3 4 13 3 0 7 0 2 7 15 4 13 10 9 7 0 9 2 16 13 1 10 9 2
68 3 2 16 1 9 13 13 10 9 1 10 9 0 1 13 10 9 1 9 2 10 9 0 13 3 0 2 9 2 9 2 9 2 9 0 2 13 1 7 1 9 2 8 2 1 10 0 7 10 9 0 2 9 1 10 9 2 9 0 2 9 1 10 9 2 8 2 2
11 1 9 15 13 12 9 16 13 10 9 2
24 10 0 9 1 11 11 13 10 0 9 1 10 9 0 7 4 13 9 1 0 9 1 11 2
30 13 10 0 9 0 1 10 9 0 1 11 2 11 2 11 2 11 2 10 11 2 11 11 2 11 7 9 1 11 2
18 10 9 1 9 13 10 9 1 2 10 9 1 10 9 1 9 2 2
11 13 1 9 1 10 9 1 11 2 8 2
38 9 1 9 2 11 11 11 2 9 1 11 2 10 9 16 13 10 9 1 10 9 1 11 2 13 0 1 12 9 1 9 7 10 9 1 12 9 2
53 11 4 4 13 1 10 9 0 1 11 11 1 10 9 11 11 2 1 9 13 10 9 1 13 15 1 12 2 10 9 13 9 7 9 0 1 11 11 2 11 11 2 10 15 15 13 1 9 0 1 11 11 2
35 13 10 9 2 11 11 11 2 16 13 10 9 0 2 7 1 10 9 3 11 13 1 10 0 9 1 10 9 1 10 9 1 10 11 2
30 10 9 15 13 0 1 10 0 9 1 10 9 1 11 2 1 9 12 2 0 1 10 9 0 1 10 11 1 11 2
31 1 10 9 13 10 9 11 11 1 10 11 11 2 11 11 7 10 9 7 10 11 1 10 11 7 10 9 11 7 11 2
24 9 13 9 3 13 1 10 9 1 9 2 1 15 10 3 9 13 2 10 8 2 1 9 2
42 10 0 9 2 15 13 1 10 9 1 15 1 10 3 0 9 1 10 9 0 2 10 11 2 1 10 0 9 16 15 13 10 9 11 1 9 7 10 11 1 11 2
19 13 13 15 16 10 9 16 13 9 1 10 9 13 1 9 1 13 15 2
12 15 13 1 10 0 9 13 1 10 0 9 2
23 1 9 0 2 15 13 10 9 2 10 9 0 16 13 10 9 1 10 9 1 10 9 2
26 12 9 0 4 13 1 11 11 2 11 11 2 7 10 9 11 11 11 2 11 11 2 1 10 9 2
16 4 13 7 13 1 11 11 2 1 15 13 10 0 0 9 2
25 10 9 4 13 3 1 9 1 9 1 10 9 1 10 9 7 1 10 9 1 10 11 1 11 2
20 10 9 2 11 11 4 13 1 10 11 11 1 10 9 9 1 12 9 8 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
25 1 10 9 2 10 9 13 16 10 9 0 13 2 9 1 10 9 0 16 15 4 7 13 2 2
17 13 9 1 10 9 13 10 0 9 16 13 9 0 1 10 9 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
51 3 1 13 15 1 10 9 0 1 9 7 9 16 4 13 13 10 9 1 10 0 9 2 13 1 10 2 11 2 2 13 1 9 1 9 2 9 7 9 1 15 16 3 15 13 1 13 15 1 9 2
17 1 10 9 1 10 9 2 10 9 15 13 2 13 3 12 9 2
35 3 13 10 9 1 10 9 3 1 10 9 2 10 9 1 10 0 9 1 10 9 1 10 3 2 7 10 1 9 1 10 9 1 11 2
14 2 11 11 11 2 3 15 13 11 11 11 3 0 2
9 10 9 4 13 1 10 9 12 2
29 7 2 16 13 13 10 9 2 4 13 10 0 9 1 10 9 16 3 13 10 9 1 10 9 13 1 10 9 2
44 10 9 0 13 1 10 9 2 16 15 13 1 9 0 1 10 9 16 13 2 10 11 2 2 13 13 2 16 13 10 9 7 10 11 1 10 9 1 11 1 10 0 9 2
18 1 10 9 12 15 13 10 9 1 10 10 9 2 4 13 10 9 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
12 2 10 9 15 4 13 1 10 9 0 0 2
28 3 13 1 10 9 1 9 1 9 7 13 10 0 9 7 10 9 1 10 9 13 3 0 7 10 15 0 2
12 3 15 2 10 9 11 7 11 13 13 15 2
40 10 9 0 1 10 9 13 16 10 9 0 1 10 9 0 1 10 10 9 1 10 9 3 13 10 12 5 12 5 8 15 15 4 13 2 10 0 9 2 2
28 10 0 9 1 10 9 11 2 12 13 10 9 1 9 2 13 15 0 1 10 9 1 9 1 12 7 12 2
21 10 9 7 11 11 2 13 10 9 1 9 1 9 0 1 10 9 1 10 9 2
30 3 15 4 13 10 9 1 10 9 1 10 9 0 1 10 9 1 9 1 9 7 1 9 2 3 16 4 4 13 2
11 3 13 9 7 3 13 10 9 16 13 2
18 10 9 7 9 2 11 11 2 13 10 9 1 10 9 1 10 9 2
27 1 10 9 15 4 13 1 11 13 10 9 7 13 1 10 9 1 10 9 2 0 1 10 9 1 9 2
24 11 13 10 9 10 9 1 13 1 11 7 1 13 1 10 0 9 1 10 9 1 11 11 2
48 10 9 13 10 9 1 10 9 16 13 1 8 2 8 1 10 9 1 10 9 2 16 9 3 15 13 7 15 13 16 10 9 13 10 11 11 2 7 11 4 13 10 9 1 8 2 8 2
59 1 10 9 0 7 9 15 13 1 10 9 7 15 13 1 10 9 1 10 9 1 10 9 2 7 10 9 1 10 9 1 10 9 0 1 10 9 1 10 9 15 13 0 1 10 13 10 9 1 10 9 1 10 9 1 10 11 0 2
23 11 3 13 16 10 9 1 9 16 13 15 13 1 10 9 1 9 1 9 7 1 9 2
52 11 2 8 2 9 1 9 2 2 13 10 9 13 1 10 0 9 1 9 0 0 0 2 16 13 1 9 1 10 9 0 2 13 15 3 1 12 9 1 9 2 1 10 11 2 1 15 15 13 3 11 2
13 13 0 1 15 1 11 2 3 15 13 1 12 2
36 3 2 11 4 13 15 1 10 9 1 9 1 11 2 1 10 16 15 13 10 9 1 11 7 15 1 11 2 1 10 9 1 11 7 11 2
32 15 13 10 9 1 9 7 10 9 2 7 10 9 13 16 4 13 3 0 2 1 15 13 1 10 9 16 15 4 13 3 2
34 11 13 10 9 1 9 0 0 0 16 13 1 9 1 10 9 11 2 13 3 12 9 1 9 1 10 11 2 1 15 15 3 11 2
7 4 4 13 1 0 9 2
37 16 10 9 13 1 13 3 2 10 9 13 3 4 13 1 10 9 10 9 4 13 1 16 3 4 1 13 15 7 15 13 10 9 1 10 9 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
35 10 9 13 3 1 10 9 16 13 10 12 9 1 9 7 2 1 10 9 2 10 9 4 4 13 1 10 9 1 11 1 10 9 0 2
11 1 10 9 1 10 9 15 15 13 3 2
30 7 10 9 1 11 3 13 1 9 2 7 13 10 9 1 13 1 10 9 7 13 15 1 15 10 16 15 4 13 2
49 15 13 3 1 10 2 9 2 10 9 0 11 11 2 10 9 11 11 2 10 9 11 2 11 2 3 7 10 9 11 11 2 10 9 0 1 11 11 7 10 9 0 11 11 11 2 1 15 2
48 1 9 1 13 10 9 1 10 9 2 10 9 1 10 9 2 9 2 1 13 10 9 1 10 11 4 4 13 1 10 9 2 11 11 2 2 16 1 9 0 4 13 13 1 2 9 2 2
21 10 0 9 1 9 13 0 2 3 3 13 1 9 1 9 13 1 9 1 9 2
27 9 1 10 11 1 10 11 2 13 1 10 9 1 11 1 10 11 1 11 11 1 11 2 9 1 11 2
47 7 15 2 10 10 11 11 2 16 4 13 1 10 9 1 1 10 0 0 9 1 10 11 1 10 11 1 12 2 4 13 10 9 1 11 11 1 9 1 10 0 0 9 1 10 9 2
13 10 9 13 1 9 1 9 0 1 9 7 9 2
16 11 4 13 10 9 3 0 7 3 13 1 10 9 1 11 2
50 10 9 0 1 11 11 13 10 9 1 10 9 1 9 0 2 13 10 9 1 10 9 1 10 0 11 2 1 10 9 1 10 11 11 1 11 2 1 10 9 16 13 1 9 1 10 9 0 0 2
59 10 9 1 10 11 11 1 11 1 11 1 10 9 1 11 2 11 11 2 13 16 10 9 1 11 13 9 1 13 9 1 10 11 1 10 11 1 3 1 12 9 1 9 10 0 12 1 11 2 16 3 13 10 9 1 13 10 9 2
12 11 13 1 10 9 13 9 0 1 10 9 2
20 10 0 9 4 13 3 1 10 0 9 0 1 10 9 0 1 10 9 0 2
41 1 11 1 12 2 1 9 1 10 9 1 9 1 10 9 2 10 9 1 10 9 0 11 2 13 10 9 1 13 10 9 13 1 9 1 9 0 1 10 9 2
6 15 13 1 9 0 2
16 10 9 1 10 9 0 4 13 10 9 1 10 9 1 11 2
54 10 9 0 1 10 0 9 13 13 10 9 2 1 13 1 10 9 1 9 2 2 7 1 3 7 1 10 9 1 10 9 15 13 10 9 1 12 9 2 7 3 15 13 1 10 9 0 2 12 7 12 9 2 2
27 3 13 9 1 13 3 10 9 1 10 9 7 1 13 10 15 3 3 1 10 12 2 9 1 9 2 2
51 3 2 10 9 1 11 13 0 1 10 9 1 10 9 0 8 12 1 10 11 2 3 7 11 3 13 1 9 1 13 1 11 1 9 1 16 10 9 2 0 2 3 13 10 0 9 2 15 15 0 2
17 10 9 1 10 9 1 9 0 7 1 9 4 13 1 10 9 2
19 11 11 11 2 11 2 12 1 11 12 2 13 10 9 7 9 1 11 2
14 1 9 1 10 9 8 11 13 11 2 11 7 11 2
11 13 9 1 11 1 11 2 9 1 11 2
11 13 0 16 3 15 13 10 9 0 0 2
7 9 1 11 2 12 2 2
31 1 10 9 11 11 2 4 13 1 10 9 0 1 10 10 9 0 2 13 15 3 1 10 9 1 10 9 1 10 9 2
45 10 9 0 2 15 13 10 11 1 11 2 13 10 11 10 9 1 10 13 10 9 0 1 10 11 1 10 11 2 1 15 15 15 13 1 10 9 1 9 3 4 13 1 11 2
24 11 13 10 9 0 16 13 1 10 9 1 11 7 11 1 13 1 10 9 8 1 10 11 2
21 10 9 13 10 9 3 13 2 7 3 13 10 12 9 1 10 9 1 10 9 2
20 3 15 13 10 9 1 9 2 9 7 9 1 7 10 9 13 10 0 9 2
21 3 1 10 9 1 10 11 2 13 1 10 9 1 4 1 13 1 10 9 0 2
27 10 11 11 11 0 15 13 1 10 9 0 2 0 3 1 10 9 7 10 9 0 1 10 9 1 11 2
17 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
25 10 9 13 9 1 9 2 13 10 9 1 13 9 1 9 13 15 3 1 10 9 0 1 9 2
24 3 13 10 9 0 1 10 9 0 1 10 9 1 9 0 1 10 9 16 13 1 10 9 2
18 10 9 13 10 9 0 1 9 12 9 1 10 9 12 1 10 9 2
23 3 1 10 9 15 13 10 9 3 0 1 10 9 2 1 10 9 1 9 0 7 0 2
18 10 11 12 11 13 10 9 0 0 1 9 0 13 1 10 11 11 2
16 10 9 13 10 9 1 10 9 1 11 7 11 0 11 11 2
12 11 11 11 13 3 10 9 1 9 7 9 2
25 10 11 2 11 11 13 10 9 0 1 9 1 11 1 10 9 1 11 2 9 1 10 11 2 2
30 3 3 1 12 2 11 11 4 13 1 10 9 1 10 9 10 9 13 13 3 10 9 0 15 13 1 10 9 0 2
18 10 9 13 10 9 0 1 5 12 9 1 10 5 12 1 10 9 2
13 3 4 13 10 11 12 2 10 9 1 12 9 2
29 1 10 9 2 10 9 1 11 13 1 10 9 1 13 10 9 0 1 10 9 1 15 1 10 9 1 10 9 2
8 10 9 2 13 3 0 2 2
10 10 9 15 4 13 3 1 10 9 2
15 11 11 2 13 10 9 1 9 0 0 1 10 9 11 2
21 11 13 15 1 10 9 3 0 1 10 9 2 7 13 0 1 0 9 13 0 2
20 11 11 11 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 0 2
26 15 4 13 3 4 13 10 9 1 9 1 9 2 7 15 0 15 15 4 13 1 10 9 3 0 2
12 10 9 1 9 1 10 9 13 1 5 12 2
35 9 2 9 7 9 13 10 9 0 1 10 9 3 0 2 10 9 13 13 1 3 10 9 1 10 9 2 16 10 9 15 13 10 9 2
22 10 9 13 10 9 3 0 2 11 15 13 1 9 0 1 10 9 7 1 10 9 2
41 10 0 9 2 13 10 9 1 12 5 1 10 9 0 2 15 15 9 15 7 13 10 9 2 2 7 1 11 15 15 13 1 10 12 5 2 13 3 15 9 2
23 7 3 13 1 13 1 10 9 1 10 9 2 16 13 10 9 3 0 1 13 10 9 2
21 15 13 1 10 9 1 11 2 11 2 3 1 10 9 0 2 2 11 7 11 2
30 1 10 11 1 11 13 1 10 9 1 10 9 1 11 11 1 11 2 1 10 9 1 11 7 1 10 9 1 11 2
47 11 11 2 3 3 13 1 2 11 11 2 2 13 1 10 9 1 11 2 10 11 2 10 12 1 11 1 12 2 13 1 10 9 0 0 16 13 1 10 11 1 9 1 10 9 12 2
14 10 9 4 13 1 11 1 10 9 0 1 11 11 2
8 15 15 13 3 3 13 3 2
27 10 9 0 1 10 11 11 13 1 12 12 1 9 1 10 9 16 13 1 11 1 12 1 11 1 12 2
28 10 0 9 0 15 11 13 13 1 10 11 1 10 11 1 10 12 1 10 9 1 10 9 1 9 1 11 2
24 1 10 9 2 15 13 1 10 9 11 11 1 10 0 9 1 10 9 1 9 1 9 0 2
12 1 10 9 1 12 10 9 13 1 12 9 2
8 13 10 9 1 9 1 12 2
32 1 15 10 9 3 9 4 13 1 10 9 0 16 13 9 2 9 0 7 0 7 10 9 1 9 1 10 9 1 10 9 2
54 3 15 13 9 7 9 2 15 13 10 9 2 10 9 13 0 2 10 9 13 0 2 13 10 9 1 9 16 3 15 4 13 2 4 7 13 15 2 13 10 0 9 1 10 9 16 10 9 15 13 1 10 9 2
50 10 9 0 1 9 2 11 11 2 13 16 10 9 0 4 13 10 9 1 16 10 9 15 13 1 10 9 1 10 9 1 9 1 9 1 11 2 10 9 16 4 13 10 2 9 2 1 10 9 2
25 1 12 2 10 9 1 10 0 9 11 11 11 1 10 9 13 9 1 10 9 0 7 10 9 2
47 16 15 4 13 16 15 10 11 2 1 10 9 13 1 10 9 0 2 7 10 11 13 1 2 9 0 2 16 10 9 15 13 1 9 2 7 1 0 9 2 9 7 9 2 3 2 2
45 10 0 9 13 1 10 9 0 1 10 11 1 11 1 11 7 13 10 9 1 9 1 9 7 0 0 9 0 1 10 9 2 10 9 4 13 1 12 9 0 7 12 9 2 2
65 1 9 2 13 10 9 3 0 1 10 9 13 1 10 9 16 13 9 2 10 11 1 11 1 10 11 1 11 11 1 10 11 11 2 13 1 12 9 2 15 13 1 10 9 2 13 15 1 15 9 1 10 0 11 11 1 11 11 7 11 1 11 2 11 2
45 10 11 11 15 13 1 10 9 1 10 9 1 11 2 15 1 10 9 0 16 13 10 9 11 2 7 1 10 9 1 10 9 1 10 11 2 1 10 7 15 13 10 12 9 2
13 10 0 9 1 9 1 10 9 7 3 3 0 2
23 1 10 9 15 13 1 10 0 12 9 0 1 9 0 15 4 4 13 1 10 9 0 2
15 3 13 0 13 10 9 0 1 13 10 9 1 9 0 2
30 4 13 12 9 1 10 9 1 9 0 7 12 1 9 1 9 1 12 1 9 7 12 1 9 7 9 1 10 9 2
46 10 11 1 11 4 13 13 10 9 1 10 9 0 7 13 2 1 13 1 3 2 1 10 9 7 10 9 0 1 10 0 9 0 2 1 10 16 13 13 10 9 0 1 10 9 2
47 11 10 11 4 13 13 10 9 1 10 9 7 1 10 0 9 7 3 4 13 13 1 10 9 1 11 2 3 15 4 13 10 0 9 1 11 11 2 16 15 13 1 10 9 1 9 2
32 10 9 13 10 9 0 10 12 1 11 1 12 2 1 10 9 1 10 9 1 9 0 2 9 0 2 9 0 7 9 0 2
26 11 15 13 16 13 10 11 11 2 3 2 3 2 1 10 2 9 2 1 10 9 1 10 11 11 2
41 11 2 11 2 1 11 11 11 2 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 1 11 2 1 10 9 1 9 7 9 1 11 2 10 2 11 2
17 10 9 0 13 10 9 16 13 10 10 9 0 1 10 9 13 2
33 10 9 13 9 1 9 1 9 7 13 10 9 1 9 13 1 10 9 1 10 9 3 1 13 10 9 1 9 0 1 10 9 2
35 1 4 13 15 3 2 11 13 10 9 1 10 9 7 2 1 10 9 1 9 2 4 1 13 10 9 2 16 13 10 9 11 11 11 2
62 1 10 12 9 2 10 9 1 11 13 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
81 2 13 15 0 2 10 9 1 9 13 1 13 1 3 1 12 8 1 12 8 2 10 9 1 10 11 11 4 13 1 10 11 11 2 9 1 10 9 11 2 15 4 9 1 10 9 12 9 2 12 1 9 7 12 1 9 2 10 9 1 10 11 13 3 0 1 10 9 1 10 9 7 1 10 9 0 2 2 13 11 2
24 1 10 9 1 9 9 0 2 4 13 15 1 9 10 9 1 9 7 10 9 1 10 9 2
14 10 11 11 11 13 10 9 3 1 10 9 1 11 2
17 10 9 9 1 9 1 10 9 0 7 9 0 1 12 9 0 2
46 1 10 12 9 2 12 13 1 10 11 2 12 1 10 9 1 10 11 11 11 2 12 1 10 9 1 11 11 1 11 2 12 1 10 11 1 11 7 3 15 1 10 9 1 11 2
38 0 11 1 11 2 1 9 2 0 11 1 11 2 7 3 11 2 13 10 9 0 1 10 9 1 11 2 1 10 9 1 11 2 11 2 11 2 2
24 10 9 15 10 9 1 11 13 10 9 2 15 13 13 1 10 9 7 4 13 1 10 9 2
24 11 13 10 15 9 2 13 0 7 0 2 7 3 4 13 1 10 9 7 9 15 13 11 2
33 10 9 15 13 3 1 10 9 1 10 11 1 10 9 2 2 9 7 9 1 10 9 2 2 9 0 7 0 1 10 9 0 2
46 1 12 2 16 3 13 0 1 10 9 0 2 15 13 10 9 0 14 1 13 3 15 4 13 10 9 0 2 10 9 4 13 1 9 1 10 10 9 13 1 11 2 11 7 11 2
