489 11
8 11 11 1 9 12 1 9 12
14 10 12 4 1 3 13 10 9 7 4 13 10 9 2
14 10 10 9 0 13 1 4 13 3 1 15 15 13 2
26 1 10 0 9 3 2 3 2 13 9 1 13 16 15 0 13 3 3 0 2 13 9 7 9 0 2
9 15 13 9 1 9 1 10 9 2
8 13 0 2 15 4 4 13 2
7 10 9 13 1 10 11 2
5 9 1 10 9 2
10 2 15 13 10 0 9 1 9 2 2
37 1 13 11 2 15 15 4 3 13 0 2 4 13 3 10 9 1 10 9 2 1 11 11 2 13 1 10 9 1 10 2 11 1 10 9 2 2
24 10 9 0 2 16 15 13 2 13 1 11 7 1 11 2 1 13 10 9 1 13 10 9 2
43 10 9 0 1 10 0 11 13 9 1 10 0 9 2 13 1 10 9 1 10 9 7 3 1 10 9 0 16 10 9 1 10 10 0 9 0 4 13 1 10 9 0 2
60 11 2 1 10 11 2 12 9 3 2 3 15 13 11 2 2 4 13 12 9 0 1 11 3 4 4 13 1 9 7 9 1 9 1 10 11 15 4 13 1 9 0 10 9 0 16 4 13 2 10 12 9 12 2 10 9 1 10 11 2
73 11 11 11 2 11 2 2 4 4 13 0 7 0 12 9 2 12 9 2 12 9 7 12 9 2 15 13 1 10 11 11 1 10 11 11 2 15 4 4 13 1 10 9 0 2 16 15 13 1 10 9 1 10 0 9 0 1 11 2 1 12 9 1 11 11 11 2 1 10 11 9 0 2
35 1 11 2 1 10 9 11 13 0 3 11 2 12 9 2 10 0 9 1 11 15 13 1 11 7 3 4 3 13 10 9 1 10 11 2
58 10 9 1 10 9 1 11 11 4 13 1 10 9 1 10 10 9 9 1 0 9 2 1 10 9 1 10 9 7 10 9 7 1 10 9 1 9 1 10 9 0 1 9 1 10 9 7 1 10 2 9 2 15 4 3 13 15 2
21 3 4 3 4 13 15 13 10 10 9 2 7 10 9 15 15 4 13 13 15 2
34 2 1 9 10 2 4 3 13 2 13 1 13 1 9 10 9 1 10 9 0 2 1 13 13 16 13 10 11 15 3 13 9 2 2
27 10 9 15 10 9 0 13 1 11 11 2 10 9 1 10 11 3 1 9 13 10 9 0 2 13 0 2
23 1 10 0 9 10 9 1 10 9 4 4 13 1 0 9 1 10 9 1 10 9 11 2
8 11 2 10 9 1 10 9 2
63 13 1 9 1 10 9 2 13 0 1 10 9 1 10 11 7 1 10 11 2 3 15 13 16 13 10 9 1 10 9 2 13 10 9 7 2 13 1 10 9 2 10 9 0 13 10 9 1 9 7 9 0 1 13 13 16 10 9 4 1 9 13 2
20 1 10 9 0 10 9 13 1 9 7 10 9 0 15 13 1 10 9 0 2
19 3 9 0 1 11 2 13 10 9 1 10 9 0 13 1 10 9 0 2
20 13 10 9 1 10 12 2 7 15 13 1 9 0 1 13 9 1 11 11 2
19 10 9 1 11 2 3 2 4 13 3 1 0 1 10 9 0 1 11 2
16 2 11 16 13 15 13 1 9 2 4 13 15 1 13 15 2
17 3 1 11 13 16 15 4 13 1 3 1 10 9 3 2 2 2
51 10 2 9 2 1 11 15 15 13 1 11 11 2 15 10 9 3 2 9 1 10 9 1 10 11 12 2 4 13 10 9 1 11 13 15 1 10 9 1 10 9 1 9 2 3 3 0 1 10 9 2
22 2 16 15 13 15 15 13 7 15 13 2 15 13 1 13 15 3 2 2 13 11 2
6 13 1 9 10 3 2
7 3 10 9 1 11 11 2
12 2 10 11 4 13 3 1 13 1 9 10 2
12 13 1 15 10 9 0 2 10 11 11 11 2
9 13 10 9 1 10 2 9 2 2
9 7 10 2 9 2 1 11 11 2
41 16 3 13 9 13 1 10 9 16 10 9 4 13 12 9 3 9 0 2 16 13 0 13 16 10 9 9 1 9 4 13 2 3 2 1 10 0 9 0 2 2
12 2 7 6 2 3 13 3 2 13 11 2 2
10 7 3 6 2 3 6 2 0 11 2
14 2 15 3 4 3 13 1 9 1 13 10 9 0 2
20 10 12 12 13 1 9 1 10 9 0 1 10 9 1 11 3 1 9 0 2
5 4 13 10 9 2
27 10 0 9 11 4 1 3 13 10 10 9 7 15 13 3 1 13 10 9 15 13 10 9 1 10 9 2
32 3 1 10 9 11 4 4 13 1 11 2 3 3 3 1 13 15 1 10 9 1 9 1 10 9 4 4 13 1 10 9 2
22 10 9 1 11 1 10 12 9 1 10 9 1 11 7 11 15 13 3 10 9 0 2
6 10 9 13 15 9 2
11 10 9 9 2 3 2 3 4 13 2 2
11 15 13 1 10 0 9 12 9 1 11 2
31 10 9 13 10 0 9 1 9 7 10 9 15 13 10 9 2 11 11 2 12 9 2 1 11 11 11 3 15 4 13 2
5 9 13 1 11 2
17 1 9 1 11 7 11 4 4 13 12 9 1 9 7 9 0 2
32 4 3 13 10 9 1 13 10 9 7 15 4 13 1 15 3 1 4 13 10 9 1 9 0 2 16 13 9 0 1 9 2
40 3 2 10 9 4 13 1 9 1 9 10 9 0 2 11 11 11 2 12 9 2 7 11 11 2 12 2 1 10 9 3 1 13 9 7 9 1 13 9 2
16 4 13 1 12 1 10 9 0 2 3 10 11 2 13 2 2
15 15 4 13 10 9 1 10 9 2 3 15 4 3 13 2
5 10 0 9 0 2
15 2 3 10 9 13 10 9 13 10 9 1 10 9 2 2
11 2 15 13 16 13 9 0 7 0 2 2
16 2 15 13 16 4 3 13 1 9 11 11 7 1 9 11 2
22 3 2 16 10 9 3 13 10 9 1 9 2 13 13 0 16 15 13 10 9 0 2
14 10 9 1 10 10 9 13 3 3 0 7 0 2 2
12 2 10 9 0 13 1 11 13 3 3 0 2
28 10 9 15 13 1 10 11 2 13 1 10 9 2 4 13 1 11 15 15 13 1 10 2 11 2 2 3 2
8 9 10 3 0 7 9 0 2
33 10 0 2 9 0 2 3 3 16 0 2 13 1 4 13 2 9 2 10 9 1 9 15 13 11 2 11 2 11 2 11 11 2
9 1 10 12 13 10 11 1 11 2
14 9 1 9 13 3 15 1 10 0 9 1 11 11 2
33 11 1 10 9 7 11 1 10 9 13 10 0 9 2 9 0 1 10 9 1 10 9 2 1 10 0 9 1 11 7 10 11 2
8 0 9 2 3 1 9 0 2
11 11 2 10 9 13 1 10 9 1 9 2
7 15 4 13 10 9 11 2
8 4 13 1 13 10 9 0 2
16 3 4 13 1 9 1 15 7 10 9 1 10 10 9 2 2
15 13 1 9 2 4 13 3 3 0 9 3 1 10 9 2
17 7 10 9 1 10 9 0 3 15 13 10 9 2 10 10 9 2
5 10 0 9 0 2
14 10 11 3 13 10 9 16 10 2 9 2 15 13 2
35 1 10 9 2 1 12 9 3 2 13 9 12 2 13 3 10 9 16 10 9 13 1 3 0 1 10 9 1 10 9 13 1 10 9 2
28 1 10 0 9 1 9 10 9 1 10 10 9 13 10 9 0 2 1 15 9 7 9 15 13 1 10 9 2
45 1 11 7 1 9 2 9 2 1 10 11 1 11 2 3 11 3 3 2 9 12 2 9 11 1 11 12 2 10 11 13 10 11 11 3 13 1 10 11 1 10 0 9 11 2
14 2 15 13 9 15 3 15 13 2 13 3 11 2 2
16 15 15 13 2 1 11 2 1 13 2 0 2 13 9 2 2
5 3 3 2 3 2
21 12 9 1 11 7 11 2 10 10 9 2 10 10 9 2 13 3 10 0 9 2
14 4 13 10 10 9 1 10 9 1 10 0 9 0 2
16 10 9 0 13 0 7 13 1 13 1 10 9 2 13 15 2
20 10 3 1 13 9 1 10 9 15 10 9 0 13 10 9 1 13 10 11 2
31 10 9 15 13 3 10 15 9 2 7 10 0 9 1 10 11 15 4 13 10 9 7 10 9 1 10 9 13 0 2 2
22 2 10 9 13 3 0 1 10 9 1 13 10 9 7 1 3 13 15 1 9 2 2
5 3 13 9 9 2
8 4 13 15 15 15 15 13 2
5 13 3 0 9 2
13 15 13 9 0 1 3 1 9 2 15 13 0 2
10 3 15 4 13 7 4 13 10 9 2
23 13 10 9 13 1 13 3 2 3 10 9 13 3 3 1 10 9 2 13 12 9 3 2
12 0 10 9 1 11 1 10 9 2 12 2 2
39 10 9 1 10 9 2 3 13 1 9 2 9 7 9 0 2 7 3 13 1 9 7 9 0 2 3 16 13 2 13 0 9 1 10 9 1 10 9 2
21 15 4 13 1 11 11 2 12 9 2 0 9 1 12 2 13 1 10 11 11 2
25 2 3 1 10 0 9 2 13 11 2 4 13 10 9 2 10 9 13 13 1 9 3 1 15 2
27 7 16 1 9 1 3 2 1 9 1 10 0 9 1 10 9 2 4 13 15 3 2 13 3 10 9 2
39 15 13 16 1 10 9 13 3 13 15 1 10 9 7 13 15 1 9 1 13 2 16 3 15 13 10 9 0 0 16 15 13 10 9 1 13 10 9 2
10 2 11 2 11 7 11 4 13 3 2
34 1 11 4 13 15 1 10 0 9 2 7 10 11 1 10 0 9 2 15 2 0 2 2 4 13 15 1 3 1 10 9 3 0 2
42 3 0 10 9 2 1 12 9 0 10 9 2 15 4 13 9 1 10 2 9 1 10 9 2 1 11 7 11 2 10 9 0 7 0 13 1 10 9 0 3 0 2
12 1 10 9 3 10 9 7 10 12 9 0 2
18 9 2 1 10 9 2 1 10 9 13 3 3 1 13 15 1 9 2
43 3 4 4 13 9 11 2 9 1 10 9 1 10 11 2 3 3 2 2 15 1 10 12 9 1 10 9 13 1 10 9 11 11 2 3 1 9 1 10 9 1 11 2
30 1 10 9 1 10 0 9 15 13 10 2 9 0 2 2 10 9 1 9 2 10 9 1 9 2 10 9 0 0 2
24 1 15 2 11 13 1 10 12 9 11 2 3 15 13 3 2 16 15 13 1 10 9 0 2
15 1 10 9 15 13 9 0 2 9 7 13 1 0 9 2
7 9 7 9 13 1 9 2
19 1 9 2 13 3 10 11 1 11 2 13 1 9 3 12 9 1 12 2
21 9 9 0 1 10 9 1 9 11 11 3 4 13 9 10 9 1 10 9 11 2
27 2 4 13 1 10 9 3 1 10 9 2 2 15 13 10 9 11 11 11 2 10 0 9 1 10 11 2
16 1 9 15 13 12 9 1 10 15 12 13 3 1 12 9 2
7 10 0 9 1 11 11 2
17 1 10 9 11 13 3 2 3 2 13 10 10 9 1 0 9 2
14 1 10 9 2 10 9 7 12 9 1 0 9 0 2
35 10 9 2 10 10 9 4 13 12 9 1 9 2 3 12 9 1 9 2 2 15 13 1 10 9 1 12 9 0 7 15 13 16 13 2
24 10 10 9 13 2 1 9 3 0 2 1 10 9 1 12 9 0 2 11 11 7 11 11 2
18 10 0 11 1 11 2 10 0 11 1 11 2 10 0 11 1 11 2
14 7 1 9 13 3 10 9 1 9 2 1 9 0 2
9 10 9 13 0 9 1 9 0 2
37 0 13 10 9 0 7 3 3 10 9 2 3 1 9 2 0 1 9 13 2 1 10 9 0 1 9 7 12 9 0 15 4 13 1 10 9 2
13 10 15 15 13 3 13 1 10 9 9 1 9 2
32 10 9 15 15 13 10 10 9 2 13 1 11 1 11 1 10 9 1 9 0 2 15 13 13 10 9 1 9 1 10 11 2
40 1 10 9 1 11 7 1 11 2 1 10 9 1 10 11 1 11 2 1 10 9 0 2 1 10 9 1 10 9 1 9 1 10 9 2 2 1 10 9 2
19 9 2 11 11 2 2 2 13 1 11 2 1 9 0 2 13 1 9 2
5 9 12 10 9 2
9 9 12 7 10 9 1 9 12 2
14 2 11 2 2 1 11 11 2 1 9 1 9 0 2
14 1 9 12 1 9 12 10 9 2 9 0 0 2 2
54 1 10 9 16 10 9 13 13 7 13 2 15 4 13 3 9 2 13 2 2 7 13 1 9 10 9 13 1 10 9 7 13 10 9 1 9 2 9 3 13 1 10 9 0 15 3 13 3 13 10 10 9 0 2
25 10 0 13 10 9 1 10 9 7 4 13 3 1 13 9 7 13 1 12 10 9 1 10 9 2
20 13 10 9 1 12 9 2 3 13 3 3 2 13 3 10 9 2 13 2 2
41 1 10 9 1 13 2 9 2 9 2 9 2 4 13 9 15 2 13 2 13 10 9 1 12 9 2 13 10 9 1 10 9 0 7 1 10 9 1 10 9 2
29 13 2 13 2 13 1 9 2 13 10 0 9 2 13 10 9 0 1 13 10 0 9 1 0 9 0 7 0 2
10 1 9 2 1 15 2 10 0 9 2
18 16 13 1 10 9 3 1 10 9 2 13 1 10 9 1 10 9 2
33 16 10 9 0 3 13 3 0 2 10 0 1 13 15 10 9 13 3 10 9 15 2 13 1 3 2 1 9 1 10 9 0 2
27 1 10 9 0 2 13 10 9 0 2 0 1 9 7 0 1 9 0 7 9 0 15 13 10 9 0 2
54 13 15 10 10 9 1 10 9 1 9 7 13 10 9 2 3 3 1 12 9 10 9 1 10 9 2 1 10 9 13 1 11 11 1 11 11 1 10 9 13 2 7 16 13 10 9 15 13 15 0 1 11 0 2
30 13 3 2 3 13 2 0 1 13 15 1 9 7 9 2 3 10 9 2 1 13 10 9 0 1 10 9 1 3 2
7 2 11 11 2 1 11 2
7 13 3 1 15 10 9 2
23 10 9 11 2 9 0 1 11 2 15 13 3 2 12 9 3 2 16 11 15 4 13 2
19 1 10 9 2 2 4 13 11 2 2 13 3 13 2 16 13 15 2 2
5 0 9 1 9 2
64 15 3 13 1 10 9 13 15 2 13 1 10 9 1 10 9 2 1 10 11 11 15 13 3 0 1 10 9 0 1 10 9 7 15 13 2 3 2 1 13 9 1 10 9 1 10 0 9 1 10 9 15 13 1 10 9 7 13 10 9 1 10 9 2
24 1 9 2 7 1 12 9 2 1 3 9 7 3 1 9 1 9 2 9 9 2 2 9 2
25 1 15 13 10 0 9 15 13 3 2 1 9 1 9 7 9 0 2 10 9 1 9 3 0 2
52 13 3 3 0 10 0 9 2 1 11 12 7 11 12 2 15 13 1 10 11 0 1 10 11 2 0 1 13 9 7 9 1 9 2 1 15 10 9 1 9 3 0 13 3 1 10 9 1 10 10 9 2
16 11 2 3 1 10 9 2 4 13 12 9 7 13 12 9 2
20 13 10 9 1 10 9 1 9 2 15 13 10 9 1 13 2 13 12 9 2
21 1 9 2 10 9 1 9 2 3 10 9 1 10 9 4 13 1 12 9 2 2
8 9 2 9 2 9 2 9 2
23 11 11 2 9 1 10 9 1 10 9 2 4 13 10 9 0 3 12 9 1 9 0 2
10 10 9 1 11 11 13 10 9 0 2
29 2 12 9 1 10 11 2 11 11 11 7 11 11 11 2 4 13 1 10 12 10 9 11 1 4 13 10 9 2
14 10 9 15 2 1 15 13 2 4 13 10 10 9 2
14 2 1 9 13 1 13 1 15 1 10 10 9 2 2
31 3 2 13 10 9 2 1 15 13 0 16 10 11 13 1 10 9 0 1 15 1 11 1 10 9 4 13 10 13 9 2
21 12 2 12 9 1 11 1 10 9 0 2 1 10 10 9 2 1 3 12 9 2
80 11 9 2 9 12 2 11 2 9 12 2 11 2 9 12 2 11 2 9 12 2 11 2 9 12 2 11 0 2 9 12 2 11 2 9 12 2 11 2 9 12 2 11 2 9 12 2 11 2 9 12 2 11 9 9 0 2 9 12 2 9 1 10 9 2 9 12 2 9 2 9 12 2 0 0 0 2 9 12 2
53 3 1 9 2 1 10 9 7 1 10 9 1 9 0 2 7 3 1 10 9 1 10 9 0 7 1 10 9 1 10 9 1 9 16 3 13 1 10 0 9 2 7 2 1 10 10 9 2 1 3 0 9 2
16 2 12 2 10 9 4 13 15 0 1 10 9 1 10 9 2
18 3 13 0 16 1 10 0 9 13 10 9 1 9 2 13 12 2 2
20 3 0 13 10 9 1 10 9 0 1 10 9 15 4 4 13 1 12 9 2
23 10 9 0 1 10 9 1 9 1 0 9 2 12 2 4 13 1 9 0 2 12 2 2
18 15 4 3 13 15 1 15 3 13 0 1 10 9 13 1 10 9 2
61 10 9 1 10 9 3 4 13 10 9 1 9 7 1 9 2 10 9 2 10 9 2 10 9 7 0 9 2 12 2 13 1 10 9 2 12 2 1 10 9 2 12 2 2 16 3 13 10 0 9 2 13 3 9 1 10 9 1 10 9 2
6 12 2 10 9 0 2
12 10 9 0 4 13 1 9 1 10 9 0 2
11 12 2 9 1 9 7 9 1 10 9 2
16 4 3 13 10 9 15 13 1 3 13 10 9 2 12 2 2
15 1 10 9 10 9 1 10 9 13 1 10 10 0 9 2
25 15 4 13 9 1 10 9 4 13 10 9 13 1 10 9 7 2 1 9 2 1 10 9 0 2
11 12 2 12 9 1 10 9 1 0 9 2
19 9 7 9 2 16 13 1 13 15 7 1 13 1 9 2 3 7 3 2
10 12 2 9 1 10 9 1 10 9 2
67 10 9 1 10 9 13 7 13 1 10 9 3 0 2 15 13 3 7 1 10 15 15 3 13 9 2 4 2 16 15 13 2 13 15 9 1 10 9 1 10 10 9 7 1 10 9 1 10 10 9 2 7 4 13 10 9 7 10 9 1 10 9 0 2 12 2 2
7 12 2 9 1 10 9 2
31 10 9 13 16 10 9 13 1 10 9 1 9 1 10 9 15 13 1 10 9 7 3 1 9 1 10 9 1 10 9 2
7 12 2 9 0 1 9 2
5 12 2 9 0 2
38 10 9 13 0 10 9 2 12 2 1 9 1 9 1 10 9 0 1 10 9 2 1 13 15 1 12 9 0 7 1 13 13 1 12 9 10 9 2
16 10 9 7 10 9 1 10 9 1 16 15 4 13 10 9 2
27 10 9 4 13 1 10 9 1 13 15 10 9 1 10 9 13 16 10 9 1 10 9 3 15 4 13 2
21 15 13 10 9 1 13 1 10 15 10 9 1 10 9 15 15 4 13 7 13 2
17 12 2 9 1 10 9 1 10 9 13 1 9 1 10 10 9 2
39 10 9 1 10 9 12 3 15 13 1 10 9 1 15 10 9 13 1 9 1 10 9 1 10 9 2 1 9 7 1 0 9 0 13 1 10 9 0 2
30 1 10 9 4 13 10 9 1 10 9 3 13 2 3 1 10 9 1 10 9 2 12 2 2 12 2 2 12 2 2
45 0 1 0 9 0 7 0 2 10 3 0 7 0 9 1 10 9 0 0 2 2 10 9 1 10 12 4 13 1 13 2 1 10 0 9 2 10 9 0 1 10 9 1 9 2
50 16 10 9 1 10 9 4 4 13 1 10 9 0 2 1 10 13 1 10 9 2 12 2 10 9 1 9 15 13 7 10 9 1 10 9 13 9 1 10 9 2 12 2 2 12 2 2 12 2 2
23 10 9 1 10 9 3 13 2 0 9 0 2 10 9 1 10 9 1 9 2 12 2 2
27 10 9 4 13 1 10 9 1 10 12 1 13 3 1 10 9 0 3 13 1 10 9 0 1 10 11 2
30 10 9 1 9 1 10 9 7 10 9 1 10 9 3 4 13 2 13 10 9 1 10 13 9 2 12 7 0 2 2
9 12 2 9 13 1 10 9 0 2
24 15 4 13 1 10 9 10 9 15 15 4 13 2 12 2 2 0 10 9 13 1 10 9 2
8 12 2 9 2 9 7 9 2
11 10 9 4 3 13 0 9 2 12 2 2
13 12 2 9 1 10 9 7 9 0 1 10 9 2
15 10 0 9 15 13 16 10 9 4 13 3 1 10 9 2
10 12 2 9 1 9 13 1 10 9 2
50 15 13 3 10 9 0 2 12 7 0 2 2 10 9 0 13 2 12 7 0 2 7 10 9 2 12 7 0 2 2 3 16 10 9 2 10 9 7 10 9 4 13 3 16 10 9 4 3 13 2
7 12 2 9 1 10 9 2
10 12 2 9 1 10 9 1 10 9 2
41 7 1 10 9 0 10 9 1 10 9 13 4 13 9 7 13 7 13 10 9 13 2 16 15 13 1 9 1 10 9 2 1 10 10 9 7 1 10 10 9 2
10 1 10 9 7 1 10 9 1 9 2
60 15 13 9 1 13 9 1 9 2 9 2 9 2 9 2 9 7 9 4 2 16 13 0 2 13 7 13 10 9 1 10 9 2 1 10 9 3 1 13 10 9 7 1 13 7 13 10 9 0 1 13 10 9 1 10 9 2 12 2 2
26 16 15 13 10 9 1 10 9 0 2 10 9 4 4 13 1 9 1 10 0 7 1 10 0 9 2
26 7 10 9 0 4 13 10 9 1 10 9 2 13 9 1 10 9 1 10 9 7 1 10 9 13 2
37 1 10 9 1 10 9 7 10 9 1 9 2 10 9 4 13 15 13 1 9 1 13 10 9 1 10 9 13 1 10 0 9 1 10 9 13 2
30 10 9 15 13 2 12 2 12 2 2 16 1 10 0 9 15 13 10 9 1 10 9 13 1 15 1 10 9 13 2
12 10 9 13 10 9 1 9 1 10 9 0 2
27 3 15 13 9 1 10 13 9 1 9 1 10 9 7 9 1 9 2 15 4 4 13 1 10 9 0 2
13 1 10 9 1 10 9 7 1 10 9 1 9 2
18 1 10 9 10 9 13 1 10 9 1 15 4 4 15 13 10 9 2
26 15 4 13 10 9 4 13 1 10 9 1 10 0 9 2 1 10 9 13 1 10 9 1 10 9 2
19 10 9 15 13 1 9 9 1 9 4 13 15 3 1 10 9 1 9 2
35 0 0 9 1 10 9 2 10 9 15 1 10 9 1 10 9 15 13 1 10 9 1 15 2 13 3 1 10 9 0 7 0 1 15 2
22 1 9 1 0 9 1 10 9 2 15 13 10 9 1 10 0 9 1 10 9 0 2
31 10 0 9 15 13 16 2 4 13 10 9 0 2 15 4 13 10 9 2 7 16 13 15 1 10 9 0 1 10 9 2
38 10 0 15 2 1 9 1 10 9 2 15 13 1 10 9 10 9 2 4 13 1 9 1 10 9 0 2 16 10 9 3 13 3 1 13 10 15 2
16 10 9 0 0 15 13 1 10 9 1 10 9 0 3 13 2
25 10 9 7 10 9 1 9 1 9 7 1 9 0 7 1 9 0 7 0 4 13 1 9 0 2
52 15 4 13 1 9 3 1 9 0 1 10 9 0 1 10 9 1 9 2 1 10 15 10 9 1 10 9 3 15 13 2 7 1 10 9 1 9 1 10 9 15 10 9 0 13 1 10 9 1 10 9 2
18 13 10 9 2 10 9 7 10 9 2 13 10 9 0 1 10 9 2
20 9 7 9 13 10 9 1 13 9 7 9 1 9 2 1 9 1 10 9 2
20 13 7 13 10 9 7 10 9 0 13 1 13 7 13 10 9 1 10 9 2
8 13 10 0 7 10 0 9 2
22 13 0 1 9 10 10 9 15 1 10 9 1 10 9 4 13 10 12 9 1 9 2
24 10 9 1 10 9 13 10 9 1 10 9 1 10 9 7 2 1 9 1 15 2 10 9 2
26 10 9 13 1 10 9 1 10 9 1 10 9 7 13 10 9 2 10 9 7 10 9 1 10 9 2
10 10 9 4 13 1 9 1 10 9 2
5 10 9 13 0 2
8 10 9 15 13 10 0 9 2
60 10 9 2 16 13 16 10 9 7 10 9 13 9 1 9 1 10 9 7 1 10 0 9 13 10 10 9 1 9 2 4 13 10 9 1 9 0 3 1 10 9 0 1 12 9 1 10 9 1 10 9 7 1 10 9 13 9 1 9 2
43 3 1 16 3 13 1 9 10 9 0 2 10 9 1 10 9 13 1 10 9 12 13 9 1 10 9 7 1 10 9 1 10 9 0 1 10 9 1 9 1 10 9 2
46 1 9 1 10 9 12 2 4 13 1 9 2 1 3 3 10 9 1 10 9 1 9 1 10 9 2 9 0 1 10 9 1 9 7 1 10 9 1 10 9 0 1 10 9 0 2
58 2 12 2 10 9 15 13 9 7 13 1 10 9 1 10 9 0 13 1 10 9 1 9 1 10 0 9 4 4 13 1 10 9 11 7 1 10 13 9 2 1 10 9 1 13 10 10 9 1 10 9 0 7 10 10 0 9 2
68 9 1 9 1 10 9 15 13 1 10 9 9 3 13 10 9 1 10 9 1 10 9 15 13 7 13 10 9 1 10 9 1 10 12 9 12 2 15 13 10 9 1 9 1 9 1 9 2 9 7 9 1 10 9 1 10 9 1 10 9 0 2 9 2 11 2 2 2
27 15 1 10 9 4 13 1 10 9 1 10 9 2 1 9 1 10 9 9 2 1 10 9 1 10 9 2
38 10 9 1 9 13 1 3 12 9 1 10 9 7 1 10 0 12 1 9 0 1 11 7 10 9 1 10 11 15 13 10 10 9 1 10 9 0 2
42 15 4 13 1 10 9 1 11 11 2 12 9 2 15 1 10 12 9 1 10 9 1 9 2 16 1 10 9 1 10 9 1 9 4 13 10 9 1 10 9 0 2
10 10 9 15 13 2 7 3 15 13 2
27 13 10 9 1 10 12 9 16 1 3 4 13 10 9 13 1 10 9 0 1 12 9 1 9 1 9 2
53 16 10 9 1 9 1 10 9 1 10 9 4 13 10 9 1 10 9 2 13 13 3 3 1 10 9 1 10 9 2 10 9 15 4 13 1 9 7 9 1 10 9 1 11 3 15 4 13 3 12 9 13 2
33 1 10 9 1 10 9 1 9 2 13 1 11 3 12 9 3 2 10 9 1 9 4 13 10 0 9 1 9 1 9 7 9 2
23 1 10 9 10 9 1 10 9 1 10 0 9 13 3 10 9 1 13 9 7 13 9 2
12 3 10 9 13 1 10 9 1 10 10 9 2
38 10 9 4 13 16 4 13 10 9 0 7 0 1 13 0 9 1 9 2 0 1 15 15 1 10 9 0 2 1 10 9 1 10 9 1 10 9 2
13 1 15 4 13 15 10 9 1 2 9 0 2 2
27 15 3 4 13 9 0 3 1 15 7 1 10 9 11 11 7 0 9 1 10 9 7 1 10 9 0 2
16 3 10 9 1 12 13 3 1 10 9 1 10 9 1 11 2
12 10 9 1 10 11 13 1 13 10 0 9 2
12 13 1 12 9 10 9 1 10 9 1 9 2
44 10 9 11 11 2 15 1 10 9 1 10 10 9 0 13 1 9 1 10 9 1 10 9 11 2 4 13 3 10 9 0 1 13 3 1 3 10 9 1 10 0 9 0 2
77 10 9 2 13 1 10 9 1 10 0 9 1 11 11 2 7 13 3 1 10 10 9 1 10 9 0 2 4 13 1 10 0 9 1 10 9 1 3 16 10 9 1 10 9 0 0 11 11 4 13 10 9 1 11 1 1 9 10 9 2 3 15 1 12 2 7 10 9 1 10 9 9 1 9 11 11 2
59 16 10 12 9 4 13 10 9 13 2 10 9 1 9 1 10 9 15 4 13 1 9 7 4 13 10 9 0 1 11 2 13 2 1 10 9 1 10 9 1 10 11 11 2 10 9 1 9 7 9 15 4 4 3 13 1 10 9 2
10 10 10 9 4 4 3 13 1 11 2
43 13 15 1 10 9 10 10 9 4 13 3 1 10 9 0 10 9 1 9 0 7 1 0 9 15 15 13 1 0 9 1 9 1 9 1 10 9 0 2 3 3 0 2
23 10 11 11 13 3 1 13 10 10 0 9 0 9 0 2 16 15 13 10 10 9 0 2
52 1 15 4 13 13 1 10 0 9 10 9 2 9 1 10 9 7 10 0 9 15 4 13 3 1 10 9 3 1 9 0 2 3 1 10 9 1 10 9 0 2 3 10 9 13 9 10 9 11 2 11 2
26 10 9 13 10 0 9 1 10 9 7 13 1 9 1 9 10 9 1 9 0 13 13 10 10 9 2
21 1 15 4 13 10 9 1 0 9 0 0 15 4 13 10 9 13 1 10 9 2
34 10 15 13 3 1 16 13 3 3 0 10 9 2 15 10 9 1 10 9 13 3 1 13 1 10 9 2 2 1 10 9 1 9 2
13 15 15 13 10 11 1 10 11 13 3 10 9 2
12 10 11 15 4 13 16 1 13 13 3 13 2
32 10 9 1 9 1 10 9 1 9 1 10 9 11 4 13 1 10 9 1 10 9 7 4 13 10 9 1 3 1 10 9 2
21 10 9 13 10 9 13 1 10 9 1 10 9 1 10 9 13 1 10 9 0 2
10 3 11 7 11 4 13 1 10 9 2
15 13 1 13 15 2 3 2 10 9 1 10 9 1 9 2
41 10 9 11 11 4 13 10 9 1 10 11 10 9 1 10 11 11 11 2 1 10 15 15 4 2 3 2 13 2 1 10 9 1 10 0 9 2 1 10 0 2
28 11 11 4 13 10 12 5 1 10 9 1 10 0 9 2 13 1 10 0 11 11 15 4 13 10 12 5 2
16 1 10 11 2 10 0 9 13 1 9 1 10 9 15 13 2
14 16 13 1 10 9 2 16 15 13 3 13 1 13 2
23 7 1 10 9 2 1 10 0 9 1 10 9 1 10 10 9 11 2 15 13 9 0 2
15 7 15 13 3 15 13 10 0 9 1 10 10 9 0 2
26 1 10 9 1 9 0 3 10 9 0 3 15 13 3 1 9 1 10 9 0 7 1 10 9 0 2
32 10 9 1 10 9 0 2 13 16 11 11 2 10 9 0 1 10 11 11 2 13 3 1 9 10 0 9 1 10 10 9 2
16 2 10 9 13 15 2 3 11 7 3 13 10 9 0 2 2
36 10 9 13 16 3 10 9 0 4 13 1 9 15 3 13 15 1 16 13 1 10 9 1 10 9 7 13 10 9 15 3 10 9 4 13 2
36 1 11 1 9 2 10 11 11 4 13 10 0 9 1 10 11 2 12 2 12 2 2 13 10 9 15 15 13 0 3 3 9 1 10 9 2
14 9 1 9 1 10 9 1 10 11 1 10 9 0 2
14 10 9 0 13 9 1 10 2 11 2 15 15 13 2
25 1 13 10 9 4 13 10 9 1 10 9 10 15 4 13 13 12 9 1 10 9 1 10 9 2
13 1 10 9 1 9 0 10 9 13 2 7 3 2
46 7 10 9 13 13 2 13 10 9 1 10 9 1 10 0 9 1 10 11 13 3 1 11 11 7 2 1 9 3 0 2 1 11 2 1 10 9 1 9 7 9 1 10 0 9 2
42 1 12 9 15 13 10 9 0 1 10 9 1 11 2 10 9 3 0 1 10 0 9 13 1 9 1 10 10 0 9 1 10 3 0 9 1 10 9 2 15 0 2
6 2 0 15 15 13 2
24 10 9 1 9 4 13 2 1 9 2 1 10 0 9 1 10 9 15 4 13 1 10 9 2
31 9 4 13 10 9 1 10 9 1 10 9 11 11 1 13 11 7 9 2 3 2 11 4 13 10 9 1 10 11 11 2
52 10 9 7 10 9 1 10 13 13 1 10 9 1 13 1 10 9 0 10 9 2 15 1 10 9 13 0 7 1 10 9 13 1 10 9 7 1 10 9 2 0 9 1 10 9 1 10 9 13 1 9 2
50 10 9 1 9 1 10 0 9 0 4 13 3 1 13 1 10 12 9 1 0 9 7 10 12 9 1 0 9 10 9 0 2 13 1 13 10 9 1 9 1 12 9 1 9 0 1 11 7 11 2
7 13 10 9 1 10 9 2
11 1 0 2 10 9 13 1 10 9 0 2
14 1 10 10 9 13 1 10 15 11 11 7 10 11 2
32 3 1 10 0 9 0 2 9 0 2 0 7 0 2 7 3 0 2 13 1 13 10 9 1 9 1 9 1 10 9 0 2
18 10 9 2 9 2 9 2 15 13 10 9 1 9 1 10 0 9 2
40 10 9 13 0 1 10 9 1 10 9 7 1 10 9 0 2 13 1 10 9 7 1 10 9 0 7 3 0 2 7 3 1 10 9 7 1 10 9 0 2
32 9 1 10 9 2 10 9 2 10 9 1 9 7 10 9 2 4 13 1 10 9 1 10 9 1 10 9 3 13 10 9 2
12 10 9 1 10 9 1 10 9 13 3 0 2
35 1 10 12 10 9 0 1 10 9 2 15 13 1 10 9 1 11 1 15 1 11 2 4 13 7 13 10 9 1 11 11 2 11 2 2
53 10 9 4 13 1 10 12 1 10 9 1 10 9 1 10 9 1 11 7 10 9 1 11 2 13 10 9 15 13 1 10 9 1 10 9 1 10 9 13 1 10 9 0 1 11 7 1 10 9 1 10 9 2
30 1 10 0 9 4 13 3 10 9 0 1 10 9 9 1 10 9 2 1 11 7 11 2 13 1 10 9 1 9 2
33 1 10 9 2 10 9 11 13 10 9 3 0 2 16 13 1 10 9 10 9 13 10 9 1 9 1 11 2 3 1 13 11 2
29 10 9 11 11 13 10 9 1 9 0 15 13 13 11 7 11 11 1 10 9 0 7 1 10 9 1 10 9 2
43 0 1 10 9 13 2 11 1 10 9 12 13 1 10 3 9 1 10 9 11 11 2 10 9 1 13 1 9 10 9 1 9 7 9 3 0 1 10 9 3 15 0 2
62 10 0 9 0 1 10 9 1 10 11 11 12 1 10 9 0 13 10 9 1 10 11 1 10 3 3 0 9 1 10 11 15 13 1 10 9 1 10 9 1 10 9 1 9 1 10 9 1 9 11 1 13 1 10 12 9 12 1 10 11 12 2
13 10 9 15 13 1 10 9 1 9 1 10 9 2
27 1 1 10 9 2 10 9 1 10 9 4 13 1 10 9 1 9 7 9 7 1 10 9 1 10 9 2
36 10 9 1 9 3 3 13 1 10 9 7 3 1 10 9 2 10 9 0 15 13 1 9 1 13 15 1 10 9 7 10 9 1 10 9 2
11 10 9 13 10 9 15 15 13 3 3 2
36 9 2 10 9 16 13 10 9 0 1 9 1 13 10 9 15 13 7 2 1 10 9 2 10 9 9 1 9 1 10 9 1 9 1 9 2
47 0 2 9 2 9 7 9 1 9 1 10 9 0 1 10 9 7 1 10 9 7 2 16 3 13 2 9 2 9 7 9 1 9 1 10 9 0 0 1 13 10 9 1 9 1 9 2
39 0 2 10 9 13 1 10 9 1 9 15 13 1 10 9 1 10 9 1 9 7 9 2 3 1 10 9 16 15 13 1 10 9 1 9 7 1 9 2
59 10 9 13 1 10 9 1 15 1 10 9 12 3 1 10 9 1 10 9 1 9 2 16 10 9 4 4 13 1 9 1 10 9 13 10 9 1 9 1 9 15 3 13 1 13 10 9 0 7 10 9 1 10 9 1 10 9 12 2
47 10 9 1 10 9 1 15 1 10 9 0 3 13 10 9 7 10 9 1 10 9 1 9 2 10 15 13 3 9 1 10 9 1 10 0 9 2 3 0 15 13 10 9 1 10 9 2
13 9 2 10 9 13 1 10 9 7 1 9 0 2
13 13 10 9 1 10 11 0 7 0 2 12 2 2
13 10 9 0 1 10 9 13 3 13 1 10 11 2
11 10 9 4 13 1 4 13 10 9 0 2
6 3 4 13 11 11 2
8 10 15 4 13 10 9 11 2
8 15 13 10 0 9 1 11 2
14 15 4 13 10 9 2 9 0 1 10 0 9 2 2
9 10 15 13 10 2 9 11 2 2
9 1 10 9 4 13 10 9 9 2
9 3 4 13 10 9 1 10 11 2
15 1 10 9 10 9 0 4 13 10 2 11 11 11 2 2
7 13 10 9 1 10 9 2
11 1 10 9 1 9 0 13 9 11 11 2
5 3 13 11 11 2
11 15 13 10 3 0 9 1 10 9 0 2
8 15 4 13 10 11 1 11 2
6 10 15 13 10 11 2
8 15 13 10 9 1 10 11 2
11 3 13 10 9 0 1 10 11 11 11 2
9 15 13 10 9 1 10 9 0 2
10 10 9 15 13 1 13 10 9 0 2
13 3 4 13 10 9 0 1 10 9 1 10 11 2
8 1 10 9 15 13 11 11 2
8 15 13 10 9 1 10 11 2
9 1 15 13 10 9 1 10 11 2
5 15 13 11 11 2
10 10 9 4 13 10 9 1 10 11 2
11 10 9 0 13 1 10 11 11 1 11 2
11 1 10 9 1 11 15 13 10 11 11 2
12 15 13 10 9 1 10 9 0 11 1 11 2
11 15 13 10 9 0 1 9 1 10 9 2
7 15 13 0 10 9 11 2
10 1 10 9 15 13 10 11 1 11 2
6 15 13 0 10 11 2
18 15 4 13 10 9 9 1 10 9 1 11 1 13 9 1 9 0 2
11 1 10 9 1 9 13 10 9 11 11 2
10 13 10 9 1 15 4 13 11 11 2
5 3 15 13 11 2
7 1 10 9 13 11 11 2
5 3 13 11 11 2
13 15 13 10 11 1 2 10 11 7 10 11 2 2
11 15 13 10 9 1 10 11 11 11 0 2
9 15 13 10 9 0 1 10 11 2
6 15 13 1 11 11 2
9 15 13 10 9 1 10 11 11 2
6 10 9 13 10 0 2
16 10 9 13 11 11 1 10 9 15 15 13 1 13 10 9 2
5 3 13 11 11 2
9 3 15 13 10 11 1 10 9 2
9 10 9 0 15 13 1 10 9 2
10 3 15 13 10 9 1 11 11 11 2
13 3 13 11 2 11 11 2 1 11 2 11 11 2
22 1 10 9 10 9 11 13 10 9 1 10 9 1 10 9 1 10 9 1 11 11 2
10 3 4 13 10 9 1 10 11 0 2
6 10 9 13 11 11 2
12 10 9 13 11 11 3 1 13 1 13 9 2
9 10 9 0 15 13 1 10 9 2
11 3 4 13 10 9 1 13 1 10 9 2
8 1 10 15 4 13 10 11 2
24 10 2 8 8 2 4 13 11 2 11 2 11 1 10 9 1 10 10 9 1 10 9 0 2
14 10 9 4 13 10 9 1 9 1 15 13 10 9 2
6 15 13 10 9 0 2
10 10 0 4 13 10 9 0 1 9 2
19 10 9 13 10 9 1 10 10 9 0 1 10 9 2 11 1 3 2 2
5 15 13 11 11 2
17 3 15 13 10 9 15 13 3 0 1 4 13 1 10 9 0 2
11 10 9 13 10 11 11 11 1 11 11 2
17 10 9 0 13 1 10 9 0 15 13 1 10 9 1 10 9 2
6 3 4 13 10 11 2
5 15 13 11 11 2
8 3 4 4 13 10 11 11 2
7 1 15 4 13 10 9 2
7 1 15 4 13 10 9 2
17 10 9 1 10 9 11 7 11 4 13 3 9 1 10 11 11 2
37 13 15 1 10 9 1 10 9 1 9 13 1 10 11 1 11 1 9 1 11 11 11 2 10 9 1 10 11 3 1 9 1 9 1 9 0 2
24 10 9 1 9 1 9 1 9 4 4 13 1 10 9 1 11 1 10 9 1 10 9 11 2
24 10 9 1 11 2 9 0 1 9 1 11 11 2 10 0 9 1 11 11 7 9 1 11 2
29 10 9 15 15 13 13 9 1 10 9 1 10 9 1 9 0 13 15 1 11 11 2 3 1 10 9 1 11 2
13 1 10 12 4 4 13 9 0 1 10 0 11 2
22 1 9 1 11 11 11 11 3 11 11 2 15 13 10 9 1 9 1 10 9 0 2
14 10 9 1 11 11 15 4 13 10 9 4 4 13 2
26 11 11 2 15 1 10 9 4 13 1 10 11 11 11 2 13 3 3 7 0 3 1 10 0 11 2
30 10 9 4 13 3 1 10 9 1 0 9 0 1 11 11 11 7 1 11 7 2 3 4 13 3 1 10 9 2 2
28 15 1 10 9 7 9 1 11 11 2 11 11 2 13 13 1 13 10 0 9 1 9 13 1 10 10 9 2
25 11 13 0 1 9 15 13 2 7 3 1 9 15 3 13 9 7 13 9 0 7 1 9 0 2
26 15 4 13 1 13 12 9 2 15 4 13 13 2 13 2 15 4 13 10 9 7 13 1 10 12 2
21 10 9 3 13 1 4 13 1 9 7 13 3 10 9 2 2 13 9 11 11 2
25 10 9 11 11 2 1 9 2 11 11 2 2 3 13 10 9 0 7 3 13 9 1 9 0 2
37 10 9 2 1 3 13 2 4 13 1 9 1 10 9 1 10 9 1 10 0 9 2 11 11 11 11 2 2 2 11 2 7 2 9 2 2 2
5 9 1 9 9 2
58 1 10 9 1 13 9 2 4 13 16 10 11 13 1 10 9 0 1 13 10 9 1 15 13 1 10 9 0 1 10 9 1 9 2 1 9 2 1 10 9 1 10 9 1 10 9 1 9 0 0 9 12 9 12 5 12 2 2
23 10 9 1 10 9 13 7 13 10 9 1 10 9 1 15 15 13 1 9 7 9 0 2
19 3 2 10 9 1 10 10 9 4 4 13 1 9 0 1 9 3 0 2
23 4 13 16 15 13 10 9 1 10 9 1 10 0 9 2 1 10 9 1 10 0 9 2
68 10 9 11 1 10 9 1 9 0 4 13 1 10 9 1 10 9 1 10 11 1 9 7 1 10 9 12 13 10 9 13 1 13 10 9 1 9 1 9 1 10 9 1 10 9 15 3 13 1 13 10 10 9 1 9 0 1 10 9 2 1 10 9 1 10 9 0 2
12 13 1 9 16 4 13 0 3 10 9 0 2
10 0 9 2 13 10 9 13 10 9 2
19 0 9 11 11 2 15 3 4 4 13 9 0 1 10 9 1 10 9 2
15 2 9 1 10 9 1 10 9 1 10 11 2 11 2 2
13 3 2 15 13 10 0 9 1 9 1 10 9 2
9 4 3 13 15 1 10 0 9 2
13 9 9 2 0 9 2 0 9 7 0 0 9 2
27 4 13 3 10 9 13 1 10 9 1 9 1 10 9 1 10 9 1 10 9 1 9 1 10 9 0 2
16 1 10 9 11 13 10 10 9 1 10 9 13 1 10 9 2
25 1 10 9 1 10 9 15 13 9 1 10 9 16 1 10 9 0 1 10 9 4 13 3 0 2
50 4 13 1 10 9 16 3 13 1 9 1 13 15 15 1 10 9 1 9 1 10 9 1 9 1 9 1 10 12 9 0 7 16 10 11 11 13 10 9 1 13 10 9 13 9 10 3 0 0 2
40 15 13 15 16 10 9 0 1 9 2 11 2 3 4 13 1 13 1 10 9 13 10 9 1 10 9 0 1 13 1 10 9 0 1 9 1 10 11 11 2
15 10 9 13 3 10 12 9 1 10 9 1 10 9 0 2
23 13 16 10 9 1 10 9 13 1 9 1 10 9 0 1 10 9 7 1 10 10 9 2
33 10 9 1 10 9 2 13 1 10 9 1 10 9 2 4 4 3 13 1 9 1 10 9 1 10 9 0 7 1 10 9 0 2
42 10 9 13 1 9 1 10 9 1 9 13 1 10 9 1 9 7 1 9 1 10 11 10 9 0 1 10 9 1 11 7 13 3 1 10 9 1 10 9 1 9 2
21 10 0 9 13 1 10 9 2 15 3 13 9 0 7 1 9 1 9 7 0 2
11 10 9 0 4 13 3 1 13 10 9 2
44 13 16 10 9 1 10 9 0 1 10 10 9 1 10 9 0 7 1 10 10 9 2 0 7 0 2 13 10 9 1 10 9 2 1 10 9 7 1 10 9 1 10 9 2
8 10 9 13 9 1 10 9 2
47 3 2 16 13 1 13 11 1 10 0 9 2 13 0 16 13 15 1 4 13 10 0 9 13 1 10 9 1 11 7 5 7 1 10 9 1 9 1 15 13 1 10 9 1 9 0 2
27 1 13 15 1 10 0 9 2 13 10 10 9 2 9 1 9 2 9 7 9 9 1 10 9 0 3 2
17 11 1 9 1 10 12 5 1 10 9 13 1 10 9 1 11 2
13 13 0 1 10 10 9 0 2 15 13 3 0 2
16 11 13 9 1 13 15 1 10 9 0 1 10 9 1 9 2
34 1 10 9 1 10 10 9 11 15 13 13 1 10 9 1 13 13 12 9 2 12 11 2 1 9 1 11 1 13 7 13 1 11 2
16 16 15 13 10 9 2 13 1 10 9 1 10 9 7 13 2
34 1 11 13 10 9 1 10 9 2 11 13 10 3 2 9 1 9 0 2 3 16 13 1 10 9 1 10 9 3 0 1 10 9 2
26 11 11 11 2 12 2 7 11 11 11 2 12 2 13 10 9 1 11 11 11 2 10 9 0 2 2
16 10 10 9 13 13 10 0 9 1 9 2 0 9 7 9 2
30 16 13 7 13 9 1 10 9 0 1 10 9 0 11 11 2 11 13 1 13 10 9 0 1 10 9 1 10 9 2
37 10 9 13 10 9 1 11 10 9 1 10 9 2 10 9 3 0 7 0 1 10 9 2 15 13 1 13 10 9 0 1 3 13 1 10 9 2
16 2 1 10 0 9 2 10 9 13 10 9 0 1 9 0 2
31 1 9 1 10 9 1 10 0 9 1 10 9 1 2 9 0 0 2 2 11 13 16 2 10 9 4 13 1 15 2 2
18 1 10 9 1 12 9 2 13 11 11 2 1 10 15 13 12 9 2
27 11 13 10 9 7 10 9 13 1 10 10 9 7 10 10 9 3 13 10 9 0 1 1 10 0 9 2
24 10 10 9 0 1 9 13 9 2 7 3 15 15 13 10 12 9 2 10 9 1 0 11 2
28 1 10 12 2 10 9 1 9 1 10 9 13 10 10 9 2 15 13 11 1 10 9 9 1 10 9 11 2
20 9 1 10 9 0 7 1 10 9 1 11 13 16 10 9 15 4 13 9 2
30 1 10 12 2 15 13 1 0 1 9 1 10 9 2 1 10 9 1 9 1 10 9 1 11 11 1 10 9 0 2
21 3 13 9 1 10 9 0 13 11 11 2 10 9 1 9 1 9 7 0 9 2
28 1 10 12 2 4 13 1 9 1 11 1 11 2 10 9 15 13 10 9 0 1 10 9 1 11 2 11 2
26 10 15 0 12 9 0 13 10 9 2 3 1 11 11 2 15 15 13 1 9 0 1 10 11 11 2
12 2 13 7 3 13 2 15 13 10 9 2 2
24 1 10 12 2 11 11 11 13 16 10 11 0 2 4 13 1 0 9 1 9 7 9 2 2
11 10 9 13 12 9 2 1 15 12 0 2
11 15 13 1 11 11 2 10 9 1 11 2
26 15 13 12 9 13 1 11 11 2 11 7 11 2 10 10 9 0 13 0 1 15 1 10 9 0 2
40 1 10 9 1 11 2 10 9 0 2 10 9 7 10 9 13 3 0 1 15 3 15 13 3 2 7 10 10 9 1 10 9 4 13 1 13 10 9 0 2
29 1 10 9 12 2 10 9 1 0 9 0 13 10 9 7 13 10 9 1 10 9 2 0 2 0 2 1 11 2
13 1 12 9 13 10 0 11 11 2 15 13 0 2
36 1 10 0 0 9 2 11 11 13 12 1 10 0 9 1 11 1 9 2 7 1 10 9 13 13 15 9 2 10 9 1 11 4 3 13 2
5 3 2 13 15 2
36 10 9 1 11 2 11 2 11 2 1 10 15 2 4 13 10 9 1 9 0 7 13 16 4 4 13 0 9 2 1 10 11 1 10 11 2
13 1 0 9 2 10 9 1 9 13 13 9 0 2
29 13 0 1 9 1 10 9 1 10 9 13 13 16 10 0 9 0 13 10 10 9 1 9 1 9 0 13 3 2
34 7 10 9 13 16 10 9 13 1 10 9 1 9 0 13 10 9 1 10 9 7 1 10 9 0 7 1 10 9 1 9 1 9 2
29 13 3 16 10 9 0 13 10 9 0 15 10 9 0 4 13 1 10 13 10 9 7 13 10 9 1 10 9 2
43 11 11 2 15 1 10 9 1 10 11 13 1 11 2 4 13 10 9 0 1 10 9 0 2 13 10 2 10 9 7 1 13 7 1 13 0 9 1 9 3 0 2 2
20 10 9 1 10 9 3 13 0 1 13 2 7 10 9 1 10 9 13 0 2
19 10 9 13 10 9 1 13 9 0 16 10 9 0 4 13 9 3 0 2
38 7 16 10 9 13 1 13 15 10 9 0 1 10 9 0 7 10 9 2 4 13 3 0 0 1 10 12 2 7 3 3 9 0 2 9 1 3 2
14 1 11 2 10 9 0 4 13 15 1 9 7 9 2
38 10 11 4 13 10 0 9 1 9 2 13 15 1 10 9 1 9 1 13 15 1 10 9 0 1 10 9 7 1 10 9 1 9 2 9 7 9 2
37 3 4 13 10 9 1 10 9 1 10 9 2 3 1 10 9 1 9 0 3 10 9 0 0 7 10 9 1 10 9 1 10 0 13 3 0 2
23 10 9 0 1 10 9 13 10 9 1 10 9 13 1 10 9 10 9 0 1 10 9 2
19 7 16 10 9 13 1 10 9 1 10 9 2 10 9 13 3 3 0 2
27 10 9 15 13 10 9 0 7 0 13 7 13 1 10 9 1 10 9 3 3 1 10 10 9 3 0 2
62 1 9 2 10 10 9 0 1 10 9 0 2 13 1 10 9 1 9 2 13 1 13 10 9 1 9 0 1 1 10 12 5 1 10 12 2 1 9 1 10 9 1 9 1 10 9 1 0 9 7 1 9 0 7 10 9 1 10 9 0 13 2
19 10 11 15 13 1 10 9 1 13 10 9 1 10 10 9 1 10 9 2
35 10 0 9 10 9 1 10 11 4 13 1 13 3 10 0 9 2 10 0 9 0 1 10 9 0 1 10 10 13 9 1 13 10 9 2
27 1 9 1 10 9 2 15 13 3 12 12 9 1 9 0 1 10 9 15 13 12 12 9 1 9 0 2
29 3 1 10 9 0 7 0 1 10 9 10 9 4 13 1 9 10 9 1 10 9 0 1 10 9 1 10 9 2
27 13 10 11 1 10 9 0 0 1 13 3 10 11 2 10 10 9 4 13 3 13 9 1 10 9 0 2
