26491 17
40 10 3 1 15 7 10 3 0 3 3 13 1 9 9 0 13 2 1 7 9 15 1 0 13 15 13 13 3 0 13 13 3 1 10 9 7 1 10 15 2
23 1 3 9 9 10 3 9 15 0 13 9 13 1 15 13 2 7 3 1 0 3 13 2
18 10 3 9 1 10 1 0 1 10 0 0 13 9 13 10 0 3 2
18 3 9 0 10 9 3 0 13 1 10 9 1 10 15 3 3 13 2
47 1 3 10 0 9 10 9 7 9 13 1 9 10 0 3 0 13 13 2 7 9 13 3 1 0 0 3 13 9 9 10 9 2 16 3 1 9 0 3 3 0 13 10 9 9 13 2
11 13 3 15 3 15 10 0 9 3 0 2
12 1 3 10 0 15 13 0 3 13 10 9 2
5 13 3 3 9 2
21 3 3 3 9 13 1 10 3 9 3 2 16 15 13 2 0 1 9 9 13 2
28 10 3 3 3 0 9 1 9 3 0 15 13 7 0 9 13 15 1 10 0 1 9 7 9 15 0 13 2
11 3 3 0 10 9 9 3 0 13 13 2
22 10 3 0 2 16 13 2 13 1 10 9 1 0 13 2 10 10 9 3 13 15 2
7 13 3 3 1 9 15 2
24 3 1 15 0 10 9 10 0 9 13 1 3 9 10 9 3 9 3 9 7 10 3 9 2
12 10 3 13 0 10 9 1 10 0 9 13 2
17 9 3 13 15 10 9 3 3 13 10 3 3 1 0 0 9 2
18 1 10 0 3 9 10 3 9 13 7 13 10 9 1 10 0 13 2
30 3 10 0 15 10 0 1 10 0 3 0 9 16 9 3 0 13 13 7 0 9 9 9 13 10 1 10 9 9 2
16 1 15 3 9 10 0 1 10 0 1 0 0 10 9 13 2
27 0 3 3 9 3 1 10 3 9 0 9 13 3 1 10 15 1 10 0 10 10 0 13 0 3 13 2
14 13 3 0 7 1 10 0 13 9 1 10 13 13 2
24 10 3 3 3 1 10 0 9 9 13 1 10 9 10 9 13 2 7 3 0 9 16 13 2
26 3 3 3 1 10 9 13 15 3 2 7 3 10 0 2 9 7 9 9 13 2 7 13 15 13 2
16 0 3 3 7 15 15 13 10 0 0 0 10 3 0 13 2
14 3 3 0 9 13 10 9 2 9 3 13 7 9 2
9 15 3 3 10 0 10 9 13 2
41 9 3 13 1 9 1 0 10 9 7 10 9 13 0 13 10 13 1 10 9 2 1 0 9 13 2 13 10 3 9 10 9 13 7 10 9 15 3 3 13 2
14 3 1 0 10 9 3 3 13 0 9 1 9 13 2
23 9 3 15 13 10 3 9 13 7 3 15 10 9 9 13 10 9 9 13 10 9 13 2
21 13 3 9 3 0 15 13 7 9 13 2 16 9 15 13 2 16 15 0 13 2
16 3 1 10 9 3 10 9 13 15 0 9 7 9 0 13 2
13 13 3 13 3 0 10 9 0 13 10 1 15 2
41 3 16 3 9 0 13 2 7 16 0 10 3 9 3 3 0 13 13 2 3 0 3 15 9 13 13 3 13 10 9 0 0 10 3 9 13 7 10 9 13 2
60 3 13 13 2 3 10 9 10 9 3 13 16 10 9 2 13 7 10 9 0 0 3 13 10 1 15 2 13 7 10 3 2 10 9 3 9 16 15 13 3 3 13 2 15 13 1 10 0 3 9 13 13 2 3 7 13 3 3 0 2
10 15 3 9 1 1 9 9 3 13 2
14 9 3 16 13 3 0 0 2 1 10 9 9 13 2
7 9 3 0 13 10 0 2
39 9 3 3 13 0 13 1 10 9 7 10 3 1 9 2 3 3 7 13 9 13 1 9 0 2 3 3 10 9 0 13 2 7 10 0 9 0 13 2
24 1 10 0 3 3 7 0 9 10 0 13 3 0 13 13 2 3 1 0 10 9 3 13 2
11 0 3 13 3 10 9 15 0 10 9 2
19 15 3 3 10 9 15 13 10 0 9 13 9 2 10 3 13 0 13 2
51 9 3 16 13 13 9 7 13 0 1 9 7 9 3 10 9 13 2 3 3 9 13 13 2 10 3 3 3 0 2 7 9 10 3 13 13 2 9 7 3 13 1 0 3 9 7 0 10 9 13 2
38 3 1 9 10 3 1 15 0 13 7 0 3 3 15 2 0 10 3 13 2 13 10 9 0 13 10 9 7 10 3 1 15 1 10 9 9 13 2
18 3 3 1 10 0 10 9 3 13 3 7 13 2 16 3 13 13 2
30 10 3 3 9 10 9 1 9 0 13 0 13 2 7 9 1 10 9 3 1 0 13 2 1 15 13 10 9 13 2
40 3 3 1 0 9 13 10 9 3 7 3 13 9 13 2 7 9 3 9 7 9 10 0 13 2 9 7 7 9 10 0 9 10 7 0 9 13 0 9 2
8 0 3 15 9 10 0 13 2
23 0 3 9 13 0 10 3 9 13 10 1 10 9 2 7 9 1 9 0 10 9 13 2
11 13 3 3 9 9 0 9 9 13 9 2
16 9 3 13 3 0 1 10 9 0 10 9 16 9 9 13 2
10 9 3 0 15 13 13 9 1 9 2
14 9 3 3 3 15 0 7 0 13 1 10 0 9 2
6 0 3 13 10 9 2
25 16 3 10 9 3 13 2 10 9 13 10 0 13 2 7 9 13 0 0 13 9 9 10 9 2
28 3 9 9 0 13 0 1 9 9 0 13 7 9 10 9 15 2 10 7 1 15 9 9 13 13 0 9 2
23 3 9 9 13 1 9 0 13 15 3 10 9 0 13 7 9 13 13 10 9 10 0 2
8 9 3 9 13 9 13 13 2
7 0 3 15 10 0 13 2
25 13 3 3 15 0 9 9 13 10 0 9 3 0 13 2 9 7 3 7 9 0 13 16 15 2
28 0 3 1 10 0 7 10 9 9 2 15 1 9 9 13 2 9 1 3 9 10 9 1 9 13 7 9 2
14 15 3 0 1 10 9 9 0 0 1 10 9 13 2
19 9 3 7 9 2 3 16 0 15 2 0 13 2 7 15 10 0 9 2
24 3 3 1 15 9 9 13 9 13 2 7 3 10 0 0 13 2 10 9 13 15 3 13 2
8 3 15 3 13 1 0 9 2
17 10 3 3 0 10 9 15 13 2 10 3 0 7 10 0 13 2
16 9 3 13 3 3 0 10 13 15 9 3 9 7 15 9 2
14 13 3 10 9 13 2 3 3 0 3 0 13 9 2
14 1 9 3 9 2 3 0 3 9 13 2 0 13 2
29 0 3 13 2 0 3 13 2 1 0 10 0 0 2 7 0 9 0 1 10 15 1 15 9 3 13 10 9 2
20 3 3 1 10 3 3 13 9 9 7 0 3 10 0 0 1 9 0 13 2
52 9 3 0 13 1 10 0 9 2 10 1 15 0 13 1 3 10 9 7 1 10 10 0 9 13 1 9 0 13 3 10 9 13 2 13 7 0 1 15 9 0 2 16 3 7 15 1 0 10 15 0 2
9 10 3 1 9 1 0 13 9 2
20 3 3 10 9 1 0 9 13 3 3 0 15 13 2 1 9 7 0 13 2
17 0 3 9 1 15 3 10 0 10 0 9 1 10 9 13 13 2
33 3 0 9 13 10 3 9 10 13 9 13 9 13 2 7 10 9 13 10 9 13 13 10 9 7 13 1 10 9 13 0 13 2
24 3 3 13 10 0 2 0 3 0 13 1 3 9 7 9 10 3 13 9 9 7 10 13 2
6 9 3 15 0 13 2
11 13 3 10 3 1 9 2 10 7 9 2
21 3 0 3 9 13 10 9 2 16 13 10 9 7 9 13 1 10 0 1 15 2
14 3 10 0 9 16 15 3 13 2 1 15 3 13 2
44 3 10 3 9 3 0 13 9 10 0 13 2 1 9 7 15 0 0 3 16 13 13 2 9 7 9 3 10 9 10 9 13 1 9 7 9 2 7 9 10 0 13 13 2
22 3 13 15 1 0 10 9 10 0 9 0 16 3 10 0 3 1 0 10 9 13 2
14 10 3 3 0 0 13 2 0 13 0 3 9 13 2
20 10 3 9 10 9 10 13 2 3 16 0 15 13 2 3 3 1 15 13 2
46 0 3 7 15 3 3 3 9 7 3 9 13 3 10 0 9 3 3 13 2 16 10 3 9 9 3 0 9 13 0 2 7 0 2 7 10 9 9 15 13 2 15 3 13 3 2
16 3 0 10 0 10 9 10 9 2 7 1 10 0 3 13 2
68 1 3 10 13 9 3 15 3 15 13 3 15 13 3 13 2 7 3 16 9 13 1 15 1 10 0 13 3 13 2 7 16 9 13 1 10 0 10 9 16 0 2 13 0 7 10 0 1 9 15 3 1 10 0 13 2 13 7 13 1 10 0 9 16 0 13 3 2
37 3 10 9 0 2 3 10 9 1 15 3 3 13 10 13 3 0 13 2 13 7 10 0 3 13 2 1 0 10 9 13 13 3 0 13 15 2
35 3 0 3 9 13 0 3 13 13 7 1 15 3 13 2 0 10 9 0 10 13 13 13 15 3 15 15 13 7 10 3 3 15 13 2
28 3 3 3 13 15 0 1 10 3 13 10 13 3 13 2 13 16 0 10 0 9 10 3 13 2 3 13 2
37 10 3 9 10 13 1 10 9 3 1 10 13 13 13 13 2 7 16 15 13 2 7 15 3 15 13 7 1 10 15 0 0 9 1 0 13 2
27 3 3 13 2 16 10 13 10 9 0 3 10 15 1 10 15 13 2 7 16 0 15 9 7 9 13 2
12 3 1 3 9 3 10 3 0 15 0 13 2
28 0 3 13 10 3 13 10 0 13 7 10 13 3 3 1 10 0 15 3 0 13 2 0 13 15 3 13 2
13 9 3 1 3 3 16 9 1 10 3 13 13 2
21 10 3 0 9 0 13 10 0 2 7 15 3 0 9 7 9 0 10 9 13 2
24 0 3 10 9 9 3 0 13 2 9 7 13 13 1 15 10 9 0 3 0 1 0 9 2
70 10 7 0 9 3 13 2 9 7 0 13 3 0 13 2 9 3 1 2 15 1 0 3 9 9 7 0 10 0 13 2 9 3 9 2 15 0 1 10 1 10 3 9 13 13 2 9 7 13 1 15 0 3 1 15 3 9 7 10 3 0 13 7 9 0 13 10 0 9 2
10 15 3 0 1 0 10 9 3 13 2
17 13 3 15 9 7 9 13 10 0 9 15 15 13 1 9 9 2
25 16 3 13 2 10 9 13 0 7 10 9 2 10 3 15 13 3 1 15 0 9 10 9 13 2
25 10 3 3 0 9 2 0 7 9 2 10 9 13 0 13 7 9 13 10 9 13 1 10 13 2
21 10 3 1 10 0 13 9 15 13 0 2 1 15 13 10 9 1 10 9 13 2
11 9 13 9 1 9 13 1 10 0 9 2
26 15 13 3 9 2 9 7 13 9 9 0 9 10 1 9 2 1 3 10 0 9 1 10 9 13 2
11 13 3 3 9 15 7 10 0 0 9 2
13 13 3 10 9 13 10 10 9 9 0 7 0 2
24 13 3 1 15 9 0 2 16 13 2 1 9 0 10 0 9 13 7 10 9 10 0 13 2
32 10 3 0 1 0 10 9 10 9 15 13 10 0 2 10 7 13 1 10 9 13 10 1 10 9 1 3 9 7 1 9 2
38 10 3 1 10 9 13 9 16 13 2 13 1 10 9 9 3 9 13 2 13 3 15 13 13 2 7 10 3 13 13 15 7 10 10 9 9 13 2
12 10 3 9 10 9 3 13 2 7 0 13 2
39 13 3 10 9 0 15 1 9 9 13 1 0 13 13 10 13 2 7 13 1 9 10 9 13 16 13 9 10 9 3 9 7 9 0 13 1 15 13 2
9 10 3 15 13 13 7 9 13 2
37 13 3 10 9 1 10 9 1 10 9 13 10 9 2 10 3 9 13 15 1 9 13 7 10 9 13 2 13 7 3 15 13 13 2 7 13 2
33 9 3 1 3 10 0 13 10 9 2 13 3 0 15 13 10 9 16 9 2 3 3 7 9 10 9 2 16 15 13 13 0 2
21 13 3 0 1 9 2 9 13 9 2 9 10 9 16 13 1 15 1 9 13 2
21 9 3 16 13 10 3 9 7 9 13 1 10 9 10 7 9 9 13 2 13 2
26 10 3 9 15 15 13 2 7 13 1 15 10 9 0 9 1 10 9 3 13 2 7 10 9 13 2
15 13 3 10 9 13 9 3 10 13 7 10 9 0 13 2
12 13 3 3 10 13 0 7 10 10 9 13 2
16 13 3 3 10 9 9 15 13 2 16 3 13 1 9 13 2
13 10 3 13 15 0 9 13 2 7 9 9 9 2
22 3 9 13 2 15 13 0 2 9 7 0 7 9 0 2 9 7 0 7 9 0 2
15 9 3 9 13 7 9 2 9 7 9 3 0 7 9 2
10 0 3 9 9 13 0 7 0 9 2
37 16 3 13 10 9 10 9 2 13 1 9 1 0 7 0 9 2 15 13 2 13 9 10 1 9 9 3 7 9 13 2 16 3 13 15 9 2
17 16 3 15 13 2 9 13 13 1 9 1 9 15 3 0 13 2
9 13 3 3 10 1 9 9 13 2
6 9 3 3 13 13 2
25 16 3 3 2 3 15 13 13 2 15 13 2 9 13 15 3 13 0 10 3 13 3 9 1 2
19 10 3 9 13 15 2 16 10 3 9 7 10 9 1 9 13 2 13 2
15 9 3 13 2 16 3 15 10 1 9 13 2 13 15 2
41 9 3 15 15 13 2 7 16 0 15 13 10 9 7 10 0 13 2 13 9 0 9 13 9 2 13 0 9 7 0 0 7 9 13 1 10 9 9 0 13 2
29 13 3 10 3 9 9 10 9 3 9 10 9 7 9 10 9 2 10 7 0 9 3 10 9 7 9 10 9 2
54 16 3 13 1 9 10 0 9 2 3 10 9 10 9 13 2 1 10 9 10 0 9 2 10 9 9 3 13 15 1 9 13 16 13 1 15 7 10 9 3 13 2 13 3 10 0 16 0 13 7 10 15 13 2
15 3 13 10 9 1 0 7 9 0 7 0 13 10 9 2
29 10 3 0 9 15 13 3 10 10 9 13 13 9 16 10 3 9 13 2 9 7 13 13 16 3 0 15 13 2
27 1 3 10 9 10 9 0 13 1 10 9 10 9 9 10 3 0 15 13 0 13 2 9 7 13 13 2
52 0 3 2 16 10 9 7 10 0 13 10 9 13 1 9 2 10 9 0 13 10 1 0 10 9 10 9 2 3 13 1 9 10 9 9 10 9 13 7 9 10 9 9 13 2 16 9 7 9 13 9 2
59 10 3 9 10 0 1 10 9 13 10 9 7 10 10 9 0 13 13 2 1 15 9 13 10 9 13 9 7 9 2 16 15 10 0 13 2 13 1 9 7 1 10 9 10 9 9 1 10 3 9 7 10 0 9 0 15 0 13 2
13 13 3 3 10 9 1 10 9 9 3 7 0 2
17 13 3 0 15 2 7 10 9 0 13 9 3 13 1 9 0 2
32 10 3 9 13 15 13 7 0 1 10 9 13 2 16 3 15 1 10 9 0 3 10 15 13 0 13 13 10 9 15 13 2
14 13 3 9 1 9 13 2 7 10 3 9 13 15 2
16 9 3 1 10 9 10 9 3 15 13 0 15 13 13 15 2
23 13 3 10 0 9 1 3 15 1 10 9 15 0 7 1 10 0 15 1 10 13 0 2
11 10 3 3 13 9 15 1 0 13 9 2
9 0 3 13 1 10 1 15 0 2
3 3 13 2
52 0 9 0 7 15 10 0 0 2 16 0 15 3 1 0 9 7 9 13 9 15 13 2 15 13 0 1 9 7 9 13 15 2 3 3 13 1 3 10 0 9 2 15 3 13 9 2 15 7 0 9 2
27 15 1 10 0 9 0 3 3 0 13 2 7 0 9 13 15 13 9 7 9 3 0 13 16 13 13 2
27 16 3 13 16 3 0 10 0 0 15 13 2 13 16 0 9 3 3 13 13 10 9 2 13 7 13 2
15 3 3 1 10 0 2 7 1 10 0 10 13 13 13 2
6 16 3 13 0 13 2
16 13 3 1 9 1 9 9 3 16 10 0 13 10 9 13 2
15 10 3 0 10 9 1 10 13 10 0 13 0 3 13 2
12 13 3 3 10 9 9 13 15 0 13 0 2
19 13 3 1 15 2 10 9 9 15 0 13 2 13 1 0 3 13 13 2
52 3 0 16 15 3 1 3 10 0 13 13 10 9 3 3 3 1 10 0 9 7 3 0 1 10 0 0 2 15 7 1 10 13 3 9 13 7 1 10 3 3 9 2 7 1 9 13 13 15 15 13 2
11 0 3 1 0 9 15 3 13 15 13 2
31 15 3 3 13 7 3 0 13 13 2 15 7 3 3 9 0 13 7 13 13 2 7 3 1 10 0 9 9 13 13 2
37 0 3 2 16 1 9 13 2 10 13 13 2 7 0 16 10 3 15 0 15 13 2 15 0 9 2 7 15 3 0 2 7 0 10 13 13 2
90 3 15 15 13 3 13 13 2 13 7 16 1 15 13 10 9 13 2 13 10 3 13 15 9 13 10 0 3 13 2 10 7 13 3 13 0 13 1 13 10 0 0 13 2 7 3 3 1 10 9 3 10 0 16 3 10 9 13 2 7 3 10 0 15 13 2 16 1 10 13 7 0 3 13 9 10 3 13 13 9 13 15 1 0 9 13 3 7 13 2
32 10 3 3 9 7 9 3 9 13 2 16 3 3 0 13 9 13 10 7 3 1 10 3 13 2 7 1 10 15 0 13 2
19 0 3 3 0 2 10 7 0 3 1 0 2 15 3 3 13 15 13 2
33 15 3 16 13 10 0 1 0 13 7 9 15 13 2 9 3 7 9 3 13 2 13 7 15 13 1 15 0 9 10 0 13 2
6 15 3 10 9 13 2
55 0 9 0 3 0 1 10 13 15 10 9 13 2 7 16 3 15 3 13 7 15 3 3 13 2 13 0 3 15 1 0 3 3 1 10 0 9 13 2 16 10 1 15 3 9 0 13 7 10 15 9 3 3 13 2
10 13 3 9 1 10 0 15 3 13 2
23 10 3 1 9 7 3 9 13 2 0 3 0 13 1 10 9 7 9 13 7 13 13 2
34 3 10 9 15 3 0 9 13 13 15 9 15 13 15 3 16 1 9 13 2 1 10 0 1 10 3 13 3 10 15 9 13 13 2
40 3 0 10 0 0 3 16 3 13 0 13 2 7 16 1 0 13 7 16 1 15 3 3 13 13 2 3 3 16 13 0 13 2 16 7 3 15 13 13 2
30 3 16 13 9 2 16 13 2 0 2 0 0 13 10 3 2 0 3 0 13 15 10 9 13 7 13 10 0 13 2
31 3 3 1 10 15 7 1 15 15 13 2 0 7 13 13 3 1 0 7 3 13 2 13 16 3 1 10 3 13 13 2
23 15 3 3 15 13 1 10 1 15 13 13 2 7 1 10 9 3 13 7 10 13 13 2
13 10 3 0 9 13 15 2 7 3 1 0 13 2
26 3 0 16 2 16 10 0 13 13 2 15 3 0 3 3 13 2 7 13 3 3 3 3 15 13 2
23 0 3 13 2 16 3 13 2 15 3 13 10 0 9 2 15 7 0 13 10 15 9 2
29 9 3 7 9 9 0 1 15 15 3 13 7 9 0 13 13 3 3 13 2 13 7 15 1 9 13 9 13 2
38 3 13 3 9 0 13 13 2 15 3 3 10 13 7 1 10 0 13 13 15 13 13 2 7 10 1 0 10 3 9 3 7 10 9 3 13 13 2
23 15 3 3 16 13 10 9 2 7 16 13 15 3 13 2 3 3 10 0 10 9 13 2
27 3 3 13 3 10 3 0 15 13 2 7 3 15 3 13 3 13 2 7 13 7 0 13 15 13 15 2
60 15 13 2 16 0 13 2 3 13 2 7 3 1 15 15 3 13 2 15 7 13 2 7 1 15 15 10 3 9 15 3 3 13 10 9 3 13 7 10 9 13 10 1 15 9 10 0 13 2 3 7 13 10 9 0 3 10 13 13 2
17 16 3 3 15 3 1 13 9 13 7 15 0 7 9 13 13 2
10 16 3 3 3 3 15 13 13 13 2
48 16 3 13 1 10 9 13 1 0 15 13 10 0 9 13 2 3 10 1 9 0 13 10 9 13 2 7 15 3 15 15 13 9 13 7 15 3 10 13 2 16 13 2 9 1 9 13 2
9 15 3 15 3 13 15 13 3 2
15 3 3 15 0 9 3 13 2 7 3 15 1 0 0 2
15 9 3 2 16 13 1 15 2 3 13 3 1 15 15 2
31 16 3 10 0 15 13 13 13 2 13 3 15 10 0 3 0 15 13 2 7 10 9 1 15 0 3 16 1 15 13 2
40 9 3 3 0 1 15 13 0 1 10 9 9 2 9 7 7 9 9 0 2 15 3 0 13 16 13 7 3 0 16 13 2 13 15 1 10 13 13 13 2
18 9 3 0 13 3 1 10 9 1 10 0 9 1 9 0 9 13 2
35 0 3 3 13 10 13 2 16 3 0 0 13 2 0 7 10 13 2 16 3 13 0 13 2 16 3 10 0 0 13 9 1 10 3 2
19 10 3 3 13 10 0 0 9 16 10 3 0 13 1 9 10 0 13 2
23 10 3 0 13 2 13 15 0 13 10 9 1 15 10 3 13 0 3 7 10 13 0 2
13 3 9 0 3 0 13 9 15 7 13 15 13 2
14 3 15 13 10 13 3 13 7 10 0 13 15 0 2
7 15 3 3 10 9 13 2
49 13 3 10 1 9 9 3 3 13 15 2 7 10 9 13 3 13 10 9 9 13 0 2 13 7 16 3 15 15 2 16 0 13 2 16 15 13 2 9 3 7 10 15 9 13 1 9 13 2
16 3 3 10 3 9 7 9 3 13 15 10 9 1 9 13 2
22 0 3 9 10 9 10 9 13 2 7 10 9 13 3 0 0 0 9 15 13 0 2
16 13 3 15 9 3 10 9 3 9 10 9 7 9 10 9 2
10 13 3 15 10 3 13 1 10 9 2
18 9 3 0 13 3 3 1 9 0 2 9 7 9 10 9 0 0 2
18 16 3 13 10 1 9 9 1 9 13 2 13 1 9 10 9 9 2
18 13 3 9 2 7 9 1 15 13 1 9 1 10 9 10 9 9 2
9 13 3 1 15 9 9 1 9 2
18 1 3 10 9 9 9 13 13 1 15 2 1 15 3 10 9 13 2
20 13 3 3 9 9 2 13 10 9 7 9 2 15 1 10 9 13 10 9 2
13 10 3 3 9 10 9 3 13 3 7 9 13 2
31 10 3 9 16 13 15 13 2 13 0 7 0 9 2 15 13 9 3 9 7 9 2 13 1 0 10 9 15 13 9 2
6 3 10 0 0 13 2
16 1 3 10 9 15 10 9 10 0 13 7 9 0 9 13 2
13 13 3 3 10 9 1 10 9 0 10 9 13 2
10 10 3 3 9 3 3 15 0 13 2
35 16 3 13 10 9 2 13 0 9 9 13 16 1 9 1 10 9 9 2 7 3 9 13 13 10 10 9 9 0 3 7 1 15 13 2
21 0 3 9 0 10 9 10 0 10 9 13 1 10 9 7 10 0 10 9 13 2
34 13 3 2 16 10 9 0 13 2 13 2 0 3 9 13 0 1 10 9 2 0 7 9 3 7 9 2 10 0 9 0 3 13 2
19 13 3 10 9 0 2 10 3 9 3 3 2 9 7 10 0 0 13 2
37 16 3 13 15 2 3 3 13 1 3 10 9 7 9 10 9 2 3 3 15 13 10 1 10 9 9 1 10 9 2 15 13 13 13 10 9 2
15 9 3 3 13 2 7 9 7 9 10 0 13 16 9 2
42 3 3 3 0 9 7 0 13 10 9 2 1 15 10 0 9 13 10 9 2 16 3 13 2 9 3 13 10 0 2 9 7 3 13 13 10 9 10 9 10 9 2
9 3 3 10 0 9 10 9 13 2
17 3 3 3 10 9 7 10 0 13 2 3 2 7 10 9 13 2
21 10 3 9 13 10 9 13 3 3 3 13 2 10 3 0 13 16 3 13 15 2
35 16 3 10 9 13 3 7 13 10 9 2 3 3 9 0 13 3 7 13 15 3 2 7 13 1 15 9 16 13 15 10 9 7 9 2
46 10 3 9 13 10 9 10 9 3 3 13 13 10 9 15 13 2 1 7 10 9 13 13 13 3 16 13 2 10 7 15 9 2 3 13 16 13 10 1 10 0 9 2 13 13 2
15 9 3 0 9 1 9 9 9 0 3 10 1 15 13 2
41 16 3 13 10 9 10 9 1 10 9 2 1 10 9 7 10 9 10 0 13 2 7 10 0 13 16 13 1 10 9 2 3 15 10 1 9 9 10 9 13 2
9 13 3 10 9 10 9 9 0 2
9 15 7 13 3 13 13 10 9 2
25 10 3 10 0 3 0 13 0 1 10 0 9 7 15 13 2 13 16 1 10 9 15 13 13 2
17 15 3 13 10 9 7 13 1 9 13 3 0 13 7 0 13 2
6 3 3 3 15 13 2
12 13 3 3 2 7 10 9 13 10 9 13 2
14 3 3 10 9 13 15 2 7 10 9 13 1 9 2
45 10 3 9 13 1 10 9 10 0 9 10 1 10 9 0 2 15 13 9 3 10 9 7 2 9 10 9 2 2 1 10 9 7 9 13 13 1 10 9 3 0 0 16 13 2
3 3 13 2
34 10 3 0 13 10 3 0 0 9 7 10 9 0 0 13 13 1 10 1 10 9 9 2 1 15 10 9 13 2 13 13 16 13 2
28 10 3 3 9 3 13 3 13 2 13 16 10 9 13 13 10 9 2 16 1 9 13 2 3 13 15 13 2
16 13 3 15 9 1 9 13 1 9 13 10 9 7 13 13 2
5 13 3 13 15 2
11 15 3 0 10 0 13 3 13 9 13 2
29 16 3 15 9 13 13 3 15 1 9 7 3 16 3 13 13 7 10 9 13 2 15 0 0 13 13 16 0 2
6 10 3 3 15 13 2
22 10 3 9 10 3 9 0 13 13 3 13 3 15 7 13 2 10 7 9 15 13 2
11 16 3 3 3 3 13 13 2 3 13 2
18 16 3 1 9 13 7 1 10 15 15 9 2 3 13 1 10 0 2
24 15 10 9 13 10 3 9 10 3 9 10 1 9 13 7 9 13 1 10 1 10 9 9 2
40 10 3 9 10 3 9 7 9 13 10 1 15 13 1 3 10 9 7 9 2 15 13 10 9 13 15 3 2 7 9 13 1 10 1 10 9 9 3 13 2
8 9 3 0 0 10 9 13 2
31 9 3 13 10 9 1 9 2 16 3 9 0 7 9 13 2 3 9 13 0 3 0 0 9 7 13 1 0 13 9 2
6 3 3 0 13 13 2
12 13 3 3 9 15 10 0 0 13 10 9 2
17 1 15 3 3 3 0 13 13 10 9 7 9 9 1 10 13 2
15 15 3 1 10 9 10 9 13 3 1 10 1 9 9 2
22 10 3 3 9 3 3 0 13 2 9 7 10 9 9 9 13 0 0 7 0 13 2
18 13 3 16 9 10 15 9 7 9 3 1 15 13 10 9 9 13 2
24 13 3 13 1 7 10 9 13 16 9 13 15 1 9 2 7 10 9 13 10 9 1 9 2
31 13 3 9 3 10 1 9 9 7 9 13 2 13 2 16 0 15 13 0 13 10 9 2 0 3 10 9 1 15 13 2
21 3 9 13 9 10 1 9 9 13 7 13 13 1 9 0 7 9 0 0 13 2
24 10 3 13 15 10 15 9 10 9 1 10 9 9 13 13 2 16 3 10 1 9 9 13 2
13 3 10 3 13 3 13 10 9 7 1 9 13 2
22 10 3 0 9 10 9 13 1 10 1 9 2 7 13 10 3 9 7 10 15 13 2
42 13 3 10 9 0 13 1 3 9 13 10 13 9 7 10 13 9 13 1 10 9 2 1 15 3 10 0 13 2 7 13 13 1 9 7 10 9 9 3 9 13 2
21 13 3 15 9 10 9 2 1 9 7 15 3 0 10 0 1 9 9 9 13 2
8 13 3 10 9 3 3 0 2
11 3 13 0 9 9 1 9 16 9 13 2
79 13 3 3 15 10 9 13 3 2 3 7 9 13 7 9 0 1 10 9 2 16 15 13 10 9 7 10 9 13 2 13 1 10 9 2 7 13 1 9 3 3 1 9 3 13 0 10 9 7 3 13 13 1 9 1 10 9 2 0 3 9 15 2 3 3 10 0 0 2 9 7 0 9 10 1 9 7 9 2
6 3 3 9 13 0 2
11 1 0 3 13 0 13 1 9 7 13 2
17 13 3 3 3 10 9 7 13 10 9 2 9 1 15 13 13 2
38 9 3 6 10 10 9 9 7 10 13 10 3 9 9 7 10 9 0 1 9 13 2 16 13 10 3 13 2 15 7 13 10 9 13 1 10 9 2
25 3 16 1 10 9 13 7 13 10 0 13 3 1 9 2 13 3 15 2 7 3 0 0 13 2
28 3 0 3 10 10 9 9 7 0 1 15 13 9 3 7 10 0 9 13 10 1 15 7 13 13 1 0 2
17 10 3 0 9 9 7 9 13 1 10 9 7 1 10 9 13 2
40 13 3 3 13 10 1 15 3 1 0 9 9 13 1 10 9 2 7 13 1 10 9 1 10 9 13 3 7 3 2 0 3 15 13 2 10 7 0 13 2
26 16 3 1 9 10 9 10 9 13 7 10 9 13 2 3 13 1 10 9 7 10 9 1 10 9 2
5 9 3 0 13 2
16 1 3 10 9 0 13 10 9 7 10 9 0 13 10 9 2
22 13 3 9 3 7 10 9 0 0 0 2 9 7 0 0 7 0 7 9 10 9 2
8 10 3 1 10 9 0 13 2
29 3 3 0 13 13 1 3 10 9 13 7 1 10 9 13 13 2 13 16 15 10 9 7 10 9 13 3 13 2
26 3 13 10 1 10 9 9 10 9 0 13 2 9 0 13 0 7 0 9 15 7 9 10 9 9 2
16 3 3 3 1 9 10 9 3 13 7 1 9 9 3 13 2
45 9 3 13 15 7 9 0 13 9 2 16 3 15 1 9 7 15 1 9 13 2 13 3 1 0 9 13 10 15 13 2 16 1 0 10 9 13 2 7 15 13 10 13 13 2
26 16 3 3 13 2 13 10 1 15 13 7 16 10 3 13 3 0 2 9 13 13 10 9 10 9 2
27 3 13 1 9 10 3 15 13 7 9 13 1 10 9 0 13 2 1 7 10 9 13 3 9 0 13 2
25 1 3 10 9 10 9 9 3 13 10 0 7 0 10 9 7 9 13 7 13 15 3 9 13 2
13 3 3 10 3 9 3 13 2 7 3 9 13 2
7 0 3 15 10 9 13 2
18 13 3 10 9 3 13 2 9 3 15 13 7 3 1 10 9 13 2
23 13 3 3 1 10 9 10 9 7 13 13 10 9 16 9 3 13 13 7 13 10 9 2
29 9 3 3 3 3 13 2 13 10 9 2 3 7 3 0 1 15 13 10 9 2 13 3 13 0 1 10 9 2
26 10 3 9 13 10 9 3 7 16 15 15 0 13 13 1 9 2 9 15 0 13 10 13 13 13 2
37 3 15 3 13 9 13 3 0 7 9 2 13 3 3 0 3 0 9 2 3 7 9 3 13 10 1 10 9 9 7 10 9 9 1 10 9 2
15 13 3 0 9 7 10 15 13 0 13 10 9 13 15 2
16 3 1 15 9 3 13 2 9 7 0 1 10 1 9 13 2
32 3 3 13 15 15 13 1 9 13 2 3 1 15 13 3 10 9 13 2 7 10 13 3 13 16 1 10 15 0 0 13 2
42 3 1 15 3 16 13 2 7 16 1 10 9 13 2 10 9 0 13 2 1 15 13 15 3 0 13 2 0 3 0 9 13 1 3 9 13 2 1 7 15 13 2
17 3 16 3 0 3 13 13 10 9 2 9 3 3 3 13 13 2
32 3 3 3 9 3 13 9 15 13 7 9 13 2 15 10 3 0 9 1 10 1 9 13 2 10 7 0 3 0 13 9 2
43 3 15 15 0 2 10 3 0 13 15 10 9 1 10 0 13 7 0 10 0 13 9 2 1 15 7 3 13 3 0 10 1 15 13 9 2 7 3 10 0 3 9 2
28 3 3 10 13 2 7 10 13 3 13 13 7 0 15 13 2 16 3 10 9 10 9 3 13 10 9 13 2
11 3 3 3 3 13 3 7 3 1 0 2
13 13 3 3 16 13 3 13 2 7 1 15 13 2
13 10 3 13 13 1 3 13 3 7 3 13 13 2
15 3 13 0 9 10 9 7 15 1 0 13 1 10 3 2
18 3 13 3 13 1 10 0 15 0 13 2 13 7 13 13 3 13 2
13 3 15 15 1 9 10 0 7 9 13 15 13 2
13 9 3 3 0 9 13 13 2 9 7 0 13 2
51 3 3 2 16 15 3 0 2 0 13 13 10 3 9 13 2 3 3 3 0 10 13 13 2 1 15 3 13 15 3 13 2 7 13 3 1 0 15 9 13 7 0 15 7 3 0 13 10 9 13 2
14 10 3 3 0 7 13 0 7 13 9 15 3 13 2
18 3 3 10 3 3 1 9 9 3 1 9 9 7 1 10 0 9 2
22 10 3 0 10 3 9 0 13 10 3 9 3 10 0 13 10 7 0 3 13 13 2
12 3 3 3 0 1 0 9 7 9 1 0 2
20 13 3 10 3 10 9 3 15 13 2 15 7 10 13 3 10 0 3 13 2
13 13 3 10 0 1 0 13 7 13 1 0 13 2
22 3 3 10 3 9 0 1 10 9 13 2 10 7 9 0 1 10 13 15 1 15 2
25 3 15 3 3 13 3 13 2 0 13 13 2 15 7 3 13 13 2 0 1 10 13 13 13 2
14 16 3 3 15 3 9 13 2 13 15 13 10 9 2
20 0 3 13 3 3 7 13 15 3 13 1 10 0 10 9 13 15 3 13 2
23 3 16 15 15 13 13 13 1 10 3 15 13 9 7 10 0 9 13 2 3 3 13 2
9 3 3 3 9 0 13 13 15 2
16 3 3 2 15 3 3 13 2 0 15 10 9 1 15 13 2
20 3 13 3 9 10 0 0 0 2 1 0 7 13 13 0 3 10 9 13 2
14 1 15 3 10 10 9 1 10 9 1 0 15 13 2
9 1 3 3 15 13 15 10 9 2
40 3 3 10 3 15 7 9 2 16 13 2 13 1 9 13 1 10 9 2 16 3 9 3 0 7 0 10 0 13 7 15 10 0 9 1 0 0 9 13 2
16 13 3 3 0 15 3 1 9 10 9 7 1 9 10 13 2
18 13 3 9 3 10 1 9 15 13 2 7 10 3 13 15 3 13 2
7 13 3 15 0 13 13 2
12 3 3 0 3 13 13 7 0 3 15 13 2
17 1 15 13 3 7 10 9 13 3 0 13 16 10 9 15 13 2
6 15 3 10 9 13 2
56 10 3 9 13 3 9 0 1 10 9 1 15 13 2 7 16 13 10 9 2 13 15 0 1 10 9 13 2 10 3 9 1 15 13 15 10 9 13 2 13 7 1 10 0 16 3 3 15 0 13 2 7 1 0 0 2
19 13 3 10 9 13 13 3 15 1 10 9 15 13 2 16 15 3 13 2
13 10 3 13 3 13 2 7 13 10 9 13 15 2
19 10 3 9 15 3 1 9 10 0 9 13 2 7 1 15 10 9 13 2
28 3 3 16 13 2 1 9 13 2 15 10 3 9 9 13 2 10 7 9 3 0 2 16 15 13 2 13 2
21 13 3 3 9 3 1 16 9 7 9 1 0 15 9 3 3 13 10 9 13 2
50 13 3 9 3 0 13 10 9 7 16 10 0 13 2 3 0 13 1 9 13 2 13 1 10 9 3 1 9 13 2 15 13 3 1 9 15 13 10 9 13 2 0 3 13 1 9 0 15 13 2
6 9 3 0 15 13 2
19 13 3 10 9 3 3 15 0 13 10 9 1 9 10 0 10 9 13 2
45 9 3 3 1 10 0 0 0 10 0 9 2 9 7 13 2 15 0 1 10 0 13 13 2 15 0 13 10 9 2 3 0 1 15 15 13 3 3 9 0 10 1 15 13 2
59 9 3 3 0 0 13 2 10 3 2 16 15 1 9 15 13 2 10 15 3 1 15 13 13 13 10 9 7 10 0 13 3 3 10 10 0 9 0 13 7 13 0 15 13 2 7 13 1 10 9 13 7 3 13 16 15 3 13 2
11 3 13 3 0 15 13 15 16 13 15 2
26 15 3 1 3 10 3 13 3 13 7 1 10 1 0 9 13 13 13 15 3 10 9 7 15 0 2
49 16 3 13 0 10 9 13 2 16 3 15 2 1 10 9 2 7 3 13 0 13 1 10 9 3 13 2 15 3 13 3 15 3 13 9 0 13 2 7 1 9 3 15 13 10 9 3 13 2
31 3 3 0 15 13 3 13 2 7 15 3 3 13 13 1 10 0 10 9 2 15 7 13 10 9 7 15 13 9 13 2
26 1 0 3 10 9 13 10 0 13 15 1 15 2 3 3 1 9 2 3 3 9 2 0 7 9 2
33 3 3 0 3 13 13 10 0 13 2 7 15 3 3 13 13 2 15 7 15 3 3 0 2 7 0 7 0 13 2 13 13 2
9 3 3 3 10 9 1 15 13 2
12 0 3 0 10 13 10 0 1 9 3 13 2
34 3 16 3 13 1 0 13 1 10 9 2 16 15 2 3 13 3 3 0 15 0 13 10 9 7 13 3 3 13 3 7 15 13 2
19 13 3 0 15 13 10 0 9 16 0 13 0 16 1 10 13 9 13 2
15 15 3 3 3 13 10 0 13 13 3 3 16 15 13 2
15 15 3 3 1 10 0 9 10 0 16 9 3 3 13 2
24 3 13 3 1 10 0 1 10 9 9 7 1 15 0 1 10 0 9 13 10 9 13 13 2
23 3 15 13 15 10 3 3 3 9 13 7 0 15 1 10 0 0 13 16 15 3 13 2
10 13 3 15 3 13 2 13 15 13 2
52 10 3 13 1 15 1 10 0 13 2 16 15 1 10 3 13 13 3 9 7 9 10 1 10 9 7 3 13 2 3 10 0 3 13 9 13 2 7 10 0 0 13 16 16 1 0 13 10 9 3 13 2
13 13 3 2 16 13 2 10 9 3 13 16 13 2
16 10 3 3 1 10 0 13 13 2 10 7 1 10 0 13 2
8 10 13 3 3 0 10 0 2
38 15 3 3 3 16 13 15 13 2 3 3 10 9 15 1 10 0 9 13 13 2 16 0 3 3 1 10 9 1 0 13 13 2 0 3 3 13 2
26 0 3 10 3 1 15 0 0 10 15 13 7 3 9 0 13 3 15 13 7 15 10 0 9 13 2
19 13 3 3 16 3 1 0 2 7 3 0 9 7 9 13 0 9 13 2
20 13 3 13 1 9 10 0 13 2 15 0 3 13 7 3 13 1 0 13 2
24 13 3 10 9 1 10 9 10 9 0 13 2 15 13 0 13 2 13 7 3 10 9 13 2
40 15 3 1 0 3 0 9 13 3 0 7 15 13 13 15 2 16 3 0 0 10 9 2 9 3 13 7 13 10 9 2 10 7 9 9 13 1 10 9 2
18 16 3 3 2 9 10 0 9 13 13 13 9 13 3 3 3 13 2
6 15 3 10 9 13 2
30 16 3 10 3 9 13 10 9 10 9 10 1 10 9 7 10 9 15 13 2 13 0 13 1 15 0 1 10 13 2
19 13 3 3 15 1 15 3 13 3 3 0 13 2 16 3 15 15 13 2
21 1 3 3 9 7 10 0 0 15 10 9 2 7 1 0 0 3 1 0 13 2
4 3 0 13 2
18 3 0 0 3 15 13 3 3 1 0 13 7 3 1 10 0 13 2
19 3 3 15 13 16 10 9 15 7 10 9 13 2 16 10 9 13 13 2
16 10 3 0 9 13 0 15 13 2 7 1 9 15 13 13 2
18 16 3 3 10 9 13 13 2 13 3 15 9 13 10 0 13 9 2
7 0 3 13 15 10 9 2
20 16 3 3 3 9 13 7 10 9 13 1 15 10 0 13 2 13 10 0 2
20 3 3 3 0 3 10 9 13 16 0 13 10 9 2 16 10 9 15 13 2
10 13 3 3 16 3 10 9 15 13 2
15 3 13 9 9 3 10 9 13 7 3 0 13 10 9 2
20 16 3 3 2 13 9 0 7 0 0 3 2 16 13 2 13 13 1 15 2
32 3 3 13 15 3 10 3 9 7 10 9 15 0 13 3 3 13 2 3 9 3 0 13 7 1 13 0 7 3 13 13 2
18 3 3 0 15 13 10 9 15 16 9 13 3 3 0 0 0 13 2
16 15 13 13 3 1 0 2 7 3 1 9 13 15 0 13 2
21 16 3 0 10 10 9 9 13 13 15 2 13 16 3 0 7 0 10 9 13 2
11 9 3 3 3 9 7 9 0 3 13 2
21 9 3 0 13 1 10 0 2 15 3 13 13 1 15 13 2 3 0 3 13 2
12 3 9 0 0 0 9 3 0 13 13 13 2
34 13 3 3 15 3 0 9 13 9 2 7 13 10 9 3 9 10 0 7 9 2 1 15 10 9 13 2 3 3 7 9 1 0 2
35 13 3 0 15 2 3 3 10 10 9 9 0 13 2 15 3 3 10 13 10 0 1 0 10 9 13 2 15 7 1 9 15 15 13 2
14 3 10 0 7 13 2 15 13 3 15 2 3 13 2
21 13 3 3 0 3 13 1 10 0 13 2 7 3 0 7 0 9 1 0 13 2
8 3 13 3 9 0 15 13 2
14 0 3 1 15 9 3 3 13 7 9 0 0 13 2
31 10 3 1 9 13 15 1 10 0 1 10 13 15 3 13 9 2 7 16 15 3 1 9 13 2 15 3 3 13 13 2
11 3 3 3 1 3 13 10 0 9 13 2
18 3 3 1 15 3 13 13 13 10 9 2 7 3 15 0 3 13 2
18 0 3 13 3 13 13 9 9 2 0 7 13 15 1 10 0 13 2
39 0 3 15 10 9 3 15 13 9 7 15 1 0 13 13 3 13 2 7 13 1 0 9 9 1 0 9 3 9 3 9 7 9 13 2 7 1 9 2
8 13 3 15 3 0 1 9 2
12 1 3 10 13 3 0 0 16 1 13 13 2
10 15 3 3 0 13 7 10 0 0 2
7 3 10 3 9 15 13 2
18 13 3 9 0 2 9 10 9 3 13 2 13 2 10 9 2 3 2
10 10 3 9 10 0 10 9 3 13 2
16 13 3 0 15 3 13 16 3 13 10 0 9 7 10 9 2
26 3 16 1 10 9 13 0 3 2 1 7 15 0 3 2 0 9 0 13 2 16 1 0 0 13 2
23 15 3 0 3 3 7 3 13 2 7 10 9 2 16 13 2 3 13 13 7 13 13 2
7 10 3 3 13 3 13 2
42 15 3 3 9 13 0 3 9 7 9 2 15 7 9 0 2 15 3 0 10 9 13 2 7 9 7 9 0 3 9 3 15 13 2 7 0 1 0 3 0 9 2
19 3 16 15 13 13 13 15 13 2 7 10 13 13 3 13 0 9 13 2
12 15 13 13 15 9 13 1 10 9 10 9 2
14 13 3 13 2 7 0 0 13 15 13 10 9 13 2
33 13 3 10 9 13 16 15 3 13 13 10 9 2 13 7 3 10 0 9 13 9 13 2 16 3 13 10 9 13 2 16 13 2
19 3 10 3 13 1 9 13 15 2 7 10 9 9 9 1 15 13 13 2
30 10 3 9 0 10 9 2 10 10 9 13 2 13 1 10 0 7 0 9 10 9 9 13 2 15 13 1 10 0 2
36 13 3 10 9 10 9 13 7 0 13 3 15 10 9 13 10 9 0 13 10 9 16 1 0 13 2 13 15 10 0 10 9 0 3 13 2
13 10 3 9 9 0 13 1 10 9 1 15 13 2
35 9 3 10 0 2 16 15 10 9 1 10 9 13 2 13 3 3 13 9 3 9 7 10 13 9 2 7 10 9 13 13 7 10 9 2
26 10 3 3 0 0 13 7 9 10 3 0 13 2 0 7 13 2 1 15 0 13 10 0 10 9 2
52 9 3 13 10 13 13 9 2 10 3 3 15 0 3 13 3 15 7 0 15 9 13 2 10 7 0 10 9 13 7 13 10 3 0 15 10 9 2 15 3 3 13 2 7 10 1 10 0 9 9 13 2
57 13 3 15 3 13 2 7 3 10 1 9 3 0 13 13 1 15 10 0 2 10 3 13 7 0 10 9 3 13 1 10 9 2 3 7 10 9 2 16 3 13 2 3 3 13 1 0 3 2 16 3 1 10 9 2 13 2
12 10 3 9 0 13 9 3 7 9 0 13 2
22 10 3 9 9 9 10 3 9 15 13 13 16 13 1 15 9 1 15 13 3 13 2
39 15 3 13 13 3 0 10 9 1 10 9 2 0 7 1 15 13 9 3 3 13 2 7 13 1 15 16 3 10 9 0 13 16 13 1 10 0 9 2
16 3 10 3 15 13 7 13 10 15 16 15 10 3 13 13 2
16 3 1 10 9 13 3 13 1 10 9 2 7 13 7 13 2
39 3 16 15 15 13 10 1 9 13 16 3 13 1 10 0 2 13 10 9 13 2 9 7 0 13 15 13 2 13 7 1 0 13 7 13 16 3 13 2
32 10 3 13 10 3 9 13 1 9 15 2 10 7 15 13 7 3 13 16 13 3 7 3 9 13 2 3 13 16 13 13 2
21 13 3 15 13 15 3 9 3 13 16 13 15 0 9 15 0 7 3 13 13 2
63 10 3 3 9 10 9 2 16 13 2 13 2 7 10 9 13 10 9 3 3 3 13 16 10 3 9 15 13 3 16 0 13 13 10 13 2 16 7 15 13 9 7 10 9 13 1 15 2 3 1 13 10 0 13 10 3 15 0 0 7 10 0 2
33 10 3 3 9 16 13 13 0 13 7 1 10 9 13 2 1 15 13 13 13 2 7 0 3 1 15 13 2 15 0 9 13 2
14 3 0 3 0 13 13 13 7 3 15 13 3 13 2
9 10 3 9 0 13 1 9 3 2
12 0 10 9 10 9 10 9 13 1 0 9 2
13 3 0 10 9 3 3 3 13 16 1 9 13 2
28 10 3 0 0 9 13 7 3 13 13 3 2 7 16 0 3 13 2 0 3 9 1 9 7 9 13 13 2
17 0 3 10 0 3 13 10 9 2 7 1 15 0 3 13 13 2
18 3 13 10 15 9 10 9 10 9 15 3 3 0 13 1 10 9 2
9 0 3 9 0 15 10 9 13 2
25 3 3 3 9 7 9 13 2 7 13 0 9 7 9 0 2 9 1 15 10 3 7 9 13 2
9 10 3 9 0 3 13 15 13 2
32 13 3 10 9 7 10 9 13 10 10 0 9 2 9 7 13 0 3 15 0 13 10 9 2 10 7 15 1 10 9 13 2
25 10 3 9 3 13 2 13 2 16 15 13 2 10 9 9 10 1 9 9 0 10 1 9 13 2
31 10 3 9 0 13 10 3 9 2 7 3 10 9 13 2 16 3 3 1 9 13 2 13 1 15 10 9 1 0 13 2
15 9 3 3 3 13 7 10 15 13 3 1 10 9 9 2
16 9 3 10 9 1 9 9 10 9 13 1 0 9 1 9 2
12 13 3 3 9 0 9 7 10 0 9 9 2
24 3 13 1 9 7 15 10 0 13 2 7 0 1 9 9 13 2 7 13 1 0 10 9 2
22 3 3 0 13 15 10 3 0 9 13 3 3 0 10 9 7 0 1 9 3 13 2
22 13 3 1 10 9 13 15 9 15 13 1 10 0 7 9 3 13 2 16 3 13 2
23 10 3 9 13 3 10 9 7 13 10 9 3 3 13 10 15 7 13 15 13 0 15 2
12 1 15 3 10 9 13 9 13 15 1 13 2
20 3 3 9 0 13 15 1 10 9 10 13 2 7 9 3 13 9 3 9 2
21 13 3 15 13 7 3 3 10 9 10 15 9 1 9 13 1 10 1 9 9 2
19 13 3 1 9 10 3 0 1 15 9 13 2 10 7 0 13 3 13 2
11 13 3 15 3 0 9 7 13 0 13 2
19 3 15 3 3 13 9 2 9 7 7 0 15 1 15 9 13 3 0 2
8 15 3 13 10 9 10 9 2
32 13 3 10 9 10 9 0 10 9 0 10 9 1 10 9 9 2 13 15 3 13 13 10 9 9 1 10 9 7 15 9 2
11 9 3 13 13 15 13 13 10 9 9 2
13 3 9 3 0 9 13 9 2 15 13 10 9 2
8 3 3 13 10 9 10 9 2
11 13 3 10 0 9 13 0 9 7 0 2
14 9 3 9 13 15 2 7 10 9 1 10 9 13 2
48 13 3 0 10 0 10 9 7 1 0 9 13 15 13 9 3 7 9 9 1 0 10 9 7 10 0 2 15 13 1 3 10 9 15 7 1 10 0 9 13 7 9 10 3 13 1 0 2
20 15 3 15 3 13 1 10 0 9 9 2 3 3 7 10 9 3 3 13 2
15 3 3 3 10 9 9 13 10 10 9 1 0 9 13 2
18 0 3 9 10 1 9 9 13 9 13 7 13 2 9 10 9 13 2
17 3 9 10 1 10 0 9 2 15 13 9 2 13 7 13 15 2
17 1 3 9 15 1 10 0 9 9 13 2 7 9 13 1 9 2
29 9 7 13 1 15 13 7 9 13 2 0 7 0 9 9 1 10 13 13 2 3 7 3 10 0 16 0 13 2
21 9 3 0 3 13 10 9 7 0 10 10 9 7 9 9 7 9 16 15 13 2
17 10 3 9 3 13 7 0 13 3 13 7 13 13 13 10 9 2
27 13 3 3 7 3 10 9 3 3 1 9 13 2 7 3 13 1 10 0 0 7 13 13 15 10 13 2
7 15 0 0 13 10 9 2
55 1 3 10 9 0 10 9 10 0 15 2 16 3 1 9 13 2 9 13 1 10 9 10 13 9 13 2 7 10 3 9 13 10 0 1 10 9 15 15 13 2 15 7 2 16 13 2 0 7 0 1 10 9 13 2
44 13 3 1 15 3 10 1 9 9 1 9 9 7 9 9 7 10 9 1 9 2 7 13 10 0 9 0 9 9 10 9 13 2 7 13 9 9 7 13 10 0 1 0 2
22 9 3 0 13 9 15 13 2 13 1 10 1 10 3 9 9 7 10 9 15 13 2
13 0 3 10 9 13 10 10 0 9 3 13 0 2
7 15 3 9 13 10 0 2
9 10 3 13 9 13 9 3 0 2
7 9 3 3 13 10 9 2
13 3 9 1 0 10 9 0 9 7 9 0 13 2
16 3 9 3 3 0 1 15 10 0 9 13 0 1 9 13 2
14 13 3 3 9 7 9 10 13 7 9 10 3 13 2
19 3 10 9 13 1 10 9 10 3 10 9 13 13 7 10 15 13 13 2
10 10 3 9 13 15 10 9 1 9 2
15 1 3 10 9 3 0 15 13 9 13 9 7 9 13 2
12 13 3 15 1 9 13 13 0 9 0 13 2
17 13 3 1 15 10 9 3 3 9 0 7 10 0 9 3 0 2
7 0 3 13 0 7 0 2
18 3 9 3 1 10 9 13 7 13 3 13 1 9 1 9 7 9 2
11 3 3 10 10 9 9 13 0 9 13 2
14 9 3 3 1 9 13 1 9 10 1 10 9 9 2
15 10 3 1 10 0 9 9 7 10 9 1 9 3 13 2
15 3 13 9 7 9 13 9 10 9 13 10 9 1 9 2
12 0 3 13 9 0 9 13 9 7 9 0 2
12 3 3 0 9 13 15 13 7 13 13 9 2
9 3 9 13 7 13 13 9 13 2
13 3 10 13 9 13 7 10 15 0 0 3 13 2
11 13 3 9 3 9 7 9 13 10 9 2
13 10 3 9 3 1 9 13 10 9 1 10 9 2
6 15 3 13 9 9 2
14 13 3 3 1 0 10 9 9 9 13 13 10 9 2
6 13 3 15 3 9 2
15 13 3 3 1 10 9 0 9 9 7 15 1 10 9 2
8 13 3 9 3 10 9 13 2
10 13 3 3 9 16 3 0 0 13 2
30 15 3 0 0 13 10 9 1 3 15 7 10 9 13 1 9 0 3 1 10 3 9 9 7 10 9 0 10 9 2
12 3 3 10 9 13 9 13 13 16 13 13 2
14 15 3 0 3 9 3 13 3 9 13 16 13 15 2
13 1 15 3 3 13 13 15 10 9 1 9 13 2
14 9 3 13 13 0 3 13 9 0 10 0 15 9 2
9 0 3 10 9 9 3 16 0 2
9 0 3 9 9 1 10 13 13 2
14 15 3 9 13 0 10 9 7 9 0 1 0 13 2
15 10 3 3 13 15 13 0 16 1 0 10 3 13 13 2
6 15 3 10 9 13 2
6 3 10 9 13 13 2
16 3 0 3 9 13 10 9 13 10 9 10 9 13 10 9 2
6 10 3 9 13 15 2
20 13 3 10 9 1 9 13 10 9 1 10 9 10 0 9 13 10 9 9 2
16 10 3 9 13 13 3 3 1 10 9 1 15 7 13 13 2
11 3 3 10 0 10 0 10 0 9 13 2
14 10 3 1 10 9 13 3 13 9 3 7 9 9 2
10 10 3 3 9 7 10 9 15 13 2
15 13 3 15 3 1 10 0 9 10 9 1 10 9 13 2
18 3 1 15 0 7 0 10 9 15 3 13 7 10 9 10 1 15 2
27 3 3 15 13 13 3 15 15 0 9 13 15 1 10 9 16 3 1 10 15 9 10 9 13 10 9 2
13 13 3 3 10 9 10 9 10 1 9 9 13 2
10 13 3 3 10 10 0 9 13 15 2
4 13 3 15 2
15 9 3 1 15 0 1 9 13 7 10 0 9 9 13 2
9 13 3 3 9 10 9 13 15 2
10 0 3 13 13 15 13 1 15 13 2
4 13 3 15 2
6 3 13 9 9 9 2
18 0 3 15 13 7 10 9 3 0 13 1 0 3 16 15 13 13 2
12 1 15 3 1 10 9 3 0 10 9 13 2
19 10 3 13 3 0 0 13 7 13 9 13 10 9 13 10 0 1 9 2
26 10 3 3 9 10 9 13 3 3 1 10 9 0 7 13 3 10 9 0 13 10 9 13 10 9 2
6 13 3 3 10 9 2
14 3 15 13 3 1 10 9 2 3 10 0 2 13 2
11 10 3 13 0 9 0 3 1 9 13 2
19 10 3 9 13 3 15 7 13 9 7 9 1 10 9 0 13 1 9 2
11 13 3 9 13 15 15 1 15 13 13 2
20 10 3 1 10 9 15 13 10 3 9 9 0 13 13 7 10 9 10 9 2
19 13 3 10 9 0 3 9 9 13 7 3 15 1 15 3 0 0 13 2
12 10 3 0 7 0 1 10 0 3 13 3 2
6 13 3 13 10 9 2
13 9 3 3 15 1 9 13 10 0 1 10 9 2
19 10 3 9 13 13 15 10 13 3 13 15 7 13 3 9 1 10 9 2
9 3 3 13 13 3 1 9 13 2
18 9 3 1 3 10 0 9 15 13 3 7 13 1 10 0 10 9 2
17 13 3 10 9 10 9 3 0 3 13 16 3 10 9 10 9 2
13 9 3 0 3 0 13 13 15 7 3 3 0 2
15 9 3 3 13 13 3 9 0 13 7 10 9 9 13 2
12 10 3 0 0 13 3 10 9 13 0 13 2
15 10 3 0 15 0 0 15 13 10 9 7 9 10 9 2
13 13 3 0 3 13 15 1 10 0 15 3 13 2
20 10 3 0 13 9 10 3 0 7 0 9 1 10 0 1 9 10 3 13 2
17 10 3 10 9 7 10 0 13 16 3 0 13 13 1 0 13 2
7 1 15 13 15 0 13 2
8 10 3 9 10 9 3 0 2
12 3 3 3 10 9 7 10 0 15 0 13 2
11 10 3 10 9 0 13 3 3 15 13 2
12 3 3 15 13 15 3 1 10 0 13 3 2
28 3 1 10 9 15 3 13 10 9 10 3 15 13 7 1 10 0 3 9 0 9 1 0 9 9 15 13 2
7 0 3 10 10 9 9 2
3 13 3 2
12 3 15 3 3 1 0 9 1 10 9 13 2
11 3 10 3 13 1 9 7 3 0 13 2
11 9 3 9 10 13 13 7 9 10 13 2
46 1 9 10 9 3 3 15 13 13 0 2 15 3 3 9 3 9 3 9 7 1 0 10 1 10 9 15 7 10 9 9 0 13 9 2 0 7 10 9 1 15 13 10 9 13 2
33 10 3 3 9 13 7 13 10 0 9 13 15 2 15 13 3 9 10 9 2 9 13 10 3 9 1 15 9 10 9 13 13 2
26 10 3 10 9 10 1 9 13 13 10 9 2 16 9 7 9 2 3 0 9 0 13 10 0 9 2
25 9 3 13 2 0 1 9 13 9 3 1 10 0 9 2 10 0 10 0 9 1 10 9 13 2
16 13 3 3 9 9 9 1 15 10 9 13 13 1 10 9 2
27 9 3 3 9 3 13 3 10 0 10 1 9 9 2 10 7 13 13 10 0 15 7 3 9 13 9 2
27 3 3 3 3 3 13 10 9 2 13 10 0 13 9 7 0 9 13 10 13 1 10 9 13 10 9 2
25 10 3 9 15 3 3 13 9 2 1 15 3 10 9 13 9 10 9 7 9 13 0 9 13 2
34 13 3 10 9 1 9 0 7 0 13 1 9 2 13 10 0 9 15 13 2 16 13 3 15 7 10 1 15 0 1 10 0 9 2
36 3 3 1 15 13 15 3 1 15 10 9 2 7 10 9 15 13 9 2 16 13 0 9 10 3 0 13 10 9 2 13 7 13 10 0 2
41 1 3 10 0 9 10 3 9 13 2 10 7 0 9 10 3 13 10 13 10 0 2 10 7 1 9 7 1 9 13 2 9 7 9 13 10 9 1 0 9 2
11 1 15 3 10 9 10 9 13 13 13 2
18 13 3 9 0 2 0 9 13 13 2 10 0 9 9 13 10 9 2
17 13 3 3 15 1 0 9 13 13 2 16 0 13 2 10 9 2
12 3 16 3 10 9 10 9 0 13 13 13 2
26 16 3 15 0 13 2 10 3 9 13 10 9 13 2 16 9 13 2 10 7 9 15 16 0 13 2
10 10 3 10 0 9 0 9 9 13 2
55 16 3 10 9 13 3 7 9 13 2 13 13 10 9 1 10 13 15 13 10 9 2 10 3 9 15 13 2 1 7 10 9 0 3 13 2 7 13 7 13 13 2 3 13 13 13 15 7 13 13 10 9 7 13 2
47 3 3 13 3 10 9 10 9 2 16 13 13 2 13 0 10 9 15 7 9 2 15 13 13 2 16 3 0 13 2 13 10 9 2 16 7 9 2 13 1 15 15 0 3 13 13 2
18 13 3 13 15 1 10 9 13 9 3 13 10 9 10 9 15 13 2
7 13 3 9 12 10 0 2
33 13 3 3 15 0 1 10 9 2 7 0 13 10 3 0 9 7 0 9 13 13 10 1 9 13 15 7 13 13 3 10 13 2
10 0 3 0 9 3 1 10 9 13 2
29 1 15 3 13 7 13 10 0 2 13 13 9 10 9 2 7 13 7 3 10 9 1 9 13 13 9 10 9 2
8 3 13 0 3 1 9 13 2
54 9 3 13 10 9 1 9 7 9 0 2 1 9 3 7 9 0 10 0 13 7 0 2 15 13 13 3 10 9 7 13 10 9 10 9 1 10 13 3 1 15 9 2 16 9 0 10 9 13 10 9 15 15 2
48 1 3 10 9 10 9 1 9 13 2 13 2 16 13 2 10 0 9 2 0 13 7 0 2 10 0 9 7 9 2 16 9 9 0 0 7 0 2 13 13 10 9 10 9 7 10 9 2
28 13 3 0 3 9 10 9 0 1 10 9 2 13 7 3 0 9 0 2 3 10 9 2 16 13 2 13 2
9 0 3 15 3 3 0 13 9 2
41 9 3 3 1 15 13 10 9 13 2 3 10 1 10 0 9 10 0 9 3 13 13 1 10 9 2 7 13 10 0 7 9 0 3 3 10 9 7 0 13 2
11 15 3 3 9 0 3 10 0 9 13 2
27 16 3 3 9 7 9 13 10 9 7 1 10 9 13 10 9 13 2 15 1 9 10 9 9 13 13 2
22 3 3 3 10 9 13 0 10 9 10 9 2 7 13 15 13 0 13 13 10 0 2
50 13 3 1 3 13 3 13 10 13 13 7 13 10 9 2 16 10 1 9 9 0 9 3 9 2 16 3 15 16 9 0 7 13 0 9 10 13 13 7 13 9 1 9 7 9 0 13 0 9 2
9 13 3 15 0 3 13 1 9 2
28 13 3 15 13 10 0 7 13 13 2 3 13 10 0 0 2 3 3 1 0 13 0 7 13 1 10 9 2
25 16 3 10 9 13 2 12 10 0 13 1 10 9 3 1 9 13 9 1 7 9 1 10 13 2
7 3 12 10 0 9 13 2
17 10 3 3 10 9 9 13 0 7 13 10 1 10 9 9 13 2
21 13 3 10 9 10 9 9 13 3 1 15 0 10 9 13 2 13 1 10 9 2
15 3 3 3 13 13 10 9 15 1 10 13 10 9 13 2
37 0 3 13 1 10 9 0 13 7 0 10 9 10 9 2 15 13 10 9 10 10 9 9 13 13 7 13 0 1 10 0 9 3 7 9 13 2
21 15 3 13 13 10 9 9 2 16 12 10 0 1 9 13 12 10 9 13 13 2
13 10 3 9 1 9 13 15 13 10 10 9 13 2
27 13 3 3 15 3 10 10 9 1 9 9 13 13 2 7 16 10 15 9 0 13 1 10 9 0 13 2
23 15 3 13 3 0 13 10 9 16 10 0 13 12 2 10 12 7 12 10 0 9 13 2
21 3 3 1 0 13 10 9 10 9 16 9 1 9 13 1 15 2 15 9 13 2
4 13 3 3 2
28 1 15 10 3 9 13 7 9 13 13 13 7 13 10 9 1 9 2 15 10 3 9 2 10 7 9 13 2
11 9 3 10 9 13 2 10 7 13 13 2
13 3 10 9 7 10 9 10 9 1 10 9 13 2
16 1 0 3 15 10 9 13 2 3 9 13 7 0 0 9 2
19 13 3 3 15 10 9 16 10 9 15 13 2 16 3 9 13 1 15 2
54 3 10 9 10 9 13 2 3 0 3 10 9 7 0 10 1 15 13 13 7 13 2 16 13 10 9 2 0 9 13 15 10 10 9 9 2 9 3 3 12 7 12 1 9 0 10 1 9 9 13 1 9 13 2
27 15 7 13 1 10 15 9 13 3 0 13 10 9 10 9 16 13 2 0 3 3 2 13 2 0 0 2
37 10 3 13 10 3 13 1 10 9 13 10 9 2 16 3 13 15 9 7 9 10 1 15 9 13 2 15 13 7 13 10 9 1 10 0 13 2
84 15 3 3 10 9 9 7 9 13 0 1 10 9 7 9 2 0 7 9 2 9 7 9 9 7 9 13 2 15 10 0 1 9 13 2 1 7 10 9 3 0 13 15 13 2 3 1 0 9 13 2 7 9 3 10 9 2 3 9 7 10 9 2 10 13 13 13 16 0 13 3 3 9 10 9 10 10 9 13 7 13 1 15 2
13 0 3 10 9 9 7 0 10 10 9 9 13 2
26 13 3 10 9 10 9 13 10 3 15 10 0 0 0 9 2 10 7 1 10 9 10 9 13 0 2
6 15 3 13 9 9 2
16 0 3 13 10 3 9 0 13 2 0 7 1 15 13 9 2
27 10 3 9 13 0 15 16 9 13 9 3 12 9 9 2 9 7 12 2 7 10 0 9 3 10 9 2
19 13 3 13 15 15 2 10 9 1 9 7 9 0 2 0 7 15 13 2
39 13 3 15 0 3 9 10 9 13 1 9 3 13 2 13 10 9 0 7 0 2 13 2 7 13 1 10 13 16 10 0 13 0 0 9 13 3 13 2
33 13 3 3 10 9 13 2 16 3 13 10 0 7 0 2 16 3 13 13 10 3 9 2 0 13 9 7 13 10 1 15 9 2
15 0 3 3 13 0 9 13 7 13 0 13 10 0 13 2
26 3 15 3 1 0 9 7 9 9 0 13 2 16 12 9 9 9 3 0 1 9 13 7 9 13 2
10 15 3 13 13 9 9 0 10 9 2
25 15 3 7 13 13 7 13 7 13 7 13 15 3 13 0 13 7 13 0 2 7 3 13 0 2
24 9 3 2 16 13 2 0 9 10 9 13 13 10 1 15 9 7 9 2 0 7 0 13 2
11 1 3 15 10 0 7 0 13 9 9 2
64 10 3 0 0 3 13 1 10 0 9 7 13 9 13 2 16 3 13 15 10 0 7 0 13 2 9 13 9 0 1 10 9 2 7 13 10 0 3 9 9 2 3 9 0 2 3 9 9 2 3 0 15 2 3 0 9 9 2 3 3 9 3 13 2
16 3 3 13 1 0 10 9 10 13 7 13 0 1 15 13 2
21 3 0 15 13 10 0 13 2 9 3 13 1 0 10 9 2 7 13 7 13 2
35 3 3 10 0 10 9 7 0 0 2 9 3 9 7 9 2 0 1 15 13 2 7 9 10 0 13 3 1 10 9 2 16 13 9 2
31 10 3 3 13 10 9 7 13 10 9 13 10 9 2 7 10 0 13 3 7 13 10 9 2 0 13 10 9 10 13 2
7 0 3 3 15 10 9 2
13 13 3 10 9 10 0 1 10 9 13 10 9 2
32 0 3 3 3 15 13 2 0 7 10 10 9 0 2 16 13 9 2 7 0 13 10 9 10 9 7 10 1 10 9 9 2
25 9 3 3 13 3 9 7 9 3 7 9 10 0 9 2 1 10 0 9 10 9 10 0 13 2
24 3 3 3 13 10 9 1 0 10 9 0 13 10 0 2 7 13 1 15 0 13 7 13 2
10 9 3 13 1 0 13 10 9 9 2
9 3 10 3 15 13 1 9 13 2
24 10 3 3 9 15 13 1 10 9 2 7 13 0 13 10 9 10 9 13 7 13 10 9 2
21 9 3 0 7 9 10 13 13 2 16 13 10 9 15 7 13 1 10 9 13 2
32 10 3 9 15 3 13 13 2 10 7 9 13 3 0 3 15 3 13 7 13 2 13 7 10 0 9 7 9 15 13 13 2
21 3 3 3 15 13 7 0 13 9 2 1 0 0 7 0 0 9 7 0 13 2
9 10 3 9 9 10 3 9 13 2
36 0 3 10 9 2 15 3 9 13 10 13 10 0 9 2 13 3 13 2 3 13 7 10 9 2 7 3 10 9 10 9 10 9 0 13 2
13 10 3 13 9 13 10 9 1 10 9 0 13 2
11 13 3 1 12 3 0 15 0 7 0 2
32 13 3 0 1 9 10 9 9 9 2 9 9 12 2 9 12 9 2 9 9 12 2 1 7 15 1 9 0 15 3 9 2
14 3 3 3 13 15 9 7 13 9 13 1 10 9 2
17 13 3 3 13 16 13 15 7 13 13 2 10 7 15 13 13 2
9 3 1 3 0 10 9 3 13 2
36 1 3 10 9 3 9 13 2 16 1 9 9 13 2 3 9 13 0 7 0 9 13 2 15 7 13 13 7 13 1 9 7 13 3 13 2
11 3 13 3 13 13 2 7 10 13 13 2
20 10 3 13 0 13 10 0 10 9 2 1 15 2 13 2 3 9 3 13 2
10 13 3 10 13 10 9 13 3 13 2
9 10 3 13 10 10 13 13 9 2
16 7 0 13 15 2 3 13 10 13 2 13 0 13 15 13 2
11 9 3 13 10 9 1 15 10 9 13 2
30 10 3 9 13 3 1 15 10 0 9 2 16 3 9 13 10 0 2 7 13 10 9 2 15 7 10 9 13 13 2
14 13 3 15 10 0 9 1 10 9 3 13 0 9 2
7 13 3 3 13 1 9 2
23 3 3 13 1 9 13 2 3 15 7 15 9 2 16 13 9 7 9 3 7 3 13 2
8 10 3 3 9 0 13 9 2
16 9 3 13 10 9 3 13 2 7 0 10 13 9 13 15 2
50 10 3 3 0 7 0 1 9 9 7 9 2 1 10 9 13 7 10 9 10 9 13 2 13 0 7 0 2 13 10 9 9 0 10 9 2 15 10 9 13 10 9 2 9 9 13 1 0 15 2
40 10 3 0 7 0 0 7 13 10 9 3 3 2 0 13 3 13 0 9 7 0 9 2 7 13 1 10 9 2 9 13 7 9 2 15 3 10 13 13 2
13 10 3 0 7 0 10 9 9 1 10 9 13 2
15 0 3 3 10 9 13 2 16 13 2 3 13 9 0 2
37 1 3 0 10 9 13 3 9 10 0 1 9 13 2 7 13 10 9 10 9 10 9 0 7 0 2 13 10 0 16 0 1 15 10 9 13 2
24 0 3 9 13 10 9 2 10 13 1 10 0 0 3 13 2 16 3 3 13 13 0 13 2
25 3 3 13 0 13 9 2 0 2 13 2 10 9 1 9 13 2 3 13 15 7 13 13 13 2
17 10 3 3 0 9 9 13 2 3 1 10 9 13 7 9 13 2
26 10 3 9 2 15 0 13 10 9 7 0 9 13 2 3 13 3 13 10 1 10 9 7 10 9 2
46 3 3 2 16 9 13 2 13 13 10 9 2 13 3 13 10 0 9 7 9 1 10 0 9 10 9 2 1 15 13 0 13 15 2 7 1 15 3 10 13 15 13 7 9 13 2
8 3 3 15 10 13 9 13 2
47 10 3 3 9 10 9 9 3 9 7 9 9 7 9 13 2 16 10 3 10 13 9 0 1 0 9 9 13 13 0 2 15 7 1 9 10 9 13 3 3 7 3 13 1 10 9 2
31 13 3 9 3 9 7 9 0 0 0 13 10 9 10 9 0 3 13 7 1 0 0 13 7 13 10 0 13 7 13 2
13 13 3 16 3 9 13 1 0 3 13 10 13 2
20 3 3 1 10 0 15 0 1 9 13 13 2 9 0 7 9 13 10 9 2
17 10 3 13 1 9 7 0 1 10 9 13 13 13 1 10 9 2
32 10 3 1 9 7 9 9 0 0 10 1 9 9 13 2 3 3 1 10 9 3 10 0 9 3 10 9 7 10 9 13 2
44 10 3 9 10 9 15 0 13 2 9 3 13 2 9 7 13 2 7 9 0 7 9 9 13 2 7 9 10 0 13 3 0 2 3 0 0 15 3 9 7 9 9 13 2
16 3 15 3 13 13 7 13 0 3 1 9 13 10 9 9 2
27 13 3 15 2 16 13 2 0 1 15 16 0 10 9 13 15 10 9 2 0 3 2 13 2 13 9 2
9 13 3 3 3 15 0 1 9 2
31 13 3 10 9 10 9 3 10 9 7 10 9 1 9 10 0 2 13 3 0 2 7 0 2 16 13 10 9 2 9 2
10 3 3 3 3 9 0 13 10 0 2
8 13 3 1 10 9 10 9 2
11 9 3 7 9 15 0 0 13 2 13 2
14 3 3 10 1 9 13 15 13 2 3 0 13 9 2
20 13 3 15 10 0 15 9 3 13 2 13 2 3 3 15 15 10 13 13 2
18 13 3 1 9 2 3 0 7 0 1 9 2 7 3 13 7 0 2
28 10 3 13 10 9 13 13 2 10 3 9 1 9 13 2 9 7 0 7 9 13 13 1 9 0 1 9 2
18 13 3 9 3 0 13 3 3 13 10 0 2 13 1 10 0 0 2
47 3 10 0 3 13 2 10 3 9 13 7 13 2 1 7 10 9 3 1 9 13 2 13 7 13 16 15 13 10 3 2 3 3 10 9 13 7 13 16 3 1 9 3 13 15 13 2
21 3 15 13 3 0 9 2 7 16 3 9 13 0 16 1 9 13 10 15 9 2
51 0 3 10 9 13 9 7 9 2 15 0 13 10 0 7 0 9 2 1 0 13 9 3 7 9 0 13 1 10 9 2 9 7 3 9 13 10 0 2 13 10 3 0 7 0 15 13 9 7 9 2
33 13 3 3 9 0 0 9 2 16 3 15 10 9 7 0 13 0 7 13 2 13 1 15 7 13 0 9 0 15 13 10 13 2
38 13 3 3 9 0 2 10 0 15 7 0 13 9 0 13 2 13 10 9 13 2 3 1 9 2 0 13 7 13 9 0 2 0 0 7 0 13 2
34 0 3 3 3 0 13 10 9 10 9 2 7 0 10 9 10 9 2 3 3 1 10 13 2 7 1 10 0 13 13 13 10 9 2
79 3 0 9 7 9 13 10 1 15 10 15 9 2 15 9 3 7 9 1 10 0 10 9 13 9 13 7 9 10 9 2 10 7 9 13 13 2 1 15 0 13 13 2 16 0 13 2 16 9 2 16 0 2 3 3 0 10 13 7 13 10 9 13 0 2 16 1 0 13 2 7 3 0 2 16 0 13 9 2
28 15 3 3 13 3 7 3 3 0 13 10 0 13 13 1 10 9 9 16 3 0 13 10 10 9 1 15 2
23 3 9 13 9 0 9 10 3 0 2 15 13 1 9 15 13 10 9 1 15 2 13 2
18 9 2 13 10 9 2 13 0 2 15 13 10 9 1 10 9 13 2
7 3 3 3 13 9 15 2
15 13 10 9 2 3 3 3 2 13 2 1 9 9 13 2
8 15 3 3 13 1 10 9 2
46 10 3 13 3 13 9 10 13 13 2 7 13 13 1 9 0 9 13 2 1 15 13 10 9 10 0 13 10 9 2 16 3 0 13 7 0 2 13 13 2 9 15 10 0 13 2
19 3 3 9 10 9 2 7 9 13 10 9 2 9 0 13 10 9 15 2
22 13 3 13 10 0 7 0 1 10 0 13 2 10 7 0 3 13 7 13 10 9 2
45 13 3 1 10 9 9 0 1 9 2 16 1 9 13 10 9 10 9 7 10 9 9 13 2 3 7 0 10 9 3 0 3 0 9 3 1 9 0 7 0 9 0 7 9 2
11 3 3 10 3 0 10 9 0 13 9 2
12 3 10 3 10 0 9 13 9 13 13 9 2
19 3 15 2 16 9 13 2 9 13 9 9 2 0 15 10 0 13 9 2
48 10 3 9 9 3 1 0 7 0 13 9 10 9 2 7 13 0 13 7 13 16 13 10 9 2 7 0 3 0 13 13 15 1 9 13 2 7 0 13 7 0 1 15 13 13 7 13 2
18 3 1 15 13 3 13 13 7 13 13 2 16 10 9 13 9 9 2
8 9 3 3 1 10 9 13 2
17 10 3 0 0 9 1 10 13 3 13 3 13 13 7 13 13 2
25 3 3 10 9 13 13 15 10 9 2 1 9 7 13 3 13 0 13 7 0 3 10 0 13 2
24 13 3 0 1 9 3 13 2 0 9 1 10 9 13 2 0 10 9 7 9 7 9 0 2
11 1 0 9 0 10 9 10 0 9 13 2
28 13 3 3 1 9 7 9 1 9 2 15 15 13 2 10 1 10 9 13 9 10 9 10 9 1 9 13 2
10 3 3 10 15 9 10 0 0 13 2
50 3 13 10 0 2 3 3 13 1 10 9 2 7 13 7 13 15 13 2 3 3 2 7 9 0 0 13 0 3 9 13 3 9 7 9 2 16 3 9 13 7 9 0 10 13 10 13 7 13 2
27 3 3 3 3 9 1 10 0 7 0 9 13 2 7 1 9 15 13 10 13 9 3 10 0 7 0 2
18 9 3 13 10 9 3 0 1 9 13 2 9 7 10 9 10 0 2
26 0 3 10 9 2 12 9 13 2 13 3 10 13 1 10 9 2 7 1 9 9 13 1 10 9 2
13 13 3 10 3 0 9 13 2 10 7 0 9 2
25 3 13 13 2 10 3 1 10 9 13 2 10 7 1 10 10 9 9 13 3 3 3 7 3 2
16 16 3 13 2 0 13 9 10 9 2 3 13 13 7 3 2
19 13 3 3 10 9 15 0 3 13 2 13 3 13 10 13 7 3 13 2
17 0 3 15 13 9 2 16 1 15 13 10 9 13 13 7 13 2
7 3 15 3 9 10 9 2
8 13 3 13 10 10 9 9 2
9 10 3 0 15 3 0 13 13 2
52 10 3 0 7 0 3 9 13 1 10 9 2 10 7 0 7 0 1 9 13 2 16 3 3 10 1 10 13 13 9 0 3 2 0 7 7 0 13 10 9 2 1 10 9 10 9 13 3 1 10 13 2
12 3 3 10 3 9 10 13 1 0 13 13 2
37 3 3 13 3 10 9 2 16 13 15 3 9 9 13 7 10 9 13 2 13 1 10 9 10 9 10 9 7 10 9 2 1 10 13 13 13 2
23 3 15 3 3 1 10 3 9 0 13 2 15 0 1 10 9 10 0 13 13 10 9 2
21 13 3 10 9 13 10 3 13 13 10 9 2 10 7 9 0 13 13 13 9 2
17 1 15 3 3 13 10 0 7 13 3 1 9 13 1 10 9 2
26 10 3 13 2 15 9 0 2 7 15 3 0 2 13 10 13 2 0 13 7 1 9 0 9 9 2
18 13 3 10 9 3 1 9 13 7 9 1 0 0 13 9 7 0 2
14 10 3 3 13 13 9 13 1 10 9 1 10 9 2
23 3 3 3 0 13 7 9 10 9 13 10 9 2 9 13 16 1 9 7 16 13 13 2
24 3 13 3 3 13 2 10 7 9 13 9 13 2 16 0 10 13 13 7 3 3 7 3 2
11 13 3 10 9 10 9 10 9 1 0 2
17 3 13 3 9 1 10 13 9 0 13 13 10 9 1 10 9 2
46 3 3 10 13 13 1 15 2 16 3 10 9 13 10 0 7 0 9 2 10 13 3 13 2 7 3 9 13 9 1 15 10 10 15 13 2 7 13 3 13 16 0 13 10 13 2
18 13 3 10 9 3 9 13 9 13 13 9 7 0 1 0 9 9 2
49 10 3 3 0 9 0 13 13 1 0 9 9 10 9 2 16 13 2 10 7 10 9 9 0 1 0 7 0 9 1 0 7 0 13 9 2 10 0 9 10 9 0 7 13 1 10 9 13 2
30 16 3 10 9 10 1 10 9 0 0 3 10 0 7 0 13 2 3 10 1 10 13 9 0 10 9 13 7 0 2
41 9 3 3 10 9 2 13 0 15 10 0 9 1 10 9 2 7 13 16 3 15 10 0 13 1 10 9 2 3 10 3 2 13 2 15 13 10 9 10 0 2
26 15 3 3 10 9 13 10 9 0 3 13 13 2 3 7 10 9 13 2 7 10 9 13 10 13 2
18 3 3 10 9 0 0 15 13 13 7 0 2 16 13 13 10 9 2
15 0 13 10 1 10 9 1 10 13 13 9 1 10 9 2
13 15 3 2 13 2 0 1 10 9 15 13 9 2
12 13 3 3 3 1 9 9 0 1 10 9 2
6 3 3 0 9 13 2
11 3 0 13 7 3 0 0 0 13 15 2
13 3 3 13 0 9 15 9 2 7 3 9 13 2
14 1 3 3 0 7 10 0 9 3 13 9 7 13 2
14 10 3 1 10 9 10 9 9 9 15 10 9 13 2
26 9 3 10 9 10 9 1 10 9 15 10 9 13 2 13 16 10 9 3 13 0 3 9 13 0 2
25 9 3 13 15 0 10 9 16 13 1 10 9 15 13 2 10 13 2 13 2 9 7 9 13 2
13 15 3 10 0 13 9 3 13 9 2 15 13 2
32 9 3 2 13 15 10 9 3 3 10 9 7 3 13 2 3 15 0 2 13 2 9 13 1 9 12 9 0 13 10 9 2
18 9 3 10 9 2 9 0 10 9 0 13 2 3 2 13 2 13 2
10 0 3 9 15 15 0 13 1 15 2
13 13 3 3 10 1 9 13 1 15 13 10 9 2
22 13 3 3 13 10 9 3 2 7 13 9 15 3 3 3 3 13 0 9 0 9 2
17 10 3 3 13 10 13 10 9 13 2 0 2 13 2 13 15 2
8 13 3 15 9 0 9 13 2
7 13 3 13 0 15 13 2
28 9 3 1 10 13 15 13 9 13 1 10 13 2 3 15 3 2 13 2 7 13 15 10 13 1 10 13 2
24 0 3 15 13 1 9 13 1 9 9 2 3 13 2 13 2 3 13 3 3 13 13 0 2
24 10 3 3 10 9 9 13 15 16 3 13 15 3 3 16 3 13 10 13 16 10 13 13 2
48 10 3 1 10 9 7 10 9 9 3 0 13 10 1 10 9 9 7 9 2 7 3 10 9 9 13 0 9 7 0 9 0 7 0 2 7 10 9 13 0 7 0 1 9 0 7 0 2
35 9 3 13 3 10 0 10 13 1 10 9 13 2 3 9 10 13 2 3 0 7 0 13 9 2 9 3 7 9 1 9 13 10 9 2
10 15 1 9 3 0 13 0 15 13 2
19 12 3 9 1 10 12 9 13 1 10 9 2 10 3 10 9 13 13 2
7 10 3 10 13 13 13 2
5 15 3 3 13 2
6 16 3 13 2 13 2
7 15 3 3 13 0 0 2
46 3 3 3 15 13 10 0 9 2 15 3 1 15 0 13 2 7 10 0 9 13 2 15 13 1 10 9 13 10 0 2 3 3 13 3 10 9 7 10 9 10 9 10 9 13 2
9 10 3 3 3 13 1 10 9 2
12 3 9 3 0 13 3 9 0 7 9 0 2
4 9 3 13 2
15 3 9 9 3 0 9 13 9 3 9 3 9 7 9 2
8 0 3 3 7 0 13 15 2
15 13 3 1 10 9 10 3 13 2 16 10 0 9 13 2
38 3 3 1 10 9 13 10 9 10 9 2 13 2 16 13 2 10 9 7 10 9 2 16 13 0 1 10 0 7 9 0 0 13 10 9 10 13 2
34 3 3 3 10 0 10 0 10 9 13 2 3 13 13 1 9 7 9 9 7 9 2 13 2 16 9 2 13 7 13 1 10 9 2
36 13 3 3 9 0 1 10 9 2 7 10 0 9 3 3 13 7 0 10 0 13 2 16 0 9 15 10 1 10 9 9 9 13 10 9 2
45 3 3 13 0 9 2 16 0 3 7 0 10 9 13 2 9 3 1 10 9 13 7 3 9 13 1 10 9 7 10 9 13 2 7 3 7 3 1 10 9 13 1 10 9 2
26 3 3 9 7 9 13 13 10 3 13 9 13 2 7 0 9 1 9 7 9 2 3 10 9 13 2
14 13 3 10 9 1 10 0 13 1 15 9 9 13 2
13 13 3 3 0 0 15 7 0 2 7 3 0 2
23 13 3 10 13 1 15 16 10 13 13 2 13 7 10 13 2 10 13 10 13 13 0 2
28 0 3 10 9 9 3 10 9 0 13 13 7 0 0 9 2 9 7 3 10 1 9 10 9 9 9 13 2
17 13 3 3 10 0 9 10 9 0 7 1 9 3 13 9 13 2
28 3 13 15 2 16 9 13 2 10 9 3 13 7 13 1 9 10 1 10 9 2 7 13 3 13 7 13 2
8 10 3 9 1 10 0 13 2
60 15 3 13 13 16 13 13 2 7 0 1 9 10 9 7 9 13 13 7 9 1 10 0 2 7 3 13 3 15 2 7 10 9 13 13 2 16 3 15 13 0 13 13 2 13 10 9 2 7 13 15 10 0 7 13 15 1 10 0 2
13 10 3 9 15 13 10 9 2 9 10 13 13 2
38 13 3 15 9 9 13 2 7 13 0 9 9 13 13 13 7 13 1 10 0 13 7 3 13 2 13 13 10 13 15 15 13 10 10 9 13 9 2
12 3 0 13 10 1 10 9 7 10 9 9 2
28 9 3 2 16 13 2 13 1 10 9 2 3 9 7 9 15 13 2 9 7 1 9 7 9 1 9 13 2
25 9 3 3 9 3 9 7 9 1 3 9 3 9 7 9 10 0 9 13 2 16 3 13 13 2
25 10 3 3 0 12 9 10 3 3 13 1 9 2 7 1 10 0 7 10 0 13 10 9 9 2
26 10 3 0 0 13 3 13 1 15 13 2 7 3 10 0 10 9 1 10 9 7 10 13 9 13 2
20 3 3 1 15 13 3 13 1 15 2 15 13 10 1 9 7 9 0 13 2
30 3 10 0 13 10 0 9 9 13 0 10 0 2 7 10 0 13 2 1 9 7 9 2 3 13 1 9 7 9 2
9 3 3 0 13 3 0 10 9 2
31 3 3 10 10 9 9 15 13 9 13 2 10 9 3 9 10 9 7 10 9 13 1 9 1 10 9 7 10 0 9 2
10 3 13 3 9 0 15 13 10 9 2
23 10 3 3 9 3 13 1 10 0 13 3 0 2 16 13 16 0 15 0 10 9 13 2
29 10 3 9 9 9 2 16 13 15 1 9 10 1 9 13 1 15 2 13 16 3 10 9 13 7 10 9 3 2
18 10 3 9 15 3 2 16 13 2 13 10 0 1 10 13 10 9 2
17 9 3 1 10 13 13 13 10 0 9 13 10 1 12 9 13 2
12 3 0 13 10 1 9 9 15 13 7 0 2
8 13 3 10 9 0 10 9 2
24 9 13 9 0 13 3 1 9 2 10 3 9 3 13 7 13 2 10 7 9 0 13 13 2
24 9 3 16 15 3 10 13 13 2 3 3 0 2 7 0 1 9 13 7 9 13 10 9 2
32 13 3 10 0 9 2 1 0 13 10 9 10 9 2 3 13 15 13 2 3 16 0 3 0 3 0 7 3 13 10 13 2
10 15 3 0 13 7 0 2 15 13 2
7 10 3 13 13 10 9 2
16 10 3 0 0 15 9 13 13 16 10 9 0 13 10 9 2
7 13 3 1 10 9 13 2
15 3 10 3 15 13 3 2 0 7 9 15 13 13 13 2
42 3 1 10 9 1 10 9 10 9 10 0 13 9 2 15 3 13 13 13 2 7 13 10 9 13 16 15 15 13 0 15 13 2 16 15 13 1 10 0 13 9 2
11 3 3 3 10 1 10 9 0 13 15 2
51 0 3 3 13 9 0 1 10 9 13 10 9 2 7 3 13 10 9 10 9 3 13 2 0 13 10 0 9 7 0 10 0 2 16 3 13 7 13 10 9 16 13 10 13 9 9 7 1 9 13 2
16 3 13 15 13 2 7 1 9 7 9 9 13 10 9 13 2
19 13 3 9 13 3 13 10 9 2 7 9 1 9 7 9 10 9 13 2
10 10 3 0 13 13 9 13 10 9 2
19 15 3 13 0 7 13 2 7 9 13 10 0 9 0 9 7 9 9 2
20 3 3 13 13 10 13 7 13 2 0 13 9 7 9 9 0 7 9 0 2
42 3 3 10 13 1 15 0 7 13 1 10 9 13 2 3 2 16 9 13 2 13 16 10 9 9 13 7 1 9 15 0 13 2 7 3 16 3 9 0 15 13 2
9 1 3 0 9 9 9 13 0 2
7 9 3 0 9 0 13 2
17 1 15 9 9 0 13 7 9 13 1 10 13 9 2 16 9 2
18 3 3 13 13 13 10 9 16 9 3 13 0 16 9 0 3 13 2
29 1 3 3 15 0 13 9 9 7 9 2 15 13 0 10 9 9 2 16 3 13 1 9 2 3 7 1 9 2
36 10 3 13 9 1 15 2 16 3 3 15 10 9 9 0 13 2 16 9 13 2 0 3 13 3 10 9 1 10 9 7 10 9 13 9 2
4 13 3 15 2
27 10 0 10 9 1 9 10 3 9 13 13 1 10 9 3 13 2 13 9 7 9 0 2 0 7 15 2
27 10 3 1 9 3 1 0 13 9 2 13 15 7 13 2 3 7 13 1 10 9 10 9 10 13 13 2
13 3 3 3 10 9 13 10 0 7 0 15 13 2
50 3 3 9 1 10 9 13 10 1 9 13 1 10 9 13 3 3 0 13 7 13 10 10 9 9 2 0 7 9 0 0 13 2 0 16 0 13 2 16 3 3 7 9 13 15 13 0 9 13 2
26 9 3 3 13 3 10 9 2 16 1 10 9 13 0 2 10 9 13 9 2 16 0 13 10 13 2
28 3 15 3 3 13 7 3 15 2 16 3 13 13 0 0 1 10 9 13 2 13 10 13 0 13 10 0 2
16 3 9 13 13 7 9 13 0 7 0 2 13 7 10 0 2
38 10 3 3 0 9 9 13 10 9 13 2 3 1 10 0 9 2 15 13 10 9 1 9 13 2 3 0 0 10 9 13 7 0 10 9 13 9 2
28 3 3 3 15 13 9 0 3 10 9 9 1 10 0 15 9 7 9 13 10 9 2 15 3 10 9 13 2
38 13 3 0 1 9 2 10 3 15 3 13 13 7 3 1 9 7 9 10 9 2 10 7 0 13 7 0 3 3 13 0 1 15 16 13 10 9 2
25 13 3 1 10 9 7 10 9 13 2 13 16 3 10 9 7 3 1 9 7 9 9 13 13 2
26 13 3 10 9 3 10 9 3 13 7 10 9 0 13 10 9 13 9 2 10 9 13 1 9 13 2
52 15 3 10 9 3 13 7 10 9 13 7 10 9 2 13 3 10 9 13 10 9 2 3 7 13 10 9 3 2 9 13 1 15 3 13 3 7 13 13 0 13 2 3 10 1 15 3 1 9 13 13 2
29 13 3 13 2 13 13 10 0 9 3 10 9 0 13 7 0 10 10 9 9 2 7 1 9 9 7 9 13 2
6 3 3 13 10 9 2
25 10 3 10 9 9 3 9 13 2 7 9 10 9 2 7 13 1 10 9 13 0 13 10 9 2
49 9 3 13 13 9 0 1 10 9 2 7 1 10 9 9 7 9 9 13 1 9 2 15 15 13 0 1 9 2 13 10 9 9 7 9 2 9 7 9 1 10 9 13 7 10 9 13 9 2
8 15 13 9 10 9 7 9 2
47 3 15 13 10 13 16 13 3 13 2 13 7 3 13 9 2 7 10 9 10 9 13 9 2 15 2 13 15 13 10 9 1 10 9 0 13 2 3 2 13 2 1 10 9 0 13 2
18 3 3 13 13 10 13 3 13 2 7 10 9 9 3 13 10 9 2
9 13 3 10 3 13 10 3 13 2
16 9 3 3 9 2 7 9 13 10 15 10 13 7 13 15 2
17 13 3 3 9 3 9 1 15 7 9 13 2 7 0 9 9 2
36 1 15 3 9 13 13 2 1 9 13 7 13 9 13 9 7 9 2 9 7 13 2 3 3 15 13 2 9 7 2 16 13 15 2 13 2
8 3 15 3 13 1 10 0 2
27 9 3 10 0 1 10 1 9 9 13 10 9 0 13 2 15 15 13 13 9 1 10 13 10 9 13 2
27 0 3 9 13 10 9 9 3 9 3 9 7 0 0 15 1 15 13 13 13 2 9 7 9 13 0 2
43 10 3 3 9 7 9 2 7 9 9 0 1 9 13 2 7 10 0 13 10 13 1 10 0 9 13 13 0 10 9 13 2 3 13 10 9 10 3 13 1 10 9 2
21 1 15 3 9 0 13 13 9 16 13 13 15 13 1 9 2 3 13 10 0 2
14 9 3 3 13 15 2 7 13 1 0 9 16 9 2
14 13 3 3 10 9 15 13 3 9 1 10 9 13 2
15 3 9 9 15 13 13 1 9 10 9 1 10 0 9 2
7 15 13 0 10 9 13 2
16 10 3 9 3 10 9 13 13 7 10 0 9 13 9 13 2
12 13 3 3 9 15 10 9 1 15 13 9 2
7 3 9 13 1 15 13 2
3 13 9 2
6 3 3 15 9 13 2
10 0 3 3 13 13 10 13 10 9 2
9 13 3 10 9 10 9 10 9 2
5 3 3 13 13 2
16 15 13 3 7 13 10 9 15 3 10 9 13 7 10 15 2
20 0 3 13 9 1 10 9 16 3 13 10 9 13 10 0 7 13 10 13 2
12 3 13 3 10 0 9 7 13 3 10 9 2
17 3 10 3 9 13 9 10 13 9 9 1 0 9 13 7 9 2
8 3 3 3 10 0 9 13 2
9 3 3 13 13 15 10 9 0 2
11 3 3 13 9 1 9 13 10 9 9 2
6 15 13 10 9 13 2
7 13 3 10 9 9 13 2
9 10 3 9 3 13 13 0 9 2
8 13 3 10 9 13 13 13 2
6 3 15 3 3 13 2
10 9 3 13 3 3 3 1 9 0 2
15 10 3 1 9 13 9 1 10 9 10 9 9 0 13 2
12 10 3 0 9 13 13 9 7 9 13 0 2
9 9 3 13 13 1 9 13 15 2
10 13 3 3 10 0 9 9 10 9 2
6 3 15 3 0 13 2
13 0 3 3 3 3 13 10 9 0 7 0 13 2
12 10 3 9 0 3 13 3 10 9 10 9 2
4 0 10 9 2
11 0 3 10 0 0 13 10 10 9 9 2
17 3 3 3 3 9 0 7 9 13 1 10 9 0 0 9 13 2
14 0 3 0 7 0 13 3 16 13 9 1 9 0 2
7 3 3 15 1 9 13 2
18 10 3 9 10 9 3 0 13 13 1 10 9 16 13 1 10 9 2
5 16 3 13 13 2
19 1 3 10 9 3 13 13 1 9 10 9 10 0 7 10 9 0 13 2
7 9 3 13 13 10 9 2
13 13 3 3 9 3 9 0 13 10 9 10 9 2
11 10 3 0 3 15 13 3 0 7 0 2
17 13 3 3 9 3 1 9 13 16 10 9 3 3 13 0 9 2
7 0 3 13 0 0 15 2
13 3 0 13 10 9 1 15 1 10 10 9 9 2
22 3 3 10 0 9 9 9 13 3 13 15 0 13 10 9 0 7 0 1 10 9 2
17 13 3 1 9 7 9 9 13 3 10 9 13 7 13 10 9 2
27 1 3 15 9 0 7 9 13 9 10 9 0 3 9 9 7 9 1 9 9 10 9 7 10 9 13 2
16 15 3 1 10 9 13 9 10 9 13 9 13 1 10 9 2
16 10 3 10 1 15 9 13 0 3 9 7 0 0 15 13 2
2 13 2
9 3 0 15 7 0 10 13 13 2
11 1 3 0 3 10 0 0 3 0 13 2
13 15 13 10 9 15 0 7 15 0 13 3 0 2
9 15 3 13 0 1 10 13 13 2
10 3 9 1 13 15 9 0 10 9 2
10 3 3 3 13 10 9 13 9 9 2
8 10 3 3 9 3 13 13 2
10 1 3 10 9 1 10 3 13 13 2
11 10 3 0 3 15 13 15 9 7 9 2
6 0 9 13 10 9 2
9 3 13 15 0 13 1 10 9 2
10 3 1 15 10 9 13 0 10 9 2
20 1 3 10 1 9 10 9 9 13 1 9 3 9 3 9 7 9 1 9 2
11 10 3 0 13 7 13 1 9 9 13 2
15 10 3 0 9 10 0 7 0 10 9 3 13 1 9 2
14 13 3 7 13 10 3 9 13 1 9 16 13 15 2
8 3 0 3 13 7 13 13 2
13 1 3 10 9 3 0 10 9 10 9 3 13 2
9 10 3 3 15 3 13 10 9 2
7 13 3 3 9 9 13 2
12 10 3 9 3 1 9 13 10 10 9 13 2
15 3 3 13 3 10 9 10 10 9 9 1 10 9 9 2
12 3 3 15 13 10 9 1 10 1 10 9 2
12 15 3 13 9 7 15 9 10 13 10 9 2
13 10 3 3 1 10 9 9 0 1 9 9 13 2
11 3 3 13 3 0 10 13 3 10 0 2
12 13 3 15 3 9 10 9 3 13 7 13 2
19 3 3 13 0 16 10 0 9 0 13 10 0 13 9 10 9 10 9 2
14 3 0 3 0 9 1 9 13 10 9 7 9 9 2
18 0 3 9 13 1 10 9 0 13 3 1 10 13 7 13 10 9 2
17 0 3 9 13 10 9 9 3 13 7 13 10 9 1 9 13 2
20 3 1 0 10 3 9 13 7 13 10 10 9 9 13 1 10 9 10 9 2
12 13 3 3 9 3 13 10 9 10 13 9 2
4 13 10 9 2
3 9 13 2
4 13 3 9 2
24 3 7 13 10 1 10 9 13 7 15 13 16 13 3 10 0 13 9 15 3 13 0 13 2
23 3 3 3 0 0 13 13 1 9 10 9 10 0 13 9 1 10 9 1 9 10 9 2
13 10 3 0 13 9 13 10 9 9 15 13 13 2
12 10 3 13 10 3 9 13 15 7 9 13 2
23 13 3 10 9 15 7 13 10 0 9 0 13 3 13 10 9 1 0 1 10 9 13 2
13 13 3 10 9 1 9 13 13 7 13 10 9 2
5 3 3 3 13 2
10 9 3 1 10 9 15 13 7 13 2
17 3 3 9 9 1 9 13 10 9 13 10 9 10 9 3 13 2
12 10 3 3 9 15 13 13 7 13 10 9 2
7 13 3 3 0 0 0 2
8 9 3 0 9 1 15 13 2
14 3 3 10 9 3 13 13 0 3 10 10 9 9 2
13 3 1 10 3 10 9 10 9 0 0 9 13 2
16 3 3 3 7 3 13 13 10 9 10 9 13 7 13 15 2
13 0 3 3 15 0 13 9 1 10 9 0 13 2
11 13 3 3 9 13 13 7 10 0 9 2
11 3 3 10 0 9 1 0 13 10 9 2
8 10 3 13 13 7 3 13 2
18 10 3 13 10 9 1 10 9 9 10 9 9 13 13 1 9 13 2
10 10 3 9 0 13 13 13 10 9 2
17 13 3 3 10 9 0 9 3 10 9 13 7 10 0 9 13 2
10 9 3 3 3 13 3 10 9 13 2
21 3 3 3 3 1 10 13 13 0 9 0 3 3 13 10 9 10 9 9 13 2
16 9 3 9 13 9 16 9 3 13 13 3 13 9 10 9 2
20 0 3 13 13 10 9 13 15 10 1 10 9 1 10 9 7 10 9 13 2
12 3 10 3 9 3 0 13 13 1 10 9 2
20 3 3 16 15 1 10 9 9 13 2 13 0 15 3 0 9 9 7 0 2
14 15 3 13 15 0 13 2 16 13 0 3 13 15 2
13 9 3 13 0 13 7 3 1 15 13 0 13 2
39 3 9 3 10 9 2 10 0 9 13 2 16 3 13 10 9 2 1 9 13 10 9 15 10 1 10 10 0 9 2 13 3 13 15 16 0 0 9 2
18 15 3 13 3 10 10 9 9 1 10 0 13 9 1 9 13 9 2
14 13 3 10 9 2 15 7 13 10 9 2 0 13 2
19 3 15 13 3 10 0 15 9 10 1 10 9 7 10 9 9 3 13 2
20 3 0 13 15 9 9 3 9 3 9 9 3 9 7 9 2 7 9 0 2
11 3 9 3 1 9 1 15 13 13 13 2
9 10 3 9 13 3 9 13 13 2
28 3 9 0 13 13 10 9 3 10 9 13 10 0 15 1 10 0 13 9 2 7 10 0 13 13 1 15 2
19 0 3 3 13 10 9 13 1 10 9 2 15 13 1 9 1 9 13 2
20 3 10 9 0 13 1 10 0 9 13 7 13 9 7 9 13 15 9 0 2
12 13 3 1 10 9 2 16 13 15 13 13 2
5 3 13 0 9 2
26 13 3 0 0 2 16 3 3 9 13 0 13 9 0 3 13 9 15 9 13 2 0 13 2 9 2
5 10 3 9 13 2
17 15 3 13 10 9 9 0 2 7 10 9 10 9 7 10 9 2
18 3 1 3 10 9 2 13 1 10 1 9 9 2 3 3 0 13 2
6 3 3 13 16 15 2
32 10 3 3 0 7 3 0 13 2 3 9 13 7 10 9 13 2 10 7 9 13 1 9 3 1 9 7 1 10 15 9 2
7 9 3 1 10 9 13 2
6 9 3 3 0 0 2
38 16 3 9 2 3 1 10 9 10 1 10 0 2 15 3 0 13 13 2 3 10 13 9 13 1 9 2 16 16 9 10 9 9 3 10 0 13 2
19 3 3 3 10 10 13 1 9 7 9 7 0 9 7 9 0 3 13 2
11 9 3 10 0 1 10 1 9 15 13 2
26 10 9 7 10 9 10 0 13 9 7 0 13 9 10 9 13 2 0 13 10 9 10 10 9 9 2
19 0 3 10 10 9 13 7 13 13 0 7 0 13 2 16 9 7 9 2
20 3 3 10 15 9 10 9 15 7 10 9 13 2 0 7 0 10 0 13 2
7 13 3 10 9 7 13 2
7 10 3 13 9 7 0 2
15 3 10 9 9 2 16 13 2 0 3 13 7 0 13 9
26 0 3 3 13 9 2 0 3 13 9 2 9 7 13 10 9 0 9 1 10 9 7 10 9 13 2
14 9 3 15 9 13 10 9 2 16 3 13 16 13 2
18 3 15 13 10 10 1 9 13 9 7 0 10 10 9 0 9 13 2
25 3 10 0 3 2 13 2 7 0 9 1 9 13 0 0 10 9 13 13 2 9 3 3 13 2
11 0 3 9 1 0 9 0 7 0 9 2
7 15 1 3 9 0 9 2
9 3 13 2 13 2 9 1 9 2
7 3 3 0 9 0 9 2
24 3 9 3 10 9 7 10 13 9 13 13 0 2 16 9 3 9 13 2 3 7 13 9 2
21 3 3 9 13 10 1 9 7 9 9 0 1 9 13 16 9 13 7 9 13 2
22 15 1 9 0 10 1 9 9 13 2 0 3 9 13 2 1 0 7 3 9 13 2
10 13 3 3 15 1 10 3 15 13 2
22 15 3 2 13 2 10 0 9 13 1 9 9 0 13 2 9 13 3 9 7 9 2
33 3 9 3 10 9 2 0 13 9 2 16 3 0 10 9 13 2 16 13 10 9 2 3 0 15 13 10 9 2 7 10 0 2
14 0 3 10 9 13 10 9 2 3 3 10 9 13 2
11 9 3 10 9 0 13 13 13 10 0 2
17 10 3 1 10 9 9 9 13 13 9 10 0 9 2 15 13 2
9 15 15 15 0 1 9 13 13 2
25 10 3 9 13 10 9 13 10 9 1 10 13 0 10 9 13 10 0 15 13 2 13 10 9 2
19 3 3 15 9 3 9 9 3 9 3 9 3 0 9 3 0 7 9 2
9 3 3 3 13 15 13 3 13 2
9 15 13 3 10 13 9 10 9 2
9 10 13 3 13 0 3 0 13 2
7 3 13 3 9 1 9 2
5 9 9 13 0 2
22 13 3 15 13 0 13 10 9 10 9 2 13 10 0 9 3 10 1 9 2 13 2
26 10 3 9 1 9 13 13 0 1 9 2 1 3 15 9 9 9 13 2 10 7 0 9 13 15 2
8 3 10 9 3 1 15 13 2
10 3 3 15 15 13 13 3 13 7 2
9 13 13 9 3 0 7 9 0 2
14 3 3 9 9 7 9 9 10 9 1 10 9 13 2
24 0 3 1 9 13 0 0 9 9 2 15 3 10 9 13 3 1 9 2 13 7 1 9 2
14 13 3 10 9 13 9 7 9 1 10 9 10 9 2
14 1 9 3 13 9 7 1 9 10 13 10 9 9 2
20 3 10 9 3 15 13 10 9 10 10 9 9 3 0 13 10 10 9 9 2
14 13 3 2 16 13 9 2 1 9 7 10 13 9 2
10 0 3 13 10 9 7 0 10 9 2
37 16 3 3 1 10 9 13 2 13 2 9 2 3 13 0 13 1 10 9 10 9 7 1 9 13 2 7 3 15 0 9 13 7 15 13 13 2
8 3 10 9 0 1 15 13 2
16 13 3 15 3 0 9 2 16 13 10 0 9 1 0 0 2
20 15 3 10 3 0 13 16 9 13 2 10 7 9 13 7 13 13 9 13 2
19 3 13 1 10 15 9 0 13 9 0 2 1 15 15 15 13 16 9 2
19 16 3 1 10 0 9 13 2 13 1 10 9 2 3 7 3 1 9 2
8 0 3 3 13 1 10 9 2
12 16 3 1 9 13 2 3 10 9 15 13 2
24 10 3 9 1 15 13 13 0 13 2 15 13 9 9 0 0 2 1 15 13 9 0 0 2
24 13 3 2 16 13 2 10 0 3 7 0 15 1 10 9 9 3 10 10 9 13 9 13 2
5 3 13 3 13 2
28 10 3 13 15 15 0 9 13 9 10 13 3 0 13 15 9 13 2 0 7 3 15 13 15 2 9 13 2
48 9 3 10 0 1 10 0 10 1 9 9 1 15 2 13 2 13 9 10 10 9 9 16 13 10 0 9 1 9 9 0 0 2 1 15 9 0 1 0 13 9 2 7 15 13 9 0 2
18 3 1 9 0 9 0 2 3 9 0 13 9 2 7 13 0 9 2
13 13 3 1 10 9 3 0 9 0 1 10 9 2
18 10 3 9 15 9 13 1 10 9 3 9 13 1 10 0 9 13 2
15 9 3 1 0 1 9 1 9 13 13 3 0 13 9 2
11 10 3 15 16 15 13 2 9 10 9 2
22 9 3 1 0 9 13 2 13 2 3 3 10 1 9 9 7 10 9 9 7 9 2
17 3 3 10 3 1 9 9 13 13 2 10 7 10 9 9 13 2
8 13 3 13 3 10 9 15 2
34 15 3 0 3 3 10 9 0 13 3 13 2 7 3 3 10 9 10 9 1 9 13 2 16 3 13 10 9 2 7 13 10 9 2
7 3 3 9 0 15 13 2
28 3 3 1 10 9 3 0 9 3 9 7 9 15 13 13 2 7 3 1 0 10 9 9 0 7 9 13 2
28 1 3 3 10 9 3 13 15 3 10 10 9 7 10 10 9 9 2 7 1 15 0 9 9 13 15 13 2
9 1 10 3 3 13 1 15 3 2
13 3 3 9 0 13 1 10 9 16 1 10 9 2
11 3 3 10 9 3 16 10 3 13 13 2
33 9 3 1 10 0 1 9 9 2 13 2 1 9 9 13 7 0 15 13 13 2 0 13 10 3 3 15 13 10 10 9 9 2
22 3 3 13 9 10 10 15 9 7 9 1 10 9 10 1 10 9 9 13 13 13 2
9 15 0 13 10 1 9 13 9 2
10 10 3 1 9 13 13 9 13 9 2
29 13 3 3 15 0 7 13 10 13 15 0 9 10 1 10 9 9 10 10 9 9 13 1 0 9 1 15 13 2
12 1 15 3 13 1 9 13 10 9 10 9 2
14 3 10 9 10 0 10 9 13 10 9 13 0 9 2
42 3 0 3 9 9 0 13 10 13 2 7 3 9 10 0 2 3 3 10 1 9 7 0 3 10 9 10 15 9 13 2 0 15 9 13 13 1 9 9 7 9 2
6 15 3 13 13 0 2
13 3 9 3 15 13 10 9 2 3 9 7 0 2
6 3 13 1 10 9 2
22 13 3 15 13 10 0 9 1 0 9 3 0 9 3 0 9 9 3 7 9 0 2
9 13 3 15 9 1 9 7 9 2
6 9 3 13 10 13 2
7 3 13 9 7 13 3 2
4 0 0 9 2
15 3 0 3 15 16 13 15 2 13 10 9 15 3 13 2
4 9 3 13 2
13 10 15 3 3 3 9 13 2 9 7 9 13 2
14 0 13 15 2 10 0 3 9 13 3 9 7 9 2
5 0 13 10 9 2
9 13 10 9 3 9 1 13 3 2
18 10 1 10 9 9 13 3 16 0 9 13 2 9 2 9 1 0 2
9 15 3 15 9 13 7 9 0 2
12 15 0 13 9 3 13 2 9 7 7 9 2
18 3 1 10 9 3 13 10 9 13 1 9 7 9 2 16 13 9 2
15 3 9 3 1 9 13 1 10 9 2 16 9 1 9 2
31 9 3 10 0 10 10 0 13 1 10 13 0 13 16 10 1 10 0 9 9 0 3 13 7 15 0 2 13 3 15 2
8 15 3 13 10 9 7 9 2
28 13 3 3 3 1 10 9 1 9 7 9 10 9 13 7 13 3 9 9 15 7 0 13 2 7 9 13 2
21 3 16 15 15 13 3 3 13 2 13 9 1 10 0 10 9 7 15 9 13 2
23 10 3 13 3 13 13 10 9 7 13 10 9 2 7 10 9 16 13 13 7 15 13 2
10 3 16 13 10 9 3 13 2 13 2
21 10 3 9 13 10 9 1 10 9 3 10 1 15 9 7 9 13 9 0 0 2
18 1 3 9 3 13 13 9 1 10 0 16 10 9 0 10 9 13 2
20 9 3 1 10 0 0 10 9 3 9 13 13 1 10 9 0 13 10 9 2
24 13 3 15 3 1 10 9 10 15 2 7 1 15 16 13 10 13 2 7 13 15 16 13 2
20 13 3 3 15 10 15 9 10 13 2 9 10 0 13 7 13 10 9 0 2
19 15 3 0 13 9 3 0 15 1 10 0 15 13 2 7 3 13 13 2
8 0 3 3 15 1 15 13 2
33 3 15 13 0 13 16 3 13 2 16 10 3 9 10 9 13 2 13 7 15 15 2 16 13 10 7 10 2 13 3 10 9 2
12 16 3 13 1 9 7 1 9 2 13 3 2
33 0 3 16 13 13 7 13 13 2 13 1 15 10 9 10 9 3 13 3 3 9 2 3 3 9 3 0 2 3 7 3 9 2
20 3 13 3 3 3 10 9 2 0 7 3 3 13 13 10 9 7 10 9 2
18 3 3 13 1 15 3 0 10 9 2 3 3 13 7 13 10 9 2
13 0 3 10 1 9 13 9 13 7 13 10 9 2
21 3 1 3 10 9 9 13 0 7 9 15 10 9 13 2 16 1 15 10 9 2
18 1 15 16 13 2 13 15 0 9 2 15 13 10 13 7 10 13 2
20 13 3 15 10 9 0 3 10 9 10 10 9 13 2 13 1 9 7 9 2
20 1 3 10 9 10 9 2 16 9 13 2 1 9 3 13 3 13 7 13 2
35 0 3 13 1 9 3 10 10 9 9 2 15 7 10 1 15 9 13 13 0 2 13 10 1 15 13 9 2 16 13 9 1 0 9 2
8 1 3 9 15 13 3 13 2
24 1 15 0 13 1 10 9 9 7 9 13 2 10 3 0 13 7 16 3 13 13 10 13 2
10 3 13 3 3 9 1 10 9 13 2
21 13 3 1 15 9 16 9 9 1 9 3 13 13 13 10 9 13 15 9 13 2
28 1 9 3 13 15 10 10 13 9 13 15 9 13 13 2 16 15 13 9 9 3 13 10 13 15 10 9 2
40 15 3 9 13 1 9 7 13 1 9 2 1 10 9 13 7 13 1 15 2 0 3 13 13 10 10 9 13 9 2 3 7 13 13 15 10 15 15 13 2
20 9 3 1 15 3 10 9 1 10 10 9 9 9 3 13 7 9 13 13 2
24 1 15 7 10 0 15 9 10 10 9 9 13 2 16 13 9 1 0 9 2 13 13 9 2
9 3 0 15 15 13 1 0 9 2
10 1 15 13 1 10 13 2 13 15 2
12 10 3 15 13 3 9 10 0 1 9 3 2
29 3 3 0 0 2 13 2 13 9 13 9 2 16 13 9 2 16 9 13 7 13 3 9 7 9 2 0 0 2
32 3 9 3 1 10 1 9 7 9 9 13 10 0 0 3 7 9 13 0 9 13 3 15 1 10 9 13 1 10 9 13 2
12 3 10 9 13 10 9 9 7 9 3 9 2
10 13 3 10 9 3 9 0 9 13 2
17 13 3 10 3 1 9 9 2 10 7 3 10 9 16 9 13 2
21 10 3 0 15 16 1 9 13 2 3 1 9 13 10 0 9 1 0 9 13 2
13 13 3 15 15 3 10 1 10 9 13 9 0 2
36 10 3 0 15 13 9 3 10 9 2 1 15 1 9 10 9 1 10 9 13 10 3 1 10 9 13 2 10 7 1 10 9 10 9 13 2
37 13 3 3 3 0 7 0 9 3 10 3 13 0 9 13 7 15 13 1 10 0 9 7 10 9 2 13 3 9 2 7 10 1 10 9 9 2
11 1 9 3 13 3 9 1 15 13 13 2
12 0 3 3 9 13 2 15 13 1 10 9 2
18 13 3 10 13 1 10 9 15 13 1 10 13 1 10 10 9 9 2
48 13 3 0 10 9 0 13 16 1 10 9 2 0 10 9 13 7 10 9 3 0 1 10 9 13 2 10 3 10 9 9 7 10 1 10 9 9 13 0 13 7 13 13 1 10 9 3 2
27 10 3 9 15 1 0 13 10 3 9 3 3 7 1 9 9 13 13 2 10 7 0 10 9 9 0 2
19 13 3 3 3 1 9 10 13 2 15 13 9 9 2 13 1 15 13 2
5 3 10 9 13 2
18 16 3 3 0 0 9 9 13 2 3 15 9 3 7 0 9 13 2
12 15 13 13 13 15 10 9 16 3 13 13 2
21 13 3 15 10 9 10 9 16 15 10 9 15 13 15 13 1 10 0 3 13 2
15 16 3 10 0 13 1 10 10 9 15 9 2 13 13 2
19 13 3 13 1 15 9 2 3 10 9 7 1 0 10 15 13 1 9 2
19 3 3 3 0 13 15 9 0 10 9 2 1 15 3 13 13 2 13 2
18 1 15 3 13 9 13 16 3 1 10 9 10 9 13 1 9 13 2
25 15 3 13 10 9 16 15 13 2 16 3 9 13 1 10 9 15 2 13 10 9 10 0 9 2
9 13 3 15 3 9 1 0 9 2
20 3 3 13 13 10 9 3 0 13 2 7 3 10 9 13 13 1 10 9 2
15 10 0 13 3 1 9 10 0 9 1 0 9 13 3 2
7 9 1 9 13 7 13 2
8 9 3 10 9 13 10 9 2
15 15 3 9 13 1 10 9 13 7 0 9 13 9 13 2
20 9 3 9 13 16 9 13 1 15 2 7 0 1 15 13 1 10 9 13 2
20 3 13 1 10 9 1 10 9 10 9 13 1 10 9 13 9 1 10 9 2
30 10 3 9 0 10 9 13 1 10 9 13 1 10 9 2 7 1 10 0 9 13 10 0 16 13 13 13 10 9 2
22 15 3 13 10 9 13 1 10 9 9 2 7 13 10 9 1 10 9 13 0 9 2
17 3 16 10 9 13 2 13 13 10 9 0 10 9 10 9 13 2
14 10 3 9 10 9 1 10 9 13 2 7 3 13 2
29 9 3 15 1 9 3 13 13 1 10 9 0 13 9 2 1 15 3 13 7 13 0 7 1 15 10 9 13 2
14 10 3 3 13 13 3 10 9 7 13 10 9 13 2
19 3 15 10 13 13 13 15 2 13 16 13 10 9 16 1 10 9 13 2
21 10 3 13 16 3 3 15 13 16 1 10 9 13 13 7 3 1 10 9 13 2
47 9 2 13 2 13 1 9 13 9 10 9 1 10 9 13 7 10 1 10 9 13 1 9 10 9 13 2 16 3 13 10 9 10 9 10 3 9 7 10 0 9 13 3 1 10 9 2
29 3 3 3 10 10 9 13 9 13 7 10 13 2 10 0 9 3 10 10 9 10 0 13 7 10 13 0 13 2
27 3 3 13 1 9 10 0 1 9 9 13 0 15 13 7 1 10 9 10 9 13 7 1 9 13 13 2
12 15 3 15 3 10 9 13 9 13 10 9 2
18 13 3 1 0 9 0 15 10 9 10 15 13 9 1 10 15 9 2
10 13 3 3 9 9 1 10 9 15 2
12 3 3 3 13 10 9 16 0 1 9 13 2
10 9 3 10 0 1 10 1 9 13 2
34 3 1 10 9 15 13 3 10 10 9 9 2 10 7 9 13 9 9 2 16 10 3 0 9 13 9 2 13 13 10 10 9 9 2
18 3 0 13 7 13 0 2 10 3 10 10 9 10 3 9 13 13 2
16 3 9 3 2 16 13 9 2 1 10 13 9 13 1 9 2
15 10 3 3 1 9 13 15 13 2 7 1 9 10 9 2
30 15 10 3 9 13 9 2 9 7 10 9 9 13 7 1 10 15 9 13 1 9 13 1 9 2 9 10 9 13 2
6 3 13 13 1 9 2
15 1 15 3 0 13 9 13 10 0 10 9 1 10 9 2
25 0 3 3 10 9 2 13 10 9 2 13 10 0 9 13 2 10 0 9 13 0 3 0 9 2
7 10 3 9 15 13 13 2
28 9 3 13 9 1 0 9 9 7 9 13 1 15 9 13 16 10 0 9 13 7 10 9 0 10 0 13 2
18 13 3 2 13 2 3 9 0 0 2 15 3 10 10 9 13 9 2
14 3 3 10 9 13 16 9 10 1 9 13 13 0 2
22 3 3 3 3 1 9 0 10 9 0 13 10 1 9 13 0 13 9 1 10 9 2
21 1 15 1 0 13 9 3 13 10 13 7 10 0 13 9 2 7 13 9 9 2
56 9 3 3 10 9 1 9 13 1 9 9 13 7 13 2 10 1 15 9 13 10 9 1 10 9 9 1 15 9 2 3 0 9 13 16 0 10 9 13 7 9 0 13 9 3 0 13 2 10 7 13 7 13 0 13 2
12 3 1 9 13 9 7 9 15 13 10 9 2
11 0 3 13 3 3 13 10 1 9 9 2
23 3 0 10 1 15 3 3 1 9 13 7 0 9 13 13 2 0 10 3 13 0 13 2
21 9 3 3 1 0 9 7 0 13 7 9 0 13 15 13 10 1 10 9 9 2
12 9 3 13 10 10 15 9 10 9 13 9 2
13 13 3 1 10 1 10 9 9 2 1 9 13 2
32 3 10 10 9 3 13 2 15 0 13 10 1 9 13 2 0 3 9 2 16 13 9 7 9 2 1 9 13 3 0 9 2
31 3 3 3 1 15 13 13 0 9 2 15 13 9 0 2 7 13 1 15 1 10 0 9 2 16 9 10 0 9 13 2
14 3 9 3 10 9 13 10 9 10 9 1 10 9 2
15 3 3 15 0 9 3 0 7 0 2 0 1 9 9 2
20 13 3 10 9 2 16 3 9 13 7 9 1 9 9 2 1 9 0 9 2
13 3 3 0 9 13 0 3 10 1 10 9 9 2
36 9 3 16 3 3 13 2 13 9 2 16 13 9 2 7 10 3 1 9 9 13 7 10 0 9 13 9 0 2 7 0 1 10 9 13 2
10 9 3 10 0 1 0 1 9 13 2
12 10 9 9 13 9 1 9 9 7 0 9 2
11 10 10 0 3 13 1 9 13 10 0 2
14 3 3 10 0 13 0 15 9 13 1 10 9 13 2
14 15 13 13 15 3 0 13 9 7 9 0 0 13 2
18 3 10 9 1 0 9 13 15 10 9 7 13 1 0 9 13 13 2
15 3 15 9 3 9 13 0 0 3 9 7 9 3 0 2
22 9 3 1 0 9 13 13 10 9 10 9 9 13 3 10 0 2 3 13 13 15 2
10 3 10 0 0 7 3 1 10 0 2
10 3 1 9 3 3 10 9 15 13 2
10 0 3 9 0 0 9 13 10 9 2
10 3 3 13 0 0 9 1 10 9 2
19 13 3 3 16 15 0 2 10 0 9 3 9 7 10 0 15 9 13 2
29 13 3 3 3 3 7 0 0 10 9 1 10 13 13 1 15 13 9 16 0 10 9 1 15 13 13 10 9 2
14 15 10 0 13 3 7 3 1 10 9 13 10 9 2
21 10 3 9 15 10 9 10 1 9 7 9 0 9 13 10 9 2 9 9 13 2
37 3 0 9 0 10 13 10 9 9 3 13 10 9 13 10 0 10 9 2 16 10 10 9 7 10 9 1 15 9 1 9 13 9 9 9 13 2
25 0 3 3 3 13 16 15 0 10 10 9 9 13 13 1 10 13 10 1 9 9 0 15 13 2
35 1 10 9 3 10 13 15 9 2 16 1 10 9 3 10 3 10 9 9 7 10 9 13 2 0 9 10 3 10 1 9 9 13 13 2
12 10 3 0 9 13 9 7 9 1 9 13 2
16 10 3 1 9 3 13 1 9 2 9 3 0 13 3 9 2
35 3 0 13 0 9 13 7 13 13 2 16 13 10 9 13 1 9 2 0 3 16 1 9 2 0 3 16 1 9 2 10 7 1 9 2
5 13 3 0 7 2
55 16 13 1 10 0 2 13 1 15 10 15 9 13 13 1 9 2 3 9 0 15 13 0 7 9 15 1 2 7 10 15 9 7 9 10 9 0 9 9 13 1 10 1 9 9 2 16 1 10 0 9 13 13 15 2
22 13 3 3 9 10 1 10 9 1 10 0 13 2 16 13 9 1 10 0 7 9 2
5 13 3 1 9 2
31 3 1 0 3 10 9 9 10 0 1 10 0 1 10 1 9 9 13 1 10 9 15 7 15 13 0 9 13 3 15 2
12 10 3 10 9 0 3 0 7 0 9 0 2
8 10 3 9 1 0 13 9 2
15 13 3 10 3 0 15 2 10 3 0 2 10 7 0 2
9 13 3 3 15 3 0 7 0 2
11 13 3 3 0 9 2 15 13 0 0 2
21 13 3 3 15 2 13 2 3 10 13 0 2 15 13 3 0 1 10 0 9 2
15 10 3 9 9 0 0 1 10 3 9 9 13 1 0 2
10 15 0 13 13 10 0 13 1 9 2
9 13 3 10 10 9 9 3 13 2
22 10 3 3 13 16 9 13 1 9 9 2 13 9 0 2 0 9 9 9 0 13 2
24 9 3 10 0 1 10 1 9 9 13 1 9 13 1 10 1 15 9 16 9 10 9 13 2
38 9 3 2 16 13 9 2 10 9 13 0 1 10 9 2 16 1 9 13 1 9 9 7 9 13 2 13 13 10 9 0 9 2 16 3 9 13 2
18 3 3 13 1 10 0 9 16 15 15 3 13 10 9 7 13 13 2
11 1 3 15 10 0 9 13 1 10 13 2
14 9 3 1 0 9 0 13 9 15 0 13 9 13 2
10 15 3 3 9 0 3 13 7 0 2
14 3 1 10 0 9 1 9 7 9 13 0 9 13 2
14 15 13 1 15 3 9 10 0 1 10 0 10 9 2
12 0 3 1 0 9 9 9 1 9 15 13 2
12 3 9 2 7 15 9 0 0 0 9 13 2
18 9 3 1 10 1 9 7 3 3 10 9 13 1 10 9 10 9 2
7 3 3 3 10 0 9 13
13 3 10 9 3 15 13 9 1 0 9 0 13 2
11 1 3 9 7 9 10 15 13 9 15 2
39 13 3 10 9 3 1 10 13 0 3 9 3 10 9 1 9 13 13 7 10 9 0 1 10 9 7 10 9 13 0 7 13 7 13 13 1 10 9 2
43 9 3 16 3 13 15 10 9 0 1 9 7 9 0 13 13 2 16 7 10 9 10 9 13 2 13 1 9 2 3 10 1 9 9 1 0 7 0 9 7 0 13 2
50 1 3 9 13 1 10 0 13 16 13 10 3 1 10 9 7 10 9 13 2 10 7 1 9 3 9 7 10 15 9 13 2 7 3 13 16 9 0 10 9 13 0 3 10 15 9 16 13 13 2
12 9 3 0 2 13 2 9 13 0 7 0 2
22 13 3 10 9 2 16 3 9 13 2 0 9 0 13 1 3 10 9 7 10 9 2
18 15 15 0 13 1 10 9 13 10 9 2 13 10 15 9 7 9 2
23 1 3 9 9 3 1 0 9 13 16 1 10 10 9 9 7 10 10 9 9 0 13 2
25 9 3 1 0 9 9 2 13 2 15 10 0 0 13 1 9 0 3 13 3 0 13 10 15 2
17 0 3 13 1 9 9 3 7 9 2 16 3 9 13 1 9 2
26 3 3 3 13 15 15 13 2 7 3 13 2 7 13 3 2 0 9 0 15 9 7 0 1 9 2
7 9 3 1 10 9 13 2
15 15 3 10 9 13 1 9 3 7 9 13 16 0 13 2
29 1 3 15 10 9 3 3 0 15 3 13 10 1 10 9 9 1 0 13 13 2 0 7 3 3 13 3 13 2
7 1 0 3 9 13 3 2
20 13 3 3 0 9 0 13 9 13 3 9 13 7 0 9 10 13 13 9 2
17 9 3 0 9 1 10 1 10 9 9 13 16 13 13 3 15 2
18 1 3 10 0 9 13 0 13 9 1 10 1 9 7 9 13 13 2
14 3 13 3 2 13 2 13 10 13 9 13 10 9 2
6 3 1 9 0 13 2
6 3 13 9 9 13 2
36 3 9 3 10 1 9 2 16 13 9 7 10 13 10 1 15 13 0 2 13 13 3 0 9 13 7 1 9 1 10 9 13 1 9 13 2
10 1 3 3 9 7 9 9 15 13 2
8 1 3 10 1 9 15 13 2
17 15 3 13 3 9 2 15 10 3 9 13 9 2 10 7 9 2
20 10 3 0 2 15 13 3 9 2 13 1 15 13 16 15 15 13 13 13 2
44 9 3 13 1 9 15 13 3 13 0 9 7 13 1 10 9 13 15 13 1 10 0 2 9 13 9 0 9 2 1 15 13 0 9 0 7 0 7 0 9 7 0 0 2
29 13 3 1 10 9 3 9 0 1 9 3 9 13 7 13 15 3 1 3 10 9 7 10 9 1 10 0 9 2
25 10 3 0 9 7 0 9 13 10 9 13 13 1 9 1 10 3 9 2 13 15 0 0 9 2
24 13 3 10 9 9 0 3 7 0 2 7 1 9 13 0 9 7 0 2 16 3 13 9 2
11 3 13 13 10 9 2 7 13 0 9 2
12 10 3 13 13 10 9 7 13 15 9 13 2
7 15 3 0 13 10 9 2
11 10 3 3 9 3 13 16 13 3 13 2
47 3 10 0 0 9 2 10 1 0 10 9 13 10 9 2 7 13 13 1 10 10 9 9 10 9 13 0 9 13 0 10 10 9 9 2 3 0 13 9 9 15 13 13 3 1 9 2
7 13 3 3 0 13 9 2
7 3 3 13 15 10 9 2
13 9 9 9 13 7 9 0 9 2 7 3 13 2
8 3 15 9 0 13 15 13 2
19 9 3 1 10 0 10 1 9 9 13 13 9 1 10 9 10 9 9 2
18 9 3 1 9 2 15 13 2 13 2 9 2 9 13 1 9 13 2
25 3 13 3 3 10 10 9 9 2 1 15 13 9 0 13 10 0 9 10 9 2 3 3 13 2
10 9 9 9 9 7 9 13 9 0 2
6 13 2 13 2 13 2
10 16 15 15 3 0 10 9 13 13 2
18 3 3 15 13 0 9 7 9 0 13 2 16 9 13 1 0 9 2
36 9 3 1 0 9 9 13 10 0 1 9 13 3 1 9 1 10 10 9 9 2 16 3 13 13 2 3 3 7 10 9 3 10 9 13 2
17 3 3 9 9 10 0 13 16 13 3 13 10 9 10 9 13 2
10 9 3 0 2 9 7 13 9 0 2
35 9 3 13 9 10 9 9 7 10 9 13 9 13 0 7 9 2 7 16 9 9 13 15 1 10 9 13 12 7 12 13 7 13 9 2
15 9 3 10 0 9 1 9 13 1 10 0 10 9 13 2
11 9 9 0 13 2 16 15 13 2 0 2
11 15 13 9 9 2 9 0 0 0 9 2
22 15 3 13 9 3 13 13 7 1 9 9 0 13 2 16 9 2 9 10 9 13 2
31 3 9 2 3 9 15 2 7 13 13 2 7 13 2 7 13 0 13 3 7 13 13 2 10 7 15 0 1 9 13 2
18 13 2 3 9 7 7 9 13 3 9 7 1 10 3 9 9 9 2
5 3 3 3 13 2
9 13 3 0 13 0 13 0 13 2
14 15 3 1 9 3 9 3 9 7 0 9 13 13 2
7 9 3 0 10 0 13 2
18 9 3 1 0 0 9 9 13 10 0 9 13 9 7 9 0 9 2
25 0 3 10 9 9 13 13 13 3 13 7 9 7 9 13 2 15 3 10 9 13 13 0 9 2
40 3 15 3 15 13 1 10 9 0 10 3 9 2 16 13 9 2 1 10 0 9 7 9 13 10 9 2 10 7 9 1 9 3 9 7 9 13 10 9 2
17 13 3 3 13 1 15 7 13 0 0 0 7 0 13 10 9 2
36 10 3 13 1 0 9 2 16 15 13 2 16 13 1 10 13 10 3 9 10 9 7 10 9 10 9 10 1 0 13 13 13 10 15 15 2
8 13 3 13 0 13 7 0 2
16 3 3 1 3 10 10 9 9 13 2 7 0 0 9 13 2
12 1 3 10 0 10 0 9 1 9 13 13 2
41 13 3 3 10 1 9 13 2 15 0 10 9 10 1 10 9 13 3 1 9 7 9 13 2 7 13 10 9 3 13 9 9 0 7 0 9 2 15 13 9 2
30 3 13 1 0 3 13 9 3 10 9 13 7 13 1 10 9 2 0 7 0 13 16 1 10 9 13 7 13 13 2
23 13 3 3 10 9 16 9 13 10 9 3 13 15 10 9 7 9 13 13 13 10 9 2
17 3 3 0 13 13 15 10 0 13 16 13 10 9 1 10 9 2
33 13 3 15 7 13 15 13 1 10 9 2 13 15 13 7 15 0 1 10 15 2 7 10 0 13 13 13 3 10 9 15 13 2
21 10 3 9 0 3 3 13 10 15 9 10 15 9 13 10 9 1 10 9 13 2
13 1 3 10 0 10 0 1 9 10 0 13 13 2
5 0 3 13 0 2
11 3 1 10 9 1 10 0 7 0 13 2
45 15 3 13 13 9 3 9 7 0 9 2 7 10 9 10 13 1 10 9 10 3 1 15 10 9 13 2 10 7 15 13 3 10 3 13 3 10 9 13 7 10 9 10 13 2
23 1 15 10 9 10 10 9 3 13 2 7 1 15 3 3 15 13 10 9 2 7 3 2
54 3 3 15 15 10 9 13 2 16 10 3 9 1 10 9 7 1 10 9 13 2 10 3 0 15 0 1 9 3 9 7 10 15 9 2 10 7 9 0 0 13 1 10 0 9 7 9 16 1 10 10 9 9 2
24 1 3 10 13 10 9 9 1 10 1 9 13 9 9 2 13 2 10 0 1 9 9 12 2
18 1 15 13 9 1 10 9 13 10 0 10 13 9 1 10 9 9 2
8 15 13 3 9 10 9 13 2
11 1 15 3 9 10 10 9 9 13 3 2
11 9 10 10 9 13 3 13 7 13 13 2
6 3 3 13 3 9 2
9 9 13 3 0 13 9 9 3 2
4 3 0 13 2
6 10 15 13 3 9 2
14 9 3 13 3 10 9 9 7 9 13 9 7 9 2
10 3 10 9 15 9 3 13 10 9 2
32 3 3 1 10 9 7 1 10 9 9 13 2 16 9 13 1 10 0 7 0 2 7 13 10 13 13 13 7 13 15 13 2
8 15 0 13 3 9 13 15 2
14 1 15 3 3 13 1 10 0 10 0 10 9 13 2
32 9 10 0 1 10 9 7 10 9 0 10 9 13 9 2 16 10 13 10 9 13 13 7 13 16 15 13 10 1 10 9 2
7 3 10 9 13 0 0 2
34 13 3 3 10 1 0 9 15 15 13 2 7 13 16 13 3 3 9 0 7 0 13 9 15 7 13 13 2 16 15 13 15 13 2
11 1 3 15 0 13 7 0 13 10 9 2
21 10 3 9 3 1 0 0 13 2 16 3 10 3 10 9 9 15 15 13 9 2
43 9 3 10 0 13 9 10 0 1 10 1 9 16 13 1 10 9 10 9 7 10 1 9 9 13 13 3 1 9 10 1 9 9 7 10 0 9 10 9 1 15 13 2
19 9 3 3 9 13 7 9 13 3 0 13 9 1 10 9 13 0 13 2
32 9 3 1 0 0 10 9 13 1 9 10 0 9 13 13 9 3 10 9 0 13 7 9 9 13 3 10 9 9 3 13 2
13 3 3 9 15 1 9 1 9 13 13 1 15 2
12 10 3 15 9 13 7 0 13 15 0 0 2
23 0 3 13 10 9 9 3 13 1 0 10 9 7 9 13 13 2 15 1 15 9 13 2
23 7 3 13 13 1 9 13 1 10 9 2 13 3 0 1 10 9 7 3 1 10 9 2
28 3 3 9 10 0 3 3 15 9 13 10 9 0 15 3 0 3 0 3 0 7 0 1 9 0 13 13 2
15 1 3 10 9 16 13 2 0 10 0 9 16 9 13 2
40 9 3 3 15 0 13 0 2 9 3 10 9 15 0 13 2 9 3 13 1 10 9 7 9 0 2 0 7 9 13 7 10 15 10 1 10 1 9 9 2
29 15 10 3 13 9 7 9 13 15 2 1 3 0 9 13 13 7 1 10 9 15 9 2 0 13 10 0 9 2
8 3 13 3 3 0 13 13 2
17 9 3 13 1 9 7 9 13 2 1 15 13 9 9 9 13 2
7 3 3 13 10 9 13 2
9 13 3 9 0 13 10 0 13 2
11 9 3 10 9 1 10 9 15 13 13 2
13 3 15 13 9 2 15 3 13 13 13 0 13 2
23 16 3 13 9 0 2 13 3 15 2 7 16 3 13 7 13 9 2 9 13 13 9 2
13 13 3 3 1 9 16 0 1 9 1 9 3 2
6 9 1 10 9 13 2
3 15 13 2
8 3 3 13 10 15 13 9 2
5 3 9 3 13 2
16 3 13 9 3 9 2 16 13 2 9 0 10 9 13 3 2
12 1 9 3 13 13 10 9 10 9 9 9 2
31 13 3 15 15 3 9 1 13 13 2 7 16 10 13 1 15 13 3 10 9 7 3 13 10 9 1 9 7 1 9 2
17 13 3 13 15 10 3 9 10 0 9 9 7 9 10 0 9 2
17 10 3 9 1 15 15 13 1 3 10 9 10 9 13 0 9 2
33 16 3 3 13 7 10 9 13 10 9 2 9 3 13 10 0 13 10 0 9 2 9 7 10 9 13 10 1 10 9 9 13 2
6 3 3 3 13 15 2
13 3 3 0 9 13 10 9 7 3 0 9 9 2
23 13 3 9 10 9 9 7 13 9 10 0 13 9 7 10 0 13 9 2 3 3 9 2
27 9 3 1 10 0 7 0 10 9 9 3 2 13 2 10 10 9 9 13 10 0 9 10 0 13 9 2
16 10 3 9 9 9 9 7 0 9 2 3 7 9 13 0 2
10 9 3 16 10 9 13 0 13 9 2
5 9 3 0 13 2
11 10 3 3 9 15 13 13 1 0 9 2
16 13 3 1 3 10 9 10 9 3 9 9 13 10 0 9 2
13 15 3 9 0 13 9 3 7 3 13 10 9 2
24 10 3 9 15 13 0 13 10 9 10 9 2 10 7 0 13 0 9 13 7 10 0 9 2
21 9 3 0 13 2 10 9 0 13 13 2 1 10 9 13 10 0 9 10 9 2
14 13 3 10 9 3 13 1 10 9 1 10 9 13 2
71 9 3 10 0 1 0 10 1 10 9 9 2 13 2 10 1 9 13 9 2 10 10 9 13 0 7 1 9 13 1 9 13 10 0 9 10 13 10 9 10 1 10 9 13 2 15 3 3 3 13 13 2 13 13 2 3 15 13 2 0 10 9 2 1 10 9 7 9 13 15 2
14 13 3 3 9 10 0 2 16 9 1 10 0 13 2
18 1 3 10 0 13 16 9 10 9 13 10 0 9 13 3 7 3 2
16 3 3 13 10 3 9 13 2 7 13 3 1 9 3 13 2
10 3 0 13 1 9 13 13 15 0 2
25 3 13 7 1 10 9 13 3 9 13 2 3 9 0 9 13 10 0 1 10 13 15 10 9 2
23 9 3 1 10 0 10 9 0 13 10 13 9 9 13 9 2 9 0 10 1 15 13 2
7 13 3 3 0 7 0 2
35 13 3 1 9 0 9 2 16 3 3 13 7 13 1 0 9 10 0 1 10 9 13 3 10 13 13 1 7 10 9 3 13 2 13 2
12 1 3 9 7 10 15 9 13 3 0 13 2
18 3 16 3 9 10 0 1 10 1 9 13 1 15 2 3 13 13 2
25 16 10 0 1 9 13 10 9 2 3 2 16 13 2 9 9 9 9 13 10 10 9 9 2 2
18 13 3 1 10 9 10 15 13 7 10 9 1 9 0 13 10 9 2
10 13 3 0 13 13 10 9 10 9 2
25 16 3 3 10 10 9 9 13 1 10 9 9 2 13 0 13 10 9 2 3 13 15 9 13 2
36 10 3 13 10 10 9 9 1 9 10 9 10 9 13 13 10 9 1 10 9 2 7 13 1 10 9 0 10 0 13 15 10 9 0 13 2
34 3 9 10 1 15 13 10 10 9 13 13 9 3 1 9 9 16 13 10 9 3 13 2 13 3 3 0 1 0 9 0 9 13 2
4 3 13 0 2
7 13 3 1 10 0 13 2
15 10 3 9 2 13 2 10 3 9 7 10 9 15 13 2
40 1 3 10 9 10 3 9 9 3 10 0 1 10 1 10 9 7 9 9 13 16 1 10 9 13 15 0 9 7 9 0 2 1 15 13 13 1 10 9 2
41 9 3 13 16 1 10 9 0 10 9 13 13 10 9 7 16 1 10 0 9 0 10 9 0 15 13 1 10 9 9 13 7 10 0 3 13 3 10 15 13 2
39 15 3 0 16 3 1 15 9 10 9 1 10 9 13 13 10 0 9 13 15 9 7 9 13 13 2 9 10 0 15 15 13 9 2 7 3 10 9 2
13 13 3 10 9 3 9 0 7 9 0 10 9 2
9 13 3 15 9 7 10 0 9 2
11 9 3 7 9 13 0 1 9 10 13 2
6 0 3 13 7 0 2
5 13 3 13 0 2
20 13 3 0 1 10 9 2 13 10 9 2 9 13 0 7 10 0 9 0 2
35 9 3 1 10 0 10 1 9 9 16 2 13 2 13 9 2 9 13 15 3 7 10 0 0 2 0 7 0 9 13 1 10 0 9 2
18 13 3 10 9 0 2 1 15 0 13 9 13 9 0 0 9 0 2
6 10 3 15 0 13 2
37 13 3 1 10 9 3 10 0 0 7 13 0 15 3 7 10 0 9 2 10 7 0 9 0 3 7 0 7 10 9 7 10 13 1 10 9 2
14 10 3 13 10 9 13 9 0 0 3 0 7 0 2
17 13 3 1 10 0 0 9 0 7 0 2 9 13 0 7 0 2
9 10 3 9 13 10 9 9 9 2
26 13 3 10 9 1 9 3 3 1 10 9 2 3 3 7 3 16 13 13 2 16 0 13 10 9 2
38 1 0 3 9 13 10 9 2 7 13 3 0 3 0 7 0 2 7 10 1 10 0 0 13 13 2 3 7 9 0 7 9 0 9 3 10 0 2
7 1 15 13 9 9 0 2
13 13 3 3 9 9 0 2 9 0 2 9 0 2
11 13 3 9 3 10 0 7 9 10 0 2
10 9 3 13 9 10 0 2 9 0 2
21 3 3 10 0 13 9 9 13 1 10 10 9 9 2 1 15 3 13 10 9 2
7 13 3 3 9 10 9 2
18 10 3 13 2 13 2 9 1 10 9 7 10 0 9 13 0 0 2
16 9 3 1 10 1 9 1 9 13 10 13 1 10 9 13 2
30 10 9 9 13 10 10 9 15 13 1 0 10 0 13 13 10 9 7 13 15 3 13 0 16 10 9 0 13 13 2
12 15 0 13 3 9 0 9 1 10 9 13 2
17 9 3 10 0 13 16 13 13 2 1 9 9 13 10 13 13 2
20 9 3 7 9 13 13 9 0 10 9 2 1 15 13 9 1 10 9 13 2
17 13 3 15 3 9 0 10 10 9 13 1 10 1 10 9 9 2
17 9 3 7 9 0 13 9 9 0 13 2 15 13 10 9 13 2
46 10 3 0 9 7 10 0 9 1 15 10 9 9 13 3 13 2 0 9 13 7 10 0 9 0 7 0 9 13 10 9 2 0 13 10 9 13 10 1 9 3 13 1 9 9 2
15 13 3 15 10 9 9 0 2 0 7 9 0 13 15 2
13 10 3 13 9 0 9 13 0 13 10 3 9 2
16 3 0 3 9 0 0 1 15 3 13 0 7 0 9 13 2
7 13 3 15 9 9 0 2
20 1 3 0 10 9 0 13 9 2 1 15 13 13 10 9 10 9 3 13 2
40 3 3 9 10 9 10 10 9 9 13 13 3 9 0 0 9 13 2 3 0 9 2 10 7 10 9 13 9 1 0 13 2 15 9 13 13 10 9 0 2
14 15 3 13 3 10 0 7 10 13 15 13 13 9 2
7 15 13 10 1 15 9 2
18 13 3 3 3 9 10 1 9 9 7 0 9 2 16 15 9 13 2
9 13 3 10 9 0 0 13 9 2
7 13 0 9 7 9 0 2
24 9 3 10 0 13 9 13 9 1 10 0 7 0 10 9 10 1 9 9 13 9 0 13 2
20 13 3 2 13 2 3 0 9 10 13 7 9 9 3 9 3 9 7 9 2
22 13 3 13 1 10 9 0 13 7 13 10 9 3 10 1 10 9 7 10 13 9 2
24 1 3 10 0 1 10 0 15 9 13 10 1 9 1 9 13 13 16 9 13 1 9 0 2
28 1 15 1 10 13 7 13 9 0 13 10 9 0 9 0 3 3 0 7 0 9 0 13 2 9 13 13 2
39 9 3 1 0 0 9 1 0 9 13 13 10 9 1 10 9 2 9 3 0 7 0 13 2 9 3 1 9 7 9 2 9 7 1 9 7 10 9 2
11 13 3 2 13 2 3 9 1 9 0 2
19 1 3 10 13 13 9 0 7 9 13 13 10 3 9 7 0 9 13 2
31 1 0 3 15 0 13 10 9 16 3 13 9 7 9 13 2 3 1 10 10 9 9 13 2 7 3 13 9 10 9 2
8 3 3 1 9 13 10 13 2
14 0 3 10 9 3 9 15 13 1 10 9 9 13 2
23 9 3 13 16 9 10 10 0 9 9 1 10 1 10 9 9 13 2 13 10 9 0 2
27 3 10 3 1 9 9 0 13 10 1 10 9 9 13 1 10 9 7 10 9 9 13 10 13 0 9 2
25 15 3 10 3 0 9 0 15 13 9 0 13 7 10 1 9 7 9 0 9 3 13 10 9 2
10 10 3 0 9 9 7 9 9 0 2
23 13 3 15 1 10 0 9 9 15 13 3 3 3 0 2 1 15 0 10 1 9 13 2
13 15 13 13 9 10 0 13 0 0 7 0 9 2
15 13 3 3 9 1 15 1 10 13 1 10 1 9 9 2
8 13 3 15 0 9 7 9 2
9 13 1 15 3 9 1 10 0 2
26 1 3 10 9 10 0 9 9 9 9 10 0 13 1 10 9 13 13 1 15 0 9 1 10 13 2
11 3 9 3 1 10 0 10 9 13 3 2
12 3 0 1 0 15 9 13 1 10 9 13 2
22 3 1 3 0 9 10 13 9 7 9 15 13 0 1 10 9 13 1 9 13 15 2
17 3 16 10 9 0 13 2 13 1 10 10 9 9 9 13 15 2
19 3 13 10 3 9 13 1 9 2 10 7 0 13 13 10 7 13 15 2
16 3 1 10 0 9 13 15 10 9 2 16 10 9 13 13 2
5 10 3 9 13 2
12 15 3 9 9 13 7 13 3 10 9 13 2
16 0 3 10 13 9 13 10 9 9 0 7 0 13 10 9 2
46 9 3 10 9 1 10 1 9 0 13 13 9 9 0 10 9 13 9 0 2 9 7 9 0 2 1 15 13 9 7 0 9 9 13 7 0 13 9 1 10 9 7 9 10 9 2
6 0 3 15 13 13 2
24 9 3 10 9 1 0 0 1 9 13 9 13 3 13 15 13 9 2 1 15 13 9 10 9
26 10 3 9 10 9 0 9 13 1 10 0 13 0 9 0 2 16 13 9 1 0 10 1 9 9 2
29 9 3 1 10 0 10 9 1 9 13 10 9 2 1 15 10 0 13 9 2 16 9 13 0 2 9 3 15 2
12 0 3 3 3 13 10 9 1 10 9 13 2
56 9 3 10 9 2 16 13 9 1 10 0 10 9 2 0 7 0 9 1 9 0 13 7 1 15 0 13 1 10 9 7 10 10 9 9 10 0 0 1 10 0 9 13 2 9 1 0 9 0 13 7 9 15 9 13 2
19 7 10 3 9 10 1 10 9 10 9 13 2 10 7 9 9 7 9 2
21 9 3 9 13 1 10 9 2 0 7 0 10 9 1 10 9 13 13 1 9 2
29 13 3 3 1 9 9 13 7 9 9 0 2 7 10 10 15 13 9 9 7 10 9 13 0 15 10 9 13 2
26 13 3 3 10 9 2 10 3 9 10 1 10 9 13 3 9 10 9 13 7 10 0 9 13 15 2
11 13 3 10 9 0 7 10 13 0 13 2
26 1 3 10 9 10 9 15 13 9 13 2 13 10 9 1 15 9 9 10 9 2 1 15 0 13 2
10 3 3 0 0 0 9 15 9 13 2
33 9 3 10 0 1 0 9 9 2 13 2 10 9 9 10 9 13 1 9 0 1 9 13 2 9 13 16 10 9 10 9 13 2
7 9 3 13 0 0 13 2
16 3 1 9 3 13 15 10 9 9 0 9 13 7 9 0 2
47 16 3 13 2 9 10 0 10 3 9 7 9 13 2 7 15 13 15 10 1 9 13 1 9 16 13 10 9 10 9 9 1 9 0 0 9 13 9 7 0 13 7 9 10 10 0 2
10 13 3 0 10 9 10 13 15 9 2
29 3 0 13 10 9 13 16 1 9 15 13 1 10 0 13 1 10 9 9 10 0 10 3 9 2 16 13 15 2
50 9 3 10 0 1 10 0 7 0 10 9 9 13 13 1 9 7 13 9 3 13 10 1 9 9 13 1 0 9 1 10 0 9 9 7 0 1 0 0 9 13 2 13 0 9 9 9 7 9 2
16 0 3 13 1 0 3 9 1 9 7 9 2 16 13 9 2
5 1 3 9 13 2
12 9 3 7 9 1 9 0 13 3 0 13 2
14 3 3 9 1 9 13 16 0 15 10 9 13 9 2
32 9 3 1 10 0 10 0 0 13 1 10 9 2 16 0 13 7 13 13 3 9 7 9 2 0 13 7 10 9 0 0 2
25 13 3 10 9 3 0 0 1 15 13 10 9 3 1 10 0 9 13 3 9 7 9 0 13 2
35 3 3 1 10 0 10 10 9 7 10 9 13 16 3 9 10 0 9 9 13 2 0 9 1 10 9 13 2 16 13 9 1 10 9 2
20 15 3 1 9 1 10 0 13 9 10 9 13 7 13 10 1 15 13 9 2
8 0 9 9 7 13 15 13 2
9 3 15 13 1 15 13 0 9 2
9 13 3 1 0 9 15 3 15 2
16 3 9 13 9 2 15 3 15 13 0 2 9 0 13 9 2
6 13 3 3 1 15 2
8 16 3 0 13 2 13 15 2
12 13 3 3 9 13 9 0 0 9 1 0 2
5 0 3 13 9 2
6 0 3 15 13 9 2
30 13 3 3 1 0 1 9 10 9 7 13 2 13 15 10 0 2 13 16 15 3 0 13 2 9 3 13 0 13 2
27 13 3 1 9 9 3 9 0 1 10 9 13 9 3 13 0 9 13 0 7 0 13 10 9 10 9 2
24 3 3 10 1 10 9 3 13 3 3 2 16 3 13 13 2 16 13 9 1 10 1 9 2
25 13 3 13 2 16 10 1 9 9 13 2 16 9 15 13 10 9 13 15 1 10 10 9 9 2
6 3 3 13 10 9 2
15 0 3 0 13 3 13 9 1 9 2 0 15 13 13 2
12 3 9 3 9 0 10 1 10 9 9 13 2
11 0 3 10 13 13 10 0 3 13 13 2
15 9 3 3 13 10 9 7 10 9 9 13 3 3 13 2
27 9 3 13 16 3 0 3 9 1 15 13 13 13 7 10 9 15 13 10 9 1 10 3 13 0 13 2
37 15 3 3 2 13 2 13 3 13 15 2 3 7 0 13 0 1 15 2 15 7 3 3 0 13 1 10 0 9 2 3 7 13 3 13 15 2
8 3 1 15 3 13 10 9 2
29 9 13 3 1 10 10 9 9 2 13 7 1 10 13 1 9 2 16 3 13 13 13 2 13 10 9 3 13 2
10 13 3 10 9 10 0 1 9 13 2
25 3 3 10 9 1 10 9 13 16 3 13 15 10 9 7 10 9 13 10 9 7 10 9 13 2
12 10 3 9 1 10 9 13 13 7 3 13 2
12 3 1 9 13 15 1 10 9 10 0 9 2
7 3 9 13 7 13 16 2
16 13 3 15 9 1 9 13 15 9 13 1 15 10 9 15 2
14 10 9 0 1 9 3 3 13 9 13 7 13 13 2
21 15 9 13 9 13 10 9 2 7 10 9 3 3 3 13 2 10 7 9 13 2
12 9 3 1 9 1 10 10 9 9 13 13 2
6 1 10 3 9 0 2
8 3 15 13 3 10 9 13 2
21 13 3 3 9 7 9 1 3 10 9 7 10 0 1 10 0 9 13 10 9 2
18 13 3 13 3 3 10 9 9 7 16 15 3 9 0 9 13 13 2
21 15 0 9 9 0 13 2 7 3 9 1 10 9 13 13 10 13 13 0 9 2
16 0 3 10 0 9 13 10 13 9 2 3 1 9 3 13 2
23 3 16 0 13 9 10 9 1 10 0 13 10 9 2 3 0 2 7 0 9 15 0 2
27 15 3 13 13 10 3 9 7 9 7 10 0 10 0 3 7 0 2 0 3 1 10 13 9 13 13 2
9 0 3 13 15 7 0 13 9 2
15 0 3 2 13 2 10 0 9 13 15 3 3 0 13 2
23 15 3 3 10 3 9 0 13 2 2 10 7 9 9 3 3 0 15 13 1 15 13 2
30 9 3 3 9 1 10 0 9 13 10 9 3 15 0 1 7 10 13 10 9 9 2 9 7 9 1 10 0 9 2
9 15 3 13 10 10 0 9 9 2
22 10 3 9 13 13 10 10 9 9 7 15 10 9 13 2 13 13 10 10 9 9 2
24 13 3 10 9 10 10 9 9 0 3 10 1 10 9 9 13 2 7 3 0 3 9 13 2
19 13 3 3 15 10 10 9 9 2 16 1 0 3 9 7 9 13 9 2
16 1 15 3 3 9 7 9 13 7 9 13 10 1 9 9 2
9 3 10 9 3 13 10 9 13 2
32 9 3 10 10 9 9 1 10 1 15 9 1 10 9 15 13 3 9 15 13 7 10 9 10 0 9 2 15 3 9 13 2
32 3 16 3 10 9 13 7 10 9 2 10 3 13 10 9 2 7 10 9 7 10 9 15 1 10 1 9 13 2 15 13 2
3 13 3 2
36 3 3 15 13 13 0 13 3 10 1 9 9 2 13 3 10 1 0 2 13 3 10 1 9 2 13 7 3 10 1 9 1 9 0 9 2
7 3 9 1 10 9 13 2
6 3 10 9 3 13 2
10 9 7 9 0 0 10 10 9 9 2
12 3 10 0 7 10 0 1 15 13 10 9 2
8 1 10 1 9 3 3 13 2
14 0 10 0 3 10 9 7 10 0 2 16 9 13 2
22 16 3 3 13 2 13 0 2 3 0 1 15 13 10 9 10 9 7 9 9 13 2
5 1 15 3 13 2
14 13 10 0 7 10 3 15 13 2 16 0 9 13 2
26 3 3 13 0 10 0 0 9 7 9 10 0 13 10 9 2 9 10 9 13 2 1 15 13 9 2
25 3 3 3 9 1 9 13 10 0 2 9 7 10 9 3 0 10 9 10 15 9 2 13 15 2
16 13 15 3 0 16 0 13 9 1 10 9 3 1 10 9 2
43 16 3 3 13 10 9 2 13 9 13 16 10 3 9 0 13 1 10 9 3 2 10 7 9 0 3 13 1 15 13 3 13 2 7 10 9 15 1 9 13 10 0 2
5 3 3 3 13 2
15 10 3 9 1 9 9 13 9 10 9 1 9 15 13 2
18 10 3 9 7 13 9 2 3 13 15 13 15 2 7 0 13 0 2
16 13 3 3 1 9 2 16 13 2 0 7 13 9 9 13 2
19 16 3 13 15 10 13 2 15 15 9 9 3 3 13 9 1 10 9 2
32 3 9 3 10 0 2 16 13 9 10 0 2 1 9 13 9 1 10 9 1 0 9 7 0 0 10 13 13 9 3 13 2
15 0 3 3 10 9 13 13 10 0 9 7 9 0 13 2
51 1 3 10 13 1 15 9 3 9 7 9 10 0 9 3 10 10 9 9 7 10 10 9 7 9 9 15 13 16 0 13 7 13 13 1 10 9 13 2 3 1 9 0 7 9 7 9 0 13 13 2
17 15 3 0 13 9 3 0 7 9 13 2 9 7 7 9 0 2
17 15 3 0 13 0 1 10 0 10 3 9 7 10 9 10 13 2
28 10 3 9 1 9 3 1 10 0 10 9 9 1 10 9 9 13 0 9 2 15 13 0 15 1 10 9 2
10 13 3 10 9 3 9 0 7 0 2
12 1 3 9 9 10 9 1 0 9 3 13 2
33 10 0 13 9 1 10 10 13 9 13 9 0 3 13 9 0 10 13 13 9 10 15 2 13 1 9 10 10 3 15 13 9 2
25 10 3 9 9 13 7 1 10 9 9 13 10 9 2 16 3 9 13 7 10 9 10 13 13 2
15 3 3 3 15 13 10 0 0 9 10 1 10 9 9 2
31 0 3 15 0 9 10 9 2 1 15 13 10 15 9 1 10 0 10 9 16 1 10 3 13 3 0 9 10 13 13 2
26 3 16 15 15 13 0 9 13 3 3 7 1 9 0 9 13 2 15 3 2 13 2 9 1 13 2
34 9 3 10 0 1 0 1 9 9 2 13 2 10 9 13 15 15 13 0 10 13 0 10 12 9 2 13 10 15 3 0 1 13 2
49 9 3 0 9 10 9 7 10 0 1 10 9 9 0 13 2 16 13 13 10 0 10 9 15 13 15 9 13 10 9 2 16 3 15 15 13 2 10 0 13 2 13 2 1 0 9 7 9 2
38 9 3 10 0 1 0 9 9 2 13 2 10 0 9 10 0 9 9 13 9 13 0 3 10 9 0 2 1 15 13 2 9 7 0 7 9 0 2
15 9 3 1 10 9 1 9 13 3 10 9 1 9 13 2
18 3 9 3 10 15 9 13 13 1 10 9 2 0 13 10 9 9 2
30 0 3 3 15 0 10 9 13 1 10 0 9 2 10 7 3 1 9 9 13 2 15 7 3 1 9 1 0 9 2
26 3 13 10 9 13 9 0 10 9 13 2 15 1 10 9 7 10 9 13 16 1 9 13 0 13 2
16 1 3 3 15 1 10 13 1 10 9 9 3 13 10 9 2
14 16 3 1 10 0 9 10 9 13 13 2 3 13 2
26 10 3 9 13 10 13 13 9 10 9 16 10 3 0 9 13 2 10 7 9 0 13 13 10 13 2
21 13 3 15 9 0 3 13 0 1 10 9 2 10 9 13 1 15 9 1 9 2
7 0 3 9 13 1 9 2
8 13 2 16 3 0 13 9 2
25 13 3 13 9 0 1 10 0 2 15 13 0 7 0 2 0 10 1 15 9 9 7 9 13 2
23 9 3 10 0 2 13 9 10 9 13 1 9 7 13 15 2 13 1 0 10 9 3 2
17 1 3 9 13 10 9 1 9 7 9 9 2 15 0 13 13 2
9 13 3 3 0 16 3 1 9 2
41 16 3 9 3 13 0 10 9 15 2 15 1 15 13 1 10 0 10 9 13 16 3 9 13 10 1 9 9 7 16 9 13 10 1 15 13 9 2 13 3 2
38 15 3 13 0 9 13 3 0 9 2 1 15 0 3 10 0 13 13 2 0 3 13 16 3 10 0 9 2 3 7 0 9 9 3 0 0 9 2
8 3 3 15 3 0 9 13 2
18 1 9 3 13 3 10 9 15 9 2 10 10 15 9 13 13 15 2
36 10 3 10 9 9 13 3 1 10 9 2 13 3 1 10 1 15 2 1 0 7 9 13 2 3 13 0 3 13 2 16 3 0 13 13 2
18 1 3 10 1 10 9 9 1 0 9 13 0 0 15 10 13 13 2
42 1 3 0 10 15 13 1 10 0 7 0 3 10 13 9 13 2 16 15 3 10 9 0 13 7 10 9 10 9 0 13 2 0 1 0 9 13 10 9 10 0 2
19 13 3 10 9 3 1 0 9 3 10 1 10 9 7 10 9 10 0 2
13 3 3 9 13 1 0 9 9 2 15 7 15 2
20 3 9 3 10 0 9 2 16 9 13 10 9 0 2 3 13 0 10 9 2
12 3 10 9 3 13 1 15 13 1 9 13 2
8 3 3 9 13 0 15 0 2
11 16 3 13 2 3 10 13 15 9 13 2
12 13 3 3 10 9 1 10 9 10 9 13 2
14 10 3 13 0 15 13 3 9 2 9 0 7 9 2
10 3 15 9 9 7 9 9 13 13 2
19 9 3 1 0 9 13 0 13 9 2 15 13 13 9 7 3 3 13 2
8 13 3 0 9 1 15 9 2
3 0 13 2
5 3 15 3 13 2
4 3 3 13 2
8 3 3 1 0 9 13 3 2
10 1 3 10 9 3 9 1 9 13 2
11 1 3 9 0 10 9 1 9 13 3 2
32 13 3 3 0 7 0 10 9 2 1 15 3 0 9 13 9 2 9 9 15 13 1 10 1 10 15 9 3 10 9 13 2
10 13 3 1 10 9 15 13 9 9 2
29 15 3 15 2 16 3 9 2 3 13 0 9 1 10 9 13 9 13 16 3 13 1 3 10 9 7 10 9 2
32 16 3 13 10 9 0 7 0 15 9 10 9 1 10 1 9 0 13 9 13 2 13 15 13 10 9 13 7 1 15 13 2
27 16 3 10 9 13 7 3 0 2 3 15 13 13 1 10 3 1 9 13 13 7 1 10 9 15 13 2
6 13 3 3 10 9 2
25 13 3 16 3 3 13 16 9 13 10 10 9 0 2 15 15 0 13 0 0 7 0 9 13 2
25 3 15 13 10 15 1 9 13 15 10 3 15 0 13 3 13 2 10 9 7 13 1 0 9 2
32 3 1 15 3 9 3 9 7 9 13 2 0 9 13 10 9 2 1 7 9 9 15 0 9 13 2 13 3 10 15 9 2
20 3 3 16 15 13 10 9 13 2 7 16 13 10 9 7 10 9 10 0 2
39 10 3 3 13 7 13 3 0 15 0 13 2 10 7 3 13 0 9 13 7 1 0 9 13 3 13 13 10 9 15 0 13 10 10 15 15 15 13 2
9 1 3 3 9 15 10 9 13 2
30 0 3 13 3 9 10 0 9 2 15 3 1 10 10 9 9 9 1 9 13 13 1 10 9 16 3 1 9 13 2
24 9 3 10 9 1 10 1 9 9 13 10 9 13 1 0 7 1 9 13 9 9 13 13 2
30 10 3 15 13 16 3 9 9 3 0 13 2 9 7 13 10 9 2 7 16 13 9 10 9 9 0 10 9 13 2
7 13 3 0 2 0 13 2
13 13 3 0 10 9 1 9 2 16 10 9 13 2
6 9 3 1 9 13 2
8 1 9 0 0 15 13 9 2
7 3 1 9 0 9 13 2
11 9 15 10 0 15 13 9 0 13 9 2
12 16 3 3 13 13 10 13 9 1 9 13 2
10 3 13 2 9 0 1 9 13 13 2
6 3 15 3 15 13 2
4 0 3 13 2
16 0 3 0 13 15 0 13 10 9 16 7 13 9 1 9 2
36 9 3 10 0 1 10 1 9 9 13 10 9 1 9 1 9 13 7 0 9 13 2 16 1 10 9 13 2 1 9 13 13 15 10 9 2
19 9 3 13 9 3 10 9 10 13 13 9 2 16 9 3 1 9 13 2
8 3 10 9 3 13 15 9 2
17 1 3 9 15 9 0 2 0 3 7 0 2 10 9 13 0 2
21 1 3 9 13 15 3 13 13 10 10 9 9 16 1 9 10 9 10 9 13 2
6 3 13 3 10 9 2
12 3 3 13 10 0 9 2 3 7 13 9 2
7 3 9 15 13 9 9 2
9 3 10 9 13 15 10 0 9 2
14 16 0 10 9 3 13 15 10 9 13 7 2 13 2
13 3 3 3 13 9 15 7 10 9 3 0 13 2
21 15 3 15 0 15 15 13 13 2 0 0 7 9 13 9 2 3 3 0 13 2
4 13 3 3 2
13 3 10 1 9 3 9 9 1 9 0 13 13 2
12 9 3 1 9 10 9 13 10 10 0 13 2
16 1 15 3 16 9 10 9 10 0 1 9 13 7 13 15 2
6 3 0 1 15 13 2
18 10 3 10 0 9 7 9 9 1 9 10 10 9 9 13 10 13 2
18 3 10 15 9 9 7 9 10 1 10 13 9 10 9 13 13 15 2
18 3 3 0 13 10 0 9 2 16 3 1 9 13 10 0 9 13 2
13 13 3 10 10 0 13 7 1 10 0 3 13 2
15 3 0 10 13 0 13 1 10 9 7 13 10 0 13 2
19 3 10 3 1 10 9 13 13 2 7 9 13 13 9 13 9 3 0 2
17 3 3 13 10 9 10 3 16 3 9 9 9 13 1 15 9 2
7 9 0 13 0 9 9 2
14 15 13 3 1 15 13 1 10 0 13 0 13 0 2
14 3 3 13 9 9 9 7 0 13 13 15 3 15 2
7 3 15 13 13 10 0 2
20 15 3 1 9 13 13 1 9 0 13 7 13 10 13 10 9 15 13 0 2
30 10 3 9 16 13 15 0 13 9 3 13 2 13 1 10 9 10 9 15 2 13 15 10 9 2 7 13 10 9 2
19 15 3 1 10 9 9 13 2 16 3 10 9 9 1 10 9 13 13 2
6 13 9 9 1 9 2
21 15 3 13 9 0 13 9 9 13 9 10 9 2 16 13 3 9 1 10 9 2
19 1 9 3 9 0 13 3 3 10 0 9 13 1 10 1 9 3 13 2
45 10 9 9 10 9 13 3 1 9 15 16 0 10 9 10 1 10 9 13 13 15 13 2 7 13 15 3 13 3 13 7 13 13 1 9 0 0 3 15 13 15 9 9 13 2
17 3 10 3 13 15 13 2 10 7 13 13 7 13 1 0 9 2
34 16 3 10 9 15 9 1 9 13 13 15 13 9 7 10 9 13 2 13 3 1 10 1 9 9 2 3 13 1 10 9 13 0 2
34 3 3 10 9 10 0 15 9 13 9 13 1 10 1 9 13 16 1 9 1 9 15 0 0 13 10 9 2 13 3 10 0 9 2
9 3 0 15 13 2 15 13 0 2
13 3 3 9 13 16 13 10 0 0 13 0 13 2
42 9 3 10 0 1 10 1 9 1 9 2 13 2 10 0 10 9 1 9 15 1 10 9 13 13 2 16 10 1 10 9 9 13 13 3 7 1 9 13 10 9 2
19 1 3 9 0 9 0 9 13 2 3 10 0 13 10 9 7 9 13 2
17 3 3 13 15 0 13 2 3 13 10 0 1 10 9 10 9 2
25 13 3 9 2 9 10 0 2 9 10 0 2 9 2 15 10 0 9 13 13 15 10 1 9 2
17 13 3 1 10 9 9 9 10 0 2 15 15 13 13 10 9 2
12 13 3 10 13 1 10 9 9 9 10 0 2
40 1 3 9 13 10 9 10 9 10 9 1 10 16 9 13 10 9 10 9 2 3 7 3 1 10 10 9 2 16 13 9 1 10 0 2 1 10 9 13 2
13 3 10 9 3 0 13 9 7 10 9 3 13 2
5 13 3 10 9 2
15 1 3 10 9 3 13 10 10 9 9 10 10 9 9 2
25 9 3 3 13 10 9 16 13 0 3 13 3 15 10 9 9 2 3 1 10 0 7 0 13 2
28 3 10 9 3 0 13 10 9 1 15 10 9 13 2 15 1 10 9 10 9 13 2 1 9 13 0 9 2
22 13 3 3 15 2 13 9 2 16 0 10 9 9 13 9 13 9 2 0 13 9 2
33 3 3 13 15 13 10 9 1 10 10 9 9 3 1 9 3 1 0 7 3 1 10 1 10 9 9 2 16 3 13 10 9 2
17 13 3 10 9 13 9 13 10 9 2 1 15 3 10 9 13 2
7 3 13 10 1 15 9 2
9 10 3 9 16 9 1 9 13 2
19 0 15 9 9 2 0 7 9 13 1 9 0 2 15 15 9 0 13 2
20 3 3 13 2 13 10 9 2 1 9 13 10 9 10 9 2 7 1 9 2
10 3 3 10 0 9 1 10 13 13 2
10 1 15 3 10 10 9 15 9 13 2
14 1 0 3 3 9 0 13 9 9 2 16 9 13 2
6 9 3 13 3 9 2
14 0 3 3 13 10 9 9 2 1 15 10 9 0 2
9 13 3 0 0 13 0 1 9 2
10 3 10 9 13 9 2 1 15 9 2
9 9 3 9 13 3 3 9 13 2
32 9 3 1 10 0 10 0 13 10 10 9 13 9 13 10 3 15 1 9 13 2 10 3 1 9 2 15 7 1 0 9 2
21 9 3 13 3 9 7 9 2 1 15 3 10 1 9 9 13 2 16 13 9 2
6 9 3 13 3 9 2
10 1 3 10 9 3 1 9 13 9 2
7 1 3 10 9 9 13 2
40 9 3 10 9 3 13 3 1 10 9 9 2 16 9 10 1 9 13 2 15 1 10 0 9 0 0 13 9 2 16 13 9 1 0 1 10 10 9 9 2
8 10 3 9 3 1 9 13 2
28 1 9 3 0 7 0 15 13 2 16 13 9 1 10 1 10 9 15 2 9 9 13 13 1 15 9 9 2
9 13 3 3 9 9 9 7 9 2
16 13 3 3 10 9 9 13 9 2 1 15 13 9 7 9 2
23 3 10 9 3 16 13 2 13 1 15 9 10 10 9 9 13 9 10 9 7 9 0 2
8 13 3 3 15 13 10 9 2
15 1 0 3 13 9 13 10 9 3 9 2 9 7 9 2
12 3 15 13 10 9 0 10 9 10 15 13 2
21 3 3 1 15 10 9 10 3 9 3 3 0 2 13 2 7 3 0 9 13 2
19 3 10 9 13 13 15 1 9 13 9 10 9 2 7 15 15 10 9 2
14 3 1 15 9 3 1 9 13 2 9 7 1 9 2
12 3 10 9 3 13 10 9 9 10 13 9 2
8 9 3 13 3 9 10 9 2
8 9 3 1 0 9 13 3 2
17 13 9 15 16 9 13 9 2 1 3 10 9 2 13 10 9 2
14 10 3 9 15 9 3 13 15 0 9 13 1 9 2
39 16 13 10 9 2 1 10 3 9 9 0 13 0 2 1 3 10 9 9 1 10 9 9 0 13 2 1 10 9 7 10 9 13 13 9 2 0 9 2
19 9 3 1 9 13 15 9 9 13 3 2 15 3 9 13 3 0 13 2
3 3 13 2
7 15 3 0 13 10 9 2
18 13 3 13 1 9 0 3 10 9 2 15 16 10 9 13 10 0 2
10 9 0 3 9 15 15 10 9 13 2
10 10 9 3 3 13 3 9 13 3 2
17 9 3 15 2 13 7 10 9 3 2 16 13 15 13 0 0 2
9 10 3 9 15 3 13 9 13 2
16 3 0 13 9 10 0 13 3 13 2 7 13 9 0 9 2
18 10 3 9 10 9 3 3 3 13 2 10 7 9 13 13 15 9 2
8 10 9 3 3 9 13 13 2
10 9 7 9 9 2 10 9 7 9 2
28 9 0 3 0 13 10 9 13 2 15 13 3 3 15 2 7 1 9 15 2 16 13 3 13 7 13 3 2
23 3 0 15 13 2 13 2 9 7 9 2 7 3 9 0 2 7 2 13 2 9 0 2
20 3 10 3 13 15 13 3 16 9 2 3 13 13 15 2 13 7 0 0 2
13 10 3 13 13 3 13 13 7 13 3 1 9 2
12 13 3 3 9 13 9 0 3 13 9 0 2
22 15 0 10 9 13 10 9 13 10 10 9 9 10 1 10 9 9 13 15 10 9 2
8 16 13 9 2 3 9 13 2
9 10 10 3 9 13 1 15 9 2
14 10 3 3 9 13 13 2 15 7 13 3 13 3 2
22 15 3 13 13 2 15 7 13 13 13 2 13 2 3 9 0 13 7 13 13 3 2
6 9 3 1 9 13 2
15 3 13 10 9 3 0 2 15 10 9 3 3 9 1 2
8 3 3 9 13 0 9 9 2
23 10 3 9 3 13 3 13 2 10 7 13 16 3 10 9 0 9 13 7 1 15 0 2
8 0 3 13 15 9 0 13 2
7 10 3 0 3 13 3 2
4 3 13 13 2
6 13 15 7 9 0 2
4 9 13 0 2
7 3 3 9 13 3 15 2
20 6 0 2 3 3 15 10 0 9 13 2 10 7 3 0 3 13 0 13 2
8 0 3 13 10 13 0 0 2
7 10 3 3 0 15 13 2
10 3 3 13 15 0 13 0 13 9 2
11 10 3 0 13 1 0 13 15 13 0 2
3 13 3 2
4 15 15 13 2
10 3 13 2 15 15 13 13 7 13 2
12 3 13 2 16 9 13 2 15 13 10 9 2
4 13 3 15 2
7 1 15 15 13 3 13 2
3 13 9 2
5 13 2 13 3 2
7 13 3 3 9 13 3 2
25 0 13 15 3 10 0 13 13 2 3 10 0 2 3 10 0 2 3 10 0 2 7 10 9 2
14 9 3 10 0 1 9 2 15 9 6 9 2 13 2
8 13 3 13 16 9 13 0 2
23 3 13 3 3 10 1 9 0 13 9 1 0 0 15 13 2 3 10 0 9 13 15 2
9 3 3 0 13 9 0 9 9 2
11 3 3 9 13 16 9 2 7 9 13 2
10 13 3 9 3 1 9 0 13 9 2
7 3 9 3 1 9 13 2
7 3 0 0 13 9 9 2
20 16 3 9 3 0 13 9 9 2 10 9 13 7 1 9 0 9 13 13 2
13 0 3 3 15 13 10 0 9 9 13 9 13 2
8 3 3 13 10 9 10 9 2
44 3 10 0 3 9 13 2 16 13 9 1 10 1 10 0 9 2 16 9 1 9 13 2 0 13 2 13 9 10 9 10 9 9 9 7 10 9 9 13 1 10 0 9 2
8 0 3 9 13 3 10 9 2
8 13 3 3 0 9 1 9 2
27 10 3 9 13 10 0 9 1 10 9 13 10 15 13 1 9 10 9 9 2 0 13 1 9 10 9 2
17 10 3 10 3 15 3 13 2 13 3 9 13 15 9 7 9 2
7 13 3 10 9 9 9 2
18 10 3 9 13 10 9 9 1 10 13 9 1 9 7 13 1 9 2
20 9 3 1 10 0 7 9 10 9 1 0 0 10 9 9 13 13 1 9 2
16 9 3 10 0 3 0 13 9 13 0 9 10 9 7 9 2
20 1 15 10 9 13 10 13 10 9 1 10 9 3 15 15 13 7 1 9 2
6 3 13 9 0 0 2
16 1 15 15 3 13 10 0 9 9 9 2 15 13 3 15 2
19 9 3 9 9 2 9 0 13 2 7 13 15 10 9 0 0 13 0 2
10 3 3 0 9 15 13 1 9 13 2
13 10 3 0 10 15 9 3 13 1 7 0 13 9
16 10 3 13 13 10 0 3 3 13 2 13 7 3 16 13 2
9 3 1 10 9 3 15 15 13 2
9 13 3 13 7 9 13 1 9 2
8 0 3 15 13 10 9 15 2
22 3 15 3 13 0 0 13 2 3 13 7 1 15 10 13 13 13 9 15 13 15 2
18 3 3 1 10 9 13 10 9 9 13 0 13 1 10 10 9 9 2
18 15 13 9 3 7 9 13 2 1 15 10 0 9 10 15 13 13 2
25 9 3 15 13 10 9 0 13 13 10 9 16 10 9 3 10 9 13 3 10 9 13 13 15 2
12 3 1 10 0 3 9 7 3 10 9 13 2
21 9 3 1 10 9 9 13 2 3 1 10 10 13 9 13 10 9 3 7 9 2
21 3 9 3 1 10 9 10 0 10 9 13 1 15 13 10 9 2 16 9 13 2
28 10 3 1 9 0 9 13 13 1 0 7 13 2 10 10 9 9 13 2 13 9 0 1 0 7 0 9 2
22 1 15 9 3 9 9 13 2 7 10 9 13 13 13 0 10 1 10 9 15 9 2
10 15 13 10 9 13 10 1 9 9 2
14 13 3 1 9 1 10 0 7 10 9 13 13 15 2
30 13 3 3 0 7 9 2 3 3 9 7 9 2 3 0 7 3 0 2 7 13 3 2 9 9 7 0 9 13 2
29 3 15 15 2 3 10 9 7 9 2 3 13 15 15 13 2 7 3 13 3 15 15 2 3 7 13 10 9 2
12 15 13 10 13 0 9 3 7 13 9 0 2
16 3 15 13 1 9 13 2 7 13 0 10 9 10 10 9 2
16 13 3 3 0 7 0 13 10 13 10 9 2 0 7 3 2
8 3 3 3 13 9 15 9 2
6 9 2 16 13 15 2
24 9 3 1 10 0 9 13 10 0 13 16 10 9 10 13 10 9 13 2 3 3 10 9 2
12 15 13 3 13 9 2 13 7 7 13 0 2
16 10 3 0 0 9 3 1 10 13 1 10 13 9 13 3 2
8 15 3 13 10 13 13 9 2
33 15 13 3 0 3 0 13 13 3 13 10 9 3 13 7 0 10 9 2 0 2 0 2 0 2 0 1 10 0 2 13 0 2
8 15 13 10 13 3 9 13 2
8 3 3 15 13 10 9 0 2
15 16 3 13 15 10 9 10 9 2 13 15 0 1 13 2
9 9 0 2 9 0 2 9 0 2
12 15 13 13 0 7 10 0 13 15 13 3 2
14 3 3 3 13 13 1 10 9 10 0 3 7 9 2
10 13 15 3 13 9 16 13 1 15 2
9 1 3 10 13 9 1 9 13 2
3 15 13 2
16 3 15 13 7 16 9 9 13 3 10 13 3 13 15 13 2
12 13 3 16 13 3 10 9 7 10 9 13 2
36 3 15 13 9 10 0 10 0 3 3 13 1 10 0 1 10 0 0 1 15 9 2 0 15 1 10 9 13 16 0 2 15 9 13 9 2
15 10 1 9 15 2 13 2 13 1 9 9 1 15 13 2
9 3 3 3 3 0 9 13 9 2
18 9 3 1 10 9 10 9 13 13 0 2 3 10 9 7 10 9 2
20 13 3 15 15 3 3 13 10 9 7 10 9 7 13 10 0 7 10 0 2
21 3 3 10 0 9 13 2 16 3 10 9 13 2 3 3 13 10 13 13 9 2
6 10 3 9 9 13 2
25 3 10 9 3 13 10 9 1 15 15 10 9 10 13 13 7 10 9 2 1 15 10 9 13 2
14 9 3 3 1 10 9 10 9 13 13 10 9 13 2
21 15 13 3 15 2 13 7 15 2 0 13 9 2 16 9 1 9 13 13 9 2
34 9 3 10 0 10 9 13 13 10 9 3 13 15 13 10 9 2 7 13 10 9 13 10 13 2 16 1 0 13 10 10 13 9 2
4 13 3 3 2
10 9 3 13 9 9 0 9 13 9 2
6 10 3 9 15 13 2
30 10 3 10 0 9 9 13 10 9 7 13 15 10 9 2 13 10 9 0 3 15 13 7 10 9 13 2 13 3 2
13 9 3 1 10 9 13 13 1 0 9 9 9 2
9 15 3 13 10 9 13 10 13 2
12 3 3 3 2 16 15 13 2 13 10 9 2
15 13 3 3 10 9 1 3 10 9 7 10 10 9 9 2
6 13 3 3 10 9 2
14 10 13 10 9 1 9 13 2 10 0 3 13 15 2
24 3 3 9 10 9 9 0 13 13 2 7 1 9 13 3 3 0 10 0 13 9 13 9 2
6 3 3 9 13 3 2
13 16 13 15 7 13 13 2 0 15 13 15 0 2
20 3 3 13 13 15 13 7 0 10 9 13 0 2 7 0 15 15 13 0 2
14 1 15 9 0 15 13 2 16 3 15 15 13 13 2
10 9 3 13 15 3 13 10 9 13 2
14 3 15 13 13 10 9 16 9 15 13 7 3 9 2
28 0 3 15 1 9 13 3 13 3 13 7 15 3 13 2 0 3 13 13 15 13 10 9 2 3 7 13 2
17 1 9 3 9 13 3 13 3 10 13 15 13 1 10 0 13 2
15 1 9 3 9 13 10 13 9 9 15 0 0 13 15 2
8 3 15 3 10 0 13 9 2
51 10 3 0 0 9 2 16 13 9 10 0 2 13 15 2 3 10 13 2 1 10 9 7 10 0 9 13 16 10 13 15 10 9 7 3 13 13 0 7 0 2 16 10 10 9 13 9 0 7 0 2
38 13 3 13 10 9 7 10 9 13 1 10 10 9 9 3 13 3 9 13 0 3 9 13 10 9 7 9 13 10 3 9 13 7 0 0 13 9 2
7 13 3 3 15 10 9 2
13 3 3 1 10 9 10 0 13 7 15 13 13 2
32 1 9 3 3 9 13 9 2 7 10 0 10 10 9 13 9 13 2 10 3 0 10 9 13 2 10 7 0 10 9 13 2
26 9 3 10 9 13 16 1 10 9 13 0 3 10 0 7 9 10 0 2 0 13 10 9 10 9 2
40 3 3 13 1 9 10 9 2 9 15 0 13 2 0 7 0 7 0 2 16 13 1 10 0 2 13 10 9 15 2 13 16 9 1 9 10 9 13 13 2
4 9 3 13 2
13 3 10 1 9 3 9 13 10 9 10 9 13 2
7 3 0 9 1 9 13 2
17 13 3 3 15 10 9 1 10 9 10 9 2 3 1 0 13 2
9 13 3 1 9 10 9 15 13 2
12 0 3 3 15 3 3 13 9 7 3 0 2
5 9 3 9 13 2
22 13 3 3 0 10 0 9 2 16 3 3 10 0 13 9 2 16 13 9 1 0 2
10 16 13 3 2 10 9 9 0 13 2
25 9 1 9 13 1 15 2 7 1 9 10 9 13 9 9 10 9 9 1 15 2 16 0 13 2
6 10 9 3 15 13 2
4 15 3 13 2
25 1 9 3 3 10 0 10 9 1 9 9 13 2 9 13 2 9 13 3 2 16 3 1 9 2
14 9 3 10 9 10 0 13 10 9 9 3 0 13 2
10 15 3 3 3 10 0 10 0 13 2
13 13 3 10 9 10 9 10 13 10 9 10 9 2
23 1 9 3 10 9 3 13 0 13 1 10 9 7 10 9 7 13 13 10 0 10 9 2
19 15 1 10 9 7 10 9 3 13 2 3 9 10 9 1 10 0 13 2
12 1 9 3 13 7 13 15 3 16 9 13 2
7 13 3 13 2 3 13 2
25 9 3 1 10 1 9 2 16 0 10 9 2 10 9 13 13 15 1 9 13 13 1 0 9 2
19 15 3 13 9 10 0 2 15 9 1 10 0 1 10 9 0 13 13 2
20 3 3 13 3 15 15 3 0 13 2 16 9 3 9 3 7 9 10 9 2
16 13 3 15 3 15 3 13 9 1 10 1 10 1 9 9 2
3 9 13 2
9 3 3 3 9 15 13 9 13 2
5 3 13 10 9 2
16 0 3 10 10 9 9 2 10 10 9 13 16 9 9 9 2
36 3 3 13 0 10 9 2 16 1 9 13 16 13 2 16 9 13 10 10 9 1 10 1 9 10 9 9 2 10 0 15 9 13 13 9 2
14 13 3 9 2 16 9 13 1 0 2 10 13 9 2
7 13 3 0 13 3 0 2
11 3 3 13 15 15 13 1 9 1 9 2
25 3 15 10 0 9 13 16 3 10 9 13 3 7 13 0 3 13 0 13 1 0 10 9 13 2
11 3 1 10 13 3 9 10 0 9 13 2
10 15 10 9 3 9 13 1 9 13 2
34 0 10 9 13 15 13 2 15 3 1 15 3 3 13 2 1 7 9 3 9 3 9 0 7 15 9 10 9 3 13 0 7 13 2
20 9 3 1 10 13 9 0 10 0 9 7 10 1 9 9 10 9 3 13 2
13 16 3 13 3 2 13 0 9 2 0 10 9 2
16 3 13 15 2 16 3 10 9 7 10 9 0 13 13 3 2
5 13 0 15 13 2
6 9 1 10 9 13 2
3 0 15 2
12 9 0 13 10 7 9 1 10 9 13 13 2
5 15 10 9 13 2
5 3 13 15 9 2
11 13 13 15 2 16 10 9 13 10 13 2
4 9 0 13 2
9 9 13 15 15 15 13 10 0 2
14 0 13 15 0 10 9 16 9 15 1 10 3 13 2
6 10 9 0 13 15 2
3 13 0 2
4 13 13 9 2
3 13 9 2
5 3 3 15 13 2
3 9 13 2
6 0 13 10 9 15 2
4 15 0 13 2
4 0 9 13 2
33 16 3 3 13 13 2 13 10 9 3 2 16 10 9 10 13 3 2 16 3 13 9 9 2 9 9 13 0 0 1 10 9 2
12 3 10 9 13 2 16 3 13 16 7 3 2
7 9 1 0 13 10 9 2
18 3 3 9 0 13 2 10 9 9 15 0 15 13 7 13 9 13 2
8 3 3 13 1 10 9 9 2
13 1 15 3 3 7 13 15 0 13 9 10 9 2
13 3 1 9 16 9 10 9 7 3 9 2 13 2
13 15 9 3 0 13 3 2 3 3 0 13 0 2
11 9 15 10 0 13 2 15 9 9 13 2
24 13 3 3 9 1 9 10 3 15 13 7 13 1 10 0 9 7 10 0 10 9 15 13 2
12 0 2 0 3 0 1 10 9 13 10 0 2
43 15 13 13 15 15 13 2 0 2 0 2 0 2 0 2 0 2 0 2 0 2 0 2 0 2 3 9 13 13 3 2 3 1 9 3 13 9 7 1 9 13 9 2
19 15 13 3 13 7 10 3 9 13 13 9 2 10 7 9 2 10 0 2
17 3 15 0 13 3 2 3 2 1 9 2 1 9 2 0 9 2
7 3 10 3 9 3 13 2
8 15 3 1 0 13 9 9 2
6 13 0 2 16 13 2
3 0 13 2
6 3 3 15 13 13 2
4 13 13 15 2
6 3 10 9 13 13 2
2 13 2
11 3 13 3 0 9 7 9 2 7 13 2
2 13 2
7 13 13 2 0 13 15 2
48 3 9 3 10 0 13 9 0 9 2 7 13 1 10 15 9 10 9 2 16 3 10 0 9 13 2 13 10 0 9 16 9 1 10 9 9 7 10 13 1 15 9 1 9 13 10 0 2
9 9 3 9 13 3 9 13 0 2
10 3 10 9 9 13 13 9 9 0 2
11 3 9 10 9 13 9 0 1 0 9 2
23 15 3 0 13 9 9 2 9 13 1 9 2 1 15 9 3 1 10 0 9 15 13 2
25 0 3 9 0 13 7 9 2 10 1 9 13 13 7 13 0 2 13 7 0 15 13 10 9 2
18 15 3 16 13 0 1 10 9 9 13 7 9 0 13 1 10 9 2
14 16 3 13 3 2 3 9 1 10 9 13 13 3 2
6 3 15 13 13 9 2
8 3 9 3 3 13 3 9 2
23 15 3 16 13 3 9 7 0 2 1 10 9 13 13 2 13 7 3 15 9 0 3 2
22 16 3 0 10 9 3 13 10 9 7 13 10 9 2 13 3 15 0 13 16 13 2
20 13 7 3 3 13 2 13 3 3 9 7 9 2 13 7 3 9 7 0 2
16 13 3 10 9 3 9 1 9 7 0 9 15 13 1 15 2
6 10 1 9 9 13 2
6 13 15 15 0 9 2
6 3 15 0 13 9 2
8 13 2 9 13 2 10 9 2
15 3 13 16 3 13 0 13 13 3 2 16 13 13 9 2
11 7 0 13 15 2 16 1 9 13 9 2
13 3 3 13 9 16 0 9 13 2 13 10 9 2
7 3 0 13 7 0 13 2
18 13 3 15 15 9 13 15 13 0 9 9 2 16 15 13 10 0 2
12 1 15 13 10 0 9 1 10 1 9 3 2
5 15 3 13 0 2
22 13 3 3 10 0 9 3 7 3 7 10 9 10 0 7 0 9 2 16 10 9 2
9 15 3 9 10 0 0 3 13 2
9 9 7 9 3 3 0 13 9 2
39 13 3 3 10 13 9 7 10 1 9 13 13 2 3 3 1 10 0 13 2 7 1 10 0 2 3 3 7 9 1 9 1 10 9 10 9 13 13 2
11 0 3 13 9 10 9 3 3 0 13 2
13 3 3 13 2 16 13 13 15 15 2 13 3 2
30 13 3 13 10 9 16 0 2 7 10 9 13 3 2 13 2 13 13 3 0 3 7 13 0 15 10 13 13 0 2
9 9 3 1 9 0 9 13 13 2
30 3 3 13 3 2 3 16 15 10 9 13 9 13 10 9 7 10 9 13 3 2 7 0 0 3 13 16 9 0 2
12 10 3 15 9 13 10 9 3 3 13 0 2
20 16 3 15 3 13 9 10 13 15 13 1 9 2 1 10 9 9 9 13 2
15 3 15 3 3 16 13 9 2 9 7 1 9 13 13 2
8 3 3 3 13 3 0 15 2
13 1 15 10 9 0 3 10 9 3 13 1 15 2
11 15 3 13 16 3 15 13 10 0 13 2
10 3 3 1 10 15 9 1 9 13 2
23 16 3 13 0 0 13 15 9 13 0 7 9 13 13 2 13 13 15 15 10 9 9 2
12 10 15 13 3 9 10 9 1 10 1 9 2
11 1 3 10 9 3 9 1 9 15 13 2
14 3 3 9 9 13 3 2 7 3 9 0 10 9 2
26 13 3 3 9 9 13 1 9 3 1 10 9 2 7 1 0 9 2 15 13 9 1 9 13 3 2
7 10 10 9 9 13 9 2
18 13 3 0 9 10 9 13 10 9 9 9 13 7 10 9 9 13 2
9 13 3 3 10 9 9 10 9 2
12 9 3 9 9 13 1 9 2 16 13 9 2
45 9 3 10 0 1 0 9 0 10 1 9 9 2 15 10 3 1 9 13 2 10 7 1 9 2 0 2 13 2 9 13 10 13 9 16 13 10 9 2 13 3 1 10 9 2
14 9 3 1 10 9 3 1 9 13 9 13 9 9 2
79 9 3 1 0 0 9 2 13 2 10 9 9 3 0 1 13 10 13 0 13 2 13 15 3 7 10 9 15 0 2 7 3 13 13 10 1 10 9 9 0 13 10 3 3 13 10 9 9 2 1 9 13 2 16 13 15 10 1 10 9 9 2 3 16 13 13 2 13 10 9 7 0 10 10 9 13 0 13 2
20 9 2 3 10 9 1 10 1 9 9 2 16 0 2 15 9 13 2 13 2
28 10 3 9 9 1 13 2 10 3 9 10 1 9 9 2 10 7 9 10 13 3 7 10 3 9 0 13 2
47 0 13 0 1 9 2 16 3 9 10 9 13 1 10 1 9 2 16 10 9 13 1 0 10 9 2 13 1 10 9 10 9 3 0 2 3 15 13 10 9 7 0 1 10 0 13 2
38 3 16 3 1 10 9 10 9 13 10 9 2 16 3 9 13 7 9 1 10 0 2 10 0 9 13 1 10 10 9 9 1 10 10 9 13 9 2
35 3 3 9 13 10 9 9 10 9 10 3 3 3 13 7 10 9 0 13 10 3 13 10 9 7 0 13 1 10 9 13 0 10 9 2
12 15 1 9 3 7 0 9 13 13 9 0 2
11 3 3 0 13 0 9 9 9 9 13 2
20 3 10 9 3 13 10 9 13 1 15 3 13 10 9 13 15 3 10 9 2
26 13 3 10 0 0 1 10 9 9 10 0 13 1 9 1 10 9 3 15 13 9 13 10 9 13 2
45 9 3 10 3 0 13 1 15 0 15 10 9 9 13 9 2 0 7 3 9 10 1 10 9 13 2 1 15 10 9 3 13 1 10 9 15 13 10 9 7 13 10 9 13 2
3 3 13 2
6 13 3 3 10 9 2
6 13 3 3 3 13 2
17 3 13 15 15 13 9 9 0 0 9 13 0 2 0 0 9 2
16 0 3 16 1 10 9 13 13 0 15 13 10 9 10 9 2
11 13 3 2 16 13 2 15 15 13 3 2
5 13 9 0 9 2
15 16 3 3 9 0 13 3 10 9 2 9 1 13 13 2
16 10 9 0 3 13 9 13 9 7 10 9 3 13 1 15 2
34 1 3 9 2 16 13 9 10 9 1 10 1 10 1 9 9 2 9 13 10 0 9 9 2 15 13 3 9 13 0 2 13 3 2
16 9 3 15 13 1 10 10 9 9 0 0 7 10 13 9 2
15 9 15 3 13 13 1 9 9 10 9 2 13 1 9 2
16 13 3 3 15 10 1 9 10 9 9 1 9 1 9 13 2
16 1 15 3 1 9 13 9 2 13 15 10 0 0 9 9 2
12 15 3 13 1 10 9 0 9 9 10 9 2
35 3 13 3 13 16 1 9 15 13 15 2 16 9 10 0 1 10 9 10 9 10 1 9 13 0 9 13 15 15 3 0 13 13 15 2
4 13 3 3 2
18 9 0 13 9 9 2 1 15 13 10 0 16 1 9 7 9 13 2
22 13 3 10 3 9 9 7 10 3 9 2 10 7 9 10 3 0 9 1 10 9 2
13 10 3 3 10 9 9 9 9 9 13 9 9 2
26 1 15 1 10 9 13 16 3 1 10 9 13 10 9 13 2 10 7 0 0 15 9 13 1 15 2
11 13 3 15 13 1 10 1 10 9 9 2
18 13 3 10 9 0 10 1 10 9 9 2 3 10 9 7 13 0 2
10 13 3 15 13 9 10 1 15 0 2
29 3 1 3 0 9 10 9 13 10 1 10 9 9 3 0 7 0 13 10 9 2 3 13 15 13 13 10 9 2
17 13 3 10 9 13 10 9 10 9 1 10 9 13 13 10 9 2
15 13 3 7 13 0 13 0 9 7 13 13 15 13 13 2
5 15 3 13 9 2
11 15 13 0 13 13 2 13 10 9 13 2
9 13 3 15 16 13 10 9 13 2
31 10 3 13 1 10 9 13 10 9 13 1 0 10 9 7 9 13 1 10 9 13 1 9 0 2 13 1 10 0 9 2
24 3 3 10 9 13 1 15 10 9 13 7 13 1 0 9 0 9 10 9 13 13 9 0 2
26 7 13 1 10 9 7 13 10 9 13 1 10 9 3 13 13 7 3 10 9 13 3 13 1 15 2
14 3 15 13 15 13 1 10 9 7 13 13 10 9 2
34 13 3 10 9 0 1 10 10 9 13 0 7 3 13 0 2 7 10 9 0 13 1 10 9 7 10 9 2 3 7 10 0 9 2
12 3 10 15 9 10 0 10 9 9 13 9 2
13 10 0 13 13 3 9 1 10 9 9 13 3 2
9 9 10 1 9 9 13 13 9 2
17 0 10 9 13 9 10 9 1 9 13 10 9 13 1 10 9 2
8 10 3 9 13 0 10 9 2
16 13 1 10 9 13 10 9 9 13 15 13 13 10 13 9 2
17 10 3 9 13 13 3 1 9 7 3 1 0 0 9 10 9 2
7 9 3 13 10 9 9 2
13 3 13 9 1 9 1 10 9 3 3 9 13 2
9 9 3 13 9 9 7 10 9 2
18 9 3 2 16 13 9 2 3 9 13 9 13 9 13 1 10 9 2
10 13 15 9 3 9 3 9 7 9 2
11 3 3 0 9 1 9 13 13 9 9 2
10 3 9 13 1 10 1 0 9 9 2
5 9 0 9 9 2
8 3 13 10 0 9 13 9 2
18 9 3 10 0 1 10 0 7 0 10 0 9 9 15 13 13 9 2
20 9 3 10 1 10 9 13 3 9 13 10 9 10 0 7 0 13 13 13 2
9 15 9 13 0 9 13 9 13 2
8 13 3 15 3 10 0 9 2
13 10 3 0 9 3 9 13 1 15 10 0 9 2
14 1 15 13 9 3 9 13 10 13 10 1 9 9 2
36 0 3 10 9 1 10 9 9 3 9 13 10 0 13 9 7 13 15 9 7 9 2 9 7 9 2 15 13 9 10 9 10 1 9 9 2
16 10 3 0 10 9 2 13 2 3 9 3 9 7 9 13 2
21 3 9 3 13 9 2 13 3 3 9 9 2 9 7 0 10 13 7 0 9 2
18 10 3 9 9 9 3 9 10 9 13 2 10 3 0 13 10 9 2
19 9 3 10 13 9 3 9 13 9 0 10 9 2 0 7 3 10 9 2
14 13 3 10 15 1 10 0 10 1 15 13 13 0 2
26 10 3 9 3 13 3 16 0 13 9 3 9 3 15 2 13 2 13 2 16 1 15 9 13 9 2
18 9 3 10 9 3 3 13 9 10 9 2 1 15 13 3 9 9 2
26 10 3 9 9 13 1 10 1 10 1 9 9 9 9 3 13 9 0 2 13 7 9 10 13 9 2
15 13 3 3 9 3 0 9 0 10 9 7 15 3 0 2
11 9 3 10 9 1 10 13 9 13 3 2
5 10 3 15 13 2
10 1 15 3 9 2 16 13 2 13 2
20 13 3 10 9 3 0 7 0 1 10 9 2 16 3 9 2 1 15 13 2
10 3 3 1 10 9 10 9 3 13 2
12 9 3 10 9 9 9 9 1 9 0 13 2
15 10 9 3 13 9 15 3 3 13 13 13 7 10 9 2
4 9 3 13 2
16 9 3 10 10 9 1 10 1 10 9 9 9 9 13 13 2
18 9 3 10 9 1 10 0 7 0 10 9 9 13 9 13 10 9 2
12 1 3 10 13 10 9 9 10 9 15 13 2
20 3 3 3 13 15 3 3 3 10 3 9 16 0 0 9 13 7 13 9 2
11 10 9 3 13 10 3 9 0 15 0 2
27 16 15 13 3 2 9 3 0 9 13 2 15 7 16 13 15 7 13 3 2 1 0 13 9 10 9 2
14 3 10 9 10 9 13 13 13 15 15 10 0 9 2
7 3 10 9 13 16 9 2
10 13 3 13 2 16 13 2 10 9 2
14 9 3 1 10 9 16 13 2 13 15 3 1 9 2
15 16 3 13 3 0 15 13 2 15 1 15 10 9 13 2
15 10 9 13 9 3 10 9 7 13 15 0 9 9 9 2
10 1 3 9 13 13 15 0 3 13 2
17 13 3 13 7 3 9 9 9 0 9 1 9 15 13 3 13 2
15 13 13 10 9 3 1 10 9 9 9 13 9 0 0 2
17 13 13 0 9 9 3 13 3 3 10 9 13 2 0 13 13 2
20 1 10 9 3 13 13 15 1 10 9 10 13 13 0 10 13 3 1 9 2
10 10 3 9 1 15 3 13 13 15 2
17 1 9 3 2 16 13 2 1 10 9 13 15 10 0 15 3 2
12 3 3 13 0 3 13 13 3 13 7 3 2
11 1 15 3 13 15 16 15 13 9 13 2
18 3 0 3 9 9 10 9 13 2 15 3 0 13 1 10 3 13 2
15 10 3 13 10 0 9 3 3 1 15 3 10 9 13 2
11 9 9 0 13 1 10 9 1 9 13 2
18 15 15 3 13 16 9 3 13 13 1 9 16 13 1 0 9 13 2
28 16 13 10 9 10 9 7 3 3 13 13 9 2 1 10 9 13 15 13 3 9 13 7 13 0 13 0 2
2 13 2
9 10 3 13 3 2 13 2 9 2
34 9 0 9 9 13 10 0 9 7 0 13 2 13 3 9 13 3 1 10 3 10 13 13 10 0 2 0 7 13 1 10 9 9 2
22 9 3 15 13 1 9 0 13 13 1 10 9 2 9 1 9 2 13 2 9 13 2
28 13 9 10 9 0 3 7 0 0 7 2 16 13 2 9 7 0 2 3 7 10 9 0 2 13 1 9 2
17 3 3 3 10 9 7 0 15 13 13 10 9 1 15 13 13 2
10 3 9 3 3 10 9 0 15 13 2
41 1 10 9 13 9 9 3 9 2 3 0 13 9 2 9 13 13 10 9 1 10 9 1 0 0 2 10 7 9 15 10 9 3 13 13 9 13 0 10 9 2
14 10 9 3 1 10 9 7 10 9 13 9 0 13 2
12 9 13 3 0 10 9 13 7 13 15 3 2
26 1 10 9 9 3 0 2 13 10 9 3 3 7 13 13 1 10 3 10 9 3 15 13 10 9 2
31 3 3 13 1 9 2 1 15 13 13 9 15 9 2 3 13 10 9 13 9 2 13 7 7 13 0 13 13 15 9 2
29 0 13 3 7 0 3 1 9 1 15 13 13 10 9 13 2 0 9 3 13 0 2 3 13 7 1 15 3 2
6 3 13 13 10 9 2
21 1 15 13 0 13 9 2 13 7 2 16 9 3 3 7 0 15 13 10 9 2
10 10 9 3 13 0 2 13 2 9 2
10 13 2 13 2 7 13 2 16 13 2
32 9 13 3 10 9 1 9 13 1 9 0 0 0 3 1 9 2 10 0 13 9 1 15 9 3 0 9 7 0 9 0 2
18 3 15 1 0 0 9 0 9 13 0 10 3 1 10 9 3 13 2
7 3 3 15 13 15 13 2
6 3 3 3 15 13 2
16 9 13 10 0 3 9 13 1 9 0 9 7 9 13 13 2
5 10 3 13 13 2
10 15 3 0 2 16 3 10 13 13 2
14 10 9 13 1 9 0 0 9 0 0 13 1 9 2
16 3 16 9 13 13 2 13 10 9 10 9 13 13 13 9 2
5 10 9 3 13 2
13 16 3 9 9 15 2 13 2 13 0 2 13 2
7 10 13 3 13 15 15 2
17 10 10 9 9 13 10 9 9 0 13 3 0 13 3 0 13 2
13 13 3 9 2 16 10 0 3 13 9 3 9 2
13 13 3 1 10 9 13 0 9 0 7 13 9 2
19 13 3 15 13 15 3 2 13 2 0 16 15 10 9 2 0 0 13 2
14 9 13 10 9 9 13 9 10 1 10 9 3 13 2
14 15 3 3 10 9 3 13 1 9 1 10 9 9 2
6 13 3 13 3 15 2
7 13 3 3 13 1 0 2
10 3 13 15 0 9 13 1 10 0 2
5 3 10 9 13 2
6 9 13 9 10 0 2
11 3 13 15 9 0 10 9 0 2 13 2
9 3 0 0 0 13 13 9 0 2
16 13 3 3 15 2 13 2 16 3 15 13 2 7 15 13 2
33 9 13 10 9 2 9 0 15 3 13 2 9 7 10 0 13 2 7 0 13 3 2 16 13 2 15 2 13 1 10 13 9 2
18 9 2 13 2 16 3 0 10 0 13 2 1 0 0 13 13 3 2
10 1 3 15 13 10 1 10 9 13 2
24 10 3 0 15 9 0 9 13 9 2 1 15 13 0 3 13 2 0 9 13 9 3 13 2
6 15 3 13 9 9 2
25 10 3 9 13 3 2 16 3 0 13 2 9 10 9 2 16 7 9 10 0 1 10 9 13 2
20 1 9 3 3 15 13 3 13 1 10 9 13 7 15 0 13 1 10 9 2
22 13 3 10 9 13 10 9 15 10 9 2 10 3 15 3 2 13 2 3 13 13 2
10 3 3 13 0 1 10 9 10 9 2
17 3 0 3 9 0 13 1 15 2 9 13 7 10 9 9 13 2
8 3 3 0 1 10 9 13 2
12 9 3 9 1 9 9 9 3 3 0 13 2
8 9 3 0 9 13 10 9 2
8 15 3 13 2 16 3 13 2
8 10 9 3 2 13 2 13 2
21 9 3 10 9 13 7 1 9 0 13 2 10 9 2 13 2 1 10 9 13 2
21 13 3 15 9 1 9 0 7 13 16 9 2 0 3 2 13 2 3 0 9 2
10 3 3 9 10 9 13 2 7 9 2
18 9 3 0 13 15 16 3 9 2 13 2 13 2 13 3 15 13 2
14 13 3 10 3 0 13 13 2 10 7 9 0 13 2
28 10 3 13 1 15 13 1 9 7 10 9 1 10 13 1 10 9 13 10 9 2 10 9 13 9 13 13 2
23 1 3 9 0 13 16 13 1 9 3 3 2 13 2 1 10 0 9 3 13 10 3 2
10 15 3 13 1 0 2 1 9 13 2
13 15 3 3 2 13 10 9 2 15 3 13 13 2
21 9 3 10 9 13 2 13 10 9 2 9 0 13 0 1 9 2 3 0 13 2
9 15 3 13 15 1 0 9 13 2
10 3 10 9 2 13 2 7 10 9 2
27 9 3 10 9 2 9 10 9 9 3 13 1 0 9 2 3 3 15 2 13 2 15 13 3 9 13 2
14 13 3 15 1 10 3 9 13 2 13 2 16 13 2
4 15 13 9 2
11 0 3 10 9 9 15 13 3 2 13 2
21 13 3 9 7 9 2 16 15 13 15 13 10 9 2 9 13 10 9 3 13 2
11 0 3 13 3 10 9 7 3 0 13 2
26 15 3 9 0 13 2 1 15 13 10 9 1 15 7 10 9 13 2 1 9 10 10 15 13 9 2
16 13 3 15 9 1 10 0 9 10 9 7 9 15 0 13 2
13 0 10 9 0 13 7 0 2 9 0 0 0 2
8 9 3 10 13 9 9 13 2
2 13 2
15 9 10 9 13 7 13 1 10 9 9 13 9 13 13 2
6 13 3 13 9 15 2
11 10 3 13 2 13 2 7 10 3 13 2
27 9 9 0 15 9 1 0 9 13 7 13 13 15 13 2 15 7 13 2 13 2 13 2 0 10 0 2
21 9 13 1 9 2 13 1 10 9 9 7 10 9 15 15 3 13 2 0 13 2
16 16 3 13 10 0 15 13 15 13 2 10 0 15 13 13 2
10 1 9 10 0 9 9 13 13 13 2
6 10 3 3 13 13 2
3 9 13 2
15 9 1 9 13 9 2 16 15 15 13 3 13 2 13 2
14 9 13 3 9 13 9 13 2 13 2 7 15 13 2
16 13 3 1 0 9 1 0 9 10 9 13 2 13 16 13 2
15 9 3 0 13 1 15 7 13 0 13 2 1 9 13 2
13 13 3 10 9 13 15 2 13 2 7 0 13 2
11 0 3 0 9 13 15 13 9 13 9 2
12 9 3 3 1 10 1 9 9 13 7 9 2
28 13 3 15 9 1 9 7 1 9 2 1 9 2 1 13 2 1 9 2 3 9 1 9 7 9 1 9 2
23 1 3 10 9 9 13 1 10 1 10 3 9 16 9 13 2 16 1 10 9 13 13 2
8 9 3 1 10 1 9 13 2
10 3 3 10 9 13 10 0 9 13 2
14 15 9 13 2 16 0 7 0 13 10 9 0 13 2
15 9 3 1 10 1 9 9 13 9 13 1 10 0 9 2
8 0 16 15 13 10 9 13 2
24 1 15 13 9 1 10 1 10 0 9 2 16 1 10 10 9 9 10 9 13 10 9 3 2
12 10 0 3 13 3 9 1 10 1 9 9 2
17 3 3 13 9 10 9 15 10 9 3 0 9 13 7 9 13 2
6 9 10 9 15 13 2
10 13 3 3 15 9 7 3 9 9 2
16 9 3 1 10 1 9 2 16 3 0 10 9 2 15 13 2
21 9 3 3 13 13 3 0 13 3 9 3 9 3 9 3 9 3 9 7 9 2
9 3 3 13 13 1 10 9 9 2
26 3 3 13 1 15 9 13 9 2 1 7 9 3 0 9 13 2 16 13 2 9 7 9 9 13 2
11 3 10 10 1 9 3 9 13 13 15 2
28 1 3 10 1 9 0 10 9 2 16 0 10 9 2 3 9 10 9 13 2 7 1 10 1 9 9 9 2
6 0 3 13 15 9 2
41 10 3 0 13 9 2 16 9 13 1 10 1 9 2 9 15 13 13 3 16 13 13 7 13 7 16 15 13 10 9 9 13 13 15 0 9 2 0 7 15 2
14 3 9 1 10 1 9 9 9 13 3 13 10 9 2
14 15 3 16 9 13 13 2 1 10 9 10 9 13 2
25 16 3 9 13 10 9 2 16 3 1 9 13 10 9 7 3 9 13 1 15 2 0 13 9 2
13 3 10 3 9 1 9 16 13 10 9 13 3 2
18 3 3 2 16 15 9 13 2 9 9 13 0 13 9 13 0 9 2
9 13 10 9 3 9 1 9 3 2
9 9 3 1 9 13 3 13 9 2
31 9 3 1 10 1 9 9 2 13 2 13 10 9 2 16 9 3 0 13 7 13 9 7 9 0 2 13 7 13 0 2
15 13 3 9 10 9 9 2 10 10 9 13 1 9 9 2
12 3 9 3 10 9 9 13 1 10 1 9 2
17 1 15 0 13 3 13 9 3 13 10 9 2 9 0 9 13 2
25 13 3 10 0 13 9 3 0 10 13 2 7 3 10 0 9 2 16 13 9 1 10 1 9 2
19 3 10 0 9 1 9 13 13 9 15 13 2 13 2 7 1 9 9 2
8 9 3 1 9 0 13 9 2
14 9 2 9 2 9 2 9 2 7 9 13 0 3 2
16 3 9 3 3 13 9 0 2 10 7 9 0 9 0 0 2
10 9 3 3 13 15 16 10 0 13 2
15 3 9 3 13 13 13 2 9 7 3 9 13 7 9 2
9 9 3 3 9 7 9 3 13 2
5 1 3 9 13 2
5 9 3 3 13 2
35 15 13 1 0 9 10 9 3 15 15 15 10 9 2 13 2 10 3 1 10 0 13 3 10 10 9 9 13 2 16 3 10 9 13 2
11 15 3 10 0 10 9 9 13 1 15 2
7 1 0 3 9 13 9 2
8 3 0 3 13 10 0 9 2
18 15 0 9 0 13 13 3 10 3 15 1 9 13 2 0 9 13 2
11 3 15 3 10 9 13 0 2 0 13 2
14 0 3 10 9 3 9 13 13 10 1 9 0 13 2
23 10 3 3 16 13 13 13 13 2 0 3 10 0 13 1 10 9 2 9 7 3 3 2
25 9 3 10 9 3 9 13 10 9 13 1 10 9 13 7 13 10 9 13 3 15 1 0 9 2
19 13 3 15 10 9 16 1 9 9 1 10 9 13 2 3 13 2 13 2
13 15 3 15 13 1 9 1 3 0 9 0 13 2
17 10 3 15 3 9 13 1 9 10 9 2 16 13 9 1 9 2
21 16 3 0 13 7 9 0 9 0 13 13 15 0 15 2 13 2 13 10 9 2
9 3 3 3 13 13 13 10 9 2
22 3 3 13 10 9 0 16 3 10 9 13 1 15 13 10 9 10 9 7 10 9 2
22 13 3 3 10 9 10 9 0 0 13 9 2 3 13 0 7 9 7 3 15 13 2
14 9 3 1 9 12 9 2 13 15 1 9 10 9 2
22 3 13 1 9 16 15 3 15 0 9 13 2 10 7 9 9 10 9 13 2 13 2
4 3 3 13 2
4 3 15 13 2
11 3 3 3 9 13 0 13 15 0 13 2
13 9 3 1 9 7 9 0 15 13 13 1 15 2
9 13 3 3 10 9 0 7 15 2
9 3 3 13 3 2 13 7 0 2
5 9 3 0 9 2
30 3 3 9 13 2 13 13 15 1 0 9 1 9 2 13 0 9 9 2 1 9 7 9 0 9 13 1 9 9 2
8 15 13 9 2 13 7 9 2
7 13 3 1 0 0 9 2
12 13 3 10 13 15 1 9 13 1 10 9 2
37 9 3 10 9 3 1 9 10 9 13 9 7 13 15 1 9 2 16 13 9 1 10 1 9 0 2 9 13 10 13 13 1 10 10 9 9 2
12 10 3 0 15 9 3 9 10 0 9 13 2
15 9 13 10 1 9 9 2 15 3 1 9 0 13 9 2
41 9 3 10 0 2 16 13 9 1 0 0 2 3 1 9 2 3 10 0 7 10 9 10 0 13 2 3 0 9 9 7 0 9 13 2 3 13 0 10 9 2
9 13 3 0 9 1 0 3 0 2
34 15 3 10 10 9 9 13 2 16 9 10 0 13 2 1 10 0 15 9 13 7 13 15 2 1 10 13 1 9 3 9 7 9 2
41 9 3 10 0 13 13 0 9 3 10 9 13 7 13 1 15 13 10 9 2 3 13 3 15 9 9 13 1 15 0 13 16 16 1 10 9 7 10 9 13 2
28 3 9 3 9 10 9 3 13 2 7 0 13 9 2 7 13 9 13 10 9 15 10 9 10 10 9 13 2
22 9 3 10 9 9 2 15 13 0 1 9 10 1 9 13 2 13 13 9 10 0 2
9 15 9 10 10 9 9 9 13 2
21 3 10 9 2 16 9 0 2 3 13 10 9 13 2 16 13 3 13 10 9 2
8 9 3 13 15 13 1 9 2
22 16 9 3 13 10 9 2 15 13 15 2 10 9 3 13 15 0 1 15 13 9 2
6 3 3 13 15 3 2
6 1 15 10 9 13 2
12 13 3 16 3 13 10 9 9 1 9 3 2
6 13 2 13 10 9 2
18 13 3 3 0 9 13 10 3 2 16 3 13 10 10 0 9 9 2
7 9 3 1 9 13 3 2
29 9 3 10 0 0 3 15 2 3 3 7 1 10 9 13 10 9 2 16 15 13 10 13 15 1 10 9 9 2
53 9 3 10 9 1 10 0 9 10 9 13 9 9 10 0 9 13 2 7 15 3 1 9 13 2 1 9 3 9 2 9 7 1 9 2 15 0 13 9 13 13 2 0 7 3 0 15 13 2 16 9 13 2
24 1 3 10 1 9 9 9 13 13 10 9 7 3 10 9 13 10 13 9 1 10 9 13 2
7 13 3 10 9 1 9 2
9 13 3 1 9 10 1 9 13 2
14 3 13 10 9 3 3 13 0 9 2 16 13 9 2
12 13 3 3 3 10 9 0 1 10 3 13 2
8 3 3 3 13 15 13 0 2
11 0 3 9 13 7 10 0 3 13 9 2
24 10 3 10 0 9 7 10 10 0 1 9 10 9 0 13 9 7 13 10 9 13 10 9 2
9 3 1 15 9 10 9 9 13 2
27 3 9 3 10 9 13 15 10 0 9 1 15 13 7 1 10 10 9 9 10 1 10 9 10 9 13 2
18 9 15 13 13 9 2 1 0 13 0 9 2 9 9 15 13 15 2
9 9 3 13 3 13 2 7 13 2
10 10 3 13 10 9 13 15 1 9 2
16 0 3 10 9 10 9 9 13 13 1 9 0 1 9 0 2
5 13 3 15 9 2
13 15 3 13 9 10 0 13 10 10 9 9 9 2
27 9 3 1 0 13 10 3 1 10 9 13 13 9 13 1 10 13 7 13 10 13 15 2 10 7 0 2
33 13 3 3 10 9 7 13 13 10 9 2 16 13 9 16 9 3 13 2 13 7 9 10 9 2 16 13 9 1 10 1 9 2
18 13 3 10 9 9 9 13 10 9 2 16 3 9 10 0 9 9 2
14 9 3 1 10 1 9 10 0 13 15 13 9 9 2
17 3 13 3 16 10 13 1 15 9 9 9 10 9 9 13 13 2
11 9 3 10 0 1 9 15 13 1 15 2
9 9 3 15 13 0 0 10 9 2
14 3 3 16 0 10 3 9 13 2 10 3 9 13 2
26 13 13 10 9 0 9 10 9 13 1 10 9 2 7 10 9 1 9 13 1 9 13 10 9 3 2
13 13 3 16 3 9 10 9 1 9 9 13 9 2
10 15 13 3 1 10 9 13 9 13 2
23 3 9 3 10 9 9 9 13 9 9 9 2 16 13 9 10 0 1 10 10 9 9 2
6 13 3 10 9 13 2
26 13 3 9 0 0 3 13 9 7 9 2 10 7 13 0 9 2 15 9 3 13 2 9 7 13 2
9 15 3 13 1 10 1 9 13 2
10 10 3 9 13 13 1 0 9 3 2
21 1 3 9 13 10 9 2 16 13 9 2 9 13 10 9 7 10 9 9 13 2
24 16 3 0 13 10 9 13 10 9 2 10 0 15 9 9 13 1 15 15 13 9 3 13 2
7 16 10 9 1 9 13 2
21 3 3 3 9 10 10 9 0 9 13 13 7 9 2 16 9 13 1 10 9 2
14 9 3 1 10 1 9 10 9 10 9 13 13 13 2
16 13 3 3 10 9 9 10 9 2 15 13 9 9 10 9 2
16 3 3 9 10 9 10 9 9 13 3 15 9 9 10 9 2
23 10 3 9 0 9 1 10 1 9 0 2 16 0 10 9 2 13 13 13 9 13 3 2
23 13 3 9 9 9 9 2 15 9 9 13 2 10 3 9 0 2 10 9 7 13 13 2
8 13 15 3 9 1 10 9 2
8 13 3 9 3 1 15 9 2
6 0 9 7 3 9 2
27 9 3 1 10 1 9 13 13 10 9 10 9 13 9 10 9 1 10 9 2 1 15 3 13 15 9 2
23 3 9 3 1 10 1 9 2 16 0 10 9 2 13 15 2 13 3 0 9 1 15 2
23 9 3 3 13 13 3 0 13 3 9 3 9 3 9 3 9 3 9 3 9 7 9 2
11 9 3 10 9 3 13 1 9 13 9 2
31 15 3 1 10 1 9 9 13 10 9 1 10 9 3 1 15 9 13 1 10 9 2 7 9 13 10 13 10 9 13 2
13 0 3 13 10 9 1 10 0 2 16 13 9 2
16 9 3 0 13 9 7 1 15 13 1 9 13 15 10 9 2
13 13 3 3 1 9 3 1 0 7 1 9 0 2
8 3 3 10 9 3 15 13 2
9 15 3 3 15 1 9 13 13 2
15 13 3 3 1 10 9 13 0 9 9 2 3 9 13 2
28 9 3 10 0 9 9 13 10 9 10 10 9 0 7 1 10 9 9 13 10 9 2 16 13 9 10 9 2
35 9 3 10 10 1 9 13 9 9 13 10 0 9 9 13 10 9 2 15 1 9 1 9 13 10 9 7 13 1 10 10 9 9 13 2
24 3 13 15 15 10 9 13 10 9 10 9 10 9 13 10 9 10 9 2 16 3 15 13 2
17 9 3 10 9 10 0 9 13 3 0 9 13 10 1 10 9 2
22 1 15 15 3 13 13 1 9 2 10 7 13 2 16 13 9 1 10 0 13 15 2
45 10 0 10 9 9 2 13 1 15 10 0 2 9 3 13 10 1 9 10 0 13 9 2 9 7 13 0 9 2 13 16 13 13 10 9 10 9 13 10 9 2 13 10 9 2
15 10 3 13 7 13 13 1 15 13 0 9 13 1 9 2
7 3 13 9 13 1 9 2
21 13 3 10 9 10 13 1 10 9 13 10 9 2 15 10 13 0 1 9 13 2
21 10 3 9 13 2 16 13 10 13 15 9 2 13 1 10 9 3 9 15 13 2
13 10 3 0 9 3 1 9 13 1 10 0 3 2
7 9 9 10 9 9 13 2
13 3 13 15 15 13 3 1 10 0 10 9 13 2
20 9 3 10 9 9 10 0 9 13 3 1 15 3 9 13 2 16 13 9 2
5 13 3 3 0 2
16 9 3 10 9 9 13 9 10 9 2 9 7 10 9 9 2
27 10 3 9 13 9 9 10 0 3 9 10 9 7 9 10 9 2 15 13 9 3 9 2 9 7 9 2
18 10 3 9 13 9 1 9 2 9 13 0 2 9 7 9 10 9 2
27 15 3 10 10 9 9 9 10 0 9 13 16 0 9 13 9 10 9 2 16 13 9 1 10 1 9 2
9 15 3 1 9 10 9 15 13 2
18 9 10 9 13 1 10 9 3 13 7 13 1 10 0 10 9 13 2
43 3 15 3 13 15 7 16 9 10 9 0 1 10 9 10 1 10 9 3 13 9 13 2 0 13 1 0 10 9 9 3 13 2 3 15 13 10 9 2 7 10 9 2
9 0 3 9 13 3 10 0 9 2
14 15 0 13 13 0 0 9 2 9 13 9 10 0 2
38 9 3 13 10 9 1 15 10 9 13 10 9 10 9 7 13 13 10 9 10 1 15 9 2 16 0 13 2 13 10 9 9 10 9 9 0 13 2
12 10 3 3 13 13 10 9 3 13 15 13 2
11 3 10 9 10 9 13 10 9 2 13 2
16 9 3 10 0 13 10 9 10 3 13 15 2 10 7 13 2
11 3 10 0 0 13 2 3 13 10 9 2
18 1 15 9 13 2 16 13 9 1 10 1 9 2 9 13 10 9 2
9 13 3 3 9 1 15 1 15 2
11 9 0 0 13 9 2 0 9 9 9 2
10 16 3 3 9 10 9 13 9 0 2
3 13 3 2
19 9 3 9 13 7 0 15 13 1 10 9 2 13 9 3 15 13 0 2
23 9 3 10 9 10 10 9 0 9 13 7 13 1 9 13 9 0 1 15 13 9 13 2
6 3 13 0 9 13 2
32 13 3 15 1 10 9 2 16 13 9 1 10 0 7 0 10 9 2 9 10 0 9 0 3 0 9 7 9 13 10 9 2
11 9 3 1 10 1 10 1 9 9 13 2
19 15 3 13 15 3 1 10 9 9 13 1 10 1 9 10 9 9 13 2
35 3 3 3 13 3 3 13 10 0 10 10 9 13 9 3 10 9 2 13 1 10 9 0 13 9 0 3 0 3 3 15 13 10 9 2
15 3 3 16 13 9 10 9 13 2 0 13 9 13 15 2
13 9 3 1 10 1 9 9 10 9 13 9 13 2
15 13 3 7 13 3 1 10 1 9 0 9 9 13 13 2
11 1 0 3 9 16 0 0 9 13 15 2
46 15 3 0 13 0 9 0 10 13 13 2 15 13 10 0 13 15 13 9 7 9 13 7 13 10 9 7 10 9 0 9 2 3 10 3 1 9 9 13 7 10 0 9 13 13 2
7 13 15 3 9 1 0 2
8 9 13 9 2 16 3 13 2
7 10 9 13 7 10 9 2
8 13 3 15 3 9 1 9 2
34 1 3 10 9 9 10 9 9 13 3 0 9 2 16 10 9 13 2 13 13 10 9 3 13 15 2 16 3 15 13 3 10 9 2
19 13 3 9 0 10 9 1 9 10 9 2 3 3 15 7 15 13 13 2
36 13 3 15 13 1 10 9 10 1 9 7 13 1 10 9 13 3 9 13 7 10 0 9 13 2 15 13 13 10 0 9 7 10 15 13 2
34 13 3 15 3 10 10 9 10 0 9 13 2 15 13 9 13 1 10 9 9 2 16 9 13 10 0 7 0 7 3 0 10 9 2
13 13 3 10 9 3 13 10 9 1 9 7 13 2
29 3 10 3 9 3 13 13 2 10 7 9 3 13 1 15 7 10 9 9 13 10 9 13 1 9 2 13 3 2
13 13 3 2 3 3 10 9 13 0 2 9 0 2
20 1 0 3 0 9 10 0 9 2 15 3 9 13 13 1 10 9 15 9 2
19 3 3 10 0 0 9 13 15 3 13 13 16 13 10 9 3 10 9 2
7 9 3 3 13 10 9 2
10 1 3 10 3 10 9 13 15 13 2
17 13 3 15 13 0 13 3 2 9 9 0 9 13 7 13 15 2
10 16 3 13 0 13 9 2 0 13 2
15 3 3 10 9 0 7 10 9 13 2 9 7 3 3 2
17 3 3 13 9 10 9 15 10 9 3 0 9 13 7 9 13 2
6 9 10 9 0 13 2
9 13 3 3 15 9 3 9 9 2
12 0 3 9 7 1 9 13 13 3 10 9 2
18 1 3 10 9 0 13 9 9 2 3 3 1 10 9 3 15 13 2
4 13 3 15 2
13 0 3 13 0 3 7 13 9 10 0 13 9 2
16 9 0 0 2 15 9 3 13 13 16 13 9 9 0 9 2
12 3 9 3 13 1 10 9 7 15 9 0 2
16 13 3 3 10 9 2 16 10 9 13 2 0 13 10 9 2
24 3 10 1 9 3 10 9 0 9 9 10 0 9 13 0 13 2 16 13 9 1 0 9 2
25 9 3 10 9 3 0 13 9 2 7 3 9 1 7 1 9 0 13 2 13 7 9 10 9 2
23 9 3 10 0 9 3 15 0 2 10 9 1 10 9 13 2 16 10 10 0 13 13 2
15 15 3 13 1 10 1 9 10 9 15 13 13 10 9 2
34 9 3 10 9 9 13 10 13 9 9 2 10 13 9 7 0 1 10 3 0 9 13 1 10 13 2 16 13 9 1 10 1 9 2
14 13 3 3 10 9 9 9 7 10 9 10 0 9 2
23 1 3 15 9 15 13 13 0 0 9 2 15 1 10 0 9 13 0 2 3 3 13 2
27 13 3 0 7 0 9 2 3 9 0 13 1 9 9 13 2 9 7 1 0 13 9 1 0 13 9 2
13 3 13 1 9 0 13 9 2 0 7 13 9 2
31 9 3 0 1 9 13 13 2 7 0 9 13 9 2 1 9 3 9 13 2 1 9 7 9 0 2 0 9 13 9 2
11 3 13 0 13 9 9 0 9 13 9 2
18 10 3 0 9 9 1 9 9 0 13 9 2 0 9 9 13 9 2
7 0 3 13 3 1 9 2
21 3 10 3 9 13 0 0 13 2 0 7 9 13 9 13 2 1 0 9 13 2
14 15 1 0 13 0 13 9 2 0 1 0 13 9 2
15 13 3 9 3 9 3 9 9 7 9 2 9 13 9 2
19 9 3 10 0 15 13 0 13 9 7 0 9 1 0 2 13 3 9 2
11 0 3 1 3 9 13 9 13 1 9 2
15 13 3 9 10 3 0 7 9 0 2 13 0 13 9 2
13 0 3 9 9 1 3 9 13 9 9 13 9 2
17 9 3 13 1 0 13 9 13 2 13 7 13 13 0 1 9 2
11 9 3 13 9 0 2 1 0 13 9 2
15 0 9 3 2 0 13 9 2 9 13 0 9 2 13 2
11 10 3 9 9 13 9 0 13 9 9 2
12 3 3 10 10 0 13 9 13 0 3 9 2
19 13 3 3 3 13 9 2 3 7 15 0 9 13 9 2 9 1 0 2
10 10 3 0 13 9 3 0 9 3 2
25 9 3 0 9 9 9 13 1 0 13 9 9 7 10 9 9 9 7 15 3 0 9 13 9 2
26 13 3 3 0 10 3 13 9 7 0 9 13 1 9 0 1 9 1 0 13 9 0 3 13 9 2
12 3 9 0 13 9 13 2 13 7 9 9 2
27 13 3 3 10 9 2 15 9 9 0 0 13 1 9 9 13 0 2 1 0 9 9 7 0 13 9 2
41 3 3 3 0 0 9 13 9 2 0 13 9 2 15 15 1 0 9 13 9 7 0 9 9 13 9 2 3 15 0 9 13 9 13 2 0 7 13 1 9 2
24 0 3 0 9 13 9 9 2 9 0 9 13 2 7 9 0 13 9 0 1 9 0 13 2
17 0 3 13 15 0 13 9 9 13 9 1 9 9 13 9 9 2
13 1 3 0 9 0 13 9 2 9 1 9 13 2
27 9 3 0 1 9 13 9 0 2 16 0 9 13 0 9 2 0 7 13 9 13 2 0 7 13 9 2
27 1 15 10 9 13 13 13 9 7 9 2 10 3 1 9 7 9 13 2 10 7 1 9 10 9 9 2
17 9 3 1 10 1 9 3 13 15 13 1 15 13 1 9 15 2
12 9 3 15 0 13 9 9 9 0 13 13 2
10 3 10 9 3 1 15 15 13 13 2
11 15 3 13 13 10 9 1 0 10 9 2
15 3 3 9 10 9 13 1 9 9 9 9 9 7 9 2
7 9 13 10 9 1 9 2
14 0 3 13 9 10 3 10 0 9 13 2 9 0 2
25 13 3 0 13 9 7 0 10 9 2 3 3 7 10 9 10 0 2 10 9 1 9 13 13 2
14 15 3 3 13 7 13 3 0 13 7 1 0 13 2
8 15 13 15 15 7 0 9 2
13 13 3 10 0 9 13 9 13 1 9 9 1 2
23 16 3 13 1 15 0 2 13 15 0 7 13 3 2 1 15 0 13 3 7 13 9 2
14 3 10 0 3 9 1 10 9 0 13 10 9 13 2
14 13 3 0 9 13 9 2 9 7 9 13 9 13 2
9 9 3 1 0 9 13 13 9 2
11 10 3 13 9 9 3 9 7 9 0 2
9 9 9 3 1 13 9 0 13 2
5 10 3 15 0 2
8 1 9 0 3 10 9 13 2
27 0 3 9 9 7 0 13 3 9 13 9 2 10 3 13 0 13 9 2 13 7 0 13 1 15 0 2
17 3 3 10 9 10 3 13 7 10 0 9 15 7 9 13 15 2
22 15 3 9 3 0 13 9 2 3 0 13 7 0 0 13 3 13 10 0 9 9 2
12 15 10 0 13 3 3 9 0 13 1 9 2
10 13 3 1 15 3 10 0 9 15 2
44 3 3 15 9 13 7 13 2 1 3 3 9 9 13 9 9 13 2 9 1 0 13 2 9 3 9 0 9 13 2 9 7 10 9 9 1 9 13 9 0 9 9 9 2
10 9 15 3 9 3 0 13 9 13 2
24 13 3 3 16 10 9 3 3 13 2 9 3 13 2 13 7 3 1 10 9 10 9 13 2
6 13 3 3 1 15 2
11 0 0 9 13 9 0 9 10 0 9 2
15 3 9 3 3 3 0 13 13 3 0 10 9 10 9 2
10 15 3 3 10 0 13 0 7 9 2
8 3 3 9 15 13 10 9 2
8 3 13 10 15 0 10 9 2
9 3 10 9 3 9 13 7 13 2
20 3 1 9 13 0 9 2 13 1 9 0 9 0 0 3 3 13 0 9 2
9 3 9 3 3 3 13 0 13 2
9 13 3 13 7 9 13 1 9 2
9 3 3 10 9 1 10 9 13 2
25 9 13 2 9 3 13 2 9 7 13 2 7 3 13 13 16 15 15 13 1 10 0 0 9 2
8 16 13 13 2 3 13 13 2
17 13 3 3 10 0 9 10 9 2 15 13 15 9 2 15 13 2
42 10 3 9 9 3 9 13 13 15 3 9 13 2 1 0 7 9 13 9 9 0 9 2 1 7 9 13 0 3 1 9 13 3 7 0 9 9 13 0 9 13 2
20 3 15 9 3 9 3 13 9 0 9 13 2 16 3 13 9 0 1 9 2
12 3 3 10 0 9 10 1 10 0 13 0 2
17 9 3 2 16 13 2 7 10 1 9 9 1 10 9 3 13 2
15 9 3 1 10 0 3 10 9 13 13 10 9 7 9 2
27 10 3 13 9 1 15 13 13 10 9 1 10 9 7 10 9 13 9 13 2 1 15 3 9 0 13 2
39 3 10 1 9 3 9 13 9 2 3 1 9 9 13 2 9 13 7 10 9 15 9 13 9 2 16 9 7 9 13 10 0 1 10 1 10 9 9 2
27 9 3 10 0 0 13 13 10 10 9 9 16 3 10 10 0 9 7 10 1 15 0 13 0 9 13 2
17 9 3 13 9 0 3 13 3 13 16 0 9 13 1 10 9 2
34 9 3 15 13 10 13 3 1 9 0 9 7 10 1 10 9 9 1 9 7 9 13 2 1 9 7 1 9 10 9 7 9 9 2
16 9 3 13 10 9 2 16 13 9 10 0 1 10 1 0 2
24 3 3 10 9 13 1 15 9 10 9 10 9 13 2 15 13 10 13 10 9 16 15 13 2
29 13 3 3 1 10 1 10 9 2 13 10 0 10 0 2 3 0 7 9 10 0 13 10 13 0 1 10 9 2
6 13 3 10 9 15 2
11 0 3 13 3 10 1 9 10 9 13 2
35 15 9 13 0 2 9 13 10 9 0 9 1 0 9 0 2 16 13 9 10 0 1 0 1 9 2 0 15 13 10 9 1 10 13 2
13 15 3 13 10 9 9 2 9 7 13 10 0 2
16 13 3 15 3 10 9 3 9 10 0 9 13 3 7 13 2
7 3 13 9 10 0 9 2
21 1 3 9 2 16 9 13 10 0 2 1 10 9 10 9 16 0 9 13 13 2
7 3 3 10 9 9 13 2
21 3 13 3 16 10 1 9 7 9 13 13 9 10 9 1 10 1 10 9 9 2
29 15 3 13 10 0 9 13 9 13 1 9 7 13 10 9 0 9 2 15 3 13 7 13 1 9 1 9 13 2
11 9 3 10 0 1 9 13 13 10 9 2
13 3 9 3 10 0 3 0 13 9 0 3 13 2
11 9 3 1 9 13 9 13 10 9 13 2
9 9 3 13 3 3 9 10 9 2
37 9 3 1 10 1 10 1 9 9 9 10 9 3 15 13 13 16 1 9 9 0 13 15 13 2 7 10 9 13 1 9 3 13 3 13 13 2
20 9 3 1 0 9 9 2 13 2 10 9 9 0 13 7 13 3 1 15 2
19 16 3 9 1 9 15 13 13 9 2 10 9 13 10 9 13 10 9 2
15 3 15 3 2 13 2 3 3 3 15 13 16 15 13 2
38 0 3 13 10 9 9 7 10 9 9 0 13 3 0 13 2 7 3 15 13 13 16 13 0 2 7 3 3 9 1 10 9 13 0 15 13 13 2
17 3 3 9 15 13 13 10 9 10 9 13 3 15 13 7 9 2
10 9 3 10 0 9 9 13 13 9 2
17 9 3 1 10 9 9 13 9 13 0 2 3 7 10 9 13 2
12 9 3 9 13 9 2 13 1 10 9 13 2
12 9 3 10 0 1 9 9 13 9 9 13 2
22 9 3 10 9 9 13 9 10 9 2 1 15 9 10 0 1 10 9 9 13 3 2
7 9 10 9 13 10 9 2
29 3 3 3 1 9 13 1 0 9 7 13 1 10 9 13 15 13 15 1 9 10 9 2 15 3 13 10 9 2
10 9 3 13 10 9 2 16 9 9 2
11 9 3 10 9 1 10 13 9 13 3 2
5 13 15 3 13 2
13 13 3 15 3 3 3 13 15 7 13 10 9 2
11 3 0 3 13 10 9 13 1 10 13 2
6 3 3 9 13 13 2
8 13 3 1 0 9 9 9 2
14 3 3 3 3 3 13 9 0 13 10 9 10 0 2
19 16 3 10 9 9 0 13 0 10 9 10 9 2 3 3 3 0 13 2
11 3 3 13 10 0 10 3 0 13 13 2
18 0 1 9 13 9 9 2 7 10 9 2 13 2 10 13 9 9 2
20 0 3 16 13 10 9 10 10 9 9 7 3 0 2 0 3 13 10 9 2
19 16 3 15 1 0 9 13 10 9 2 9 9 7 3 9 0 13 3 2
18 13 3 10 3 9 13 10 9 2 10 7 3 10 9 10 9 13 2
17 13 3 15 1 10 9 9 10 0 9 13 2 16 13 10 9 2
25 13 3 15 10 9 1 10 9 3 10 9 10 15 9 13 2 16 3 10 9 10 9 0 13 2
12 16 3 13 15 3 3 2 13 10 9 13 2
12 3 9 13 3 15 13 2 13 7 3 13 2
10 3 3 3 1 0 15 13 10 9 2
12 15 0 3 13 3 7 13 16 13 7 13 2
18 10 3 0 3 0 7 0 13 2 7 16 3 0 9 10 0 9 2
20 3 9 3 10 0 1 10 0 9 13 16 9 0 9 1 9 13 13 15 2
19 10 3 3 9 10 0 9 1 10 9 13 2 10 7 10 9 9 13 2
20 1 3 10 9 10 9 13 10 10 9 9 13 2 13 10 9 10 0 9 2
33 0 3 13 13 10 13 9 13 7 13 10 13 3 15 3 13 0 13 10 9 2 7 15 13 2 10 7 9 1 10 9 13 2
27 3 10 9 13 13 1 15 10 0 9 2 13 10 1 10 9 7 9 9 2 7 15 1 9 15 13 2
7 15 3 13 0 9 13 2
39 9 3 1 10 1 10 13 1 9 9 9 13 10 9 9 10 0 9 13 13 1 10 9 7 3 15 13 2 13 7 10 9 0 1 9 1 10 9 2
19 1 3 10 0 9 9 0 3 13 13 9 10 9 9 2 9 7 9 2
18 15 3 2 13 2 3 13 10 9 13 2 16 3 1 10 9 13 2
16 0 10 9 1 9 13 1 10 9 7 3 13 15 13 13 2
51 0 10 9 1 9 1 15 1 10 9 9 2 13 9 1 10 9 10 0 15 13 9 1 10 9 10 9 9 2 16 13 1 9 13 2 16 0 13 1 10 9 13 2 0 13 10 9 13 1 15 2
15 3 10 9 0 13 10 9 13 1 10 10 9 9 13 2
23 3 3 3 10 9 13 0 2 16 9 13 10 9 2 0 13 9 9 2 16 13 9 2
18 15 3 1 10 9 9 0 13 0 3 9 2 9 2 9 2 9 2
8 13 10 9 2 16 13 9 2
11 10 3 3 1 10 9 0 9 9 13 2
12 13 3 0 15 0 13 2 16 9 10 9 2
18 15 3 10 1 9 0 9 13 13 15 1 10 9 2 3 13 13 2
23 3 16 13 1 3 10 9 7 10 0 10 9 2 3 10 9 13 7 13 0 9 13 2
17 10 9 0 13 3 9 10 9 1 10 13 9 9 2 13 3 2
11 13 3 2 16 13 2 1 9 15 0 2
10 0 13 9 9 13 7 15 10 9 2
7 3 9 10 15 13 13 2
12 3 1 9 3 10 0 9 3 9 13 0 2
7 3 1 10 9 13 15 2
17 9 3 13 9 10 9 2 16 13 9 10 0 1 10 1 9 2
39 9 3 7 10 13 10 13 0 1 9 2 13 2 1 10 9 9 9 13 0 12 2 15 10 0 9 13 10 13 13 15 13 7 10 9 9 13 9 2
7 3 0 3 9 9 13 2
24 13 3 10 3 9 9 2 10 7 9 13 9 9 10 9 9 2 16 13 9 1 0 9 2
14 1 9 3 9 13 9 2 16 9 13 1 0 0 2
17 10 3 9 0 9 1 10 0 9 13 13 7 10 9 0 13 2
16 1 3 9 13 9 3 13 9 9 16 3 10 9 13 13 2
15 9 3 1 9 9 13 9 2 16 13 9 1 10 0 2
11 10 3 9 13 15 1 9 7 13 3 2
9 13 3 3 10 1 10 9 9 2
22 1 3 10 9 0 9 0 13 9 2 15 1 10 15 1 9 13 1 10 9 13 2
24 9 3 1 15 1 10 9 13 3 13 1 10 9 13 1 0 13 7 3 13 1 10 9 2
13 0 3 13 7 0 9 10 9 9 7 13 13 2
29 9 3 1 10 0 9 2 13 2 10 0 13 9 10 9 13 9 7 13 13 9 13 7 13 13 1 10 9 2
17 3 1 15 9 13 1 9 7 0 13 0 1 9 13 10 9 2
44 13 3 15 0 1 10 9 7 10 9 1 10 9 13 1 9 1 10 9 2 1 10 9 9 9 13 1 10 9 0 0 3 10 13 10 9 2 3 13 7 13 10 9 2
17 10 3 0 13 9 1 10 9 0 9 10 9 9 13 1 9 2
4 13 3 3 2
11 0 3 10 9 13 0 9 15 9 13 2
12 15 13 10 10 13 9 9 9 15 0 13 2
14 13 3 10 9 0 0 9 13 10 9 1 10 9 2
18 3 3 1 15 13 10 9 13 2 10 7 16 3 13 10 9 13 2
19 16 3 10 9 13 15 9 2 1 0 10 9 10 9 13 15 1 9 2
12 16 3 3 15 13 2 9 3 13 10 9 2
21 3 1 15 1 0 10 9 10 9 13 1 10 13 9 13 10 9 10 9 13 2
13 16 3 13 2 10 9 10 9 13 7 13 15 2
10 10 3 15 13 3 10 9 9 3 2
20 3 3 10 3 3 3 7 3 15 13 13 13 2 10 7 3 7 3 13 2
30 3 16 0 13 1 9 1 9 13 2 3 3 15 13 15 13 10 13 9 2 16 3 10 0 7 0 9 13 3 2
15 10 3 13 0 13 3 1 15 13 1 10 9 10 15 2
11 3 16 13 10 9 2 10 0 9 13 2
13 15 3 3 13 1 10 1 9 9 1 9 13 2
21 15 3 13 3 3 7 3 2 16 13 2 3 3 15 15 13 2 7 3 15 2
47 16 3 10 9 13 7 13 0 3 9 7 10 0 0 9 2 16 15 9 13 2 1 10 9 0 13 2 3 3 13 15 10 9 2 7 1 10 9 13 7 13 3 0 0 9 13 2
21 3 0 10 9 13 16 13 15 15 13 2 7 0 15 0 3 0 10 0 13 2
36 3 0 13 10 9 2 16 9 13 1 10 9 13 2 1 10 13 3 0 13 3 10 13 2 0 15 0 13 2 13 7 3 13 15 13 2
19 3 9 1 9 13 10 0 0 9 3 1 9 3 3 13 13 10 9 2
11 3 15 13 10 9 10 1 10 9 13 2
12 13 3 9 10 9 1 10 1 9 13 3 2
22 13 3 3 9 10 0 2 9 7 9 2 10 13 0 2 16 10 9 10 9 13 2
33 13 3 3 10 9 1 10 0 2 16 0 13 9 1 10 1 9 9 15 13 15 1 10 9 13 7 10 9 10 9 0 13 2
8 13 3 10 0 13 3 15 2
36 9 13 0 10 9 0 12 12 2 9 9 12 7 12 2 9 0 12 9 2 9 12 12 2 0 12 2 0 12 2 9 12 2 9 12 2
18 10 3 10 0 9 9 1 9 0 13 15 13 13 1 10 0 9 2
21 13 3 10 3 0 1 9 13 9 13 9 2 10 7 3 9 9 10 0 13 2
8 0 3 9 9 13 9 13 2
9 9 3 9 0 0 9 13 9 2
11 15 3 13 0 9 2 15 13 0 9 2
16 10 3 13 9 1 9 13 9 2 13 9 13 3 9 9 2
33 13 3 13 9 1 2 9 3 0 13 9 9 7 2 15 0 1 9 9 9 9 13 2 9 7 0 13 9 9 0 13 9 2
14 0 3 13 10 9 0 1 10 9 3 1 9 13 2
11 3 9 3 9 13 13 0 9 7 0 2
9 9 3 13 0 9 0 13 9 2
10 1 3 10 9 9 9 13 10 9 2
17 3 10 3 15 1 0 9 9 0 13 2 9 13 13 9 9 2
8 1 3 9 1 9 13 3 2
15 9 3 1 10 0 9 13 10 9 9 0 9 13 9 2
13 15 3 13 9 10 10 9 9 9 10 9 9 2
25 13 3 15 9 7 10 9 15 9 2 16 3 10 9 0 13 9 10 9 13 13 13 1 9 2
11 3 16 13 0 10 9 2 13 10 9 2
27 3 10 13 3 9 1 10 9 2 3 9 9 9 13 2 0 13 13 2 15 3 10 9 13 10 9 2
4 9 3 13 2
29 13 3 3 9 10 9 10 13 15 9 9 10 9 9 2 7 9 10 13 9 13 9 0 13 10 1 15 13 2
24 13 3 2 16 13 2 10 9 9 10 9 13 7 10 1 9 9 13 0 2 1 15 13 2
12 9 3 1 0 9 10 1 9 9 9 13 2
11 0 3 3 13 9 2 16 3 9 13 2
21 3 9 3 1 10 10 9 9 0 13 13 9 10 3 9 1 9 10 0 9 2
10 13 3 3 1 9 9 9 3 13 2
21 1 15 13 9 1 10 0 13 13 15 9 2 9 13 1 10 9 1 10 9 2
16 13 3 3 3 3 10 9 0 2 7 10 13 9 0 13 2
22 9 3 9 9 13 13 1 9 2 7 10 9 13 1 9 13 7 10 13 9 9 2
23 15 13 13 9 10 0 10 9 2 10 7 13 13 1 10 9 7 13 1 10 9 13 2
12 10 9 3 15 13 9 13 9 1 0 0 2
20 3 3 13 10 0 9 3 9 9 1 9 13 7 9 2 16 1 10 9 2
15 10 9 3 3 0 2 16 7 3 2 9 13 1 9 2
16 15 10 9 3 13 7 0 15 1 10 9 13 10 9 13 2
12 9 2 15 3 0 15 2 9 13 10 0 2
7 3 3 9 10 0 13 2
6 9 9 13 3 13 2
6 3 10 9 3 13 2
22 3 16 3 15 15 13 15 13 10 1 10 0 9 13 2 9 7 0 3 13 9 2
19 3 3 15 1 10 9 2 13 3 2 7 1 10 9 10 0 9 9 2
6 15 3 0 15 13 2
30 3 3 3 10 9 9 13 3 3 3 13 10 9 3 15 10 1 10 9 15 13 7 1 10 9 7 16 3 13 2
7 15 3 3 13 10 9 2
7 13 3 15 0 10 9 2
12 13 3 1 10 0 7 0 2 10 9 13 2
12 3 3 15 3 0 15 10 9 13 0 13 2
24 15 3 0 9 10 9 13 10 0 9 13 2 16 10 9 13 1 0 9 2 7 3 9 2
6 9 3 1 9 13 2
7 15 13 9 2 15 9 2
30 0 0 13 10 9 9 7 10 9 2 16 10 10 10 9 2 16 13 2 9 13 10 0 1 9 13 1 10 9 2
30 3 9 3 0 9 13 0 9 10 9 2 1 15 9 13 9 10 9 0 2 9 1 10 9 9 13 10 9 9 2
16 3 9 3 10 0 0 13 10 9 10 9 3 13 10 0 2
6 3 3 13 3 13 2
14 13 3 15 3 10 0 9 10 9 1 13 13 3 2
4 6 2 13 2
19 3 10 3 9 1 10 9 13 13 0 2 1 10 7 9 13 0 13 2
19 1 15 9 3 13 10 1 10 1 10 9 13 13 1 10 0 0 13 2
12 13 3 1 15 3 9 10 0 7 9 13 2
6 3 3 13 9 13 2
24 9 3 10 13 10 1 9 9 1 9 10 0 13 13 2 16 13 9 10 9 1 10 0 2
18 13 3 13 1 10 9 9 3 0 9 13 2 0 7 10 13 13 2
28 9 3 3 10 1 9 7 1 10 0 7 0 0 7 10 13 0 13 7 0 10 10 3 13 9 0 0 2
10 15 0 13 15 10 10 0 9 13 2
18 3 3 13 7 13 15 10 13 2 9 7 0 13 3 7 3 13 2
16 1 15 0 0 3 9 2 0 7 13 1 10 10 9 0 2
8 15 3 13 10 13 9 0 2
21 15 3 13 9 10 0 15 13 10 9 0 13 9 10 9 1 10 10 9 9 2
6 13 3 3 10 9 2
8 13 3 2 13 2 9 0 2
13 9 3 13 2 13 7 15 0 9 10 9 9 2
27 3 3 9 1 9 7 9 13 3 13 15 13 9 13 13 3 1 9 2 13 9 10 9 13 1 9 2
4 3 3 13 2
8 3 3 15 10 9 15 13 2
38 3 10 3 9 10 3 13 2 1 15 9 13 3 13 2 13 15 13 10 9 2 10 7 9 3 1 15 0 13 16 13 10 15 9 0 3 13 2
22 0 3 9 13 2 10 3 0 9 3 13 2 7 1 0 10 9 16 1 9 13 2
23 15 3 1 10 9 3 10 9 13 10 13 13 16 13 10 13 1 9 15 13 15 13 2
20 3 3 10 1 10 9 13 16 0 0 13 13 1 10 9 13 16 15 13 2
16 0 3 3 15 3 13 15 13 13 16 15 10 9 15 13 2
17 3 3 3 10 9 13 9 10 9 2 10 9 13 12 9 13 2
23 15 13 13 3 13 16 10 3 9 15 7 10 9 0 13 2 15 7 1 9 9 13 2
26 3 3 10 9 13 10 9 15 13 2 15 0 10 9 13 2 0 0 13 2 16 10 9 10 9 2
6 3 15 13 15 9 2
8 10 3 3 9 10 9 15 2
26 15 3 1 10 9 10 0 9 15 3 13 2 7 13 2 13 10 1 15 7 10 0 9 3 9 2
38 15 3 10 0 2 7 16 1 9 13 2 13 13 0 3 7 0 2 15 9 3 1 9 9 13 3 1 9 0 9 0 13 2 16 15 0 9 2
9 1 3 0 9 9 13 0 0 2
15 15 15 9 13 0 3 13 13 2 16 15 9 13 3 2
18 9 3 1 0 3 2 0 3 15 2 10 0 13 9 9 3 9 2
9 15 1 9 15 13 9 13 15 2
9 7 9 3 3 9 3 3 13 2
4 3 3 13 2
12 7 15 13 13 0 10 9 2 15 3 13 2
13 15 3 13 13 9 7 15 10 9 9 13 3 2
11 9 3 13 9 0 3 2 16 3 3 2
15 9 3 9 0 13 3 15 1 9 9 13 2 0 13 2
9 9 3 13 7 9 13 13 9 2
20 13 3 9 2 15 0 3 2 9 16 9 0 13 2 13 0 13 13 3 2
14 0 9 1 9 3 1 9 3 10 9 13 13 15 2
14 3 3 3 9 15 0 13 2 3 3 3 13 13 2
26 1 15 3 13 0 9 9 2 15 3 1 9 15 0 0 1 9 13 2 0 3 3 13 0 13 2
8 3 3 13 15 9 13 15 2
15 9 3 3 0 2 7 3 12 9 1 0 12 0 13 2
5 13 15 0 9 2
15 0 15 9 13 13 2 15 15 3 9 13 9 1 13 2
17 3 3 2 16 0 10 0 13 9 0 2 15 13 13 10 0 2
25 3 3 15 0 9 13 9 2 16 16 15 15 1 9 13 13 2 13 13 9 10 3 0 9 2
11 15 3 9 9 3 2 13 3 0 9 2
9 7 13 2 9 16 15 13 9 2
14 10 3 13 9 3 9 9 0 9 13 15 9 13 2
12 0 3 2 16 7 0 13 2 13 15 3 2
9 7 13 15 3 2 3 15 13 2
8 3 3 3 13 7 13 13 2
5 10 9 3 13 2
12 16 3 0 15 9 13 15 2 3 3 13 2
15 3 3 10 0 9 3 13 9 15 13 3 3 13 3 2
16 3 3 3 13 2 0 13 10 7 3 0 13 15 9 1 2
14 7 3 0 10 3 3 13 2 16 13 2 9 13 2
36 13 3 9 13 10 0 9 3 2 0 15 0 9 2 3 13 0 9 9 2 7 0 9 9 13 9 0 9 0 13 2 0 0 13 9 2
34 0 3 16 0 7 9 7 9 15 9 3 0 9 13 13 3 13 2 3 3 10 0 13 2 10 3 13 2 9 0 3 9 0 2
10 7 15 9 3 0 9 15 9 13 2
10 15 13 15 0 3 2 0 3 13 2
10 13 3 3 13 9 10 0 13 15 2
12 0 3 3 3 10 0 13 9 13 0 9 2
13 7 1 9 7 9 0 13 2 0 9 9 9 2
26 13 3 3 3 0 9 9 3 3 9 3 3 9 2 7 3 13 2 15 3 13 13 3 7 13 2
11 15 7 15 10 9 9 13 15 3 13 2
10 13 3 2 3 13 2 13 9 0 2
13 7 3 15 13 2 3 13 13 3 3 0 13 2
50 10 3 13 1 15 13 9 0 2 7 15 3 9 9 3 3 9 3 3 9 0 13 2 7 9 0 13 9 1 0 16 15 1 9 9 13 13 3 1 9 9 9 2 3 1 9 7 9 13 2
15 3 3 15 13 2 10 0 13 9 2 0 15 15 13 2
8 9 3 3 3 0 15 13 2
10 9 3 2 0 3 3 2 3 13 2
41 9 3 3 10 0 9 13 1 9 9 2 3 1 9 13 0 9 13 9 2 15 3 3 13 3 2 0 9 13 2 3 13 2 7 7 15 13 13 3 13 2
56 3 3 7 3 3 13 13 3 9 10 15 13 15 13 9 13 3 15 9 9 0 9 0 13 2 9 13 16 0 3 9 13 0 13 2 3 7 13 13 15 15 10 9 7 0 13 10 9 9 10 0 3 13 0 9 2
22 0 13 1 9 13 10 0 13 9 2 3 10 0 9 13 3 9 0 1 9 13 2
13 7 15 9 13 9 10 3 13 2 16 13 9 2
4 9 3 13 2
17 10 3 9 9 7 13 13 7 13 1 9 13 9 9 10 0 2
9 7 15 15 9 7 9 13 13 2
11 1 0 9 1 0 13 9 10 9 0 2
18 15 15 13 13 2 16 3 0 13 15 1 15 15 13 7 13 9 2
8 0 3 3 13 2 16 13 2
15 9 3 0 9 0 9 13 13 2 3 3 13 13 3 2
15 15 3 13 0 13 13 3 3 13 2 16 1 9 13 2
9 3 0 3 0 2 0 3 13 2
6 13 3 0 3 0 2
18 13 9 0 9 10 0 2 3 3 0 0 13 9 10 9 9 9 2
16 13 3 10 9 13 2 9 0 13 2 0 16 15 7 13 2
14 15 3 15 13 13 3 7 13 7 13 3 9 0 2
2 13 2
14 9 15 13 0 2 3 13 9 9 3 0 0 9 2
12 0 0 9 13 9 13 0 9 7 9 0 2
13 3 1 0 10 9 10 0 9 13 13 9 0 2
21 3 2 7 10 3 0 3 0 9 13 2 3 13 0 2 3 0 2 7 13 2
13 0 3 13 9 10 0 9 13 2 3 0 13 2
25 3 13 0 9 13 3 9 0 13 13 2 3 3 10 9 15 10 9 1 9 3 9 13 3 2
17 3 13 9 2 7 16 0 13 2 9 13 0 13 9 10 0 2
10 15 3 0 0 9 13 15 13 9 2
44 15 0 13 1 9 0 2 9 0 13 2 0 3 9 13 2 0 3 0 9 2 13 9 3 16 0 13 9 10 0 9 13 1 9 9 2 13 3 0 9 16 0 13 2
10 9 3 3 13 13 2 13 3 0 2
32 15 13 9 2 16 13 3 9 0 1 9 2 9 9 13 2 3 3 0 9 2 0 3 9 13 2 1 0 13 0 9 2
26 9 3 3 15 13 9 10 10 0 9 9 0 0 15 13 3 3 13 2 16 0 0 9 9 13 2
12 16 3 3 13 2 9 3 13 1 9 13 2
8 9 3 3 13 3 3 9 2
13 15 3 15 13 1 0 0 13 9 13 1 15 2
14 0 3 9 3 0 13 2 15 3 0 13 0 13 2
19 0 3 0 2 16 3 0 9 13 0 9 10 9 2 13 15 7 13 2
16 3 3 3 15 13 3 2 9 0 13 9 15 2 0 9 2
15 7 3 13 10 3 13 13 10 3 13 2 16 13 3 2
6 3 15 13 15 13 2
2 13 2
12 15 3 13 15 2 15 3 3 15 7 13 2
5 9 9 15 13 2
3 3 13 2
7 7 3 3 3 13 3 2
9 3 3 9 1 15 10 9 13 2
5 9 0 9 13 2
36 3 3 10 3 3 0 1 0 9 13 9 2 15 0 13 3 3 0 3 3 0 2 7 3 13 9 9 13 0 2 1 15 9 0 13 2
13 10 3 3 9 0 3 0 3 2 7 9 13 2
20 1 3 9 13 3 0 2 16 15 3 3 13 13 2 15 3 3 0 13 2
7 0 13 3 0 9 15 2
4 15 3 13 2
6 15 15 15 13 9 2
3 13 13 2
15 3 3 3 3 10 3 9 3 13 2 3 3 3 13 2
10 15 15 3 0 13 2 0 3 13 2
8 7 3 13 2 10 9 13 2
22 9 15 0 15 13 3 13 9 1 0 2 7 7 3 0 7 3 3 0 9 13 2
3 15 13 2
7 3 15 13 0 0 13 2
8 15 3 3 13 9 15 13 2
49 0 13 9 13 15 2 0 13 9 2 16 10 9 0 1 0 9 3 13 10 3 0 9 2 9 3 15 0 9 13 13 15 2 3 1 0 3 3 1 9 9 9 3 3 10 0 9 9 2
7 15 3 13 0 3 13 2
43 7 3 3 13 10 0 10 9 13 2 0 16 13 9 2 9 0 9 3 13 13 9 10 0 2 1 15 10 9 15 13 13 9 2 13 3 9 9 15 7 9 13 2
5 3 3 13 15 2
14 7 0 0 1 0 0 9 13 3 15 2 16 13 2
15 16 3 7 13 0 2 3 13 2 10 3 0 13 3 2
6 15 13 9 0 0 2
8 3 0 13 2 3 13 13 2
18 13 2 7 15 0 10 0 2 10 3 0 15 13 7 13 0 0 2
17 13 13 9 2 16 3 3 0 13 2 16 15 1 9 13 13 2
3 7 13 2
7 7 3 3 1 9 13 2
4 15 3 13 2
5 7 15 13 13 2
16 13 2 16 15 9 3 0 1 9 2 7 0 1 9 13 2
10 13 2 7 13 2 3 13 2 15 2
14 6 1 0 1 9 0 13 13 2 16 15 13 9 2
9 7 16 15 13 13 2 13 15 2
8 3 7 10 0 10 9 13 2
10 13 0 9 2 15 3 3 13 13 2
9 15 10 9 3 13 15 13 13 2
7 15 3 13 3 13 13 2
5 1 15 13 13 2
10 15 3 1 15 3 15 0 13 13 2
10 13 13 2 16 13 2 15 15 13 2
6 13 9 13 15 0 2
13 0 13 13 9 2 16 13 1 15 7 0 13 2
5 15 3 13 13 2
7 15 3 3 15 13 13 2
2 13 2
7 0 3 13 3 13 15 2
6 13 2 16 15 13 2
6 7 3 3 0 13 2
11 10 0 2 15 13 1 9 2 13 3 2
2 13 2
5 1 15 3 13 2
10 15 3 13 15 13 0 15 13 1 2
11 1 0 0 9 0 15 0 3 13 9 2
4 13 3 13 2
9 0 3 3 13 9 13 13 9 2
9 3 0 13 9 13 9 0 13 2
15 7 2 1 15 10 1 0 0 9 9 13 2 13 9 2
14 9 3 3 15 13 9 16 1 9 2 3 3 13 2
11 0 3 13 7 9 16 13 2 15 3 2
4 3 13 0 2
13 7 16 3 1 0 13 13 2 9 3 0 13 2
15 16 3 0 0 3 13 2 16 13 13 0 2 13 0 2
5 7 13 0 0 2
18 16 3 13 2 3 3 13 2 16 10 7 13 2 0 15 13 3 2
13 3 15 0 1 3 15 9 0 13 3 3 9 2
7 7 0 3 13 1 9 2
15 15 3 15 13 0 1 0 13 2 1 3 15 13 3 2
14 13 13 0 2 3 13 9 9 15 1 15 13 9 2
7 13 3 3 3 0 13 2
18 0 10 0 9 3 9 13 2 7 15 1 10 0 13 0 9 9 2
32 16 3 3 3 0 13 9 2 0 3 7 0 1 0 0 9 7 13 10 9 7 13 9 2 15 13 1 15 2 3 13 2
17 7 3 7 13 16 0 13 2 3 9 3 0 13 2 9 13 2
23 7 1 9 13 2 16 9 3 9 13 2 15 3 1 9 9 13 13 2 7 0 13 2
10 0 15 9 10 9 2 13 9 3 2
19 7 1 15 3 9 15 0 13 1 9 2 15 0 0 3 13 9 9 2
9 15 3 0 13 1 0 13 9 2
9 0 3 0 1 0 9 13 13 2
14 3 13 9 2 13 3 9 9 2 0 3 3 9 2
15 13 3 0 9 2 13 3 9 0 9 2 7 9 0 2
14 10 3 9 0 0 1 9 13 2 10 0 13 9 2
7 15 3 9 3 0 13 2
8 10 3 0 9 9 0 13 2
9 1 9 3 13 2 16 9 0 2
10 7 3 12 13 13 0 1 9 9 2
15 15 9 2 10 0 15 0 13 2 0 13 10 0 9 2
13 15 3 13 3 3 13 13 0 0 15 10 9 2
16 10 3 3 13 15 3 15 3 9 13 2 13 10 0 9 2
12 13 3 9 10 3 13 3 2 10 3 13 2
11 15 13 13 9 9 2 15 3 13 9 2
15 0 3 13 16 9 3 9 0 13 2 10 0 3 9 2
27 15 15 2 10 0 3 9 1 9 10 0 9 13 2 13 1 9 2 3 13 0 9 2 13 0 9 2
6 1 3 9 9 13 2
7 13 3 10 9 0 13 2
14 0 3 9 3 13 15 3 13 2 15 3 13 13 2
24 9 3 16 3 15 13 10 9 7 9 10 1 9 2 13 9 2 16 15 3 13 13 0 2
6 16 3 7 2 13 2
16 7 16 15 13 9 1 10 13 2 13 1 15 3 13 3 2
18 3 13 3 10 9 2 16 10 3 13 13 2 9 3 3 13 3 2
19 7 13 13 13 2 16 3 3 16 13 13 2 13 3 9 2 7 13 2
10 7 3 13 2 15 3 13 0 3 2
5 1 9 3 13 2
6 0 1 15 3 13 2
4 15 13 13 2
37 13 3 15 13 16 9 9 0 1 13 9 2 3 3 13 15 3 9 9 3 9 0 3 0 9 2 16 0 0 0 3 13 13 9 9 0 2
27 3 3 13 2 16 3 0 1 9 13 13 7 13 3 2 13 9 15 7 13 9 9 0 0 1 9 2
14 7 15 13 9 2 15 0 0 9 9 15 13 13 2
34 7 16 9 15 13 9 0 2 3 15 7 13 3 1 15 3 2 10 3 3 15 9 3 13 13 13 2 9 3 9 15 13 13 2
4 13 3 3 2
11 7 3 13 15 3 1 9 3 13 13 2
6 13 3 7 13 13 2
7 15 3 3 0 3 13 2
16 10 9 3 15 9 3 0 13 9 13 2 7 9 0 9 2
13 10 3 9 9 9 13 0 9 9 13 1 9 2
14 15 0 13 3 2 0 13 9 2 0 2 9 0 2
12 10 3 15 0 9 0 0 9 0 3 13 2
8 3 3 9 13 13 0 9 2
3 13 13 2
21 7 13 0 9 9 0 2 16 15 1 9 13 2 9 9 13 2 3 13 9 2
12 3 13 0 2 10 9 0 13 1 9 9 2
3 3 13 2
13 13 3 2 16 13 3 0 0 13 1 9 0 2
27 15 3 15 10 9 15 9 2 13 9 0 9 2 13 13 9 0 2 7 13 0 16 0 1 9 9 2
9 7 15 15 13 0 7 0 13 2
3 13 0 2
32 3 3 2 3 13 0 2 13 3 1 9 1 9 3 9 2 13 0 9 9 2 13 13 0 9 0 9 9 2 3 13 2
11 3 3 13 13 9 0 2 0 9 13 2
20 10 3 9 13 13 3 10 9 2 15 13 2 1 0 9 2 9 1 9 2
4 15 13 0 2
23 1 3 9 2 3 13 2 13 0 9 2 0 9 16 0 0 13 1 9 0 1 9 2
7 13 3 15 9 0 13 2
18 3 3 3 3 2 1 15 13 10 9 15 13 9 2 15 13 1 2
11 3 13 2 7 10 13 13 13 13 15 2
12 15 15 0 2 16 3 13 2 10 9 13 2
14 0 3 0 2 16 15 7 13 9 2 15 0 13 2
19 10 3 13 9 13 7 9 9 13 2 15 3 13 2 13 15 0 9 2
15 1 3 15 15 9 13 9 9 0 3 3 13 7 15 2
14 3 13 2 0 16 13 2 0 1 9 15 13 3 2
17 13 3 9 0 3 13 2 10 3 9 3 13 10 9 13 1 2
17 3 13 1 10 7 0 9 3 3 9 2 15 7 9 15 13 2
17 0 3 3 13 3 10 10 0 9 2 7 15 9 13 3 0 2
16 13 3 13 15 10 0 9 2 16 7 15 13 9 10 15 2
10 10 3 13 15 3 13 3 0 13 2
11 15 1 9 13 0 3 9 13 15 13 2
7 3 3 13 9 7 13 2
8 3 15 10 0 13 0 9 2
17 15 0 13 2 16 15 13 2 13 3 12 0 13 9 9 9 2
9 3 10 0 3 12 13 0 9 2
15 7 0 3 0 0 9 2 9 3 13 7 9 2 13 2
28 16 3 0 9 13 9 0 1 0 9 2 9 13 9 2 7 13 9 0 2 16 9 2 9 0 1 9 2
6 13 3 9 9 0 2
8 3 0 0 9 9 3 13 2
15 15 3 0 13 0 10 0 0 9 13 2 3 13 13 2
25 0 16 13 7 0 9 0 9 13 2 13 9 15 2 9 3 13 2 13 1 0 1 9 9 2
13 9 3 0 9 13 2 0 9 13 9 3 3 2
14 0 3 13 9 9 2 15 3 13 2 15 3 13 2
6 0 13 9 0 13 2
13 3 3 13 9 2 0 3 0 9 9 3 9 2
17 7 13 3 2 7 3 3 15 13 3 3 15 7 15 13 9 2
20 16 3 9 13 2 7 15 1 3 15 9 13 7 0 2 3 3 3 13 2
16 0 13 2 1 0 9 13 15 1 9 15 13 3 13 9 2
10 7 15 3 7 13 13 7 13 3 2
6 16 9 3 2 13 2
4 15 3 13 2
8 3 13 16 13 13 10 0 2
3 13 13 2
9 9 9 0 0 13 3 13 0 2
15 9 3 3 9 15 13 13 0 2 15 9 7 13 13 2
4 7 13 13 2
12 10 3 9 15 0 13 9 2 15 0 13 2
6 7 15 3 0 13 2
15 3 3 3 10 3 13 3 1 3 0 9 13 13 9 2
38 16 3 15 9 0 9 13 0 9 9 2 13 9 2 15 13 9 2 13 3 0 9 2 3 15 3 9 0 16 3 13 2 0 3 9 13 9 2
11 9 3 3 15 13 9 0 0 9 13 2
38 15 15 10 9 0 0 13 9 9 0 13 9 10 3 0 13 2 10 3 1 0 9 13 0 9 3 3 0 13 2 3 3 0 0 13 9 9 2
10 10 3 13 9 13 0 7 0 9 2
4 13 9 9 2
10 10 3 0 9 0 0 15 13 9 2
13 0 15 0 2 7 13 15 9 1 9 3 13 2
3 15 13 2
15 13 15 3 0 2 7 0 9 3 2 7 15 13 9 2
10 13 9 10 0 9 0 1 0 9 2
3 0 13 2
4 13 10 0 2
3 0 13 2
6 15 9 13 15 13 2
3 0 13 2
11 15 9 7 15 9 15 9 9 0 13 2
8 3 13 1 9 9 13 0 2
7 13 2 3 3 0 9 2
3 15 13 2
3 13 13 2
6 0 1 0 13 15 2
3 15 13 2
12 13 13 3 0 10 0 15 9 9 15 9 2
14 3 3 2 16 13 0 13 0 13 2 3 3 13 2
8 7 0 13 15 9 0 13 2
7 13 3 2 16 13 15 2
31 3 3 3 9 13 2 16 15 0 13 9 9 2 13 10 0 13 2 0 10 0 9 13 7 10 9 1 10 0 9 2
13 16 3 15 13 2 3 15 13 10 0 9 13 2
6 15 0 9 13 13 2
11 13 3 10 9 9 10 0 0 13 9 2
24 0 13 0 9 13 10 0 9 2 3 0 13 9 9 2 1 3 13 9 0 9 3 0 2
14 15 0 13 2 0 13 2 10 9 13 10 13 15 2
19 1 15 10 3 3 3 13 2 13 0 0 9 9 1 9 7 9 13 2
6 13 3 10 9 13 2
23 13 3 0 9 1 9 16 13 15 2 3 13 15 1 9 16 0 1 10 9 13 15 2
4 0 3 13 2
15 3 3 13 10 3 3 2 16 3 13 15 10 13 9 2
12 15 3 13 13 9 2 15 3 13 1 9 2
26 6 0 15 13 0 9 9 2 15 15 13 1 9 2 16 10 0 0 9 7 0 13 0 13 3 2
11 3 3 3 3 3 13 2 0 3 9 2
6 15 3 3 13 15 2
8 3 0 13 0 0 13 9 2
3 15 13 2
4 15 3 13 2
4 13 3 0 2
6 7 13 13 9 0 2
3 3 13 2
3 13 9 2
8 1 15 9 13 13 0 9 2
6 15 3 3 0 13 2
18 3 13 15 0 13 9 9 13 7 3 13 15 1 9 9 3 9 2
10 3 3 13 3 3 13 0 15 13 2
8 0 15 3 13 9 2 0 2
16 15 7 3 15 13 10 0 13 9 2 15 0 9 9 13 2
5 9 3 3 13 2
5 15 15 15 13 2
3 3 13 2
5 13 15 2 13 2
6 13 15 15 7 13 2
18 13 3 15 2 0 3 9 3 3 3 3 3 3 13 15 13 9 2
4 0 13 9 2
7 15 15 15 15 13 13 2
12 13 3 3 2 13 0 13 15 0 0 9 2
23 13 3 9 2 15 15 13 0 9 0 2 15 3 13 13 3 2 3 3 3 15 13 2
31 3 0 3 3 9 10 9 13 3 10 0 9 15 2 0 15 10 9 9 9 13 9 10 0 9 0 9 2 15 13 2
34 9 3 13 1 3 0 13 9 2 9 3 9 13 13 2 1 3 0 9 15 13 3 2 7 13 9 10 0 2 0 15 13 9 2
30 3 0 9 9 2 3 10 0 9 9 3 3 0 9 2 3 9 3 3 0 3 0 15 9 13 13 2 13 3 2
16 9 3 2 0 13 3 9 9 2 0 15 3 13 9 3 2
32 13 3 15 0 0 2 15 16 9 13 13 2 7 15 3 3 3 9 3 15 9 13 3 13 13 2 7 0 3 13 0 2
15 7 3 13 13 3 9 2 13 3 0 0 9 1 13 2
6 13 3 15 1 9 2
9 13 3 3 3 2 13 2 13 2
13 0 3 9 0 13 2 0 0 13 15 0 9 2
23 7 3 3 3 15 13 2 16 10 9 13 7 9 13 2 10 3 13 15 13 1 15 2
16 13 0 2 16 13 0 13 16 7 13 0 3 7 13 13 2
7 13 3 15 15 0 13 2
11 13 15 15 2 7 0 3 13 9 0 2
13 3 3 3 13 1 15 13 13 1 15 13 3 2
5 13 15 13 13 2
8 13 3 3 16 7 13 13 2
11 7 3 3 3 3 15 3 1 9 13 2
9 13 2 13 3 16 13 0 13 2
2 13 2
4 13 3 0 2
6 9 3 1 0 13 2
10 3 15 13 9 2 16 10 0 13 2
4 0 9 13 2
5 13 3 3 13 2
7 0 10 9 13 0 13 2
13 9 3 13 13 15 13 2 16 13 10 3 9 2
12 9 3 9 13 15 15 9 10 0 13 9 2
8 13 13 2 9 3 13 15 2
14 7 3 3 9 3 2 7 0 9 13 16 13 9 2
17 9 3 15 3 13 0 13 2 15 3 3 10 9 9 13 13 2
10 13 3 3 13 0 13 9 0 13 2
21 15 3 13 0 1 9 3 2 10 13 15 13 1 2 7 15 9 13 9 13 2
18 15 3 10 9 9 2 3 10 0 13 0 2 3 13 15 13 13 2
46 13 3 15 0 13 0 9 0 2 10 3 0 2 15 15 0 7 9 15 9 13 9 13 1 10 0 7 0 9 2 15 15 9 10 13 7 13 3 13 9 10 13 15 9 13 2
4 13 13 3 2
10 15 3 13 3 0 0 1 13 15 2
7 10 3 13 9 3 13 2
6 13 9 0 0 15 2
8 3 1 15 9 15 3 13 2
8 3 0 13 3 3 13 15 2
8 13 9 3 10 15 13 9 2
4 7 15 13 2
7 13 15 2 9 13 0 2
9 16 3 3 13 2 9 13 13 2
4 3 7 13 2
3 13 3 2
4 13 3 3 2
8 13 3 10 9 9 0 9 2
41 3 3 13 0 13 15 9 9 7 1 15 13 0 2 0 3 9 10 0 9 13 2 0 3 9 13 3 0 9 2 9 0 13 2 7 0 13 9 9 13 2
14 16 3 7 2 13 15 15 7 1 13 0 3 0 2
4 0 15 13 2
14 16 3 7 2 9 0 13 15 3 3 0 13 3 2
9 7 3 13 9 3 13 15 0 2
10 7 16 13 1 0 2 0 3 13 2
7 9 3 3 9 3 13 2
9 10 3 0 13 3 13 0 9 2
5 7 13 7 0 2
10 13 3 15 9 0 1 0 0 13 2
6 10 0 13 3 9 2
8 9 13 2 16 3 13 15 2
2 13 2
20 0 15 13 2 16 13 13 2 0 9 13 2 13 9 2 3 3 13 9 2
2 13 2
13 10 3 3 0 13 15 0 13 10 3 13 9 2
16 10 3 13 13 0 2 10 3 3 13 13 15 3 3 13 2
7 7 13 0 15 13 13 2
12 9 15 2 3 13 2 3 13 15 13 9 2
11 7 3 9 9 13 15 13 10 0 9 2
8 15 3 15 1 13 13 0 2
7 3 3 13 10 13 13 2
7 13 13 3 15 3 15 2
5 0 9 13 9 2
11 3 13 3 13 2 10 0 9 13 9 2
14 7 3 15 0 3 13 0 9 9 13 10 9 3 2
4 13 15 13 2
11 7 15 13 1 10 0 13 10 0 0 2
23 16 3 0 13 0 9 1 9 10 3 2 0 13 0 2 3 3 13 3 3 3 13 2
4 15 3 13 2
6 13 3 15 13 9 2
16 3 3 9 15 10 9 9 15 3 13 2 15 3 13 13 2
20 9 3 2 16 13 2 1 9 9 0 7 9 1 9 13 10 3 0 0 2
32 10 3 3 13 9 9 9 13 13 10 7 9 13 3 3 13 15 2 13 3 0 2 0 2 9 0 9 13 1 9 9 2
15 3 13 15 0 2 7 13 3 7 0 13 7 0 0 2
6 16 13 7 13 13 2
5 3 9 3 13 2
9 3 3 13 13 15 2 0 9 2
6 3 3 3 13 13 2
9 7 0 0 10 0 15 13 1 2
16 0 3 9 12 0 1 9 13 10 0 9 0 13 0 9 2
21 3 3 3 0 3 15 13 13 0 0 13 2 16 9 9 9 9 7 9 13 2
15 7 13 13 15 3 9 16 13 2 3 1 9 3 13 2
20 15 3 3 13 15 1 9 9 13 2 16 13 15 2 10 1 9 13 13 2
9 10 3 0 13 3 13 9 0 2
20 3 3 3 13 3 3 3 2 16 13 3 13 2 15 3 3 3 13 1 2
11 7 13 0 15 13 2 0 3 15 13 2
5 3 3 3 13 2
13 15 3 2 16 13 2 10 10 9 0 13 13 2
14 15 3 3 0 13 2 10 3 9 9 13 13 0 2
6 15 3 15 3 13 2
9 15 3 3 9 13 9 0 13 2
5 10 0 13 9 2
17 7 3 13 3 0 15 9 2 3 3 13 2 1 3 3 15 2
11 0 0 13 13 2 16 7 0 13 15 2
6 0 1 0 9 13 2
9 7 13 13 15 3 13 15 13 2
4 7 0 13 2
9 3 2 16 3 7 13 2 13 2
7 9 3 13 3 13 0 2
16 16 0 13 2 13 3 1 15 2 0 3 10 13 13 9 2
13 7 13 15 7 10 1 15 9 13 10 0 0 2
11 13 3 3 0 0 16 7 3 3 13 2
7 7 16 13 15 2 13 2
30 15 1 0 9 9 13 9 1 0 0 13 9 1 9 3 13 2 0 9 9 0 2 0 1 9 1 3 0 9 2
26 13 3 1 9 13 13 9 9 0 9 13 2 16 3 0 9 9 13 3 7 9 9 0 9 13 2
11 0 1 9 13 9 9 2 0 9 9 2
28 9 3 0 9 9 13 2 7 15 13 0 9 13 9 9 9 2 0 13 9 9 1 0 3 9 13 13 2
19 0 3 1 9 13 13 0 2 15 3 13 1 9 13 13 9 0 9 2
16 13 3 0 15 3 2 0 3 1 0 13 13 0 9 9 2
38 12 9 3 1 12 9 13 0 1 0 13 9 0 0 9 2 1 10 0 2 15 9 9 9 3 0 13 1 0 0 9 13 13 0 9 9 0 2
35 7 3 10 0 13 9 10 0 13 9 2 1 3 3 9 10 3 13 9 2 9 3 9 9 0 0 13 2 10 9 3 0 0 13 2
40 15 3 15 9 1 0 3 13 13 0 3 10 9 13 13 3 9 3 9 2 0 3 2 3 9 13 9 2 16 13 2 1 10 0 3 9 13 0 9 2
31 16 3 0 1 0 9 0 1 9 13 13 3 7 13 0 1 9 2 15 9 3 0 7 9 13 9 1 9 10 13 2
26 15 3 15 0 13 9 7 10 0 13 9 7 1 9 15 9 13 13 0 13 3 3 7 3 13 2
14 7 0 15 1 10 0 9 0 13 2 0 3 13 2
20 15 15 9 15 13 9 2 7 3 0 15 13 13 9 9 10 1 9 1 2
15 15 0 9 2 3 1 3 15 9 13 10 0 10 0 2
15 7 15 0 15 10 9 2 13 7 13 3 1 15 13 2
14 9 3 13 0 3 13 15 7 15 13 0 13 1 2
6 0 15 0 13 13 2
8 7 13 0 10 0 3 9 2
8 15 3 3 0 0 13 3 2
8 3 13 3 0 15 13 13 2
9 7 1 9 9 10 9 3 13 2
12 0 3 13 9 9 2 9 13 15 1 9 2
7 9 3 13 0 15 13 2
6 3 15 3 3 13 2
6 0 13 13 9 0 2
6 3 9 0 13 0 2
8 9 3 3 3 13 13 15 2
9 16 10 9 13 2 13 3 3 2
15 10 9 3 13 13 2 10 7 13 3 0 1 15 0 2
9 15 3 13 1 15 15 13 9 2
6 13 13 15 0 15 2
23 10 3 9 3 3 13 3 3 13 15 13 10 13 2 3 3 3 3 1 0 13 15 2
8 3 3 13 13 9 15 9 2
7 13 3 7 15 13 0 2
8 10 0 3 3 13 9 0 2
8 3 13 3 2 3 13 13 2
5 7 3 13 15 2
15 10 0 15 3 13 13 1 9 0 9 13 13 15 13 2
3 15 13 2
7 15 9 13 10 13 15 2
3 3 13 2
18 0 3 9 7 9 2 9 3 3 13 9 2 7 0 9 15 13 2
13 16 3 10 0 15 9 13 2 0 9 0 13 2
15 9 3 15 13 0 13 2 0 0 2 7 13 7 13 2
27 13 3 0 7 9 13 9 7 9 13 7 9 13 2 10 3 13 3 15 13 10 9 13 3 3 13 2
21 9 3 16 0 13 13 0 2 13 15 9 2 15 0 1 9 9 13 9 13 2
12 3 3 13 3 3 13 3 16 13 3 13 2
13 13 3 10 9 16 0 15 9 13 15 3 0 2
7 13 3 0 9 0 9 2
13 13 3 3 0 9 13 9 13 15 10 0 1 2
20 0 13 3 9 13 0 2 15 0 9 13 13 9 7 9 0 7 9 13 2
7 7 10 0 13 13 9 2
3 3 13 2
27 7 0 7 3 9 9 3 13 13 15 2 3 9 13 2 3 3 1 9 9 3 13 2 3 13 15 2
10 1 15 0 13 3 13 9 13 15 2
9 0 3 9 0 9 0 9 13 2
10 0 7 9 13 2 15 9 13 9 2
12 15 13 7 13 9 0 1 0 9 13 9 2
11 9 3 13 9 13 7 0 9 9 13 2
13 0 3 13 13 15 2 9 3 13 16 13 9 2
18 7 16 13 9 3 1 15 9 2 3 0 13 2 0 3 15 13 2
13 1 10 3 0 9 10 0 13 13 3 7 13 2
8 13 15 13 7 13 3 13 2
8 3 13 7 3 16 3 13 2
12 10 13 15 13 10 9 2 10 3 9 15 2
5 13 3 10 9 2
17 16 3 0 7 13 15 10 13 2 13 16 10 0 9 9 13 2
5 7 13 3 3 2
15 7 3 3 1 9 9 3 0 13 13 10 9 0 9 2
8 0 10 0 0 9 0 13 2
14 0 7 0 3 9 0 9 13 2 0 13 1 9 2
20 0 3 9 9 13 13 7 9 0 9 9 3 0 9 9 0 2 0 9 2
19 13 3 9 0 9 9 2 9 3 9 13 1 9 13 0 3 9 9 2
19 7 9 7 0 9 7 9 9 13 7 0 9 0 7 0 13 9 0 2
7 0 1 0 13 15 13 2
6 9 0 9 3 13 2
6 9 3 0 9 13 2
11 3 15 0 13 3 0 13 15 15 13 2
6 1 0 9 13 15 2
9 3 13 13 15 3 13 9 9 2
15 3 3 3 15 3 13 10 0 13 9 7 1 9 13 2
4 15 13 13 2
8 15 1 9 0 1 13 13 2
4 15 3 13 2
5 0 0 13 9 2
15 9 3 3 13 2 7 13 0 9 2 3 0 2 15 2
9 15 3 0 0 13 15 13 0 2
8 13 3 15 15 9 3 13 2
5 0 10 9 13 2
3 0 13 2
9 3 7 13 7 13 3 15 13 2
6 3 0 7 0 13 2
6 7 3 13 0 13 2
5 0 13 10 9 2
17 9 15 13 0 2 16 1 9 0 13 0 9 9 7 9 13 2
6 13 3 13 0 9 2
21 3 3 0 2 0 16 13 9 2 9 13 2 1 3 9 0 13 10 9 13 2
22 15 13 13 2 1 3 15 13 3 0 13 2 7 15 3 3 10 3 3 13 9 2
11 0 3 15 13 2 3 3 15 3 3 2
11 7 0 0 0 13 15 13 10 0 9 2
8 7 13 13 3 13 10 7 2
12 15 3 13 3 15 3 13 1 0 9 0 2
2 13 2
5 15 3 3 13 2
4 0 3 13 2
7 7 3 13 15 13 9 2
24 3 3 15 15 9 13 10 13 15 2 3 3 10 0 10 3 9 9 15 1 9 13 9 2
19 3 3 13 0 13 10 0 9 2 16 0 0 9 0 13 0 13 13 2
16 0 15 3 13 2 9 0 9 13 2 1 9 10 9 13 2
8 13 3 13 2 15 3 3 2
12 16 3 10 9 1 13 2 9 0 15 13 2
16 15 3 1 0 3 15 0 13 2 3 15 3 13 9 13 2
17 7 3 2 16 15 1 0 9 13 0 13 9 2 0 3 13 2
5 15 3 3 13 2
15 15 3 16 13 3 0 13 13 2 3 15 0 9 13 2
10 13 10 9 0 1 0 9 10 9 2
6 13 3 3 13 0 2
25 7 13 3 15 0 3 9 13 3 2 7 10 0 9 0 1 9 0 13 7 13 0 3 13 2
9 0 9 3 13 10 13 9 13 2
11 3 3 13 13 0 15 9 13 15 3 2
12 0 3 13 3 3 13 2 9 13 10 13 2
21 7 7 9 7 0 10 0 15 9 0 13 2 0 3 10 0 3 13 9 0 2
10 7 3 3 0 0 13 15 13 9 2
4 7 15 13 2
11 1 3 13 3 13 0 3 3 0 9 2
13 13 3 3 16 1 0 15 13 3 0 13 13 2
8 13 15 0 16 13 15 13 2
5 0 13 0 13 2
4 15 3 13 2
8 3 3 7 15 0 13 13 2
14 3 3 9 3 3 0 13 16 10 0 1 9 13 2
13 0 0 0 13 13 3 2 16 7 9 13 9 2
15 7 10 9 0 3 0 13 13 0 13 13 3 15 13 2
7 15 0 0 15 0 13 2
8 13 0 2 15 3 13 9 2
10 15 3 3 13 2 15 3 16 13 2
7 3 3 0 0 13 9 2
7 3 13 0 10 13 9 2
9 3 3 15 9 2 7 9 13 2
9 3 10 3 9 10 9 0 13 2
7 15 13 16 3 0 15 2
7 3 13 2 7 13 13 2
10 3 3 13 2 16 0 2 13 0 2
7 15 3 13 3 13 9 2
12 9 3 9 1 0 9 13 2 13 9 9 2
13 13 9 2 16 15 13 7 13 7 13 10 0 2
13 7 1 0 10 0 3 13 0 15 10 9 13 2
8 9 3 15 13 3 13 0 2
4 13 13 15 2
3 9 13 2
8 15 0 13 15 2 0 13 2
10 13 3 3 16 13 3 1 15 13 2
10 15 3 3 7 3 15 3 13 15 2
3 13 15 2
5 3 13 15 13 2
10 15 3 3 13 13 2 15 3 13 2
2 13 2
18 10 9 13 15 10 3 3 0 13 2 15 3 1 15 15 0 13 2
5 3 3 13 3 2
7 7 13 0 10 15 9 2
6 0 3 0 13 9 2
6 0 15 9 9 13 2
10 3 3 13 7 15 7 10 0 9 2
8 3 3 13 15 10 15 9 2
8 9 10 13 15 10 9 13 2
11 1 3 15 13 9 13 15 3 3 13 2
15 13 3 3 10 0 2 16 3 3 10 9 13 10 9 2
15 15 3 3 13 3 9 2 9 0 13 9 1 9 13 2
24 0 16 0 9 0 16 0 9 0 13 9 2 13 3 0 9 2 7 0 9 13 9 9 2
27 0 10 9 9 13 9 0 1 9 13 2 3 3 13 9 9 2 7 13 9 15 2 3 3 13 9 2
28 3 3 0 1 9 15 13 9 1 9 9 2 1 3 15 0 9 10 0 13 9 9 3 9 7 9 9 2
24 15 3 9 13 3 10 0 13 2 3 3 9 0 9 2 0 3 9 9 13 9 0 9 2
12 13 3 0 13 2 16 9 0 9 15 13 2
8 9 3 1 15 0 9 13 2
7 13 3 0 9 1 9 2
11 3 13 9 13 9 9 2 9 9 13 2
5 3 13 9 0 2
11 15 3 0 13 9 0 13 15 3 13 2
10 15 3 13 3 9 0 16 0 0 2
14 7 13 3 3 0 13 10 9 1 9 15 13 15 2
22 16 3 0 13 3 15 9 13 1 0 0 2 0 3 15 3 13 9 2 7 13 2
6 1 0 13 9 0 2
15 1 10 3 0 15 13 9 0 2 13 1 9 0 13 2
20 15 3 13 7 9 13 7 13 10 13 13 2 3 13 9 0 1 15 13 2
14 7 15 9 13 15 13 13 7 0 7 0 7 0 2
28 7 0 3 10 9 13 15 3 3 13 2 3 3 3 13 13 2 9 3 3 1 9 13 13 0 0 9 2
7 9 3 0 3 13 0 2
15 0 9 13 2 15 0 9 13 2 15 0 9 9 13 2
10 10 3 13 13 10 0 9 10 9 2
11 3 0 13 10 13 2 3 9 3 0 2
17 0 3 2 16 13 2 1 9 13 2 3 3 9 0 13 3 2
16 15 3 2 16 7 10 9 13 2 13 3 15 13 13 1 2
17 15 3 16 15 7 13 3 15 2 3 3 3 13 3 13 13 2
6 13 3 0 3 13 2
16 15 3 3 13 0 13 0 13 15 7 13 15 7 13 13 2
19 15 10 0 0 1 9 13 0 3 1 9 9 13 13 3 1 9 15 2
6 15 0 3 13 9 2
24 15 3 0 7 13 0 13 2 7 9 2 15 3 0 2 7 9 13 2 0 13 13 0 2
18 13 1 9 0 0 9 13 2 9 3 13 2 10 3 13 0 13 2
18 3 3 9 15 0 9 13 13 9 2 0 3 13 10 0 9 13 2
7 7 13 7 9 9 13 2
20 9 3 16 15 1 15 0 13 2 13 15 13 0 13 10 9 0 9 0 2
5 3 3 13 3 2
12 10 0 7 13 3 13 1 9 0 10 9 2
14 16 3 15 0 2 3 10 9 13 3 16 9 13 2
7 9 3 13 10 13 13 2
9 3 3 3 13 13 1 10 0 2
7 3 15 3 15 13 9 2
7 3 13 9 15 9 9 2
8 9 3 15 15 13 13 13 2
8 13 15 3 13 3 3 0 2
9 9 3 3 13 15 9 13 9 2
7 3 10 13 10 9 13 2
9 3 3 0 3 15 9 13 0 2
9 15 2 3 13 2 10 9 13 2
5 15 3 3 13 2
7 3 3 0 15 13 13 2
7 13 3 10 0 9 13 2
9 3 3 13 9 3 10 9 13 2
9 3 3 13 0 3 10 0 15 2
9 0 3 3 13 16 3 13 13 2
9 15 3 3 13 7 13 13 15 2
6 7 13 3 13 0 2
9 15 3 13 9 1 0 9 13 2
8 13 13 2 13 9 0 0 2
12 16 7 9 13 2 13 3 15 3 3 13 2
7 9 13 9 7 13 15 2
8 13 13 15 7 13 9 13 2
13 13 10 9 16 1 9 3 13 13 0 10 9 2
7 9 3 13 0 13 0 2
2 13 2
7 13 0 16 1 9 13 2
9 10 3 3 9 15 3 13 9 2
7 0 3 0 7 13 13 2
5 3 3 3 13 2
8 9 3 0 7 15 13 13 2
26 13 0 3 3 13 9 9 13 0 13 1 9 2 9 0 16 9 0 13 2 16 9 0 13 9 2
29 3 10 9 2 15 0 13 9 2 13 3 13 10 7 13 2 7 13 3 7 3 16 9 0 13 1 9 13 2
5 10 3 13 13 2
15 13 3 0 9 9 0 9 2 10 0 0 1 9 9 2
28 7 15 10 9 9 13 13 10 9 9 2 3 9 0 2 3 3 0 3 15 15 9 13 2 7 9 13 2
31 3 0 7 9 13 1 15 13 9 9 2 3 3 9 13 9 3 3 9 9 13 2 7 0 13 0 3 0 9 13 2
41 13 3 0 13 10 0 0 9 9 1 0 2 15 9 3 0 0 9 13 2 7 15 9 13 2 3 9 9 2 9 3 0 13 2 13 3 1 9 0 9 2
6 15 15 9 0 13 2
14 15 15 2 1 9 0 2 3 13 13 2 7 0 2
6 0 3 13 15 9 2
16 13 0 15 9 2 9 0 9 10 3 0 0 9 0 9 2
9 1 15 0 0 15 15 9 13 2
14 13 3 9 15 2 9 3 15 9 13 0 0 13 2
6 15 3 0 13 9 2
9 10 3 0 9 0 0 0 13 2
21 3 13 2 9 7 9 1 10 13 16 3 3 3 9 13 3 2 16 13 13 2
5 3 13 3 0 2
23 7 0 9 13 2 3 13 15 2 13 0 0 2 3 13 13 7 1 0 13 13 9 2
14 15 3 0 1 15 10 9 9 3 3 10 3 13 2
27 3 3 3 3 3 3 2 16 9 9 13 2 3 3 16 9 15 13 13 2 9 9 15 3 13 9 2
8 15 9 3 0 1 9 13 2
33 9 3 3 15 13 0 13 2 7 9 1 0 9 2 16 15 13 2 9 3 1 9 7 9 13 3 13 9 15 3 13 3 2
36 7 3 13 15 1 9 3 13 0 2 0 2 3 3 15 9 9 13 3 3 0 9 2 7 3 0 1 0 10 0 13 1 13 13 9 2
10 15 13 15 10 0 1 9 3 13 2
15 7 16 3 3 15 13 1 9 0 2 13 3 13 13 2
15 16 3 15 13 2 7 0 0 13 16 7 13 3 15 2
11 3 10 0 9 0 9 9 15 3 13 2
9 3 0 10 13 9 13 9 1 2
9 13 0 13 7 3 15 3 13 2
11 13 7 9 0 9 13 9 1 0 9 2
7 13 3 1 0 9 13 2
9 3 10 9 0 13 0 3 9 2
10 0 13 9 13 10 9 1 0 9 2
14 13 3 3 0 9 0 3 9 2 0 3 13 9 2
13 1 3 13 0 0 9 13 2 9 13 0 9 2
24 15 3 9 3 0 13 9 2 0 3 1 9 13 9 1 0 0 0 9 1 9 9 9 2
9 10 0 3 0 9 1 9 13 2
7 3 3 3 0 13 9 2
7 3 1 0 15 13 9 2
5 13 13 13 0 2
8 13 13 3 3 1 9 9 2
4 15 3 13 2
7 3 15 10 0 13 9 2
8 13 2 9 9 10 0 13 2
25 1 3 0 9 0 13 2 7 13 15 0 9 9 2 9 13 9 9 2 0 13 9 7 13 2
8 7 13 1 9 0 9 13 2
7 9 3 9 3 0 13 2
8 3 3 13 0 13 9 0 2
11 0 9 15 13 1 2 13 0 9 9 2
9 7 0 10 0 1 9 13 9 2
25 3 3 13 0 9 3 9 1 15 3 3 9 9 2 3 3 9 0 13 9 0 13 9 9 2
8 9 3 10 0 0 13 13 2
23 16 3 13 2 0 3 13 9 0 3 3 0 2 15 1 0 13 13 3 3 0 13 2
5 9 3 9 13 2
9 7 13 10 13 3 3 13 13 2
6 3 15 13 3 13 2
8 15 3 1 9 13 13 3 2
10 3 3 13 16 9 13 0 9 13 2
8 3 13 9 15 2 3 13 2
5 0 0 0 13 2
8 0 15 3 10 9 0 13 2
7 3 13 10 9 13 3 2
9 7 3 13 2 0 15 13 13 2
7 15 3 1 9 9 13 2
8 3 13 9 13 15 13 13 2
2 13 2
8 1 15 3 15 13 13 9 2
7 13 15 0 1 9 13 2
9 3 3 3 7 13 10 0 9 2
56 7 3 3 3 13 7 0 3 9 9 9 13 2 1 15 10 0 0 1 9 9 9 0 9 13 13 2 1 15 13 3 15 3 13 3 9 3 3 1 9 13 2 13 3 10 3 3 3 9 0 2 0 2 0 9 2
17 0 15 9 0 13 9 7 9 9 2 1 10 0 15 13 0 2
7 7 0 13 16 13 13 2
12 13 3 3 0 9 9 9 9 0 9 9 2
25 0 3 0 13 9 2 0 9 7 9 13 7 9 7 15 0 9 2 13 0 9 0 1 9 2
22 13 3 2 1 15 0 15 15 1 9 13 9 2 7 3 3 0 9 1 9 13 2
6 13 0 7 13 9 2
15 10 3 13 3 0 2 13 3 9 13 9 1 0 1 2
5 15 3 13 13 2
2 13 2
4 13 3 15 2
14 13 9 3 1 9 9 13 2 13 3 10 13 9 2
7 7 0 13 7 13 13 2
8 13 3 9 0 10 0 9 2
9 3 3 2 9 3 13 10 13 2
10 13 3 15 13 7 3 1 0 13 2
6 3 3 13 13 3 2
15 15 3 2 16 9 3 13 2 0 3 13 7 13 13 2
13 13 3 16 10 13 9 0 13 13 10 9 13 2
19 15 3 1 0 9 9 13 9 2 3 0 13 9 9 2 9 3 9 2
19 7 15 0 9 0 9 0 3 9 0 13 2 0 9 13 0 13 9 2
10 10 1 0 13 0 9 9 1 0 2
28 9 3 13 0 2 3 15 2 3 2 13 3 0 15 0 9 13 3 9 0 9 13 2 13 0 9 9 2
5 7 3 13 0 2
18 10 3 9 16 13 9 2 3 13 15 13 0 2 7 0 13 9 2
16 13 3 3 1 9 2 16 13 2 0 7 13 0 9 13 2
19 16 3 13 0 10 13 2 0 15 9 9 3 3 13 9 1 10 9 2
9 15 3 3 15 9 9 13 13 2
2 13 2
4 7 15 13 2
2 13 2
3 9 13 2
4 9 3 13 2
7 3 3 13 0 13 1 2
10 7 3 13 0 9 3 9 10 9 2
10 1 3 9 3 13 9 7 9 1 2
7 0 3 3 0 13 13 2
11 15 3 15 13 3 15 1 9 9 13 2
18 15 3 0 9 13 9 9 1 0 2 3 13 0 0 9 9 3 2
16 15 3 0 0 13 9 13 3 3 2 13 3 9 13 0 2
8 3 0 9 13 10 13 9 2
5 9 15 13 9 2
7 15 1 0 9 9 13 2
4 15 9 13 2
5 1 15 9 13 2
18 15 3 0 9 13 10 9 2 13 9 0 13 2 9 13 0 9 2
7 1 3 13 9 9 13 2
24 3 10 0 0 13 2 3 13 2 13 13 9 0 9 2 1 3 0 9 3 0 9 13 2
10 7 13 0 13 9 0 9 0 9 2
5 15 0 3 13 2
3 0 13 2
22 9 3 13 9 9 13 1 9 9 3 13 2 7 1 9 1 9 13 9 0 13 2
3 3 13 2
15 15 3 3 10 3 3 9 0 13 13 10 3 0 9 2
15 7 13 2 7 15 7 0 3 13 9 13 2 9 13 2
14 3 3 3 13 2 7 10 3 3 13 3 9 9 2
9 15 3 13 3 0 1 0 3 2
3 13 13 2
9 15 3 2 15 15 9 3 13 2
32 15 3 0 0 1 9 13 0 9 2 13 3 10 3 13 9 0 9 2 3 3 15 2 0 3 15 0 9 13 10 0 2
9 15 15 3 0 13 15 0 9 2
12 3 9 3 15 0 13 1 10 13 15 13 9
7 0 3 13 1 9 9 2
9 9 13 2 16 15 9 1 0 2
14 13 13 2 13 9 10 0 13 15 0 13 9 0 2
9 13 13 2 16 3 9 0 13 2
7 10 13 15 13 13 13 2
6 13 3 15 15 13 13
7 7 15 13 2 0 13 2
5 7 3 13 9 2
15 0 3 0 1 9 2 15 3 1 9 15 9 0 13 2
7 0 10 13 9 0 13 2
9 13 3 15 3 1 9 9 13 2
13 0 3 9 0 9 10 0 13 9 10 13 13 2
31 7 3 1 9 15 0 13 9 2 3 9 0 13 2 3 13 7 13 9 10 0 0 2 16 13 3 3 3 3 3 2
11 3 3 15 13 9 9 3 15 0 9 2
13 3 3 9 3 13 2 9 13 9 7 9 0 2
9 0 3 2 0 0 2 13 3 2
13 9 3 15 15 9 0 13 13 2 16 13 15 2
8 13 3 0 0 2 7 13 2
7 15 2 9 15 13 9 2
14 13 3 3 13 9 0 7 13 1 9 0 9 9 2
8 15 3 0 0 15 9 13 2
4 9 3 13 2
13 0 3 10 3 3 3 10 3 3 0 13 9 2
8 7 1 15 0 3 13 9 2
7 15 3 9 15 13 9 2
10 3 3 10 9 7 1 0 15 13 2
7 3 13 2 16 13 15 2
7 3 1 15 0 13 0 2
7 3 3 13 1 9 13 2
9 3 3 2 1 0 13 0 9 2
7 3 3 13 9 13 9 2
25 15 15 13 2 0 1 9 9 13 10 0 9 2 7 1 3 9 13 0 3 9 0 9 9 2
8 3 13 13 0 9 9 13 2
16 13 3 13 3 0 9 9 13 13 2 3 3 0 13 9 2
35 3 16 15 13 9 2 10 13 3 9 13 9 9 3 0 1 9 13 2 3 9 2 3 3 0 9 13 2 7 3 1 9 0 13 2
14 13 3 3 15 15 0 9 2 16 0 0 13 13 2
10 13 3 13 3 3 9 13 10 9 2
10 15 3 9 0 9 13 0 9 13 2
3 9 13 2
4 13 9 1 2
5 3 15 3 13 2
8 3 3 13 3 3 9 13 2
9 3 1 9 2 7 3 13 13 2
4 15 3 13 2
6 3 3 9 15 13 2
8 15 3 13 0 1 9 13 2
6 13 9 3 13 13 2
8 13 3 15 3 3 13 9 2
10 7 3 3 3 15 3 13 13 3 2
6 15 13 9 7 13 2
6 13 3 0 9 13 2
9 13 3 13 3 13 3 13 13 2
3 13 3 2
7 13 3 3 3 13 13 2
7 15 0 3 13 10 0 2
11 3 15 0 15 13 9 15 10 9 9 2
3 3 13 2
12 7 0 15 13 2 13 9 3 1 0 9 2
7 9 13 3 13 15 3 2
7 3 3 1 9 13 9 2
9 13 9 2 3 10 0 13 15 2
6 13 3 0 13 9 2
15 3 2 15 3 3 9 10 10 9 2 3 9 9 13 2
4 7 13 15 2
7 3 0 9 13 15 3 2
8 13 3 0 3 15 3 13 2
7 15 3 10 0 13 0 2
8 3 3 10 0 3 3 13 2
8 0 3 13 15 3 0 9 2
4 13 1 9 2
14 0 15 3 15 9 7 0 7 13 0 13 10 0 2
5 15 3 0 13 2
23 13 3 15 0 3 2 3 13 0 2 7 9 13 0 2 0 15 0 3 7 0 13 2
14 13 3 15 0 13 0 1 9 0 13 7 0 9 2
29 0 3 13 0 9 3 13 0 1 9 9 2 3 3 9 13 9 2 16 15 0 7 9 13 7 0 9 9 2
9 3 9 13 3 13 3 0 0 2
10 10 3 0 9 13 7 13 10 0 2
23 15 3 7 9 9 7 0 9 1 9 0 13 2 0 9 13 7 13 0 7 9 9 2
34 3 3 10 3 13 9 0 9 13 15 1 9 2 15 10 0 9 13 13 9 9 7 9 2 15 0 3 13 0 2 13 9 9 2
14 15 9 0 13 1 9 13 0 9 2 7 3 13 2
20 1 3 15 3 0 13 2 7 0 15 13 15 13 13 3 10 0 9 13 2
9 10 3 0 9 13 3 3 13 2
11 1 3 3 15 0 0 13 3 3 13 2
8 1 3 15 13 10 9 13 2
9 3 0 0 1 0 9 9 13 2
12 1 3 0 0 0 3 7 0 13 1 0 2
14 7 3 3 3 10 0 9 13 2 13 15 0 9 2
16 0 9 3 13 3 3 3 2 16 15 13 2 9 13 0 2
14 7 9 3 15 9 9 13 0 9 0 9 13 9 2
6 13 3 3 0 9 2
10 7 13 7 9 0 7 9 0 9 2
15 0 3 9 3 0 13 1 0 9 2 0 13 9 0 2
5 15 3 9 13 2
12 3 3 10 0 0 0 9 0 13 9 13 2
9 15 3 13 10 9 9 15 9 2
6 3 3 13 9 0 2
6 9 3 0 9 13 2
10 9 3 13 15 10 0 0 9 13 2
22 0 13 9 0 9 0 3 3 0 2 10 0 9 1 13 2 15 10 0 9 13 2
5 6 13 10 13 2
14 0 9 13 2 0 9 13 0 9 9 7 9 0 2
9 3 3 3 15 0 13 13 9 2
14 15 15 3 3 13 1 9 2 15 3 13 3 13 2
8 0 13 9 0 9 1 0 2
13 13 0 9 13 1 15 13 2 15 9 0 13 2
17 0 3 1 9 13 0 9 3 13 2 7 3 0 0 9 13 2
14 10 3 13 0 9 2 15 0 13 2 0 9 13 2
9 7 16 13 2 3 3 13 13 2
24 0 3 3 2 16 13 15 9 2 13 2 0 13 0 9 13 2 7 0 1 0 13 13 2
7 15 3 3 13 13 3 2
4 3 0 13 2
5 3 13 3 13 2
24 9 0 2 3 13 1 10 9 2 0 3 13 15 13 1 0 2 15 3 10 13 13 13 2
22 3 3 3 13 13 10 9 2 0 3 9 0 13 0 15 3 3 0 0 16 3 2
9 3 13 0 3 0 1 0 0 2
13 13 3 15 7 13 16 2 1 9 9 15 13 2
8 3 3 13 15 13 15 13 2
8 15 3 3 9 10 0 13 2
6 13 15 10 13 9 2
7 0 13 9 3 9 13 2
19 0 3 0 9 2 3 0 9 3 13 2 0 13 13 9 9 13 0 2
6 15 2 13 7 13 2
15 15 15 0 3 1 9 13 13 9 3 3 15 13 9 2
7 7 3 3 0 13 9 2
11 15 3 13 1 15 0 2 3 3 13 2
9 15 13 13 2 15 3 13 0 2
9 7 10 3 3 3 13 13 9 2
15 3 3 13 0 13 3 9 2 9 9 2 0 3 9 2
31 9 3 13 1 9 9 15 9 13 2 10 3 9 1 2 10 3 1 9 2 13 9 0 2 0 1 0 9 13 13 2
26 3 13 3 1 9 3 2 0 3 3 1 9 13 2 7 0 9 7 13 9 2 13 9 2 13 2
15 1 3 9 9 13 13 0 9 2 9 3 9 13 9 2
8 7 10 3 13 0 0 9 2
22 3 15 10 0 13 9 2 16 3 13 0 10 13 9 2 13 1 15 9 13 3 2
14 15 3 3 13 9 0 2 15 3 0 3 13 15 2
14 1 3 0 3 7 0 9 15 3 3 9 13 13 2
9 7 0 0 9 13 9 3 13 2
20 3 3 1 15 13 0 9 0 9 2 0 2 1 0 9 0 0 13 13 2
8 7 0 13 7 15 13 0 2
7 0 3 3 7 13 13 2
7 0 3 10 15 13 9 2
9 7 3 13 9 0 15 13 9 2
12 9 13 7 13 7 10 3 9 13 13 13 2
4 15 3 13 2
4 3 3 13 2
3 9 13 2
10 7 10 3 13 9 2 15 3 13 2
4 9 13 13 2
3 7 13 2
9 3 3 15 9 1 15 13 13 2
4 3 2 13 2
13 13 3 13 15 10 15 9 2 0 3 13 13 2
7 6 3 13 0 13 3 2
7 13 3 9 16 3 13 2
3 0 13 2
13 3 0 0 13 9 2 0 10 9 10 9 13 2
20 13 10 0 2 10 0 2 10 1 0 0 9 2 1 0 15 9 0 9 2
5 3 0 13 9 2
8 6 1 9 13 7 13 3 2
7 15 3 3 13 1 13 2
10 3 3 13 3 0 16 3 3 13 2
8 1 3 9 0 7 13 13 2
8 13 3 15 2 3 3 13 2
4 9 0 13 2
6 3 13 3 13 0 2
9 7 13 0 2 3 15 13 13 2
8 15 3 13 13 15 15 13 2
9 7 15 10 9 0 9 0 13 2
5 3 15 3 13 2
4 3 13 13 2
5 0 15 13 13 2
6 3 3 0 3 13 2
14 3 15 13 3 3 16 13 13 13 2 0 15 13 2
13 15 3 3 13 3 0 0 13 9 10 0 0 2
10 3 3 13 7 3 13 15 7 3 2
5 0 3 0 13 2
19 15 9 3 15 1 0 9 10 0 9 13 9 1 9 13 0 9 13 2
28 15 3 10 0 9 2 10 0 1 9 9 13 3 0 9 3 3 9 0 9 13 0 2 0 0 3 13 2
6 3 0 3 13 13 2
23 16 13 9 10 9 10 15 1 13 13 9 9 15 2 3 3 15 0 13 0 1 15 2
14 3 3 0 9 9 0 9 13 2 9 15 13 9 2
22 16 3 15 9 7 9 0 9 13 10 0 2 3 3 3 9 1 0 9 3 13 2
27 3 3 10 9 0 0 9 3 15 1 0 9 13 0 13 2 13 0 9 2 3 1 15 9 13 9 2
10 0 3 13 13 2 0 3 3 0 2
13 16 3 15 9 13 2 13 3 10 0 10 0 2
6 7 3 15 13 13 2
19 15 3 9 13 2 13 3 15 9 9 2 13 3 9 0 7 9 15 2
15 0 1 9 2 0 13 9 0 3 9 2 9 0 13 2
18 3 15 13 3 13 0 13 10 9 1 2 15 0 13 9 9 0 2
5 3 13 9 0 2
19 7 3 13 1 9 9 2 13 0 0 7 13 15 0 2 3 0 13 2
8 7 3 3 9 3 13 3 2
4 3 13 0 2
13 15 3 1 9 9 13 13 13 13 10 3 13 2
11 3 3 13 0 9 9 15 0 9 13 2
11 7 7 3 13 7 3 13 10 0 13 2
4 0 13 9 2
14 13 3 3 7 13 9 0 9 13 2 15 9 13 2
14 15 3 0 3 13 9 2 16 15 13 1 9 9 2
5 3 3 13 9 2
10 9 3 3 13 3 7 0 3 9 2
44 3 2 16 10 0 9 13 2 3 13 10 0 2 7 15 13 1 3 0 9 9 3 10 0 2 15 13 15 2 16 15 13 9 0 13 10 0 1 0 2 0 13 15 2
26 15 3 13 15 7 13 13 2 0 13 15 10 3 9 9 13 0 1 1 9 10 0 0 13 9 2
9 7 15 0 9 9 13 9 13 2
17 13 10 9 9 2 15 0 13 9 2 0 9 1 0 9 13 2
4 0 13 15 2
15 15 3 9 13 2 15 3 0 9 0 7 10 0 9 2
11 15 3 3 13 1 15 15 13 1 15 2
19 15 3 15 9 13 9 2 7 9 0 9 10 13 3 13 9 0 9 2
9 15 3 15 13 3 1 15 9 2
6 1 15 0 15 13 2
5 7 13 15 9 2
8 9 9 3 13 10 13 3 2
15 15 3 13 9 3 13 2 3 3 13 3 0 0 9 2
7 13 3 3 10 15 9 2
16 3 3 9 13 1 3 15 2 16 0 10 13 3 13 13 2
10 13 3 15 9 10 0 2 16 13 2
7 3 3 9 3 0 13 2
5 7 15 15 13 2
8 13 3 3 13 9 15 15 2
9 7 3 15 2 13 0 3 13 2
7 13 9 7 9 15 13 2
10 15 3 3 3 1 15 3 13 15 2
8 13 15 13 0 0 3 13 2
7 3 3 3 3 9 13 2
8 15 3 13 3 3 9 13 2
6 13 13 7 13 9 2
7 3 3 13 9 15 3 2
16 13 3 3 0 3 15 13 9 2 16 3 13 0 15 3 2
12 3 3 0 0 1 9 9 13 13 13 9 2
6 7 13 3 3 0 2
15 3 15 7 3 0 3 13 13 2 7 0 15 13 0 2
20 7 3 13 1 0 2 13 15 16 9 13 1 0 2 0 1 0 2 13 2
21 0 9 9 9 1 15 13 9 3 0 3 2 16 3 0 13 2 0 9 13 2
8 10 3 0 9 0 15 13 2
18 7 3 9 10 9 15 3 13 7 9 13 2 3 3 0 9 13 2
3 13 0 2
6 13 13 15 10 9 2
8 3 3 15 13 9 15 13 2
4 6 3 13 2
15 7 15 1 10 0 9 7 9 13 2 16 13 15 13 2
4 3 3 13 2
11 3 13 15 9 16 0 13 13 9 3 2
3 0 13 2
4 10 13 13 2
5 15 3 3 13 2
5 0 3 3 13 2
5 3 13 3 9 2
5 1 9 2 13 2
12 0 15 9 13 2 16 0 9 3 13 13 2
14 7 15 0 9 13 0 2 6 15 2 0 9 0 2
10 15 13 3 3 3 0 13 1 9 2
10 3 3 3 9 9 0 0 9 13 2
12 0 10 0 0 9 13 3 0 7 13 13 2
14 3 13 0 0 2 7 13 10 0 9 10 0 9 2
19 15 3 2 15 10 0 13 3 2 9 9 3 13 9 1 15 10 9 2
11 13 3 15 0 1 0 9 3 0 13 2
19 7 13 1 3 9 7 0 9 2 16 3 9 13 0 9 0 13 9 2
23 13 3 9 3 3 0 13 2 13 15 9 0 2 0 9 2 9 13 3 3 15 13 2
8 7 0 9 9 3 13 3 2
19 15 3 1 15 9 0 13 1 9 9 0 2 3 15 0 13 0 1 2
13 7 13 0 10 9 9 2 0 0 9 3 0 2
13 3 10 0 13 3 9 13 2 13 3 9 13 2
6 9 13 2 16 0 2
10 3 3 10 0 7 10 0 0 13 2
8 0 3 0 9 13 0 9 2
11 13 3 9 0 9 10 0 9 9 13 2
8 0 3 9 9 13 13 9 2
7 15 3 3 3 13 13 2
31 13 3 3 16 10 3 0 15 1 15 0 2 3 3 13 3 2 1 3 10 0 0 13 13 13 2 7 3 3 13 2
9 10 0 3 9 0 13 9 9 2
7 7 1 3 0 3 13 2
7 15 3 13 3 3 0 2
7 13 9 2 0 3 13 2
6 3 3 15 13 13 2
16 0 3 1 9 13 9 9 10 0 0 15 13 1 0 0 2
7 13 0 9 1 9 9 2
24 0 10 0 9 13 2 0 0 13 3 2 7 3 1 0 9 13 9 3 9 0 3 9 2
7 9 13 3 0 1 9 2
10 0 3 13 9 13 10 0 0 3 2
38 13 3 3 0 1 9 13 13 2 3 9 13 3 3 0 13 15 3 2 15 10 13 9 13 0 13 2 16 3 13 10 3 3 9 0 13 13 2
12 3 1 0 13 3 3 9 9 0 13 9 2
12 13 3 9 13 15 3 9 9 1 9 9 2
11 7 15 9 3 2 13 2 16 13 15 2
8 10 9 3 0 13 13 9 2
15 0 15 13 10 15 10 9 13 13 7 2 13 15 0 2
7 15 3 13 9 15 13 2
15 7 13 3 2 1 10 0 13 9 2 9 16 13 9 2
14 0 13 9 9 0 0 2 16 15 9 3 13 13 2
7 15 3 13 15 9 13 2
6 0 13 7 13 13 2
14 13 3 0 15 9 0 0 9 9 2 3 13 13 2
24 10 3 0 0 9 13 0 1 9 9 13 10 9 2 15 9 9 13 3 3 1 9 13 2
12 0 3 1 9 3 13 0 3 13 13 9 2
6 15 3 3 0 13 2
6 15 3 3 3 13 2
10 15 3 3 1 0 13 0 13 9 2
4 15 13 9 2
22 3 0 0 9 2 3 13 15 13 1 0 9 0 13 2 3 13 0 0 3 9 2
13 15 3 9 0 9 13 9 2 3 1 9 13 2
14 3 16 13 15 9 2 3 3 13 0 1 9 0 2
5 0 10 9 13 2
14 10 3 3 1 9 13 15 15 13 15 9 9 13 2
13 16 3 13 2 3 13 9 0 2 16 9 0 2
9 13 3 1 9 0 16 13 15 2
14 15 15 3 0 2 3 13 0 0 2 1 9 13 2
14 15 13 9 2 3 13 13 9 15 9 15 13 15 2
3 3 13 2
18 3 13 10 0 9 2 9 3 16 2 0 16 13 2 3 13 1 2
11 0 13 9 13 9 0 3 3 13 0 2
10 3 3 13 9 2 1 15 13 15 2
4 13 0 3 2
8 15 3 9 0 9 13 13 2
11 13 3 3 9 13 7 10 0 9 13 2
3 3 0 2
8 3 13 15 3 3 3 13 2
15 13 2 13 2 3 9 9 13 13 9 3 15 13 13 2
8 13 0 2 3 9 13 0 2
8 9 3 9 7 9 3 13 2
12 13 3 1 9 0 10 0 2 0 9 0 2
14 13 3 0 3 13 15 2 0 15 9 1 9 13 2
4 3 3 13 2
8 13 3 15 3 0 9 13 2
34 13 15 15 9 2 0 9 9 13 2 0 16 15 13 13 15 1 0 9 2 7 3 1 0 15 13 3 13 9 0 9 3 9 2
16 3 3 0 2 15 7 13 9 2 13 0 9 1 0 9 2
15 3 0 9 0 13 3 2 7 0 10 9 1 9 15 2
7 3 15 3 3 13 13 2
5 9 9 9 13 2
8 3 3 3 3 3 13 15 2
6 0 13 15 13 9 2
5 9 3 13 15 2
15 3 3 3 3 3 10 1 9 13 9 9 3 13 13 2
30 15 3 3 15 2 15 3 0 9 13 0 9 2 7 15 9 9 7 0 0 9 2 10 0 16 3 13 13 13 2
6 15 9 0 13 9 2
4 15 3 13 2
11 9 15 15 3 0 13 2 0 9 0 2
7 15 3 3 13 9 0 2
10 1 3 15 9 0 15 9 0 13 2
12 15 3 10 0 0 2 10 0 0 2 13 2
3 3 0 2
32 3 15 0 9 13 15 3 2 16 0 3 2 15 3 0 2 13 13 13 3 1 9 1 3 0 9 13 9 1 0 9 2
5 6 2 15 13 2
5 15 15 13 0 2
14 3 0 3 2 16 13 2 13 2 13 9 15 13 2
13 0 15 0 7 13 13 0 0 9 0 1 9 2
11 15 3 13 0 13 2 15 3 3 13 2
2 13 2
11 6 2 0 0 13 0 9 9 15 9 2
4 7 13 9 2
9 3 3 15 13 3 3 9 13 2
6 3 0 3 9 13 2
9 15 3 3 13 13 0 10 15 2
16 3 3 2 16 13 3 2 13 2 13 3 13 1 9 9 2
14 10 3 0 9 0 9 13 3 13 2 3 15 13 2
11 15 0 13 7 0 0 2 0 3 0 2
7 15 3 15 13 3 1 2
9 9 13 0 2 3 0 2 3 2
7 1 0 9 1 0 13 2
14 9 3 0 3 13 2 7 15 13 9 7 9 13 2
2 13 2
11 9 3 13 9 13 13 9 15 0 9 2
13 15 3 9 10 15 2 3 15 9 13 10 9 2
17 3 0 9 3 0 13 3 2 16 15 7 0 9 9 0 13 2
6 13 2 13 2 13 2
8 10 13 3 13 0 13 13 2
14 0 3 15 9 3 9 15 13 0 0 16 13 13 2
13 15 13 0 3 3 13 13 2 3 3 13 13 2
10 13 2 13 2 16 13 10 0 0 2
4 0 15 13 2
16 0 9 0 2 1 9 0 2 13 2 1 0 1 9 13 2
12 9 3 0 9 13 2 9 9 1 0 13 2
7 3 0 0 15 13 13 2
5 6 2 15 13 2
5 3 15 13 0 2
10 13 16 9 13 15 9 3 13 13 2
10 13 2 1 9 2 10 9 12 9 2
21 9 3 2 15 3 15 13 1 2 9 13 0 1 9 13 3 2 16 13 9 2
12 0 3 0 15 9 13 1 15 13 0 9 2
15 15 3 3 7 0 7 10 0 3 13 3 9 13 9 2
16 15 3 3 15 13 1 9 0 2 0 3 0 13 15 15 2
16 3 13 3 2 7 3 13 9 13 10 9 15 15 13 3 2
16 13 3 0 9 2 7 3 3 0 13 15 3 0 13 9 2
8 15 3 13 15 9 13 9 2
2 13 2
6 15 9 15 13 9 2
7 3 3 13 15 9 13 2
12 15 9 0 13 9 3 13 2 16 13 9 2
27 16 3 9 15 15 9 13 2 15 3 3 15 15 15 13 9 13 3 13 0 9 2 0 3 3 13 2
13 3 3 13 9 10 15 9 1 9 7 9 13 2
7 1 0 9 0 13 9 2
20 16 3 13 3 2 13 13 2 3 13 3 13 2 16 3 13 2 9 13 2
12 3 3 13 3 9 3 13 13 3 13 0 2
12 3 0 1 9 13 9 9 13 10 13 13 2
35 3 3 3 3 3 3 1 9 9 3 13 3 2 3 3 13 9 2 3 3 3 9 3 3 13 3 2 9 9 9 3 3 9 13 2
17 7 9 13 2 16 9 13 0 2 13 13 3 16 1 0 0 2
13 9 3 15 13 9 3 3 2 9 13 15 13 2
22 3 3 13 13 3 15 13 13 2 0 13 10 9 9 3 1 0 13 1 9 13 2
20 7 13 15 3 9 15 0 2 7 3 13 13 3 13 3 13 3 3 13 2
4 13 3 0 2
13 3 0 13 0 9 2 3 3 15 0 3 13 2
16 3 15 13 15 3 13 2 16 3 15 13 0 1 9 13 2
17 3 13 1 9 3 2 3 15 13 13 15 9 0 3 0 13 2
7 3 0 13 3 0 13 2
5 3 15 13 15 2
11 3 3 15 9 13 13 15 15 13 3 2
8 9 13 13 2 3 15 13 2
14 9 0 3 13 2 3 0 9 2 3 9 13 3 2
11 7 15 13 13 7 10 0 9 13 0 2
23 15 3 2 3 3 15 13 3 0 9 2 1 9 15 13 3 2 3 10 0 13 9 2
6 3 3 13 10 9 2
26 1 0 0 3 9 13 7 10 9 13 2 10 3 0 9 3 3 13 2 7 3 13 0 3 13 2
9 3 3 3 0 9 1 0 13 2
11 10 0 3 3 2 16 0 13 2 13 2
7 10 9 13 3 0 13 2
7 3 3 0 10 9 13 2
9 0 3 15 13 2 9 16 13 2
7 16 0 13 15 3 13 2
9 10 9 15 10 9 3 0 13 2
8 1 10 0 3 0 13 13 2
9 0 3 13 2 16 3 13 13 2
9 9 3 13 15 2 15 3 13 2
8 3 3 13 9 2 9 13 2
7 15 3 3 13 9 9 2
8 3 15 3 9 0 13 3 2
3 13 13 2
5 3 15 0 13 2
6 9 3 0 0 13 2
10 1 10 9 2 3 15 2 15 13 2
8 0 3 3 3 15 13 0 2
7 0 1 9 9 13 15 2
4 9 15 13 2
5 15 13 3 0 2
6 7 13 0 16 13 2
36 3 3 13 9 15 9 0 9 13 9 10 13 2 15 9 3 3 3 13 2 3 1 0 9 13 2 7 1 9 13 13 13 15 13 9 2
22 3 3 3 15 3 10 0 0 9 0 9 3 3 15 13 0 9 13 10 0 9 2
16 15 3 3 9 13 9 0 2 15 1 0 13 10 15 3 2
13 3 0 13 15 0 15 9 3 0 13 0 9 2
7 16 3 13 2 13 13 2
6 0 0 9 13 13 2
17 13 3 3 15 2 13 2 3 15 13 2 0 3 0 16 15 2
3 3 13 2
2 13 2
3 13 3 2
6 13 0 9 15 9 2
29 16 3 15 9 9 15 13 15 10 9 2 0 3 0 13 9 2 9 0 9 13 2 3 7 15 15 13 9 2
27 15 3 0 1 15 13 0 9 9 2 10 0 3 15 0 9 9 13 1 10 0 9 2 0 9 9 2
20 13 0 9 13 0 7 10 0 9 0 9 2 15 0 13 9 9 0 9 2
5 0 3 13 9 2
7 9 3 9 13 2 6 2
16 13 3 2 0 3 2 3 0 9 13 9 2 0 9 9 2
14 3 3 3 3 0 9 13 15 9 7 9 0 9 2
7 3 3 0 13 0 9 2
9 15 15 2 15 3 3 9 13 2
19 13 7 0 13 9 9 0 2 0 1 9 9 2 10 0 16 13 9 2
7 0 3 13 0 13 9 2
14 15 3 10 0 9 13 15 13 1 15 3 3 13 2
6 0 13 9 3 0 2
8 3 3 0 9 13 1 15 2
45 0 13 10 0 9 9 0 13 3 2 16 3 13 1 9 0 2 3 13 3 15 3 3 13 13 15 10 0 13 9 2 7 3 15 7 0 13 3 7 1 9 13 10 13 2
27 1 15 3 10 9 3 3 3 9 13 3 0 9 2 16 10 9 13 13 7 15 3 1 10 3 13 2
5 7 0 15 13 2
17 3 3 10 0 3 3 0 9 0 2 7 10 13 3 13 3 2
13 0 3 9 9 1 0 7 9 0 1 9 13 2
16 7 15 13 0 15 10 9 13 3 2 16 3 9 13 15 2
13 15 9 3 13 2 7 3 9 2 13 13 13 2
3 3 13 2
21 3 13 15 13 9 0 15 13 9 3 0 2 15 1 15 1 15 13 10 0 2
8 15 3 13 3 3 13 15 2
7 10 0 3 9 3 13 2
7 3 15 0 9 13 13 2
8 0 3 0 15 13 0 13 2
7 7 13 3 0 0 13 2
4 15 0 13 2
18 3 15 13 10 13 15 2 15 3 13 2 3 15 3 2 13 9 2
7 3 15 0 0 13 0 2
14 3 13 15 9 3 15 13 9 0 13 9 0 9 2
6 0 13 15 13 9 2
10 0 3 15 9 0 2 13 9 9 2
28 3 3 0 1 9 12 13 3 13 15 1 9 2 15 3 15 15 1 9 13 13 0 2 3 3 13 13 2
16 3 3 15 13 2 0 16 13 3 2 13 15 12 3 13 2
11 1 0 13 3 0 2 7 3 10 0 2
18 3 16 15 13 15 2 13 3 3 0 13 3 16 2 1 15 0 2
10 3 3 13 9 9 15 1 0 9 2
11 15 3 9 9 13 13 0 13 9 0 2
3 13 0 2
6 13 3 13 0 15 2
10 15 3 15 13 2 3 3 9 13 2
15 3 13 13 15 10 9 9 0 2 7 1 9 13 15 2
12 13 3 13 0 0 15 9 0 16 3 13 2
2 13 2
16 3 3 13 3 3 3 13 2 16 0 15 15 0 0 13 2
3 13 3 2
12 10 9 15 1 9 3 13 0 3 3 13 2
14 3 3 10 9 15 3 13 15 13 3 10 9 13 2
43 15 3 13 3 0 0 9 2 1 15 2 13 10 0 9 2 7 0 3 13 15 15 15 3 13 3 2 3 3 13 9 9 13 0 0 2 0 9 13 2 1 9 2
8 3 3 3 3 3 13 15 2
12 3 3 15 0 2 7 10 9 9 13 3 2
8 13 3 2 3 13 13 0 2
8 3 3 13 3 13 15 13 2
9 13 10 0 9 13 15 1 9 2
2 13 2
6 13 3 10 0 13 2
7 13 0 9 10 9 13 2
9 15 0 9 2 7 0 3 13 2
4 15 3 13 2
5 0 3 13 9 2
8 13 3 9 15 10 9 0 2
7 15 13 3 15 13 0 2
7 0 13 3 13 9 15 2
7 15 15 0 15 9 13 2
8 13 3 15 10 9 13 13 2
6 3 3 0 3 13 2
8 3 0 0 0 9 0 13 2
10 15 3 15 3 13 16 2 15 13 2
8 0 3 9 2 3 0 13 2
9 3 3 13 2 3 0 3 13 2
27 3 3 3 3 0 13 16 15 15 3 13 3 15 3 0 9 2 0 3 3 3 13 15 3 0 13 2
7 15 3 13 13 15 13 2
17 7 3 3 9 1 15 13 2 0 3 0 13 2 15 13 0 2
19 7 10 13 15 13 13 7 13 7 9 13 0 13 10 0 9 13 9 2
36 0 3 13 0 0 9 0 13 9 2 3 3 13 13 13 15 13 13 0 2 3 10 9 0 13 0 3 10 0 13 0 0 13 9 1 2
25 3 15 9 15 10 13 9 0 3 9 7 0 9 0 3 13 2 3 13 10 9 9 13 3 2
16 10 3 0 3 13 2 16 15 9 13 13 2 0 9 13 2
6 15 3 0 0 13 2
9 15 3 9 1 15 0 13 13 2
4 3 13 3 2
16 16 3 3 2 13 15 0 13 15 15 2 13 13 10 0 2
6 3 3 0 13 9 2
18 7 15 3 0 9 9 13 2 15 3 0 9 0 9 0 13 0 2
11 0 3 1 9 9 9 10 0 9 13 2
9 3 3 0 9 3 13 0 9 2
32 3 3 0 2 0 15 9 13 13 2 13 2 13 2 15 9 13 10 0 0 0 3 0 0 9 2 7 13 2 3 13 2
8 2 3 0 9 13 13 13 2
14 9 3 3 3 9 13 2 3 3 9 3 7 9 2
10 0 3 3 13 15 7 3 13 9 2
19 10 3 0 9 13 9 13 1 3 9 0 9 2 1 9 3 0 9 2
27 9 3 3 3 13 15 15 3 3 15 9 13 0 2 9 3 0 1 3 9 9 13 1 3 9 9 2
33 15 3 13 9 0 13 0 9 9 15 13 2 7 0 1 15 0 13 0 3 3 13 2 7 9 9 13 13 3 15 13 9 2
14 9 3 10 0 3 13 13 3 1 0 7 13 0 2
6 7 9 15 13 9 2
15 9 3 7 10 3 0 9 13 15 2 7 3 0 13 2
20 3 3 13 16 13 0 2 7 13 2 16 15 3 13 15 15 1 0 13 2
26 10 3 3 15 9 1 9 13 0 1 0 0 0 2 10 3 0 9 9 3 15 7 15 3 13 2
11 15 3 3 13 13 9 0 2 0 13 2
10 7 15 9 3 13 9 13 15 13 2
10 10 3 13 3 13 0 10 13 9 2
17 16 3 13 2 3 15 0 7 13 3 13 0 0 3 13 9 2
14 7 1 0 15 3 13 15 3 3 9 13 13 15 2
10 3 3 3 9 0 3 13 0 9 2
3 3 13 2
16 13 3 7 10 0 2 16 13 1 0 13 2 0 3 13 2
5 13 3 0 9 2
14 3 3 3 0 3 3 3 13 13 10 3 3 9 2
4 1 0 13 2
13 15 3 0 13 10 9 16 7 10 0 9 1 2
8 13 3 0 13 10 9 1 2
20 13 15 9 3 9 9 9 2 3 13 9 1 15 2 13 3 3 0 13 2
7 0 3 9 15 13 9 2
3 13 13 2
6 3 3 13 3 3 2
11 0 13 3 13 3 10 9 9 13 15 2
6 15 3 13 15 9 2
8 15 15 13 9 0 0 9 2
5 1 15 13 9 2
16 9 2 3 13 2 13 2 3 1 9 3 13 2 16 13 2
16 3 3 9 15 3 3 9 9 13 2 15 15 13 13 3 2
13 9 3 0 3 13 13 2 9 0 16 13 9 2
14 9 13 13 3 0 9 13 15 2 7 1 9 9 2
19 3 3 10 9 2 16 15 7 1 9 13 3 2 1 15 3 9 13 2
4 13 0 13 2
9 9 3 13 0 0 1 0 13 2
13 0 3 0 3 2 9 3 13 2 13 0 13 2
12 10 0 9 15 1 9 13 13 15 0 13 2
8 7 1 9 3 0 15 13 2
14 3 3 9 2 3 3 15 1 10 13 15 13 9 2
14 1 3 3 10 3 0 2 7 0 0 0 13 9 2
16 15 3 13 0 10 13 2 3 3 15 3 0 9 13 13 2
6 0 13 3 15 13 2
10 7 3 0 1 10 9 13 7 13 2
10 15 3 9 7 3 13 15 15 13 2
14 9 3 10 13 15 9 1 9 7 13 7 9 0 2
15 13 3 15 0 9 2 3 3 1 9 9 15 15 13 2
15 3 3 3 0 0 9 13 3 3 9 0 9 13 9 2
17 0 3 3 0 13 15 0 9 0 0 9 13 9 1 0 9 2
5 15 9 0 13 2
9 0 3 9 1 9 0 13 3 2
12 13 3 16 15 9 13 2 0 1 9 13 2
2 13 2
21 15 3 13 2 0 16 13 9 13 13 10 9 3 13 2 9 13 3 9 0 2
13 15 0 3 10 9 15 13 2 0 3 10 13 2
10 16 3 13 2 9 13 0 1 0 2
7 13 3 0 3 0 0 2
5 9 3 13 0 2
15 16 3 3 15 0 13 1 0 9 10 9 2 7 13 2
25 16 3 3 13 2 7 15 7 0 13 13 9 7 0 15 2 1 15 13 2 0 13 13 15 2
15 15 3 3 15 15 3 9 10 3 9 15 13 0 13 2
21 13 3 10 13 2 3 15 9 13 13 3 0 1 2 0 3 15 0 13 9 2
21 15 3 0 0 13 13 2 1 3 15 10 9 3 15 3 9 3 3 3 13 2
27 3 3 16 3 13 10 9 3 0 2 0 15 13 13 3 13 2 9 3 0 9 3 13 2 7 13 2
10 3 3 1 10 0 9 13 10 9 2
35 1 15 15 15 2 3 0 9 2 13 1 0 13 2 13 10 9 10 9 13 2 10 0 9 9 3 7 10 3 9 10 3 3 9 2
28 7 0 10 7 13 13 9 3 9 0 9 13 15 3 3 9 9 2 7 10 9 10 3 13 3 15 0 2
22 15 3 10 0 0 2 0 15 13 13 2 10 3 0 9 10 0 3 13 3 9 2
11 3 3 13 3 3 3 10 13 13 13 2
3 0 13 2
13 7 13 9 15 7 13 3 3 3 9 13 9 2
9 10 0 1 15 3 13 0 13 2
12 16 7 0 13 2 7 13 10 7 3 13 2
9 7 3 1 0 3 3 0 13 2
7 13 3 9 13 0 9 2
6 3 3 7 0 13 2
5 0 3 13 9 2
6 13 13 1 15 9 2
3 13 15 2
6 10 3 13 0 13 2
5 7 13 0 13 2
15 15 3 10 0 3 9 3 13 2 15 0 13 9 0 2
34 9 3 2 16 15 7 13 10 9 2 13 15 13 2 9 0 3 13 15 15 9 2 16 10 13 9 13 3 13 7 9 9 13 2
5 1 15 3 13 2
7 0 3 3 15 13 13 2
6 3 3 3 3 13 2
4 15 3 13 2
4 3 0 13 2
5 13 15 1 9 2
14 3 3 10 0 3 15 15 13 0 2 16 15 13 2
18 3 3 0 13 3 3 0 9 15 2 15 15 13 2 15 13 9 2
12 13 3 3 3 15 10 0 9 13 1 9 2
5 0 3 3 13 2
17 15 3 3 7 3 0 2 16 3 13 7 10 0 2 13 0 2
3 15 13 2
12 13 3 13 2 7 13 15 13 7 13 9 2
9 15 3 3 15 3 3 15 13 2
5 15 0 3 13 2
6 3 3 3 13 15 2
17 9 13 10 0 2 10 0 3 3 13 3 13 2 7 15 13 2
17 15 3 0 3 3 3 13 9 13 2 15 3 15 15 13 9 2
9 13 3 0 2 16 15 9 13 2
5 3 3 3 13 2
12 1 15 2 16 13 2 13 1 9 15 0 2
13 7 3 13 3 0 2 3 9 13 2 15 13 2
15 13 3 13 15 7 13 9 13 3 2 0 7 9 13 2
25 13 15 10 9 15 13 13 2 1 9 10 3 13 3 15 3 15 2 3 13 9 15 0 9 2
7 3 3 13 15 15 9 2
6 7 3 15 13 13 2
2 13 2
5 0 3 13 13 2
7 15 3 15 0 13 13 2
7 13 3 2 16 3 13 2
4 3 13 3 2
4 7 3 13 2
8 9 15 13 9 15 13 13 2
9 7 3 15 13 3 3 9 13 2
9 13 15 3 0 2 16 13 0 2
16 13 15 13 1 10 0 3 13 2 3 3 13 7 13 0 2
8 3 7 13 0 3 13 13 2
6 7 13 2 1 15 2
18 15 3 0 3 13 16 0 10 3 9 15 3 9 15 3 9 13 2
19 0 13 1 9 2 16 3 15 3 0 2 15 9 13 2 13 3 3 2
16 3 3 2 16 10 9 3 13 9 2 13 15 15 9 0 2
14 3 10 3 9 3 13 13 9 13 2 7 9 13 2
13 15 3 15 13 13 2 13 9 13 10 0 3 2
10 13 13 15 7 15 10 13 15 13 2
5 15 3 15 13 2
10 3 3 15 15 13 9 2 7 9 2
9 13 3 2 16 7 0 15 13 2
20 15 7 13 3 13 3 13 0 2 3 3 3 13 2 3 3 15 13 1 2
6 3 13 1 15 13 2
38 7 13 0 13 10 0 0 1 1 9 3 2 7 15 9 9 3 7 10 0 9 13 3 1 9 15 9 9 2 13 3 3 0 2 3 3 9 2
17 0 3 9 3 13 0 2 15 15 13 15 3 7 10 0 9 2
9 1 0 7 9 7 0 9 13 2
10 15 3 3 13 9 0 15 13 3 2
8 3 3 0 9 15 13 13 2
17 3 3 15 15 13 0 13 2 16 9 15 3 9 10 0 13 2
20 15 15 13 2 16 3 15 13 2 0 2 9 3 2 15 15 13 2 0 2
7 15 9 13 15 7 13 2
7 6 0 3 0 0 13 2
7 3 15 0 0 13 13 2
8 0 13 2 15 15 13 0 2
8 0 3 3 15 10 9 13 2
10 7 16 9 15 13 2 3 15 13 2
3 13 3 2
3 13 3 2
7 3 3 13 3 15 13 2
4 13 3 15 2
33 10 9 0 2 15 3 13 13 13 9 10 0 2 0 13 3 2 0 9 9 2 3 3 0 13 0 2 3 3 13 10 9 2
15 0 3 1 13 7 0 1 0 0 1 9 13 9 13 2
27 13 3 9 10 0 13 9 0 7 9 2 1 15 13 9 9 7 9 2 7 10 9 0 3 7 9 2
6 7 0 13 3 13 2
11 16 13 13 2 13 15 3 0 9 13 2
18 0 3 1 0 13 9 7 9 10 9 9 2 0 3 3 13 9 0
14 13 3 10 0 3 13 9 9 10 0 9 0 13 2
22 13 3 1 0 9 1 3 9 7 9 0 0 0 9 13 2 10 0 9 13 9 2
6 15 3 3 13 13 2
15 0 3 3 2 0 13 0 9 3 3 13 3 3 13 2
6 15 15 13 3 13 2
7 9 3 3 9 13 9 2
14 7 3 15 3 2 16 13 0 9 2 13 3 13 2
30 3 3 1 0 10 9 15 10 9 0 13 2 7 1 0 2 16 0 3 1 9 2 0 3 1 15 7 0 13 2
15 7 13 3 3 0 9 3 3 9 13 3 16 9 9 2
16 9 3 13 2 10 0 9 16 13 10 9 10 9 0 13 2
10 13 3 15 2 13 3 3 9 15 2
13 1 9 3 0 3 1 0 9 13 9 0 15 2
3 3 13 2
8 0 3 15 3 9 1 13 2
4 13 16 13 2
11 1 10 13 0 13 2 3 13 0 13 2
8 0 3 7 0 15 13 15 2
9 0 0 3 15 0 13 3 13 2
16 16 3 13 9 10 9 13 15 10 9 3 2 3 3 13 2
16 16 3 13 9 0 3 13 3 13 10 9 2 3 3 13 2
6 13 15 0 0 13 2
15 13 7 3 13 2 16 13 15 1 10 9 9 13 15 2
8 7 3 3 0 13 10 9 2
4 3 3 13 2
5 0 13 0 9 2
7 0 0 3 3 13 9 2
10 3 3 10 9 0 13 1 10 9 2
9 13 3 15 15 10 3 1 9 2
7 7 3 9 10 13 13 2
6 13 2 3 3 3 2
3 3 13 2
10 3 3 3 0 10 0 3 13 15 2
3 3 13 2
9 15 3 13 7 13 3 3 13 2
8 16 3 13 3 2 3 13 2
8 16 3 13 15 2 0 13 2
11 15 3 15 13 13 0 15 15 15 3 2
2 13 2
6 3 3 3 9 13 2
6 9 10 0 13 13 2
6 9 3 13 15 13 2
8 13 3 0 0 9 0 13 2
7 15 13 13 0 15 13 2
7 3 13 15 15 12 0 2
8 3 3 3 7 0 13 0 2
22 15 3 3 3 3 0 13 13 9 13 3 16 9 13 2 3 3 0 15 13 13 2
20 3 3 3 1 15 0 1 9 13 2 16 3 0 13 2 0 7 9 13 2
12 3 3 15 9 0 13 9 0 7 9 13 2
13 3 15 13 13 16 0 13 16 10 1 9 0 2
16 3 0 13 2 3 15 0 13 2 3 10 15 13 13 15 2
8 10 3 13 0 0 3 1 2
9 3 3 15 0 3 13 13 15 2
8 3 3 13 9 0 3 13 2
18 7 3 3 9 15 10 9 13 3 3 3 1 0 13 3 13 3 2
15 7 15 9 0 3 3 13 13 10 13 16 3 13 15 2
8 9 3 0 7 15 3 13 2
14 7 1 9 13 15 3 2 16 9 0 9 13 0 2
8 0 3 7 1 9 13 0 2
13 16 0 15 13 3 13 2 0 13 15 13 3 2
4 15 3 13 2
7 13 2 3 13 15 13 2
8 3 3 13 3 3 13 13 2
7 3 3 13 15 3 13 2
6 7 1 0 13 0 2
4 7 13 0 2
8 15 9 13 2 3 15 0 2
2 13 2
19 7 3 13 2 7 0 2 16 15 15 13 2 13 2 15 13 15 13 2
6 15 15 13 3 13 2
12 15 3 3 3 0 3 3 1 9 0 13 2
5 13 3 15 13 2
2 13 2
5 13 3 15 13 2
17 3 3 13 2 0 16 13 2 15 13 9 7 9 1 15 9 2
19 7 15 0 9 9 13 9 2 15 16 0 0 13 10 3 10 1 15 2
17 15 3 3 13 2 16 13 15 3 13 7 9 0 15 13 9 2
12 10 3 0 2 3 15 15 2 13 9 0 2
7 0 3 3 3 13 13 2
13 0 3 13 0 13 2 0 3 2 16 9 13 2
10 10 3 0 9 0 3 13 0 13 2
6 3 15 13 3 13 2
12 13 2 15 3 13 9 2 1 3 15 0 2
5 7 15 13 9 2
14 3 15 2 3 2 9 13 2 13 3 13 3 13 2
15 13 3 13 2 0 13 9 9 2 0 13 7 13 9 2
2 13 2
9 13 2 16 3 10 9 13 13 2
6 9 15 13 9 13 2
7 13 3 15 9 15 0 2
17 7 15 3 2 3 3 10 9 2 0 3 9 13 1 0 0 2
21 9 3 9 3 13 9 12 2 7 15 9 0 13 9 13 0 9 0 1 9 2
19 3 9 3 3 0 13 9 13 9 3 3 9 10 0 13 1 9 13 2
11 15 3 3 9 9 13 2 3 0 13 2
6 9 9 0 13 13 2
9 13 3 0 3 3 3 13 13 2
16 9 3 10 9 13 2 0 3 9 1 0 9 1 9 13 2
7 7 15 9 15 13 13 2
15 3 15 1 7 15 15 13 9 9 13 2 0 13 9 2
4 3 15 13 2
14 10 3 9 9 15 13 13 2 15 3 9 9 13 2
10 13 15 1 9 0 13 3 3 13 2
3 3 13 2
8 3 13 16 13 10 9 13 2
9 13 3 3 2 16 9 13 3 2
12 7 3 13 3 2 15 3 3 13 13 13 2
13 0 13 0 7 0 13 9 9 2 0 9 9 2
10 12 13 10 0 2 1 3 0 13 2
6 9 3 13 9 0 2
7 3 1 9 13 3 13 2
34 1 15 3 3 13 7 9 15 3 13 13 9 3 13 2 13 10 0 9 13 9 15 13 1 9 9 2 3 0 13 15 0 9 2
4 13 15 15 2
12 0 3 0 9 0 13 13 15 7 0 9 2
9 3 3 13 3 15 1 9 3 2
2 13 2
6 7 1 15 0 13 2
4 7 13 3 2
11 3 7 13 3 2 1 0 9 15 13 2
15 15 3 3 7 0 13 3 16 15 2 1 9 15 13 2
12 15 9 3 9 13 0 2 9 3 9 9 2
26 13 3 9 9 0 10 3 2 16 15 9 15 13 2 13 3 0 2 9 3 3 10 0 3 0 2
18 15 13 10 3 13 9 3 13 2 0 3 13 3 9 9 3 13 2
10 15 3 3 9 13 10 13 10 9 2
13 15 15 3 0 13 2 3 3 13 15 3 0 2
4 13 3 0 2
14 1 9 15 10 3 9 0 3 10 9 1 9 13 2
18 7 15 10 9 16 13 2 9 13 13 2 0 9 0 9 15 13 2
19 3 3 0 3 13 2 7 3 9 13 1 15 9 0 0 9 3 13 2
5 13 3 10 0 2
17 16 3 10 0 0 13 9 15 0 2 15 15 3 9 13 0 2
7 15 0 3 3 13 9 2
20 15 7 0 13 3 3 9 15 9 13 3 3 13 15 2 13 3 1 9 2
4 3 13 0 2
16 3 3 1 0 0 9 15 3 13 1 9 15 3 13 9 2
12 16 3 3 3 1 10 13 13 2 13 9 2
4 15 13 15 2
12 16 3 13 13 15 0 2 15 3 13 9 2
7 0 3 15 0 13 9 2
10 3 3 13 3 9 3 10 0 0 2
16 16 3 9 9 0 13 2 3 0 13 3 9 1 15 13 2
16 7 3 13 3 9 3 13 2 3 13 0 0 3 13 3 2
10 9 3 13 2 3 15 0 2 15 2
15 3 15 3 0 3 10 0 3 13 2 7 0 3 13 2
3 3 13 2
12 7 3 10 9 13 15 13 3 3 0 13 2
3 13 13 2
5 7 13 1 9 2
10 0 3 3 13 3 15 3 15 0 2
42 7 15 13 13 9 10 0 9 9 9 3 0 2 15 9 13 9 2 0 1 9 13 2 15 9 9 0 2 3 3 15 0 9 9 13 3 3 7 3 9 13 2
8 0 1 0 9 3 3 13 2
4 9 13 9 2
11 10 3 3 13 9 9 3 13 9 13 2
7 9 3 13 3 9 13 2
12 15 3 3 1 15 9 9 9 13 9 13 2
12 16 3 10 15 9 0 2 15 13 15 13 2
28 3 10 0 13 9 1 9 13 2 3 3 1 10 9 9 3 3 10 9 2 16 7 15 0 0 13 9 2
13 13 3 9 0 0 13 3 2 3 9 9 0 2
5 13 3 10 0 2
9 3 3 13 9 9 3 9 0 2
15 7 0 3 7 1 0 3 13 2 0 3 13 0 9 2
7 0 3 13 10 9 1 2
10 7 13 15 13 13 15 15 13 13 2
18 10 3 9 13 3 2 13 3 2 3 3 3 3 2 13 3 3 2
4 15 3 13 2
6 0 9 3 13 0 2
12 9 0 0 9 10 0 13 2 16 13 3 2
3 3 13 2
8 16 7 13 0 2 13 13 2
22 0 9 3 13 10 9 13 16 13 2 7 3 15 1 10 9 13 3 3 15 1 2
15 13 9 15 2 7 13 13 10 0 3 13 10 9 9 2
10 0 3 15 3 13 7 15 15 13 2
6 0 15 15 9 13 2
14 16 0 0 13 15 13 3 2 3 13 0 0 13 2
6 0 0 9 13 9 2
9 9 10 0 2 3 13 2 13 2
13 10 3 3 13 13 9 13 1 9 9 0 15 2
7 3 15 15 0 13 3 2
2 13 2
6 15 3 10 9 13 2
9 7 3 3 0 9 1 9 13 2
10 7 3 10 9 3 13 9 15 13 2
17 15 3 3 13 9 15 15 10 9 13 2 9 3 13 15 0 2
9 0 3 3 1 9 9 9 13 2
12 7 0 15 1 0 13 2 3 10 9 13 2
7 0 3 7 9 13 1 2
9 15 3 13 0 15 1 9 13 2
18 13 3 15 9 3 13 13 9 15 10 3 0 9 9 10 0 13 2
10 15 7 10 9 1 15 3 3 13 2
8 3 3 15 13 3 13 9 2
9 7 3 9 3 3 0 13 15 2
8 7 3 13 10 13 3 3 2
8 3 13 3 1 9 0 13 2
3 3 13 2
6 3 3 9 13 15 2
11 7 3 15 13 3 3 0 3 3 15 2
8 7 1 15 3 9 15 13 2
8 3 3 1 0 9 13 0 2
7 10 3 3 0 13 9 2
9 15 3 13 7 13 15 0 13 2
8 13 3 1 15 15 10 9 2
5 3 0 9 13 2
7 9 3 13 1 9 9 2
8 15 3 9 13 9 15 13 2
7 9 3 9 13 10 0 2
7 13 15 13 0 9 9 2
6 0 3 9 9 13 2
2 13 2
3 3 13 2
8 10 13 3 0 15 0 13 2
11 3 3 1 0 15 13 3 3 0 13 2
8 3 2 7 9 0 13 15 2
5 3 13 13 9 2
6 15 9 3 15 13 2
6 0 9 0 13 9 2
10 3 13 3 13 0 2 16 13 15 2
7 15 3 0 13 3 0 2
22 13 15 15 10 13 3 2 15 13 10 9 15 13 2 7 3 1 9 7 3 13 2
8 13 2 16 10 9 13 15 2
14 13 3 0 0 16 15 1 9 2 15 13 3 13 2
10 3 15 3 15 3 0 3 9 13 2
4 15 0 13 2
3 9 13 2
9 10 3 13 13 3 3 13 3 2
14 7 1 9 2 16 15 10 15 9 13 2 13 0 2
2 13 2
15 15 3 3 3 3 16 0 15 9 13 0 2 13 0 2
4 7 13 15 2
9 3 3 13 7 3 15 13 3 2
10 7 3 13 3 3 10 0 15 13 2
8 10 0 3 0 15 13 3 2
8 13 15 13 3 10 9 15 2
7 0 3 13 0 13 9 2
12 0 3 15 13 0 13 2 0 3 3 0 2
4 0 13 13 2
12 0 3 15 2 16 0 13 2 9 13 13 2
13 15 3 15 9 10 9 13 10 3 13 3 13 2
5 15 3 13 9 2
10 10 3 0 9 15 0 7 0 13 2
25 3 10 9 13 2 3 10 0 9 13 1 0 9 15 9 13 1 15 9 9 2 15 0 13 2
19 1 3 3 0 9 13 15 9 0 2 3 3 10 13 3 9 13 15 2
15 10 3 9 15 15 13 3 3 3 2 10 9 13 3 2
11 9 3 13 7 15 0 0 3 9 9 2
5 9 3 13 15 2
7 9 10 0 15 9 13 2
9 13 3 9 2 13 3 0 9 2
9 10 9 15 3 13 3 3 13 2
5 0 9 7 13 2
7 7 15 3 9 13 15 2
16 9 3 3 0 3 1 9 15 13 0 3 1 10 9 9 2
8 13 15 0 7 3 13 13 2
8 13 0 2 3 1 0 9 2
17 13 13 3 2 3 13 9 15 15 13 2 16 15 9 13 15 2
4 15 3 13 2
6 1 15 0 9 13 2
4 3 13 13 2
9 13 3 13 0 2 7 3 13 2
11 15 1 9 3 3 13 2 13 3 13 2
8 3 3 9 15 15 13 9 2
8 10 9 13 15 15 0 13 2
2 13 2
6 13 3 13 15 9 2
9 7 1 15 13 7 13 3 0 2
9 0 3 3 2 16 13 2 13 2
10 9 15 2 16 13 2 1 9 13 2
12 3 3 15 2 7 13 2 16 13 2 3 2
9 0 3 3 15 2 13 3 9 2
8 13 2 16 15 0 13 3 2
7 10 9 3 15 13 9 2
7 0 3 3 3 9 13 2
12 10 3 1 3 3 13 0 9 15 16 13 2
6 3 3 13 15 15 2
7 13 15 10 13 13 9 2
8 3 3 13 10 9 15 15 2
7 15 3 9 1 0 13 2
12 16 3 0 13 15 13 0 2 13 0 13 2
6 10 0 3 13 0 2
17 15 3 2 15 9 0 10 9 13 16 15 0 13 7 13 13 2
17 1 15 7 9 13 0 7 10 0 13 2 10 0 1 9 13 2
17 13 15 0 10 0 13 9 2 13 3 0 9 3 13 7 13 2
8 13 3 3 9 13 1 9 2
14 10 3 0 13 2 13 3 1 15 7 13 0 9 2
31 13 3 3 3 3 9 3 3 9 3 13 9 15 10 9 2 0 13 2 10 3 3 1 10 9 13 0 0 3 0 2
9 10 3 9 3 13 15 13 0 2
13 13 3 3 3 15 1 13 10 7 3 0 13 2
6 1 3 0 15 13 2
15 10 3 0 10 9 13 3 7 13 2 13 0 9 9 2
8 10 3 13 10 3 0 13 2
6 10 3 9 3 1 2
16 7 3 2 0 3 1 15 9 1 2 13 10 0 0 9 2
36 9 3 2 16 13 2 13 1 13 10 3 9 3 0 2 9 0 9 13 2 1 15 13 3 0 2 15 3 13 13 10 0 0 0 9 2
8 7 3 1 15 3 13 13 2
20 13 3 13 9 2 1 15 3 13 10 0 13 0 2 7 1 0 13 13 2
23 13 3 15 9 13 13 2 9 3 3 9 2 0 3 3 13 0 9 15 3 7 9 2
7 13 3 0 9 13 15 2
11 3 3 0 10 9 13 2 0 9 13 2
10 0 13 3 3 3 3 13 13 9 2
22 0 3 3 9 9 13 2 3 3 13 9 13 9 2 7 3 0 9 9 13 13 2
16 15 1 12 13 2 3 0 1 2 7 9 7 9 0 0 2
11 10 3 0 3 9 13 3 3 9 3 2
10 3 3 13 10 0 1 15 9 0 2
8 9 3 3 7 9 15 13 2
5 13 3 7 15 2
6 9 3 9 15 13 2
10 9 3 13 3 0 0 7 13 13 2
18 7 3 3 13 13 15 2 13 0 13 2 0 13 2 0 3 13 2
5 0 9 13 15 2
6 15 15 9 13 3 2
12 0 13 15 3 9 3 15 9 7 9 0 2
8 3 3 13 15 10 0 13 2
18 3 3 15 13 2 7 13 3 2 3 0 2 10 3 0 9 7 2
11 6 0 13 2 3 13 0 0 9 13 2
5 15 15 13 9 2
14 15 3 13 15 13 2 15 3 13 9 13 13 0 2
7 13 15 7 7 15 13 2
22 13 15 13 2 15 0 9 0 0 13 15 1 3 9 13 13 2 0 1 9 13 2
13 3 3 3 13 3 13 0 3 3 15 15 9 2
6 13 15 0 3 13 2
15 3 9 3 3 9 13 3 3 9 9 13 15 13 1 2
12 16 3 15 0 3 0 0 2 0 13 9 2
8 3 13 16 15 13 13 3 2
9 0 3 13 3 13 16 13 0 2
18 16 3 15 3 3 13 0 13 2 7 15 13 2 3 3 13 3 2
29 15 3 3 13 9 0 13 9 3 3 13 1 9 13 3 3 3 0 9 2 15 15 12 9 13 0 9 13 2
15 7 10 9 3 9 13 0 2 13 16 13 2 13 15 2
11 15 15 9 13 0 0 13 9 0 13 2
29 7 16 10 13 3 13 9 1 9 9 2 3 3 13 15 7 13 0 0 9 2 16 13 0 3 7 13 9 2
9 3 3 0 3 13 1 0 13 2
7 13 2 13 9 0 13 2
5 13 2 7 13 2
22 7 15 13 1 9 13 15 9 10 13 7 10 13 2 16 9 13 0 1 15 9 2
6 15 15 13 9 0 2
9 10 3 3 1 0 0 13 0 2
34 7 16 10 0 7 13 3 9 2 10 3 0 13 9 13 9 9 2 15 9 0 3 13 2 15 3 9 3 9 0 3 9 13 2
7 7 3 0 1 9 13 2
14 15 1 9 3 0 3 13 0 3 13 3 13 0 2
19 1 9 2 16 9 15 13 2 0 13 1 0 9 15 2 13 15 15 2
8 1 15 3 3 3 15 13 2
8 7 15 15 9 3 13 13 2
14 13 15 9 1 15 0 0 2 3 0 13 15 0 2
4 3 13 0 2
7 3 3 9 0 13 1 2
10 7 3 15 3 1 10 9 9 13 2
18 7 15 3 13 3 7 13 2 15 3 1 9 0 15 13 9 13 2
9 7 3 3 10 3 0 13 1 2
44 15 3 3 13 15 0 9 13 9 13 2 7 13 15 13 9 2 3 13 0 9 0 2 15 9 3 15 9 3 13 13 0 9 2 16 1 0 2 15 15 13 2 13 2
11 7 10 3 15 9 2 3 13 2 13 2
16 9 13 2 16 7 9 3 13 2 3 3 13 2 10 9 2
4 15 15 13 2
10 7 3 3 9 13 15 13 13 0 2
3 15 13 2
22 3 3 13 3 1 9 10 15 0 13 2 7 15 13 9 13 15 10 0 0 0 2
3 13 15 2
2 13 2
17 15 3 13 10 13 15 2 13 10 13 9 2 15 15 13 3 2
25 3 13 2 13 1 10 9 15 10 0 9 2 15 10 0 9 15 3 13 10 3 0 13 9 2
4 7 15 13 2
5 13 3 3 13 2
21 0 3 9 13 1 9 2 0 3 9 2 3 3 13 1 9 13 1 10 9 2
5 15 3 0 13 2
6 10 9 9 15 13 2
19 10 13 13 2 3 3 0 13 2 1 10 0 13 15 2 15 0 13 2
3 0 13 2
4 3 15 13 2
16 7 13 15 2 3 0 13 0 0 2 1 0 10 0 9 2
4 0 3 13 2
5 7 13 9 1 2
6 13 1 15 3 13 2
7 13 2 7 3 13 13 2
6 10 9 15 13 9 2
6 7 9 3 0 13 2
4 3 13 3 2
4 13 15 3 2
9 0 7 13 3 3 13 13 3 2
6 13 3 15 3 3 2
7 13 3 2 9 3 13 2
6 3 0 3 13 15 2
5 0 7 13 13 2
9 7 3 13 3 15 10 9 13 2
39 3 3 13 2 13 9 10 0 13 0 3 9 0 15 2 3 15 9 1 9 15 3 1 0 0 7 9 13 13 13 13 15 1 9 2 9 0 9 2
10 16 3 15 9 13 9 2 13 9 2
32 3 3 9 0 2 16 13 9 2 1 10 0 9 3 13 2 7 0 9 13 2 3 3 15 15 3 13 0 1 0 13 2
28 15 3 3 13 10 0 9 2 16 13 15 9 9 9 13 10 13 1 2 13 15 0 10 9 15 13 3 2
17 3 3 15 7 9 3 7 9 0 13 2 3 3 13 3 13 2
7 15 3 0 0 13 9 2
18 13 3 9 13 16 13 9 1 0 9 2 9 0 1 0 9 13 2
5 3 10 9 13 2
49 15 3 9 9 2 16 13 2 9 0 7 0 9 13 3 0 13 3 2 9 0 13 9 2 15 7 15 9 13 3 13 2 16 9 13 0 9 13 0 2 0 16 13 9 0 3 7 13 2
14 15 3 15 13 0 2 16 9 13 9 13 13 9 2
9 13 3 2 0 9 1 9 0 2
11 3 3 13 3 7 10 0 9 3 13 2
9 15 3 13 9 9 1 9 13 2
5 13 3 3 0 2
4 15 3 13 2
6 3 13 10 0 9 2
6 13 13 3 13 9 2
12 0 3 13 9 3 1 15 7 9 15 13 2
9 0 3 13 3 13 9 0 9 2
12 6 10 15 13 13 2 16 15 9 15 13 2
18 7 1 10 0 1 0 9 3 13 13 2 1 15 9 13 0 0 2
6 15 15 10 0 13 2
23 15 3 15 0 13 2 0 2 0 2 0 3 13 2 9 0 2 10 0 9 13 0 2
10 15 3 13 15 3 13 15 3 13 2
8 15 3 3 15 13 9 13 2
11 3 3 3 13 2 13 3 3 13 13 2
12 0 10 0 9 13 3 15 13 13 3 13 2
15 7 15 3 10 0 13 3 9 0 2 3 3 3 13 2
31 15 1 9 13 2 15 0 0 9 13 2 7 3 15 0 0 13 9 9 2 3 3 0 1 9 2 0 3 13 9 2
24 9 13 10 13 2 9 10 13 2 0 3 13 9 2 16 3 9 3 9 13 10 0 13 2
19 15 9 10 0 0 0 9 13 13 2 3 3 3 9 13 15 13 9 2
5 13 7 3 13 2
14 3 9 13 1 0 10 13 0 1 9 13 3 3 2
13 0 3 15 0 13 2 0 0 13 3 9 9 2
5 0 13 2 0 2
7 13 2 3 13 15 9 2
14 7 1 3 0 3 13 0 9 2 16 15 9 13 2
15 15 3 0 13 2 3 3 3 1 9 13 0 3 9 2
17 7 3 9 3 13 2 9 3 15 0 2 7 13 15 9 9 2
6 7 15 9 9 13 2
6 1 15 0 13 9 2
21 3 13 0 0 3 2 16 15 13 0 2 13 0 2 9 0 13 9 0 9 2
30 16 3 10 3 13 9 3 7 0 13 13 0 2 15 3 7 3 13 0 9 2 13 3 3 9 0 3 9 0 2
9 16 3 7 3 13 2 15 13 2
5 15 3 13 3 2
11 7 10 9 3 0 13 15 13 2 13 2
15 3 3 15 0 9 2 0 13 9 2 3 13 15 3 2
13 15 1 9 7 1 9 3 13 3 16 13 13 2
13 15 0 3 15 9 2 10 15 13 2 0 13 2
25 3 9 1 10 15 10 9 10 9 13 2 1 15 13 1 15 15 13 3 3 7 10 13 13 2
31 7 3 13 10 13 2 13 0 9 2 1 15 3 9 10 0 1 9 13 2 0 9 13 7 13 9 0 0 15 0 2
21 15 3 13 10 0 1 9 13 2 13 2 13 9 10 0 9 13 0 1 0 2
12 3 3 3 13 1 15 0 15 9 9 13 2
11 0 3 10 9 0 9 13 15 13 0 2
16 3 13 2 3 3 15 1 9 3 10 3 13 10 3 9 2
3 15 13 2
6 3 3 0 13 13 2
15 3 0 15 13 9 2 15 1 9 13 9 10 0 13 2
8 7 13 3 13 3 0 9 2
12 15 3 9 15 13 3 9 13 10 0 13 2
15 13 3 3 13 15 10 13 3 15 7 10 13 9 13 2
15 13 13 2 0 13 9 3 13 15 15 7 13 1 9 2
12 7 13 15 3 2 16 13 3 2 0 13 2
5 3 3 9 13 2
16 3 3 15 13 3 1 9 10 0 13 2 16 3 0 13 2
5 7 3 13 13 2
5 7 3 15 13 2
9 10 9 15 13 2 13 7 13 2
3 13 13 2
3 13 3 2
7 13 3 0 15 13 13 2
8 13 3 13 9 9 13 0 2
8 7 3 15 13 0 3 9 2
2 13 2
7 13 0 2 16 13 0 2
9 13 2 16 3 3 3 13 15 2
6 7 3 3 13 9 2
20 3 3 1 0 15 13 13 13 2 7 7 13 3 13 15 2 13 3 7 2
8 0 3 0 7 15 13 13 2
13 16 3 0 15 13 13 2 10 13 13 0 0 2
13 0 3 15 0 9 0 0 2 0 1 15 13 2
29 15 13 3 3 16 2 16 13 9 2 10 0 9 13 3 2 15 3 9 0 13 3 3 13 10 3 13 13 2
7 3 0 1 0 9 13 2
17 7 13 2 7 13 1 15 2 15 15 9 13 3 15 13 9 2
3 3 13 2
16 13 3 0 2 16 10 13 9 13 2 16 15 13 3 9 2
26 15 3 3 3 3 3 2 3 3 16 15 10 0 13 15 13 9 2 1 15 3 13 2 0 13 2
9 15 3 0 9 13 7 13 9 2
9 15 3 13 15 7 13 0 9 2
17 10 0 3 3 13 9 13 2 3 3 3 15 2 0 3 13 2
13 3 3 13 9 0 0 9 13 2 13 10 9 2
13 3 3 13 0 0 2 13 9 7 0 13 0 2
22 3 3 3 13 3 2 16 7 0 0 1 0 13 13 2 15 0 10 0 13 9 2
6 13 13 3 15 0 2
13 16 3 15 15 0 15 13 2 3 3 13 3 2
8 7 13 15 0 0 13 15 2
30 13 3 15 2 16 15 7 13 9 2 3 13 3 7 3 9 9 13 2 13 3 1 0 9 9 15 1 13 0 2
11 1 0 13 7 15 7 3 0 13 13 2
8 3 0 3 15 7 13 13 2
8 7 13 15 3 7 1 9 2
5 15 3 13 9 2
8 9 3 10 13 3 9 13 2
11 7 13 3 2 16 15 3 3 13 13 2
8 7 15 13 10 0 13 0 2
4 7 3 13 2
5 3 0 9 13 2
8 13 2 16 13 2 9 13 2
7 0 13 9 1 0 13 2
8 15 3 3 13 7 13 15 2
7 7 3 9 15 13 0 2
6 13 3 3 13 9 2
4 3 3 13 2
7 9 15 13 9 13 9 2
3 3 13 2
5 0 3 13 13 2
4 15 0 13 2
8 13 15 9 15 15 9 1 2
10 16 15 13 15 9 2 13 3 3 2
8 7 3 13 1 1 0 13 2
4 13 7 15 2
10 0 3 0 9 13 3 7 13 9 2
16 9 15 0 13 13 9 10 0 3 0 0 9 13 1 9 2
16 0 3 0 3 13 2 1 16 13 15 0 15 10 9 9 2
10 16 3 15 13 2 1 0 13 3 2
19 7 7 9 7 0 9 13 15 2 3 7 3 1 9 9 0 13 9 2
9 7 16 13 0 0 0 13 3 2
24 9 3 3 2 16 7 0 9 0 13 2 15 0 9 3 3 3 15 3 13 2 15 13 2
30 13 3 16 15 3 0 13 9 15 1 9 13 9 2 1 15 13 0 2 16 0 2 13 2 1 9 9 9 13 2
10 3 7 13 0 0 0 10 9 13 2
3 3 13 2
5 7 0 3 13 2
35 13 3 13 3 0 15 0 0 1 0 13 2 7 9 9 1 0 9 0 3 13 13 9 2 16 10 0 0 0 9 13 16 3 13 2
14 13 3 3 2 13 15 0 13 13 15 0 0 9 2
6 1 9 10 9 13 2
2 13 2
14 10 3 0 3 13 9 12 13 2 7 13 10 13 2
9 13 15 9 2 0 13 3 9 2
26 3 3 3 13 3 10 13 15 9 9 2 3 3 10 0 0 0 9 2 15 15 13 0 1 9 2
12 13 7 9 7 9 10 0 13 9 9 9 2
11 0 0 3 13 0 9 9 15 3 9 2
18 1 15 3 15 13 7 3 7 3 15 0 13 9 10 13 7 13 2
22 7 3 9 9 3 13 1 0 9 3 3 1 0 2 16 7 15 9 9 3 13 2
24 16 3 10 13 9 13 2 0 9 0 9 0 13 2 3 15 3 13 1 15 9 0 9 2
9 13 3 2 3 13 2 3 13 2
17 3 3 13 9 2 15 15 13 3 7 3 0 3 13 13 0 2
11 3 3 16 13 0 2 0 13 15 3 2
21 3 0 1 0 15 3 13 16 0 7 3 9 13 2 13 7 15 7 10 0 2
17 15 3 9 3 3 13 2 3 3 15 13 3 13 1 15 3 2
3 3 13 2
6 15 9 3 13 15 2
19 10 3 9 15 13 2 3 15 0 2 15 13 15 13 2 16 13 13 2
4 0 0 13 2
9 7 3 13 0 10 3 0 13 2
15 7 1 9 3 9 13 0 2 3 13 15 15 13 9 2
26 0 0 9 3 13 0 2 15 15 3 13 13 13 2 9 7 9 13 2 15 10 9 15 13 9 2
10 13 3 2 16 7 0 3 9 13 2
11 13 3 3 10 13 3 2 16 9 13 2
9 15 3 3 3 13 10 13 0 2
14 16 3 15 13 13 3 2 9 0 13 10 3 13 2
16 13 3 3 3 3 15 16 13 15 0 3 15 15 13 1 2
17 7 16 13 15 2 10 13 3 1 13 3 3 10 9 3 3 2
4 7 3 13 2
14 16 3 15 3 3 9 13 2 3 3 13 0 13 2
5 7 3 13 15 2
4 9 13 13 2
15 15 3 0 9 13 3 0 3 2 16 3 3 3 7 2
15 13 3 10 9 9 2 15 9 15 0 9 13 1 9 2
27 9 3 0 2 3 15 13 2 9 13 1 9 13 9 0 9 9 2 15 1 9 13 9 15 13 13 2
18 1 15 13 0 9 13 0 2 16 9 0 10 9 13 10 0 9 2
6 3 13 10 0 9 2
15 1 15 2 13 0 13 2 3 13 0 2 3 9 9 2
13 13 13 15 10 9 9 7 9 15 7 9 13 2
18 16 3 13 0 1 0 2 15 3 0 13 3 2 16 9 3 13 2
8 7 13 7 9 3 13 13 2
5 3 0 13 3 2
10 7 7 0 13 16 10 9 9 13 2
18 7 3 3 3 3 13 13 15 2 10 0 13 9 16 10 9 13 2
28 7 15 15 9 16 9 3 0 1 15 13 2 10 13 9 0 2 1 3 15 0 0 3 13 10 3 0 2
9 15 0 3 15 15 13 9 13 2
17 15 3 7 13 15 1 0 2 3 13 0 3 0 7 9 0 2
16 16 3 13 15 10 9 0 2 3 15 10 0 3 13 9 2
4 13 9 13 2
19 0 3 15 13 1 3 15 9 2 15 0 10 13 13 2 7 0 0 2
11 3 15 13 13 3 1 0 9 9 1 2
13 3 3 13 15 15 9 13 2 16 7 13 15 2
9 13 3 16 0 13 3 15 13 2
16 7 10 3 1 15 9 7 10 0 9 13 15 0 13 9 2
6 0 3 0 9 13 2
8 15 3 13 15 2 3 15 2
5 15 3 13 9 2
7 15 3 9 10 9 13 2
2 13 2
15 1 9 13 2 13 15 13 15 13 2 3 3 13 13 2
17 3 13 3 3 1 0 9 13 15 2 16 15 3 13 0 13 2
6 13 2 13 2 13 2
13 3 3 13 0 9 2 16 3 3 3 13 3 2
33 3 3 1 0 10 9 2 3 3 0 13 13 1 9 13 15 0 15 2 16 1 9 3 7 0 9 13 0 9 1 0 9 2
4 7 3 13 2
5 3 3 15 13 2
13 10 3 0 0 7 13 15 13 15 9 13 13 2
9 15 1 9 3 13 13 0 13 2
4 0 13 3 2
8 3 7 9 15 13 13 0 2
6 13 3 3 9 13 2
5 15 15 0 1 2
12 15 13 13 9 0 0 1 9 9 3 3 2
4 13 15 13 2
10 13 3 15 0 13 15 15 13 9 2
2 13 2
3 13 9 2
5 1 0 13 13 2
4 7 0 13 2
8 13 9 3 3 7 3 13 2
8 13 1 0 7 15 0 13 2
33 0 3 13 1 10 0 9 9 9 0 9 9 2 16 13 9 0 9 9 13 2 15 0 9 2 13 0 2 0 15 3 9 2
13 9 3 13 10 9 10 9 9 13 13 0 9 2
15 16 3 1 0 0 15 13 3 13 15 9 9 7 9 2
4 9 3 13 2
14 16 3 15 9 13 2 13 3 3 3 3 13 13 2
18 0 3 0 9 2 16 0 13 9 13 9 9 2 13 0 9 1 2
14 9 13 0 2 9 1 9 2 12 9 0 9 9 2
18 13 3 16 0 10 13 9 9 13 7 13 9 2 0 1 9 13 2
9 15 3 3 9 13 9 9 13 2
9 3 3 0 13 9 9 0 9 2
5 9 3 3 13 2
17 3 3 0 13 13 9 0 2 16 13 9 15 0 7 9 0 2
13 3 3 1 9 7 9 9 13 2 13 0 9 2
8 7 3 3 0 0 13 9 2
9 3 3 0 9 0 9 9 13 2
14 1 3 9 13 0 0 3 3 9 9 13 0 9 2
17 3 0 0 1 9 0 13 13 2 0 3 13 9 0 0 9 2
15 13 3 0 3 2 0 13 9 9 2 10 9 9 13 2
30 16 3 13 0 15 13 2 0 1 9 9 13 0 9 13 2 13 9 13 2 3 0 2 3 0 9 13 0 9 2
15 7 10 3 0 0 0 9 13 10 0 0 1 0 9 2
11 3 13 9 0 13 9 13 9 0 13 2
9 13 3 9 0 9 1 9 13 2
6 1 3 13 0 9 2
10 15 3 13 9 9 13 1 0 9 2
23 7 15 9 13 3 1 0 9 0 9 0 9 13 9 9 13 2 16 0 9 13 9 2
14 10 0 3 9 10 3 0 2 3 13 2 13 9 2
12 3 3 13 2 16 10 15 10 9 13 0 2
5 0 10 13 13 2
9 3 3 3 13 9 15 13 13 2
23 16 3 3 9 9 3 3 1 9 15 13 0 2 7 10 13 9 13 15 3 3 13 2
4 15 13 3 2
7 0 3 3 13 3 13 2
6 13 15 13 13 3 2
2 13 2
5 3 3 13 13 2
7 3 9 7 15 13 15 2
8 13 15 2 3 16 15 13 2
9 3 13 3 2 16 15 3 13 2
4 7 13 3 2
14 15 3 3 13 13 15 3 0 7 10 10 0 0 2
22 13 3 10 0 13 9 15 15 0 13 9 3 2 15 9 13 13 0 3 15 0 2
7 3 3 3 15 13 13 2
10 0 3 13 2 15 3 13 7 9 2
5 3 15 3 13 2
12 1 0 13 15 2 16 13 2 10 3 13 2
4 9 0 13 2
2 13 2
15 16 10 3 13 1 9 9 13 2 1 15 13 3 13 2
9 13 3 9 9 0 9 13 9 2
3 0 13 2
2 13 2
3 13 13 2
6 15 3 0 3 13 2
4 0 0 13 2
3 13 13 2
8 7 15 3 3 13 2 16 3
3 15 13 2
5 0 0 13 9 2
13 13 2 3 3 15 9 13 3 3 9 1 15 2
11 13 3 9 3 9 15 3 13 7 13 0
16 3 3 3 13 10 0 15 9 9 2 15 9 3 13 13 2
10 7 15 9 9 15 13 3 13 3 2
16 15 3 1 15 3 3 0 2 0 9 13 2 15 13 9 2
9 1 15 15 13 13 15 0 9 2
16 1 3 9 13 2 16 13 15 10 0 7 13 7 0 13 2
8 7 3 13 15 0 0 13 2
24 16 3 13 9 0 9 2 13 9 1 0 0 9 9 7 0 9 0 0 13 9 9 9 2
8 0 3 13 9 0 9 13 2
15 7 3 3 3 7 3 13 7 15 15 9 1 0 13 2
10 15 3 13 1 3 15 7 15 15 2
11 15 3 3 1 9 13 0 15 13 9 2
18 7 3 3 3 3 9 3 10 9 13 0 13 3 3 13 13 3 2
6 7 13 9 0 0 2
9 10 0 3 3 0 3 9 13 2
6 15 13 10 3 0 2
10 10 3 3 3 0 13 9 9 0 2
4 15 3 13 2
6 3 1 9 13 15 2
10 3 13 3 9 3 3 3 9 13 2
10 3 3 3 15 13 15 3 13 3 2
6 9 1 0 3 13 2
5 15 15 13 9 2
12 15 3 9 3 13 15 0 9 1 9 9 2
16 15 3 1 9 9 15 13 13 2 3 13 3 7 13 9 2
15 7 3 2 16 13 2 10 3 13 3 0 3 13 0 2
5 3 13 15 0 2
12 16 3 15 13 2 10 3 13 9 13 9 2
6 3 10 13 13 3 2
6 3 13 15 3 13 2
6 3 3 3 0 13 2
7 15 3 13 15 15 0 2
9 7 16 15 9 3 2 3 13 2
8 13 2 9 3 1 0 13 2
2 13 2
6 13 0 0 3 13 2
7 13 3 3 3 13 13 2
20 9 3 13 7 15 3 0 16 0 15 13 2 7 9 13 13 7 0 13 2
20 15 3 16 3 10 9 9 13 3 13 2 13 9 9 3 0 9 13 9 2
8 0 3 15 13 13 15 3 2
12 3 3 13 0 2 1 15 9 13 3 0 2
21 15 13 3 13 9 0 9 13 2 13 3 13 1 15 10 9 0 13 0 3 2
9 7 15 3 3 13 16 13 3 2
20 3 3 3 0 13 9 9 16 0 3 7 0 9 13 13 2 9 0 0 2
20 3 16 13 10 0 9 2 0 3 9 1 9 3 13 13 10 9 3 3 2
15 3 3 2 3 13 2 0 13 10 0 7 9 0 13 2
8 13 3 1 10 0 0 13 2
13 15 3 3 9 7 0 15 13 15 9 3 13 2
23 0 13 13 2 15 13 0 13 2 15 1 3 9 1 3 0 9 13 0 7 9 9 2
13 1 10 0 13 10 9 7 10 13 7 13 0 2
13 3 3 3 13 0 9 0 3 13 15 13 13 2
3 3 13 2
14 9 3 3 3 9 13 2 13 3 0 10 0 9 2
15 9 3 15 3 13 1 9 2 15 3 13 1 9 13 2
10 15 3 0 9 13 13 0 9 13 2
13 13 3 15 0 3 3 13 9 0 13 3 13 2
16 7 13 2 16 0 10 0 15 3 13 13 9 2 13 9 2
2 13 2
12 9 0 9 13 9 13 0 3 3 9 0 2
4 0 0 13 2
7 3 3 13 15 13 13 2
7 3 3 3 0 3 13 2
9 6 13 15 10 9 9 13 13 2
5 0 3 3 13 2
11 7 13 9 3 2 10 3 9 0 3 2
7 13 0 9 1 9 13 2
6 3 3 13 13 15 2
10 13 15 10 9 2 10 3 9 13 2
6 13 13 16 3 13 2
10 7 3 3 1 15 3 7 13 15 2
2 13 2
6 15 3 9 3 1 2
2 13 2
6 7 15 9 3 1 2
7 13 9 0 0 13 0 2
9 3 3 3 0 9 13 15 15 2
9 7 3 13 3 3 15 9 13 2
8 10 0 0 3 13 15 13 2
10 16 3 3 13 2 3 13 15 15 2
7 13 3 15 15 13 0 2
8 3 13 15 0 1 9 13 2
8 7 13 3 10 9 9 13 2
8 0 15 13 10 9 3 13 2
8 7 16 13 0 2 13 15 2
8 7 3 13 3 0 13 15 2
9 7 0 0 2 3 3 13 3 2
7 9 3 0 13 0 0 2
7 13 13 0 15 15 13 2
7 3 13 0 3 3 15 2
3 13 3 2
3 7 13 2
13 3 15 7 13 3 2 3 3 16 3 13 13 2
11 7 16 15 13 13 15 13 2 13 0 2
11 16 3 1 0 3 13 2 0 13 9 2
33 0 3 0 13 9 2 15 3 9 0 13 2 16 10 0 9 2 3 3 15 10 13 0 10 3 7 13 0 2 0 13 9 2
6 15 3 9 3 13 2
13 13 15 3 9 7 9 0 0 0 3 9 13 2
8 15 3 13 7 15 13 13 2
8 7 3 3 13 10 13 0 2
13 15 3 3 0 15 1 13 3 15 0 9 9 2
6 3 13 10 0 9 2
9 7 15 9 13 9 9 13 1 2
5 3 15 13 9 2
14 13 0 0 9 1 0 9 13 2 3 13 2 13 2
14 16 15 13 10 0 0 2 15 9 13 9 0 13 2
7 13 2 15 13 2 13 2
19 3 3 3 1 9 3 13 13 15 2 7 7 0 15 7 1 9 9 2
31 3 13 3 13 9 2 16 1 0 15 9 13 9 13 15 13 9 2 16 13 13 10 3 9 2 9 0 0 13 9 2
11 3 3 13 0 1 9 0 13 1 15 2
7 0 3 13 9 16 13 2
3 13 9 2
4 13 15 15 2
5 0 0 13 13 2
4 13 3 0 2
19 13 3 1 9 9 9 2 15 15 15 3 9 3 13 3 13 0 0 2
25 7 0 10 0 9 10 0 3 0 13 2 15 15 3 15 13 1 0 9 9 3 7 9 0 2
22 7 3 3 13 3 2 1 15 13 10 0 2 7 3 13 10 0 13 7 13 9 2
7 10 3 13 3 13 13 2
5 16 7 3 13 2
7 0 3 15 0 13 13 2
3 15 13 2
5 3 9 13 13 2
6 13 3 3 9 13 2
5 15 3 13 9 2
6 1 15 0 13 13 2
9 15 13 0 2 7 3 3 13 2
7 1 15 13 15 10 13 2
9 7 3 13 3 0 10 0 0 2
9 7 3 13 3 15 3 0 13 2
5 3 0 13 0 2
5 3 15 13 9 2
8 15 3 15 9 15 13 9 2
8 9 13 2 9 3 0 13 2
9 3 3 13 3 3 10 13 1 2
8 15 13 3 15 15 13 9 2
7 0 9 3 13 13 3 2
8 0 3 13 10 0 13 0 2
8 3 3 3 15 0 13 3 2
10 15 13 3 2 16 15 15 0 1 2
9 7 13 0 2 16 1 0 13 2
10 13 15 9 3 2 16 10 0 13 2
6 13 13 3 13 3 2
4 3 13 13 2
3 0 13 2
6 1 9 3 3 13 2
8 3 10 13 9 3 9 13 2
7 3 15 13 15 13 9 2
6 3 0 13 10 13 2
8 3 3 13 0 15 0 9 2
3 3 13 2
7 15 3 13 3 13 9 2
5 3 13 3 9 2
10 15 13 15 9 9 13 16 0 13 2
4 3 3 13 2
4 13 15 9 2
2 13 2
5 7 3 13 13 2
4 15 3 13 2
10 13 3 3 3 1 9 16 9 13 2
6 3 3 13 13 3 2
14 10 0 15 2 10 0 3 13 13 13 15 9 9 2
7 3 3 13 3 0 9 2
3 13 15 2
4 3 13 15 2
13 15 3 3 0 3 15 13 13 3 3 9 9 2
8 3 13 2 16 9 15 13 13
15 13 0 15 3 3 9 2 16 15 9 13 0 1 9 2
5 0 0 13 15 2
14 10 3 15 13 13 13 2 10 3 13 3 9 13 2
4 15 7 13 2
9 7 15 13 10 0 9 9 13 2
7 3 3 7 0 13 13 2
2 13 2
5 3 3 13 15 2
15 13 3 0 13 9 2 15 15 3 3 3 1 0 13 2
32 10 3 13 10 9 13 2 7 3 9 3 0 13 15 2 3 3 0 9 9 9 13 2 15 3 13 2 10 3 13 3 2
8 9 3 3 15 9 13 9 2
9 7 3 1 9 10 3 13 13 2
11 16 3 13 2 3 13 13 7 13 3 2
9 3 3 3 3 13 10 13 9 2
9 7 13 3 3 2 3 3 3 2
17 3 3 3 13 15 2 15 0 15 15 9 13 3 7 13 13 2
5 13 3 15 0 2
13 16 3 0 15 13 9 2 13 0 3 15 9 2
10 7 3 3 3 13 15 7 3 13 2
10 13 13 16 1 9 13 15 3 13 2
7 3 3 9 15 13 15 2
30 7 3 13 10 0 9 7 10 0 15 1 9 9 1 13 2 16 10 3 13 0 1 10 0 13 2 13 3 9 2
7 3 3 13 3 13 15 2
7 13 3 15 7 13 15 2
8 13 2 16 13 2 3 13 2
9 9 15 1 9 13 3 13 9 2
4 13 3 0 2
4 13 13 3 2
3 3 13 2
7 3 3 3 1 9 13 2
9 3 13 15 15 13 1 9 3 2
3 15 13 2
3 15 13 2
6 7 15 13 0 9 2
13 3 15 0 13 2 15 15 15 13 1 0 9 2
5 9 3 13 13 2
2 13 2
13 13 3 16 3 15 9 15 13 13 1 9 0 2
4 13 13 15 2
11 15 3 13 3 10 13 16 3 9 13 2
15 16 3 13 2 13 3 0 3 7 0 0 0 0 13 2
9 13 3 13 10 0 9 13 9 2
20 13 3 9 0 0 0 9 0 9 2 16 3 3 3 13 0 9 9 13 2
18 13 3 9 9 0 1 9 2 0 9 1 9 2 0 9 9 13 2
16 10 9 3 9 9 15 13 9 9 13 1 0 9 3 13 2
4 7 3 13 2
4 15 3 13 2
12 15 3 1 9 9 13 2 15 3 13 3 2
7 15 3 3 13 1 15 2
4 13 15 3 2
12 7 3 1 15 13 0 3 3 10 13 9 2
7 13 2 16 13 2 0 2
3 13 9 2
6 13 10 9 1 13 2
10 0 3 9 13 10 13 10 3 13 2
5 7 3 13 15 2
12 0 3 9 13 9 9 2 3 3 13 13 2
4 13 10 0 2
9 3 13 0 16 15 9 13 3 2
2 13 2
6 13 3 9 1 0 2
5 13 3 10 9 2
2 13 2
2 13 2
5 3 13 13 3 2
4 7 3 13 2
5 3 3 13 15 2
20 1 9 3 0 3 3 3 13 1 9 15 13 2 0 16 13 1 9 9 2
20 15 13 15 3 3 10 9 0 2 15 13 9 15 13 9 13 0 1 9 2
2 13 2
10 9 3 3 3 13 10 0 10 0 2
7 15 3 3 13 10 0 2
3 13 15 2
5 0 3 9 13 2
7 3 7 13 13 7 3 2
9 3 2 7 13 2 3 9 0 2
7 13 3 15 16 0 13 2
8 13 3 2 7 3 0 9 2
8 3 0 13 15 13 3 3 2
9 13 3 2 16 15 0 13 15 2
37 13 13 13 9 0 0 0 3 13 2 16 16 15 0 9 0 3 13 9 15 2 3 13 9 9 13 0 3 3 1 9 15 9 13 13 9 2
6 7 3 13 1 15 2
11 10 3 9 9 13 2 16 13 10 0 2
8 16 3 13 9 2 3 13 2
15 13 0 9 1 9 2 16 10 0 3 1 15 9 13 2
5 7 3 13 13 2
4 3 3 13 2
3 15 13 2
3 15 13 2
11 3 3 13 3 13 10 13 16 13 0 2
12 3 3 13 16 15 3 9 13 10 13 15 2
7 7 9 13 0 13 3 2
7 7 15 13 7 0 13 2
15 15 3 9 3 1 0 13 13 10 13 3 9 9 13 2
18 7 3 0 13 7 13 13 9 2 15 15 13 13 13 2 0 15 2
6 13 3 3 1 9 2
12 9 3 3 3 13 9 2 7 0 9 1 2
7 15 3 1 9 13 15 2
14 3 2 15 16 0 9 2 9 13 3 0 13 13 2
3 7 13 2
14 13 3 3 13 9 10 0 2 16 3 1 0 13 2
7 15 15 9 13 15 0 2
7 7 3 0 10 9 13 2
8 0 13 2 10 3 9 13 2
3 7 13 2
2 13 2
7 13 13 15 0 15 0 2
8 10 3 0 3 3 13 0 2
29 0 3 9 13 9 7 9 13 2 0 3 10 3 1 9 13 9 15 1 9 2 13 15 3 9 7 9 9 2
9 7 3 3 9 13 2 13 3 2
15 0 3 0 9 13 2 0 2 15 1 9 9 9 13 2
7 3 10 10 13 0 9 2
19 3 0 3 0 2 0 13 0 9 2 3 13 2 9 3 13 7 9 2
21 10 3 0 9 13 7 9 9 9 13 9 0 9 1 9 0 2 13 9 13 2
27 7 16 3 9 13 13 9 2 10 10 13 9 3 13 1 9 2 3 3 13 13 9 3 1 15 0 2
7 9 3 13 0 1 9 2
11 10 3 3 13 0 9 16 15 9 13 2
11 10 3 3 0 9 1 9 0 0 13 2
10 10 3 9 13 9 9 3 9 3 2
8 10 10 3 13 9 0 13 2
11 2 6 6 2 0 3 3 9 9 13 2
16 1 3 9 9 13 9 2 3 3 13 3 7 15 13 9 2
12 3 13 9 2 7 3 9 9 13 0 13 2
7 3 3 0 0 13 2 2
18 10 9 0 13 13 2 3 3 0 7 0 9 13 2 16 9 13 2
14 3 9 2 13 3 9 13 13 15 9 2 13 13 2
14 3 3 15 9 0 1 9 13 0 13 9 1 0 2
8 15 3 13 13 9 9 2 2
27 3 3 3 9 15 0 13 2 15 1 3 9 13 9 2 1 3 0 9 0 13 2 10 9 0 13 2
6 9 3 13 15 9 2
14 3 3 3 3 13 1 0 0 3 9 13 0 2 2
39 3 15 3 13 2 16 15 9 3 13 7 15 9 1 9 13 2 1 9 13 9 13 0 0 9 13 2 15 3 15 3 9 0 13 7 9 9 9 2
25 3 13 1 9 13 0 9 2 0 0 2 15 15 13 7 1 0 7 1 0 9 1 9 9 2
24 13 3 0 9 2 0 0 9 2 0 0 0 2 10 13 9 9 9 2 10 3 13 9 2
20 13 3 1 9 9 13 2 13 3 9 1 9 1 9 9 2 9 1 0 2
6 13 3 3 9 9 2
17 15 3 3 9 1 9 9 13 13 1 9 9 2 15 13 0 2
42 15 3 0 0 13 9 0 2 13 3 1 9 0 13 9 2 13 9 0 1 9 2 16 3 13 9 10 3 9 1 9 13 2 9 3 0 13 7 9 15 13 2
14 13 3 0 9 2 13 3 1 9 9 3 9 13 2
18 3 3 13 9 13 0 7 13 0 9 2 7 15 13 9 0 13 2
10 3 3 9 13 13 15 15 13 2 2
6 1 3 9 9 13 2
29 1 3 0 9 13 0 2 1 0 9 2 16 9 13 9 9 13 2 0 13 2 7 16 15 1 9 13 13 2
15 9 3 0 9 13 13 0 0 2 1 0 9 2 13 2
6 1 3 0 13 9 2
14 9 3 0 9 13 13 2 9 0 13 2 13 13 2
15 9 3 9 9 13 13 0 2 1 3 15 13 0 9 2
7 9 3 0 3 13 13 2
6 1 3 13 9 0 2
33 10 3 3 3 13 1 9 3 9 3 2 15 3 9 3 9 1 9 13 2 9 3 9 13 1 9 2 9 3 9 13 0 2
9 15 3 1 9 0 13 9 13 2
16 9 3 1 9 9 0 13 9 2 15 3 13 1 9 9 2
8 3 3 15 13 13 0 13 2
16 3 9 13 0 9 2 3 13 9 2 16 3 13 10 0 2
20 16 0 3 3 13 13 2 0 3 13 0 9 13 7 0 9 3 9 3 2
23 3 3 15 3 3 13 0 9 2 3 8 15 15 9 2 16 3 15 0 9 13 13 2
6 10 3 13 0 9 2
9 3 3 15 15 13 7 3 13 2
5 15 3 13 9 2
6 0 3 1 9 13 2
8 3 3 15 9 13 1 9 2
4 15 13 13 2
35 7 15 0 13 0 2 16 3 13 2 7 0 13 7 3 0 13 9 2 16 0 13 9 0 9 0 2 16 3 0 0 13 9 2 2
9 2 3 15 15 0 3 3 13 2
12 9 9 0 13 13 9 2 3 9 0 13 2
26 3 3 3 1 9 13 7 9 13 1 0 9 1 0 9 2 1 9 1 9 2 13 3 0 9 2
17 9 3 15 15 13 1 9 1 9 2 1 9 9 1 9 0 2
55 9 3 0 0 13 13 1 9 2 16 3 3 9 13 13 9 9 2 15 3 13 3 13 2 7 3 1 9 9 13 9 1 0 2 15 15 9 3 9 3 13 2 16 3 15 9 1 9 13 13 1 9 9 0 2
4 3 3 13 2
8 3 3 15 3 9 13 9 2
33 3 3 3 13 1 9 0 9 2 7 3 3 0 13 0 9 9 1 0 2 0 3 15 9 13 0 2 15 3 0 13 0 2
25 3 3 15 15 13 2 16 1 9 0 13 7 16 13 13 2 7 3 9 13 7 9 3 13 2
19 3 3 3 0 3 0 1 9 9 13 2 3 16 3 3 0 9 13 2
9 13 16 3 13 2 16 0 13 2
34 3 3 9 3 7 9 0 13 0 2 16 3 3 13 0 2 16 3 15 1 9 13 2 3 3 0 0 10 0 13 0 1 9 2
8 10 3 3 9 13 0 13 2
14 9 3 3 15 13 10 13 2 3 15 3 3 13 2
19 7 3 15 3 13 0 3 15 13 9 9 2 15 9 0 1 9 13 2
21 3 3 15 0 13 0 9 2 10 15 1 13 13 2 16 15 15 0 13 2 2
18 2 3 3 15 9 3 9 0 3 13 2 16 15 3 0 13 9 2
9 3 3 15 15 13 7 3 13 2
9 15 9 2 15 3 9 15 13 2
10 3 3 15 13 3 13 13 1 9 2
14 13 3 9 9 0 13 2 15 15 0 3 13 2 2
8 15 3 3 9 13 0 13 2
43 3 3 3 13 9 0 13 2 15 0 3 0 13 1 0 9 2 16 3 3 13 3 3 13 2 7 1 15 9 13 9 1 9 2 7 0 1 9 2 16 9 13 2
18 3 3 15 9 3 13 9 2 7 3 7 15 9 0 9 13 3 2
7 3 3 15 3 9 13 2
12 13 0 0 2 15 3 9 3 9 3 13 2
17 3 3 3 0 13 13 0 2 16 3 15 0 9 0 9 13 2
7 15 3 13 13 9 0 2
8 3 3 15 13 3 0 2 2
7 15 3 13 13 9 9 2
8 0 3 0 3 13 0 3 2
12 15 3 13 13 2 16 3 9 13 1 9 2
10 7 3 3 3 13 7 0 13 9 2
16 3 1 9 13 9 0 9 13 0 2 9 3 1 9 13 2
24 9 3 1 0 13 13 2 9 3 2 16 15 9 13 13 2 3 13 1 9 9 0 13 2
10 15 3 0 3 13 2 16 3 13 2
18 16 3 3 9 9 7 9 13 2 3 3 3 13 3 3 13 9 2
29 3 16 3 0 13 3 7 13 2 13 3 3 1 9 7 1 9 16 3 9 1 9 0 13 7 9 7 3 2
13 3 8 3 15 13 9 13 2 16 3 0 13 2
17 3 15 1 9 0 13 3 7 9 2 15 3 15 3 13 13 2
11 15 3 0 13 2 7 0 13 9 2 2
8 15 3 3 9 13 0 13 2
46 3 3 3 13 2 13 3 9 2 16 13 3 13 3 0 9 2 9 13 1 9 13 2 13 1 9 2 0 2 3 0 2 15 15 9 13 1 15 2 0 0 9 9 13 2 2
11 2 3 15 3 3 13 2 13 3 9 2
21 9 3 15 3 15 13 0 9 13 2 3 13 13 3 13 2 3 3 0 13 2
7 15 3 0 13 9 2 2
9 15 3 9 15 13 13 1 9 2
5 13 3 9 13 2
7 3 3 9 13 0 9 2
12 15 3 9 13 0 2 15 3 9 13 13 2
14 15 3 0 9 13 0 2 15 1 9 13 9 9 2
18 9 3 0 13 15 9 2 3 0 2 1 15 3 7 9 12 13 2
23 15 3 16 3 9 13 0 9 2 13 3 1 9 9 3 0 2 1 9 13 0 9 2
8 9 3 3 15 0 3 13 2
7 13 3 3 13 0 9 2
13 10 9 3 15 13 13 2 15 3 9 9 13 2
23 0 3 13 9 0 2 15 3 15 3 1 9 0 9 13 2 16 15 3 13 9 0 2
19 0 3 9 13 13 3 2 9 2 15 9 0 1 9 7 0 9 2 2
8 15 3 3 9 13 0 13 2
13 10 3 9 3 13 9 2 15 15 13 0 13 2
8 15 3 13 9 7 9 13 2
10 9 3 9 13 0 2 3 3 15 2
8 15 3 9 13 1 9 2 2
7 15 3 13 3 3 13 2
7 15 3 9 13 13 9 2
13 0 3 13 9 2 0 9 13 2 13 1 9 2
8 0 3 3 9 1 13 2 2
19 2 3 13 2 15 3 3 0 3 1 9 13 9 13 2 15 3 13 2
17 3 15 3 1 0 9 9 9 13 2 15 15 9 0 13 2 2
8 15 3 3 9 13 0 13 2
9 3 3 0 13 9 3 13 13 2
8 3 13 0 0 1 9 13 2
28 3 3 3 9 0 13 3 0 0 1 0 9 2 0 7 0 2 10 3 15 15 13 2 16 13 0 9 2
9 9 3 0 13 7 9 15 13 2
15 7 15 9 9 13 13 2 3 0 0 9 13 15 13 2
9 0 13 3 13 2 3 13 13 2
8 15 3 3 9 13 0 13 2
23 3 3 9 3 13 2 16 3 13 2 7 9 13 2 15 15 9 1 9 13 9 13 2
10 3 13 9 2 9 3 0 9 13 2
8 15 3 13 0 1 9 13 2
7 3 3 13 13 3 0 2
22 9 3 2 3 15 9 0 9 0 13 0 1 9 2 3 13 1 9 0 9 13 2
18 10 15 3 13 9 13 2 7 15 3 9 13 2 7 13 0 13 2
17 13 3 9 9 3 0 2 13 3 1 9 2 0 3 13 9 2
8 7 10 3 9 0 13 9 2
17 3 10 3 0 2 13 9 9 2 13 9 15 9 15 13 9 2
7 2 9 3 1 9 13 2
14 3 3 13 9 9 2 0 0 9 2 0 1 9 2
9 3 15 3 9 13 9 13 9 2
26 15 3 3 1 9 0 7 9 0 13 2 1 3 15 9 0 13 2 0 3 3 9 13 9 9 2
15 9 3 3 1 0 9 13 1 3 9 7 1 0 9 2
9 3 3 15 13 9 7 9 0 2
9 7 3 15 15 0 1 9 13 2
21 3 16 3 3 15 9 13 7 13 13 2 3 3 15 0 13 2 13 3 9 2
15 13 3 15 13 9 9 0 2 3 3 9 9 13 9 2
16 0 3 9 9 13 9 2 7 13 7 13 2 15 3 13 2
16 9 3 1 0 13 9 0 0 2 16 3 15 13 0 3 2
14 3 15 9 9 13 13 2 16 13 9 3 7 0 2
6 3 3 3 13 13 2
5 0 3 13 9 2
25 2 3 3 3 13 9 3 7 9 2 10 9 3 3 13 0 9 2 7 3 13 13 3 13 2
9 3 3 15 13 13 1 0 0 2
22 0 3 1 9 13 0 0 9 2 15 3 3 0 9 13 3 13 0 1 9 13 2
9 3 3 15 15 13 13 9 9 2
10 2 3 13 2 9 3 0 13 9 2
10 9 3 13 2 9 3 1 0 13 2
25 3 15 3 13 1 9 0 13 2 7 13 1 9 13 1 9 2 7 0 13 7 3 0 13 2
11 3 13 7 13 2 13 3 1 9 13 2
15 15 3 13 0 9 9 3 1 9 9 2 13 3 9 2
22 3 16 9 3 13 7 9 2 3 3 15 9 3 13 7 9 13 1 9 0 9 2
12 15 3 13 13 1 0 3 9 7 0 9 2
10 13 3 1 9 1 9 1 9 13 2
9 15 3 1 9 13 1 3 13 2
6 15 15 0 13 9 2
19 3 3 15 3 13 2 16 13 9 0 7 9 7 16 3 15 0 13 2
12 2 13 15 9 3 0 1 15 3 9 0 2
5 9 3 13 9 2
18 3 3 15 9 13 13 3 3 13 9 10 2 15 3 9 13 9 2
9 13 2 16 3 9 13 15 13 2
15 13 3 9 9 1 9 0 0 9 2 16 3 13 9 2
18 3 3 0 9 0 13 9 2 15 3 13 2 15 3 0 9 13 2
9 3 3 9 3 7 9 13 9 2
38 3 16 1 9 0 13 2 15 1 9 0 13 3 3 2 9 3 0 0 0 1 9 13 2 0 3 9 13 2 3 15 3 3 0 13 9 9 2
9 15 3 3 1 9 0 13 0 2
23 3 3 3 3 13 9 3 1 0 2 3 3 0 3 3 0 2 0 3 13 3 9 2
7 13 3 9 1 0 13 2
19 3 3 3 3 9 3 3 9 13 9 2 9 3 0 13 1 9 13 2
26 3 3 15 9 13 13 13 2 15 15 9 13 1 9 9 13 2 9 12 13 2 0 9 3 13 2
9 15 3 3 1 9 13 0 9 2
7 3 3 9 1 9 13 2
9 15 3 3 3 9 13 0 9 2
7 3 9 13 9 13 9 2
9 15 3 12 13 9 1 9 13 2
7 3 15 13 9 1 9 2
15 3 3 0 9 1 9 13 9 3 13 9 3 3 13 2
8 9 3 3 13 0 9 13 2
23 16 15 15 13 9 0 1 2 3 3 15 9 0 13 1 9 15 1 9 13 9 0 2
14 3 3 0 9 13 13 13 9 2 16 1 9 13 2
9 15 3 9 0 13 2 13 9 2
10 3 3 1 9 0 13 9 9 0 2
7 3 10 0 0 3 13 2
16 2 3 3 3 13 13 9 2 0 1 9 2 0 13 9 2
6 9 3 1 9 13 2
15 0 3 13 0 9 9 3 1 9 2 15 9 13 9 2
16 3 3 1 9 9 13 9 0 1 9 2 7 15 9 13 2
18 3 3 13 12 3 9 7 12 9 13 3 9 3 7 9 9 13 2
34 3 16 3 0 9 0 13 9 2 3 3 15 0 9 13 7 9 0 3 1 9 13 1 9 2 16 3 9 13 9 9 3 13 2
25 13 3 9 1 0 13 2 7 15 13 9 1 9 9 2 9 1 9 2 1 9 0 7 9 2
17 13 3 3 1 9 7 1 9 13 7 13 2 16 13 0 9 2
23 3 3 15 13 13 0 13 2 0 13 1 9 0 7 9 9 9 9 13 13 3 13 2
29 3 16 3 1 13 13 9 9 2 3 3 15 15 9 13 0 13 2 15 3 15 0 9 0 1 9 0 13 2
9 15 3 3 13 1 9 9 13 2
7 3 3 15 13 9 9 2
19 10 3 3 9 0 13 2 1 3 13 1 9 13 2 1 3 13 9 2
10 15 3 15 13 9 0 1 9 13 2
43 3 15 13 9 3 9 3 2 9 3 2 0 3 9 2 0 3 13 13 9 0 9 2 13 3 3 13 1 9 0 9 13 2 16 3 3 13 1 9 9 13 0 2
6 3 3 0 9 13 2
15 1 3 13 1 9 2 13 3 9 0 9 3 9 0 2
20 3 3 2 16 1 9 0 9 3 9 3 2 13 9 2 3 3 13 9 2
21 2 3 13 2 15 3 3 0 9 13 2 1 3 13 1 9 9 0 13 9 2
6 3 3 0 9 13 2
12 3 16 13 13 9 2 9 13 13 0 9 2
17 3 3 3 0 9 1 9 13 13 13 9 3 0 7 9 0 2
16 16 3 9 13 7 1 9 13 2 3 3 13 1 9 9 2
16 16 3 9 13 0 9 2 3 3 15 9 13 1 0 13 2
9 3 13 0 16 15 3 13 9 2
6 15 3 3 13 13 2
14 13 3 9 1 0 13 9 2 15 1 9 0 13 2
5 0 3 0 13 2
12 9 3 1 0 13 9 1 9 0 7 9 2
8 13 3 3 0 1 9 13 2
8 3 3 3 15 9 13 13 2
15 2 3 15 3 0 0 9 13 2 9 3 1 0 13 2
10 15 3 15 13 2 15 3 9 0 2
8 9 3 1 9 0 13 3 2
7 1 3 13 9 9 9 2
13 13 3 13 2 3 15 3 12 7 12 9 13 2
7 1 3 15 13 13 3 2
14 13 3 1 9 13 9 9 0 9 2 0 1 9 2
18 1 3 15 9 13 0 7 9 2 15 0 13 2 16 0 9 13 2
17 3 3 15 3 13 1 9 2 3 3 15 3 9 0 13 13 2
9 15 3 13 2 16 13 0 9 2
31 13 3 1 9 9 9 2 9 3 3 13 13 9 0 2 9 13 0 0 2 0 9 0 3 7 0 7 0 9 13 2
4 3 13 0 2
10 15 3 3 13 9 13 0 7 13 2
7 15 3 3 0 9 13 2
8 9 3 13 2 13 9 13 2
23 13 3 13 1 9 3 9 3 2 1 3 15 9 3 7 9 7 9 0 9 9 13 2
12 13 3 9 9 0 2 16 3 13 0 9 2
15 3 16 13 3 7 13 2 3 3 9 13 1 9 13 2
23 15 3 9 3 13 9 9 3 9 3 7 9 2 3 9 13 0 2 3 10 3 3 2
16 2 9 3 3 13 0 1 9 0 9 9 13 7 0 9 2
14 3 3 15 13 13 9 13 3 2 9 9 0 13 2
12 1 3 15 9 9 13 2 9 3 13 9 2
16 3 16 3 15 0 13 13 2 3 3 10 0 9 13 9 2
13 13 1 9 13 9 0 0 9 2 0 1 9 2
5 15 3 13 13 2
10 15 3 3 13 9 13 0 7 13 2
7 15 3 3 0 9 13 2
8 3 15 13 2 13 9 13 2
12 15 3 3 13 0 2 3 3 15 0 13 2
5 0 3 13 13 2
20 2 3 13 2 3 15 1 3 9 0 9 13 2 0 0 2 1 3 9 2
8 15 3 3 13 0 9 13 2
14 3 15 3 0 13 13 9 7 15 13 9 0 13 2
16 13 3 2 16 3 3 0 13 3 3 15 0 13 0 9 2
6 7 1 15 0 13 2
7 3 3 3 13 0 9 2
10 3 15 13 2 0 3 15 13 9 2
14 1 3 3 15 13 9 2 9 3 13 1 3 13 2
14 9 3 15 15 1 9 13 3 3 9 0 9 13 2
6 3 15 13 3 13 2
9 3 3 3 15 0 13 7 13 2
19 13 2 15 9 0 13 1 9 9 13 2 15 3 15 9 13 0 9 2
8 0 3 15 13 0 9 9 2
10 13 15 9 2 13 3 1 9 9 2
8 3 3 3 3 13 15 13 2
14 3 3 13 9 0 2 15 15 13 2 13 3 0 2
24 16 3 9 15 13 0 9 2 3 3 15 9 0 13 1 9 9 13 2 3 3 13 13 2
7 15 3 15 13 13 13 2
18 3 15 3 3 13 9 9 2 16 3 15 13 3 9 0 3 13 2
17 2 3 3 13 13 9 9 1 9 13 2 7 15 9 0 13 2
10 9 3 0 13 2 9 3 0 9 2
6 9 3 15 13 9 2
14 0 3 3 13 9 3 0 2 9 3 3 0 13 2
25 9 3 3 13 1 0 9 9 1 0 2 15 3 1 9 9 13 2 0 3 15 9 13 13 2
7 13 3 1 9 9 9 2
10 3 13 13 2 9 3 15 13 9 2
10 15 3 3 13 9 13 0 7 13 2
6 3 15 13 13 9 2
10 13 3 15 13 1 9 0 0 0 2
6 1 3 9 9 13 2
21 13 3 15 9 0 9 2 16 13 2 1 3 3 9 13 2 0 13 1 9 2
21 3 16 13 3 7 13 2 3 3 15 13 2 9 13 9 3 13 1 3 13 2
10 2 13 3 3 2 1 0 13 9 2
16 15 3 0 13 13 7 13 9 2 7 15 13 9 0 13 2
6 8 15 3 13 9 2
11 9 15 13 16 3 15 13 15 9 13 2
21 3 3 3 3 3 15 0 9 15 9 13 2 15 3 13 7 0 13 9 9 2
9 15 3 15 1 9 0 9 13 2
24 3 15 3 9 13 0 2 15 3 15 3 13 13 0 9 2 1 9 13 0 1 9 0 2
23 3 3 3 9 3 9 13 2 15 3 3 9 0 13 2 16 13 9 7 9 13 0 2
12 2 3 13 2 15 3 3 13 2 3 13 2
18 3 16 3 13 3 13 3 10 9 2 7 3 15 9 13 0 9 2
18 2 0 3 3 3 3 1 9 13 9 2 15 15 9 1 9 13 2
22 13 3 3 15 3 1 3 9 1 3 9 1 3 0 9 2 15 3 1 3 13 2
16 15 15 3 13 9 1 9 0 0 3 2 3 3 9 13 2
16 15 3 0 1 9 13 9 0 2 1 3 15 13 0 9 2
16 15 3 0 9 9 9 13 0 1 0 2 13 3 0 9 2
13 15 3 0 9 13 7 9 13 0 1 9 0 2
4 13 3 9 2
35 3 16 3 13 9 1 9 9 2 1 3 9 13 13 1 9 0 2 0 13 2 1 9 3 7 9 2 16 15 1 9 0 13 9 2
34 3 16 13 3 7 13 3 9 2 1 3 15 9 0 13 7 9 2 13 3 15 13 1 9 0 0 0 2 1 3 9 9 13 2
15 9 3 0 9 13 13 0 0 2 1 0 9 2 13 2
6 1 3 0 13 9 2
14 9 3 0 9 13 13 2 9 0 13 2 13 13 2
4 13 3 13 2
15 0 3 3 13 9 2 7 13 13 2 0 3 13 9 2
26 2 9 3 16 13 15 13 3 3 1 9 9 13 2 0 3 15 9 13 2 3 13 9 0 13 2
7 3 15 3 9 0 13 2
7 3 3 15 15 13 13 2
7 3 3 15 13 0 9 2
17 3 16 3 0 13 13 3 13 2 13 2 16 9 13 0 9 2
26 2 3 13 2 9 3 1 9 13 9 13 1 9 2 9 3 13 9 2 1 3 13 9 13 0 2
16 15 3 3 13 0 2 15 3 1 0 13 13 0 9 0 2
20 15 3 1 3 9 9 13 2 15 3 13 9 0 2 15 15 13 0 9 2
16 9 3 3 13 0 16 3 13 2 7 0 0 7 0 13 2
10 13 3 15 0 13 3 1 9 0 2
12 0 3 0 13 9 2 1 3 9 0 13 2
6 9 3 13 3 0 2
16 9 3 3 0 13 3 2 9 3 1 9 13 9 3 0 2
9 0 3 3 13 7 13 0 9 2
15 13 3 1 9 0 0 9 0 13 2 0 1 9 13 2
11 3 3 3 9 13 2 7 0 13 13 2
10 3 15 0 16 13 9 2 0 13 2
24 13 3 3 15 9 3 13 2 3 16 9 13 7 9 0 0 9 2 3 3 13 7 13 2
7 7 15 13 9 0 13 2
9 3 3 2 10 0 9 13 9 2
17 2 9 3 3 0 13 3 2 9 3 1 9 13 9 3 0 2
19 0 3 13 15 3 0 13 2 16 13 9 0 1 9 9 13 7 13 2
4 0 3 13 2
11 2 3 13 2 15 3 3 0 9 13 2
8 9 3 15 0 13 0 9 2
7 7 15 13 9 0 13 2
7 0 3 3 0 9 13 2
9 3 15 9 0 9 13 3 0 2
8 15 3 13 9 1 9 9 2
12 3 3 3 9 0 1 9 13 2 3 13 2
6 13 3 0 0 9 2
26 2 3 3 10 0 9 1 9 9 3 13 3 7 13 3 9 2 1 3 3 9 0 13 7 9 2
17 15 3 16 0 13 13 3 3 2 13 13 2 1 3 13 9 2
7 8 3 3 0 9 13 2
19 13 3 0 7 0 1 9 13 9 0 2 7 0 0 9 13 1 9 2
26 3 3 13 9 7 13 9 2 1 15 3 3 9 1 9 13 2 0 16 0 13 0 9 0 9 2
16 3 3 9 0 0 1 9 13 13 9 3 0 7 9 0 2
28 3 16 3 3 9 13 2 1 3 13 9 9 13 2 1 3 9 0 13 2 7 3 15 13 13 9 9 2
11 2 3 13 2 3 15 3 13 9 0 2
18 3 3 3 0 9 1 9 13 13 2 13 9 15 0 7 9 0 2
16 16 3 9 13 7 1 9 13 2 15 3 13 1 9 0 2
15 3 15 9 13 0 9 9 13 2 9 3 15 13 9 2
7 7 15 13 9 0 13 2
26 9 3 15 13 3 2 7 0 9 2 15 15 13 0 9 1 15 13 2 16 3 15 3 1 13 2
19 13 3 1 9 13 2 3 3 3 15 9 13 3 13 7 13 9 9 2
16 3 16 13 3 13 3 13 2 3 3 3 15 9 13 13 2
10 1 9 3 3 3 15 13 9 0 2
8 15 3 3 3 9 9 13 2
25 3 3 1 9 9 3 13 9 3 2 15 3 9 9 13 9 2 9 3 9 3 12 9 0 2
6 1 3 9 0 13 2
38 0 3 13 9 0 9 2 13 1 9 9 9 2 15 15 0 2 13 1 9 9 3 13 0 2 9 3 3 9 13 0 0 2 15 9 13 0 2
27 3 16 9 13 0 9 0 2 3 9 9 13 0 3 0 1 9 13 2 0 3 3 13 13 9 9 2
8 3 3 0 9 13 9 13 2
23 0 3 9 0 13 1 9 13 2 3 3 13 9 0 9 9 1 13 2 16 9 13 2
10 1 3 15 9 3 9 3 9 13 2
25 0 3 0 9 0 13 9 2 0 7 0 2 1 3 9 13 9 0 0 2 9 3 13 9 2
13 3 15 1 9 13 13 9 0 9 1 9 0 2
11 8 3 3 13 13 0 9 2 7 13 2
7 3 3 15 13 9 9 2
11 3 3 3 3 3 3 3 0 13 9 2
19 9 3 15 13 0 2 3 3 15 3 0 1 9 3 3 9 0 13 2
25 13 3 9 9 7 9 13 3 13 7 13 9 0 0 13 13 1 9 0 2 7 1 9 13 2
12 1 3 15 9 9 13 2 9 3 8 13 2
9 2 13 3 15 15 1 9 13 2
8 3 3 3 15 9 13 13 2
36 2 3 16 3 3 1 9 0 7 9 9 13 13 0 1 9 13 2 3 3 3 13 9 1 9 0 9 13 9 0 3 0 2 3 13 2
13 15 3 9 3 13 9 13 7 3 7 3 13 2
46 2 3 16 3 1 9 13 7 9 2 9 3 3 0 13 1 9 0 2 1 3 9 13 7 9 9 0 2 1 3 10 9 13 13 2 1 3 7 0 13 13 0 1 9 13 2
9 15 3 9 0 13 1 9 13 2
8 15 3 9 3 9 3 13 2
7 15 3 0 13 9 13 2
8 13 3 9 13 3 0 9 2
9 2 15 3 1 9 13 0 9 2
35 3 3 1 0 9 13 13 9 2 3 16 3 13 1 9 0 2 3 16 3 3 1 9 1 3 13 2 7 1 9 0 13 0 9 2
12 9 3 3 13 13 2 1 3 10 9 13 2
17 0 3 3 1 9 9 13 2 16 1 9 13 2 15 13 9 2
9 2 3 9 3 9 9 3 13 2
37 15 3 9 0 13 1 9 9 13 0 3 0 3 7 3 2 1 0 3 9 13 0 9 2 0 9 2 3 3 0 9 2 10 0 3 9 2
6 1 3 9 0 13 2
38 0 3 13 9 0 9 2 13 1 9 0 9 2 15 15 0 2 13 1 9 9 3 13 0 2 9 3 3 9 13 0 0 2 15 9 13 0 2
10 15 0 1 9 13 3 0 0 9 2
6 15 3 0 9 13 2
23 0 3 9 0 13 1 9 13 2 3 3 13 9 0 9 9 1 13 2 3 9 13 2
8 3 3 3 13 1 9 0 2
16 9 3 1 9 9 13 15 0 7 0 2 16 9 0 13 2
16 15 3 15 13 13 13 3 9 2 7 15 13 9 0 13 2
11 2 3 13 2 15 3 15 13 13 9 2
19 9 3 1 9 13 3 13 0 13 13 1 9 0 2 7 1 9 13 2
12 1 3 15 9 9 13 2 9 3 3 13 2
31 3 3 15 15 3 13 2 3 13 2 1 3 9 7 9 2 15 15 13 0 13 2 9 3 2 15 0 1 9 13 2
41 3 15 0 0 13 3 13 13 2 16 15 15 9 9 13 2 7 15 13 1 9 2 15 15 13 2 9 15 15 13 0 1 9 9 2 9 0 3 13 13 2
19 0 15 15 13 13 3 1 9 9 2 15 7 0 13 13 1 0 9 2
9 15 3 15 13 13 13 3 9 2
19 3 3 3 3 13 0 2 0 3 13 2 9 1 13 2 3 9 13 2
17 2 13 3 1 9 0 9 0 9 13 2 15 3 13 7 13 2
17 3 13 9 2 13 3 9 0 2 9 16 13 7 15 0 13 2
12 2 3 13 2 15 3 13 9 0 9 13 2
7 15 3 15 0 13 9 2
18 3 3 13 13 9 2 15 15 9 13 9 13 16 15 9 0 13 2
49 3 3 3 3 3 3 0 3 13 13 2 16 3 13 0 9 13 7 9 2 16 3 0 13 0 9 9 9 2 13 0 9 2 13 3 13 9 7 0 9 9 2 15 0 13 7 0 13 2
20 15 16 3 3 0 13 9 3 13 2 3 3 3 1 9 0 3 13 13 2
20 0 3 16 3 3 13 2 3 3 13 2 13 1 0 9 2 9 1 0 2
9 3 3 3 0 3 9 13 13 2
40 3 16 9 1 9 0 13 7 9 7 3 0 9 2 13 3 3 13 0 9 2 1 15 3 15 13 15 3 13 9 9 2 3 3 3 9 13 9 13 2
19 3 3 3 15 3 13 9 0 3 3 0 9 2 15 3 9 9 13 2
12 9 3 15 13 3 0 2 3 3 15 13 2
20 9 3 15 1 9 0 0 3 0 13 2 15 3 15 13 9 1 0 13 2
6 3 3 9 0 13 2
6 15 3 15 0 13 2
10 2 3 13 2 3 15 15 13 13 2
9 3 3 15 15 13 7 3 13 2
6 9 15 13 9 13 2
18 15 3 0 13 1 9 2 3 3 0 9 13 3 13 3 3 13 2
11 2 3 13 2 15 3 15 3 13 13 2
10 2 0 15 9 13 7 1 9 13 2
17 15 15 3 3 13 9 13 9 1 13 2 15 3 15 0 13 2
12 15 3 3 13 2 15 3 3 3 13 3 2
15 3 15 3 13 0 2 16 1 9 13 7 13 9 0 2
11 3 3 13 2 7 15 13 9 0 13 2
14 3 3 3 3 13 3 13 9 3 7 9 0 9 2
14 3 3 3 13 1 9 2 3 3 13 1 9 9 2
10 2 3 13 2 3 15 15 13 13 2
35 3 3 3 1 13 9 2 3 3 3 0 9 13 2 7 3 13 13 9 2 1 15 10 0 13 9 0 0 1 0 2 16 9 13 2
9 3 3 15 15 13 7 3 13 2
8 15 3 15 9 13 0 9 2
13 7 0 9 2 7 9 9 0 0 9 13 13 2
12 2 3 3 0 3 13 13 9 0 1 9 2
12 0 3 15 3 13 9 3 7 9 9 13 2
25 0 3 3 3 15 13 0 9 2 7 0 9 9 13 7 9 0 13 2 15 13 9 9 13 2
4 0 3 13 2
20 3 16 13 9 13 3 9 2 3 15 1 9 9 0 9 13 0 13 9 2
21 3 15 3 13 13 2 0 3 9 9 13 0 9 13 2 0 3 1 9 13 2
9 3 3 3 15 13 7 9 13 2
31 3 3 15 3 1 9 0 9 0 0 9 13 13 2 3 3 15 3 15 9 13 2 15 3 3 9 0 9 13 9 2
22 3 3 13 2 13 3 15 9 13 2 3 3 15 1 9 9 0 7 3 9 13 2
15 15 3 9 0 13 3 3 2 7 15 13 9 0 13 2
15 3 15 15 9 15 0 9 13 2 16 3 3 13 13 2
35 3 3 3 9 3 7 9 9 13 2 7 15 3 3 9 0 9 13 13 2 16 3 0 13 0 9 9 2 9 3 3 9 13 13 2
5 3 3 0 13 2
12 0 3 0 13 2 16 3 3 0 13 9 2
15 15 3 1 9 0 0 13 2 3 15 13 16 13 0 2
9 15 3 15 1 9 0 13 9 2
14 13 0 9 0 1 9 3 13 13 3 0 9 0 2
11 15 3 0 13 2 7 0 0 9 13 2
5 15 3 13 0 2
23 2 3 3 3 0 9 13 0 2 15 13 9 0 0 13 2 13 3 9 9 13 9 2
12 15 3 3 13 0 9 1 9 9 13 0 2
18 0 3 3 9 13 2 9 0 2 13 2 13 3 9 0 3 9 2
10 13 3 0 9 2 1 3 9 13 2
22 3 16 3 13 9 0 9 2 1 3 3 15 13 9 2 9 3 13 1 3 13 2
13 13 3 9 13 0 9 2 16 3 0 9 0 2
12 3 3 13 1 9 2 7 13 3 3 13 2
7 3 15 3 13 9 9 2
16 15 3 13 9 13 7 9 2 15 0 9 9 0 13 0 2
7 15 3 0 9 13 13 2
7 3 3 0 9 13 9 2
15 3 15 3 1 9 0 9 13 0 13 9 0 1 9 2
19 15 3 13 1 9 9 0 2 13 9 0 1 0 9 2 0 9 13 2
18 3 3 3 9 15 13 15 3 9 9 0 1 9 13 9 0 0 2
8 15 3 0 13 9 0 13 2
27 3 16 3 9 3 7 9 13 3 13 9 7 13 9 2 3 3 3 15 13 9 0 2 0 0 13 2
5 9 3 13 9 2
6 9 3 13 0 9 2
15 0 3 15 3 7 0 13 9 2 3 9 3 13 0 2
17 9 1 9 13 13 2 3 1 9 9 0 2 16 9 0 13 2
10 3 3 3 13 2 16 9 9 13 2
24 3 13 9 9 2 15 0 13 9 2 0 2 16 15 1 9 9 13 13 3 9 0 9 2
11 3 3 15 9 13 9 1 0 9 9 2
17 2 9 3 9 3 13 0 3 9 2 15 9 0 9 13 0 2
17 0 3 3 3 15 13 3 3 13 2 0 9 9 13 7 9 2
8 3 3 3 3 9 13 0 2
8 9 3 9 15 3 13 2 2
19 2 3 13 2 15 3 3 0 3 13 9 2 9 3 13 1 9 0 2
7 15 3 9 0 13 9 2
11 9 3 3 0 13 2 0 3 13 9 2
13 3 3 13 13 2 3 3 10 9 3 13 13 2
11 0 3 15 9 1 9 9 9 13 2 2
3 3 13 2
11 9 3 1 15 13 9 3 9 3 2 2
17 2 0 3 3 3 13 9 2 16 3 15 3 0 9 0 13 2
20 9 3 13 3 3 9 13 3 3 13 1 3 2 1 15 3 0 9 13 2
10 9 3 9 13 0 2 3 3 15 2
8 15 3 9 13 1 9 2 2
7 15 3 13 13 0 9 2
16 7 3 0 7 0 9 13 0 2 0 15 3 13 13 2 2
15 3 3 3 9 13 1 9 2 15 3 15 13 0 9 2
19 3 3 1 9 0 13 2 16 15 15 13 1 9 10 0 9 13 2 2
7 15 3 13 13 0 9 2
21 2 3 16 9 3 13 3 3 0 9 9 0 2 13 3 1 9 9 9 13 2
16 1 3 0 13 2 0 1 0 9 1 9 13 7 9 13 2
11 13 3 3 15 0 2 16 13 9 0 2
19 13 3 15 3 3 2 0 1 9 13 2 13 1 15 9 2 13 13 2
21 3 3 3 15 3 13 9 0 3 3 15 9 2 0 3 3 13 1 0 9 2
17 2 15 3 15 13 13 13 3 9 2 7 15 13 9 0 13 2
13 7 15 3 1 9 9 13 13 0 9 0 9 2
21 7 15 0 9 13 1 9 9 13 7 9 9 0 2 7 1 9 13 7 9 2
11 2 3 13 2 15 3 15 3 13 13 2
5 3 13 0 9 2
26 1 3 0 9 3 13 9 3 0 2 15 3 3 1 0 9 0 13 7 9 7 9 7 9 13 2
14 3 3 0 9 9 13 2 3 13 7 1 0 9 2
22 15 3 9 13 2 3 3 15 13 13 3 1 9 9 1 9 13 1 3 9 13 2
13 0 3 7 0 13 9 0 2 0 13 9 9 2
12 3 3 13 3 0 9 7 9 0 3 13 2
22 15 3 3 0 13 15 3 1 9 13 7 13 3 0 9 2 3 15 3 0 13 2
14 9 3 13 1 0 2 0 3 9 9 13 3 13 2
11 2 3 13 2 15 3 15 3 13 13 2
12 2 3 3 3 3 3 15 9 3 0 13 2
22 3 15 9 0 13 2 15 3 3 13 2 7 15 3 13 2 15 3 3 13 13 2
11 3 3 15 9 3 0 13 15 13 3 2
19 9 3 15 13 1 9 0 2 15 3 3 3 1 9 13 9 2 0 2
18 3 3 15 3 9 0 13 13 2 7 0 9 13 2 15 9 13 2
12 10 3 0 3 3 3 9 13 9 9 13 2
7 3 3 15 13 3 0 2
12 0 3 15 13 2 15 3 1 9 13 0 2
13 3 2 3 3 3 2 0 1 0 9 9 13 2
9 3 3 3 13 1 9 0 9 2
11 3 3 15 13 2 13 15 3 7 13 2
28 13 3 1 9 8 9 7 9 7 0 9 9 3 2 15 0 13 9 3 9 3 10 0 9 1 0 9 2
13 13 3 9 15 0 9 7 3 13 9 0 13 2
10 2 3 13 2 3 15 15 13 13 2
19 3 3 3 1 13 9 2 3 3 3 0 9 13 2 7 3 13 0 2
18 3 3 3 15 0 13 0 9 0 2 3 3 0 13 9 3 13 2
11 2 3 13 2 15 3 15 3 13 13 2
23 13 3 0 13 13 0 2 9 1 0 2 15 3 9 0 13 2 7 0 9 13 13 2
17 3 3 15 13 9 7 9 0 2 15 0 13 13 3 1 9 2
15 0 3 15 15 0 1 9 0 13 1 9 1 0 0 2
17 3 3 16 1 9 9 13 9 2 3 0 13 7 3 13 9 2
7 9 0 7 15 13 0 2
8 0 3 0 13 1 9 0 2
19 0 3 3 3 3 15 13 9 3 3 13 9 0 3 3 9 9 13 2
22 15 3 3 3 0 13 3 13 2 9 3 13 9 7 9 0 2 0 3 9 13 2
36 3 16 3 9 9 13 0 2 9 7 9 0 13 1 9 13 0 2 3 3 3 13 0 9 3 3 0 13 2 0 3 0 13 1 9 2
6 3 3 3 13 9 2
23 2 3 13 2 9 3 0 9 13 0 13 1 0 9 2 0 15 15 9 13 0 13 2
15 2 10 3 0 9 9 13 13 13 2 13 3 9 0 2
23 0 3 9 9 9 3 13 2 13 1 9 2 15 15 15 13 13 1 9 9 1 9 2
5 13 3 9 9 2
8 9 3 9 13 7 9 9 2
9 3 3 3 13 13 15 1 9 2
7 15 3 15 9 13 0 2
11 15 3 0 0 9 9 8 13 13 3 2
7 13 3 9 7 0 9 2
11 3 3 3 13 13 2 7 3 15 15 2
13 3 15 13 9 1 9 0 10 0 9 13 13 2
28 2 15 3 1 9 0 13 9 3 13 1 0 9 2 15 0 13 1 0 9 9 13 9 0 2 3 0 2
25 15 3 1 12 13 9 2 9 3 15 3 13 9 13 2 9 3 13 2 15 3 3 13 9 2
12 2 7 3 9 13 0 9 13 13 1 9 2
5 15 3 13 9 2
10 13 3 13 2 13 3 3 13 13 2
24 3 3 13 10 9 13 13 2 3 9 13 13 2 1 3 9 9 0 13 2 13 3 9 2
17 15 3 13 10 9 1 9 13 2 15 3 9 13 1 9 0 2
13 2 7 3 9 13 0 9 13 9 13 0 0 2
15 3 3 15 3 13 9 3 9 3 9 3 13 1 9 2
10 3 16 13 9 13 2 3 13 9 2
7 3 3 3 13 9 0 2
20 3 15 3 3 13 13 2 1 3 9 13 1 9 2 9 3 1 9 13 2
15 3 13 3 3 0 15 13 2 15 0 9 0 13 9 2
17 13 3 3 15 0 2 16 13 9 2 7 15 13 9 0 13 2
11 9 3 9 13 9 2 3 9 13 0 2
14 3 3 0 0 9 13 2 15 3 15 0 13 9 2
8 7 3 15 3 13 9 13 2
12 3 3 3 0 13 15 3 15 0 13 9 2
9 15 3 15 13 7 13 1 9 2
8 9 3 15 13 7 0 9 2
10 3 3 1 9 13 0 0 9 0 2
18 15 3 0 9 13 2 16 15 0 9 0 9 1 9 13 0 9 2
16 2 3 3 1 9 13 13 9 0 3 13 1 3 0 13 2
9 15 3 3 13 7 1 9 13 2
7 3 3 13 13 9 0 2
17 9 3 3 13 2 7 0 13 9 2 13 13 0 1 9 13 2
21 3 16 9 3 13 7 9 9 2 9 13 7 1 9 13 13 0 9 0 9 2
7 2 15 3 10 0 13 2
15 3 3 3 9 1 9 13 13 2 7 3 3 13 13 2
14 1 3 0 13 0 9 7 9 0 7 0 9 0 2
10 3 3 13 9 7 13 9 3 0 2
6 1 3 9 13 13 2
22 3 15 13 9 7 0 13 2 16 3 15 9 0 7 9 7 1 9 13 9 13 2
17 3 3 3 0 9 1 9 13 13 13 9 3 0 7 9 0 2
32 3 3 9 13 7 1 9 13 2 15 3 13 1 0 9 2 15 3 15 9 13 0 1 9 13 3 7 13 7 13 0 2
8 3 15 15 0 1 9 13 2
9 7 3 3 15 9 13 9 9 2
23 8 0 3 3 0 13 2 15 3 13 2 3 15 15 13 2 13 3 15 3 9 0 2
16 9 3 0 13 2 15 3 3 0 9 13 2 15 15 13 2
18 3 13 2 1 3 9 13 9 9 13 0 2 16 15 13 10 0 2
33 3 0 13 16 3 13 2 13 15 1 9 0 9 3 9 3 0 1 9 2 1 3 0 9 13 2 16 3 13 9 13 9 2
19 16 3 3 13 9 13 3 13 2 15 3 15 3 0 3 1 9 13 2
28 3 16 3 15 3 1 13 9 2 3 15 3 3 3 13 2 0 3 15 9 13 2 7 3 0 9 13 2
5 13 3 15 3 2
15 3 3 3 9 0 2 1 3 0 9 0 13 0 9 2
9 9 3 3 15 3 9 0 13 2
28 3 3 3 3 3 0 13 3 3 9 0 2 15 3 9 9 9 13 2 7 3 3 15 3 13 0 9 2
7 3 0 13 9 0 13 2
30 15 3 3 3 15 9 13 9 2 15 15 13 2 7 3 3 9 3 9 7 9 9 9 9 13 9 3 0 9 2
20 3 3 3 15 3 3 13 0 1 9 2 7 9 13 2 16 0 13 9 2
22 15 3 3 3 13 2 3 3 3 9 0 13 9 3 3 1 9 3 3 1 9 2
21 3 3 3 13 0 9 3 3 13 2 3 3 16 15 9 3 12 7 9 13 2
8 9 3 0 13 2 0 13 2
14 3 3 3 1 9 0 0 9 9 13 0 9 13 2
8 3 3 1 9 13 0 13 2
16 15 3 3 9 3 0 9 0 13 2 0 3 3 9 0 2
34 15 3 3 9 13 12 0 0 2 12 3 3 15 9 0 2 1 3 0 0 9 2 1 3 0 9 0 7 0 2 0 0 9 2
40 0 3 3 1 9 0 13 2 1 3 13 9 0 9 2 3 3 13 2 9 13 2 9 3 9 3 2 3 16 3 0 13 9 2 15 0 13 0 9 2
12 15 3 3 3 3 9 0 13 13 1 9 2
10 13 3 3 9 0 9 13 9 0 2
4 7 3 13 2
10 15 3 1 9 13 0 2 9 13 2
9 15 3 1 0 9 13 0 9 2
13 3 3 3 3 13 1 9 2 3 3 13 0 2
9 3 15 3 3 13 2 16 13 2
11 3 3 3 13 15 1 0 3 3 9 2
24 3 3 9 9 13 3 9 3 13 2 16 3 0 0 13 12 9 1 9 13 7 3 0 2
10 2 3 13 2 3 15 15 13 13 2
6 3 3 9 13 0 2
21 15 3 3 3 0 2 7 0 0 13 2 0 3 0 3 7 0 3 3 0 2
6 3 3 15 13 9 2
23 16 3 13 13 1 9 2 13 2 16 15 3 13 13 0 9 2 0 3 1 9 13 2
8 15 15 3 13 1 9 13 2
7 2 9 3 1 9 13 2
11 9 3 3 13 0 2 3 3 3 13 2
22 15 3 3 13 13 3 9 9 9 1 9 13 3 13 2 9 13 0 7 9 9 2
21 15 16 3 3 0 13 9 3 13 2 3 3 3 3 1 9 0 3 13 13 2
16 0 3 16 3 3 13 2 3 3 13 2 13 1 0 9 2
15 3 15 1 9 13 13 9 0 3 13 1 3 0 13 2
9 15 3 3 13 7 1 9 13 2
8 3 3 13 0 9 13 9 2
9 3 3 9 0 13 1 9 13 2
8 15 3 9 3 9 3 13 2
9 2 3 3 15 9 13 13 9 2
18 3 13 3 15 2 16 13 7 3 13 7 3 13 9 7 9 13 2
11 9 3 0 13 0 9 13 7 9 0 2
6 0 15 13 9 13 2
22 3 15 9 13 1 0 2 16 0 3 13 2 0 1 9 2 1 3 0 9 13 2
17 16 3 3 13 15 13 3 13 2 15 3 0 3 1 9 13 2
9 3 3 3 13 9 0 9 9 2
5 13 3 9 0 2
15 3 3 9 3 13 7 9 13 0 2 13 3 9 9 2
24 13 3 9 9 9 13 7 15 3 1 9 0 13 2 15 3 1 9 13 13 9 0 9 2
13 3 15 9 0 9 0 9 0 13 9 0 13 2
15 3 3 13 9 2 16 13 0 9 9 3 9 9 9 2
8 3 3 9 1 9 0 13 2
21 15 3 1 9 15 13 3 9 3 9 3 0 1 9 2 1 3 0 9 13 2
8 0 3 13 0 9 13 9 2
26 3 16 0 13 0 3 13 13 2 3 13 2 15 3 3 13 0 9 3 13 2 0 3 13 9 2
27 3 3 3 15 3 13 9 0 2 16 3 15 9 1 9 9 13 2 7 15 3 13 13 7 0 13 2
24 13 3 3 0 0 1 9 0 0 9 3 9 9 13 2 13 3 2 0 13 1 9 9 2
7 2 3 13 13 9 0 2
13 3 0 9 13 13 2 13 3 13 9 9 13 2
5 15 3 13 13 2
39 3 16 3 15 3 13 2 3 3 3 3 9 9 13 3 3 3 9 2 3 1 9 13 0 0 9 2 15 15 1 9 13 2 15 3 1 9 13 2
19 2 3 16 3 10 9 13 2 3 3 9 7 0 9 13 7 9 13 2
16 15 3 3 13 1 9 13 9 2 13 3 3 0 1 9 2
12 13 3 3 9 2 16 3 9 0 9 13 2
18 3 3 3 15 0 13 0 2 16 16 9 13 1 9 0 0 9 2
12 3 3 3 2 3 7 15 13 2 13 0 2
22 15 3 9 9 9 0 13 9 13 2 16 3 3 9 13 15 3 9 13 7 13 2
11 3 1 9 13 2 16 9 0 9 13 2
25 0 3 9 7 9 1 13 9 2 15 3 9 13 2 16 15 13 3 13 7 1 0 15 13 2
16 3 3 3 9 3 9 0 13 2 16 3 15 15 13 13 2
18 3 15 13 0 9 7 12 9 0 1 9 13 1 9 9 13 9 2
16 3 3 3 13 13 2 13 3 15 9 3 13 1 0 9 2
7 2 15 3 0 13 13 2
14 3 3 9 2 3 3 0 9 0 13 9 0 9 2
25 3 16 13 9 0 9 2 0 3 13 13 2 3 3 9 0 13 2 3 3 9 13 9 0 2
6 15 3 0 9 13 2
8 15 3 1 15 13 13 9 2
19 3 3 15 9 0 1 9 9 12 13 2 15 9 3 9 3 0 13 2
19 13 3 1 9 0 3 7 1 9 3 15 13 9 7 9 3 3 13 2
37 3 3 16 1 9 9 0 9 9 10 0 9 1 9 13 1 9 13 9 9 0 2 13 3 3 13 13 3 2 3 15 3 13 13 1 9 2
14 0 3 0 0 13 9 0 2 0 13 9 9 13 2
19 2 3 16 9 13 0 3 9 9 3 2 3 3 9 1 0 9 13 2
18 3 3 15 3 9 13 1 9 0 9 3 13 9 13 9 3 9 2
8 3 3 15 9 13 13 9 2
8 3 3 0 0 13 15 13 2
8 3 1 10 9 13 9 0 2
10 2 3 13 2 15 3 13 0 9 2
8 3 3 9 0 15 13 9 2
10 1 15 9 2 3 3 15 9 13 2
45 3 3 3 15 3 0 0 13 2 15 3 9 9 13 7 7 9 3 13 9 13 2 3 3 3 9 1 0 0 13 9 2 7 3 1 9 0 13 13 9 13 1 0 9 2
23 3 3 3 3 3 13 9 0 9 3 13 0 1 9 13 2 3 3 13 13 0 9 2
17 3 3 3 13 15 3 0 13 9 2 7 15 13 9 0 13 2
9 3 3 3 15 0 13 0 9 2
24 16 3 15 7 9 9 7 9 0 9 13 2 3 3 15 9 0 7 9 7 15 9 13 2
10 7 0 13 9 2 15 0 13 9 2
31 3 16 3 13 3 13 3 10 9 2 13 1 9 0 0 9 1 9 0 2 7 13 9 9 2 3 3 9 3 13 2
24 3 16 9 7 9 1 9 13 2 13 3 3 0 13 9 2 15 13 9 0 1 9 13 2
7 13 3 15 13 0 9 2
29 16 3 3 9 13 2 1 3 9 13 2 13 1 0 9 9 9 9 0 2 1 3 9 13 9 3 7 9 2
5 13 3 3 9 2
14 16 3 9 13 0 9 2 9 3 13 0 9 13 2
9 3 3 13 9 0 9 7 9 2
9 3 3 15 9 13 1 9 13 2
21 9 3 0 0 13 9 2 3 3 15 0 13 3 9 16 3 9 3 9 3 2
17 2 15 3 16 3 9 13 7 9 0 2 3 9 13 13 9 2
18 3 3 15 1 9 13 2 16 9 13 2 16 15 15 9 13 13 2
25 3 16 3 1 9 13 13 9 2 9 13 2 3 1 9 13 9 2 13 0 9 15 9 13 2
10 15 3 3 15 0 9 1 9 13 2
7 9 3 9 0 13 9 2
15 3 3 2 9 9 13 0 13 0 2 15 9 0 13 2
14 15 3 13 3 7 13 9 2 9 13 0 9 0 2
9 3 3 13 9 0 0 1 9 2
24 3 16 3 13 7 13 7 13 2 9 3 13 1 3 9 13 0 13 2 1 0 3 13 2
16 3 3 13 9 13 1 13 0 2 7 9 13 13 9 0 2
18 3 16 1 9 13 7 9 13 2 13 3 3 0 7 1 9 13 2
18 3 3 15 9 13 0 9 2 13 3 13 1 9 0 7 9 9 2
17 3 16 3 1 13 13 9 0 2 3 3 15 9 13 0 9 2
7 13 3 9 0 0 13 2
8 10 3 9 0 9 13 13 2
7 3 3 0 13 13 9 2
17 16 3 15 3 13 9 0 9 2 13 1 9 7 1 9 13 2
17 15 3 3 15 3 9 0 9 9 0 13 13 0 1 9 9 2
8 2 0 3 15 13 9 0 2
8 15 3 13 9 9 0 13 2
27 2 3 16 3 1 9 13 7 9 2 13 3 0 3 2 3 3 15 9 13 13 2 9 3 13 3 2
8 15 3 3 3 9 9 13 2
13 2 3 3 3 0 0 9 13 9 9 13 0 2
35 3 16 3 0 9 1 9 13 9 2 3 3 3 9 3 13 9 13 2 15 3 3 13 13 0 9 2 9 13 1 3 9 0 13 2
36 2 3 16 3 10 9 13 2 3 3 15 0 13 9 2 7 9 7 9 2 3 3 0 9 13 9 9 1 0 2 13 3 9 1 0 2
9 15 3 13 3 3 0 1 9 2
18 3 3 13 13 9 0 1 9 13 2 9 3 9 13 9 9 0 2
12 9 3 3 13 2 9 3 0 1 9 13 2
18 15 3 3 0 1 9 13 9 9 2 1 3 9 13 0 3 9 2
15 15 3 3 9 13 13 1 9 2 13 3 9 9 0 2
9 9 3 3 13 7 13 9 9 2
19 15 3 13 0 9 13 9 2 1 3 9 13 2 13 3 1 9 9 2
15 15 3 9 0 1 9 0 9 13 2 9 3 13 9 2
27 3 15 1 9 13 2 16 1 9 13 9 9 2 15 3 0 13 9 2 1 3 15 9 13 1 9 2
10 3 1 0 0 13 2 9 9 13 2
28 2 3 3 3 9 3 13 9 13 2 13 3 1 9 3 2 13 0 9 9 2 16 3 10 0 13 9 2
15 0 13 2 3 3 9 13 13 1 9 9 0 3 9 2
7 15 3 13 9 0 9 2
14 3 15 1 0 9 3 13 2 15 13 13 3 9 2
13 3 3 3 13 3 3 13 9 0 3 3 13 2
19 9 3 3 13 2 0 3 13 9 2 0 3 0 3 2 13 3 9 2
12 3 3 13 2 16 13 3 9 7 9 3 2
6 13 3 15 13 3 2
21 16 3 1 9 9 3 13 13 9 0 13 0 2 3 3 10 3 9 9 13 2
24 13 3 15 3 9 7 9 13 2 0 3 13 1 0 9 2 13 3 1 15 13 9 0 2
11 9 3 3 13 9 9 3 9 3 13 2
7 3 3 3 13 0 9 2
5 15 15 15 13 2
10 0 3 15 13 3 3 13 13 2 2
18 3 13 2 15 3 3 0 3 13 9 2 9 3 13 1 9 0 2
22 15 3 9 0 13 15 13 2 0 1 9 0 0 9 3 13 0 2 13 3 9 2
22 9 3 3 9 0 1 9 13 7 9 0 0 3 0 9 2 0 9 0 3 13 2
10 3 3 15 13 9 0 7 9 3 2
8 15 3 3 13 1 9 13 2
9 3 13 9 2 15 3 13 9 2
22 15 3 13 13 3 0 2 3 3 9 13 0 9 2 3 13 2 13 3 0 9 2
9 15 3 1 9 13 7 9 13 2
15 15 3 9 13 0 9 9 9 0 9 2 15 0 13 2
12 3 9 0 1 9 9 13 13 2 13 13 2
5 3 3 13 13 2
7 3 9 0 13 9 9 2
13 3 3 9 0 13 2 9 3 3 13 13 9 2
10 0 3 3 9 13 13 1 0 0 2
10 15 3 3 13 13 9 0 7 9 2
14 9 3 9 13 0 2 7 3 15 0 0 13 2 2
19 3 13 2 15 3 3 0 13 7 13 13 10 9 2 16 1 9 13 2
7 3 3 9 13 9 9 2
15 3 13 2 9 3 9 9 13 2 13 3 3 0 3 2
15 15 3 9 13 0 2 15 9 0 13 2 3 1 9 2
21 1 3 13 0 9 2 9 3 1 9 13 9 0 2 7 15 13 9 0 13 2
4 3 15 13 2
15 15 3 13 15 1 9 9 3 7 9 7 9 9 2 2
24 3 13 1 9 13 0 9 2 15 3 1 9 13 9 9 2 13 1 9 0 7 9 9 2
26 9 3 3 15 9 1 13 9 2 15 3 9 13 0 7 9 2 15 3 0 9 0 3 13 13 2
10 15 3 0 9 3 13 7 9 0 2
20 1 3 3 9 13 9 3 9 3 9 1 9 0 2 16 0 13 2 0 2
23 16 15 13 13 9 9 2 3 15 0 9 1 9 13 2 0 2 0 2 9 0 13 2
7 15 3 3 3 13 3 2
15 3 15 3 13 9 9 13 2 9 13 9 0 9 13 2
28 15 3 3 3 0 13 9 0 1 9 9 3 9 0 3 9 13 2 3 3 3 3 13 2 13 0 13 2
21 16 9 13 0 2 15 3 3 13 13 9 9 0 2 3 3 9 13 0 9 2
15 3 3 3 1 9 13 9 0 2 16 3 9 9 13 2
9 1 3 9 3 7 9 13 0 2
6 3 3 3 13 9 2
12 3 3 15 0 9 13 2 7 0 9 13 2
8 3 15 3 13 2 3 13 2
6 3 3 13 9 9 2
46 15 3 1 9 13 0 3 0 9 0 1 9 13 0 1 3 9 7 9 0 2 1 3 3 1 9 13 13 9 2 1 3 9 13 2 15 15 9 0 13 3 13 1 0 9 2
26 7 15 3 3 1 9 9 0 13 1 9 2 16 3 15 9 9 2 3 3 9 13 2 13 13 2
7 0 3 3 3 3 13 2
17 3 3 9 13 9 2 15 0 9 0 13 2 9 3 13 9 2
11 7 3 3 9 13 0 0 13 3 13 2
15 9 3 15 3 3 13 3 2 16 15 0 13 7 13 2
6 3 15 15 13 9 2
10 0 3 3 13 0 7 0 9 13 2
8 15 3 13 3 3 9 3 2
10 13 16 13 7 15 0 13 9 2 2
7 15 3 13 3 9 9 2
8 3 0 3 9 13 7 13 2
33 3 3 9 13 0 9 2 1 9 13 2 1 0 9 13 2 16 3 13 2 13 3 9 9 2 0 3 15 9 9 13 2 2
7 15 3 13 13 9 9 2
3 3 13 2
17 15 3 1 13 9 2 15 15 9 13 7 13 3 9 0 13 2
5 15 3 3 13 2
9 3 3 15 13 13 1 0 0 2
6 3 3 13 0 2 2
5 3 3 15 13 2
26 2 6 6 2 3 3 3 15 0 0 13 9 0 2 15 13 9 13 15 2 16 9 0 13 0 2
24 13 3 9 9 0 2 9 2 1 9 13 2 1 0 9 13 2 0 3 15 9 9 13 2
5 3 13 10 9 2
7 15 3 3 3 0 13 2
13 9 3 13 9 2 16 3 15 13 0 1 9 2
20 9 3 9 12 13 13 2 16 3 13 2 3 3 15 0 9 9 13 2 2
11 3 13 2 15 3 13 2 13 3 9 2
10 13 3 3 13 7 3 13 0 9 2
16 13 3 3 3 7 0 13 9 9 0 2 13 3 9 13 2
7 15 3 9 0 13 15 2
6 15 3 3 0 13 2
7 6 13 13 1 9 3 2
16 15 3 3 0 0 9 13 2 15 3 15 13 7 13 13 2
22 3 3 3 3 3 3 13 13 2 3 3 3 3 13 2 16 3 15 9 0 13 2
17 9 15 13 0 2 15 3 3 0 9 13 7 13 15 15 13 2
19 3 3 3 10 9 13 7 13 2 16 15 15 13 0 1 9 13 2 2
14 15 3 13 0 9 13 1 9 0 9 2 0 13 2
29 3 3 15 13 9 2 9 9 13 0 2 9 9 2 0 2 0 3 9 9 13 2 0 1 9 13 0 9 2
11 9 3 1 0 9 13 2 9 3 9 2
16 15 3 9 13 13 7 0 13 2 7 15 13 9 0 13 2
14 15 3 15 3 13 3 3 9 7 15 0 9 13 2
10 3 15 0 13 0 2 16 3 13 2
10 15 9 2 15 9 2 15 9 13 2
15 7 3 15 9 0 2 7 15 9 13 9 13 9 9 2
8 3 3 15 3 3 0 13 2
20 3 3 3 0 7 3 0 13 2 3 3 3 0 2 3 3 3 0 13 2
8 3 3 9 13 13 3 9 2
7 7 15 13 9 0 13 2
21 3 3 15 3 0 13 2 3 3 15 3 13 9 2 3 1 9 9 0 13 2
13 2 13 9 3 3 1 9 0 2 3 1 9 2
9 3 3 13 3 0 9 1 15 2
15 15 3 15 13 13 0 9 3 2 3 9 13 1 9 2
20 9 3 3 0 13 9 2 3 3 15 15 9 13 2 13 3 15 9 13 2
24 3 16 3 15 3 13 0 9 2 3 15 1 9 13 9 0 13 2 7 15 0 9 13 2
16 3 3 3 15 3 13 9 9 0 0 2 3 3 13 13 2
7 3 3 13 13 3 9 2
26 9 3 1 9 13 2 3 3 15 15 9 9 13 2 3 3 13 13 2 7 3 13 13 9 0 2
25 3 15 3 0 9 13 13 2 15 3 9 0 0 1 9 13 13 2 3 3 0 1 9 13 2
9 15 3 1 0 3 13 13 13 2
7 3 15 13 13 9 2 2
13 9 3 13 9 0 3 0 3 7 0 9 13 2
7 7 15 13 9 0 13 2
18 2 0 3 13 7 0 15 15 13 1 0 9 2 3 16 9 13 2
34 3 3 2 3 0 13 2 13 0 9 2 16 15 3 13 9 3 0 0 9 7 9 2 15 3 1 0 9 9 3 13 7 9 2
33 15 3 13 3 9 2 3 3 15 13 3 9 3 9 2 0 2 16 3 13 13 2 7 9 13 9 0 2 9 13 9 2 2
7 15 3 13 13 0 9 2
6 15 3 0 0 13 2
15 3 3 9 0 13 13 9 13 2 16 15 9 9 13 2
21 3 3 15 1 9 13 2 3 3 13 13 1 9 0 2 7 15 0 9 13 2
17 3 15 3 3 13 13 0 13 2 16 9 13 7 0 7 0 2
16 3 3 3 0 9 13 13 13 1 9 13 9 3 9 3 2
38 15 3 3 3 0 13 13 3 3 13 2 16 3 3 0 9 13 2 15 3 3 3 13 1 9 2 0 3 15 3 13 9 3 7 9 9 13 2
20 3 15 15 3 3 3 13 2 7 1 9 13 2 15 13 13 1 0 9 2
10 3 3 15 13 9 9 2 16 13 2
15 0 3 3 9 13 0 2 3 15 0 13 9 0 9 2
9 0 3 9 13 9 13 9 2 2
10 3 13 9 13 9 2 13 3 9 2
17 13 3 3 3 0 0 9 2 13 0 9 2 13 3 0 9 2
8 3 3 9 13 2 9 13 2
6 3 3 9 0 13 2
28 3 3 9 13 2 3 10 3 3 2 16 3 13 0 15 9 9 9 0 3 13 7 15 0 9 13 2 2
11 2 13 2 3 15 0 1 9 0 13 2
17 3 9 3 9 9 0 13 3 3 2 16 3 15 15 0 13 2
9 0 3 13 16 3 9 13 2 2
12 3 13 9 13 9 0 2 13 9 1 9 2
12 15 3 13 0 1 9 9 13 9 0 9 2
27 15 3 0 3 9 13 1 9 0 3 3 13 7 13 9 0 2 9 13 2 9 3 15 0 13 2 2
7 15 3 13 13 0 9 2
9 3 3 9 13 2 16 13 0 2
17 1 3 15 0 13 2 9 0 13 2 0 16 9 13 0 9 2
19 2 3 3 15 15 3 13 2 3 3 15 13 2 16 3 3 0 13 2
18 7 15 13 9 3 9 3 13 0 9 9 9 2 15 15 9 13 2
8 3 3 15 0 13 0 9 2
51 13 3 9 0 1 0 9 2 0 3 1 9 13 9 2 1 3 9 13 15 3 13 13 9 13 2 13 3 15 9 3 0 13 2 16 3 0 0 9 13 0 3 9 7 9 2 15 1 9 13 2
25 0 3 0 9 13 2 15 15 9 9 2 3 3 15 0 13 2 9 3 0 13 7 0 9 2
6 13 15 3 9 13 2
26 15 3 13 1 9 9 1 3 9 9 2 13 9 0 7 0 9 13 2 15 3 9 13 13 9 2
7 15 3 13 13 0 9 2
13 2 3 3 3 3 15 13 2 1 9 0 13 2
6 9 3 15 0 13 2
10 2 3 3 15 0 3 3 0 13 2
11 0 15 13 2 16 9 0 13 3 13 2
18 3 3 15 13 9 2 7 0 13 1 9 9 2 1 3 0 13 2
17 3 3 15 13 0 1 9 0 2 13 13 2 16 0 9 13 2
20 3 15 3 3 13 2 16 3 15 9 13 9 9 2 15 15 9 13 2 2
8 3 3 15 13 9 13 9 2
32 13 3 9 0 1 0 9 2 0 3 1 9 13 9 2 1 3 9 0 9 0 13 9 2 13 3 15 9 3 0 13 2
11 1 3 15 0 9 0 13 9 2 0 2
11 13 3 15 9 7 0 9 2 0 0 2
6 1 3 9 13 9 2
6 15 3 3 13 13 2
11 15 3 3 1 9 0 13 1 9 9 2
32 3 15 1 9 13 0 9 9 1 0 1 9 2 3 15 9 13 0 9 2 15 15 9 3 13 9 2 15 13 0 9 2
25 15 3 3 1 9 13 13 2 3 15 9 0 13 2 0 1 9 2 0 3 0 3 2 0 2
18 9 3 3 13 3 3 7 3 2 0 7 0 2 10 0 9 13 2
12 1 3 9 9 12 13 1 0 2 9 9 2
9 10 3 9 3 13 2 0 0 2
17 15 3 13 13 0 9 2 16 13 9 3 0 9 10 0 0 2
8 15 3 0 3 7 12 13 2
13 0 3 1 9 0 13 9 2 13 9 0 0 2
17 10 3 0 13 3 9 13 9 0 9 2 16 13 9 13 9 2
7 3 3 9 13 9 0 2
5 15 3 13 13 2
11 3 9 13 9 2 9 3 15 13 9 2
9 3 3 0 1 9 0 13 9 2
16 3 9 3 9 0 13 13 1 9 2 9 3 15 13 9 2
10 10 3 13 13 9 3 0 0 9 2
5 15 3 13 9 2
11 3 3 15 0 9 13 9 3 9 3 2
15 0 3 9 13 7 13 13 2 0 3 9 9 13 13 2
23 3 15 13 3 9 13 1 0 9 9 3 9 3 2 16 3 3 13 7 13 9 9 2
31 3 13 3 13 0 9 2 13 3 13 2 9 3 13 0 2 13 3 1 9 0 0 9 2 0 0 2 0 7 0 2
15 13 3 9 16 15 3 13 2 9 3 13 1 3 13 2
10 1 3 9 13 0 9 3 9 3 2
9 9 3 0 3 0 3 13 0 2
14 15 3 9 9 13 3 13 2 16 13 9 10 0 2
11 3 3 15 0 13 9 2 16 3 13 2
18 3 13 2 3 13 9 1 9 13 3 2 16 0 9 1 9 13 2
16 3 3 15 13 9 1 9 9 1 0 2 16 9 13 2 2
18 3 13 9 3 13 9 2 13 3 13 1 9 2 3 9 13 9 2
17 3 13 12 13 7 0 13 2 13 3 13 3 7 1 9 13 2
11 13 3 3 0 13 13 9 0 0 9 2
6 15 3 9 0 13 2
17 1 3 3 9 13 0 9 2 0 3 0 13 2 13 3 13 2
16 3 0 3 9 9 13 2 3 9 13 1 9 3 3 9 2
16 3 3 0 9 9 0 13 2 7 9 13 7 0 9 9 2
6 9 3 13 0 13 2
8 3 3 15 9 3 13 0 2
6 15 3 3 15 13 2
20 0 9 9 2 0 9 9 2 0 9 0 9 13 9 3 7 0 9 9 2
16 3 3 9 0 9 12 0 9 13 2 1 3 9 0 13 2
16 15 3 15 0 1 9 9 13 2 0 9 15 15 13 0 2
19 3 15 9 15 13 3 13 3 2 7 15 9 10 0 3 13 13 2 2
21 3 16 13 7 13 9 9 2 3 15 13 13 9 2 15 3 13 2 9 0 2
15 15 3 13 2 13 3 9 2 7 15 13 9 0 13 2
8 13 3 0 13 9 1 9 2
10 13 15 2 16 3 3 13 0 13 2
6 1 0 3 13 2 2
16 15 3 3 13 9 1 9 13 2 13 1 9 0 0 13 2
27 15 3 3 13 13 7 0 13 2 7 15 13 9 1 9 13 2 15 9 13 9 2 16 9 3 13 2
17 15 3 3 13 9 0 15 9 9 1 9 13 2 9 3 13 2
18 3 15 3 3 13 2 0 3 9 3 0 2 15 3 3 2 13 2
31 3 3 3 0 0 3 9 13 2 3 13 2 3 3 16 3 9 7 9 3 13 9 2 3 3 13 7 15 13 0 2
17 3 3 3 15 3 0 13 2 13 3 9 13 13 1 0 9 2
7 3 15 9 9 13 13 2
8 1 3 15 13 7 13 9 2
9 3 15 0 13 3 3 13 2 2
8 15 3 3 13 0 0 9 2
14 3 15 3 3 13 2 7 1 9 2 16 13 9 2
15 9 3 15 13 3 2 16 3 15 13 10 0 9 13 2
13 3 3 3 2 3 3 3 13 2 3 15 13 2
15 0 3 15 0 1 9 9 13 2 15 9 13 0 13 2
18 13 3 9 0 9 2 0 3 9 2 9 3 9 0 2 15 13 2
9 3 3 3 15 0 13 3 13 2
7 15 0 9 13 3 9 2
15 3 0 13 2 7 0 3 13 2 3 3 15 0 13 2
14 3 3 9 1 9 0 13 2 16 15 13 0 9 2
37 15 16 13 9 9 0 2 7 15 13 13 1 9 3 15 9 9 0 0 2 9 7 9 0 2 15 3 15 0 13 9 3 0 7 15 9 2
10 15 3 13 1 9 9 1 9 0 2
18 15 3 9 0 3 13 13 2 16 1 9 13 0 1 9 9 0 2
20 3 3 3 0 3 13 2 7 3 13 7 3 13 7 3 15 13 9 9 2
6 0 3 1 9 13 2
8 3 3 15 9 13 1 9 2
4 15 13 13 2
11 3 3 3 15 15 0 13 3 13 2 2
24 13 3 3 15 1 9 7 9 7 9 0 9 1 13 2 13 0 2 0 3 1 9 13 2
23 3 3 3 3 1 9 0 3 15 13 13 0 9 9 2 0 3 3 0 9 9 13 2
36 15 3 0 13 9 9 2 7 15 0 0 13 9 9 2 15 15 9 13 13 15 3 1 9 9 7 13 9 9 3 9 3 7 9 0 2
12 3 3 3 15 9 13 9 13 1 9 9 2
17 13 3 9 0 9 1 0 9 2 16 3 0 13 3 3 0 2
14 3 3 3 0 13 7 3 9 3 15 13 13 13 2
8 3 3 15 9 13 3 0 2
13 3 3 3 9 15 9 3 13 7 9 7 9 2
32 16 13 3 9 9 2 0 0 13 2 3 3 15 9 13 9 0 2 7 0 0 13 9 13 9 0 15 3 15 13 9 2
5 0 13 1 9 2
12 3 15 15 0 13 15 3 9 1 9 13 2
8 0 3 3 0 9 13 9 2
23 16 3 3 9 13 9 0 3 9 13 7 0 9 9 1 0 2 7 15 3 13 0 2
9 15 13 0 2 0 3 3 13 2
16 3 3 9 13 2 7 3 3 0 3 0 3 1 9 13 2
31 2 3 16 3 10 3 0 9 0 9 13 2 15 0 9 1 9 13 2 3 3 15 13 7 0 9 9 13 1 9 2
13 3 3 15 9 13 13 2 0 3 13 9 9 2
23 3 3 0 13 9 0 2 10 0 3 9 9 13 13 3 1 9 2 9 3 13 0 2
8 3 15 0 0 13 9 9 2
12 9 3 0 13 13 9 0 3 9 7 9 2
15 3 3 3 15 9 13 13 2 9 3 13 1 0 9 2
9 12 9 13 2 3 3 13 9 2
8 3 3 3 0 9 9 13 2
13 3 15 9 0 13 9 3 13 0 3 9 13 2
22 3 3 15 3 15 9 13 2 7 0 7 0 13 2 15 3 9 3 9 3 13 2
23 3 3 3 3 15 13 9 9 3 1 9 13 7 9 13 2 9 3 1 9 13 13 2
7 3 3 1 9 13 9 2
9 15 3 9 13 1 9 13 13 2
12 13 3 0 9 0 3 7 9 9 3 9 2
17 1 3 9 0 9 0 9 0 13 2 3 3 15 13 13 0 2
6 1 3 0 3 13 2
17 3 15 0 3 13 0 9 2 15 3 13 0 2 15 13 9 2
11 3 15 9 3 13 9 7 13 9 13 2
16 15 13 7 15 13 2 1 9 3 15 13 13 3 9 13 2
15 2 3 3 0 13 3 2 0 3 13 9 1 0 9 2
4 13 3 0 2
8 3 1 0 13 0 1 9 2
41 3 16 3 9 3 7 9 13 3 13 9 7 13 9 2 1 9 15 1 9 13 0 9 13 2 16 15 1 9 13 2 3 3 15 16 13 7 0 9 13 2
10 15 13 1 9 2 13 3 2 9 2
12 15 3 13 9 9 0 0 2 0 1 9 2
6 9 3 15 13 9 2
35 3 16 3 9 3 13 2 3 3 15 0 13 9 2 7 9 7 9 2 3 3 0 9 13 9 9 1 0 2 13 3 9 1 0 2
13 15 3 13 0 9 13 9 2 1 3 9 13 2
6 13 3 1 9 0 2
10 15 3 9 0 1 9 0 9 13 2
5 9 3 13 9 2
23 3 15 9 0 2 13 3 9 9 2 9 0 9 0 1 9 13 2 16 3 9 13 2
7 15 3 13 13 0 9 2
15 3 13 2 0 3 15 9 0 9 9 13 0 9 13 2
21 15 3 0 9 13 9 7 9 13 13 1 9 2 9 13 2 16 13 9 9 2
10 1 3 15 9 3 9 3 9 13 2
6 2 3 9 15 13 2
10 3 3 1 0 9 0 3 3 13 2
8 0 15 1 9 9 13 9 2
31 15 3 1 9 13 13 2 16 9 1 9 0 9 9 13 2 16 13 9 1 0 9 3 3 13 2 7 3 7 3 2
26 13 3 1 15 0 2 13 1 9 2 9 13 7 0 13 9 2 15 3 15 13 0 1 0 9 2
5 3 15 3 13 2
10 13 3 13 9 9 9 1 9 0 2
10 3 15 3 15 13 13 9 9 3 2
17 15 3 0 9 13 9 1 15 2 16 3 3 9 1 9 13 2
14 3 16 9 0 13 0 9 2 3 0 9 15 13 2
7 0 3 9 0 9 13 2
21 3 15 3 13 0 1 9 9 0 3 2 0 3 13 3 1 9 9 9 13 2
9 3 15 9 3 13 9 0 3 2
28 9 3 1 9 13 2 0 9 13 13 9 9 2 3 3 9 13 0 13 2 3 3 3 3 13 1 0 2
13 3 13 2 3 3 9 13 0 9 2 13 13 2
6 15 3 0 13 13 2
19 3 3 3 15 13 0 13 13 3 2 15 3 3 3 13 9 1 0 2
15 15 3 13 9 0 3 2 7 15 9 13 13 9 13 2
24 3 3 15 9 3 13 9 2 7 3 3 0 9 0 9 13 3 3 3 15 3 9 13 2
19 3 3 3 13 2 16 3 3 15 0 9 13 13 2 16 9 3 13 2
22 3 15 3 10 0 13 13 2 7 15 13 3 13 9 2 7 15 13 9 0 13 2
33 3 15 3 0 13 13 7 13 2 1 15 3 15 0 9 13 9 2 15 3 9 13 2 0 1 9 13 2 13 0 1 9 2
5 15 3 15 13 2
18 7 13 13 7 1 9 7 1 9 2 0 9 13 2 1 0 9 2
19 3 3 3 15 15 13 3 3 13 2 7 9 0 13 0 3 13 2 2
6 3 3 3 9 13 2
27 16 3 3 13 9 0 1 15 9 2 13 15 9 3 9 3 9 13 3 13 2 3 15 0 13 9 2
25 16 3 3 3 13 9 0 7 13 2 9 13 13 0 1 9 2 16 3 0 9 13 13 2 2
7 15 3 13 13 0 9 2
14 0 15 3 9 13 2 16 1 9 0 13 9 2 2
17 3 15 3 0 1 0 13 2 0 3 9 3 7 9 13 9 2
11 2 13 9 10 0 2 16 9 13 0 2
15 3 3 0 13 2 15 3 9 3 13 13 9 1 0 2
8 0 3 0 9 0 13 2 2
16 3 3 13 13 9 0 9 2 15 3 9 13 3 9 0 2
7 15 3 3 13 1 9 2
7 3 3 9 13 3 0 2
5 9 3 13 0 2
10 13 3 13 9 9 2 15 13 13 2
5 15 3 13 9 2
5 3 3 15 13 2
6 1 3 9 13 13 2
6 1 3 9 0 13 2
8 7 15 3 3 0 13 13 2
13 9 3 9 0 13 0 9 2 13 3 9 9 2
7 7 15 13 13 0 9 2
5 13 3 0 2 2
18 13 3 3 9 13 9 0 2 13 3 0 9 9 0 1 9 13 2
7 15 3 13 0 1 9 2
21 9 3 15 13 9 2 15 3 9 0 13 0 13 9 2 1 9 7 9 9 2
9 1 3 3 15 9 13 9 0 2
9 15 3 1 9 0 13 9 13 2
25 3 16 9 7 9 1 9 13 2 9 3 15 13 9 2 15 3 1 9 9 7 9 13 13 2
20 9 3 3 13 0 0 2 13 3 3 9 0 2 7 13 9 0 3 0 2
26 15 3 9 13 2 9 13 2 16 3 15 13 9 13 2 7 15 9 0 13 2 16 15 13 3 2
15 2 13 3 2 9 7 0 0 9 2 13 15 9 13 2
32 9 3 13 0 2 15 3 13 9 3 3 13 7 3 0 13 2 7 3 13 13 2 7 15 9 13 15 3 3 0 0 2
10 3 16 3 10 0 13 2 3 13 2
17 6 3 13 9 3 15 0 13 2 3 16 1 9 9 13 13 2
15 13 3 9 3 7 9 9 2 15 3 1 0 13 15 2
4 0 3 13 2
29 3 16 3 3 13 1 9 0 3 9 2 15 3 1 9 1 9 0 2 1 9 7 9 2 1 9 13 13 2
10 9 3 3 13 0 9 13 2 0 2
16 3 0 0 9 13 7 9 2 13 3 0 2 9 13 9 2
24 3 15 9 3 13 9 13 9 2 16 3 13 13 3 2 7 13 9 0 13 7 9 0 2
22 3 16 3 3 9 13 2 1 3 9 13 2 3 3 15 9 13 3 13 9 13 2
6 15 3 3 3 13 2
5 3 3 13 9 2
7 1 15 13 9 9 13 2
7 3 3 3 0 13 2 2
20 2 3 13 2 15 3 3 9 13 15 1 9 2 0 0 13 13 7 13 2
9 13 3 0 9 15 1 9 13 2
12 2 13 3 2 16 15 15 0 0 13 2 2
11 2 13 3 1 9 9 13 13 3 9 2
6 0 15 0 13 9 2
6 3 3 9 1 13 2
13 15 3 1 9 0 13 3 2 13 3 0 9 2
9 3 3 13 9 3 15 0 13 2
16 13 3 15 9 1 9 9 2 0 2 9 7 9 9 0 2
10 3 3 15 13 0 9 9 13 2 2
18 3 3 3 9 13 3 3 15 0 2 15 13 9 0 13 2 3 2
8 3 3 3 10 0 9 13 2
26 3 16 13 9 0 9 2 0 15 9 3 9 3 9 13 2 13 3 3 15 9 9 3 13 2 2
4 3 9 13 2
21 1 3 9 13 0 0 7 0 2 15 15 13 9 2 13 16 15 9 0 13 2
12 13 3 9 2 16 3 15 9 13 3 13 2
17 13 3 13 13 3 3 9 0 9 1 0 13 2 9 1 9 2
17 9 3 3 9 13 0 2 7 1 9 9 1 0 9 9 13 2
7 3 3 13 13 0 9 2
15 3 13 0 9 0 9 13 2 16 3 3 0 9 13 2
11 3 3 3 9 3 9 3 13 9 13 2
10 15 3 13 0 9 9 7 13 9 2
10 3 3 15 15 3 9 1 9 13 2
8 13 3 0 9 1 9 9 2
21 0 13 9 13 15 3 13 2 9 3 0 7 0 0 3 13 13 3 3 13 2
24 3 15 3 13 0 13 0 9 15 15 15 0 13 13 2 1 15 3 15 13 9 0 9 2
12 0 3 15 15 9 13 2 15 3 13 9 2
13 9 15 3 9 13 1 9 9 3 9 3 0 2
6 3 15 3 3 13 2
13 3 3 15 9 13 9 9 2 15 3 9 13 2
12 3 3 9 13 0 9 2 9 3 3 13 2
14 13 3 15 9 3 0 15 15 15 13 3 13 3 2
33 3 16 0 9 9 13 2 9 3 1 9 13 7 0 9 2 0 3 0 9 13 2 15 15 9 9 2 3 3 15 0 13 2
5 3 3 9 13 2
20 15 3 13 9 1 9 13 9 9 2 16 15 0 13 7 1 9 13 2 2
27 15 3 3 3 13 13 1 0 9 2 3 15 9 1 0 9 13 3 9 13 2 7 15 1 9 13 2
5 3 3 13 9 2
9 3 13 2 3 3 0 13 9 2
9 3 3 15 9 13 3 13 2 2
8 15 3 13 3 9 0 9 2
17 13 3 3 0 9 9 2 15 3 3 3 13 2 3 3 13 2
17 0 3 0 13 2 15 3 3 13 13 9 13 7 15 13 13 2
9 13 9 13 13 2 13 3 13 2
27 3 13 1 15 3 9 13 0 13 0 2 15 3 9 13 2 13 3 9 9 1 9 13 3 3 13 2
25 16 3 13 13 1 9 7 0 9 2 16 15 0 13 2 13 3 15 9 2 9 3 9 13 2
8 15 3 3 9 13 3 13 2
10 3 3 3 9 13 13 1 9 0 2
17 7 9 0 13 0 13 2 7 15 15 1 9 9 0 13 2 2
11 15 9 13 13 9 0 9 13 3 9 2
7 15 3 3 3 13 13 2
18 0 3 1 9 13 0 2 3 0 2 1 15 3 9 13 7 9 2
15 9 3 13 9 2 3 13 15 9 0 2 15 13 0 2
5 13 3 0 0 2
11 13 3 13 3 1 9 2 16 13 9 2
6 15 3 13 0 9 2
17 9 3 2 0 1 0 9 9 13 2 13 15 0 7 0 13 2
5 13 15 9 13 2
15 0 3 13 0 2 9 3 1 9 13 2 9 3 9 2
7 15 3 13 15 13 2 2
10 3 13 1 9 13 9 0 9 9 2
16 9 3 13 0 9 13 1 9 2 9 3 13 1 3 13 2
9 3 3 0 1 9 13 1 9 2
14 15 3 15 13 13 9 0 7 0 1 0 9 2 2
11 3 13 1 9 13 2 15 3 13 13 2
16 7 15 3 1 9 13 9 9 13 2 7 0 0 13 9 2
9 15 3 13 1 9 9 0 9 2
10 13 3 3 3 1 9 3 9 3 2
15 9 3 0 9 13 13 0 0 2 1 0 9 2 13 2
6 1 3 0 13 9 2
7 9 3 0 9 13 13 2
6 13 3 9 9 0 2
9 15 3 1 9 0 13 9 13 2
23 15 3 1 9 13 0 9 2 9 13 1 9 9 0 2 1 9 0 2 16 13 13 2
9 13 3 9 1 2 13 3 13 2
17 3 3 15 3 9 7 0 13 2 16 1 9 13 9 0 2 2
8 15 3 3 9 13 9 13 2
29 7 3 15 3 13 3 2 13 9 1 9 2 13 16 1 15 13 9 0 13 2 3 13 9 0 7 0 2 2
12 15 3 13 13 2 7 0 1 9 9 13 2
7 15 3 9 9 13 9 2
15 3 13 2 13 3 0 9 2 16 15 1 9 13 13 2
8 15 3 9 0 13 13 9 2
4 2 13 15 2
14 3 15 13 2 3 1 9 0 13 7 3 13 13 2
8 15 3 3 9 13 9 13 2
10 3 3 15 3 3 9 3 13 2 2
7 13 7 1 9 9 13 2
10 15 3 3 3 13 3 1 9 13 2
8 15 3 0 13 9 3 13 2
8 13 3 9 13 3 0 9 2
11 3 3 9 13 15 3 15 1 0 13 2
24 16 3 0 13 0 9 2 9 3 13 1 3 9 0 13 2 1 3 13 9 7 9 0 2
10 13 3 13 2 15 3 3 0 13 2
8 3 3 3 13 9 0 9 2
7 7 3 9 13 9 9 2
14 9 3 3 13 13 1 9 9 2 3 3 9 13 2
8 15 3 9 3 3 9 13 2
18 2 3 13 2 9 3 3 0 13 9 2 16 15 1 9 13 13 2
8 3 3 15 13 13 0 13 2
7 7 15 13 9 0 13 2
17 2 9 3 13 13 3 0 9 2 16 15 3 13 13 3 9 2
11 3 3 15 15 13 1 9 7 1 9 2
23 0 0 9 0 2 3 15 13 2 3 0 13 3 13 2 3 3 15 13 3 13 0 2
6 3 3 13 3 2 2
17 3 3 13 13 9 9 3 0 1 9 2 3 3 3 9 13 2
6 9 3 9 13 13 2
23 2 3 13 2 15 3 3 15 3 3 13 7 13 2 3 3 3 13 7 1 9 13 2
16 3 3 15 3 15 13 7 13 2 13 3 9 9 1 0 2
26 3 3 3 0 9 13 2 9 13 9 3 0 2 0 13 2 15 15 9 0 0 1 9 13 9 2
27 3 15 3 13 9 7 13 9 0 1 9 1 9 7 13 9 0 0 9 2 9 3 9 13 1 9 2
23 9 3 13 9 0 2 3 9 0 9 2 15 1 9 13 9 3 0 7 9 0 9 2
14 3 3 13 9 9 2 7 13 1 9 0 1 9 2
8 9 3 13 9 3 9 3 2
15 3 3 3 9 0 13 9 9 1 0 2 16 0 13 2
14 3 0 9 9 9 13 9 3 0 2 16 13 9 2
17 15 3 3 9 13 2 9 3 9 13 2 15 3 9 1 13 2
18 15 3 13 13 13 3 0 1 9 0 2 7 15 13 9 0 13 2
5 15 3 13 9 2
8 15 3 3 9 13 9 13 2
15 1 9 9 13 2 9 3 15 13 9 2 16 3 13 2
7 3 3 3 13 0 9 2
15 3 3 9 3 13 7 9 0 13 13 9 3 13 2 2
7 15 3 3 13 9 0 2
16 15 13 9 7 9 0 13 2 16 3 15 9 1 9 13 2
14 3 15 9 13 2 16 15 13 13 2 16 15 13 2
5 13 3 13 2 2
8 15 3 3 9 13 9 13 2
14 2 3 3 3 15 13 3 13 9 0 2 7 13 2
9 3 3 13 2 0 3 13 2 2
17 3 3 13 15 13 0 9 2 7 15 3 1 9 13 9 0 2
8 1 3 3 0 9 13 0 2
14 1 9 3 3 3 13 2 1 3 15 0 13 9 2
5 15 3 0 13 2
8 9 3 9 13 13 9 13 2
5 15 3 3 13 2
21 9 3 0 0 1 9 13 13 2 1 3 9 13 2 13 3 9 0 0 9 2
22 15 3 0 9 13 0 9 2 0 13 1 9 2 16 0 9 13 13 9 0 9 2
8 13 3 1 9 7 9 0 2
8 13 3 9 13 3 0 9 2
16 3 3 3 9 13 0 2 13 7 3 9 13 7 3 13 2
7 1 3 15 13 9 0 2
33 3 16 9 7 9 1 9 13 2 15 3 9 13 2 9 13 2 7 15 3 3 13 13 3 13 3 1 9 2 7 13 3 2
14 3 1 9 13 13 13 2 16 3 15 13 7 9 2
16 3 15 3 3 13 7 3 9 0 13 15 3 15 3 13 2
15 1 3 9 0 9 13 2 16 3 15 9 7 9 13 2
26 7 3 13 1 9 9 0 9 13 9 9 2 7 3 9 0 13 2 16 15 9 13 9 0 13 2
9 3 3 3 13 1 15 15 13 2
12 1 3 15 13 2 15 3 13 7 15 13 2
8 3 15 3 3 13 3 13 2
28 3 3 15 13 9 0 2 7 0 2 9 3 13 7 9 2 3 3 0 9 7 0 9 2 15 15 13 2
10 0 3 9 9 7 9 7 9 13 2
3 3 13 2
8 15 3 13 3 0 0 9 2
8 9 3 3 13 0 0 9 2
18 3 1 0 9 0 9 13 9 2 15 15 13 9 7 9 7 9 2
17 9 3 3 13 2 9 3 13 3 9 1 9 13 0 1 9 2
21 3 3 9 13 13 0 3 9 0 2 15 15 3 13 13 7 1 0 9 13 2
11 15 3 13 2 0 3 15 15 0 13 2
6 13 3 15 3 3 2
6 3 3 3 0 13 2
10 3 15 0 9 13 0 9 15 13 2
9 15 13 3 13 3 7 0 13 2
30 0 3 9 13 9 9 13 7 0 13 7 13 13 3 2 3 3 3 15 13 3 2 0 3 9 3 9 13 2 2
7 15 3 13 13 0 9 2
9 13 3 13 2 13 3 13 13 2
11 3 3 15 15 13 2 16 9 2 13 2
12 10 3 0 15 9 7 9 13 2 13 13 2
10 1 3 9 13 13 1 9 0 13 2
15 15 3 1 9 13 3 13 3 9 0 13 0 2 13 2
18 1 3 3 3 9 13 9 2 15 15 3 3 0 13 7 0 13 2
10 0 3 15 13 15 15 13 7 13 2
35 2 9 15 9 13 2 16 3 13 2 9 1 2 3 9 9 2 3 15 0 3 0 2 7 0 3 2 0 2 0 2 0 2 0 2
18 9 3 3 3 9 13 2 3 3 15 0 9 1 0 13 0 9 2
19 3 16 13 9 1 9 9 2 13 0 9 9 1 0 0 9 13 13 2
10 3 12 9 2 3 3 15 0 13 2
18 13 3 9 0 9 9 1 9 2 0 3 0 3 7 0 9 13 2
7 15 3 3 9 0 13 2
24 13 15 0 13 0 1 9 9 7 9 2 15 3 9 13 0 9 2 3 15 3 0 13 2
9 13 3 3 15 13 7 3 13 2
9 15 3 3 3 9 13 0 9 2
16 2 1 3 9 0 13 13 2 9 3 13 9 15 3 0 2
19 3 15 13 9 9 9 3 13 2 13 3 3 3 13 15 9 1 9 2
7 15 3 0 9 13 2 2
11 2 15 3 3 13 9 2 15 13 3 2
22 2 3 3 3 3 3 3 1 15 3 13 2 16 13 9 7 9 0 9 0 3 2
8 3 3 3 13 7 0 13 2
19 3 16 3 13 3 13 3 10 9 2 15 3 3 13 9 7 13 9 2
22 2 13 3 2 3 15 15 13 9 0 9 2 13 7 1 9 2 7 3 1 9 2
11 3 13 1 9 9 2 13 3 9 0 2
17 3 16 3 3 9 0 9 13 2 9 15 3 3 1 9 13 2
10 13 3 3 9 2 15 3 0 13 2
10 3 3 3 0 9 15 13 3 13 2
16 9 3 9 0 1 9 13 2 0 3 0 2 3 13 3 2
20 15 3 13 1 9 2 15 3 15 0 9 13 2 3 13 1 0 9 2 2
26 2 15 3 3 3 13 13 1 9 0 2 15 3 9 0 1 15 3 13 1 9 0 9 0 13 2
19 3 16 3 0 9 13 15 13 2 3 3 3 9 13 2 15 13 9 2
16 13 9 9 0 1 9 9 0 9 13 2 1 3 9 13 2
6 15 3 15 13 9 2
18 3 3 15 13 0 1 9 13 2 15 3 15 9 13 9 13 3 2
16 13 3 1 9 7 9 7 9 9 9 2 15 15 9 13 2
21 15 3 3 1 9 13 2 9 3 9 2 15 3 3 12 9 13 1 9 13 2
5 3 15 13 9 2
9 13 3 9 2 13 3 0 9 2
17 15 3 1 9 0 13 3 13 2 3 3 9 9 13 0 9 2
11 15 3 3 13 13 0 9 2 15 13 2
6 1 3 9 9 13 2
9 3 3 3 13 9 3 7 9 2
26 3 16 3 0 9 1 9 13 9 2 10 3 3 9 13 9 0 2 9 3 13 13 3 0 9 2
10 7 15 3 9 7 9 9 13 13 2
6 3 15 13 13 9 2
17 15 3 9 13 13 9 3 7 9 2 3 15 9 13 9 0 2
9 3 15 3 9 15 13 9 2 2
8 15 3 3 0 9 13 9 2
35 3 3 3 15 3 1 3 0 0 13 9 2 16 9 9 13 0 13 0 2 15 3 15 13 9 3 9 3 3 2 13 3 0 9 2
12 3 15 3 0 9 1 9 13 3 13 2 2
18 3 15 3 0 1 0 13 2 13 3 3 0 1 9 2 7 3 2
6 3 3 9 13 0 2
10 1 3 9 13 2 1 3 0 13 2
17 1 3 3 0 13 1 9 9 2 9 3 13 13 3 0 9 2
16 3 16 9 7 9 1 9 13 2 15 3 9 13 13 9 2
16 2 15 3 3 3 13 9 0 2 3 15 9 13 7 9 2
9 0 3 1 9 13 0 9 13 2
7 15 3 3 13 9 0 2
9 3 3 0 9 13 7 0 9 2
8 15 3 3 9 13 9 13 2
12 2 3 3 15 3 15 3 3 3 13 13 2
17 3 3 3 15 3 9 1 9 13 2 7 1 15 9 9 13 2
16 3 3 0 0 9 13 3 3 9 0 13 7 9 9 13 2
20 3 15 3 9 13 0 2 9 13 2 16 3 15 1 9 13 0 9 2 2
19 1 3 9 13 9 13 2 1 3 9 13 3 1 9 3 7 0 9 2
17 0 3 3 13 9 0 0 1 9 9 2 3 15 0 3 2 2
8 15 3 3 9 13 9 13 2
20 3 3 3 13 9 3 0 3 9 1 15 2 16 3 15 15 13 13 2 2
20 3 3 15 10 9 13 1 9 0 3 13 7 13 2 1 15 3 13 2 2
8 15 3 3 9 0 9 13 2
17 3 13 1 9 13 2 13 3 9 0 3 13 1 3 0 13 2
9 15 3 3 13 7 1 9 13 2
21 9 3 1 9 13 0 9 2 13 3 0 9 2 0 0 9 2 9 1 9 2
5 15 3 0 13 2
28 15 3 3 13 9 13 2 16 13 9 2 3 15 13 9 3 0 2 15 9 0 13 13 2 9 0 13 2
11 9 3 13 9 0 2 3 3 13 13 2
14 13 3 0 9 13 3 9 2 1 3 9 13 9 2
8 3 3 3 9 9 0 13 2
7 9 3 1 9 13 2 2
14 3 3 0 13 9 2 16 15 0 9 13 1 9 2
20 13 3 13 9 2 1 3 3 15 9 13 9 2 15 13 2 13 0 9 2
19 15 3 0 13 9 2 13 3 15 9 3 7 0 9 0 9 3 0 2
6 0 3 15 13 9 2
7 7 3 13 9 0 13 2
13 3 15 3 15 3 13 13 2 16 13 9 3 2
14 3 3 3 15 3 9 13 3 3 9 2 7 13 2
14 3 3 3 15 13 9 2 9 9 13 0 9 2 2
8 15 3 3 9 13 3 13 2
12 2 3 3 0 3 13 13 9 0 1 9 2
13 0 3 15 3 13 9 3 7 9 9 13 2 2
8 3 3 13 15 13 0 9 2
10 3 15 3 3 13 7 13 0 9 2
10 15 3 3 3 13 9 9 1 0 2
11 3 13 2 15 3 3 13 1 3 13 2
8 13 1 0 9 7 9 3 2
7 3 13 3 9 0 9 2
31 15 3 3 9 9 13 9 0 2 15 3 10 0 13 13 2 9 3 3 13 1 9 2 1 3 3 9 13 0 9 2
9 15 3 1 9 0 13 9 13 2
16 3 16 9 7 9 1 9 13 2 3 3 9 13 0 9 2
8 3 3 15 9 13 1 9 2
4 15 13 13 2
11 3 3 3 15 15 0 13 3 13 2 2
16 1 3 9 9 13 0 2 13 3 0 9 1 9 13 13 2
8 3 3 15 13 15 3 9 2
17 3 3 9 9 1 9 13 13 0 1 9 2 15 3 15 13 2
4 13 16 13 2
7 9 3 15 13 13 2 2
8 15 3 3 9 13 3 13 2
9 3 3 3 10 9 15 13 9 2
17 0 3 0 13 7 3 3 9 13 9 13 2 16 15 0 13 2
10 16 3 13 2 15 13 1 9 13 2
18 9 3 3 15 13 7 9 0 13 2 16 3 3 15 13 7 9 2
12 3 3 3 3 15 15 3 1 9 13 13 2
6 3 3 0 9 13 2
8 15 3 3 13 0 0 9 2
35 13 15 7 0 13 2 7 15 3 9 13 1 9 2 13 9 9 2 7 15 9 13 2 15 3 9 13 13 2 3 16 0 9 13 2
23 3 3 1 15 9 13 0 9 2 16 3 15 0 0 0 13 2 13 1 9 9 9 2
8 15 3 3 9 13 3 13 2
26 3 3 15 15 0 9 13 13 2 3 3 9 13 2 15 3 9 13 13 2 3 16 0 9 13 2
7 3 3 0 9 13 9 2
13 0 9 9 9 13 2 0 3 3 9 9 13 2
12 3 9 0 15 1 9 13 13 3 3 13 2
9 3 3 0 3 0 13 1 9 2
7 15 3 13 13 9 0 2
7 3 3 15 13 3 0 2
10 3 3 3 3 0 9 1 9 13 2
13 3 15 3 13 2 15 3 3 13 2 0 13 2
8 10 3 0 3 15 0 13 2
7 0 3 15 0 13 2 2
5 2 13 2 13 2
6 15 3 3 13 13 2
8 15 3 3 9 13 3 13 2
11 2 0 2 7 3 15 13 2 13 3 2
16 16 3 3 13 0 0 9 2 0 3 10 9 13 0 9 2
15 3 15 3 13 3 13 2 3 3 1 9 13 1 0 2
11 3 1 9 13 0 9 13 16 0 3 2
7 0 3 3 13 9 2 2
6 13 3 7 13 9 2
13 15 3 13 9 9 2 13 3 1 9 3 13 2
13 9 3 13 9 0 3 0 3 7 0 9 13 2
8 13 3 1 0 9 9 13 2
7 15 3 3 1 9 13 2
19 13 3 0 9 2 1 3 13 9 1 0 9 9 2 13 3 1 0 2
5 15 3 13 9 2
22 3 3 0 9 9 13 3 3 13 2 16 3 9 9 7 9 13 13 1 9 0 2
12 3 3 15 0 0 1 15 13 13 13 2 2
7 13 3 0 9 13 9 2
17 9 3 15 0 0 7 9 13 1 9 2 9 3 13 7 9 2
16 3 3 0 13 2 9 3 13 2 0 3 13 9 1 9 2
8 15 3 3 3 13 3 13 2
6 3 9 13 1 9 2
23 13 3 15 0 9 2 13 3 3 13 9 2 16 9 13 2 7 15 13 9 0 13 2
11 3 3 15 9 13 2 15 9 0 13 2
14 3 13 2 16 15 13 13 0 7 0 9 2 13 2
4 13 3 15 2
8 15 3 13 3 9 0 9 2
7 2 3 15 3 9 13 2
5 15 15 0 13 2
18 3 9 0 13 2 15 1 15 13 13 9 0 2 9 13 9 2 2
13 3 3 13 9 13 2 1 3 9 9 13 3 2
6 3 3 13 3 3 2
25 3 3 3 3 0 9 15 13 0 0 3 9 2 16 3 9 0 13 3 13 13 0 7 9 2
10 3 3 3 0 13 9 7 0 13 2
11 3 3 9 13 2 15 9 0 13 2 2
7 15 3 13 13 9 9 2
29 3 3 3 3 3 0 13 3 9 2 7 15 15 15 2 13 0 2 0 3 13 2 13 0 9 1 0 9 2
25 3 3 13 1 3 13 2 9 3 13 9 0 13 2 9 13 2 0 3 15 1 9 13 9 2
10 3 3 15 3 0 1 9 9 13 2
16 7 3 3 13 13 9 9 2 16 3 9 13 0 9 3 2
4 15 13 13 2
11 3 3 3 15 15 0 13 3 13 2 2
8 15 3 3 13 9 0 9 2
16 9 15 13 0 2 15 3 3 0 9 13 2 15 15 13 2
9 3 15 3 1 9 9 9 13 2
14 3 3 3 13 9 9 2 16 3 0 9 3 13 2
17 3 3 15 9 13 13 2 16 13 0 3 7 15 15 9 13 2
24 3 3 0 1 9 0 13 13 2 7 3 15 13 13 0 1 0 2 7 3 13 0 2 2
8 15 3 3 9 13 3 13 2
5 3 3 0 13 2
4 9 15 13 2
11 3 3 3 13 9 12 0 7 0 13 2
6 3 3 13 3 9 2
14 1 3 9 12 7 12 9 13 2 12 3 9 13 2
16 15 16 3 0 13 3 13 2 3 0 7 0 9 13 13 2
21 3 15 3 2 16 13 15 9 13 2 13 2 15 3 15 15 13 0 9 2 2
8 15 3 3 13 0 0 9 2
12 2 3 15 13 2 15 3 13 7 15 13 2
18 7 13 7 3 15 9 1 9 9 13 2 7 15 0 9 13 2 2
8 15 3 3 9 13 3 13 2
12 15 3 3 0 9 3 13 7 0 9 2 2
8 15 3 3 13 9 0 9 2
24 2 3 3 3 0 3 0 9 1 13 9 0 2 3 9 7 15 1 9 0 9 13 9 2
15 3 15 3 3 13 1 9 13 3 2 7 9 0 13 2
14 3 15 1 9 9 0 13 2 0 0 0 7 9 2
5 15 3 13 13 2
11 3 3 3 13 13 9 2 0 9 13 2
7 15 3 3 3 15 13 2
7 3 3 15 13 0 9 2
12 0 3 15 13 2 15 3 1 9 13 0 2
34 3 3 0 1 9 13 9 2 13 3 15 15 9 2 15 3 3 13 0 15 1 9 0 9 13 1 9 0 9 13 13 0 3 2
12 3 9 0 9 13 2 16 3 15 13 13 2
24 2 1 9 13 2 16 3 15 13 0 3 3 13 13 9 2 7 13 2 0 9 13 9 2
7 0 3 13 9 9 2 2
21 2 15 3 0 12 9 7 12 9 13 7 0 9 9 13 2 16 3 13 13 2
11 15 3 3 3 9 9 13 7 9 9 2
12 0 3 15 13 2 15 3 1 9 13 0 2
42 16 0 3 0 13 7 9 0 2 3 15 3 9 13 3 13 2 3 3 9 13 15 3 3 9 3 15 9 3 0 9 2 7 0 15 3 15 3 9 13 9 2
9 3 3 3 15 9 3 15 13 2
11 3 3 3 15 9 15 13 13 15 0 2
5 15 3 13 13 2
10 3 3 3 13 0 13 2 9 13 2
13 15 3 1 9 0 9 13 0 3 3 1 9 2
18 3 3 3 15 9 15 13 13 2 15 3 15 13 7 15 9 13 2
27 9 3 3 3 15 3 1 9 13 15 13 2 7 0 0 13 2 16 0 3 15 13 9 9 0 2 2
33 15 3 16 3 9 0 1 13 2 9 3 15 3 0 1 9 13 2 9 3 15 13 0 9 2 3 3 1 9 13 0 9 2
17 3 16 3 3 13 9 0 9 2 9 3 3 0 1 9 13 2
14 9 3 13 9 3 13 0 0 15 0 9 13 13 2
20 3 16 3 0 9 13 2 13 3 13 1 9 2 13 3 9 3 9 3 2
6 13 3 15 3 13 2
25 3 3 9 0 13 15 15 0 2 1 3 9 9 13 2 15 3 0 0 13 3 3 13 2 2
27 3 3 0 13 2 16 3 9 13 9 2 13 1 9 2 9 0 1 2 9 3 13 9 3 9 13 2
8 0 3 3 13 13 0 9 2
7 2 3 15 3 9 13 2
20 7 15 15 15 13 9 2 7 13 0 9 13 2 15 3 3 13 13 2 2
26 3 13 2 15 3 13 13 1 9 9 2 3 3 9 0 1 9 13 2 9 3 15 13 0 9 2
20 0 3 1 9 13 0 2 3 3 15 0 13 3 3 0 13 3 3 9 2
10 9 3 9 13 1 9 0 3 0 2
29 1 3 9 13 3 3 1 9 9 13 2 7 1 9 9 0 13 13 9 0 2 9 13 2 16 13 13 0 2
10 3 3 13 0 3 13 13 15 9 2
8 15 3 3 13 13 0 9 2
15 7 15 0 13 7 15 13 9 0 2 0 3 13 9 2
24 9 3 0 7 9 13 2 13 1 9 1 15 2 9 3 3 0 9 13 13 7 15 13 2
35 16 3 15 15 9 13 2 7 13 0 3 13 7 13 0 0 2 3 15 9 3 3 0 13 3 13 2 7 1 9 0 13 9 13 2
14 15 3 3 3 13 15 3 0 13 7 0 13 2 2
11 3 13 2 15 3 3 0 3 13 9 2
5 9 3 13 0 2
7 15 15 0 13 7 13 2
7 0 3 9 0 13 13 2
6 3 0 9 13 9 2
17 16 3 3 13 9 0 9 2 0 3 13 15 3 0 0 13 2
10 16 3 3 13 9 2 13 13 2 2
9 3 13 9 2 15 3 13 9 2
15 3 3 13 13 9 1 9 2 13 3 13 1 0 9 2
8 13 3 0 9 1 9 9 2
8 13 3 13 3 1 0 9 2
32 3 16 3 9 13 0 9 2 13 3 1 9 9 3 0 2 3 9 13 0 9 2 9 3 13 9 3 13 1 3 13 2
7 15 3 3 3 0 13 2
13 3 3 13 16 3 9 0 13 13 2 9 13 2
12 3 3 13 3 2 16 9 13 9 13 9 2
6 15 3 15 0 13 2
15 15 3 13 13 7 13 0 9 7 1 9 13 0 0 2
8 3 9 13 7 13 13 3 2
18 15 3 9 0 13 2 13 3 9 9 3 13 2 15 3 3 13 2
9 3 15 13 13 7 13 0 2 2
8 3 15 0 1 9 0 13 2
9 3 3 13 2 7 3 13 13 2
30 3 15 9 0 13 1 9 0 2 16 3 3 15 0 9 3 9 15 13 9 0 1 9 13 2 13 3 9 0 2
20 3 15 9 0 0 0 13 9 2 3 3 15 15 9 13 13 1 3 9 2
10 3 13 13 2 15 3 13 0 9 2
9 0 3 9 7 9 0 9 13 2
11 15 3 3 9 3 13 2 9 13 0 2
8 15 7 9 0 1 9 13 2
7 15 3 9 13 1 9 2
18 3 3 3 9 0 3 13 1 9 2 7 3 15 3 13 3 13 2
11 2 3 13 15 0 13 7 13 9 13 2
10 0 15 9 13 9 13 3 3 13 2
7 0 3 3 10 3 13 2
5 15 3 13 9 2
22 3 1 9 2 3 3 0 9 13 2 13 13 2 16 9 0 13 13 1 9 0 2
14 0 3 13 9 1 0 2 13 3 9 7 9 0 2
12 7 15 13 15 13 2 3 3 15 13 2 2
17 3 13 2 13 3 0 9 9 1 9 9 13 2 13 3 9 2
20 15 3 16 3 13 9 13 3 9 2 13 2 3 3 15 9 13 9 0 2
17 3 16 9 7 9 1 9 13 2 9 3 13 7 9 9 13 2
19 3 3 15 3 13 13 9 3 0 9 3 0 2 3 3 0 15 13 2
6 3 15 3 3 13 2
13 10 9 0 13 1 9 2 16 3 3 9 13 2
10 13 3 15 15 3 13 9 7 9 2
14 15 3 3 3 13 0 9 13 2 13 3 9 9 2
12 10 9 3 16 3 3 13 2 0 0 13 2
7 15 3 13 13 0 9 2
11 0 0 13 1 9 16 1 9 9 13 2
7 13 3 15 15 3 13 2
15 3 3 1 9 13 3 0 13 2 16 13 9 0 13 2
3 3 13 2
19 15 3 13 9 15 2 15 15 13 2 3 16 3 9 13 9 3 13 2
7 3 3 15 9 13 0 2
8 3 3 3 9 13 13 2 2
18 3 13 2 9 3 1 9 13 2 0 9 13 2 0 3 9 13 2
26 3 16 3 13 9 3 13 2 9 3 3 13 13 1 9 0 2 0 3 3 13 7 13 0 9 2
20 15 3 0 0 13 9 9 2 9 13 9 1 0 2 13 3 3 3 13 2
17 1 3 3 0 9 9 0 13 2 7 13 13 9 3 7 9 2
22 3 15 3 15 3 13 13 2 16 13 9 3 3 2 15 3 2 0 1 9 9 2
9 3 3 15 13 16 13 9 2 2
8 15 3 3 9 13 9 13 2
29 3 13 2 0 9 9 13 2 1 9 13 1 0 9 13 0 9 0 9 13 2 16 3 3 9 0 9 13 2
17 3 15 9 13 2 16 13 9 2 15 15 3 1 13 3 13 2
26 15 3 15 13 1 0 9 2 9 3 15 13 1 9 13 3 13 7 13 2 1 15 3 13 2 2
10 3 3 13 2 15 3 0 13 9 2
24 15 3 13 2 0 9 9 13 2 13 0 9 0 9 13 2 16 3 3 9 0 9 13 2
10 9 3 3 3 1 9 13 9 13 2
8 1 15 3 12 9 0 13 2
9 0 3 3 15 3 9 13 9 2
8 15 3 3 0 9 13 13 2
14 1 3 15 9 9 13 0 13 2 0 3 9 13 2
31 3 15 15 3 3 13 0 9 2 7 3 9 13 7 9 7 9 2 15 3 15 1 9 0 13 9 2 3 13 13 2
5 15 3 13 0 2
12 15 3 9 0 3 13 9 13 3 1 9 2
13 3 3 3 3 3 9 9 1 13 2 7 13 2
8 15 7 9 0 1 9 13 2
8 15 3 3 9 13 9 13 2
23 16 3 15 9 0 1 9 3 13 0 0 13 2 0 13 15 13 13 2 7 15 15 2
20 16 3 3 15 0 9 7 9 13 2 3 3 15 13 13 1 9 13 2 2
8 3 13 9 0 13 1 9 2
24 3 16 3 13 9 3 13 2 9 3 13 1 9 3 9 3 2 1 3 9 13 0 13 2
27 15 3 16 3 9 13 7 13 9 2 1 3 3 9 0 13 7 9 2 1 3 9 13 1 9 13 2
15 9 3 0 9 13 13 0 0 2 1 0 9 2 13 2
6 1 3 0 13 9 2
14 9 3 0 9 13 13 2 9 0 13 2 13 13 2
14 9 3 9 13 1 9 9 9 13 2 0 9 13 2
25 15 3 1 9 0 13 9 13 2 3 16 9 7 9 1 9 13 2 15 3 9 13 9 9 2
24 3 3 15 13 2 16 13 9 0 1 15 9 2 9 15 9 3 13 2 16 3 13 2 2
8 15 3 3 9 13 9 13 2
21 13 3 15 15 1 0 9 3 13 2 7 16 3 9 0 9 13 0 0 3 2
9 3 15 15 3 13 1 9 0 2
16 3 9 0 3 3 13 2 0 3 3 13 2 0 15 13 2
15 3 13 0 9 2 15 1 0 0 9 3 9 9 13 2
13 13 3 3 3 9 0 9 15 13 13 9 0 2
7 3 15 15 0 9 13 2
8 3 3 3 15 9 13 13 2
8 0 3 0 3 13 0 3 2
39 0 3 15 15 13 7 13 2 3 3 15 3 0 1 13 3 3 3 13 2 7 15 3 15 13 9 0 0 2 15 0 15 15 13 9 3 3 13 2
9 15 3 3 13 0 0 9 13 2
4 0 13 13 2
15 13 3 15 9 0 2 15 15 3 0 1 9 13 2 2
11 3 13 2 15 3 3 9 1 9 13 2
7 15 3 3 13 9 0 2
8 3 3 15 13 3 3 13 2
43 13 3 9 0 9 2 0 3 9 9 3 9 0 2 15 13 2 16 3 3 9 3 1 0 9 2 13 7 13 2 15 13 0 9 2 13 2 3 9 0 0 13 2
13 0 15 9 0 1 9 13 13 7 9 13 2 2
7 15 3 3 13 0 9 2
20 3 3 3 13 9 3 0 3 9 1 15 2 16 3 15 15 13 13 2 2
29 3 15 3 0 1 0 13 2 9 3 1 9 9 9 13 7 9 13 2 1 0 9 2 3 3 3 9 13 2
27 3 16 3 9 13 7 13 9 3 1 9 2 15 3 13 15 10 3 3 2 3 3 3 15 13 9 2
11 3 13 2 15 3 13 13 13 3 9 2
11 3 15 13 7 13 2 16 15 3 13 2
15 3 3 13 3 9 2 3 3 3 1 0 0 13 2 2
7 15 3 13 13 0 9 2
5 2 13 2 13 2
6 15 3 3 13 13 2
9 3 13 2 15 3 3 3 13 2
21 13 3 15 2 16 3 15 9 13 13 2 13 2 16 3 13 0 13 9 2 2
12 13 3 7 1 9 0 13 9 2 0 0 2
6 1 3 9 13 9 2
8 9 3 3 15 9 0 13 2
13 15 13 2 9 3 9 7 9 9 13 3 13 2
14 15 3 1 9 13 9 9 0 0 7 9 2 13 2
8 10 3 0 1 9 9 13 2
20 3 3 3 9 0 13 9 2 3 0 2 1 3 0 13 9 3 1 9 2
11 9 3 3 13 9 2 3 0 13 9 2
6 12 3 3 13 9 2
15 15 3 13 13 9 3 13 1 3 13 2 0 7 0 2
5 13 3 9 9 2
20 2 3 3 3 3 3 0 0 13 2 16 3 10 0 13 9 3 10 0 2
24 3 16 3 3 9 0 13 2 3 13 9 13 2 7 13 1 9 13 13 13 0 9 0 2
11 3 1 15 13 2 15 3 3 13 13 2
23 16 3 13 1 9 9 0 2 0 15 1 9 9 9 1 9 9 13 9 0 13 2 2
10 3 13 2 7 13 3 13 9 9 2
11 3 3 15 1 9 13 2 7 13 3 2
7 3 13 2 9 3 13 2
13 15 3 9 13 3 13 2 0 3 13 9 13 2
18 3 3 15 9 3 13 0 2 15 3 13 13 2 13 3 9 1 2
7 3 9 0 13 9 2 2
24 6 3 9 13 0 9 3 1 9 2 7 1 9 13 2 16 9 3 3 13 0 9 2 2
20 3 13 15 3 13 3 3 13 2 3 15 13 2 3 3 3 9 13 9 2
13 3 3 3 13 2 1 3 9 13 2 1 9 2
5 15 3 13 3 2
17 15 1 3 9 9 13 15 13 2 9 3 0 9 13 13 13 2
17 0 3 9 7 0 9 13 13 2 1 3 15 13 9 9 0 2
7 1 3 15 13 13 9 2
7 3 15 9 13 13 9 2
19 1 0 0 13 2 13 3 15 9 9 7 9 2 9 3 0 13 9 2
7 3 3 15 15 9 13 2
29 13 3 16 0 1 0 9 13 9 2 16 9 3 13 2 1 3 3 9 13 2 15 3 9 9 13 9 2 2
14 2 3 13 2 16 3 3 10 3 0 3 13 0 2
9 3 3 3 13 16 13 15 9 2
11 16 3 13 2 13 2 15 3 13 3 2
15 3 3 15 13 2 16 15 15 3 13 7 13 7 13 2
7 15 3 15 13 13 2 2
8 15 3 13 3 0 0 9 2
4 13 2 13 2
6 15 3 3 13 13 2
9 3 13 3 2 15 3 13 3 2
6 1 3 15 15 13 2
31 9 3 3 3 13 13 13 2 0 2 15 0 0 9 13 2 15 1 3 9 0 13 9 1 0 2 0 0 13 2 2
8 3 15 3 0 1 0 13 2
14 15 3 3 13 0 9 9 1 0 7 9 7 9 2
31 3 3 13 0 13 9 2 1 0 9 2 15 15 1 9 9 3 9 3 3 13 2 16 3 13 9 9 9 0 13 2
30 3 3 3 2 16 13 9 3 13 2 9 3 3 15 3 13 7 9 13 0 2 1 3 3 3 13 0 9 13 2
16 3 15 3 13 13 9 2 3 13 9 2 3 3 13 9 2
7 9 3 1 13 9 2 2
24 16 15 13 7 9 7 3 9 2 0 15 3 13 13 9 2 3 3 13 13 9 7 9 2
13 3 3 3 15 13 0 9 9 9 2 15 13 2
5 7 9 3 13 2
19 3 3 13 9 2 9 3 15 1 9 13 2 15 3 9 0 3 13 2
15 9 3 2 16 3 3 13 9 2 3 3 13 0 13 2
18 0 3 3 9 13 0 9 9 2 16 3 15 1 0 9 13 2 2
15 3 13 13 9 3 13 2 13 3 0 9 1 9 0 2
15 9 3 3 1 9 13 0 9 2 3 13 9 0 9 2
19 15 3 13 13 9 13 2 3 3 9 13 9 0 13 9 9 1 13 2
14 15 13 13 1 9 9 0 2 3 3 3 0 13 2
16 0 3 1 0 13 9 9 2 0 0 0 7 9 2 13 2
8 10 3 0 1 9 9 13 2
22 13 3 1 0 9 1 9 2 13 9 0 2 15 3 9 13 3 7 1 9 13 2
24 9 3 1 15 13 13 9 2 9 3 0 13 0 1 9 7 9 2 3 15 9 13 13 2
15 2 13 10 9 0 13 0 3 13 13 3 0 13 9 2
19 3 13 2 13 3 9 2 16 10 9 13 2 3 3 13 9 0 13 2
10 9 3 3 0 13 13 9 9 2 2
7 15 3 13 13 0 9 2
23 3 3 3 0 13 7 13 3 9 1 2 0 1 9 2 13 3 16 9 1 9 13 2
6 9 3 13 1 9 2
26 3 9 2 3 13 9 9 13 2 16 3 9 1 9 13 2 13 3 15 15 13 0 15 3 0 2
9 3 3 3 3 15 13 13 9 2
18 13 3 13 13 0 9 0 2 3 9 13 2 3 16 9 3 13 2
18 15 3 13 13 2 7 13 0 2 0 3 13 15 13 7 3 13 2
6 3 3 15 3 13 2
9 3 13 2 9 3 9 13 9 2
17 3 13 16 15 9 13 9 3 13 2 15 3 3 1 15 13 2
10 9 3 3 3 15 13 13 15 0 2
18 3 15 3 3 13 2 16 15 0 9 13 1 9 7 9 0 2 2
8 15 3 3 9 13 9 13 2
10 2 13 2 7 15 0 13 0 9 2
15 9 3 13 3 13 3 9 0 2 13 3 3 0 2 2
8 13 3 7 9 9 0 13 2
5 3 0 9 13 2
4 13 15 13 2
4 3 15 13 2
5 13 3 15 3 2
10 0 3 13 0 13 7 13 0 2 2
7 15 3 3 9 13 13 2
17 16 15 0 0 13 9 2 3 3 15 12 9 3 9 13 2 2
18 3 3 13 2 7 9 13 13 9 13 2 15 3 13 0 9 13 2
14 15 3 0 0 13 2 13 3 3 9 9 7 9 2
13 3 3 3 13 9 3 1 9 13 9 13 0 2
11 13 3 1 9 2 7 15 1 9 13 2
11 3 15 13 13 3 0 16 3 0 9 2
9 15 3 3 15 13 1 0 9 2
23 3 3 15 3 9 1 9 13 0 0 7 3 13 9 2 0 0 13 7 15 13 13 2
16 13 3 9 3 0 0 3 0 15 3 3 13 7 0 13 2
8 13 3 1 9 9 9 9 2
23 3 3 3 3 15 13 0 9 3 1 9 13 7 9 13 2 9 3 1 9 13 13 2
29 15 3 9 13 2 13 9 0 2 3 3 0 9 0 9 13 2 1 3 9 13 7 0 9 2 0 3 13 2
7 3 3 1 9 13 9 2
9 15 3 9 13 1 9 13 13 2
12 13 3 0 9 0 3 7 9 9 3 9 2
17 1 3 9 0 9 0 9 0 13 2 3 3 15 13 13 0 2
6 1 3 0 3 13 2
17 3 15 0 3 13 0 9 2 15 3 13 0 2 15 13 9 2
10 3 3 3 3 15 13 9 13 2 2
10 2 15 9 15 9 13 2 9 9 2
17 13 3 1 0 2 0 1 9 2 16 3 0 9 7 9 13 2
4 3 0 13 2
7 15 3 13 13 0 9 2
25 3 15 3 3 1 9 0 9 3 3 9 13 2 15 3 0 13 3 15 15 13 9 13 13 2
6 15 3 0 13 2 2
17 3 13 2 9 3 13 3 3 2 7 15 3 13 9 0 13 2
20 2 3 3 15 3 0 1 9 3 13 3 13 2 16 3 3 9 13 2 2
23 15 3 13 3 9 0 2 3 3 3 15 13 9 9 2 7 0 13 9 2 0 13 2
23 3 3 15 3 1 9 13 1 3 13 2 1 3 3 9 13 0 2 1 3 9 13 2
16 3 15 9 13 9 1 0 2 0 2 15 0 0 9 13 2
18 3 16 3 9 3 9 7 9 13 2 9 1 9 9 9 13 2 2
10 3 13 2 15 3 3 0 3 13 2
7 3 3 15 13 0 9 2
21 7 3 9 9 13 0 2 0 13 2 13 9 2 9 9 3 7 9 13 2 2
11 3 3 13 9 2 15 3 3 13 9 2
27 9 3 1 3 9 0 9 13 13 2 3 3 3 9 3 13 1 9 2 7 0 13 9 2 0 13 2
16 15 3 16 3 13 0 9 13 1 9 2 1 3 9 13 2
10 2 6 3 0 15 13 0 9 2 2
9 15 3 3 9 9 1 9 13 2
9 2 6 3 1 9 9 0 13 2
10 3 3 15 0 3 0 9 13 2 2
7 15 3 3 13 0 9 2
7 9 3 3 0 9 13 2
9 9 15 0 13 1 9 9 13 2
4 9 3 13 2
18 3 0 3 0 13 3 13 3 2 0 3 9 0 13 0 9 2 2
13 15 3 3 3 13 1 9 9 2 13 1 9 2
9 15 3 1 15 13 13 0 9 2
5 0 3 13 2 2
11 0 15 3 13 2 13 3 15 0 9 2
14 12 3 3 15 9 13 2 12 3 9 13 1 9 2
7 0 3 15 13 9 13 2
8 3 3 3 9 13 0 13 2
8 3 15 15 13 13 1 9 2
15 13 3 9 9 0 13 2 9 13 2 3 9 9 13 2
11 3 3 3 3 15 13 9 13 2 13 2
8 0 3 13 9 0 3 2 2
7 15 3 3 13 0 9 2
11 2 13 2 3 13 2 16 9 0 13 2
5 15 3 0 13 2
20 16 3 9 13 7 13 1 0 9 2 3 3 1 0 9 9 13 9 2 2
14 3 13 2 9 3 0 13 2 3 3 9 0 13 2
12 13 3 9 2 3 3 3 9 9 0 13 2
10 2 13 15 2 10 9 3 3 13 2
9 3 13 15 15 9 13 0 9 2
20 3 3 7 3 0 9 9 13 0 3 2 3 3 3 15 9 7 9 13 2
12 0 3 15 13 2 15 3 1 9 13 0 2
12 3 13 2 13 3 9 2 16 10 9 13 2
7 3 3 13 9 0 13 2
13 13 15 15 9 1 9 13 2 3 9 3 13 2
21 16 3 3 15 13 0 0 13 2 13 15 9 3 9 3 2 15 15 3 13 2
9 9 3 3 13 1 9 9 13 2
8 13 3 15 15 3 13 2 2
8 15 3 3 13 0 0 9 2
11 13 3 3 1 0 2 0 3 13 9 2
15 3 9 0 13 9 2 15 9 3 9 3 0 9 13 2
31 3 3 3 2 16 15 0 9 1 9 13 3 15 0 13 13 9 13 2 3 3 15 9 15 3 13 3 3 15 0 2
15 3 3 9 1 9 13 13 2 13 3 2 1 9 13 2
14 3 3 15 13 9 1 0 9 2 3 13 1 9 2
6 9 3 3 0 13 2
10 13 3 0 2 16 15 0 13 2 2
12 3 13 2 13 3 9 2 16 10 9 13 2
8 15 3 1 9 13 13 9 2
12 7 15 3 13 0 7 3 3 13 1 9 2
17 2 13 1 9 2 15 3 3 13 3 0 2 9 13 9 9 2
8 3 15 13 13 1 9 13 2
7 15 3 3 13 0 9 2
7 13 2 16 3 3 13 2
13 3 3 3 15 3 0 9 9 13 0 13 2 2
17 3 3 9 9 0 13 2 3 13 9 2 16 3 13 10 0 2
6 15 3 3 0 13 2
13 0 3 15 0 13 2 7 13 9 16 15 13 2
15 0 3 0 13 0 2 15 9 13 16 15 9 13 2 2
8 15 3 3 9 13 9 13 2
5 15 3 13 13 2
9 3 15 15 0 7 0 13 2 2
35 3 13 2 15 3 3 3 13 0 1 9 2 13 3 3 9 9 7 9 13 3 13 1 9 2 13 3 9 3 9 3 2 0 9 2
7 15 3 9 7 9 13 2
7 3 3 3 13 0 9 2
22 13 3 1 0 0 2 15 1 9 13 9 2 1 3 13 9 0 0 13 7 13 2
16 3 3 15 13 9 3 3 9 2 9 3 3 0 13 13 2
5 9 3 9 13 2
8 15 3 13 9 9 1 9 2
15 9 3 0 13 0 2 16 13 13 2 16 3 15 13 2
12 3 13 16 3 15 13 0 2 13 3 13 2
5 15 3 13 3 2
14 9 3 0 15 13 2 3 3 15 15 13 0 13 2
15 13 3 15 13 9 3 3 15 2 9 3 9 13 13 2
22 9 3 7 15 3 13 2 16 15 13 2 16 15 9 3 13 9 7 9 13 9 2
10 9 3 3 15 3 3 3 13 3 2
14 3 3 3 15 15 13 13 0 1 9 9 9 2 2
7 15 3 13 13 9 9 2
18 15 3 0 13 13 0 2 3 3 3 0 9 9 13 9 3 9 2
10 13 3 2 16 0 13 3 15 13 2
8 3 3 3 15 0 9 13 2
12 3 15 3 1 9 0 9 1 0 3 13 2
14 15 3 13 0 9 9 2 0 3 3 13 13 9 2
10 10 9 3 7 9 13 0 9 13 2
5 3 13 3 2 2
17 3 13 2 15 3 3 0 13 13 2 1 3 3 0 0 13 2
17 9 15 9 13 1 9 2 15 1 9 13 9 3 7 9 13 2
16 0 3 3 13 0 3 13 2 15 15 3 13 13 0 13 2
9 3 13 9 2 15 3 13 9 2
7 15 3 13 13 0 9 2
10 3 15 9 13 0 2 16 9 13 2
11 3 13 2 15 3 3 0 13 3 13 2
18 3 16 3 13 3 13 3 10 9 2 15 3 3 13 0 9 9 2
9 3 13 2 15 3 3 0 13 2
27 3 9 13 3 9 1 9 2 13 3 9 0 3 0 3 2 13 3 15 0 9 9 3 0 3 9 2
9 3 9 3 13 9 13 9 9 2
7 9 3 3 0 3 13 2
9 3 3 15 13 13 1 0 0 2
18 2 3 3 9 9 0 0 13 2 0 1 9 10 9 9 13 2 2
10 3 3 13 2 9 3 3 13 9 2
9 3 3 3 9 13 13 9 13 2
5 9 3 13 9 2
10 9 3 13 9 3 13 1 3 13 2
11 3 1 15 13 2 15 3 3 13 13 2
12 3 13 2 15 3 3 3 1 9 13 9 2
5 1 0 3 13 2
6 15 3 0 9 13 2
24 3 3 13 0 0 9 7 13 16 15 9 13 3 13 2 7 15 3 13 13 3 1 9 2
17 3 3 15 13 13 0 13 2 3 13 2 16 3 15 13 0 2
23 3 3 13 1 9 0 9 2 1 3 13 1 9 13 2 1 3 13 9 13 9 9 2
8 3 9 0 9 13 0 13 2
16 3 9 13 1 9 13 9 2 16 13 9 2 9 3 9 2
8 7 15 1 9 9 13 13 2
13 9 3 15 13 9 2 7 15 13 9 0 13 2
31 2 3 3 13 9 3 9 3 13 2 3 3 15 3 9 7 0 9 13 0 13 2 16 3 15 0 3 0 13 2 2
12 13 3 7 1 9 0 13 9 2 0 0 2
6 1 3 9 13 9 2
11 3 3 15 3 1 9 13 1 3 13 2
10 15 3 13 3 0 13 7 13 9 2
10 3 3 13 2 13 3 9 0 9 2
15 9 3 3 15 0 1 9 13 2 0 9 3 7 9 2
16 9 3 9 1 9 12 13 13 7 9 0 13 2 13 3 2
9 3 3 3 3 0 13 0 2 2
7 15 3 13 13 9 9 2
11 15 15 1 13 13 2 9 3 9 13 2
11 3 15 13 2 15 3 13 7 15 13 2
16 0 0 9 13 9 2 0 0 3 9 1 13 3 7 13 2
17 3 3 3 3 13 0 13 3 2 16 9 13 9 7 9 13 2
16 3 16 3 3 0 9 0 13 2 3 15 13 0 13 9 2
16 0 3 9 13 0 9 0 1 9 13 9 9 3 9 3 2
27 3 3 15 3 13 1 9 0 13 2 0 3 0 13 9 7 9 13 2 9 3 0 0 7 0 9 2
20 3 3 15 3 3 9 0 13 2 7 15 3 9 9 9 13 2 15 13 2
18 3 15 9 3 13 2 3 3 13 0 2 16 13 0 1 0 9 2
16 3 3 3 3 13 13 9 7 0 2 16 3 9 13 2 2
18 3 13 2 7 13 13 0 9 2 3 3 1 9 13 9 9 9 2
12 3 15 13 1 9 0 13 9 2 13 9 2
6 3 3 0 13 9 2
7 3 3 3 3 13 9 2
13 13 3 3 15 9 9 1 9 7 9 3 13 2
11 3 3 3 1 3 13 1 9 3 13 2
10 0 3 13 9 3 13 1 3 13 2
9 15 3 3 9 9 1 9 13 2
7 15 3 3 13 0 9 2
20 9 3 15 3 9 2 15 9 13 2 13 2 1 15 0 13 0 1 9 2
16 3 15 9 3 7 9 13 13 2 16 3 15 13 1 9 2
7 0 3 3 13 1 9 2
4 13 3 2 2
20 9 0 1 0 9 13 2 13 3 13 2 13 3 15 9 0 3 1 9 2
14 3 3 3 0 9 0 9 13 2 16 15 13 0 2
22 9 3 15 0 9 0 13 0 2 0 3 0 9 13 2 16 3 13 9 9 0 2
16 7 15 0 7 0 13 13 2 0 3 3 15 13 0 9 2
14 15 3 0 9 13 2 7 3 13 9 9 13 3 2
10 2 3 15 3 0 0 1 9 13 2
31 7 15 3 0 9 13 9 0 3 3 2 16 3 13 1 9 9 13 2 9 13 0 0 9 2 16 0 13 0 2 2
9 3 13 13 9 0 2 3 0 2
8 1 15 3 3 0 12 13 2
8 9 3 3 15 0 3 13 2
19 15 3 3 13 9 2 9 3 3 9 13 2 0 3 13 1 9 13 2
10 9 3 13 3 3 1 9 9 13 2
10 15 3 9 9 3 1 9 13 2 2
8 15 3 3 9 13 9 13 2
6 3 3 3 0 13 2
8 3 3 3 13 13 0 13 2
17 1 3 15 13 13 3 0 15 0 13 2 15 3 3 13 0 2
19 3 3 3 9 3 7 9 9 13 9 9 2 9 3 15 3 0 13 2
8 3 15 3 0 1 0 13 2
6 9 3 9 13 9 2
7 15 3 13 3 9 9 2
18 16 0 3 13 10 0 9 13 2 0 3 9 13 0 7 0 3 2
4 3 3 13 2
7 0 3 15 13 0 9 2
19 3 3 3 16 3 13 13 1 0 9 2 0 1 9 13 15 9 13 2
16 3 3 13 7 3 15 13 9 2 7 3 13 3 1 9 2
6 15 3 3 0 13 2
16 13 9 7 9 1 9 3 3 2 7 3 3 15 3 13 2
17 3 16 3 9 13 13 2 13 15 3 13 2 0 1 9 13 2
5 2 0 3 13 2
6 15 3 3 0 13 2
17 9 3 13 16 3 0 9 13 0 15 2 15 3 9 9 13 2
9 3 15 0 9 9 7 9 13 2
8 9 3 15 9 10 3 13 2
32 15 3 0 3 9 7 0 9 13 13 7 0 13 2 0 15 3 13 9 7 0 9 2 9 9 0 2 7 0 9 13 2
8 3 3 0 9 0 13 2 2
27 3 13 2 13 3 9 0 9 2 16 15 3 9 13 2 13 3 9 0 9 2 9 3 15 0 13 2
7 3 3 0 13 9 13 2
9 3 13 9 2 15 3 13 9 2
8 9 3 3 13 13 9 0 2
9 9 3 13 0 0 9 2 0 2
7 9 3 9 0 3 13 2
5 9 3 13 0 2
9 0 3 3 0 9 0 0 13 2
8 15 3 13 0 1 0 13 2
10 3 9 12 13 1 9 2 16 13 2
19 1 3 9 0 13 2 0 3 2 0 2 0 13 9 2 7 9 13 2
7 3 3 13 9 9 0 2
18 15 3 1 9 13 2 13 3 0 13 1 9 2 7 9 13 9 2
7 3 15 0 9 0 13 2
14 16 3 3 3 13 0 9 13 2 3 15 15 13 2
6 9 3 3 13 2 2
12 3 13 2 15 3 13 2 1 0 3 13 2
27 15 3 3 13 9 0 2 15 9 3 13 2 13 3 9 2 9 3 3 13 2 13 3 3 9 9 2
18 3 3 3 3 13 9 1 9 9 2 7 15 3 9 13 7 13 2
7 15 3 9 13 0 9 2
15 3 3 15 9 13 9 2 7 3 15 3 0 9 13 2
25 3 15 15 3 9 0 0 13 2 15 15 15 1 9 13 9 0 9 13 2 13 9 0 2 2
9 15 3 3 3 13 13 0 9 2
6 3 13 9 13 9 2
13 13 3 13 1 9 2 13 3 1 9 0 9 2
6 13 3 15 0 13 2
11 3 15 1 9 13 13 13 1 0 13 2
14 0 3 15 9 13 9 0 2 15 3 3 0 13 2
20 9 3 3 3 0 13 9 9 13 0 2 16 3 3 13 9 9 9 9 2
5 9 3 9 13 2
9 3 3 15 9 0 1 9 13 2
20 3 15 13 9 9 13 0 1 9 2 16 3 15 1 9 3 3 0 2 2
9 13 3 2 3 3 13 9 0 2
16 3 3 15 9 3 0 13 2 9 3 13 9 3 9 13 2
28 3 16 3 3 9 0 13 2 3 13 9 13 2 7 13 1 9 13 2 16 3 13 13 0 9 0 2 2
7 15 3 13 13 0 9 2
40 6 3 3 3 9 13 13 2 15 3 0 2 9 2 0 2 0 13 9 2 9 2 0 2 15 3 9 3 0 2 0 3 13 2 13 3 1 9 9 2
43 16 3 3 3 9 3 13 9 3 2 3 15 9 13 7 12 9 7 9 0 2 1 9 13 2 3 3 15 13 0 1 0 13 2 3 3 3 15 10 9 13 13 2
10 3 3 13 2 7 15 9 13 0 2
17 7 3 15 13 0 13 7 0 2 16 1 0 7 3 0 13 2
29 16 3 9 13 7 13 1 0 9 2 3 3 15 10 9 2 3 0 3 3 13 2 13 13 1 9 3 2 2
17 3 13 2 9 3 13 3 3 2 7 15 3 13 9 0 13 2
15 3 3 15 9 13 9 2 7 3 15 3 0 9 13 2
6 3 3 13 9 13 2
11 3 9 9 1 9 13 9 2 9 13 2
8 15 3 3 9 13 9 0 2
15 9 3 3 13 13 2 3 15 3 13 13 0 1 9 2
16 9 3 13 1 9 0 2 3 3 15 13 13 1 0 0 2
11 2 6 13 10 9 13 3 13 16 13 2
7 3 3 15 0 9 13 2
6 9 3 15 15 13 2
11 3 3 13 13 3 13 2 16 9 13 2
8 13 3 3 15 15 3 2 2
18 3 13 2 15 3 3 0 3 1 9 13 9 13 2 15 3 13 2
14 3 3 2 9 3 13 9 2 16 13 13 3 13 2
10 10 9 3 13 1 9 9 9 13 2
7 15 3 0 13 9 2 2
10 3 13 2 15 3 0 13 9 13 2
5 9 3 13 9 2
6 13 3 3 0 3 2
9 15 3 9 13 9 13 0 9 2
19 3 16 13 3 13 3 0 13 9 2 13 3 13 13 0 1 9 0 2
14 3 10 1 9 13 0 9 2 9 9 1 9 13 2
7 3 3 9 9 0 13 2
12 3 9 0 9 13 2 16 3 15 13 13 2
24 2 1 9 13 2 16 3 15 13 0 3 3 13 13 9 2 3 13 2 0 9 13 9 2
27 1 3 3 3 15 0 1 9 13 9 16 3 13 2 9 13 1 15 2 0 13 13 3 9 7 9 2
6 0 3 13 9 9 2
6 15 3 3 0 13 2
12 3 3 13 13 2 16 3 9 13 9 2 2
8 15 3 3 13 0 9 9 2
10 3 3 2 15 15 3 13 9 13 2
11 9 3 3 13 13 2 15 3 13 2 2
8 15 3 3 9 13 9 13 2
16 3 3 0 13 15 3 0 3 9 13 2 3 3 13 2 2
10 3 3 13 2 15 3 0 13 9 2
7 13 3 9 9 3 13 2
18 15 3 3 13 9 7 0 9 13 9 3 7 9 0 9 3 0 2
13 1 3 9 9 2 0 9 13 2 9 0 13 2
8 3 3 9 13 15 9 3 2
7 15 3 13 13 9 9 2
11 2 13 7 1 0 9 13 3 3 13 2
10 0 3 9 13 9 2 15 9 13 2
19 3 15 3 13 2 15 3 13 3 2 16 3 3 9 7 9 0 13 2
9 15 3 15 13 13 3 0 2 2
26 3 13 2 9 3 1 9 13 13 1 9 2 9 1 13 2 3 3 13 2 16 15 0 9 13 2
10 3 3 3 3 13 7 9 0 13 2
14 3 10 1 9 13 0 9 2 9 9 1 9 13 2
14 10 3 13 1 9 0 9 2 9 0 7 0 9 2
16 15 1 3 9 9 13 2 3 3 13 2 0 9 7 9 2
21 15 3 9 13 9 2 7 1 9 9 13 0 1 0 2 3 1 0 13 9 2
6 3 13 3 0 9 2
7 13 3 9 0 1 9 2
18 15 3 1 3 9 0 13 7 9 7 9 2 3 3 9 9 13 2
20 9 3 1 9 3 13 2 0 3 1 0 13 9 0 2 9 13 7 13 2
8 10 3 9 13 9 0 3 2
9 7 3 3 9 13 13 3 2 2
9 15 3 3 3 13 13 9 9 2
4 9 3 13 2
29 0 0 7 9 9 13 7 3 15 3 9 1 9 13 0 0 7 3 13 9 2 0 0 13 7 15 13 13 2
17 13 3 9 3 0 2 0 3 0 15 3 3 13 7 0 13 2
5 3 9 13 9 2
4 13 3 3 2
16 15 3 3 15 1 9 9 13 13 2 16 3 0 13 2 2
26 0 3 3 13 2 16 1 15 13 0 16 10 9 13 1 9 0 1 9 13 2 16 3 13 2 2
9 3 3 3 9 9 1 9 13 2
6 13 3 15 13 2 2
17 3 13 2 15 3 3 3 13 13 9 0 7 1 0 9 13 2
7 3 13 3 9 0 9 2
7 15 3 9 13 0 9 2
5 15 3 13 9 2
7 15 3 13 13 9 9 2
32 3 15 3 10 3 0 13 0 1 9 2 3 3 0 13 9 7 0 9 2 16 15 3 9 13 9 13 3 3 13 0 2
20 3 3 15 15 13 9 1 0 13 3 13 3 13 2 16 0 13 0 3 2
20 3 15 15 9 13 2 7 15 3 0 2 13 3 13 13 15 9 9 2 2
7 15 3 13 3 9 9 2
4 3 3 13 2
7 0 3 15 13 0 9 2
16 3 3 3 9 13 3 9 3 3 15 9 2 15 9 13 2
7 3 9 13 0 13 9 2
5 15 3 9 13 2
5 15 3 9 13 2
20 9 3 15 0 13 9 9 2 13 0 9 2 1 9 13 2 0 7 0 2
5 3 3 0 13 2
10 2 3 13 2 15 3 13 9 0 2
16 3 3 0 3 13 0 9 2 9 3 13 2 16 9 13 2
9 3 0 3 13 15 7 13 0 2
12 3 15 3 13 2 3 3 13 2 1 9 2
11 3 3 3 15 13 0 9 2 3 13 2
12 3 3 1 9 13 0 3 3 1 9 2 2
7 15 3 13 13 9 9 2
5 3 1 15 13 2
10 3 3 15 9 3 13 0 16 13 2
10 3 3 3 13 15 15 13 7 13 2
16 9 15 9 13 2 0 1 9 9 2 0 7 9 2 0 2
21 3 15 3 1 9 9 9 1 13 3 9 2 15 3 9 0 9 2 0 9 2
8 3 9 15 13 7 0 13 2
13 3 3 15 3 13 9 9 2 13 3 13 9 2
19 13 3 1 9 2 3 3 9 9 2 1 9 0 2 3 3 13 9 2
7 3 3 9 13 3 13 2
10 9 3 15 13 0 3 13 0 3 2
15 15 3 3 0 7 0 13 9 13 1 9 9 9 1 2
17 15 3 15 1 9 13 3 13 2 3 13 2 0 1 9 13 2
26 7 15 10 0 9 2 15 1 0 13 2 3 9 13 7 9 9 13 7 9 13 2 16 13 9 2
8 3 12 3 13 9 0 0 2
18 13 3 9 9 0 3 3 1 9 13 13 2 0 3 15 13 9 2
7 13 9 0 13 0 0 2
17 3 3 9 13 1 0 9 2 15 3 9 13 2 16 9 13 2
8 13 3 3 15 9 13 13 2
13 3 15 13 0 9 9 13 2 13 0 9 13 2
21 3 9 9 3 13 0 13 9 2 9 3 3 16 9 13 7 9 3 1 9 2
7 9 3 15 3 9 13 2
14 15 3 16 3 13 0 9 2 3 15 9 13 13 2
22 13 15 0 15 1 9 9 13 2 0 3 0 13 2 7 9 2 15 15 13 2 2
7 15 3 13 13 9 9 2
15 3 3 15 0 9 13 1 15 3 13 7 0 13 9 2
8 3 15 13 3 15 13 9 2
9 9 0 0 13 0 9 2 0 2
8 3 15 9 9 13 9 0 2
5 3 3 0 13 2
11 1 0 9 9 13 0 9 2 13 13 2
15 10 3 9 13 1 9 0 2 0 3 9 9 1 0 2
11 3 3 13 0 2 0 3 13 9 3 2
8 3 3 0 3 0 13 9 2
31 3 13 7 15 13 1 9 3 9 2 3 15 9 13 0 1 9 13 2 7 15 3 3 9 2 16 0 9 13 0 2
6 0 3 0 13 0 2
21 7 15 15 0 9 7 9 13 0 0 7 0 9 2 3 3 13 0 1 9 2
9 7 3 15 9 0 0 0 13 2
9 7 15 15 13 2 0 13 3 2
13 0 1 9 2 0 2 0 2 9 3 9 13 2
16 13 3 15 0 0 15 9 9 2 16 15 9 0 13 2 2
7 3 3 15 9 13 13 2
22 0 3 15 9 15 13 2 0 13 2 13 1 9 2 9 3 13 0 0 9 13 2
12 15 3 3 13 3 3 13 0 1 0 9 2
15 3 3 0 9 0 1 9 9 13 13 9 3 0 2 2
7 15 3 13 13 9 9 2
5 13 3 3 0 2
25 3 3 15 3 0 13 9 13 0 2 15 9 13 9 13 2 16 9 2 15 13 9 0 13 2
10 3 9 3 13 2 15 3 13 9 2
24 3 3 15 13 3 3 13 16 3 9 15 1 9 13 3 2 9 9 1 9 9 2 0 2
10 3 13 9 0 7 0 13 1 9 2
16 3 9 9 13 7 9 0 1 9 9 2 9 1 9 13 2
8 13 3 0 9 3 7 9 2
6 15 3 9 13 9 2
8 10 3 0 13 0 1 9 2
39 15 3 3 1 9 9 13 9 1 9 2 9 1 9 2 15 0 13 2 15 3 15 1 9 9 3 13 7 15 0 13 13 3 15 13 0 3 0 2
7 3 3 3 3 9 13 2
17 3 1 9 0 0 9 13 9 2 3 3 3 15 13 9 0 2
26 13 3 1 15 0 2 13 1 9 2 9 13 7 0 13 9 2 15 3 15 13 0 1 9 9 2
5 3 15 3 13 2
10 13 3 13 9 9 9 1 9 0 2
9 7 15 9 13 2 0 13 9 2
19 3 3 3 1 0 9 0 3 3 13 2 0 15 1 9 9 13 9 2
31 15 3 1 9 13 13 2 16 9 1 9 0 9 9 13 2 16 13 0 1 0 9 3 3 13 2 7 3 7 3 2
24 2 3 15 3 3 13 0 7 13 3 3 3 2 3 3 3 1 0 7 0 9 0 13 2
6 3 3 15 9 13 2
18 13 3 9 0 2 9 0 7 0 2 9 3 9 0 2 15 13 2
9 3 3 15 15 0 13 3 13 2
17 15 0 9 13 3 9 2 10 3 13 9 2 15 3 13 2 2
7 15 3 3 13 0 9 2
19 3 3 3 13 9 3 0 3 9 1 15 2 16 3 15 15 13 13 2
11 3 15 3 1 9 13 2 16 13 3 2
37 3 3 9 3 9 13 2 3 3 15 9 13 2 16 3 0 9 13 1 9 0 9 13 1 9 2 16 3 13 3 2 9 0 13 7 13 2
13 3 3 15 9 3 3 13 2 3 3 13 3 2
5 9 3 0 13 2
24 15 3 0 0 13 7 0 13 2 15 3 13 0 9 9 3 0 2 3 13 3 13 0 2
7 15 3 13 13 9 9 2
15 0 3 3 9 0 1 9 13 7 3 13 0 9 0 2
10 3 3 15 15 9 9 0 9 13 2
35 3 3 9 9 13 0 15 15 15 9 1 9 13 2 16 3 15 9 13 0 2 0 13 2 15 15 3 13 0 9 0 3 15 3 2
10 15 3 3 3 13 9 13 15 2 2
7 15 3 3 13 0 9 2
22 3 3 3 15 9 13 3 9 0 0 0 13 9 2 16 15 3 3 13 0 13 2
34 13 3 15 9 0 9 9 13 15 0 0 3 13 7 13 2 13 9 2 16 15 0 13 9 2 15 15 9 13 2 13 3 3 2
11 3 3 9 3 15 13 9 15 3 9 2
8 3 3 1 9 9 13 2 2
20 3 3 13 2 9 3 13 9 9 2 9 3 13 0 2 9 3 0 13 2
10 3 15 1 9 9 13 0 9 13 2
32 3 3 3 15 0 9 9 0 0 9 13 3 3 0 9 2 0 15 15 13 2 13 16 13 9 3 0 13 3 0 9 2
9 3 3 15 0 3 13 0 9 2
35 3 3 3 0 13 9 9 0 2 16 15 0 9 13 2 3 15 10 9 15 13 0 2 15 3 9 3 7 9 0 13 3 13 13 2
19 3 15 9 13 3 3 0 9 7 15 1 2 16 15 13 3 9 9 2
10 3 3 3 13 9 2 15 3 13 2
26 0 3 9 0 3 13 2 3 3 3 15 13 13 3 13 3 15 9 9 3 9 3 9 13 2 2
7 15 3 13 13 9 9 2
24 3 3 13 2 9 3 9 13 13 15 9 13 2 9 3 13 0 0 2 3 3 0 13 2
12 3 9 13 1 9 2 1 3 9 13 3 2
16 3 3 1 9 13 2 16 15 13 9 13 7 3 9 13 2
8 13 3 3 3 13 9 0 2
7 9 3 15 0 13 9 2
9 15 3 13 9 13 9 7 9 2
7 15 3 15 0 3 13 2
14 9 3 13 9 1 0 9 9 0 13 13 9 15 2
18 15 3 15 9 0 1 9 13 13 9 2 9 3 13 1 3 13 2
6 0 3 3 13 2 2
7 3 3 9 9 13 0 2
30 3 15 3 2 16 3 13 0 1 0 9 13 3 2 3 3 15 9 13 2 15 15 15 13 7 15 13 13 2 2
11 15 1 13 9 2 16 15 13 0 9 2
15 15 3 3 9 3 7 9 9 9 3 13 9 3 0 2
16 9 3 9 9 13 9 13 3 15 9 3 7 0 9 0 2
8 9 3 9 13 0 9 13 2
27 15 13 1 3 13 2 7 15 13 0 2 13 3 3 3 13 3 9 2 13 3 3 2 13 3 9 2
18 3 3 3 0 9 1 9 13 13 2 3 3 15 9 13 9 0 2
21 3 3 9 13 0 9 2 13 3 13 1 9 2 7 9 7 7 0 9 9 2
7 1 15 3 0 9 13 2
18 9 3 3 0 13 9 1 9 0 9 2 10 3 1 9 13 9 2
13 1 15 3 0 9 13 1 9 2 13 0 9 2
10 3 3 3 1 9 0 13 0 9 2
25 15 3 3 3 3 9 13 9 0 13 2 3 3 15 9 13 9 13 2 3 3 9 13 3 2
12 3 3 0 13 2 3 9 13 9 3 0 2
15 15 3 9 3 9 3 1 9 13 9 2 16 13 13 2
19 15 3 0 1 9 13 3 9 2 9 3 9 13 2 13 3 0 3 2
15 10 3 3 0 9 13 13 0 9 9 0 2 13 13 2
30 15 3 3 9 9 0 13 2 9 3 9 0 0 13 3 2 9 3 9 0 13 2 3 3 13 0 1 9 9 2
23 15 3 3 9 3 7 9 9 3 13 7 0 9 13 3 13 0 1 9 13 1 9 2
20 15 3 3 15 3 13 16 15 13 13 9 0 9 2 3 13 1 9 9 2
14 15 9 9 0 13 13 3 13 2 9 3 13 13 2
7 10 3 1 9 13 9 2
6 13 3 9 9 13 2
15 3 3 15 15 3 3 13 2 16 0 9 0 13 2 2
13 13 7 9 13 9 2 13 13 0 9 3 13 2
11 15 3 3 3 13 13 0 3 3 13 2
6 15 3 9 9 13 2
17 3 9 9 13 9 13 0 2 10 3 0 15 1 13 13 3 2
10 15 3 15 13 0 15 0 1 9 2
12 3 3 9 0 13 13 0 9 1 0 9 2
19 3 16 13 7 15 9 13 9 2 13 2 16 15 3 0 1 9 13 2
9 3 3 13 2 7 3 13 13 2
28 16 3 1 15 3 9 13 9 0 2 3 3 9 13 15 13 2 3 3 0 9 1 9 0 13 9 2 2
7 15 3 3 13 0 9 2
20 13 3 0 0 9 0 3 3 0 2 13 3 3 16 15 0 9 7 9 2
28 16 3 1 15 3 9 13 9 0 2 3 3 15 13 1 9 9 2 15 3 15 13 7 15 9 13 2 2
6 3 3 15 15 13 2
10 3 3 3 0 15 13 7 13 0 2
10 3 13 9 9 2 13 3 9 2 2
12 3 3 13 2 9 3 1 9 13 13 9 2
6 10 3 0 13 0 2
24 3 16 13 3 7 13 3 9 2 3 3 3 9 13 9 9 13 2 9 3 1 9 13 2
7 15 3 9 13 0 9 2
20 3 3 3 9 3 13 0 9 2 15 15 3 9 13 0 2 3 13 3 2
8 3 15 3 9 0 13 9 2
18 9 3 3 13 13 2 13 2 1 3 0 9 13 7 0 1 9 2
25 3 16 9 13 2 13 3 9 0 2 13 1 9 2 0 3 15 1 0 9 0 9 13 13 2
19 9 3 0 16 13 3 0 7 9 2 13 3 15 13 9 1 9 13 2
28 3 3 16 3 0 13 7 9 9 13 2 3 3 15 13 3 13 1 9 2 9 13 2 15 10 13 0 2
9 3 3 15 10 9 13 7 13 2
16 9 15 1 9 12 9 13 1 9 2 7 3 15 13 13 2
24 3 15 13 7 13 1 3 9 2 1 3 15 13 9 0 2 0 13 15 15 9 13 9 2
25 9 3 9 2 15 3 15 9 9 13 3 2 3 3 0 9 13 2 15 0 9 0 9 13 2
11 2 2 3 13 2 3 15 0 9 13 2
16 13 3 9 1 9 13 9 13 1 9 2 3 3 3 2 2
7 15 3 13 13 9 9 2
7 15 3 3 13 0 9 2
8 0 3 3 9 0 13 9 2
10 15 3 3 9 13 2 15 3 9 2
17 15 15 3 3 13 1 0 9 2 15 3 13 2 9 0 13 2
19 15 3 1 0 9 13 3 2 15 3 0 13 2 9 16 3 15 13 2
9 3 15 3 3 13 0 9 13 2
8 3 3 0 15 7 9 13 2
12 15 3 9 13 0 2 15 15 9 9 13 2
22 3 3 13 9 2 10 9 2 15 0 1 9 0 13 3 2 9 3 2 12 0 2
9 13 3 15 3 0 3 13 9 2
7 3 3 9 9 0 13 2
30 15 3 3 0 13 9 1 9 7 13 9 12 0 2 15 3 1 13 2 13 15 9 0 2 3 0 2 0 9 2
9 15 3 13 13 1 3 9 2 2
22 3 3 3 9 13 3 9 2 16 0 15 9 0 13 9 3 13 13 3 9 2 2
7 15 3 3 13 0 9 2
10 3 3 3 3 13 0 13 3 9 2
12 1 3 3 0 9 13 0 0 1 0 9 2
30 3 3 3 3 15 9 13 13 1 9 2 15 15 0 13 2 3 9 0 13 2 1 15 9 13 13 9 3 0 2
4 3 3 13 2
17 15 3 13 15 1 9 2 7 3 13 7 15 1 9 13 2 2
17 3 13 13 9 0 2 3 0 2 1 15 3 7 0 13 0 2
11 3 3 9 0 13 13 3 9 13 0 2
10 15 3 13 2 15 3 13 3 3 2
9 0 3 3 15 3 9 13 9 2
8 15 3 3 0 9 13 13 2
10 13 3 1 9 9 2 13 3 9 2
17 15 3 3 9 0 13 13 2 15 3 9 0 13 7 0 13 2
14 15 3 0 13 9 1 9 0 2 0 3 13 9 2
9 7 3 3 15 13 13 7 13 2
9 15 15 3 9 13 13 7 13 2
16 3 3 0 9 13 3 9 1 15 9 0 13 0 1 9 2
6 3 3 15 3 13 2
12 15 9 0 13 7 0 9 7 15 0 13 2
18 7 15 9 9 13 13 2 15 3 15 3 13 2 16 0 3 13 2
7 0 15 13 13 2 13 2
25 3 13 2 13 3 9 9 0 9 2 3 3 3 3 13 2 13 3 13 2 13 3 0 9 2
11 9 3 15 13 9 9 9 13 9 13 2
6 0 3 9 13 13 2
6 3 3 15 9 13 2
19 15 3 9 0 13 2 15 3 1 15 15 13 2 9 3 16 0 13 2
5 10 3 0 13 2
11 3 3 3 0 3 13 7 3 13 9 2
11 3 3 3 13 2 16 15 9 3 13 2
12 9 3 13 9 2 16 3 13 13 0 9 2
16 13 7 9 0 7 9 2 15 3 9 9 7 13 7 13 2
12 15 3 3 0 13 15 13 9 3 9 3 2
13 16 3 15 3 13 2 3 3 3 3 9 13 2
9 3 3 15 0 9 13 9 2 2
12 3 13 13 2 1 3 9 13 9 9 13 2
6 9 3 13 9 0 2
16 3 0 3 0 3 13 2 3 8 15 13 9 9 13 0 2
7 9 3 15 0 13 13 2
6 13 3 3 9 13 2
19 3 3 0 13 9 2 3 3 13 0 2 1 3 13 9 1 9 0 2
17 0 3 3 13 7 13 9 0 9 13 2 9 3 15 0 13 2
9 15 3 9 15 0 1 9 13 2
11 13 0 9 1 9 13 2 0 7 0 2
5 3 3 15 13 2
11 2 3 13 2 15 3 3 13 9 0 2
16 3 3 0 3 13 0 9 2 9 3 13 2 16 9 13 2
28 3 16 0 13 9 7 13 9 2 3 3 3 15 13 9 2 15 3 13 2 7 15 3 13 13 0 9 2
10 3 15 3 13 3 3 13 1 9 2
17 15 3 3 9 13 2 16 13 0 0 9 2 13 3 0 0 2
17 9 0 13 2 13 3 15 13 10 15 3 9 13 7 13 0 2
8 15 3 15 0 9 9 13 2
8 3 3 0 3 0 3 13 2
8 15 3 3 9 13 0 13 2
20 1 3 10 9 0 13 2 0 3 9 13 2 16 9 0 13 9 9 13 2
7 9 3 15 1 9 13 2
8 3 3 0 15 3 9 13 2
23 0 3 16 3 9 13 0 2 13 15 9 2 0 3 13 9 0 9 13 13 1 9 2
16 15 3 9 13 3 13 2 16 3 3 9 13 0 9 13 2
8 0 3 3 9 1 13 2 2
14 15 3 3 3 3 13 1 9 9 0 0 13 9 2
24 7 16 3 0 9 0 13 2 3 13 13 9 0 2 1 3 13 0 9 2 13 3 9 2
16 13 3 9 9 3 3 9 0 13 1 3 9 7 9 0 2
8 13 3 9 2 16 13 9 2
9 13 3 1 9 15 3 13 13 2
9 15 3 3 13 9 9 9 9 2
8 15 15 3 13 13 7 13 2
7 9 3 3 13 15 13 2
6 15 3 0 9 13 2
21 3 3 9 3 1 0 15 13 2 7 3 3 3 13 15 9 7 9 13 0 2
12 0 3 3 0 0 13 2 15 13 9 0 2
9 3 0 3 13 2 16 3 13 2
6 15 3 3 0 13 2
8 3 3 15 3 15 0 13 2
17 13 0 0 13 2 13 1 0 9 2 0 0 0 9 3 13 2
15 9 3 3 0 1 9 9 13 2 3 3 3 0 0 2
13 3 9 13 3 2 3 3 15 13 1 0 13 2
23 3 3 0 13 13 2 3 3 3 9 13 3 13 2 0 9 9 13 2 16 3 13 2
11 3 1 15 13 2 15 3 3 13 13 2
30 16 3 0 9 0 3 0 3 13 13 9 13 13 2 0 3 15 0 0 13 2 13 3 3 3 15 13 1 15 2
6 0 3 15 13 9 2
8 9 3 1 0 15 13 0 2
7 9 15 1 9 13 13 2
21 9 3 3 3 13 2 3 8 3 0 13 2 16 3 15 3 13 0 15 9 2
24 15 3 3 13 9 0 1 15 9 13 2 3 3 1 0 13 2 15 0 13 13 0 2 2
8 15 3 3 9 13 0 13 2
9 3 3 15 13 9 7 0 0 2
19 3 3 15 13 9 0 7 12 9 2 15 3 15 3 7 3 13 9 2
33 13 3 1 9 3 7 1 9 0 9 13 9 3 13 2 16 15 15 13 9 7 9 13 1 9 2 15 3 3 13 9 9 2
20 16 3 3 9 9 7 9 13 2 3 3 3 2 13 3 2 3 13 9 2
37 16 3 3 13 13 3 8 3 13 2 13 3 3 0 1 9 9 9 3 15 13 7 1 9 13 0 3 2 0 13 2 7 9 9 13 2 2
39 3 3 15 3 3 13 1 3 13 2 15 3 13 9 2 15 3 9 0 13 9 2 7 15 13 1 9 13 9 0 2 13 3 9 7 0 0 13 2
8 15 15 3 13 13 7 13 2
26 3 15 3 0 0 7 0 13 0 9 2 3 8 9 0 13 2 7 3 0 3 13 7 0 13 2
16 7 3 15 13 9 0 9 15 13 2 9 3 3 0 13 2
14 3 3 3 9 0 3 3 13 13 9 0 9 9 2
23 3 3 0 9 13 2 0 0 13 3 2 3 3 3 13 9 0 9 13 0 13 2 2
7 15 3 9 9 0 13 2
43 16 3 3 3 9 0 0 13 13 1 9 0 9 0 13 9 13 1 9 2 3 3 15 13 9 2 3 3 13 2 13 2 7 3 3 0 9 13 2 16 0 13 2
7 15 3 3 1 9 13 2
27 3 3 2 9 3 13 1 9 0 2 0 3 13 9 9 7 9 2 15 3 15 1 9 0 13 9 2
19 3 13 2 3 3 13 9 13 1 9 2 13 3 9 3 3 0 2 2
9 3 3 13 2 13 3 9 0 2
17 15 3 3 13 0 1 9 0 2 9 3 1 9 13 0 9 2
15 9 3 3 13 1 9 9 2 9 13 0 9 13 9 2
25 2 13 15 2 10 0 9 13 0 9 7 15 1 9 13 1 0 9 9 13 9 3 13 13 2
25 3 13 13 2 3 3 15 13 9 2 9 13 7 9 7 3 9 2 7 15 13 9 0 13 2
10 3 15 3 0 9 13 3 3 0 2
20 16 3 3 0 3 13 9 7 9 2 3 15 3 3 13 13 2 15 13 2
10 15 3 9 3 0 13 15 15 13 2
18 0 3 3 9 15 0 13 2 15 15 9 0 13 7 3 13 0 2
9 15 3 1 9 9 3 9 13 2
12 13 3 9 0 1 0 9 2 0 7 0 2
13 3 8 3 3 3 9 13 2 16 9 13 9 2
26 13 3 13 1 9 2 0 13 9 2 13 3 3 9 0 1 9 2 9 13 9 3 13 1 9 2
8 15 3 3 9 13 0 13 2
13 13 3 2 3 3 0 9 13 15 13 2 0 2
9 3 3 3 15 13 0 13 2 2
11 13 3 2 7 1 9 9 13 9 3 2
7 9 3 9 1 9 13 2
7 3 3 15 13 0 0 2
8 2 3 3 9 9 15 13 2
19 7 15 1 9 13 9 0 7 10 3 3 3 2 16 3 3 13 3 2
7 0 3 3 13 0 0 2
21 2 15 3 13 2 16 3 3 0 13 0 1 9 1 0 13 13 3 3 9 2
8 3 3 3 3 13 9 15 2
29 1 3 9 9 0 0 13 2 0 0 0 3 13 2 3 1 9 13 2 16 3 9 3 13 3 9 0 13 2
9 0 3 13 9 3 13 2 9 2
7 15 3 9 13 3 13 2
8 12 3 13 7 9 13 0 2
8 1 3 15 9 13 0 9 2
8 12 3 13 9 0 9 9 2
5 0 3 0 13 2
6 15 3 0 0 13 2
16 0 3 15 13 2 3 3 3 9 1 9 13 9 3 13 2
19 13 3 1 9 3 7 1 9 0 9 13 9 0 2 16 3 13 2 2
11 3 3 13 13 0 1 9 0 13 0 2
20 15 3 15 3 13 0 13 3 2 16 3 9 13 2 15 3 0 0 13 2
7 3 13 3 1 0 13 2
8 15 3 3 9 13 0 13 2
35 3 13 3 9 0 15 13 2 16 3 16 3 0 3 0 3 13 2 7 0 13 7 13 13 2 16 3 3 13 1 9 0 13 2 2
11 3 3 13 2 9 3 9 0 9 13 2
26 3 16 3 13 3 13 3 10 9 2 3 3 15 9 1 9 13 2 1 3 15 9 13 0 9 2
8 9 3 1 9 13 9 13 2
23 9 13 1 9 13 3 2 7 3 0 9 13 13 9 2 0 3 1 9 0 13 13 2
6 15 3 15 0 13 2
28 13 3 9 13 3 0 9 2 7 3 9 0 3 13 2 0 3 1 0 9 13 2 15 3 9 0 13 2
13 13 3 1 9 9 2 1 3 0 9 0 13 2
5 9 3 13 0 2
8 13 3 13 1 9 9 0 2
16 3 9 1 0 9 13 2 13 3 13 2 9 3 13 9 2
21 15 3 13 13 1 9 2 3 3 3 3 3 13 2 16 15 9 1 9 13 2
18 3 9 13 9 9 13 9 3 13 2 9 13 7 9 7 3 9 2
9 3 13 2 16 3 13 9 2 2
8 3 3 13 13 9 9 3 2
8 15 3 3 1 9 13 9 2
17 3 16 3 1 9 13 7 9 2 13 3 1 9 9 13 9 2
8 15 3 3 13 0 9 9 2
19 9 3 0 3 3 13 2 3 3 0 9 2 0 3 0 9 13 2 2
10 3 3 13 13 2 15 3 3 13 2
16 15 3 3 0 13 0 1 9 13 2 3 13 9 0 9 2
19 1 3 3 9 9 13 2 13 3 9 2 9 3 1 0 1 3 13 2
7 1 3 3 0 13 9 2
14 15 3 0 13 2 1 3 3 0 13 1 9 13 2
8 9 3 9 13 13 9 13 2
5 15 3 13 13 2
21 9 3 0 0 1 9 13 13 2 1 3 9 13 2 13 3 9 0 0 9 2
16 13 3 9 0 9 2 1 3 9 9 0 0 13 9 13 2
8 15 3 13 1 9 13 9 2
27 13 3 3 9 0 1 9 0 13 9 0 9 2 13 3 0 9 9 2 1 0 3 3 9 9 9 2
10 0 3 3 15 3 7 9 13 9 2
16 1 3 0 9 13 2 3 1 9 0 9 2 15 13 0 2
8 9 3 3 1 9 13 13 2
10 3 9 9 0 13 1 9 13 13 2
8 15 3 13 9 1 9 0 2
31 0 3 13 1 9 7 1 9 2 7 13 9 13 0 2 7 3 13 9 0 13 0 7 0 2 9 3 15 3 13 2
7 9 3 13 9 13 9 2
6 3 0 0 3 13 2
14 15 3 13 2 16 15 9 13 1 9 13 13 2 2
9 3 13 2 1 9 13 0 9 2
10 15 3 3 1 9 9 13 13 3 2
7 3 0 13 3 7 3 2
8 3 3 15 13 9 3 13 2
5 9 3 13 9 2
11 13 3 3 1 9 7 15 1 9 13 2
7 15 3 13 13 0 9 2
10 1 3 3 3 15 0 1 9 13 2
14 16 3 3 13 9 3 15 3 3 2 15 3 13 2
6 15 15 13 13 2 2
13 3 15 9 13 2 3 15 15 13 1 0 9 2
5 13 3 15 3 2
6 3 13 15 3 9 2
13 9 3 10 13 0 13 2 0 3 13 3 2 2
20 3 13 2 7 3 15 9 1 9 13 2 0 3 3 1 9 13 0 9 2
18 16 15 9 13 2 13 9 9 2 0 2 9 3 3 13 0 13 2
8 13 3 3 1 9 13 0 2
14 3 16 13 13 0 1 9 2 9 0 13 0 9 2
25 15 9 3 13 9 2 15 3 13 0 1 9 2 13 3 0 9 9 7 9 0 7 0 9 2
24 9 3 0 1 0 13 9 9 7 9 2 9 3 13 9 0 2 9 3 9 13 0 13 2
30 3 15 13 0 9 13 2 7 15 0 13 9 2 16 9 13 3 9 1 0 13 2 3 3 15 0 9 13 9 2
16 15 3 3 15 9 13 0 0 2 0 13 0 13 1 9 2
9 3 13 2 3 3 0 13 9 2
9 15 3 3 13 9 13 0 9 2
14 13 3 3 2 13 3 15 1 9 3 13 13 9 2
28 9 3 13 7 9 2 15 13 2 1 9 13 1 9 2 1 3 9 13 3 13 2 9 3 13 9 13 2
4 3 13 13 2
5 13 3 0 9 2
21 10 3 3 0 13 2 16 1 9 13 2 15 3 0 3 13 2 0 3 13 2
6 9 3 15 15 13 2
11 13 3 3 15 0 9 2 15 3 13 2
5 3 0 13 2 2
13 3 3 13 2 13 3 9 0 9 9 3 9 2
5 13 3 13 9 2
15 10 3 0 9 1 9 0 9 13 13 1 9 0 9 2
7 1 3 9 0 13 9 2
16 9 3 1 0 13 0 9 2 13 3 0 9 2 0 0 2
12 13 3 3 1 9 13 2 1 3 9 13 2
6 3 0 3 13 9 9
7 15 3 3 13 0 9 2
16 9 3 3 13 13 2 16 13 0 2 9 3 3 13 13 2
4 13 3 15 2
46 3 16 3 9 7 9 13 2 15 3 9 13 13 9 2 3 15 3 2 3 15 3 0 7 0 2 3 13 1 9 7 1 9 13 2 7 1 0 9 7 9 9 13 1 9 2
6 9 3 13 15 2 2
19 3 13 2 9 3 1 9 13 9 13 2 1 15 3 12 9 0 13 2
9 13 3 13 1 9 1 0 0 2
20 2 13 2 15 3 9 13 13 2 13 3 2 1 3 9 0 9 13 0 2
15 15 3 9 9 0 13 2 13 3 9 7 9 0 13 2
12 15 3 1 9 13 3 2 7 13 0 13 2
18 3 3 3 9 13 9 2 7 3 3 13 2 16 3 0 9 2 2
13 3 13 2 15 3 3 15 3 3 13 7 13 2
16 15 3 12 13 1 9 0 2 15 3 3 1 9 3 13 2
6 1 3 13 9 0 2
16 15 3 3 3 7 3 13 9 2 10 3 9 13 1 9 2
15 1 3 15 13 9 12 9 13 2 15 13 1 0 0 2
17 7 15 3 3 13 1 9 0 13 2 0 3 3 9 13 0 2
7 15 3 13 13 0 9 2
6 12 3 3 13 9 2
15 7 15 3 13 1 9 0 2 0 3 3 9 13 0 2
17 3 3 15 13 13 16 9 13 2 16 15 3 3 1 9 13 2
8 13 3 3 0 9 0 2 2
19 3 13 2 15 3 3 15 13 0 9 2 7 0 13 9 2 0 13 2
18 9 3 3 15 3 13 2 15 3 3 0 9 13 2 15 15 13 2
17 7 15 3 3 13 1 9 0 2 0 3 3 13 9 3 13 2
9 0 2 3 3 13 9 9 9 2
13 3 9 13 0 9 2 16 3 9 13 9 2 2
14 3 7 0 13 9 13 2 7 15 13 9 0 13 2
7 13 15 1 3 3 9 2
8 3 3 3 3 0 13 0 2
15 3 13 9 2 16 3 13 0 2 13 9 7 9 0 2
32 13 2 16 13 2 13 3 15 9 13 9 2 16 3 0 13 15 9 13 1 9 13 2 16 3 3 13 7 13 9 9 2
10 15 3 0 15 13 13 15 0 13 2
14 3 3 15 9 1 9 13 2 3 3 9 13 9 2
9 13 3 3 9 13 3 13 9 2
10 3 15 15 9 1 9 0 0 13 2
15 3 3 3 3 0 0 9 13 13 2 16 3 0 13 2
17 3 3 15 0 13 2 16 3 13 9 9 9 1 9 13 2 2
7 15 3 13 13 0 9 2
24 13 3 9 0 9 0 3 9 9 3 9 0 2 15 13 2 3 15 3 13 13 3 9 2
17 0 3 9 13 2 16 3 13 2 13 9 2 15 3 13 2 2
8 15 3 3 13 9 9 9 2
10 13 3 0 0 9 7 9 13 2 2
13 3 3 3 9 13 0 9 13 9 9 0 3 2
18 3 15 3 0 1 0 13 2 9 3 3 9 9 3 9 3 13 2
7 15 3 9 13 7 13 2
5 3 13 9 2 2
9 3 13 9 2 15 3 13 9 2
32 13 3 1 9 9 0 9 3 13 1 9 3 9 3 2 15 3 13 9 0 7 9 9 2 13 3 9 9 7 9 0 2
13 9 3 3 13 13 2 1 3 3 9 9 13 2
5 9 3 13 9 2
9 15 3 1 9 0 13 9 13 2
23 9 3 9 13 2 9 13 2 1 0 9 2 1 0 9 2 9 0 13 0 3 9 2
20 1 3 13 9 9 2 1 3 9 13 1 9 0 2 7 15 1 9 13 2
8 2 3 3 13 1 9 13 2
27 9 3 15 0 15 7 9 13 0 9 2 16 3 3 0 13 9 15 2 7 9 2 15 3 13 0 2
6 3 3 15 13 13 2
6 3 3 9 13 9 2
14 3 3 15 3 13 1 9 2 0 3 13 9 2 2
4 3 13 9 2
7 15 3 3 3 13 9 2
9 9 3 1 9 9 0 9 13 2
20 9 3 3 3 9 13 9 9 13 0 2 16 3 3 13 9 9 9 9 2
20 13 3 15 1 9 9 0 13 2 9 3 9 13 2 9 3 1 9 13 2
12 15 3 3 9 13 0 13 9 3 13 9 2
7 15 3 3 9 0 13 2
12 9 3 3 9 13 3 2 7 13 2 0 2
8 3 13 13 9 9 9 0 2
6 15 3 0 13 9 2
7 9 3 3 9 13 9 2
5 3 13 10 9 2
5 13 3 9 0 2
19 3 3 3 15 0 13 9 0 2 7 3 15 1 9 9 9 13 3 2
9 3 3 15 15 9 1 9 13 2
6 3 3 3 0 13 2
16 3 3 15 3 3 13 13 2 9 13 9 3 13 7 9 2
8 3 3 3 15 0 13 13 2
11 3 13 2 15 3 3 0 3 13 9 2
7 3 3 3 13 9 9 2
16 9 3 3 9 15 7 9 13 0 2 16 15 9 13 0 2
39 16 3 15 9 1 9 13 13 9 9 0 3 2 3 3 15 9 13 3 13 13 3 9 1 9 2 16 15 0 13 2 16 13 9 7 0 13 9 2
8 15 3 3 9 13 9 13 2
9 13 3 0 1 9 13 9 0 2
6 3 0 9 13 2 2
4 3 13 9 2
12 9 3 9 9 0 9 13 2 13 3 9 2
13 15 3 3 9 13 0 2 0 3 3 9 13 2
12 9 3 3 15 9 13 2 9 3 13 9 2
7 15 3 3 13 9 0 2
12 9 3 0 13 9 3 9 3 3 3 9 2
16 9 3 13 2 13 3 9 2 9 3 13 9 0 3 9 2
11 9 3 9 13 2 0 3 13 9 2 2
12 3 13 2 15 3 3 0 1 0 0 13 2
7 2 13 9 0 3 13 2
7 15 3 3 13 9 0 2
17 13 15 9 3 7 9 7 9 0 7 9 1 9 13 0 0 2
31 15 13 3 2 16 13 0 15 13 2 15 3 3 15 13 3 3 13 9 2 15 9 1 0 9 9 13 0 13 2 2
17 3 13 13 9 3 13 2 13 3 1 9 2 15 15 0 13 2
14 9 3 3 0 1 0 13 9 13 2 1 0 13 2
7 3 3 15 13 0 9 2
27 0 3 15 0 9 0 9 2 9 7 9 13 2 3 3 15 9 0 3 3 9 2 7 3 9 9 2
8 0 3 3 15 0 13 13 2
12 3 16 15 15 13 2 15 3 0 0 13 2
17 10 9 1 9 9 13 1 0 13 2 3 3 15 0 13 2 2
4 3 13 9 2
21 15 3 3 13 9 2 7 0 9 13 2 13 3 2 16 3 9 0 9 13 2
17 9 3 3 15 3 13 13 0 3 7 0 2 16 3 0 13 2
19 9 3 3 3 3 0 0 13 2 0 3 3 13 9 7 0 9 13 2
5 0 3 0 13 2
16 9 3 0 13 0 9 2 13 3 9 0 9 0 0 0 2
5 9 3 9 13 2
9 13 3 13 3 1 0 9 0 2
11 15 3 1 9 13 0 9 1 9 0 2
14 3 3 9 13 1 9 2 15 3 15 0 9 13 2
13 9 3 1 9 9 9 13 9 9 0 7 9 2
10 15 1 9 0 9 13 9 0 13 2
8 1 3 13 9 0 3 9 2
14 3 3 13 7 0 2 9 3 0 13 9 1 9 2
26 15 13 9 13 2 13 3 9 2 15 3 3 3 13 0 9 2 3 15 9 13 13 1 9 0 2
14 15 3 9 9 0 7 0 9 13 2 9 9 0 2
6 3 3 9 13 0 2
16 3 3 9 9 13 9 9 2 0 0 2 15 15 9 13 2
29 15 3 3 3 0 9 13 3 0 1 9 13 2 7 3 9 9 0 13 1 9 2 13 3 15 0 1 9 2
8 15 3 13 3 9 13 9 2
12 0 13 0 9 13 9 2 13 3 15 3 2
8 15 3 3 1 0 9 13 2
13 3 3 9 13 2 1 3 3 15 0 9 13 2
14 3 13 1 9 13 9 0 9 2 15 15 13 0 2
20 13 3 1 3 2 0 1 9 13 2 13 3 3 2 1 3 13 9 9 2
24 15 3 16 3 13 0 9 2 13 3 13 3 1 9 0 9 13 1 9 0 7 9 0 2
6 0 3 13 0 9 2
8 0 3 3 15 0 3 13 2
8 3 3 9 13 7 13 9 2
17 3 3 15 0 9 13 9 13 2 7 15 13 13 13 3 9 2
7 13 3 0 9 9 0 2
39 15 3 3 0 13 9 1 9 7 13 9 12 0 2 15 3 1 13 2 13 15 9 0 2 3 0 2 0 9 2 15 3 13 13 1 3 9 2 2
7 13 3 9 13 7 13 2
10 13 3 9 3 2 16 13 9 9 2
10 9 3 13 9 3 13 1 3 13 2
19 3 0 13 13 2 7 3 13 13 2 1 3 9 13 2 9 9 0 2
9 3 3 13 3 15 9 0 13 2
18 15 3 15 0 13 2 7 3 0 13 2 9 3 3 0 13 2 2
16 3 13 2 15 3 3 9 1 9 13 9 13 13 3 9 2
25 3 3 9 3 0 13 13 1 9 9 0 2 15 3 13 13 1 9 2 1 3 13 0 9 2
8 15 3 3 13 0 9 9 2
17 9 3 15 13 0 2 0 3 13 2 0 1 13 13 15 9 2
8 3 15 13 7 13 0 9 2
17 13 3 1 9 9 13 0 0 13 2 1 3 9 0 13 9 2
22 0 3 9 13 2 1 9 13 0 0 0 2 7 1 9 13 2 3 3 9 13 2
10 9 3 13 0 13 2 16 3 13 2
7 3 3 3 3 3 13 2
10 13 3 3 1 9 13 7 9 13 2
19 3 3 3 3 3 13 9 15 0 13 2 7 9 13 7 13 13 3 2
8 15 3 3 13 0 9 9 2
29 2 6 6 2 7 3 3 0 3 13 7 9 2 7 0 13 7 3 3 9 13 9 13 2 16 15 0 13 2
33 3 13 9 3 1 15 13 3 2 13 0 0 9 2 3 3 0 9 0 13 9 2 3 3 3 1 3 13 1 9 3 13 2
9 3 13 9 2 15 3 13 9 2
12 9 3 15 0 0 13 2 0 3 13 9 2
15 13 3 3 1 9 13 7 9 13 2 3 3 15 13 2
8 3 3 13 9 13 0 0 2
5 1 3 9 13 2
30 0 3 15 9 9 13 9 7 9 2 16 3 0 0 13 13 16 13 13 2 15 1 3 3 13 2 13 9 0 2
17 3 16 9 13 7 13 2 0 3 15 3 9 0 13 9 13 2
14 15 3 3 3 13 15 3 0 13 7 0 13 2 2
33 3 3 13 7 1 15 9 13 2 13 0 0 9 2 3 3 0 9 0 13 9 2 3 3 3 1 3 13 1 9 3 13 2
10 9 3 13 9 3 13 1 3 13 2
18 3 3 3 15 3 0 13 0 9 0 3 9 9 3 13 7 9 2
8 3 0 13 3 9 0 2 2
6 15 3 0 13 13 2
11 3 3 13 13 2 0 3 9 0 13 2
6 9 3 13 3 0 2
10 1 3 0 1 15 9 13 0 9 2
17 3 16 3 3 1 9 13 7 3 9 2 13 15 9 13 0 2
6 13 3 15 9 13 2
18 0 3 13 9 13 2 16 3 13 3 3 3 7 15 9 0 13 2
7 7 3 9 13 7 9 2
9 13 16 15 9 9 3 13 2 2
8 15 3 3 13 9 9 9 2
10 13 3 0 0 9 7 9 13 2 2
13 3 3 3 9 13 0 9 13 9 9 0 3 2
15 3 16 3 15 3 9 0 13 2 3 15 9 13 13 2
18 2 3 3 3 15 0 15 2 0 0 13 13 0 9 1 0 9 2
9 13 3 16 15 13 13 0 9 2
13 10 3 0 3 15 13 13 15 3 0 3 13 2
10 15 3 2 3 13 3 2 9 13 2
22 16 3 1 15 3 9 13 9 0 2 13 0 9 7 9 13 9 3 1 15 13 2
10 3 15 3 9 9 3 9 3 13 2
7 3 13 9 0 13 9 2
33 15 3 16 13 3 3 13 0 2 13 3 1 9 0 9 13 2 7 13 13 9 3 7 9 3 3 3 9 9 7 9 13 2
16 3 3 3 13 13 9 9 2 16 3 9 0 13 13 3 2
17 2 13 9 9 3 2 16 15 13 13 9 2 3 13 3 3 2
5 3 15 9 13 2
17 0 3 3 0 2 0 9 0 2 3 13 15 13 9 7 9 2
7 3 13 13 9 3 13 2
10 13 3 1 9 13 2 3 3 13 2
10 1 3 3 3 10 9 13 0 9 2
15 9 3 3 9 1 9 13 2 13 3 7 3 9 9 2
14 3 15 3 3 3 13 13 2 0 3 13 0 9 2
9 3 15 9 0 13 2 13 3 2
5 13 3 3 0 2
6 15 3 3 9 13 2
4 3 0 13 2
10 3 9 3 3 16 3 13 0 13 2
13 3 3 3 15 13 13 2 13 1 9 9 9 2
14 3 3 2 9 3 13 9 2 16 13 13 0 9 2
9 3 13 9 2 15 3 13 9 2
22 15 3 9 3 9 1 9 13 2 9 3 9 13 0 2 13 3 3 0 13 9 2
19 15 3 16 3 13 3 13 3 0 13 9 2 15 3 13 13 9 9 2
9 3 3 9 13 9 15 3 13 2
38 3 3 15 13 9 0 2 16 1 15 9 7 9 13 2 7 15 3 13 9 2 0 3 13 1 0 9 2 7 3 15 13 9 3 9 3 2 2
16 3 13 2 15 3 3 0 3 13 2 13 16 9 0 13 2
10 9 3 13 9 3 13 1 3 13 2
22 3 13 15 0 0 1 15 13 2 3 3 15 9 13 2 3 13 9 0 7 9 2
21 9 15 13 0 2 15 3 3 0 13 2 15 3 15 3 13 3 3 0 13 2
14 15 3 16 9 13 9 2 13 0 13 9 1 9 2
20 9 3 9 13 2 1 9 3 3 13 13 2 1 9 0 9 9 3 13 2
12 15 3 9 15 13 13 0 9 13 0 9 2
16 1 15 9 7 9 9 13 2 15 3 0 0 0 13 9 2
13 3 3 15 0 9 13 2 16 3 10 9 13 2
6 3 3 3 15 13 2
13 3 0 13 3 2 3 3 13 1 9 0 2 2
7 15 3 3 13 0 9 2
25 13 2 16 3 10 9 9 0 9 13 9 3 9 3 0 13 2 3 15 13 7 0 13 9 2
10 3 3 0 3 0 3 1 9 13 2
21 3 3 15 15 15 3 1 9 13 3 13 2 16 3 3 3 3 3 13 2 2
4 3 3 13 2
16 3 0 15 0 9 13 13 3 13 9 2 1 3 13 9 2
11 3 13 2 15 3 3 9 0 13 2 2
7 15 3 3 13 0 9 2
6 15 3 9 0 13 2
18 0 3 9 3 3 0 7 0 2 9 3 1 0 9 13 13 9 2
10 3 3 15 13 9 0 2 16 13 2
10 3 3 13 2 15 3 3 13 13 2
8 15 3 3 9 13 9 13 2
18 15 3 15 15 0 13 2 16 3 13 3 3 9 13 15 9 13 2
10 9 3 9 13 0 2 3 3 15 2
8 15 3 9 13 1 9 2 2
7 15 3 13 3 3 13 2
7 9 3 9 13 13 9 2
8 9 3 3 0 13 1 9 2
7 3 3 15 13 0 0 2
26 3 3 15 1 9 9 0 13 0 1 9 2 15 13 2 16 3 9 15 13 7 0 9 0 2 2
20 3 13 2 3 2 15 13 13 0 1 9 2 13 2 16 0 13 1 9 2
6 9 3 3 13 13 2
17 3 3 3 0 13 16 15 3 0 3 13 3 13 2 13 9 2
5 9 3 0 13 2
18 6 3 0 0 2 0 1 9 13 2 9 9 3 9 3 0 13 2
17 3 3 3 3 15 15 13 13 0 1 9 2 16 0 13 2 2
14 10 3 9 13 1 9 9 1 9 9 0 13 13 2
7 1 3 13 13 9 9 2
17 3 3 13 2 15 3 0 13 9 2 13 3 9 9 3 13 2
16 9 3 1 9 9 13 3 2 13 3 3 3 9 0 9 2
19 13 3 1 9 9 9 9 0 2 15 3 13 9 2 1 3 13 0 2
13 13 3 1 9 13 2 3 3 13 2 13 9 2
20 15 3 3 9 13 3 13 2 13 3 7 3 2 16 9 9 13 13 9 2
8 3 15 13 13 1 0 0 2
9 2 3 15 9 7 0 13 9 2
27 7 3 3 3 0 3 0 3 13 7 15 3 13 13 2 16 1 9 13 3 7 3 0 0 9 2 2
15 2 6 3 3 0 9 13 7 0 3 0 13 13 2 2
5 3 3 13 9 2
42 3 0 9 2 3 16 0 9 13 7 13 3 2 7 16 9 9 13 7 9 3 13 0 1 9 9 2 13 3 0 9 9 2 3 3 1 9 13 0 9 9 2
7 0 3 9 13 13 9 2
10 15 3 1 0 13 2 9 0 9 2
13 9 3 3 9 13 0 2 0 3 3 9 13 2
7 9 3 0 13 9 13 2
8 13 3 3 3 0 0 9 2
11 13 3 0 9 2 15 15 13 9 0 2
14 10 3 0 0 1 9 13 2 15 3 13 0 13 2
37 15 3 1 9 13 13 9 9 3 2 3 1 9 13 2 13 3 9 3 13 2 9 3 3 13 0 0 9 2 1 3 3 13 3 9 0 2
5 15 3 9 13 2
13 3 15 9 0 13 2 3 3 15 9 13 13 2
6 13 7 1 9 13 2
8 2 0 3 3 9 0 13 2
25 3 3 9 0 2 15 3 3 15 13 9 2 13 2 16 3 13 2 13 3 15 9 9 2 2
8 13 7 1 9 13 0 9 2
21 3 3 15 0 9 13 13 2 0 0 2 7 3 1 9 13 2 16 13 9 2
8 9 3 15 3 1 9 13 2
25 15 3 13 1 9 9 0 1 0 2 3 16 3 0 13 2 15 13 9 3 0 7 9 0 2
17 15 3 9 1 9 13 13 9 2 3 3 0 1 9 13 9 2
21 13 3 3 2 9 3 15 13 9 13 2 3 3 9 1 9 0 13 9 0 2
7 9 3 9 3 0 13 2
6 13 3 9 0 9 2
5 3 9 0 13 2
13 3 3 3 3 9 13 15 0 0 9 1 9 2
7 3 15 3 9 13 2 2
12 13 0 9 2 16 3 13 3 13 9 13 2
9 15 3 3 3 13 13 0 9 2
9 3 15 3 0 9 9 13 2 2
12 3 13 2 15 3 3 0 1 0 9 13 2
8 13 3 0 3 13 0 9 2
7 9 3 15 0 13 13 2
34 3 15 3 13 1 9 2 0 15 13 7 13 1 9 2 9 3 13 0 0 2 9 3 9 3 13 2 1 15 3 0 9 13 2
9 15 3 3 3 13 13 0 9 2
16 3 15 13 3 7 13 7 13 2 15 3 9 7 9 13 2
9 3 15 3 13 13 0 9 2 2
12 3 13 2 15 3 3 13 9 7 0 9 2
7 15 3 9 13 0 3 2
4 3 13 9 2
9 9 3 13 7 13 9 9 0 2
25 1 3 0 0 13 0 2 16 3 15 9 13 7 9 2 13 3 1 9 2 9 3 3 13 2
10 3 3 3 0 9 3 0 13 2 2
18 3 3 13 13 9 0 0 2 3 0 2 13 3 1 0 0 13 2
23 1 3 3 9 9 13 3 2 0 3 9 13 13 2 1 3 9 13 3 7 9 0 2
15 15 3 9 13 9 9 13 2 9 3 9 0 13 13 2
6 1 9 3 13 9 2
19 9 3 9 13 0 0 13 2 13 3 9 0 2 16 3 15 13 9 2
17 3 3 15 13 9 3 13 0 9 9 1 2 1 3 9 13 2
10 13 3 13 2 9 3 13 0 9 2
11 9 3 13 2 13 0 9 3 1 9 2
17 1 3 13 16 15 0 9 13 0 7 13 9 13 7 0 13 2
18 13 3 13 2 3 3 3 0 9 13 2 3 3 13 9 0 13 2
7 15 3 13 13 0 9 2
18 2 13 13 2 16 15 13 13 9 2 16 15 13 9 0 13 2 2
20 3 13 2 9 3 0 13 9 2 13 3 13 3 2 3 15 0 9 13 2
15 3 9 3 9 13 2 9 3 12 7 9 9 0 0 2
19 13 3 13 2 3 3 3 0 9 13 2 0 3 0 1 9 13 9 2
16 3 3 3 10 9 13 9 0 2 13 3 1 9 0 0 2
11 3 9 9 3 3 0 1 9 13 13 2
5 15 3 0 13 2
44 3 16 13 9 13 9 2 9 3 1 9 0 9 13 13 2 1 9 13 2 0 3 1 9 9 13 0 2 9 3 1 0 9 0 13 2 9 2 0 3 9 3 13 2
8 13 3 0 9 12 13 9 2
25 9 3 15 13 0 1 9 2 0 3 1 9 0 9 13 9 1 9 2 9 3 13 3 13 2
11 15 3 9 13 13 0 9 13 1 0 2
6 0 3 0 13 9 2
9 15 3 9 13 2 9 0 13 2
10 3 3 3 0 9 3 0 13 2 2
12 7 3 9 0 13 9 2 15 3 0 13 2
10 3 3 2 15 9 13 13 1 9 2
15 3 12 3 9 13 2 0 3 9 7 0 9 0 0 2
11 13 3 13 2 3 3 3 13 9 13 2
19 3 3 9 13 9 7 0 9 2 16 13 13 9 9 3 9 0 13 2
6 0 3 0 13 9 2
7 3 3 9 9 0 13 2
8 15 3 3 9 13 0 13 2
6 15 3 9 13 0 2
12 13 3 0 9 2 3 3 9 13 3 13 2
34 15 3 15 0 13 2 7 15 13 2 16 3 0 3 13 2 7 15 3 13 2 16 9 13 0 2 0 0 13 0 1 9 2 2
7 15 3 13 13 0 9 2
16 2 3 3 15 7 9 9 0 13 1 9 2 3 3 13 2
18 3 3 15 3 9 9 1 9 13 2 15 3 13 3 1 9 13 2
11 3 3 3 3 13 2 9 3 13 9 2
22 3 3 15 3 9 1 9 9 13 13 0 2 3 13 9 9 9 1 9 13 2 2
11 3 15 3 3 13 2 13 0 1 9 2
17 15 3 1 9 13 2 9 13 0 2 13 1 9 0 2 0 2
20 3 9 13 13 2 15 3 1 9 9 2 15 3 1 9 0 3 7 0 2
9 15 3 9 13 13 7 9 13 2
6 9 3 15 13 2 2
8 3 13 2 13 0 13 9 2
7 9 3 3 13 1 9 2
8 3 3 0 3 9 13 13 2
6 0 3 0 9 13 2
15 3 13 2 9 3 13 3 3 2 13 3 9 0 9 2
18 3 3 3 2 16 0 3 9 7 9 13 2 1 9 13 0 13 2
13 0 3 0 1 9 9 13 13 2 9 0 3 2
20 9 3 13 9 9 2 9 3 7 9 9 3 2 9 3 9 9 3 0 2
16 15 3 9 9 13 3 0 2 0 3 13 1 3 9 13 2
9 15 3 3 13 9 7 0 9 2
9 15 3 9 13 2 9 0 13 2
18 3 3 15 9 3 13 0 9 13 2 15 3 0 13 1 0 9 2
27 3 3 3 3 0 13 9 0 2 7 3 10 12 0 13 2 16 3 3 9 13 9 13 7 9 13 2
13 3 13 2 15 3 3 0 13 7 13 2 13 2
16 3 16 3 9 13 9 2 15 3 3 9 13 0 0 9 2
13 3 13 2 15 3 3 0 13 0 9 3 13 2
21 9 3 9 2 9 3 3 9 2 9 3 9 2 9 3 3 13 9 9 9 2
16 15 3 3 3 0 3 13 0 9 2 9 3 13 9 3 2
11 15 3 3 13 2 9 3 1 9 13 2
8 3 3 9 13 0 9 13 2
7 15 3 0 0 13 9 2
14 15 0 3 9 0 9 13 2 0 3 9 3 13 2
8 0 3 1 9 9 13 9 2
16 9 3 3 9 13 9 1 9 3 2 0 3 9 13 9 2
10 9 3 9 1 9 9 0 9 13 2
8 15 3 13 2 13 3 3 2
15 15 3 3 1 9 0 0 2 9 1 9 13 0 9 2
15 3 3 9 13 0 9 2 9 3 9 2 9 3 9 2
15 9 3 3 3 9 9 9 13 1 9 2 13 3 13 2
6 13 3 9 9 9 2
8 3 9 13 9 3 9 0 2
14 9 3 9 9 13 9 0 9 2 3 3 9 13 2
10 13 3 0 2 9 3 13 0 9 2
10 3 3 9 0 9 13 3 1 9 2
5 15 3 9 13 2
9 15 3 13 1 9 9 3 0 2
6 13 3 3 9 9 2
10 3 3 15 9 13 1 9 13 3 2
14 15 3 9 13 0 9 13 2 9 3 0 9 13 2
15 3 3 3 15 13 9 1 9 13 3 3 15 13 0 2
11 3 3 0 13 9 2 15 0 3 13 2
9 3 15 3 13 0 1 9 13 2
7 3 3 9 0 9 13 2
17 3 15 1 15 9 0 13 13 2 16 3 13 9 3 0 2 2
9 15 3 3 3 13 13 0 9 2
33 2 16 3 3 1 15 9 13 13 2 3 3 13 13 1 9 3 15 9 9 0 13 2 15 3 9 3 0 13 7 9 13 2
9 3 3 3 9 3 0 13 2 2
16 3 3 13 9 13 9 0 13 2 15 3 9 13 3 13 2
8 15 15 3 1 9 0 13 2
9 13 3 3 15 3 9 9 13 2
11 13 3 1 9 13 9 0 3 1 9 2
33 3 3 9 13 2 7 13 9 9 0 1 9 0 13 13 2 3 3 0 9 9 3 9 1 9 13 2 7 9 13 13 9 2
13 3 3 15 13 13 0 13 2 9 13 9 9 2
28 3 3 15 9 0 13 3 1 9 7 9 0 2 0 3 3 9 13 13 9 2 7 15 13 9 0 13 2
18 0 15 3 9 13 2 16 3 9 13 2 15 3 9 7 9 13 2
13 0 3 13 2 9 3 15 1 9 9 0 13 2
8 13 3 15 13 7 3 9 2
5 3 15 13 13 2
18 3 13 2 15 3 13 0 9 9 2 3 3 0 9 13 3 13 2
10 2 13 3 3 15 0 0 13 9 2
33 3 9 9 13 2 15 3 15 3 9 1 0 13 9 13 2 16 3 3 15 13 9 7 9 2 7 15 13 13 1 9 2 2
10 3 13 2 15 3 13 9 13 13 2
17 13 3 13 1 9 2 1 3 9 13 9 0 2 13 9 0 2
25 3 3 1 9 13 2 3 3 13 9 9 3 3 3 13 13 9 2 7 15 13 9 0 13 2
7 15 3 13 13 0 9 2
27 2 13 2 16 3 15 0 13 7 13 2 16 13 1 9 2 3 13 3 0 2 16 9 9 0 0 2
27 3 13 9 13 3 1 9 1 9 2 15 3 7 0 9 2 16 3 15 1 9 13 15 15 13 2 2
27 3 13 2 15 3 1 13 9 13 2 13 3 3 15 3 9 0 1 9 2 3 13 2 9 13 3 2
18 13 3 9 1 0 9 2 16 15 3 9 0 13 2 13 9 0 2
28 15 3 13 3 0 1 9 7 9 13 0 2 3 9 2 15 3 9 0 1 9 0 3 9 9 13 0 2
11 15 3 3 0 9 9 13 1 9 13 2
8 15 3 3 9 13 13 9 2
8 3 3 3 9 1 0 13 2
7 3 3 9 13 0 9 2
16 3 13 2 9 3 0 13 9 2 13 3 9 13 9 9 2
2 13 2
10 13 15 9 0 2 16 15 13 2 2
21 3 3 13 2 15 3 0 13 9 2 13 3 9 9 3 13 2 13 3 13 2
5 3 9 3 13 2
22 13 3 9 1 13 9 2 9 7 9 13 3 9 2 15 3 3 13 9 13 0 2
18 0 3 3 15 9 3 9 3 3 0 13 2 0 3 1 9 13 2
8 3 9 13 9 7 9 3 2
20 15 3 16 3 9 3 7 0 13 9 2 13 3 13 2 16 0 13 9 2
15 3 9 13 7 13 13 3 2 7 15 13 9 0 13 2
9 15 3 9 13 9 7 0 9 2
18 3 15 3 13 0 9 2 3 0 3 3 3 0 2 15 15 13 2
7 3 3 9 0 9 13 2
19 3 3 15 15 9 1 9 13 2 15 3 15 13 7 15 9 13 2 2
8 15 3 3 13 0 9 9 2
15 15 12 0 9 13 2 3 3 15 13 3 3 0 9 2
16 9 3 0 3 13 2 3 3 15 9 13 13 1 9 9 2
17 3 3 15 13 9 0 13 0 9 2 15 15 9 9 13 2 2
14 15 3 3 13 9 13 2 15 3 3 0 13 2 2
16 2 3 3 13 2 9 3 1 9 13 13 9 7 13 13 2
14 3 15 9 7 9 7 9 1 15 13 9 0 13 2
9 2 13 3 9 13 7 13 9 2
12 3 3 9 0 7 9 9 7 9 0 13 2
44 3 16 3 0 9 13 2 9 13 0 9 2 1 3 9 7 0 9 9 2 13 9 0 2 1 15 3 0 9 13 7 13 9 2 15 3 1 9 13 13 3 3 2 2
19 2 3 13 2 10 3 9 0 13 0 2 3 13 2 0 1 9 13 2
19 0 3 3 9 13 13 2 1 3 3 1 9 13 0 9 2 0 13 2
6 13 3 9 0 13 2
6 15 3 13 3 9 2
12 3 3 9 0 7 9 9 7 9 0 13 2
13 3 9 7 9 7 9 9 9 3 0 9 13 2
30 3 16 0 9 13 2 9 3 13 0 9 2 1 3 9 7 0 9 9 2 13 1 9 2 3 3 3 13 13 2
7 15 3 9 13 13 13 2
27 2 3 3 3 0 9 1 9 13 15 2 15 3 0 9 1 9 13 9 3 0 1 3 9 13 2 2
23 3 3 13 2 7 9 9 0 9 13 0 13 9 2 3 13 2 16 15 9 9 13 2
10 13 3 9 3 3 3 15 3 3 2
10 1 3 9 13 1 9 3 7 9 2
28 15 3 1 3 9 3 7 9 0 9 13 2 9 3 13 2 9 0 13 2 9 3 7 9 13 13 9 2
17 15 3 3 13 9 3 9 3 1 9 3 13 2 13 3 9 2
8 3 15 3 13 0 9 9 2
10 15 3 9 13 3 13 1 0 9 2
9 0 3 13 9 1 9 13 2 2
8 15 3 3 13 0 9 9 2
21 3 3 15 9 3 9 3 9 13 2 3 3 3 9 13 0 9 13 1 9 2
6 0 3 3 13 2 2
7 15 3 13 13 0 9 2
10 2 9 3 15 0 1 9 13 2 2
17 3 13 2 3 3 13 0 9 9 2 13 3 3 9 7 9 2
10 3 9 3 13 9 7 9 7 9 2
14 9 3 3 13 1 9 0 9 13 9 7 13 13 2
10 15 3 13 1 9 9 1 9 13 2
19 15 3 3 13 7 13 9 2 7 13 13 9 3 7 9 9 3 13 2
15 15 3 0 9 13 9 7 9 2 13 3 3 9 0 2
14 9 3 1 9 13 13 2 9 13 0 9 3 13 2
8 9 3 13 2 9 3 13 2
11 13 3 3 1 9 7 15 1 9 13 2
10 13 9 7 9 13 2 3 3 13 2
18 9 3 13 0 2 15 3 0 9 13 7 9 13 13 3 9 2 2
7 15 3 3 13 0 9 2
5 15 15 3 13 2
6 3 3 9 0 13 2
23 3 15 13 0 9 13 0 3 13 7 1 9 15 13 0 2 15 15 13 0 9 13 2
15 3 3 3 15 13 2 1 15 9 13 13 9 3 0 2
9 3 3 3 13 7 3 13 3 2
32 16 3 15 15 0 3 9 2 15 15 13 2 0 13 13 7 1 9 13 2 3 3 3 3 15 15 13 13 3 1 9 2
8 15 3 0 3 9 13 2 2
8 15 3 3 13 0 9 9 2
22 9 3 3 15 3 13 3 13 2 7 9 9 9 13 2 16 9 13 9 9 2 2
19 3 13 2 15 3 13 7 1 9 13 9 13 2 9 3 1 9 13 2
7 7 15 13 9 0 13 2
8 15 3 3 13 0 9 9 2
13 2 3 13 2 3 13 2 7 9 0 13 13 2
7 15 3 3 9 13 13 2
8 13 3 9 1 13 9 13 2
13 15 3 15 1 2 0 9 13 2 13 1 0 2
5 13 3 9 13 2
6 15 3 15 13 13 2
16 3 13 2 16 15 9 13 0 0 9 2 16 0 0 13 2
8 3 3 3 15 0 9 13 2
15 13 3 0 0 0 2 13 3 7 15 7 9 1 9 2
7 15 3 3 13 0 9 2
20 13 3 16 3 0 1 9 13 0 2 3 3 15 3 7 9 2 15 13 2
24 3 3 13 15 9 0 2 3 13 2 7 15 0 13 9 0 2 9 13 0 7 0 9 2
6 3 1 9 13 0 2
12 3 9 13 3 9 9 2 13 3 0 2 2
8 15 3 13 3 0 9 9 2
10 15 13 13 2 13 3 15 0 13 2
13 3 15 15 13 1 9 9 3 13 13 9 9 2
3 3 13 2
17 3 15 15 13 0 2 16 3 15 13 2 13 15 0 9 2 2
7 15 3 13 3 0 9 2
18 3 3 13 1 9 0 2 16 13 9 9 13 2 7 15 13 2 2
5 3 13 13 9 2
20 0 3 15 9 13 2 7 3 0 9 13 2 7 13 13 9 7 9 13 2
22 15 3 16 13 7 13 0 9 2 13 3 9 0 2 1 9 9 2 9 10 0 2
22 15 3 3 1 9 0 13 3 13 2 13 16 15 15 13 0 9 2 16 13 9 2
12 15 3 3 3 13 2 9 3 15 9 13 2
16 9 3 3 3 15 3 13 2 3 3 13 0 9 9 13 2
24 3 3 3 0 3 3 9 13 9 9 13 2 15 15 0 0 13 13 0 9 1 0 9 2
9 15 3 3 9 0 13 9 2 2
7 15 3 3 13 0 9 2
18 16 3 0 3 13 9 7 9 13 2 3 3 15 13 0 3 0 2
15 13 3 15 9 2 15 3 3 15 13 13 1 0 2 2
16 3 13 2 13 3 0 0 9 2 3 3 9 9 0 13 2
6 3 3 13 3 0 2
21 3 3 16 13 2 0 3 9 9 13 2 3 13 15 7 3 3 13 15 13 2
8 15 3 13 16 3 0 13 2
25 3 3 15 3 9 9 13 1 9 2 15 3 0 13 9 3 2 13 9 3 13 7 0 9 2
13 15 3 9 9 13 2 15 0 0 9 1 9 2
7 15 3 15 13 13 2 2
8 15 3 3 9 13 9 13 2
20 0 3 0 9 1 9 13 13 2 3 3 3 15 15 0 9 13 0 9 2
19 15 3 13 3 13 2 3 3 15 13 9 13 2 0 9 3 13 2 2
16 0 3 3 13 7 13 9 2 9 3 1 9 13 9 13 2
29 3 0 9 13 9 0 15 13 0 9 2 16 3 15 13 9 13 3 13 2 7 1 9 13 2 7 15 13 2
21 3 3 9 0 9 1 9 13 9 9 2 3 3 15 13 3 9 1 0 0 2
11 3 3 3 13 15 3 9 0 13 2 2
20 10 3 13 0 9 9 0 2 1 3 15 9 13 9 3 0 7 0 9 2
12 15 3 0 9 13 9 9 13 9 3 9 2
8 3 3 15 13 9 3 13 2
9 2 3 3 3 15 13 0 9 2
22 3 9 0 0 1 9 9 9 13 7 13 9 2 1 3 15 9 0 13 7 9 2
13 3 1 9 9 0 13 9 0 3 13 7 0 2
11 1 3 9 0 13 9 2 0 9 0 2
10 3 3 15 13 9 9 3 7 9 2
8 1 3 9 13 9 0 0 2
21 3 3 3 1 3 13 1 9 3 13 2 9 0 9 2 7 15 1 9 13 2
24 3 3 3 0 3 3 9 13 9 9 13 2 15 15 0 0 13 13 0 9 1 0 9 2
7 15 3 3 13 0 9 2
6 3 3 13 9 13 2
8 3 9 13 9 13 0 13 2
7 15 3 15 3 13 9 2
20 0 3 3 13 3 3 13 2 16 3 9 0 13 3 13 13 0 1 9 2
24 9 3 3 3 15 0 9 2 3 3 3 13 2 3 13 2 16 0 9 13 1 9 0 2
9 15 3 15 13 3 3 15 0 2
10 9 13 0 9 9 1 2 0 13 2
6 0 3 13 3 9 2
26 15 3 15 13 9 13 2 16 13 2 0 9 2 7 3 3 13 2 0 3 13 9 2 3 13 2
32 7 3 3 13 9 0 9 2 9 3 1 9 13 13 9 3 7 3 2 7 1 9 13 2 9 13 2 13 3 0 9 2
18 1 3 15 13 9 13 2 16 13 2 13 9 3 7 9 7 9 2
8 1 3 13 9 9 9 0 2
6 3 15 15 9 13 2
20 3 13 2 15 3 3 13 9 7 0 9 2 9 13 15 15 0 13 9 2
19 13 3 3 3 13 2 1 3 9 9 13 9 2 9 3 13 7 13 2
18 9 3 13 9 2 15 15 13 1 0 13 9 13 7 9 9 13 2
22 3 3 3 15 15 13 3 3 13 2 16 15 3 10 0 2 16 13 2 3 13 2
16 3 3 15 9 1 9 0 13 16 15 15 9 13 9 13 2
6 0 3 0 9 13 2
10 15 3 3 3 13 9 13 9 0 2
18 10 3 9 3 3 0 13 9 0 2 1 15 0 3 15 13 9 2
12 3 13 2 15 3 3 3 1 9 13 9 2
9 13 3 13 9 0 2 0 13 2
17 3 3 15 0 13 9 13 2 9 3 3 3 3 13 9 0 2
22 3 3 15 9 13 9 9 15 16 3 13 9 9 1 2 9 9 13 7 15 0 2
7 15 3 3 13 0 9 2
27 2 9 3 3 15 3 3 13 16 9 0 13 2 16 3 15 9 13 13 9 0 7 0 1 0 9 2
7 15 3 13 13 0 9 2
7 3 15 13 3 3 13 2
6 3 3 15 9 13 2
20 3 3 3 15 3 13 9 0 2 3 3 0 9 2 15 3 9 9 13 2
12 9 3 15 15 13 0 2 3 3 15 13 2
20 9 3 15 1 9 0 0 3 0 13 2 15 3 15 13 9 1 0 13 2
6 3 3 9 0 13 2
8 15 3 15 13 0 13 2 2
7 15 3 3 13 0 9 2
8 3 15 3 0 1 0 13 2
16 3 3 3 9 3 7 9 13 9 9 0 2 9 1 13 2
27 3 16 13 0 9 13 2 9 3 13 3 3 13 2 15 3 9 9 13 13 3 2 9 1 9 13 2
7 1 9 3 13 3 13 2
9 15 3 3 0 9 0 9 13 2
17 3 10 0 9 0 9 13 9 0 3 0 13 13 2 3 13 2
17 15 3 3 13 13 2 3 3 15 9 13 1 9 16 13 0 2
16 13 3 16 0 9 13 2 3 3 13 1 9 9 0 9 2
38 7 9 13 9 9 3 2 7 16 1 9 9 13 0 2 9 13 0 9 2 9 9 2 7 13 0 9 9 3 2 15 15 13 7 13 0 13 2
17 0 3 0 13 9 2 16 15 0 9 0 13 2 13 9 9 2
28 16 3 3 9 13 0 1 9 9 0 9 13 7 3 9 2 3 1 9 0 9 13 2 16 9 9 13 2
13 13 3 9 9 1 0 2 9 3 1 9 13 2
14 3 15 9 9 7 9 0 13 13 0 1 0 9 2
44 3 3 7 0 0 13 9 2 9 3 15 15 13 2 13 1 9 2 9 3 15 15 9 0 13 2 0 3 0 15 13 2 0 3 0 13 2 1 15 3 0 13 9 2
18 3 3 3 3 15 0 9 13 2 13 9 0 2 15 15 3 13 2
15 3 3 9 13 1 9 13 9 9 2 15 13 1 9 2
17 1 9 13 1 0 9 13 2 3 3 15 13 3 3 13 2 2
25 13 3 7 1 9 13 9 0 2 13 3 9 7 9 7 9 2 0 3 9 13 0 9 13 2
18 15 3 15 3 13 2 13 3 9 2 13 3 9 2 1 3 13 2
4 13 3 9 2
17 3 3 9 13 1 9 2 15 3 3 9 9 13 3 13 9 2
8 9 3 9 0 13 9 9 2
10 15 3 13 13 2 15 3 13 13 2
29 3 3 16 9 9 9 0 13 13 2 16 3 15 13 9 1 9 2 1 3 0 13 2 3 15 13 3 13 2
10 13 3 3 15 9 0 1 0 9 2
19 1 3 13 9 3 9 7 9 9 2 7 1 9 9 7 9 9 13 2
9 0 3 13 1 9 9 9 13 2
16 1 3 0 13 2 0 1 0 9 1 9 13 7 9 13 2
6 15 0 9 13 9 2
19 3 3 3 3 15 3 13 13 9 0 2 15 3 15 13 15 3 13 2
17 7 13 9 13 2 15 3 13 2 9 1 9 9 7 9 13 2
18 3 3 15 9 3 13 9 2 7 3 3 0 9 0 9 13 3 2
10 3 3 3 15 0 9 13 13 2 2
7 15 3 3 9 13 9 2
12 15 3 1 9 9 13 0 3 2 13 9 2
6 15 3 0 9 13 2
13 3 3 3 3 13 9 2 16 3 9 9 13 2
22 3 16 15 1 9 13 1 9 2 13 1 9 2 13 9 0 9 3 0 7 9 2
11 9 3 1 9 13 1 0 0 9 13 2
14 9 3 1 9 13 0 2 1 3 9 13 0 0 2
7 15 15 0 13 7 13 2
15 9 1 9 15 1 0 0 13 2 0 9 13 13 2 2
16 1 3 15 13 9 0 9 0 13 2 1 3 0 9 13 2
9 9 3 12 0 13 9 0 13 2
9 3 3 3 15 0 3 13 0 2
6 0 3 13 9 0 2
17 0 3 13 9 2 0 3 15 1 9 13 3 0 7 0 9 2
13 13 3 1 3 9 9 7 9 0 7 9 0 2
6 13 3 9 0 9 2
11 9 3 9 13 13 2 9 3 0 9 2
37 1 0 3 3 0 7 0 9 13 0 0 9 9 9 1 13 2 1 0 9 2 16 3 0 1 9 9 13 15 15 3 13 7 15 3 13 2
13 9 3 13 9 0 9 13 0 1 9 9 0 2
20 3 3 0 9 9 13 9 2 16 3 3 13 9 13 3 0 7 13 9 2
6 3 3 0 13 9 2
16 1 9 3 15 9 13 0 9 9 1 9 7 0 9 2 2
31 3 15 3 0 1 0 13 2 0 3 15 13 9 9 2 9 9 13 9 13 2 15 3 3 13 3 13 2 16 13 2
9 9 3 15 13 9 1 9 13 2
6 15 0 9 13 9 2
11 3 3 3 3 13 13 1 9 9 0 2
14 3 15 1 9 9 13 2 13 0 9 7 9 0 2
21 3 3 0 9 13 1 9 9 13 7 9 9 0 2 7 1 9 13 7 9 2
4 13 15 13 2
6 9 3 15 13 13 2
22 3 3 13 16 3 13 0 9 2 13 9 1 0 9 9 1 3 13 0 1 9 2
15 9 3 3 0 0 13 0 9 2 9 13 9 0 2 2
7 15 3 3 9 13 9 2
6 13 9 3 13 9 2
26 15 3 3 3 13 0 9 3 3 13 2 15 13 9 7 9 0 2 7 9 15 0 1 9 13 2
11 13 0 9 1 9 13 2 0 7 0 2
5 3 3 15 13 2
11 2 3 13 2 15 3 3 13 9 0 2
16 3 3 0 3 13 0 9 2 9 3 13 2 16 9 13 2
9 3 0 3 13 9 7 13 0 2
37 3 16 0 13 9 7 13 9 2 9 13 2 1 3 9 0 13 2 3 3 3 15 13 9 2 15 3 13 2 7 15 3 13 13 0 9 2
11 3 15 3 13 3 3 13 2 1 9 2
35 2 16 15 9 13 2 13 0 9 2 13 2 9 0 7 9 2 3 3 3 3 9 0 3 13 9 9 1 9 2 3 9 13 9 2
15 3 13 0 9 9 0 2 1 9 0 13 1 9 0 2
21 15 3 9 9 0 13 13 1 9 0 2 3 3 9 0 2 3 9 3 13 2
16 15 3 9 13 0 9 9 13 2 0 0 0 7 0 13 2
8 15 3 0 1 9 9 13 2
13 3 15 3 13 1 9 0 13 7 13 13 9 2
25 3 16 9 13 9 0 9 2 3 15 3 0 13 9 9 3 13 2 3 3 16 3 0 13 2
7 9 3 15 0 13 13 2
10 3 3 0 13 9 0 2 3 13 2
5 15 3 0 13 2
11 0 3 13 15 3 15 15 9 9 13 2
24 3 3 1 9 13 9 0 13 3 2 15 3 9 13 0 9 13 2 9 3 0 9 13 2
19 3 3 3 13 0 1 9 0 2 15 3 13 0 9 1 9 13 13 2
7 15 3 9 13 13 2 2
7 15 3 3 9 13 9 2
10 3 0 9 13 0 9 2 9 9 2
17 3 15 3 0 1 0 13 2 13 1 9 9 2 1 9 9 2
26 3 15 9 13 2 1 3 9 13 3 2 1 15 13 7 13 7 13 9 0 2 15 15 9 13 2
18 1 3 9 0 9 13 2 15 3 9 3 13 1 9 2 1 9 2
8 3 9 9 7 9 9 13 2
18 2 15 3 3 13 0 9 1 2 9 3 3 9 13 15 15 0 2
24 3 15 9 13 0 2 16 3 15 13 7 13 9 2 7 3 13 2 0 9 3 13 2 2
7 3 13 9 0 9 13 2
15 15 3 3 3 3 13 2 3 9 1 13 0 9 13 2
12 10 3 0 9 13 0 1 9 2 13 9 2
25 13 3 13 9 0 0 2 1 3 9 0 9 0 13 2 9 13 2 9 3 1 9 9 1 2
10 3 3 0 9 9 13 2 9 13 2
13 3 3 15 13 13 0 13 2 0 0 9 13 2
8 15 13 3 13 3 0 9 2
9 3 3 15 3 13 9 9 13 2
7 15 3 13 13 0 9 2
21 3 3 9 3 9 1 3 15 13 2 3 3 15 15 0 13 13 9 7 9 2
12 0 3 13 2 16 13 13 3 2 13 3 2
6 15 3 9 13 9 2
5 15 3 9 13 2
12 1 3 15 13 2 15 3 13 7 15 13 2
23 9 3 13 0 1 0 9 3 13 2 7 3 3 15 9 0 9 0 0 0 13 9 2
15 13 3 1 9 9 13 2 3 13 9 9 9 13 0 2
53 9 3 15 13 0 12 9 2 13 3 15 9 0 0 2 12 3 0 9 2 0 3 9 2 0 3 9 0 2 0 3 1 15 9 2 3 3 3 9 2 0 9 13 2 9 0 2 15 13 0 13 2 2
9 15 3 13 3 9 1 9 13 2
9 9 3 0 0 13 2 0 13 2
13 3 3 15 9 13 13 9 3 2 15 15 13 2
6 15 3 9 13 13 2
10 3 15 0 13 0 2 16 3 13 2
5 15 3 13 9 2
14 3 3 9 13 0 2 15 15 13 3 0 3 9 2
7 15 3 13 13 0 9 2
9 2 3 15 15 0 3 3 13 2
15 13 3 1 8 2 3 0 9 13 2 9 9 9 9 2
7 3 15 3 9 13 9 2
11 3 15 9 13 1 9 3 13 3 13 2
10 9 3 15 15 13 1 9 1 9 2
19 3 9 15 3 0 9 13 2 1 15 3 13 7 0 13 9 2 0 2
22 3 3 15 0 13 9 13 2 0 2 15 13 3 15 13 0 2 13 3 0 13 2
13 9 3 3 15 13 13 9 7 0 9 13 2 2
10 3 13 2 15 3 9 9 13 0 2
14 0 3 9 13 9 0 13 1 9 0 2 0 13 2
17 15 3 13 9 2 1 9 3 15 3 0 9 13 0 9 13 2
9 13 3 15 13 13 2 7 13 2
7 3 13 9 9 3 0 2
5 1 3 15 13 2
6 3 3 13 13 3 2
14 9 13 1 0 9 2 9 13 0 7 0 9 2 2
7 15 3 13 13 0 9 2
18 2 9 3 0 15 13 9 2 15 1 9 15 13 9 0 9 13 2
26 15 3 15 13 7 0 9 1 9 9 9 0 2 16 7 13 9 2 15 3 13 15 13 7 13 2
28 6 3 3 15 3 9 0 1 9 13 2 15 15 3 13 2 15 3 13 15 0 0 13 2 1 9 13 2
12 1 3 0 13 2 15 3 13 7 13 0 2
11 9 15 13 12 7 12 9 2 9 12 2
13 9 3 15 3 13 13 12 2 0 3 0 13 2
15 3 3 1 9 0 13 2 16 3 9 9 13 3 2 2
20 3 13 2 15 3 0 13 9 7 0 9 2 9 13 15 15 3 13 9 2
7 1 3 9 0 13 9 2
10 15 3 1 15 13 13 0 0 9 2
15 3 16 3 13 7 1 9 9 13 2 3 9 13 13 2
21 3 3 3 13 1 9 16 3 0 3 13 0 2 9 3 3 13 9 9 2 2
7 15 3 13 13 0 9 2
11 2 13 2 3 3 0 1 9 0 13 2
10 3 13 1 9 2 15 9 1 13 2
16 3 3 9 7 9 7 9 13 2 16 3 9 13 0 2 2
8 3 3 13 13 1 9 0 2
18 3 9 3 13 9 13 9 9 2 0 3 16 3 7 0 13 13 2
5 1 3 9 13 2
13 13 3 15 0 9 2 16 13 0 9 0 3 2
7 7 15 13 9 0 13 2
8 15 3 3 9 13 9 13 2
16 3 3 15 9 13 0 1 9 2 15 3 9 3 13 2 2
18 15 3 16 3 13 9 13 3 9 2 3 13 1 9 3 9 3 2
15 15 3 16 3 9 13 13 3 9 2 13 1 9 13 2
7 3 9 0 9 13 13 2
14 0 3 9 13 13 13 1 9 2 15 13 3 2 2
27 3 3 13 2 9 3 3 13 9 13 0 2 9 3 13 13 9 1 9 2 7 15 13 9 0 13 2
12 3 13 2 15 3 3 3 13 0 1 9 2
9 3 15 3 1 9 1 9 13 2
17 9 3 3 9 3 1 9 13 3 2 9 0 9 7 9 13 2
10 0 3 1 9 13 0 2 13 9 2
9 15 15 3 9 13 13 7 13 2
19 15 3 1 9 13 0 3 7 0 13 3 9 0 2 1 3 13 9 2
7 3 3 3 0 13 3 2
19 9 3 15 3 13 3 13 13 2 16 3 3 9 3 9 3 9 13 2
16 3 3 15 3 1 9 0 13 13 2 7 0 13 13 13 2
9 3 13 2 16 13 13 0 2 2
11 3 13 9 13 2 9 3 13 0 0 2
6 9 3 13 9 0 2
8 15 3 3 13 9 13 13 2
10 3 3 9 0 3 9 15 13 9 2
16 0 15 13 9 0 2 15 3 9 1 13 7 9 0 13 2
18 0 3 9 3 3 1 9 13 13 2 3 3 9 13 13 1 9 2
6 15 3 0 13 2 2
12 3 13 2 15 3 3 0 1 0 9 13 2
8 15 3 0 13 3 7 3 2
7 15 15 0 13 7 13 2
6 15 3 3 13 13 2
5 3 3 3 13 2
5 13 15 3 13 2
11 3 13 2 16 3 15 0 0 13 2 2
12 3 13 2 15 3 3 13 0 9 0 0 2
6 15 3 0 3 13 2
12 3 3 15 13 9 1 9 2 7 9 13 2
7 3 3 3 1 9 13 2
15 3 16 3 13 1 9 0 9 2 0 13 1 9 0 2
6 15 3 9 13 9 2
6 3 9 9 9 13 2
16 7 3 9 3 0 7 9 0 13 2 7 9 1 0 13 2
7 15 3 13 13 9 9 2
4 13 7 13 2
6 13 3 15 3 13 2
26 16 3 9 13 0 9 2 9 0 13 15 3 13 3 2 15 3 3 9 3 9 3 9 9 13 2
16 15 3 0 13 7 10 3 2 9 3 7 9 3 13 2 2
14 3 13 13 3 13 9 2 13 3 1 9 9 13 2
19 15 3 16 3 9 0 1 9 13 2 15 3 3 9 13 0 0 9 2
11 2 13 15 13 16 3 3 13 13 2 2
3 3 13 2
9 1 3 9 9 13 2 3 13 2
13 13 3 3 1 9 13 2 15 3 3 13 0 2
7 3 3 9 9 0 13 2
6 2 15 3 3 13 2
5 3 13 0 2 2
21 3 16 3 13 1 9 0 9 2 13 3 9 2 1 3 13 2 13 3 9 2
8 15 3 13 13 0 0 9 2
8 15 3 3 9 13 3 13 2
10 3 13 2 9 3 13 7 9 13 2
4 3 3 13 2
10 9 3 9 3 9 1 9 13 2 2
7 15 3 13 13 0 9 2
21 15 3 3 9 13 2 1 3 13 9 2 13 3 13 2 13 3 9 1 0 2
17 1 3 13 0 9 7 0 9 2 13 3 9 3 7 9 0 2
10 3 13 9 2 15 3 0 9 13 2
19 15 3 3 13 1 9 13 9 2 0 3 1 9 13 2 9 9 13 2
7 1 3 9 13 13 9 2
15 0 3 13 0 0 9 2 13 3 13 3 3 9 0 2
15 7 3 3 9 13 0 9 2 1 3 13 1 0 0 2
7 3 3 9 13 0 9 2
12 3 13 9 2 15 3 13 2 13 3 9 2
22 9 3 13 2 13 0 9 2 9 1 0 2 16 0 13 7 0 9 1 0 9 2
16 12 3 9 13 2 0 3 1 0 13 7 13 3 12 9 2
11 1 3 3 9 9 13 2 13 3 9 2
19 3 3 3 9 13 2 16 13 9 2 3 13 9 7 15 15 9 13 2
8 3 3 3 3 13 9 0 2
8 13 15 15 9 1 9 13 2
9 13 3 15 0 2 16 0 13 2
5 9 3 3 13 2
6 3 3 13 13 2 2
6 3 3 3 13 15 2
8 3 3 3 3 9 13 0 2
13 3 3 13 3 15 9 3 13 3 13 3 2 2
8 7 3 13 13 9 9 3 2
29 13 3 1 0 9 9 3 7 9 2 3 3 9 13 1 9 2 1 3 9 9 13 9 3 13 0 3 13 2
26 0 9 9 3 13 0 13 9 7 13 1 9 9 1 0 1 9 0 1 3 9 9 7 9 0 2
13 13 3 3 9 9 2 1 3 9 13 0 9 2
27 3 16 13 3 7 13 2 15 9 13 2 13 3 0 3 9 0 9 13 2 16 3 0 13 0 13 2
6 0 3 9 13 9 2
9 3 0 13 2 9 3 15 0 2
8 3 15 0 13 0 9 2 2
9 3 13 1 9 13 9 0 9 2
14 13 3 9 13 9 0 2 16 15 0 13 0 9 2
7 3 3 13 0 9 9 2
19 9 3 0 7 9 9 13 2 3 3 0 13 0 9 0 9 0 9 2
18 13 3 3 9 7 15 13 13 2 16 3 13 0 1 9 0 2 2
9 3 3 3 13 7 0 0 13 2
7 13 3 9 0 9 0 2
8 3 3 3 13 9 0 9 2
15 15 3 16 13 9 0 7 13 2 9 13 13 0 9 2
18 2 3 3 0 13 13 7 13 9 2 10 15 13 2 16 13 9 2
5 3 13 0 9 2
22 7 15 1 9 7 3 13 0 3 9 1 9 2 15 3 13 9 13 0 0 13 2
23 0 3 1 9 9 9 13 2 16 15 1 9 13 13 7 16 15 9 0 1 9 13 2
6 15 3 3 15 13 2
6 15 1 9 0 13 2
26 3 3 10 0 9 13 2 16 3 13 0 0 9 13 2 16 3 13 9 0 7 0 9 13 13 2
7 1 3 15 0 13 9 2
8 0 3 0 1 15 13 0 2
9 15 3 0 0 3 13 0 9 2
8 3 3 13 0 0 9 13 2
14 0 3 15 0 13 13 0 9 2 3 3 13 9 2
5 9 15 13 13 2
17 3 3 3 9 3 13 2 3 3 3 13 9 0 3 13 13 2
38 3 16 9 9 13 0 2 13 3 1 9 2 9 3 13 0 2 3 3 3 9 0 1 9 13 9 0 2 16 3 3 0 3 3 0 0 13 2
12 3 15 0 0 9 13 9 1 0 9 9 2
8 15 3 9 9 1 0 13 2
20 3 3 3 9 13 0 0 9 13 1 0 9 9 2 3 3 9 3 13 2
10 3 3 3 3 9 13 9 3 13 2
8 7 15 3 0 13 9 13 2
8 9 3 13 0 9 13 0 2
7 1 3 9 13 9 0 2
5 0 3 13 13 2
12 15 3 3 3 13 2 13 3 9 0 9 2
11 1 9 3 13 13 0 9 2 3 13 2
18 9 3 3 3 13 9 2 0 2 15 3 9 13 0 1 0 3 2
10 13 3 9 9 0 2 13 3 9 2
40 3 3 3 1 15 13 0 9 2 1 9 3 13 0 9 13 2 7 1 9 13 0 2 9 1 9 2 0 1 0 13 2 7 1 9 2 1 0 9 2
6 13 3 9 13 9 2
7 13 3 1 0 9 13 2
14 15 3 3 3 0 9 13 2 1 3 9 0 13 2
12 9 3 9 0 1 9 13 2 9 0 13 2
15 0 9 13 2 16 1 9 9 0 9 9 9 0 13 2
19 0 3 9 9 13 9 2 15 13 1 9 2 9 3 15 3 15 13 2
8 3 3 3 0 3 3 13 2
8 15 3 3 9 13 0 13 2
14 3 3 15 0 13 9 9 2 9 3 0 7 15 2
7 3 3 13 13 3 2 2
19 13 15 2 7 0 13 2 7 15 3 9 13 1 9 2 13 9 9 2
21 15 3 13 16 3 3 15 9 13 13 2 7 15 3 0 13 7 3 0 0 2
8 15 3 3 9 13 0 13 2
5 3 3 0 13 2
4 9 15 13 2
16 3 3 15 3 13 15 13 2 3 3 16 9 3 13 2 2
9 3 9 3 13 3 3 9 13 2
32 13 3 3 15 3 3 9 0 13 3 3 13 7 0 9 13 2 7 13 13 0 2 3 9 13 1 9 9 7 15 9 2
8 15 3 3 9 13 0 13 2
16 0 3 3 9 0 2 7 15 3 13 0 9 7 9 0 2
18 3 3 13 9 0 13 7 13 9 2 16 1 13 9 7 9 0 2
9 3 3 3 15 13 13 9 9 2
7 3 13 9 0 9 9 2
4 3 9 13 2
13 15 3 0 13 9 9 0 2 16 13 0 0 2
34 3 3 15 3 3 13 0 1 9 13 2 7 3 15 3 9 3 7 9 13 13 1 9 1 9 2 3 3 3 15 15 13 9 2
6 3 3 0 13 9 2
9 15 3 3 3 0 13 9 13 2
12 15 3 0 9 9 0 0 0 9 13 9 2
5 9 3 13 0 2
17 1 3 3 13 3 9 9 2 15 0 13 9 3 13 13 9 2
33 3 16 3 15 9 9 13 13 2 3 3 10 3 9 13 1 9 0 13 9 9 7 9 13 2 15 3 13 13 13 0 3 2
18 3 15 3 3 13 2 13 3 9 2 16 9 13 7 1 9 13 2
41 3 16 3 3 0 13 1 9 9 1 9 0 9 9 0 13 13 2 3 3 0 9 0 9 13 2 0 3 9 1 9 13 2 9 3 13 0 2 0 9 2
14 3 13 15 3 9 13 2 3 9 13 9 1 9 2
15 13 3 15 0 0 3 1 9 9 9 9 1 0 9 2
19 3 9 0 9 1 0 9 13 2 1 9 2 0 3 9 0 9 13 2
20 15 3 3 3 13 2 9 3 13 9 9 2 3 9 3 1 9 13 9 2
13 3 10 12 9 0 9 13 13 9 3 7 9 2
16 3 15 3 3 0 9 7 9 13 13 1 9 1 0 9 2
8 3 3 0 9 13 3 0 2
15 0 3 13 0 9 2 13 9 2 13 3 9 1 0 2
15 3 3 15 15 13 13 9 0 9 3 0 7 0 9 2
17 3 3 15 13 9 0 9 0 9 13 2 0 15 9 9 13 2
10 3 1 3 9 15 13 7 13 13 2
42 0 3 0 3 13 2 1 10 9 2 3 3 13 3 9 13 2 15 15 0 13 9 1 9 0 0 2 3 3 3 3 3 9 0 13 2 16 0 3 0 3 2
11 3 13 3 1 9 3 0 7 0 9 2
9 13 3 15 0 2 16 0 13 2
5 9 3 3 13 2
12 3 13 2 9 3 3 13 7 1 9 13 2
19 3 3 13 3 9 2 13 3 9 2 16 9 7 0 0 13 9 13 2
10 3 9 1 9 13 2 7 13 2 2
10 13 3 9 9 2 15 3 13 13 2
22 15 3 9 3 9 1 9 13 2 9 3 9 13 0 2 13 3 3 0 13 9 2
10 9 3 1 9 13 2 13 3 13 2
24 3 16 13 3 13 3 2 0 13 9 2 3 3 9 7 9 0 0 13 0 1 9 13 2
7 9 3 3 13 13 9 2
11 15 3 13 9 13 2 16 0 0 3 2
15 3 0 3 3 0 3 13 2 16 3 13 0 1 9 2
15 15 3 1 9 0 13 2 16 13 3 9 13 3 0 2
8 0 3 1 15 0 13 13 2
13 10 3 0 9 0 9 13 2 0 9 0 9 2
9 3 3 13 0 1 9 0 3 2
19 3 3 1 9 0 13 3 9 15 13 2 3 3 0 3 3 3 0 2
16 15 3 0 2 16 0 13 9 2 13 1 9 3 7 9 2
14 13 3 15 9 2 15 15 0 13 7 9 0 2 2
9 3 3 13 13 0 9 9 13 2
6 9 3 13 0 13 2
9 13 3 10 0 2 16 13 9 2
12 9 3 13 9 2 9 3 13 1 3 13 2
18 15 3 3 15 13 9 9 0 0 2 15 3 3 1 9 13 9 2
9 15 15 15 13 9 9 13 2 2
10 3 13 13 2 15 3 13 9 9 2
16 3 16 9 13 0 10 9 2 3 13 1 9 3 9 3 2
21 15 3 10 9 13 1 9 13 9 0 2 15 0 9 13 9 7 1 9 13 2
17 0 3 3 13 9 9 0 2 15 3 9 9 9 13 7 9 2
16 15 3 3 0 9 13 9 2 1 3 3 9 0 13 13 2
20 3 3 15 3 3 1 9 2 13 2 16 0 13 2 13 3 9 9 9 2
17 9 3 1 9 0 9 0 0 13 9 13 2 13 3 12 0 2
15 9 3 3 9 9 3 13 13 2 16 9 9 9 13 2
28 10 3 0 13 3 0 2 13 3 3 9 1 9 0 9 13 2 9 3 9 3 3 7 0 13 9 2 2
9 3 13 2 15 3 3 0 13 2
6 13 3 9 0 13 2
7 9 3 9 9 9 13 2
14 15 3 3 9 9 13 13 2 16 9 9 13 13 2
9 9 3 13 9 9 7 0 9 2
30 9 3 15 9 1 0 9 13 1 9 13 2 0 3 13 9 1 9 9 3 0 9 0 13 1 9 13 9 13 2
5 9 3 9 13 2
22 9 3 9 9 9 3 9 3 13 2 0 3 9 13 13 2 9 9 1 9 13 2
11 9 3 13 9 0 2 13 3 9 9 2
9 15 3 3 13 1 9 9 13 2
39 15 3 16 1 0 9 13 2 13 3 9 9 2 3 3 15 13 2 3 3 1 9 13 0 1 9 2 1 3 9 13 0 13 2 1 0 3 13 2
13 13 3 1 9 10 9 2 1 3 9 9 13 2
8 0 3 1 0 13 9 9 2
26 3 16 1 9 13 7 9 13 2 13 3 3 0 7 1 9 13 2 13 3 0 9 1 9 13 2
26 3 16 13 3 7 13 3 9 2 1 3 15 9 0 13 7 9 2 1 3 9 13 9 0 0 2
12 15 3 16 13 9 0 7 13 2 13 13 2
11 1 3 9 0 13 9 13 1 0 9 2
16 1 3 9 9 9 7 9 13 9 3 2 0 13 0 9 2
8 1 3 3 9 0 13 9 2
8 15 3 0 13 9 3 13 2
12 3 3 9 13 2 15 3 15 1 0 13 2
16 16 3 9 13 0 9 2 9 3 13 1 3 9 0 13 2
8 1 3 13 9 7 9 0 2
10 13 3 13 2 15 3 3 0 13 2
12 13 3 1 9 0 2 3 3 3 13 9 2
6 0 3 13 0 9 2
8 13 3 9 13 3 0 9 2
15 15 3 13 0 9 0 2 1 3 3 9 13 9 0 2
15 15 3 13 13 9 0 9 9 7 9 0 0 1 9 2
7 15 3 9 9 9 13 2
18 15 3 15 3 3 9 7 9 13 13 9 1 9 0 2 15 13 2
21 1 3 15 13 0 9 13 2 0 3 9 1 0 2 9 9 2 13 1 0 2
19 3 13 2 7 15 13 0 9 2 7 0 13 13 2 15 3 13 2 2
8 15 3 0 13 13 0 9 2
9 3 3 3 3 9 3 0 13 2
21 3 3 3 15 9 0 13 0 9 3 13 2 16 3 3 9 3 3 13 9 2
13 3 13 9 9 2 1 3 0 3 13 13 2 2
18 3 13 2 15 3 9 13 2 13 3 0 0 9 3 13 15 0 2
41 15 3 9 3 13 1 9 13 2 7 15 3 13 1 0 9 2 1 3 13 9 2 1 3 9 0 13 2 9 3 13 1 9 13 2 15 3 13 0 9 2
9 15 3 13 13 1 9 0 9 2
14 3 3 3 9 9 13 7 9 9 1 0 9 0 2
13 3 16 13 13 9 2 1 3 9 13 0 13 2
27 15 3 16 3 9 13 7 13 9 2 1 3 3 9 0 13 7 9 2 1 3 9 13 1 9 9 2
14 9 3 0 9 13 13 0 0 1 0 9 2 13 2
6 1 3 0 13 9 2
14 9 3 0 9 13 13 2 9 0 13 2 13 13 2
15 9 3 9 9 13 13 0 2 1 3 15 13 0 9 2
7 15 3 13 13 0 9 2
7 2 9 3 13 7 13 2
11 3 3 9 13 13 2 15 15 13 9 2
22 3 13 2 7 15 9 9 1 0 13 0 1 9 13 2 15 3 15 9 13 0 2
9 15 3 1 9 0 13 9 13 2
26 3 16 9 7 9 1 9 13 2 3 3 9 13 9 9 2 3 13 9 2 16 3 13 10 0 2
6 9 15 13 13 2 2
14 15 3 13 13 0 9 2 7 15 13 9 0 13 2
9 0 3 15 3 9 7 9 13 2
39 3 3 0 13 7 0 13 13 1 9 7 0 9 13 2 9 9 3 7 0 13 2 9 3 13 7 0 7 9 7 9 2 3 3 9 3 0 13 2
8 3 3 13 9 0 1 9 2
22 16 15 1 0 0 9 13 13 2 3 15 9 0 13 3 2 3 2 9 0 9 2
8 3 3 3 13 15 9 13 2
28 3 9 15 13 13 2 15 15 15 13 2 16 3 0 13 2 7 13 9 3 3 13 2 13 0 7 0 2
26 15 13 0 3 13 1 9 9 13 2 10 3 9 0 13 2 15 3 13 9 1 0 1 9 0 2
31 15 3 3 13 0 9 13 2 15 3 9 3 0 0 2 16 3 0 13 2 3 3 15 13 2 13 15 3 7 13 2
12 3 13 2 15 3 3 9 1 9 13 9 2
17 9 3 1 9 3 13 9 13 2 9 0 1 9 13 0 9 2
27 13 3 15 9 2 13 3 3 1 9 7 1 9 2 7 15 0 9 13 13 7 0 13 0 3 13 2
21 16 15 0 13 1 9 7 1 9 2 1 3 9 9 0 0 13 9 0 13 2
16 15 9 13 12 0 9 2 0 3 9 2 12 3 9 9 2
9 3 3 3 9 9 13 0 9 2
15 0 3 9 9 3 0 13 0 2 9 3 1 9 13 2
11 15 3 15 0 9 13 13 9 0 13 2
9 3 1 0 9 13 0 9 13 2
11 13 3 1 9 2 1 3 9 9 13 2
9 3 3 15 3 9 9 13 0 2
5 13 7 0 13 2
5 13 3 15 9 2
7 15 3 13 13 0 9 2
8 15 3 3 9 9 0 13 2
15 13 3 15 13 2 16 15 7 15 9 13 7 15 9 2
36 0 3 9 13 9 9 13 1 9 2 15 3 0 9 13 2 3 3 9 15 3 13 2 3 3 15 0 13 15 3 1 9 13 9 2 2
7 15 3 13 13 0 9 2
22 7 15 13 13 13 0 0 0 2 16 15 1 9 9 13 9 0 13 0 0 9 2
7 7 3 3 3 13 13 2
20 3 3 3 15 0 13 13 3 13 3 2 16 3 16 3 9 0 9 13 2
11 3 13 2 15 3 0 1 9 13 9 2
25 13 3 0 9 2 9 13 2 13 3 9 3 7 9 9 2 3 3 3 9 9 0 13 9 2
15 13 3 1 9 0 9 2 15 3 9 13 0 0 9 2
8 15 15 3 13 9 0 13 2
11 3 3 2 16 3 3 13 2 13 15 2
14 3 3 15 3 13 13 0 2 7 3 9 13 9 2
13 13 3 3 0 13 15 3 13 9 7 9 13 2
11 3 3 0 13 9 2 3 3 0 0 2
5 13 3 15 13 2
7 15 3 13 13 0 9 2
21 15 3 9 3 13 2 15 3 13 2 9 3 3 13 2 9 3 1 9 13 2
13 9 3 3 3 3 13 9 7 15 13 0 2 2
9 15 3 1 9 0 13 9 13 2
8 3 3 0 13 9 9 13 2
19 3 3 1 9 13 9 2 3 13 2 0 3 0 3 2 0 0 0 2
44 15 15 13 2 16 9 13 2 3 3 0 3 13 1 9 9 2 3 3 16 15 13 9 3 9 3 2 3 3 16 15 1 9 7 0 9 9 13 2 15 3 9 13 2
6 3 3 9 13 9 2
13 3 16 3 13 13 3 13 2 3 9 13 13 2
4 13 3 0 2
11 3 3 3 13 13 1 9 7 9 13 2
4 13 3 13 2
16 0 3 3 3 15 13 3 3 13 2 0 9 9 13 9 2
17 3 0 15 13 7 13 0 9 9 1 9 2 3 13 9 0 2
21 0 15 9 0 13 2 9 0 1 9 13 2 9 13 2 9 0 13 9 0 2
11 15 0 13 9 9 2 15 3 13 0 2
12 15 3 15 0 13 0 13 2 7 15 13 2
5 15 3 9 13 2
16 0 3 9 13 0 9 13 1 0 2 1 3 9 13 0 2
6 3 0 0 3 13 2
53 3 0 9 13 2 16 3 15 9 13 13 3 3 2 9 3 13 2 15 9 13 2 16 15 13 3 0 1 9 9 2 9 3 0 13 9 3 9 3 3 15 13 2 3 3 3 9 3 3 15 9 2 2
7 15 3 13 13 0 9 2
16 3 3 0 13 9 3 9 3 9 9 2 0 3 13 9 2
15 3 3 3 0 15 13 9 2 0 9 0 13 0 9 2
23 0 3 15 13 7 13 0 9 9 1 0 2 7 13 0 0 0 9 9 7 9 13 2
5 13 3 15 3 2
12 13 3 15 13 9 2 15 9 13 9 13 2
7 7 15 8 0 13 13 2
20 3 3 13 0 9 13 2 1 3 3 9 13 0 2 0 0 9 13 9 2
14 3 15 7 8 7 0 9 13 1 0 13 7 13 2
13 15 3 0 13 13 7 13 2 7 3 3 13 2
8 3 9 13 7 13 13 3 2
18 3 0 3 0 3 13 9 0 2 9 3 15 3 0 13 9 13 2
14 3 9 1 9 9 13 3 0 2 13 3 0 0 2
12 3 3 13 2 16 15 3 13 9 9 2 2
8 15 3 3 9 13 0 13 2
19 3 3 15 15 15 13 0 9 2 3 3 16 15 9 3 0 3 13 2
17 3 3 1 9 13 15 2 16 3 3 9 1 0 13 13 2 2
29 3 13 2 0 3 9 9 13 9 1 9 13 7 9 0 0 13 13 3 3 9 2 9 3 13 0 3 13 2
14 15 3 13 1 9 9 1 9 13 2 9 3 13 2
6 1 3 9 13 9 2
52 16 3 9 13 0 9 2 13 3 1 9 9 0 9 9 13 2 1 3 9 0 13 9 2 9 3 1 0 13 0 9 2 13 3 13 1 9 9 0 3 2 9 3 13 2 9 3 13 1 3 13 2
6 15 15 0 13 2 2
8 15 3 3 9 13 0 13 2
26 3 3 10 0 9 13 2 16 3 13 0 0 9 13 2 16 3 13 9 0 7 0 9 13 13 2
7 1 3 15 0 13 9 2
18 3 3 15 15 13 13 3 3 13 2 7 3 15 13 3 13 9 2
8 15 3 0 13 13 0 9 2
8 0 3 0 3 13 0 3 2
17 2 9 15 3 3 9 13 13 13 2 16 3 15 13 0 9 2
8 10 3 3 13 9 13 9 2
30 9 3 15 13 0 1 9 9 1 2 9 3 15 13 2 0 3 0 3 0 0 9 13 2 15 0 9 13 3 2
26 3 15 12 9 13 9 2 3 3 3 9 13 13 0 2 15 3 3 9 9 13 1 0 9 9 2
8 15 3 3 3 3 9 13 2
8 15 15 0 13 13 1 9 2
31 2 1 3 15 13 2 15 15 15 3 13 9 2 16 15 3 15 0 13 2 7 3 13 0 13 2 15 9 0 13 2
10 15 3 3 0 13 9 13 7 13 2
17 2 0 3 13 15 9 0 9 2 16 3 15 13 7 13 13 2
9 0 3 3 13 9 9 9 13 2
11 2 3 13 2 15 3 3 13 0 9 2
30 16 3 9 0 9 13 2 3 3 1 9 13 9 0 0 9 1 9 0 9 13 2 1 3 13 13 1 9 0 2
10 3 15 15 13 1 9 13 13 3 2
8 0 3 15 13 0 10 9 2
8 9 3 3 0 13 7 13 2
15 3 16 0 13 7 13 2 13 1 0 9 3 9 9 2
27 15 3 16 3 0 13 13 2 3 3 3 15 13 9 3 9 3 2 3 3 13 13 7 0 3 13 2
17 0 3 13 13 2 0 1 9 9 13 2 7 9 7 0 9 2
7 0 3 15 9 13 13 2
7 3 3 13 1 9 9 2
19 16 3 9 13 0 9 2 3 3 3 1 9 9 0 13 0 9 13 2
5 0 3 13 0 2
5 9 3 13 9 2
9 9 3 1 9 13 0 13 13 2
7 15 3 3 1 13 0 2
10 3 3 13 2 13 3 1 9 0 2
6 3 3 0 9 13 2
8 13 3 3 9 0 0 9 2
8 15 3 3 0 1 9 13 2
8 3 0 13 7 13 0 9 2
15 9 1 9 0 13 13 0 3 13 2 13 3 9 9 2
7 0 3 0 13 13 9 2
7 9 3 1 9 13 0 2
9 15 3 3 3 13 1 9 9 2
22 0 3 10 9 13 1 9 2 13 3 9 0 2 0 3 3 13 2 13 3 9 2
15 1 3 15 0 13 9 2 3 3 15 9 13 9 13 2
10 15 3 13 13 2 1 3 9 13 2
25 3 3 10 9 0 13 9 2 7 3 3 0 9 13 0 2 3 3 9 7 9 7 0 9 2
8 13 3 0 9 7 9 0 2
7 15 3 3 13 13 9 2
18 3 16 3 3 13 10 9 0 13 2 3 3 3 15 9 13 13 2
10 2 3 13 2 3 15 15 13 13 2
25 2 3 3 13 9 3 0 3 9 13 0 0 13 2 16 0 0 1 9 13 13 1 9 9 2
11 7 3 15 13 9 9 2 15 15 13 2
7 3 3 3 9 13 13 2
11 2 3 13 2 15 3 15 3 13 13 2
13 3 3 15 15 13 13 2 3 3 13 0 9 2
13 3 3 15 13 3 0 13 2 16 3 0 13 2
11 9 3 3 12 0 0 9 1 9 13 2
7 9 3 3 3 15 13 2
9 9 3 3 3 0 13 0 9 2
8 2 9 3 1 9 13 0 2
11 9 15 0 9 13 9 0 7 13 9 2
19 3 3 3 13 9 3 13 3 9 2 16 3 0 9 13 7 0 13 2
9 13 3 3 9 13 0 9 9 2
7 15 3 9 0 13 13 2
15 3 3 9 13 9 0 13 0 9 2 1 3 13 0 2
21 3 10 3 3 13 2 10 3 9 13 9 2 15 3 9 10 0 13 0 13 2
8 15 3 13 1 9 0 13 2
11 3 15 3 3 13 2 16 13 0 9 2
5 13 3 9 9 2
39 3 16 3 3 13 9 9 0 13 2 3 3 15 13 9 9 1 0 13 0 13 2 9 1 9 2 3 9 13 9 10 3 2 3 3 13 9 9 2
33 3 16 3 3 3 13 9 0 2 3 3 9 9 13 2 7 3 13 2 3 3 15 3 13 13 0 9 7 13 13 0 9 2
13 0 3 1 0 9 0 13 2 16 3 13 9 2
23 15 3 3 1 9 13 9 2 15 3 13 9 9 13 2 1 3 13 9 9 0 9 2
17 13 3 15 3 1 9 2 16 15 13 13 2 13 3 9 9 2
9 13 3 13 13 1 9 9 9 2
7 3 3 9 0 13 9 2
15 13 1 9 12 9 0 13 9 2 3 3 13 9 13 2
21 3 3 15 9 9 13 15 15 13 2 3 3 15 9 2 3 13 1 9 2 2
30 2 3 13 2 3 15 3 13 0 9 2 13 3 1 9 13 2 3 3 3 15 9 13 3 13 7 13 9 9 2
16 3 16 13 3 13 3 13 2 3 3 15 13 9 0 0 2
11 3 0 13 16 3 3 0 0 9 13 2
6 8 0 3 3 13 2
16 15 3 0 9 13 2 15 15 3 0 13 0 9 7 13 2
8 13 3 3 13 3 13 2 2
11 2 3 13 2 15 3 15 3 13 13 2
20 15 3 13 1 9 0 1 9 13 2 9 1 9 9 2 15 15 9 13 2
9 15 3 3 13 0 0 9 13 2
24 3 9 2 3 3 3 9 0 3 3 3 9 2 7 3 9 0 13 9 9 13 13 9 2
8 2 3 13 1 9 13 13 2
16 3 15 1 9 1 0 9 13 2 0 3 15 9 13 13 2
26 3 16 3 1 9 13 7 9 2 9 3 13 2 1 3 13 0 9 2 3 3 13 1 9 9 2
33 16 3 9 13 0 9 2 9 3 0 13 1 9 0 2 1 3 9 13 7 9 9 0 2 1 3 3 0 13 1 9 13 2
8 3 3 13 0 9 13 9 2
14 3 3 1 9 0 9 13 9 2 7 13 0 9 2
17 3 16 13 9 9 3 13 2 13 9 9 2 16 0 9 13 2
18 0 13 13 2 13 3 15 9 0 2 15 15 3 0 1 9 13 2
16 3 3 3 13 1 9 0 2 16 3 0 3 0 3 13 2
16 3 3 13 0 9 2 16 13 9 0 15 13 9 0 2 2
8 15 3 3 9 13 0 13 2
9 3 3 9 9 3 0 13 13 2
9 3 3 15 13 9 1 9 0 2
7 15 3 15 9 3 13 2
10 9 3 15 3 15 13 2 9 13 2
14 9 3 1 9 3 13 2 7 15 0 3 13 9 2
24 15 3 9 13 0 2 15 1 3 9 0 2 1 3 9 9 3 9 3 7 0 9 0 2
20 3 13 2 13 3 9 0 9 2 9 3 15 13 9 3 13 1 3 13 2
6 3 15 15 0 13 2
3 13 3 2
16 9 3 0 1 0 9 9 13 2 13 15 0 7 0 13 2
5 13 15 9 13 2
14 0 3 13 0 2 9 3 9 13 2 9 3 9 2
7 15 3 13 15 13 2 2
16 3 15 3 0 1 0 13 2 9 3 1 9 13 0 9 2
11 15 3 13 3 9 2 13 3 9 9 2
7 9 3 15 9 9 13 2
9 3 15 3 1 9 1 9 13 2
21 9 3 1 9 9 9 13 7 9 13 1 0 9 2 3 3 3 2 9 13 2
5 9 15 13 13 2
7 15 3 15 13 13 2 2
9 3 13 2 15 3 1 9 13 2
18 3 3 13 1 9 13 0 2 7 3 0 9 7 9 13 7 9 2
13 2 0 15 13 2 15 13 7 15 0 9 13 2
6 13 3 3 15 13 2
28 3 15 0 13 0 2 16 3 13 2 7 15 9 0 13 9 0 2 7 0 15 13 2 16 13 9 2 2
6 2 0 0 15 13 2
14 15 3 13 3 0 2 16 9 0 13 9 9 13 2
6 0 3 13 9 13 2
17 1 3 9 15 13 13 9 2 7 9 2 15 3 0 0 13 2
4 3 15 13 2
14 13 3 9 0 0 0 2 3 3 13 9 3 2 2
15 3 3 13 13 1 9 9 2 15 3 0 13 9 0 2
8 9 3 3 13 7 13 9 2
14 9 3 0 9 0 13 2 9 3 15 9 13 13 2
6 13 3 15 3 13 2
16 1 15 3 0 9 13 3 9 13 2 13 3 1 9 0 2
6 13 3 3 0 13 2
12 3 15 0 9 13 9 2 16 9 9 13 2
33 3 3 15 13 9 0 7 12 9 2 16 15 0 13 13 7 13 1 9 9 3 9 3 0 2 16 3 3 13 1 9 2 2
12 2 3 13 2 15 3 3 0 13 7 13 2
8 3 3 13 13 9 1 9 2
16 3 3 3 9 0 9 13 0 9 2 15 9 1 9 13 2
13 9 3 15 13 9 2 15 13 9 9 1 13 2
6 15 3 3 9 13 2
8 13 3 13 13 1 9 9 2
8 15 3 1 9 13 13 9 2
13 3 13 3 3 3 13 0 7 0 3 3 13 2
38 3 3 15 9 0 10 3 13 2 9 13 2 0 9 13 1 0 9 2 3 3 15 13 0 3 3 15 13 1 9 2 15 3 13 9 0 9 2
9 0 3 13 9 2 0 3 13 2
9 0 3 3 3 3 0 9 13 2
19 3 10 3 0 9 7 0 9 13 2 3 3 15 13 9 3 0 2 2
8 15 3 3 13 9 13 13 2
15 3 0 0 3 7 0 0 9 13 2 15 3 13 9 2
8 9 13 13 0 9 3 13 2
15 15 3 13 1 9 9 1 9 0 7 1 9 0 2 2
19 3 13 2 15 3 3 13 9 7 0 9 2 3 3 15 9 9 13 2
13 10 3 15 9 9 13 2 0 3 15 13 9 2
8 3 3 3 15 9 13 13 2
8 15 3 13 3 9 13 13 2
31 2 3 13 7 15 15 9 13 2 7 3 0 9 13 13 1 9 2 16 13 9 0 7 9 7 15 15 9 13 2 2
8 3 3 13 13 1 9 9 2
28 15 3 9 13 0 2 3 3 3 3 13 9 13 0 1 9 13 2 7 3 1 9 13 0 9 0 13 2
14 1 3 9 13 0 2 0 1 9 13 0 7 0 2
7 15 3 0 13 13 9 2
16 1 3 15 0 9 13 1 0 2 0 15 3 13 7 13 2
15 3 3 9 0 13 9 9 1 9 2 3 3 13 13 2
8 15 3 3 13 0 9 9 2
6 9 3 15 3 13 2
31 15 3 13 0 9 7 3 15 13 2 16 0 3 13 7 15 0 13 7 13 13 2 16 3 3 13 1 9 0 13 2
10 15 3 3 15 3 3 1 9 13 2
6 3 3 9 13 13 2
13 3 13 2 15 3 13 9 2 13 3 9 9 2
25 15 3 13 2 0 9 9 13 1 9 13 1 0 9 2 1 3 13 9 9 2 13 3 9 2
10 3 13 13 2 9 3 15 13 9 2
7 9 3 13 1 9 0 2
7 3 3 15 13 0 9 2
21 2 3 3 3 9 15 9 9 13 2 3 3 15 13 15 15 9 9 13 2 2
18 3 3 9 0 13 13 9 2 15 3 3 0 1 9 13 15 2 2
17 3 13 13 12 9 0 2 13 3 13 1 9 0 7 9 9 2
7 9 3 15 13 0 9 2
13 3 3 1 0 15 3 13 2 1 3 13 0 2
11 3 3 9 13 2 13 3 1 0 13 2
23 0 3 13 9 9 1 9 13 2 7 15 0 1 9 13 2 0 15 13 13 0 9 2
10 13 3 13 2 13 3 15 9 0 2
18 13 3 15 1 9 9 0 2 16 9 13 13 13 9 9 3 0 2
20 1 9 3 13 1 9 9 2 13 3 3 1 9 2 7 15 1 9 13 2
22 3 3 15 3 3 13 9 3 13 13 3 3 13 2 16 3 3 0 13 0 9 2
9 3 3 3 15 9 13 13 2 2
14 15 3 13 3 9 9 2 0 3 13 1 0 9 2
13 3 15 3 3 13 2 16 3 0 3 9 13 2
43 7 15 13 13 9 7 9 0 2 15 15 13 1 9 7 1 9 2 15 3 3 9 0 13 9 2 0 9 13 1 9 2 0 2 15 9 0 1 9 7 0 9 2
10 15 3 15 3 3 13 7 3 0 2
15 0 3 0 1 0 13 2 13 13 16 0 9 13 2 2
7 15 3 13 13 9 0 2
12 2 13 2 3 3 15 3 1 9 13 3 2
5 15 3 13 13 2
7 15 3 3 13 9 9 2
7 15 3 13 13 9 0 2
10 3 13 9 1 9 13 1 9 9 2
14 0 3 15 9 13 2 16 15 0 9 13 9 9 2
13 9 3 13 13 0 9 9 9 0 1 9 13 2
7 3 15 3 13 13 0 2
16 9 3 1 9 1 0 9 13 2 16 0 9 13 7 9 2
9 15 3 9 13 9 0 9 13 2
8 13 3 15 13 1 9 9 2
16 7 3 15 13 9 0 9 15 13 2 9 3 3 0 13 2
19 3 15 3 1 9 13 0 9 13 9 1 9 9 2 15 15 9 13 2
9 15 3 3 13 0 0 9 13 2
9 3 3 9 0 13 13 3 13 2
15 15 3 13 1 9 9 1 9 0 7 1 9 0 2 2
7 15 3 13 13 9 9 2
17 3 3 3 0 3 13 9 0 2 16 3 3 0 9 13 13 2
20 3 3 15 9 13 0 3 13 7 13 9 1 0 7 0 1 0 9 2 2
9 3 13 2 3 3 13 9 9 2
25 3 3 1 9 13 0 9 2 0 0 2 15 15 13 7 1 0 7 1 0 9 1 9 9 2
8 15 1 9 13 13 0 9 2
8 9 3 13 1 9 13 9 2
22 13 3 1 9 9 9 13 2 15 3 1 0 9 9 0 9 13 0 9 13 9 2
7 15 0 0 13 9 9 2
28 3 16 3 10 9 13 3 13 2 3 1 9 13 0 3 13 2 16 0 9 13 2 15 1 9 13 0 2
6 15 3 3 13 13 2
20 9 3 1 9 0 13 2 3 3 9 9 3 0 9 3 1 9 13 13 2
12 15 3 3 13 9 0 9 13 0 9 13 2
14 9 3 3 9 13 9 0 2 0 0 13 3 0 2
9 3 3 9 0 9 7 9 13 2
14 3 3 3 3 0 3 13 13 13 7 13 9 15 2
6 3 13 13 9 9 2
15 3 16 3 0 0 13 9 2 3 3 1 0 9 13 2
17 3 3 3 9 9 0 13 0 2 3 3 16 15 3 9 13 2
28 3 3 3 9 9 3 13 2 3 15 3 1 9 13 13 2 3 3 3 2 9 7 9 7 9 9 13 2
7 9 1 0 13 9 13 2
7 3 3 3 3 15 13 2
5 13 15 15 13 2
15 13 3 15 9 13 2 16 13 13 3 7 16 13 13 2
11 3 13 3 2 16 15 1 0 13 2 2
14 3 3 13 9 13 9 9 13 2 13 3 9 0 2
16 3 16 13 7 13 9 9 2 3 3 3 15 9 13 13 2
7 2 13 15 13 9 9 2
8 3 15 15 3 10 9 13 2
3 13 3 2
9 9 15 3 13 3 13 3 13 2
10 15 3 3 0 15 13 0 9 0 2
16 3 3 3 3 13 9 9 0 3 3 13 0 9 7 13 2
24 13 15 9 13 0 0 2 10 9 2 15 9 1 9 13 0 2 0 3 9 13 13 3 2
16 3 1 9 9 13 2 15 15 13 9 3 0 7 9 0 2
19 3 0 3 0 13 0 9 2 15 3 3 3 9 3 13 7 9 13 2
8 15 3 15 13 13 7 0 2
29 3 3 15 3 9 0 1 13 2 7 3 15 9 13 0 3 13 7 13 9 1 0 7 0 1 0 9 2 2
27 3 3 16 9 13 0 9 2 3 15 13 9 3 13 2 16 1 9 0 9 0 0 0 9 13 13 2
14 3 3 3 13 0 9 2 15 15 13 13 9 9 2
23 15 3 15 13 1 9 13 0 2 16 15 9 0 9 9 9 13 13 0 1 9 9 2
19 3 0 3 0 13 0 9 2 15 3 3 3 9 3 13 7 9 13 2
17 15 3 15 13 3 7 13 2 7 13 13 0 7 0 9 0 2
29 3 16 3 3 13 9 9 0 3 3 13 0 9 7 13 2 13 2 16 15 15 13 7 13 2 9 1 0 2
8 13 3 15 3 3 15 3 2
19 3 15 0 13 2 3 3 13 2 16 3 3 0 0 0 9 13 2 2
7 15 3 3 13 9 9 2
18 2 3 3 13 2 9 3 13 9 2 16 3 15 3 13 13 2 2
7 3 3 13 13 0 9 2
8 15 3 3 1 9 13 13 2
16 3 3 3 9 3 13 3 9 1 9 0 1 3 13 13 2
21 9 3 1 9 7 9 13 9 7 9 7 9 9 13 9 1 0 13 9 13 2
7 3 3 13 13 0 9 2
7 3 3 15 3 0 13 2
10 3 3 9 0 13 13 9 0 9 2
14 3 9 13 1 0 3 2 16 15 13 1 0 9 2
21 3 15 9 7 9 7 9 0 13 0 2 15 3 15 9 13 2 9 3 13 2
36 13 3 15 9 3 2 16 3 3 0 0 0 9 13 2 16 3 9 3 13 2 15 9 0 13 2 15 15 0 13 13 3 13 3 2 2
16 3 13 2 13 3 9 0 9 2 7 15 13 9 0 13 2
14 15 3 3 3 1 9 0 0 13 2 13 9 9 2
18 2 3 3 0 3 13 7 3 0 13 2 0 3 10 9 13 13 2
20 3 15 3 13 7 13 2 15 3 15 3 0 13 2 16 15 9 0 13 2
20 3 3 15 9 13 0 2 3 3 15 0 9 1 9 0 2 7 0 2 2
8 3 3 13 13 0 9 3 2
8 15 3 3 1 9 13 9 2
37 13 3 9 0 9 7 3 9 2 7 3 15 3 3 13 1 9 3 13 9 2 9 3 13 1 0 9 2 13 7 13 2 0 9 9 13 2
16 0 3 1 13 9 0 2 15 3 1 9 9 7 9 13 2
9 15 3 1 9 0 13 9 13 2
6 15 3 13 3 3 2
43 16 3 3 13 0 9 0 15 9 9 13 2 16 0 9 13 2 3 3 3 13 1 15 15 9 13 0 3 13 2 13 3 13 0 9 2 15 3 3 13 9 0 2
29 3 3 3 0 3 9 13 13 2 3 9 3 3 9 2 16 3 3 3 3 13 0 0 9 7 9 13 2 2
7 15 3 13 13 9 9 2
17 13 3 0 0 3 2 16 15 9 9 9 0 9 3 3 13 2
12 15 3 3 9 13 2 15 3 0 7 0 2
17 16 3 3 15 13 9 1 9 9 2 13 1 9 13 0 9 2
7 1 3 15 10 13 2 2
15 13 3 3 15 3 9 9 0 13 9 2 1 0 13 2
42 3 3 9 13 0 9 2 3 10 3 9 3 9 3 13 9 2 0 3 0 9 0 13 9 2 0 7 0 2 1 3 9 13 9 0 0 2 9 3 3 9 2
7 7 3 9 9 13 9 2
14 13 15 9 0 2 13 1 9 2 0 2 3 0 2
6 13 3 3 9 0 2
6 3 3 15 13 9 2
18 12 3 13 0 2 13 3 3 9 2 13 3 3 7 1 9 13 2
17 13 3 3 0 7 13 0 2 9 3 3 15 3 7 9 13 2
21 0 15 3 9 9 13 9 9 0 2 3 13 9 2 0 1 0 9 13 9 2
10 9 3 13 2 13 0 9 2 13 2
5 3 0 9 13 2
9 1 3 9 13 7 9 13 0 2
9 1 3 3 9 13 2 16 13 2
10 13 3 15 9 3 0 9 9 13 2
5 0 3 13 9 2
7 15 3 3 13 3 15 2
22 1 3 9 3 9 3 9 3 13 1 0 2 9 3 3 15 3 13 1 9 0 2
9 0 9 13 2 7 15 13 0 2
17 10 3 3 0 13 1 9 0 9 2 9 3 13 0 7 13 2
8 1 3 15 9 13 0 0 2
8 9 3 13 0 3 0 3 2
8 0 3 9 13 9 0 9 2
46 3 15 9 13 3 13 2 3 3 15 9 1 9 13 9 3 13 7 3 13 9 9 3 2 15 3 9 9 13 2 15 3 3 13 7 3 9 13 2 0 3 0 13 9 9 2
13 15 3 1 9 13 9 9 3 1 9 9 13 2
6 13 3 15 9 13 2
10 3 3 3 15 13 9 13 9 2 2
12 3 13 13 9 2 13 3 9 9 9 13 2
16 0 3 13 9 0 9 2 1 3 9 13 9 3 7 9 2
5 13 3 3 9 2
18 1 3 9 3 9 3 13 9 3 0 7 9 9 2 0 9 13 2
18 7 3 9 13 9 7 0 9 2 13 3 3 13 1 0 9 9 2
22 13 16 3 0 9 0 13 2 15 15 13 1 9 2 16 0 9 13 2 9 13 2
7 15 3 3 3 0 13 2
17 0 9 13 9 0 9 2 13 3 9 2 13 3 9 0 9 2
22 7 3 15 3 13 13 7 9 13 9 10 16 15 0 0 9 9 13 1 9 13 2
11 3 3 13 9 2 7 15 9 13 0 2
8 3 3 0 9 13 13 2 2
17 3 3 15 13 13 0 9 1 9 0 13 2 1 3 9 13 2
13 3 3 1 9 0 13 2 9 3 1 9 13 2
19 0 3 15 9 13 0 13 9 13 9 2 3 3 9 7 9 13 9 2
19 15 3 3 3 13 0 9 2 3 3 13 3 3 13 0 1 9 9 2
11 9 3 3 13 2 15 15 13 0 9 2
19 3 3 3 3 13 2 9 3 13 9 0 2 15 15 0 1 9 13 2
25 3 3 3 3 9 13 2 13 3 2 7 13 1 9 13 0 2 1 0 3 13 9 9 13 2
11 15 3 13 0 9 1 9 3 7 3 2
26 7 3 16 0 9 13 9 1 9 2 0 3 1 0 13 2 3 15 1 9 9 13 3 7 3 2
16 3 3 3 9 9 13 13 2 3 3 3 9 9 13 13 2
25 15 3 9 13 13 2 9 13 2 9 3 13 9 13 9 2 13 3 1 9 0 13 3 9 2
9 3 3 3 15 13 3 3 13 2
11 3 3 3 13 2 13 3 15 3 13 2
10 13 3 2 15 9 1 9 13 0 2
22 3 16 9 13 9 2 3 13 13 1 0 9 0 1 9 2 0 3 3 13 2 2
17 3 3 13 9 9 13 2 0 3 3 1 9 13 13 9 13 2
6 0 3 15 9 13 2
19 3 3 3 3 13 2 16 3 9 9 15 13 2 3 15 13 0 13 2
11 3 3 3 13 2 13 3 15 13 0 2
17 16 3 3 3 9 1 9 13 2 3 3 13 7 13 9 13 2
20 3 16 3 15 9 1 9 13 2 13 2 16 3 3 15 1 13 0 2 2
29 16 15 0 13 1 9 7 1 9 2 13 3 1 0 9 9 9 2 0 3 0 3 2 0 2 13 3 0 2
8 15 3 3 3 13 3 3 2
6 3 15 9 0 13 2
22 3 9 1 9 9 13 2 9 7 9 13 2 9 3 13 2 15 15 13 0 9 2
19 3 3 9 1 9 13 2 0 3 0 9 13 2 9 13 2 13 13 2
13 13 3 9 9 2 13 3 9 1 0 13 9 2
17 2 3 3 0 0 13 13 1 9 2 1 15 3 9 0 13 2
10 3 3 3 3 15 13 13 9 2 2
18 3 3 13 13 9 9 2 13 3 1 9 2 3 15 0 9 13 2
15 3 3 10 0 9 13 9 2 13 3 13 7 13 0 2
23 13 3 1 0 9 2 1 3 9 13 2 16 15 9 0 13 0 9 9 7 9 13 2
17 3 12 9 12 3 9 9 0 13 2 0 3 15 9 13 9 2
20 3 16 3 0 9 0 13 9 2 3 3 3 9 3 13 7 9 13 0 2
15 15 3 3 3 13 9 0 3 13 2 0 1 9 13 2
17 3 16 0 13 0 3 13 13 2 3 3 9 13 1 9 9 2
16 13 3 0 9 1 9 9 0 13 2 13 3 0 9 9 2
9 7 9 9 13 9 3 9 3 2
18 3 3 9 13 9 7 0 9 2 13 3 3 13 1 0 9 9 2
27 2 6 15 2 16 3 9 0 13 13 9 2 7 3 15 9 13 13 2 9 3 3 13 9 0 3 2
32 3 3 3 9 0 2 3 3 9 13 0 2 0 3 13 9 2 0 3 9 2 7 3 3 13 9 13 0 7 13 9 2
12 3 3 15 13 13 9 1 9 9 0 13 2
6 0 3 15 13 9 2
48 16 3 3 3 3 13 2 16 3 13 9 3 9 9 3 9 2 13 16 15 3 13 9 9 1 0 13 0 13 2 7 15 15 3 9 13 0 9 1 9 2 0 3 0 13 0 9 2
10 13 3 2 16 15 13 0 9 2 2
20 16 15 0 13 1 9 7 1 9 2 3 3 15 0 9 13 0 1 9 2
16 0 3 9 13 13 9 2 15 13 13 2 16 0 9 13 2
19 3 15 3 3 13 2 0 3 15 3 13 13 2 3 3 15 13 9 2
6 15 3 0 9 13 2
16 3 3 3 0 1 9 13 9 2 16 3 9 13 0 9 2
25 9 13 2 15 3 13 3 2 13 3 2 1 9 13 2 16 3 13 9 3 9 9 3 9 2
35 3 16 3 9 1 9 0 13 13 2 3 3 15 13 9 0 2 0 9 2 7 1 9 13 9 2 13 3 13 7 13 0 1 9 2
11 0 3 15 13 2 13 1 9 9 9 2
27 0 3 3 13 3 0 9 9 15 15 13 13 2 3 3 15 3 0 3 9 0 3 9 13 0 13 2
7 9 3 15 13 13 2 2
27 3 13 2 15 3 3 13 0 9 2 13 3 9 2 3 3 15 13 9 2 15 3 13 1 9 9 2
10 15 3 3 0 9 13 9 3 0 2
15 13 3 9 0 2 9 3 13 0 1 9 3 9 3 2
15 15 3 3 0 7 0 13 13 2 9 3 15 0 13 2
20 3 16 3 3 13 7 1 9 9 13 2 3 3 3 9 1 15 13 9 2
24 7 15 3 1 9 0 13 2 3 3 13 0 9 1 9 2 3 3 3 9 13 9 0 2
13 15 3 1 9 13 9 13 2 13 3 0 9 2
9 13 3 3 13 1 0 0 9 2
6 15 3 15 0 13 2
24 16 3 3 1 9 0 9 13 2 3 15 3 9 3 0 7 0 9 1 9 13 13 9 2
9 9 3 1 9 0 13 9 1 2
37 16 3 3 1 9 13 7 0 9 9 1 0 13 2 16 15 13 9 7 9 2 0 3 15 9 13 2 13 2 16 9 9 7 9 13 2 2
8 3 3 15 13 13 0 13 2
6 13 3 13 1 9 2
8 15 3 1 9 13 1 13 2
10 0 3 3 13 9 2 1 3 13 2
25 15 3 3 3 3 9 13 9 0 13 2 3 3 3 9 13 9 13 2 3 3 9 13 3 2
7 3 3 0 0 13 3 2
5 15 1 9 13 2
8 3 3 9 13 9 0 0 2
33 7 3 16 15 9 9 13 0 9 1 9 2 15 3 13 9 0 2 9 9 13 2 16 3 3 3 13 2 3 9 9 13 2
19 15 3 3 9 9 1 9 13 2 16 15 13 0 0 9 0 9 13 2
13 3 15 3 3 13 9 0 9 9 7 9 13 2
33 3 13 13 9 0 2 13 3 9 2 3 9 9 2 1 3 9 13 9 2 7 13 9 2 7 9 13 9 2 7 13 9 2
19 3 15 3 3 9 13 3 13 2 9 3 3 13 2 9 1 9 13 2
5 9 3 13 0 2
36 15 3 9 3 9 13 9 9 2 13 3 3 1 9 2 7 15 1 9 13 2 13 9 0 9 2 15 15 9 3 13 2 13 3 9 2
7 15 15 13 13 0 9 2
30 9 3 15 13 0 0 2 15 3 9 3 13 2 3 13 0 3 0 13 2 15 3 15 13 2 15 3 15 13 2
16 1 3 3 0 9 9 13 0 2 13 3 9 7 0 9 2
7 3 13 13 1 9 13 2
19 3 15 15 9 3 13 2 16 0 13 2 16 3 3 3 3 9 13 2
17 3 3 15 13 9 1 9 0 9 2 3 15 9 13 3 0 2
23 3 3 13 9 0 9 1 9 7 9 13 2 15 3 13 9 3 7 9 7 9 0 2
18 10 3 3 3 13 13 0 9 3 2 3 13 9 9 0 3 13 2
25 3 3 9 13 3 3 3 9 13 3 3 9 13 2 7 3 9 13 0 2 0 3 13 9 2
8 15 1 13 9 9 9 0 2
8 3 13 9 2 16 13 9 2
5 13 3 3 13 2
12 15 3 1 9 13 1 0 9 9 13 0 2
17 15 3 3 13 13 1 0 9 1 9 2 3 15 13 9 0 2
9 15 3 3 3 13 0 9 13 2
9 3 3 15 0 13 1 0 13 2
11 15 3 3 13 0 9 13 1 9 13 2
3 3 13 2
8 13 3 0 9 13 9 0 2
8 15 3 0 13 7 13 9 2
2 13 2
9 3 13 9 13 2 15 3 13 2
17 15 3 3 3 9 0 0 13 2 9 3 13 13 3 1 9 2
8 9 3 1 9 13 9 0 2
30 7 15 3 13 0 1 9 2 9 3 1 9 13 0 9 0 2 1 3 9 13 2 1 3 9 13 9 1 0 2
5 9 3 13 9 2
14 13 3 0 1 9 0 9 2 16 13 1 0 9 2
12 15 3 13 9 7 9 0 2 13 3 13 2
5 9 3 13 9 2
22 15 3 3 13 2 13 3 9 7 0 2 3 0 2 1 15 3 3 0 13 0 2
34 15 3 16 3 9 9 0 13 2 3 3 3 9 13 0 2 0 3 9 0 13 3 3 13 13 2 3 10 3 9 3 13 9 2
11 7 15 3 13 9 1 0 13 9 0 2
20 15 3 1 9 9 9 13 7 13 0 9 2 13 3 1 9 3 9 13 2
23 3 16 13 3 13 3 9 0 2 3 13 1 9 9 2 3 3 9 1 9 13 9 2
19 3 16 9 13 9 3 7 0 2 9 15 3 3 13 2 1 9 13 2
7 15 3 9 0 13 9 2
8 3 10 3 0 13 9 9 2
7 9 3 13 1 0 9 2
9 0 3 13 2 0 3 13 9 2
6 15 3 1 0 13 2
15 15 3 13 0 9 2 13 3 13 1 9 7 1 9 2
8 3 3 3 9 13 1 0 2
24 3 13 9 13 0 9 2 1 0 3 9 9 13 9 0 9 2 16 13 1 9 9 9 2
23 13 3 13 3 3 9 0 9 13 2 15 3 13 13 7 13 2 1 3 15 9 13 2
11 3 9 9 0 13 13 2 0 3 13 2
4 9 3 13 2
15 0 3 0 13 13 9 2 13 3 3 0 1 9 13 2
6 0 3 9 9 13 2
13 15 3 9 9 1 9 13 7 1 9 13 9 2
5 13 3 3 13 2
26 15 3 13 9 2 7 9 13 13 9 9 2 7 3 9 3 0 13 2 16 13 9 7 9 13 2
21 3 3 15 13 13 0 13 2 13 9 3 0 2 16 15 9 13 13 9 9 2
7 3 0 7 0 13 9 2
8 9 3 15 2 7 9 13 2
16 3 3 15 9 3 9 13 1 15 2 13 15 9 9 13 2
5 9 15 13 13 2
13 9 3 3 0 9 1 9 9 0 9 13 13 2
21 13 3 3 3 2 0 3 15 13 9 2 15 9 3 3 13 15 0 9 13 2
6 0 3 15 9 13 2
7 0 0 13 9 9 9 2
13 3 3 15 3 9 13 0 3 9 9 1 9 2
14 3 3 3 13 9 2 16 3 3 3 3 13 0 2
12 3 3 13 13 2 7 3 0 9 13 3 2
24 15 3 0 0 13 1 0 13 2 15 3 0 3 15 13 9 2 15 15 9 7 9 13 2
19 9 3 15 13 2 13 3 9 13 2 16 15 3 9 9 13 3 13 2
8 15 3 3 9 0 0 13 2
12 3 3 15 15 13 2 15 3 13 13 3 2
27 3 3 2 16 0 3 9 7 9 13 2 3 3 3 9 13 3 3 15 0 2 15 13 9 0 13 2
11 9 3 15 13 2 13 3 15 9 9 2
7 13 3 7 0 0 13 2
5 3 13 9 13 2
9 3 3 3 15 0 13 13 9 2
20 3 13 0 9 0 9 3 3 13 2 15 3 9 9 1 9 13 9 13 2
17 13 3 3 0 1 9 2 0 2 3 3 15 15 9 13 0 2
13 3 15 15 0 13 3 13 2 15 3 13 13 2
17 1 3 9 13 0 9 3 0 3 2 9 3 0 3 0 3 2
27 1 3 3 15 9 3 9 3 9 13 2 13 3 0 1 9 0 9 2 13 3 3 15 13 9 9 2
8 3 3 3 0 13 0 9 2
8 3 3 0 1 9 13 9 2
8 3 3 3 3 15 3 13 2
13 3 13 2 15 3 3 13 2 13 3 3 9 2
26 3 10 1 9 9 13 0 9 9 2 15 15 9 7 0 13 9 2 1 9 3 13 9 9 0 2
42 3 16 3 0 13 7 3 13 2 1 3 9 13 15 15 13 9 9 2 15 3 9 13 9 13 0 3 13 7 0 2 1 3 9 0 13 9 2 0 9 0 2
34 3 3 3 15 9 13 9 9 9 2 15 9 13 7 9 9 9 0 2 0 3 9 13 2 3 3 15 13 9 9 3 7 9 2
13 13 3 3 13 1 9 9 2 9 7 9 13 2
4 13 3 9 2
7 3 3 3 0 0 13 2
15 3 0 3 9 2 15 9 13 2 9 15 9 13 0 2
19 3 3 3 3 15 0 13 13 2 3 3 9 13 2 15 9 0 13 2
16 6 3 15 15 9 13 13 3 13 2 7 15 13 3 13 2
23 3 13 2 15 3 3 15 3 3 13 7 13 2 1 3 3 9 13 9 3 9 3 2
11 3 3 15 13 7 13 9 0 9 3 2
6 0 3 9 13 0 2
6 3 9 0 0 13 2
29 9 3 13 13 0 1 9 2 13 3 9 9 2 1 3 13 0 2 13 3 9 2 9 3 13 1 3 13 2
11 3 3 3 13 2 13 3 15 3 13 2
20 3 1 3 3 9 13 7 9 9 2 3 1 0 1 9 7 9 3 13 2
5 15 3 9 13 2
6 9 3 9 9 13 2
6 0 3 9 13 0 2
24 3 3 9 13 9 3 3 9 2 7 9 7 9 9 7 9 0 2 15 13 0 13 9 2
10 15 13 9 0 2 16 15 3 13 2
7 3 3 13 0 1 9 2
8 7 3 15 3 13 0 13 2
5 3 3 15 13 2
6 9 3 15 13 0 2
17 3 15 3 13 13 0 1 9 9 0 2 16 3 15 3 13 2
16 7 15 15 13 0 9 13 3 13 2 13 3 15 9 0 2
17 3 3 15 3 13 1 9 9 2 15 15 13 0 3 7 0 2
29 3 3 0 13 2 15 15 0 3 13 2 15 3 3 0 9 7 9 13 2 9 13 2 16 3 0 9 13 2
8 13 0 9 9 1 9 9 2
9 1 3 9 13 2 3 3 9 2
16 3 13 13 9 2 1 15 3 15 3 13 7 13 9 9 2
11 3 3 0 13 2 3 3 9 13 0 2
15 3 3 3 15 13 15 13 9 9 2 0 9 9 9 2
20 3 16 3 15 9 13 7 9 2 3 3 9 13 2 16 3 13 9 0 2
6 9 3 15 13 3 2
16 3 3 9 0 9 13 0 2 15 15 3 13 13 0 3 2
22 15 13 9 1 9 9 13 0 2 16 0 9 13 13 3 2 16 3 3 3 13 2
8 3 3 13 13 9 0 9 2
7 15 3 3 13 9 9 2
11 15 3 3 3 13 2 3 3 13 9 2
19 15 3 3 13 2 16 3 13 0 0 3 9 3 2 9 3 13 9 2
17 13 3 9 7 15 0 9 13 0 9 2 3 3 13 0 9 2
7 3 3 13 9 9 0 2
19 3 3 3 15 13 2 16 3 3 3 13 13 2 3 15 13 0 9 2
10 3 13 13 2 15 3 13 9 9 2
7 0 3 3 3 13 0 2
5 13 3 3 9 2
11 15 3 3 13 0 9 16 0 9 13 2
34 15 3 16 3 0 9 0 9 13 2 13 3 1 9 2 9 3 15 1 13 0 0 2 15 3 1 9 9 13 9 3 13 3 2
7 0 3 1 9 0 13 2
17 9 3 0 9 13 2 16 0 9 13 2 9 3 3 9 13 2
9 15 15 9 13 7 3 9 13 2
7 3 3 9 13 3 13 2
23 3 3 9 0 9 13 0 13 9 2 16 15 9 0 13 13 3 9 7 13 15 13 2
12 3 3 15 9 0 3 13 3 1 0 9 2
14 3 3 15 13 9 2 15 15 9 7 9 13 2 2
19 3 13 9 0 2 15 3 9 13 2 3 3 15 9 13 3 3 13 2
17 3 3 0 15 3 9 13 2 3 3 13 13 15 3 3 13 2
15 9 0 15 3 13 0 9 0 13 2 16 15 13 9 2
8 3 3 13 13 9 9 3 2
8 15 3 3 1 9 13 9 2
13 15 3 3 9 0 3 13 13 1 9 1 15 2
7 13 3 0 9 9 13 2
11 15 3 3 13 2 3 3 15 9 13 2
15 0 3 9 1 0 0 9 13 2 16 3 3 3 13 2
7 9 3 0 13 1 9 2
17 9 3 9 13 0 2 1 3 9 10 0 15 3 13 9 9 2
11 3 15 3 13 9 0 2 13 3 0 2
8 9 3 13 9 3 9 3 2
27 15 3 9 13 9 2 7 15 13 2 16 3 15 1 9 13 0 2 0 3 3 9 1 9 9 13 2
33 3 0 1 9 13 3 7 13 1 3 0 9 1 3 0 9 7 9 2 15 15 3 9 3 13 13 9 2 16 13 1 9 2
11 3 3 3 15 9 3 3 0 13 0 2
9 15 3 3 13 3 9 9 13 2
29 3 3 13 13 0 9 9 1 0 2 13 3 9 0 2 13 3 1 9 7 0 9 2 13 3 9 0 9 2
8 3 9 9 1 9 13 0 2
12 0 3 15 9 13 13 2 16 0 9 13 2
14 3 3 3 9 9 13 7 9 9 1 0 0 9 2
8 0 3 9 0 9 3 13 2
17 9 3 0 1 0 13 9 2 0 3 1 9 2 0 3 9 2
25 0 3 3 7 0 9 13 2 15 9 13 13 9 9 13 0 9 2 0 13 7 0 9 0 2
9 3 3 9 9 13 13 7 13 2
4 0 3 13 2
20 0 3 3 9 0 1 9 13 13 9 1 9 13 2 13 9 1 9 9 2
7 0 3 9 13 0 9 2
13 1 3 15 13 9 9 3 13 0 7 9 0 2
6 1 3 9 13 3 2
13 3 3 3 9 13 15 3 13 2 0 3 13 2
12 3 3 3 9 13 9 13 2 0 3 13 2
13 3 3 0 9 1 0 9 0 13 2 0 13 2
9 0 3 1 9 9 13 0 9 2
7 3 13 13 9 0 9 2
15 3 16 3 0 0 13 9 2 3 1 9 13 9 1 2
19 13 3 9 9 7 9 13 9 0 9 2 15 0 13 2 16 13 9 2
19 1 3 3 9 13 9 9 9 2 7 3 3 3 0 3 13 0 9 2
10 15 3 3 13 2 9 1 9 13 2
4 13 3 13 2
20 15 9 0 13 13 2 7 9 13 0 9 1 9 9 3 15 15 9 13 2
17 3 15 9 13 9 13 0 2 16 3 3 0 1 9 13 2 2
12 3 13 1 3 13 1 9 1 9 1 9 2
8 15 3 3 0 3 13 9 2
8 15 15 3 13 13 7 13 2
31 3 3 3 9 3 1 9 0 13 13 2 15 3 9 13 9 13 2 16 3 9 0 13 2 15 3 9 3 0 13 2
9 9 3 9 9 13 3 13 2 2
14 9 3 0 9 13 13 0 0 1 0 9 2 13 2
6 1 3 0 13 9 2
14 9 3 0 9 13 13 2 9 0 13 2 13 13 2
7 3 3 9 13 9 9 2
16 3 13 2 9 3 9 9 13 2 13 3 3 0 13 9 2
18 3 16 13 3 13 3 2 0 13 9 2 15 3 9 13 7 13 2
7 3 3 13 13 3 13 2
64 3 3 9 1 0 13 9 1 9 13 7 9 13 9 0 2 3 3 3 1 9 13 2 16 3 10 9 1 9 7 9 9 1 0 0 0 9 13 13 3 2 16 3 3 3 13 2 3 3 15 3 3 0 7 9 13 2 16 3 15 0 9 13 2
21 3 3 3 13 2 15 15 9 1 9 3 0 13 13 9 2 16 15 13 9 2
17 16 3 15 0 3 1 9 13 2 0 15 3 15 3 9 13 2
24 3 3 10 3 3 9 13 0 15 2 16 13 0 9 2 13 3 1 15 13 3 3 15 2
29 16 3 3 15 3 0 13 13 9 2 3 15 13 2 16 15 1 13 2 7 3 9 3 7 0 9 9 2 2
7 15 3 13 13 9 9 2
22 3 3 15 3 0 13 2 15 9 0 13 2 3 9 3 3 9 2 7 0 9 2
15 15 15 15 13 3 13 9 9 2 15 3 1 9 13 2
18 3 3 3 3 3 3 15 0 13 2 0 3 3 0 9 9 13 2
8 3 15 3 13 13 13 3 2
54 3 3 15 0 1 9 0 0 13 2 15 3 13 15 13 9 7 3 13 7 1 9 9 13 2 7 3 15 9 3 13 9 2 15 3 3 3 13 13 7 13 2 1 3 15 0 13 0 13 2 7 13 13 2
16 13 15 3 13 9 9 0 2 9 3 7 0 0 9 2 2
19 3 13 2 10 3 3 0 13 7 13 13 10 9 2 16 1 9 13 2
6 0 3 13 9 9 2
7 15 3 9 0 13 9 2
18 13 3 9 3 9 3 9 13 0 2 15 3 0 13 1 0 9 2
7 7 15 13 9 0 13 2
6 15 15 15 9 13 2
9 3 3 13 1 9 13 3 13 2
7 15 3 13 13 9 9 2
10 0 3 15 13 15 15 13 7 13 2
13 3 3 15 0 13 3 3 9 3 3 0 9 2
18 3 0 3 0 13 0 9 2 3 15 9 3 13 9 9 3 13 2
9 3 0 3 3 9 1 9 13 2
18 3 3 0 13 0 2 9 3 3 9 13 2 15 15 0 13 9 2
26 3 16 3 0 15 13 9 13 2 3 3 3 15 13 13 13 9 1 9 2 7 3 9 13 0 2
24 12 3 7 12 3 13 9 13 2 0 3 13 9 0 9 0 2 13 3 15 0 9 0 2
37 3 3 13 3 13 9 0 2 15 15 13 9 9 2 15 15 13 9 13 9 2 13 3 9 0 2 3 3 15 9 13 1 9 0 13 13 2
6 15 3 3 9 13 2
19 3 15 3 13 15 9 13 2 16 15 9 0 13 13 9 3 7 9 2
17 3 3 15 13 13 9 1 9 2 9 1 0 13 7 0 9 2
26 3 13 13 3 2 16 13 1 9 2 3 3 15 13 9 0 2 0 9 2 7 1 9 13 9 2
11 1 3 13 13 2 1 3 0 9 13 2
15 15 3 3 0 9 13 1 9 13 2 3 3 9 13 2
7 9 3 9 1 0 13 2
16 3 3 1 9 0 13 9 13 0 7 1 9 7 0 9 2
9 13 3 9 7 15 0 9 13 2
16 0 3 1 9 0 13 9 13 2 1 3 0 13 13 9 2
3 15 13 2
16 15 3 3 15 9 13 0 2 7 3 3 13 0 13 13 2
6 3 3 3 0 13 2
18 15 15 9 13 3 7 0 9 7 13 1 9 7 15 15 9 13 2
8 0 15 13 3 9 13 2 2
7 15 3 13 13 9 9 2
25 15 3 3 15 13 1 0 13 2 7 15 3 13 13 13 3 2 16 3 3 15 9 13 13 2
10 0 3 3 13 1 9 9 9 2 2
14 9 3 3 15 7 9 13 2 16 3 13 3 13 2
8 0 3 15 3 15 13 9 2
7 3 0 0 9 9 13 2
17 7 3 15 3 13 7 1 9 13 9 10 0 7 13 3 3 2
17 13 3 3 0 1 9 0 0 9 0 7 9 13 9 9 2 2
21 3 13 2 13 3 9 0 9 2 13 3 3 13 2 9 3 13 1 3 13 2
17 15 3 3 1 0 9 0 9 13 2 15 3 3 9 13 2 2
8 3 15 3 0 1 0 13 2
26 13 3 9 0 0 9 1 9 13 7 9 0 0 13 2 13 3 3 9 9 3 13 0 3 13 2
10 15 3 13 1 9 9 1 9 13 2
6 13 3 15 9 2 2
9 3 13 2 15 3 0 13 13 2
17 9 3 3 13 9 9 0 2 1 3 9 9 9 13 7 9 2
23 3 3 9 13 0 9 2 13 3 1 9 9 9 9 2 3 3 3 0 13 0 9 2
8 13 3 13 1 0 9 0 2
8 3 13 13 9 7 9 0 2
10 3 3 13 9 9 3 7 9 13 2
9 0 3 3 13 13 9 9 0 2
39 15 3 3 9 0 13 9 9 3 7 9 7 15 0 7 0 13 13 2 16 3 9 0 0 13 0 3 0 3 7 13 9 0 2 15 9 13 9 2
20 9 15 2 3 13 15 15 2 13 13 0 9 2 7 1 0 7 0 9 2
9 9 3 13 2 7 13 0 13 2
11 15 3 2 3 10 3 3 2 13 9 2
21 3 3 3 3 3 15 0 2 15 3 0 9 13 2 3 13 0 13 1 9 2
24 3 3 9 0 13 1 9 0 0 2 9 3 12 7 12 13 1 9 2 0 3 13 0 2
8 3 3 0 13 9 3 13 2
6 15 3 3 0 13 2
5 9 3 0 13 2
22 3 10 0 0 9 0 1 9 0 13 2 16 9 1 9 13 2 3 3 15 13 2
15 15 3 3 9 1 13 9 13 2 3 9 13 13 2 2
11 3 3 13 13 2 15 3 3 13 0 2
6 9 3 13 0 9 2
8 3 3 1 0 15 3 13 2
11 3 3 13 3 13 9 0 1 0 9 2
12 13 3 3 9 3 7 9 7 9 9 13 2
17 15 3 9 12 9 13 2 12 3 0 9 2 12 3 9 9 2
11 15 13 1 3 13 2 13 3 9 0 2
20 9 3 3 13 13 0 9 2 15 1 9 13 2 13 3 0 3 0 3 2
9 9 3 13 2 13 3 0 9 2
15 15 3 3 9 13 9 0 0 9 2 1 9 0 13 2
16 1 3 1 9 13 9 0 0 1 9 7 13 9 13 9 2
18 1 3 13 9 0 3 9 2 1 3 9 9 2 13 16 9 13 2
9 15 3 1 9 0 13 9 13 2
17 3 3 15 13 13 9 9 9 1 0 2 16 13 0 9 13 2
15 3 3 3 13 9 9 9 3 7 9 9 0 1 9 2
6 0 3 9 13 0 2
17 3 9 0 0 9 13 9 0 1 9 13 2 13 3 0 9 2
8 13 3 9 1 9 9 13 2
21 3 3 16 13 13 9 9 2 9 13 9 1 9 13 7 9 0 13 13 9 2
22 3 16 3 13 7 13 13 9 10 0 2 16 13 9 2 3 9 1 9 13 13 2
6 3 3 9 0 13 2
15 3 3 9 13 9 0 9 3 2 15 9 0 13 9 2
10 3 3 13 13 2 15 3 3 13 2
18 1 3 1 9 13 9 0 2 9 3 13 9 7 13 1 9 9 2
16 13 3 15 0 9 15 3 10 0 9 10 0 2 0 13 2
14 13 3 13 1 9 2 3 3 13 0 9 2 0 2
9 1 3 13 0 0 3 7 0 2
9 15 3 3 3 0 3 13 9 2
7 15 3 1 9 13 9 2
9 15 3 3 0 3 13 13 9 2
9 15 3 13 3 0 13 9 0 2
17 0 3 1 9 9 13 9 2 0 13 9 13 2 15 3 13 2
6 15 3 9 0 13 2
8 15 3 3 9 13 0 0 2
7 9 3 9 0 0 13 2
11 3 3 15 9 13 2 7 0 13 0 2
20 3 3 15 3 15 13 0 0 9 9 3 13 2 16 3 3 0 13 2 2
9 0 3 13 13 7 13 9 2 2
18 3 16 10 3 13 0 9 9 2 13 3 1 0 13 7 9 13 2
6 13 3 15 13 9 2
10 3 3 13 2 13 3 1 9 9 2
19 15 3 9 3 0 13 2 7 3 3 9 3 13 7 0 13 9 2 2
7 15 3 13 13 9 9 2
6 3 3 9 13 2 2
9 15 3 3 3 13 13 0 9 2
4 0 9 13 2
23 0 3 3 3 9 0 13 9 2 3 9 9 9 13 2 15 3 3 1 0 13 13 2
20 15 3 3 13 9 0 2 1 3 13 13 2 13 3 1 9 9 3 13 2
11 13 15 9 1 9 0 13 3 1 9 2
25 15 3 3 9 9 2 3 15 3 13 2 7 1 0 13 13 2 16 9 3 13 9 3 0 2
7 3 3 13 9 7 9 2
11 0 3 13 9 3 9 0 3 9 13 2
11 3 3 3 2 0 0 13 2 13 9 2
10 0 3 9 2 13 3 15 13 2 2
22 13 3 7 0 9 13 13 9 0 7 0 2 0 3 0 3 16 0 9 13 0 2
12 15 3 13 13 0 1 9 2 13 3 9 2
10 15 3 13 9 0 3 13 1 9 2
15 13 3 9 9 9 9 13 2 9 3 13 1 3 13 2
7 15 3 13 15 3 9 2
12 3 15 9 15 3 13 2 3 3 13 2 2
6 7 3 3 13 9 2
6 9 3 15 15 13 2
5 15 3 13 13 2
19 0 3 0 3 7 0 13 9 2 15 15 9 9 13 9 9 1 0 2
6 15 3 0 0 13 2
18 10 3 0 3 3 15 13 3 3 13 2 7 13 13 7 13 3 2
11 0 3 3 0 13 2 1 9 0 9 2
7 3 3 9 13 0 13 2
21 0 3 9 13 13 1 9 9 0 2 16 3 3 0 9 3 13 7 13 9 2
14 0 3 15 9 13 9 9 1 9 2 16 13 0 2
18 10 3 0 15 13 0 0 13 2 0 3 9 13 1 9 9 13 2
16 3 3 3 3 13 0 9 2 3 3 1 9 13 1 9 2
10 13 3 9 13 2 16 15 13 13 2
9 9 3 13 0 3 0 15 9 2
9 0 13 9 16 15 15 13 9 2
16 3 3 3 13 9 1 0 2 16 3 9 1 9 13 0 2
7 3 15 0 9 13 2 2
11 3 13 2 15 3 3 0 3 13 9 2
7 9 3 15 0 13 13 2
36 3 3 9 13 0 3 3 9 2 7 9 3 13 7 9 0 2 3 3 15 9 3 0 9 3 9 3 9 3 0 9 3 0 7 9 2
17 9 3 15 3 13 9 0 13 2 15 3 13 1 0 9 2 2
15 3 13 9 0 2 13 3 9 13 9 0 9 1 9 2
24 9 3 0 12 0 13 0 2 15 1 9 3 13 0 2 13 3 9 2 0 3 13 9 2
9 9 3 3 13 13 9 0 9 2
7 15 3 3 13 1 0 2
15 1 3 9 9 13 2 0 9 2 13 3 9 0 9 2
10 3 9 9 13 9 2 13 3 9 2
13 3 3 15 9 13 9 2 15 15 13 13 9 2
35 9 3 16 3 0 9 13 2 13 3 13 1 9 0 9 13 2 1 3 13 9 0 9 2 13 3 9 0 0 2 16 0 3 13 2
29 3 16 3 13 9 13 9 2 13 3 13 1 9 2 3 15 0 9 13 2 1 3 3 9 13 9 9 3 2
25 0 3 3 1 9 13 2 3 9 0 2 15 3 3 3 15 3 3 13 2 3 3 9 9 2
5 1 3 0 13 2
14 3 3 9 13 0 9 2 16 13 9 9 3 13 2
12 13 3 13 1 9 0 9 13 9 0 9 2
20 15 3 1 9 13 2 1 3 3 15 13 9 2 9 3 13 1 3 13 2
9 3 13 2 15 3 0 13 13 2
7 15 3 1 9 13 13 2
18 1 3 9 0 13 9 9 2 3 3 15 13 9 13 3 3 13 2
14 0 3 15 13 0 0 2 3 13 16 9 9 13 2
9 9 3 15 9 13 13 3 9 2
9 13 3 13 1 9 0 13 9 2
11 13 3 1 9 2 9 3 15 0 13 2
9 0 3 13 2 13 3 0 9 2
19 7 13 2 3 15 3 13 1 9 1 0 9 13 2 15 3 13 13 2
14 3 3 15 3 13 3 3 13 3 3 3 3 13 2
6 3 3 13 0 13 2
11 3 13 2 10 3 13 9 1 0 9 2
14 13 9 0 2 13 9 9 2 13 3 9 0 9 2
8 0 3 9 13 9 3 0 2
12 0 3 3 13 9 9 9 9 13 9 9 2
9 3 3 15 13 13 1 0 0 2
25 13 3 0 0 2 16 3 3 9 13 0 13 9 0 3 13 9 15 9 13 2 0 13 9 2
8 3 15 3 0 1 0 13 2
10 3 13 2 1 3 9 13 0 9 2
15 3 3 9 9 13 2 13 3 3 9 0 16 13 9 2
7 7 15 13 9 0 13 2
7 15 3 3 13 0 0 2
18 15 3 15 15 13 1 0 9 2 16 3 9 13 9 7 9 13 2
7 15 3 13 3 0 0 2
11 2 3 13 3 3 13 0 9 13 2 2
7 3 13 9 13 9 9 2
29 15 3 16 1 9 13 2 0 3 13 2 3 13 15 3 3 13 2 10 3 3 9 13 0 9 2 1 9 2
6 0 3 9 13 0 2
15 9 3 9 7 9 13 3 13 2 16 15 3 15 13 2
41 15 3 16 3 9 0 1 9 13 2 0 2 15 15 9 13 0 2 15 0 13 1 9 0 13 3 2 15 3 1 9 3 13 3 13 2 16 9 9 13 2
17 3 16 3 9 1 9 13 2 13 3 3 1 9 9 0 13 2
14 9 3 13 0 13 1 9 2 0 3 1 9 13 2
8 3 3 3 9 13 0 9 2
6 9 15 13 13 2 2
15 3 13 2 13 3 0 9 9 2 3 3 9 0 13 2
8 10 9 3 15 13 13 13 2
14 12 3 1 9 0 9 9 13 2 0 3 15 0 2
13 15 15 0 9 0 7 9 7 9 9 13 0 2
18 3 3 0 13 0 2 16 1 9 9 13 1 9 13 13 1 9 2
18 9 3 15 0 13 9 7 9 2 16 3 15 9 1 9 13 2 2
7 0 3 15 0 13 2 2
14 3 13 1 9 13 9 0 7 15 13 9 0 13 2
14 9 3 16 3 15 13 0 2 3 15 13 13 9 2
20 15 3 9 9 3 13 7 9 13 13 2 16 3 3 0 1 9 13 2 2
7 15 3 13 13 0 9 2
19 3 3 15 15 9 3 9 3 13 0 2 15 3 15 13 13 9 2 2
9 13 3 3 1 9 13 9 0 2
10 13 3 9 2 7 15 0 9 13 2
9 7 15 3 1 9 13 9 0 2
13 13 3 3 9 0 9 9 1 0 13 0 9 2
14 15 3 13 0 9 9 2 13 3 13 1 0 9 2
8 3 3 3 9 13 9 9 2
9 1 3 0 13 9 0 7 9 2
36 1 3 15 9 9 13 2 13 3 9 2 16 13 3 13 3 3 13 0 9 2 15 15 9 0 3 13 2 9 3 13 7 9 9 13 2
26 3 15 15 15 9 0 0 13 2 0 2 16 15 13 9 0 13 1 9 9 3 0 3 9 2 2
16 3 13 2 9 3 1 9 13 1 9 13 9 0 7 0 2
21 15 3 0 9 13 1 9 0 2 1 3 3 9 13 2 1 3 9 13 13 2
10 9 3 9 9 13 2 13 3 9 2
16 1 3 0 9 13 0 3 9 2 7 15 13 9 0 13 2
31 2 0 3 13 9 2 3 3 1 9 13 2 16 15 15 1 9 13 2 16 3 3 13 0 9 13 1 9 0 2 2
12 3 3 3 15 9 13 13 1 3 9 13 2
23 15 3 3 3 13 9 0 9 2 16 3 15 13 3 13 2 16 3 13 9 9 0 2
10 3 3 15 9 3 9 3 0 13 2
28 15 3 16 3 9 13 7 13 9 2 1 3 15 9 0 13 7 9 2 1 3 9 13 9 1 9 13 2
28 9 3 9 1 9 13 13 3 1 9 9 3 0 2 13 3 9 1 9 13 2 7 15 13 9 0 13 2
7 15 3 13 13 0 9 2
12 3 3 15 3 3 9 3 13 3 9 0 2
10 13 3 7 1 9 13 1 9 9 2
12 13 3 3 0 0 9 2 1 9 0 13 2
6 7 15 13 13 3 2
24 0 3 9 0 9 9 0 13 7 9 2 16 3 15 9 9 13 2 13 3 9 9 2 2
13 3 3 13 2 9 3 13 1 9 13 9 9 2
8 15 3 13 2 13 3 9 2
9 15 3 1 9 0 13 9 13 2
16 3 16 9 7 9 1 9 13 2 3 3 9 13 0 9 2
31 3 3 3 13 7 9 9 13 0 2 15 0 13 1 9 2 15 3 1 9 9 13 0 9 9 13 15 3 9 13 2
25 16 3 3 15 0 1 9 13 2 3 15 0 13 9 2 16 3 15 0 9 13 9 9 2 2
8 0 3 15 9 1 9 13 2
14 3 15 3 13 2 15 3 0 0 13 13 1 0 2
23 9 3 13 13 2 16 9 13 0 0 9 2 3 13 0 0 0 9 9 7 9 13 2
14 13 3 16 9 13 9 0 3 13 2 0 9 13 2
13 3 3 0 9 13 13 13 3 3 1 0 9 2
6 0 3 9 13 0 2
11 3 9 13 2 9 3 13 1 9 9 2
8 3 9 0 1 9 9 13 2
6 3 3 9 0 13 2
15 2 13 2 9 9 7 9 2 9 3 3 13 9 0 2
8 3 3 3 0 13 15 13 2
20 1 15 13 3 7 13 9 9 2 1 15 3 3 3 13 0 9 10 9 2
7 3 3 15 9 9 13 2
16 1 9 9 3 9 3 13 9 2 15 3 0 3 13 9 2
13 3 3 3 3 15 13 9 0 15 3 15 13 2
6 13 3 15 0 13 2
32 3 3 3 15 3 0 13 9 2 3 0 3 3 3 0 2 16 15 0 13 2 7 1 0 13 2 16 3 13 2 9 2
18 3 3 9 9 13 2 3 3 15 9 13 2 15 3 0 9 13 2
27 3 0 13 9 7 9 9 2 7 0 13 9 7 9 9 9 2 7 9 0 9 13 9 7 9 13 2
21 13 3 0 9 0 9 1 9 13 1 0 9 13 2 0 3 15 9 9 13 2
5 3 13 10 9 2
16 13 3 15 15 13 7 13 1 9 0 9 7 0 9 13 2
17 15 3 9 3 13 2 13 3 9 9 2 16 13 3 13 9 2
7 15 3 13 13 0 9 2
9 0 15 15 0 1 9 13 13 2
15 0 3 0 9 9 13 0 13 2 16 3 3 13 13 2
10 15 0 15 3 2 15 3 0 13 2
27 3 3 9 0 13 2 16 3 15 13 2 15 3 7 3 13 1 0 9 15 9 13 3 3 9 13 2
16 13 9 9 2 15 0 9 9 13 2 7 15 9 9 13 2
5 13 3 9 0 2
26 0 3 0 0 1 9 13 1 9 2 15 3 3 3 1 9 3 9 3 2 0 2 7 0 9 2
11 3 3 15 3 0 9 13 0 0 13 2
18 3 3 15 3 13 9 2 0 9 2 1 9 0 2 13 9 13 2
9 7 0 3 3 9 1 9 13 2
24 3 0 0 0 9 3 3 9 13 2 16 3 3 15 3 0 9 9 1 0 13 1 9 2
18 6 3 3 15 3 9 0 0 13 2 15 15 9 13 1 3 13 2
10 3 3 15 9 13 2 13 3 0 2
18 1 9 3 9 7 9 0 13 13 2 16 3 15 15 13 13 0 2
18 3 3 3 3 15 0 9 13 15 13 2 15 3 0 0 3 13 2
11 13 3 0 9 7 9 13 9 2 0 2
15 3 3 3 0 9 9 13 15 0 2 16 9 0 13 2
14 13 3 13 9 1 9 0 2 13 3 0 0 9 2
17 16 3 9 13 7 13 0 9 2 3 3 13 13 0 3 13 2
14 3 3 9 13 3 2 3 3 3 9 13 13 0 2
9 12 3 1 0 9 0 9 13 2
9 10 3 0 13 9 3 9 3 2
16 2 3 3 3 13 13 9 2 0 1 9 2 0 13 9 2
26 3 3 3 15 3 9 13 9 2 16 15 10 0 9 3 0 13 2 15 13 1 9 9 1 13 2
19 9 3 13 9 9 9 9 9 0 2 1 3 9 13 9 3 7 9 2
5 13 3 3 9 2
17 15 3 3 13 0 2 9 3 15 3 3 7 3 13 9 9 2
16 3 15 3 1 9 13 2 13 9 2 0 3 3 13 3 2
18 3 12 9 12 3 9 0 3 13 2 3 9 3 7 9 9 13 2
26 3 16 3 0 9 0 13 9 2 9 13 1 3 9 0 13 13 2 15 3 9 3 9 3 13 2
9 3 3 3 0 13 1 0 9 2
15 3 15 9 9 3 13 9 7 9 13 2 13 3 9 2
11 2 3 3 3 13 0 9 9 1 0 2
12 3 0 13 9 9 2 15 3 0 9 13 2
18 3 3 1 9 13 7 13 9 2 3 3 9 13 0 1 9 9 2
33 3 16 9 3 13 7 9 2 3 3 15 9 13 13 13 2 15 15 9 13 1 9 9 13 9 12 13 2 0 9 3 13 2
8 15 3 3 13 13 9 9 2
15 3 3 3 9 13 9 9 0 2 7 15 13 9 13 2
18 15 3 15 1 9 13 13 9 2 9 3 1 0 1 9 13 13 2
19 3 10 0 13 0 9 13 9 13 0 2 16 3 15 9 13 9 13 2
17 15 3 3 13 7 1 9 13 2 3 3 13 0 9 13 9 2
8 2 3 3 3 13 13 9 2
33 15 3 3 3 9 0 3 3 9 2 7 15 3 0 9 13 9 1 9 0 2 13 3 0 9 7 9 2 3 3 0 13 2
19 2 9 3 0 1 9 13 2 9 9 3 3 1 3 3 3 2 0 2
7 1 3 9 0 13 0 2
23 3 3 3 9 9 13 2 3 3 15 13 9 2 15 3 1 9 9 13 9 9 13 2
26 3 3 3 9 13 3 3 9 2 7 15 3 0 7 0 9 0 9 13 2 13 3 3 0 9 2
13 3 3 3 15 0 3 2 13 3 3 0 0 2
6 3 3 0 9 13 2
5 1 3 9 13 2
16 3 13 2 7 15 9 13 9 1 0 2 3 3 13 13 2
17 9 3 1 9 0 13 2 3 3 9 3 13 2 13 3 9 2
23 3 3 15 10 9 13 9 2 3 3 3 9 0 13 1 9 13 2 16 9 0 13 2
16 13 3 9 13 9 0 2 1 3 3 0 13 1 9 9 2
7 3 3 13 13 9 0 2
14 2 16 3 9 13 0 9 2 9 13 13 1 0 2
16 3 0 9 7 9 0 13 1 9 2 1 3 3 13 13 2
7 3 3 13 9 0 9 2
13 9 3 15 13 12 2 1 3 0 12 13 9 2
6 15 3 12 13 0 2
18 2 3 3 3 0 9 1 9 13 13 13 9 15 0 7 9 0 2
11 3 3 3 9 13 9 0 2 3 13 2
18 9 3 1 9 13 3 13 2 9 3 0 3 9 9 3 7 9 2
16 3 3 9 13 7 1 9 13 2 3 3 13 1 9 9 2
16 16 3 9 13 0 9 2 3 3 15 9 13 1 0 13 2
17 15 3 3 13 7 1 9 13 2 3 3 13 0 9 13 9 2
23 3 16 3 10 9 13 3 13 2 3 3 1 9 9 13 1 9 2 0 2 9 0 2
14 1 3 9 0 13 0 9 0 3 9 7 9 0 2
14 3 3 9 13 0 2 15 3 10 9 0 13 3 2
12 3 3 1 0 13 2 7 3 13 0 13 2
26 3 3 9 13 0 2 3 3 13 9 3 0 2 7 9 0 0 9 2 15 3 13 0 1 0 2
8 13 3 1 9 0 9 9 2
7 15 3 15 13 0 9 2
8 3 3 3 3 13 0 13 2
23 3 3 15 13 9 0 9 13 0 13 9 2 0 2 3 3 9 3 13 3 3 9 2
20 2 3 3 1 9 13 2 3 3 15 3 13 2 7 13 9 1 0 9 2
7 13 3 1 9 13 0 2
12 9 3 9 13 2 13 3 9 9 7 9 2
28 3 15 3 0 9 13 9 9 13 13 3 2 3 3 3 1 9 0 9 3 7 9 9 13 13 0 9 2
9 3 3 3 13 9 13 0 13 2
23 2 3 3 9 13 13 7 3 0 9 13 13 2 13 3 15 3 13 2 16 13 13 2
19 13 3 0 9 9 0 2 16 15 0 13 2 1 3 9 13 9 13 2
8 15 3 13 13 1 9 9 2
10 3 3 13 9 0 3 13 2 0 2
14 3 3 15 3 12 7 12 9 0 0 1 9 13 2
6 0 0 9 13 9 2
30 3 3 0 3 13 0 9 0 1 9 13 13 2 0 3 3 13 1 9 2 16 15 13 13 13 7 15 0 13 2
20 3 16 3 13 13 10 0 9 2 3 3 9 13 7 13 2 13 3 15 2
5 3 13 0 9 2
24 7 15 1 9 7 3 13 2 0 3 9 2 1 9 2 15 3 13 9 13 0 0 13 2
19 2 3 13 2 15 3 3 13 0 9 2 13 9 3 0 0 3 0 2
8 3 3 3 15 9 13 13 2
23 2 2 15 3 3 13 0 0 9 1 0 9 9 2 3 13 2 0 9 0 9 13 2
6 3 3 9 13 13 2
9 0 3 13 9 7 13 9 0 2
25 15 3 3 13 10 0 9 13 2 16 15 13 9 7 3 3 13 9 2 15 3 9 9 13 2
21 9 3 15 13 2 9 3 9 9 3 9 3 2 0 2 15 9 3 0 13 2
17 3 3 9 9 0 13 3 3 9 9 2 16 3 0 0 13 2
20 3 3 3 15 9 9 13 13 3 3 15 3 9 2 16 3 9 15 13 2
19 2 3 13 13 2 15 3 3 13 13 0 2 7 15 0 13 0 9 2
19 2 2 9 3 15 13 9 9 1 9 13 0 1 9 9 2 9 13 2
6 9 3 1 9 13 2
8 3 15 1 15 13 0 9 2
10 1 3 9 3 13 2 13 3 9 2
8 15 3 1 3 13 13 9 2
16 15 3 13 13 9 9 2 0 9 13 2 9 3 13 9 2
22 3 16 9 0 13 9 0 9 13 7 1 0 9 13 2 13 1 9 13 1 9 2
28 15 3 15 13 1 9 9 3 13 2 9 0 13 1 9 2 13 1 9 2 3 9 9 13 2 9 13 2
6 0 3 15 9 13 2
9 3 3 3 3 15 13 0 9 2
14 3 3 3 13 9 0 9 13 9 0 2 15 13 2
8 3 3 3 13 13 9 0 2
20 3 16 3 13 13 10 0 9 2 1 3 15 3 3 3 12 13 13 9 2
12 13 3 9 13 0 9 2 3 13 9 0 2
10 0 3 9 1 9 13 0 9 9 2
10 2 15 3 15 1 9 0 13 9 2
11 9 3 13 0 9 1 9 2 0 0 2
8 15 3 13 2 16 13 13 2
8 0 13 9 2 0 9 13 2
16 15 3 0 3 9 15 13 13 7 13 9 2 13 3 13 2
5 15 3 0 13 2
14 15 3 13 13 9 2 3 3 13 13 1 9 0 2
18 3 15 3 3 13 13 1 9 2 15 3 1 9 13 0 3 0 2
24 3 10 0 9 13 13 2 15 15 13 15 1 9 13 13 1 9 2 16 15 0 9 13 2
20 15 3 13 15 3 3 3 13 0 13 2 9 2 3 15 0 1 15 13 2
7 0 3 13 0 9 13 2
29 3 3 1 0 9 13 0 9 0 3 2 3 3 15 13 0 1 9 2 7 15 13 2 7 3 9 3 13 2
20 3 16 3 13 13 10 0 9 2 1 3 15 3 3 3 12 13 13 9 2
15 3 3 15 9 13 3 13 2 9 1 9 13 0 9 2
12 15 3 3 9 13 2 16 15 13 3 13 2
6 15 3 13 3 3 2
10 2 3 13 2 15 3 13 7 13 2
12 13 3 3 0 0 13 7 15 13 0 3 2
24 8 13 15 3 0 2 7 15 0 9 13 3 3 2 16 15 13 0 2 15 3 15 13 2
15 3 3 9 13 0 9 9 0 2 7 15 9 9 13 2
8 7 15 9 7 9 13 9 2
12 2 3 13 2 3 15 3 15 13 0 9 2
10 3 3 13 13 2 3 3 13 9 2
16 3 16 9 1 9 13 9 2 3 3 3 15 9 13 0 2
12 9 3 15 13 9 7 9 7 0 0 9 2
14 2 9 15 0 13 1 0 9 2 10 3 0 3 2
6 15 3 15 9 13 2
21 2 13 7 13 13 0 2 3 3 13 13 0 9 2 1 3 15 9 13 9 2
8 9 3 13 9 9 3 0 2
5 15 3 13 9 2
13 3 3 15 10 9 1 9 13 0 2 16 13 2
12 9 3 0 9 13 2 16 15 15 13 13 2
33 3 16 3 3 10 9 0 1 9 13 13 2 0 3 13 2 13 3 3 2 3 3 15 3 13 1 9 2 3 3 9 13 2
6 3 9 13 0 9 2
13 15 3 9 13 0 2 0 1 9 2 9 13 2
30 15 3 3 13 13 2 3 16 15 13 9 0 9 9 2 15 3 3 3 13 9 13 3 2 15 3 13 0 3 2
16 3 15 1 9 0 9 13 13 2 15 3 9 13 0 13 2
18 0 3 15 9 3 7 9 13 9 9 13 2 13 3 15 9 9 2
15 0 3 0 13 2 1 3 13 9 2 15 3 13 13 2
9 3 15 9 13 9 13 9 0 2
26 15 3 3 13 1 15 9 13 2 3 15 9 0 13 2 15 3 15 1 13 1 9 1 9 0 2
9 3 3 15 15 9 9 0 13 2
10 3 3 15 15 0 13 9 7 9 2
10 2 15 3 3 1 9 13 0 9 2
8 2 15 3 13 9 0 13 2
27 16 3 3 3 15 15 13 0 13 2 9 3 3 3 13 9 0 13 2 7 15 3 13 9 9 9 2
32 9 3 13 3 7 13 9 9 13 1 3 9 13 9 2 0 3 1 9 13 9 13 2 16 15 3 1 9 13 13 3 2
10 3 3 3 15 13 1 9 0 13 2
19 3 15 13 2 16 3 0 13 2 16 15 9 9 9 7 15 0 13 2
6 0 3 0 3 13 2
9 15 3 15 1 9 0 13 9 2
15 15 3 1 0 9 13 2 10 3 0 3 13 13 9 2
7 12 3 0 9 9 13 2
10 3 9 9 0 3 13 13 13 9 2
8 3 3 3 13 13 9 0 2
23 2 16 3 9 13 0 9 2 3 3 3 3 13 9 9 2 0 3 13 0 1 9 2
4 9 3 13 2
12 9 3 9 0 13 0 9 13 9 0 13 2
12 0 9 9 13 3 9 13 7 15 0 13 2
7 15 3 13 13 0 9 2
31 3 15 3 3 13 13 9 2 3 0 0 13 0 9 9 0 13 2 0 3 9 9 13 2 0 3 3 13 13 0 2
13 6 3 13 0 3 13 13 3 0 0 9 13 2
28 3 3 15 9 3 1 9 3 3 13 13 1 9 2 1 3 3 0 9 13 0 2 15 15 0 13 9 2
10 2 3 13 10 9 1 15 13 3 2
17 13 3 0 1 9 3 7 9 0 1 9 13 2 13 3 9 2
18 3 3 10 9 9 2 0 9 2 0 13 13 2 16 1 9 13 2
15 0 3 0 9 13 2 15 13 9 2 15 3 13 13 2
26 3 15 3 13 2 1 3 9 13 0 2 13 2 7 13 3 0 9 0 1 9 13 13 0 9 2
17 15 3 3 13 7 1 9 13 2 3 3 13 0 9 13 9 2
17 3 16 0 13 2 0 3 13 13 2 3 3 15 9 13 0 2
8 3 15 9 13 7 9 0 2
24 3 15 9 13 0 9 13 1 2 9 3 13 13 13 9 2 16 1 9 13 2 9 13 2
5 15 3 13 13 2
15 3 16 3 3 0 9 13 13 2 3 3 3 9 13 2
9 3 3 9 0 9 13 3 0 2
20 16 3 13 15 7 13 13 2 1 3 13 15 9 7 0 9 9 0 13 2
4 0 3 13 2
18 2 3 13 2 7 3 13 0 0 9 2 7 15 0 13 13 9 2
15 3 3 15 9 0 7 0 13 3 13 2 0 13 9 2
18 3 3 15 13 0 3 7 0 7 9 9 13 2 16 15 13 9 2
12 15 3 15 9 13 2 9 3 0 13 13 2
22 0 3 2 16 3 13 2 13 2 3 3 15 0 3 3 9 0 3 3 0 9 2
10 2 3 13 13 2 15 3 13 9 2
30 3 15 3 3 0 0 9 13 13 13 2 13 3 9 0 2 1 3 13 1 9 0 0 2 13 3 9 0 13 2
7 13 3 9 13 1 9 2
11 15 3 3 13 9 2 13 3 9 13 2
43 2 3 16 3 10 9 13 2 3 3 0 9 0 13 0 2 3 3 9 13 13 2 15 13 3 2 9 3 3 13 13 1 9 2 1 3 3 0 13 1 9 9 2
17 9 3 9 0 1 9 13 13 2 16 3 15 15 13 13 0 2
11 9 3 15 0 0 9 9 13 13 3 2
16 15 3 1 9 9 0 9 2 15 0 13 2 13 9 13 2
20 15 3 3 13 0 2 7 15 3 13 16 13 0 9 0 7 0 0 9 2
18 2 3 3 3 0 9 1 9 13 13 13 9 3 0 7 9 0 2
16 16 3 9 13 7 1 9 13 2 3 3 13 1 9 9 2
21 16 3 9 13 0 9 2 3 3 15 9 13 13 0 3 13 1 3 0 13 2
17 15 3 3 13 7 1 9 13 2 3 3 13 0 9 13 9 2
16 2 3 3 3 13 13 9 2 0 1 9 2 0 13 9 2
12 9 15 3 0 13 0 7 9 7 0 9 2
8 15 7 1 9 15 9 13 2
18 13 0 9 2 0 7 9 0 3 9 7 0 13 7 0 9 9 2
12 15 7 3 13 13 9 3 3 0 9 13 2
9 13 7 0 1 0 9 13 13 2
13 13 7 3 3 9 2 13 9 9 0 7 0 2
17 15 7 1 13 9 3 0 1 9 2 13 9 0 1 0 9 2
38 16 3 3 9 7 7 9 0 13 9 7 9 0 0 9 7 9 2 3 7 13 9 0 13 3 9 9 0 2 3 15 9 13 0 9 13 3 2
11 13 7 9 9 7 9 9 9 1 0 2
6 15 7 13 9 9 2
28 3 3 3 1 9 9 9 13 13 9 1 9 13 2 7 3 9 7 9 0 13 13 2 7 9 13 9 2
12 9 3 13 2 7 3 13 9 2 15 13 2
7 15 7 3 13 0 0 2
5 7 3 13 9 2
3 7 13 2
6 15 7 9 13 9 2
12 3 3 3 15 13 7 13 13 1 9 0 2
11 15 7 1 9 0 13 9 13 3 13 2
10 7 3 15 13 3 3 0 13 9 2
19 3 7 9 13 16 10 0 3 9 13 2 10 13 2 15 13 9 13 2
5 7 13 9 13 2
12 3 7 1 9 3 13 0 9 0 16 9 2
9 15 7 9 0 7 0 13 9 2
23 13 3 3 0 9 13 9 9 7 0 9 13 1 9 9 7 0 9 9 13 0 9 2
25 7 15 9 13 13 0 7 9 2 16 3 3 3 9 0 13 9 2 15 3 9 0 9 13 2
49 13 7 1 9 0 13 9 2 9 9 2 16 13 9 2 1 9 2 16 3 13 9 9 2 9 0 0 2 15 9 13 9 7 0 9 2 0 7 9 13 0 9 9 7 9 1 9 0 2
3 3 13 2
6 0 7 9 0 13 2
7 3 7 13 9 0 13 2
25 3 9 1 9 0 0 2 16 15 3 3 7 0 13 2 15 3 15 13 7 9 7 3 9 2
3 7 13 2
7 10 7 9 13 9 9 2
5 15 7 15 13 2
6 9 15 3 9 13 2
6 15 3 13 9 9 2
19 3 3 3 1 0 9 9 13 3 13 2 9 7 0 9 9 9 13 2
24 15 3 16 9 0 3 13 2 3 9 9 13 0 7 3 15 2 9 7 13 1 0 9 2
8 7 15 3 9 0 13 9 2
20 3 7 13 1 9 0 13 0 9 2 16 3 3 15 0 13 0 13 9 2
26 7 3 9 0 1 9 13 0 13 7 9 13 7 3 9 13 9 9 0 0 7 3 9 13 9 2
4 13 3 9 2
6 3 3 3 0 13 2
17 15 3 3 15 15 1 0 9 9 13 9 13 2 7 15 13 2
5 3 3 0 13 2
32 16 7 13 2 13 2 16 1 9 9 13 7 9 0 9 13 15 0 3 2 16 3 15 13 3 13 7 7 15 9 13 2
14 0 7 15 9 1 9 0 0 13 2 0 0 7 2
18 16 15 3 13 7 9 9 13 2 3 3 15 15 13 9 0 13 2
7 0 3 15 1 0 13 2
3 7 13 2
5 15 7 13 9 2
9 15 7 0 13 9 13 9 13 2
11 15 7 3 3 13 13 13 1 0 9 2
27 15 7 16 7 9 7 9 9 9 13 1 9 13 9 9 2 3 15 13 9 9 0 13 0 1 0 2
9 1 7 9 9 13 0 9 0 2
12 13 7 1 9 0 9 2 16 3 3 13 2
8 7 3 0 1 9 9 13 2
12 15 7 3 1 0 13 9 13 1 9 13 2
9 1 7 9 0 0 9 13 9 2
6 15 7 1 15 13 2
11 15 7 9 7 9 7 7 0 9 13 2
8 13 7 15 9 7 13 13 2
6 3 13 13 9 9 2
9 15 3 15 3 3 0 13 9 2
9 15 7 9 9 13 0 9 13 2
4 15 7 13 2
9 3 3 0 15 13 13 9 0 2
12 13 7 3 9 7 9 13 13 13 9 0 2
10 15 7 9 13 9 13 2 16 13 2
15 1 3 13 9 9 7 9 2 16 7 3 3 0 9 2
11 7 9 3 9 3 13 3 9 13 9 2
6 1 3 9 9 13 2
13 3 7 2 16 13 3 2 13 0 3 15 3 2
18 9 7 15 13 15 2 15 0 7 0 13 0 2 0 7 15 13 2
18 16 15 3 13 7 9 9 13 2 3 3 15 15 13 9 0 13 2
7 0 3 15 1 0 13 2
7 15 7 3 13 0 9 2
14 13 3 0 0 0 0 2 13 7 9 0 0 9 2
9 7 3 13 0 13 9 9 0 2
5 13 7 9 9 2
18 7 15 3 9 0 0 9 9 2 15 13 0 9 2 13 1 9 2
11 9 7 13 9 9 16 9 3 0 13 2
10 15 7 0 9 13 2 16 0 13 2
5 9 3 3 13 2
22 7 3 15 13 9 7 0 7 2 16 3 3 9 0 9 9 13 0 1 9 13 2
21 13 7 7 0 13 9 13 15 1 9 7 13 3 9 7 3 13 9 0 13 2
4 7 13 13 2
6 15 7 13 0 9 2
11 3 7 3 13 16 3 9 7 9 13 2
15 9 7 0 3 13 2 16 9 0 13 7 1 9 13 2
20 9 7 3 3 3 13 9 9 0 9 7 9 0 3 1 15 13 9 0 2
15 13 7 9 0 2 15 0 0 0 7 9 7 9 13 2
15 9 7 15 15 13 2 16 3 3 3 13 0 9 13 2
7 3 7 3 7 9 13 2
5 13 7 1 9 2
11 15 3 3 9 1 9 13 0 13 9 2
6 15 7 3 9 13 2
11 15 7 13 9 0 9 13 0 1 9 2
8 13 7 15 3 13 13 13 2
6 15 7 3 13 9 2
9 0 3 3 15 13 9 7 9 2
20 7 15 3 1 9 13 0 9 13 0 9 0 9 13 7 9 1 13 9 2
6 15 7 13 9 0 2
13 7 16 13 7 13 9 2 13 3 13 3 0 2
15 7 0 9 3 13 0 1 3 0 13 9 13 0 9 2
11 0 7 9 1 9 0 13 9 7 0 2
9 0 7 0 9 3 9 13 9 2
8 0 7 0 9 0 13 9 2
13 9 7 3 0 13 13 9 0 2 0 9 13 2
3 7 13 2
19 13 7 9 9 0 2 13 7 1 9 9 0 7 15 13 9 0 13 2
4 7 13 13 2
6 15 7 3 13 9 2
10 3 3 9 0 9 3 13 0 13 2
10 7 15 13 13 9 7 9 9 13 2
5 0 7 13 9 2
24 3 3 3 3 13 0 9 16 3 13 2 3 16 9 9 13 2 16 13 9 0 0 9 2
39 7 16 15 3 13 0 0 9 2 1 9 13 0 9 2 16 9 0 13 9 0 9 1 9 0 1 9 13 1 9 2 16 15 9 9 13 13 9 2
21 13 7 10 3 9 9 3 13 2 13 1 9 1 0 9 2 3 0 9 9 2
12 15 7 3 9 9 0 2 0 2 13 9 2
7 3 7 13 13 0 9 2
21 16 0 13 9 2 13 9 0 0 9 2 9 1 9 13 2 13 7 9 0 2
3 7 13 2
13 13 7 9 9 9 9 2 7 13 9 9 9 2
6 3 7 13 0 9 2
22 10 7 13 9 13 9 0 2 15 3 3 9 0 9 13 3 13 2 0 9 13 2
3 7 13 2
11 13 7 0 9 2 3 7 13 1 9 2
26 7 10 3 15 9 9 13 13 0 3 2 1 15 13 2 16 3 13 9 0 3 1 0 9 0 2
11 9 7 3 1 0 9 13 0 0 9 2
6 3 7 3 0 13 2
6 3 7 0 9 13 2
23 7 9 7 9 9 7 9 0 9 0 7 9 13 9 2 7 1 15 0 9 13 13 2
12 15 7 13 13 2 16 9 9 1 0 9 2
10 13 2 3 13 2 16 13 0 2 2
22 7 3 3 3 13 1 0 9 2 7 1 15 7 9 0 9 2 13 0 13 0 2
30 16 7 13 2 3 3 13 1 9 9 2 13 9 0 9 1 9 2 2 10 7 12 1 15 7 7 2 15 0 2
18 2 13 7 3 15 13 1 9 0 2 7 15 15 13 9 0 9 2
8 15 7 3 9 0 0 13 2
34 16 15 9 13 9 9 0 1 9 0 7 15 9 2 13 1 9 2 16 9 13 13 0 9 7 9 0 2 3 15 13 1 9 2
5 9 7 3 13 2
7 3 7 13 9 0 0 2
11 13 7 13 1 9 1 9 0 3 0 2
6 13 7 3 3 9 2
8 15 3 13 3 0 0 13 2
17 7 3 3 0 9 0 9 13 3 3 15 9 7 9 13 13 2
5 13 7 13 9 2
7 15 7 3 13 9 0 2
8 3 7 3 13 9 9 0 2
9 1 15 15 0 7 9 13 9 2
3 7 13 2
6 7 13 9 9 9 2
9 13 7 3 9 0 9 9 9 2
24 7 3 13 3 0 13 9 9 13 2 9 7 3 0 9 13 9 2 15 7 1 9 13 2
7 3 13 0 1 9 0 2
7 15 7 3 13 9 0 2
6 2 7 3 13 13 2
5 0 7 13 9 2
7 3 7 9 13 0 9 2
3 7 13 2
6 3 7 13 0 9 2
7 3 7 9 13 9 0 2
10 0 7 9 7 7 9 0 9 13 2
8 0 3 3 9 9 13 9 2
8 0 2 15 15 13 0 9 2
18 15 7 0 9 15 7 0 2 3 13 9 13 13 3 1 9 0 2
11 3 7 13 1 9 0 0 7 0 7 2
11 3 0 2 15 15 15 3 13 0 9 2
16 3 7 15 13 3 1 0 9 9 2 15 9 9 0 13 2
9 7 15 7 15 7 15 13 9 2
12 9 3 3 10 0 9 0 13 13 10 9 2
16 10 3 9 0 10 9 13 0 10 1 10 3 9 13 9 2
20 3 3 9 1 9 13 13 9 2 3 16 9 2 7 10 9 0 15 13 2
6 13 3 3 15 9 2
30 0 3 13 9 1 15 9 10 9 2 13 15 2 13 15 1 10 9 1 9 13 9 2 13 3 16 3 13 9 2
35 0 3 3 10 1 10 9 13 9 13 10 9 9 0 13 2 9 7 0 1 9 9 0 13 7 3 13 1 10 9 10 9 9 13 2
21 10 3 9 7 10 13 9 0 13 10 9 2 10 7 9 7 10 0 13 13 2
23 3 3 9 13 13 2 7 1 10 9 9 13 15 13 10 9 10 9 10 1 10 9 2
10 1 3 10 9 3 13 9 3 9 2
22 3 3 9 15 13 13 13 15 1 9 2 7 16 1 10 9 13 10 9 10 9 2
9 15 3 3 9 3 7 9 13 2
13 15 3 10 3 0 13 2 10 0 0 15 13 2
11 15 3 1 15 13 0 2 0 13 0 2
14 10 0 3 13 9 0 1 15 13 2 13 0 3 2
37 9 13 9 3 9 2 9 3 9 2 9 7 9 10 1 9 9 2 15 13 1 9 1 9 3 7 9 13 1 9 9 1 10 9 13 9 2
21 0 10 9 0 0 15 15 13 10 3 13 9 1 9 9 2 10 7 9 13 2
18 13 3 9 3 3 9 7 9 10 1 10 9 2 0 7 13 0 2
10 1 3 10 9 9 0 9 13 0 2
22 10 3 9 9 10 1 10 9 13 9 13 0 3 9 13 10 9 7 1 9 9 2
18 10 3 9 3 13 2 13 9 1 10 9 10 9 2 13 3 9 2
18 13 9 2 10 10 9 9 13 2 9 9 2 0 7 9 10 9 2
21 9 3 3 10 9 10 9 10 9 0 9 9 13 9 2 9 7 10 9 0 2
28 10 3 0 9 13 0 10 9 13 0 9 10 9 2 1 15 10 9 0 13 10 0 0 2 0 9 13 2
20 0 3 3 10 9 13 10 15 9 2 13 7 13 15 13 9 0 0 0 2
36 3 3 15 13 2 13 3 15 10 0 9 10 9 13 3 2 0 10 9 7 10 0 10 9 13 10 9 7 3 3 10 9 10 9 13 2
10 1 3 9 13 13 3 10 9 9 2
12 3 3 10 0 9 13 2 1 15 13 13 2
16 15 3 13 15 13 0 9 0 2 7 15 13 16 13 0 2
21 10 3 3 13 15 13 2 13 16 0 15 1 15 13 0 2 10 7 13 15 2
13 9 3 15 13 3 16 3 13 15 13 1 15 2
15 15 3 15 1 10 9 1 15 13 3 10 13 9 13 2
13 1 3 15 13 13 3 10 9 10 0 1 9 2
7 13 3 1 10 9 9 2
18 1 15 10 9 1 9 0 13 13 2 7 1 9 0 13 15 13 2
27 16 3 1 10 9 13 1 10 9 1 9 7 15 13 2 15 13 10 3 16 3 15 13 13 1 9 2
11 10 3 3 16 3 13 13 2 13 0 2
27 10 3 9 2 16 13 9 10 9 13 2 13 10 9 1 10 9 2 7 1 15 3 13 3 10 9 2
10 13 3 7 13 10 9 13 10 9 2
23 16 3 1 9 13 13 10 9 1 10 9 2 13 13 3 2 7 10 9 13 15 13 2
21 13 3 10 13 1 10 9 3 13 13 7 13 13 2 1 9 13 13 10 9 2
21 1 3 10 9 2 3 3 7 1 10 0 0 3 9 13 0 1 9 0 13 2
9 3 3 3 3 15 13 9 13 2
21 16 3 9 0 13 2 15 9 10 3 13 0 13 15 2 0 13 13 10 9 2
11 10 3 15 13 15 10 13 13 13 13 2
12 13 3 3 3 2 16 10 9 13 2 13 2
11 16 3 10 9 13 2 13 10 9 15 2
35 3 3 9 13 15 3 7 10 9 13 10 9 2 7 0 15 3 3 13 13 2 16 3 3 0 13 9 10 0 13 10 3 15 13 2
21 3 3 15 3 10 15 13 13 13 2 7 15 10 15 0 13 7 13 3 13 2
20 10 3 9 3 3 13 10 13 2 3 7 13 16 15 9 13 13 0 9 2
19 3 3 13 2 7 13 9 3 13 3 10 9 13 7 15 1 15 13 2
4 13 15 13 2
5 13 3 13 15 2
18 16 15 13 9 10 0 13 3 13 2 13 13 0 3 9 13 15 2
26 15 3 13 13 1 10 0 3 9 10 9 13 3 3 3 15 15 13 0 2 13 7 10 9 13 2
33 3 1 15 13 9 13 3 7 13 15 13 3 10 9 7 10 9 9 15 3 9 10 0 1 10 0 9 13 1 9 0 13 2
12 13 3 10 9 7 13 1 10 1 9 9 2
10 13 3 3 10 9 7 13 3 9 2
17 0 10 9 9 3 7 10 9 15 9 0 13 2 16 3 13 2
58 10 3 3 9 3 13 10 9 10 9 13 2 9 7 13 13 9 1 9 3 0 2 7 0 3 9 9 2 13 15 0 1 9 2 1 7 10 9 9 0 13 0 3 7 15 3 9 0 13 13 2 9 10 9 12 0 13 2
13 13 3 15 1 10 9 9 2 9 13 12 9 2
17 0 3 9 13 3 9 10 0 13 10 9 2 7 9 10 9 2
20 0 3 10 9 0 0 15 15 13 1 9 13 9 1 9 10 9 9 9 2
16 13 3 3 3 9 10 0 9 1 15 13 13 2 13 0 2
12 13 7 10 9 0 3 3 10 10 9 9 2
21 13 3 3 9 3 15 16 13 1 3 9 7 1 9 2 7 9 10 9 13 2
34 15 3 9 3 13 1 9 7 13 2 1 15 3 13 9 9 1 9 1 9 10 9 13 13 1 10 9 7 9 1 10 9 13 2
21 9 3 13 9 13 12 9 13 9 10 9 2 7 13 9 0 2 9 7 9 2
13 1 3 3 15 3 16 13 13 2 7 13 3 2
11 0 3 9 13 13 1 10 9 0 15 2
10 13 9 2 13 10 9 1 10 9 2
8 13 3 13 10 9 9 0 2
14 16 3 13 1 10 9 9 0 2 3 13 10 9 2
14 13 3 1 9 3 7 9 7 9 0 3 7 0 2
27 16 3 1 10 9 13 2 9 3 10 1 10 9 3 13 7 13 7 9 13 2 13 7 1 9 13 2
18 10 3 10 3 9 7 10 9 10 1 10 9 16 13 2 13 3 2
15 10 3 9 10 9 13 2 16 9 3 13 9 10 9 2
33 10 3 9 3 13 10 9 15 1 2 16 13 3 13 10 9 13 3 7 13 10 9 2 15 7 15 13 13 15 3 13 13 2
24 10 3 3 12 9 10 12 9 10 9 3 9 13 2 10 3 13 3 1 10 0 10 9 2
10 9 0 3 3 10 10 9 13 13 2
31 10 3 12 10 9 10 13 10 12 9 10 9 13 2 15 13 2 16 3 0 15 13 2 1 10 9 10 9 13 3 2
14 10 3 9 0 9 10 9 0 13 16 3 9 0 2
7 15 3 10 0 13 13 2
14 3 3 3 0 10 9 10 9 10 1 0 9 13 2
15 10 3 0 9 9 13 1 10 9 13 15 0 13 9 2
20 16 13 0 10 9 2 9 13 13 9 0 9 9 2 13 7 10 9 13 2
19 3 10 3 3 9 0 13 2 1 7 10 9 13 1 9 13 10 9 2
28 0 3 15 13 10 9 13 1 9 0 2 3 3 13 15 2 7 3 15 13 13 10 9 13 1 10 9 2
26 10 3 10 9 13 1 9 3 13 13 3 16 10 9 10 0 13 2 15 13 9 10 0 1 9 2
7 9 13 15 3 13 13 2
41 9 3 15 13 15 2 9 10 9 13 9 10 3 9 13 9 1 10 3 2 13 10 9 10 10 9 13 2 13 9 13 2 16 3 15 13 1 10 13 13 2
7 9 3 3 3 13 13 2
27 9 3 2 16 15 15 13 2 3 13 9 1 9 13 9 13 9 3 7 0 9 0 3 10 9 13 2
26 10 3 3 9 1 10 9 13 2 9 7 3 13 0 9 2 7 13 15 9 13 13 2 13 15 2
34 0 13 1 10 9 9 3 15 7 0 2 15 0 13 1 10 9 13 9 2 16 15 13 2 3 13 3 0 7 9 13 1 15 2
5 10 3 3 13 2
32 16 3 3 13 3 15 10 9 7 13 1 9 10 9 10 9 13 1 10 9 2 16 15 13 2 1 15 0 13 10 9 2
35 13 3 10 9 9 3 13 0 1 10 9 7 10 9 13 1 10 0 0 2 13 10 9 13 1 10 9 10 0 9 16 3 15 13 2
38 3 3 10 3 9 15 13 1 15 3 0 15 13 7 0 2 7 12 3 1 9 9 10 9 13 10 9 1 10 9 2 15 7 1 10 9 13 2
13 1 3 10 1 9 3 7 9 9 9 3 13 2
13 9 3 13 9 9 0 10 10 9 10 9 13 2
6 13 3 10 9 9 2
30 0 10 9 13 2 10 0 10 9 13 1 9 13 13 1 9 3 7 9 2 13 7 9 0 13 3 1 9 13 2
6 13 3 13 15 13 2
16 3 10 3 13 1 9 2 10 7 9 13 13 13 1 9 2
18 9 3 10 9 10 1 0 9 13 3 13 2 13 9 12 7 12 2
17 13 3 9 13 10 9 9 10 9 2 9 13 9 12 7 12 2
7 15 3 9 0 13 0 2
22 3 3 10 9 13 1 15 13 10 9 10 9 2 13 1 10 9 9 1 10 9 2
18 13 3 1 10 3 0 9 2 15 3 13 2 7 10 9 9 0 2
39 0 3 3 15 13 10 9 2 3 7 1 9 0 9 3 7 9 2 15 15 0 13 2 15 3 13 0 13 2 0 13 2 10 7 15 3 0 13 2
22 16 3 3 10 1 10 9 9 13 1 9 9 2 10 3 13 9 13 13 10 9 2
40 9 3 15 13 13 0 16 2 16 0 13 15 13 1 15 13 9 2 13 13 9 1 9 2 16 1 10 1 10 9 13 9 13 15 2 15 15 13 13 2
10 3 3 10 10 9 13 9 9 13 2
15 1 3 9 7 9 10 15 0 1 15 13 13 10 9 2
97 13 3 15 2 9 2 9 2 9 2 9 2 9 2 9 2 9 10 9 3 7 9 2 9 2 9 2 9 2 9 2 9 13 7 15 7 13 9 9 2 13 1 9 13 9 0 3 10 0 1 10 9 9 2 15 0 10 9 13 13 2 16 0 15 13 2 7 3 3 9 9 0 2 15 9 9 13 13 13 9 12 1 9 9 13 2 16 3 3 15 10 9 13 13 10 13 2
10 0 3 3 0 3 13 15 13 9 2
14 9 3 0 13 12 9 13 9 10 3 15 9 13 2
24 15 3 3 0 7 10 9 13 10 9 1 1 9 13 1 9 7 3 3 1 9 1 9 2
10 13 3 13 1 10 9 1 10 9 2
25 1 3 9 0 7 0 13 9 10 9 9 13 1 10 9 2 7 13 0 13 0 3 7 0 2
18 13 3 15 10 0 7 13 16 15 1 9 13 2 13 10 9 15 2
14 3 3 13 15 9 13 15 16 15 3 0 13 0 2
9 10 3 13 13 9 0 15 13 2
8 13 3 9 10 13 13 3 2
7 3 3 13 9 13 0 2
26 10 3 13 9 15 3 10 9 3 13 9 13 0 7 0 2 7 15 13 0 9 13 7 0 13 2
18 15 3 10 9 3 13 2 16 10 1 15 2 9 10 9 0 13 2
33 13 3 9 9 1 10 0 1 9 2 13 7 9 13 10 0 13 0 2 7 15 9 0 3 13 3 10 3 13 7 13 3 2
30 16 3 10 1 10 9 13 10 9 10 9 13 0 3 7 0 2 13 15 0 1 15 13 2 13 3 9 3 13 2
8 10 3 13 9 3 7 9 2
17 15 3 13 9 9 9 3 13 13 2 7 1 15 9 9 15 2
14 0 3 0 3 13 2 7 3 3 13 0 10 9 2
29 13 9 10 9 10 9 13 3 10 9 15 9 13 1 10 0 2 10 7 15 9 1 10 9 3 13 1 9 2
24 13 3 10 9 10 9 13 0 1 10 9 13 10 9 2 1 10 9 7 15 13 10 9 2
11 9 3 12 7 12 13 13 1 10 0 2
30 15 3 15 13 7 13 1 10 9 9 10 9 0 13 2 13 7 1 15 10 9 16 0 13 9 13 3 16 13 2
21 9 3 3 13 13 10 9 10 9 2 10 7 9 10 9 15 2 0 9 13 2
39 10 3 9 0 13 10 3 9 7 10 9 2 13 0 10 9 13 9 3 7 9 10 15 9 2 15 15 13 3 2 10 9 13 15 9 13 0 13 2
26 1 0 3 10 9 16 13 3 7 13 2 13 1 0 10 0 10 9 3 13 7 1 9 0 13 2
12 9 3 0 9 13 13 1 9 3 0 13 2
19 1 3 10 0 9 0 3 13 13 15 3 15 13 2 0 7 3 13 2
10 1 3 12 9 9 10 9 9 13 2
17 15 13 9 12 13 9 0 3 0 7 0 2 0 9 3 13 2
42 16 3 3 13 0 10 9 9 0 13 2 16 3 10 9 13 13 1 10 13 2 9 3 1 10 12 9 10 0 13 12 12 2 9 7 1 10 9 0 0 12 2
32 0 10 0 9 10 1 10 12 9 2 13 12 3 0 3 0 7 0 2 10 0 0 10 0 9 10 3 15 0 13 9 2
13 15 3 15 3 13 0 13 7 9 0 13 9 2
18 15 3 10 13 15 2 3 15 15 13 2 16 13 3 10 9 13 2
27 3 3 15 10 0 0 3 10 1 9 13 0 13 2 16 3 15 9 13 0 0 13 3 13 10 9 2
15 0 3 3 0 9 0 13 2 0 7 3 13 9 0 2
21 10 3 3 0 0 0 3 0 13 10 0 0 2 15 7 10 0 7 0 0 2
17 10 3 9 13 7 9 0 13 13 0 2 10 7 15 13 15 2
30 9 3 7 9 3 3 0 15 13 2 15 3 10 9 15 13 2 0 7 13 2 0 2 0 9 2 9 2 0 2
27 10 0 3 3 15 13 9 13 0 13 2 16 9 0 13 0 0 13 2 7 15 3 13 0 7 13 2
10 15 3 3 10 0 13 2 15 0 2
10 3 3 3 9 9 0 0 0 13 2
10 10 3 3 13 2 15 7 0 13 2
10 0 3 3 13 9 10 9 0 13 2
33 15 13 10 9 3 3 3 13 2 7 9 15 13 0 13 2 3 13 0 13 2 15 10 13 0 13 10 9 0 9 13 13 2
22 1 3 9 13 13 1 9 9 0 9 2 16 13 2 16 13 15 13 9 0 0 2
20 3 3 15 13 13 9 2 15 15 10 9 13 10 13 13 0 1 10 9 2
6 9 3 10 13 9 2
31 10 3 16 13 7 15 9 13 2 13 10 9 13 3 10 9 9 2 13 7 13 15 10 9 3 3 1 0 9 13 2
31 9 3 3 9 7 10 15 0 15 13 1 9 9 2 1 10 9 13 1 10 9 13 2 16 15 15 13 10 9 13 2
32 13 3 15 1 9 10 9 10 9 2 13 1 10 9 9 9 13 7 3 0 9 2 13 9 3 9 2 9 7 10 0 2
20 13 3 15 1 10 9 9 1 9 10 0 0 13 13 2 9 7 15 13 2
11 13 3 0 10 9 10 9 7 10 9 2
18 16 3 10 13 13 10 9 2 13 3 3 7 15 13 2 13 15 2
7 15 3 9 7 9 13 2
6 9 3 15 13 15 2
28 9 3 0 13 0 13 7 13 1 0 2 3 13 9 0 13 1 0 2 9 7 0 3 0 13 13 0 2
8 10 3 3 9 13 1 9 2
15 1 3 10 0 9 0 1 10 0 9 9 9 13 0 2
13 13 3 15 1 10 9 0 10 10 9 9 13 2
17 3 3 10 9 1 15 13 13 3 0 15 2 13 7 1 15 2
12 9 3 13 1 10 9 10 9 9 13 15 2
6 15 13 13 3 13 2
22 3 3 13 15 10 9 3 0 9 7 9 13 15 2 16 3 15 13 1 10 9 2
17 10 3 3 15 13 2 9 7 13 10 9 10 9 13 15 0 2
9 9 3 1 10 0 3 13 3 2
6 3 3 3 15 13 2
10 0 3 3 13 7 15 10 3 13 2
24 9 3 9 7 10 9 0 13 2 7 13 10 13 13 3 0 13 15 10 9 1 10 9 2
3 15 13 2
17 13 3 15 10 9 2 13 10 10 9 9 13 10 13 10 9 2
18 3 13 3 10 9 10 3 9 15 13 2 13 1 15 10 9 15 2
30 3 3 0 15 15 13 13 2 3 0 9 15 13 7 9 3 7 0 15 13 9 1 3 9 7 1 9 13 13 2
7 0 3 15 13 9 13 2
21 15 3 15 3 13 13 1 10 9 2 7 9 13 16 15 0 13 15 3 13 2
4 13 9 15 2
31 1 3 10 9 0 10 3 9 15 0 13 7 1 10 13 3 13 2 9 13 2 16 3 13 1 10 0 15 9 13 2
8 9 3 15 0 13 13 9 2
12 10 3 3 0 13 10 9 3 13 15 13 2
5 13 10 9 15 2
16 10 3 3 13 7 13 15 10 9 2 15 15 0 13 13 2
11 13 3 10 9 1 9 0 13 15 13 2
15 9 3 0 3 13 9 2 0 7 9 0 10 15 13 2
25 16 3 3 1 9 3 13 13 15 2 7 0 15 10 15 15 13 2 13 3 15 13 15 13 2
13 16 3 3 1 9 15 13 10 9 2 13 15 2
15 3 3 13 1 15 13 2 13 7 15 13 1 10 9 2
16 13 3 15 10 9 13 10 9 9 2 13 7 15 13 15 2
24 3 3 9 0 13 13 13 1 9 3 13 13 2 3 10 13 3 2 3 7 3 13 15 2
16 15 16 15 13 9 2 13 1 15 13 0 3 9 7 9 2
19 13 3 1 10 9 10 9 13 10 9 2 13 7 7 13 15 9 13 2
29 3 3 10 9 2 0 3 10 13 10 9 2 13 7 9 2 13 10 9 10 3 13 2 13 7 10 9 9 2
37 10 3 3 13 10 9 13 10 9 10 9 2 13 7 15 13 10 9 10 13 2 13 7 1 10 9 10 3 9 7 10 10 9 9 13 15 2
19 10 3 9 10 9 10 9 13 3 15 13 16 15 13 10 15 9 13 2
57 13 3 10 9 3 13 3 9 0 13 15 1 10 9 13 13 13 7 0 3 7 0 2 10 0 0 13 9 2 10 3 0 13 2 16 3 9 13 10 0 9 10 9 13 13 2 10 7 0 2 16 9 13 15 13 0 2
17 13 3 1 15 10 9 13 10 0 2 3 7 13 15 10 9 2
40 13 3 15 1 10 9 13 15 9 13 10 9 2 13 15 13 10 0 2 13 10 3 0 15 9 2 7 16 1 15 10 13 13 13 2 3 15 13 0 2
30 13 3 3 15 15 0 10 0 0 2 16 3 0 0 13 2 7 9 3 15 2 15 15 3 3 13 10 13 13 2
11 9 3 3 13 16 13 13 10 15 9 2
43 9 3 10 9 10 9 2 0 3 10 9 3 10 0 9 13 9 7 10 13 2 16 9 10 9 13 1 10 9 2 13 9 13 15 15 13 0 2 13 10 9 15 2
13 9 3 1 12 9 1 9 0 13 10 9 13 2
44 3 3 10 9 10 9 9 13 1 9 10 9 7 10 10 9 9 13 9 3 9 13 2 13 7 1 9 2 16 3 13 2 16 0 13 10 9 2 13 15 13 10 9 2
18 10 3 15 13 1 3 9 7 1 9 2 10 7 10 0 1 9 2
8 9 3 1 9 13 15 13 2
26 13 3 13 10 9 15 0 13 2 16 16 13 10 9 13 2 13 15 0 13 16 13 1 9 13 2
15 15 0 3 3 10 0 10 9 13 2 3 13 1 0 2
27 1 3 9 16 13 0 1 10 9 10 9 13 10 9 7 13 10 13 2 10 9 1 0 9 13 15 2
19 13 3 15 9 3 9 7 9 9 2 3 0 13 2 7 3 13 13 2
23 9 15 1 9 13 0 9 13 1 9 1 0 9 2 15 9 3 13 2 9 7 13 2
13 15 10 9 13 10 0 13 13 13 1 10 9 2
20 16 3 3 15 10 13 13 13 10 9 2 3 10 9 0 13 13 10 9 2
29 10 3 16 10 1 9 13 2 3 13 3 7 13 2 13 0 13 9 10 1 9 2 16 15 13 15 15 13 2
18 16 3 3 13 1 10 9 10 0 2 13 10 0 10 9 13 15 2
24 13 10 13 0 13 3 7 13 2 9 7 9 13 3 13 15 1 9 0 2 0 9 13 2
10 10 3 3 1 9 3 10 9 13 2
11 1 3 15 9 0 10 1 9 9 13 2
37 9 3 3 10 0 0 0 13 2 9 3 0 7 0 7 9 0 7 9 0 7 9 2 13 9 0 2 13 2 13 10 9 3 15 15 13 2
14 9 3 0 13 13 0 0 15 15 15 0 13 0 2
32 16 3 1 10 9 13 2 13 9 0 9 1 15 13 2 1 3 10 0 13 0 2 1 3 10 0 0 2 9 7 0 2
12 13 3 3 9 9 9 0 13 9 9 12 2
6 13 3 15 0 9 2
6 13 3 1 9 9 2
14 13 3 15 9 9 10 0 9 13 2 7 15 13 2
9 3 3 10 13 13 15 9 13 2
37 3 9 3 0 9 13 2 15 1 10 9 9 13 2 7 9 12 13 2 0 3 7 0 2 15 10 0 13 9 13 13 9 2 3 3 13 2
22 13 3 3 15 9 2 13 7 10 15 9 9 13 13 2 15 13 10 9 3 13 2
23 3 10 3 9 2 1 15 10 9 13 10 9 2 9 13 2 3 7 10 3 9 0 2
35 0 3 9 3 0 0 13 1 15 10 9 2 3 9 0 0 2 7 3 3 9 9 0 0 2 15 9 10 9 10 9 9 13 13 2
17 3 3 3 10 15 9 10 1 10 9 13 10 9 7 10 9 2
39 15 3 1 9 13 2 10 7 9 2 13 15 10 3 9 7 10 9 2 13 9 3 0 0 3 7 9 0 0 0 2 10 9 10 9 13 3 0 2
19 10 3 3 0 1 15 13 13 1 9 7 9 1 10 9 10 0 9 2
88 10 3 13 13 10 9 0 10 9 1 10 0 13 10 9 13 10 0 16 13 1 9 9 7 16 0 9 9 13 0 2 16 7 13 1 10 13 10 9 13 10 9 2 13 10 9 13 9 10 9 3 7 0 9 9 2 13 0 9 13 0 1 9 2 15 3 0 9 13 10 9 2 7 3 15 13 16 13 1 9 7 16 0 9 9 13 0 2
28 10 3 15 13 2 10 7 9 0 1 15 10 9 13 2 13 9 2 16 13 1 9 2 0 9 15 13 2
10 10 3 9 0 13 10 13 0 13 2
41 16 3 13 10 9 13 10 9 2 13 3 10 9 2 3 7 13 13 10 9 9 2 13 3 1 9 9 13 2 13 15 10 9 2 1 9 12 9 0 9 2
26 9 3 1 15 13 9 7 9 9 3 0 7 9 2 7 13 10 13 15 13 9 1 10 3 9 2
10 13 3 10 9 10 9 13 10 0 2
11 16 3 3 13 10 9 9 2 13 15 2
7 10 3 9 15 13 15 2
32 0 13 10 9 10 9 0 15 3 0 13 2 13 9 0 1 9 13 9 2 3 3 15 7 10 1 15 13 3 10 9 2
30 1 3 15 13 13 15 3 9 0 13 13 9 2 13 7 13 0 7 9 13 10 3 10 0 9 10 7 10 0 2
17 15 3 13 10 13 2 13 10 0 10 3 0 10 7 0 9 2
12 3 10 3 3 3 13 2 10 7 0 9 2
29 1 3 3 9 9 13 9 10 9 2 1 7 9 10 9 10 1 10 9 3 7 10 9 9 2 13 3 9 2
15 1 3 10 9 16 13 1 9 2 13 1 9 0 13 2
18 3 3 3 1 10 9 13 7 1 10 9 3 1 9 13 9 13 2
12 0 3 9 13 10 9 2 3 13 3 13 2
13 16 15 13 13 13 2 13 10 9 0 9 13 2
25 16 3 13 3 0 15 10 0 2 10 0 9 13 0 1 10 9 10 1 9 3 10 9 13 2
18 13 3 16 10 13 9 9 13 1 0 10 9 2 15 13 1 9 2
18 10 3 0 9 3 16 13 3 3 10 0 13 2 16 15 13 13 2
30 13 3 1 10 0 13 0 2 1 0 15 10 9 13 13 1 9 10 9 2 9 3 13 15 7 0 9 0 0 2
17 3 3 3 15 13 3 10 0 9 2 13 0 2 0 3 13 2
25 0 3 3 10 9 10 3 0 13 3 7 13 13 10 9 1 9 10 9 0 10 9 13 9 2
12 9 3 13 9 7 13 10 0 9 13 0 2
21 13 3 15 10 0 10 9 13 7 9 3 13 0 7 9 1 9 13 7 13 2
42 9 3 10 0 13 7 13 10 9 13 9 0 3 9 3 13 0 1 10 9 2 16 7 13 13 2 0 10 9 13 2 7 16 0 15 13 13 9 2 15 13 2
12 13 3 9 7 10 9 10 0 13 13 15 2
53 13 15 3 7 9 13 1 10 9 10 9 3 13 10 0 2 10 15 13 1 9 13 13 3 2 13 7 10 9 9 0 1 15 13 2 0 13 1 10 1 9 13 9 2 9 3 13 7 0 13 0 9 2
24 10 3 9 10 10 9 13 13 15 10 9 13 9 0 15 0 3 3 13 9 2 0 7 2
8 9 3 9 13 13 15 3 2
19 1 3 3 0 9 15 13 10 3 10 9 9 7 10 10 9 13 15 2
17 3 3 9 13 10 0 9 2 7 10 9 3 9 13 13 13 2
11 10 3 13 9 3 1 9 1 15 13 2
20 13 3 10 9 10 9 13 9 2 16 13 15 10 9 13 9 1 10 9 2
59 13 3 10 9 7 13 1 15 9 2 13 3 1 10 9 9 0 2 16 15 13 2 0 2 16 3 13 1 0 10 0 9 10 0 13 3 0 7 9 0 13 3 2 16 3 3 3 15 1 9 10 0 13 13 9 9 13 15 2
23 1 10 9 10 9 13 9 15 9 13 9 2 9 1 9 9 13 0 9 3 3 0 2
28 0 10 9 13 9 2 1 9 13 7 13 9 0 0 13 0 13 13 2 13 1 10 9 2 0 9 13 2
12 10 10 13 13 13 1 10 9 2 13 15 2
7 10 3 3 15 13 13 2
33 3 3 1 3 10 9 9 13 16 9 9 13 2 7 10 1 10 9 13 10 9 13 0 10 9 13 3 10 9 7 13 9 2
22 13 3 10 9 9 10 13 10 9 1 10 9 10 1 9 13 13 10 9 10 9 2
29 0 3 9 3 15 13 9 7 13 0 13 10 9 2 3 13 15 13 1 10 0 9 9 13 15 3 1 9 2
10 9 3 16 13 13 10 9 10 9 2
24 13 3 10 9 10 13 1 15 13 1 10 9 10 3 2 13 7 1 9 13 1 10 9 2
21 9 3 9 13 13 3 10 9 2 3 13 9 1 10 9 15 15 13 3 15 2
13 0 3 0 13 9 2 9 13 10 9 10 9 2
18 3 3 2 3 0 9 13 2 9 13 7 0 15 13 1 10 9 2
30 3 3 0 0 13 1 9 2 7 0 15 9 13 9 2 15 9 13 9 2 9 0 13 2 13 3 9 7 9 2
17 1 9 3 13 1 0 9 13 3 2 7 0 10 9 13 9 2
29 1 3 0 10 9 15 13 10 3 1 10 9 9 13 15 7 1 10 9 13 2 15 10 9 1 9 13 0 2
29 15 3 3 13 2 9 7 10 1 10 9 2 16 3 9 10 9 13 2 7 3 16 13 9 2 9 0 13 2
18 16 3 13 1 10 9 15 13 1 10 9 2 3 3 13 1 15 2
37 3 15 3 9 13 1 10 13 7 10 1 9 2 16 13 1 9 13 1 10 9 2 1 15 13 13 1 9 9 0 2 7 0 13 10 9 2
22 3 0 9 13 13 9 9 10 9 0 9 2 15 10 13 13 1 0 9 15 13 2
17 13 3 10 9 2 10 3 9 13 2 9 7 13 9 1 9 2
22 10 3 3 15 13 13 15 2 9 7 13 10 0 7 13 13 10 13 13 10 9 2
9 10 3 1 9 13 10 9 13 2
19 13 3 15 9 3 0 9 13 2 16 3 13 3 10 9 13 7 13 2
28 13 10 9 1 9 13 2 10 7 13 10 13 13 10 13 1 9 2 13 3 13 7 13 0 1 10 15 2
22 1 0 9 10 9 13 2 1 0 10 9 0 13 10 9 13 1 0 9 10 9 2
25 3 9 3 13 9 2 9 7 10 3 1 10 9 13 2 10 7 15 1 9 13 1 10 0 2
29 10 3 3 9 15 10 9 0 13 10 9 13 2 10 7 9 1 0 3 0 13 7 13 3 10 9 0 9 2
19 1 3 9 13 7 9 1 9 10 0 9 13 10 9 1 9 0 13 2
19 10 3 3 0 15 3 0 13 3 0 9 1 3 15 0 7 9 0 2
6 13 3 3 1 9 2
24 9 10 9 0 9 13 1 9 1 10 9 2 16 13 1 10 9 2 3 10 9 13 15 2
8 13 3 15 9 13 7 9 2
18 10 3 3 15 1 15 13 3 13 15 10 0 10 3 13 9 9 2
22 3 3 0 9 13 2 9 13 9 2 9 3 15 13 7 9 2 1 9 13 15 2
16 16 3 13 0 2 13 10 0 0 2 7 13 15 3 13 2
23 1 3 10 1 9 13 2 9 3 9 7 9 2 1 3 15 10 9 7 9 13 9 2
14 3 3 13 13 2 10 7 9 13 0 13 13 3 2
41 0 3 1 3 9 0 7 0 3 0 9 2 3 3 13 3 7 13 2 7 3 15 3 13 9 13 2 7 13 9 0 13 13 1 9 1 0 10 9 9 2
7 10 3 9 15 13 15 2
4 9 15 13 2
4 0 15 13 2
4 3 15 13 2
11 0 1 9 0 9 13 2 10 15 13 2
6 15 3 15 3 13 2
11 13 15 9 0 13 7 0 9 9 13 2
31 15 16 13 13 10 9 2 9 3 10 0 13 2 10 7 9 13 1 9 13 2 9 0 0 2 3 3 13 10 9 2
24 13 3 10 9 2 0 15 13 2 9 3 13 15 13 15 7 9 13 10 9 10 9 13 2
23 10 3 9 0 1 15 13 3 7 1 15 13 0 1 9 1 10 9 10 9 9 13 2
41 1 3 3 10 0 9 3 3 3 13 1 10 9 2 1 7 10 1 9 9 7 10 9 3 7 9 9 1 9 3 10 9 0 10 9 13 2 9 0 13 2
23 16 3 10 9 13 1 9 2 13 0 1 9 13 15 3 9 13 3 10 9 9 13 2
12 10 3 9 15 13 10 9 10 9 9 13 2
24 16 3 13 3 0 3 13 10 9 10 9 13 3 10 1 9 13 10 9 1 15 13 9 2
10 13 3 15 10 0 13 10 9 15 2
13 3 9 13 0 9 2 15 15 13 9 9 13 2
22 10 13 0 10 9 2 10 3 13 1 10 9 2 9 10 0 13 3 13 15 15 2
14 0 3 10 9 9 13 1 9 3 9 13 7 9 2
25 13 3 0 10 9 9 1 10 9 2 13 1 0 13 9 13 2 7 1 9 13 13 10 13 2
15 15 3 1 0 13 10 9 9 13 2 13 13 9 0 2
23 1 3 9 3 3 13 0 0 9 10 3 13 15 7 13 10 0 9 0 13 10 9 2
5 13 3 13 3 2
26 10 3 3 15 13 15 3 13 2 10 7 13 10 13 13 10 9 1 10 9 15 13 2 3 13 2
45 10 9 12 13 9 10 9 13 13 2 10 3 9 7 10 9 10 3 9 7 10 0 2 10 7 13 9 10 9 1 9 13 2 1 15 0 13 2 16 1 0 9 9 13 2
13 13 3 15 7 13 1 9 13 9 0 10 9 2
10 10 3 1 9 0 13 15 9 13 2
20 10 3 13 1 9 7 13 10 15 9 1 10 9 13 1 3 13 10 9 2
20 9 3 16 13 2 13 2 13 7 10 9 7 10 9 13 13 13 1 9 2
18 3 1 0 10 9 2 16 13 15 2 0 0 10 9 13 10 9 2
11 3 3 15 3 10 0 10 9 13 13 2
24 15 3 3 0 13 10 9 13 1 9 9 9 3 13 7 13 9 2 13 3 15 13 13 2
18 10 3 13 13 13 15 9 10 9 3 7 0 9 9 2 13 15 2
32 9 3 3 15 1 9 13 2 9 7 13 3 15 10 9 10 9 13 13 3 10 9 10 9 7 13 9 9 1 7 9 2
23 13 3 10 9 1 9 9 13 2 1 9 13 13 0 15 3 10 9 1 9 13 9 2
7 9 3 15 13 13 9 2
20 15 3 3 1 10 9 10 9 13 2 7 16 1 0 15 13 9 13 0 2
32 3 15 3 15 13 0 13 2 15 7 13 9 0 9 3 3 13 1 10 9 7 9 0 9 13 13 2 9 13 13 9 2
13 0 10 9 3 13 1 9 1 9 0 13 0 2
25 10 3 9 13 16 16 13 1 10 9 10 9 13 1 10 9 2 13 9 13 15 9 0 13 2
38 0 3 9 13 16 16 13 10 13 10 9 10 9 2 13 7 9 3 7 9 13 2 13 10 9 1 9 2 9 3 9 13 13 15 1 10 9 2
15 3 3 3 3 10 13 13 13 1 9 16 13 1 9 2
8 1 3 3 10 9 3 13 2
19 9 3 13 10 9 13 9 1 9 2 13 13 9 3 7 10 9 9 2
33 13 3 9 13 1 9 2 10 15 9 13 3 3 13 0 2 1 7 0 10 9 3 10 3 9 1 9 13 2 13 9 15 2
5 9 15 13 9 2
19 1 3 3 9 13 7 13 2 3 9 7 13 13 2 3 15 0 0 2
17 15 3 3 2 16 13 2 15 15 13 2 15 3 3 13 15 2
10 13 3 10 0 0 13 7 0 13 2
17 15 3 3 9 13 9 2 15 3 1 9 13 9 13 1 9 2
7 15 13 3 13 10 9 2
14 9 3 2 16 9 13 2 13 3 0 7 0 15 2
8 10 3 9 1 9 9 13 2
18 13 3 10 9 0 10 3 0 16 9 13 9 0 2 3 7 9 2
38 10 3 9 13 10 3 0 9 7 10 0 10 9 9 2 15 13 1 0 9 1 9 2 3 7 9 3 1 0 13 13 2 1 7 10 0 9 2
20 13 3 15 7 13 3 1 9 9 3 3 0 9 13 2 1 0 7 9 2
21 3 10 9 9 13 3 0 10 9 10 3 1 9 10 3 9 1 10 9 9 2
9 13 3 9 15 10 9 0 0 2
8 9 9 0 9 12 9 13 2
24 9 3 10 9 2 13 9 3 9 9 7 9 2 9 10 9 13 13 2 13 9 9 3 2
12 9 10 9 9 9 13 13 1 9 10 0 2
20 3 3 1 0 13 15 2 9 15 13 10 9 3 13 7 10 9 10 9 2
23 9 3 13 2 3 3 13 10 9 1 9 7 3 15 13 2 3 3 13 13 15 15 2
51 10 3 15 1 9 13 2 16 0 0 15 13 2 13 10 1 15 13 9 9 13 2 13 7 15 16 13 3 10 9 13 2 9 13 13 16 9 3 2 13 7 10 0 13 1 9 10 9 1 9 2
4 15 3 13 2
21 3 3 9 7 10 13 9 10 9 0 13 2 7 10 9 15 13 9 9 13 2
23 13 3 15 1 0 10 9 10 0 9 9 13 13 16 10 9 13 10 9 3 9 13 2
26 10 3 9 0 10 9 9 10 0 10 9 13 13 2 9 13 9 0 1 15 3 3 13 10 9 2
14 15 15 3 10 9 10 13 13 13 7 9 9 13 2
12 9 3 13 13 10 9 9 9 10 9 9 2
10 1 3 9 0 9 0 3 13 13 2
28 9 3 13 0 10 9 15 3 3 9 2 7 1 15 2 16 10 9 13 1 10 9 2 10 9 13 15 2
21 0 3 3 10 9 9 13 15 9 13 13 1 9 15 15 1 10 3 9 13 2
35 10 9 13 10 9 1 3 10 9 13 16 13 1 9 2 7 3 3 13 9 0 2 13 1 15 10 9 13 2 13 1 10 9 9 2
24 3 16 3 13 0 10 9 2 0 0 13 2 10 3 7 10 3 13 3 10 0 9 13 2
6 3 15 3 3 13 2
7 3 3 3 13 13 15 2
25 3 13 3 10 9 10 9 7 13 2 13 7 10 9 15 0 2 0 7 15 13 0 0 13 2
15 9 3 13 10 15 9 7 13 10 3 13 0 13 9 2
18 16 3 13 13 10 9 2 13 9 1 10 9 13 15 1 9 13 2
6 9 3 3 3 13 2
19 9 3 16 13 7 13 9 2 3 1 10 9 9 13 1 10 0 15 2
16 9 3 0 13 7 13 0 0 2 9 0 13 13 9 13 2
25 3 10 3 15 13 2 16 13 1 10 9 2 13 9 1 10 9 13 1 0 9 13 1 9 2
29 10 3 13 7 13 9 9 2 15 13 15 0 2 0 13 13 0 13 16 3 3 13 3 3 9 13 1 9 2
9 15 13 9 10 9 0 9 13 2
12 13 3 15 10 9 13 10 9 13 13 13 2
12 13 3 15 9 2 16 3 13 13 9 13 2
9 3 3 13 0 1 10 9 9 2
13 3 3 16 3 15 13 1 10 9 13 10 9 2
21 9 3 3 15 13 9 3 13 2 15 3 13 10 13 1 9 3 7 0 9 2
46 9 3 3 13 9 1 10 9 10 13 1 10 9 2 13 16 13 13 9 13 10 9 2 13 13 9 15 13 13 16 13 0 1 10 9 2 3 16 10 0 13 10 9 10 9 2
11 16 3 15 15 13 2 3 13 1 9 2
12 13 3 10 9 1 10 9 15 9 9 13 2
26 3 9 1 9 0 13 2 16 15 1 9 13 10 9 16 16 15 13 2 3 10 9 13 1 9 2
17 13 3 0 10 9 9 0 1 10 9 3 0 7 0 10 9 2
19 10 3 9 15 13 1 9 2 9 7 13 0 2 7 15 13 13 0 2
58 0 10 9 10 15 13 0 3 7 0 9 2 15 0 13 7 13 10 9 9 1 15 13 9 9 13 2 13 3 15 13 10 0 9 13 1 10 9 9 2 10 3 9 13 10 0 9 13 2 3 7 10 0 13 10 0 9 2
30 16 3 10 0 13 2 13 10 3 0 9 3 13 13 0 10 3 13 2 9 7 0 3 13 2 3 16 13 13 2
14 15 3 13 2 10 7 9 13 0 10 9 15 1 2
17 9 9 13 2 7 3 13 3 10 9 15 13 7 10 9 13 2
24 0 3 3 15 1 13 2 7 10 9 0 13 10 0 2 10 3 15 3 13 13 10 9 2
30 16 3 3 13 1 10 9 2 3 16 13 0 10 9 10 9 7 13 15 2 3 13 2 13 7 10 9 10 9 2
25 3 3 10 3 9 10 3 0 13 2 7 16 13 10 13 2 13 1 10 9 0 10 9 13 2
6 10 3 3 13 9 2
20 9 3 13 15 9 1 0 13 10 9 13 1 10 9 0 9 1 10 9 2
24 10 3 3 0 13 1 0 9 13 13 1 9 2 15 7 13 10 0 13 13 3 13 9 2
14 1 3 3 3 10 0 13 9 7 3 3 1 9 2
21 10 3 3 0 10 9 1 0 0 10 9 13 9 13 1 9 1 9 13 9 2
13 10 3 9 15 13 10 9 9 13 13 10 9 2
27 13 3 9 10 0 13 2 3 13 1 9 13 16 0 0 13 2 0 7 3 13 2 15 13 10 9 2
10 13 15 13 2 0 7 0 13 13 2
6 13 3 15 9 13 2
36 10 3 3 0 10 9 3 13 13 1 10 9 2 10 7 10 9 9 13 10 9 0 7 13 10 9 1 10 15 9 1 10 9 13 15 2
7 9 3 0 13 13 0 2
16 9 3 1 10 9 13 13 2 13 7 3 0 0 13 9 2
8 9 3 10 0 15 13 9 2
27 10 3 9 13 10 13 10 0 9 2 13 13 1 9 10 15 9 13 2 3 15 1 10 9 13 0 2
15 0 3 10 9 13 9 13 10 0 9 13 9 13 13 2
12 10 3 3 2 16 13 10 9 2 13 13 2
23 3 15 3 13 7 9 13 0 13 0 9 2 16 13 10 9 10 9 7 13 9 13 2
9 3 3 15 3 9 13 0 13 2
5 9 3 13 3 2
23 16 0 13 9 13 9 2 9 10 9 10 15 13 9 13 10 0 13 10 9 9 13 2
33 1 3 15 13 10 9 16 3 13 2 3 10 15 13 9 9 13 13 2 15 9 13 9 2 1 15 10 9 15 0 13 9 2
10 3 3 13 0 1 15 16 13 3 2
10 0 3 3 13 3 10 9 7 0 2
30 10 3 9 10 0 9 9 0 3 13 10 9 15 15 10 9 13 2 9 13 16 13 10 9 10 9 13 9 0 2
26 10 3 9 1 10 0 9 13 2 10 13 0 10 9 10 9 2 13 15 3 13 0 3 7 0 2
31 10 3 3 9 0 10 9 13 10 0 10 15 9 1 15 10 9 13 1 9 3 13 7 13 2 13 7 1 9 13 2
13 3 3 3 15 3 13 7 1 15 15 9 13 2
14 13 3 0 3 3 9 3 13 7 0 10 9 13 2
7 1 0 3 9 15 13 2
17 13 15 9 2 15 3 0 13 2 10 3 15 0 2 0 7 2
27 1 10 3 13 9 10 9 10 0 1 15 13 2 15 3 13 2 7 3 3 1 9 1 15 13 13 2
7 10 3 9 15 13 15 2
7 13 3 1 9 0 0 2
33 13 3 10 9 2 13 3 10 15 9 13 9 3 13 2 9 3 3 13 13 1 10 13 9 13 2 7 15 15 13 13 13 2
18 15 3 3 15 0 13 2 1 7 15 3 13 10 0 9 10 9 2
31 10 3 9 10 3 3 9 13 7 0 9 13 2 13 9 0 7 0 9 13 2 1 10 9 7 13 10 15 0 9 2
9 13 3 15 10 9 13 1 9 2
11 16 3 15 0 13 2 3 13 10 13 2
60 13 3 15 7 9 13 2 13 3 16 13 3 10 9 13 0 2 7 13 0 10 15 9 13 0 3 13 2 16 7 15 0 13 10 3 15 13 2 15 0 3 1 15 13 16 3 1 0 10 0 7 3 10 1 15 0 0 13 13 2
46 3 13 1 9 9 13 10 9 9 2 16 13 0 3 9 13 10 9 2 13 7 3 13 2 13 10 9 13 2 16 15 15 13 1 15 13 2 13 7 13 15 1 10 13 0 2
11 15 3 3 0 13 15 9 1 9 13 2
18 1 3 3 10 10 9 10 9 13 2 1 7 10 10 9 10 9 2
9 3 15 9 3 0 13 3 13 2
32 10 3 15 13 2 9 7 15 13 13 3 3 15 7 3 1 0 9 13 2 13 7 13 3 15 7 10 1 15 13 0 2
7 10 3 9 13 0 13 2
10 9 3 15 13 13 13 15 0 13 2
15 10 3 15 13 13 0 10 0 9 0 15 0 9 13 2
14 10 3 13 9 3 10 0 13 7 9 10 0 13 2
7 15 3 15 3 15 3 2
8 3 13 3 7 13 10 0 2
8 9 3 0 13 15 9 13 2
15 13 3 10 15 2 13 9 15 0 15 13 1 10 13 2
20 10 3 13 16 15 9 13 0 15 2 13 2 16 15 13 0 2 13 15 2
7 9 9 13 9 13 0 2
12 3 3 13 3 2 16 15 13 15 15 13 2
25 13 10 0 1 0 10 9 9 2 10 13 1 10 13 10 9 13 16 15 3 13 13 10 9 2
20 3 15 3 15 3 13 9 13 10 9 2 7 15 13 13 15 0 0 13 2
12 15 13 10 9 13 2 16 15 13 3 13 2
18 13 3 0 2 7 13 10 0 15 9 13 13 2 13 1 9 15 2
10 9 3 13 15 0 15 15 13 13 2
27 9 3 15 13 0 10 15 9 3 10 9 10 9 3 3 10 9 2 7 16 13 10 9 13 1 9 2
13 13 3 15 13 3 13 13 15 10 9 15 13 2
50 16 3 15 13 10 9 2 13 10 9 1 9 13 13 10 9 1 10 9 10 9 13 16 3 15 13 10 9 13 9 13 1 9 3 13 10 9 9 2 1 15 15 9 15 13 2 13 10 9 2
14 13 3 10 9 7 13 10 13 10 9 13 13 15 2
9 10 13 9 0 13 13 3 9 2
27 9 3 0 9 9 13 2 15 13 0 9 2 9 0 13 13 10 9 7 13 10 15 9 15 15 13 2
27 13 3 9 16 3 1 10 9 10 9 13 10 9 9 7 3 1 0 9 2 3 0 3 13 13 9 2
11 0 3 13 15 2 13 3 7 13 15 2
7 0 3 15 13 15 13 2
11 1 3 10 9 10 13 3 3 9 13 2
15 13 3 15 9 2 16 13 1 9 2 0 9 15 13 2
19 10 3 1 15 13 3 13 13 13 13 0 10 15 7 10 9 13 9 2
11 3 13 3 10 13 7 13 15 0 13 2
14 10 3 10 0 13 13 9 1 9 2 7 15 13 2
8 13 3 3 10 9 0 9 2
31 10 3 3 13 9 7 9 9 10 9 9 2 10 7 9 3 13 7 13 1 15 7 3 13 10 0 9 10 15 13 2
17 15 3 10 9 13 10 9 2 10 7 13 1 9 7 13 9 2
13 10 3 13 13 15 13 10 9 7 3 10 9 2
15 1 3 3 10 9 3 9 7 9 10 0 9 13 3 2
15 9 3 13 0 9 1 10 9 0 7 3 10 13 0 2
40 1 3 3 9 10 9 9 0 2 10 13 10 9 10 0 2 1 3 9 10 3 9 10 0 7 10 9 10 0 2 1 7 9 10 1 9 9 0 0 2
15 15 3 3 3 1 15 13 13 2 10 7 13 10 9 2
45 10 3 3 1 3 9 7 1 10 9 13 0 3 13 7 10 0 9 9 2 10 7 0 9 1 9 13 9 0 2 15 15 3 16 13 9 13 2 13 9 13 10 9 9 2
14 10 3 9 13 9 3 9 2 9 7 9 3 0 2
14 9 3 3 1 9 13 9 9 2 9 7 1 9 2
36 16 3 13 10 9 13 10 9 10 9 2 10 9 10 13 1 9 13 13 2 10 7 9 15 3 0 13 3 9 10 13 13 1 15 13 2
7 3 1 3 9 15 13 2
25 9 3 9 10 9 1 9 3 3 13 2 0 3 3 0 9 2 1 10 1 10 9 13 9 2
15 0 3 9 0 0 13 1 10 3 9 9 7 10 9 2
23 13 3 9 10 9 9 9 2 15 10 9 3 13 9 0 2 10 7 0 9 9 9 2
14 13 3 15 10 0 9 3 10 9 7 10 13 9 2
32 9 3 0 13 3 3 1 15 13 1 10 9 3 2 3 15 9 13 15 0 13 2 7 13 13 10 10 9 9 13 0 2
21 10 3 3 9 9 10 9 13 0 2 13 15 9 2 1 15 3 13 15 13 2
5 13 3 15 15 2
22 10 3 3 9 10 9 13 9 0 7 0 9 2 10 7 9 13 9 12 7 0 2
13 9 3 13 10 9 0 2 15 13 9 0 13 2
5 13 3 15 9 2
6 15 3 3 15 13 2
36 9 3 9 3 0 13 7 9 2 3 16 16 10 0 9 13 2 0 3 9 15 15 13 9 9 7 9 13 13 2 0 7 3 9 13 2
18 13 3 0 9 3 10 9 10 3 15 3 7 9 13 15 9 13 2
17 3 3 15 3 13 1 15 13 7 9 13 2 3 1 15 13 2
7 9 3 3 1 9 13 2
27 13 3 3 10 3 15 10 9 10 3 9 15 13 10 9 9 13 2 7 10 9 15 9 13 10 9 2
37 9 13 10 3 9 1 9 0 7 0 2 0 1 15 9 13 13 2 3 3 15 1 10 9 13 10 9 13 9 0 2 7 13 10 9 13 2
12 1 3 15 3 10 0 9 13 15 10 9 2
14 13 3 0 0 1 10 9 2 3 3 1 9 13 2
16 9 1 10 9 13 0 15 9 13 9 2 9 7 13 9 2
8 0 10 9 13 9 13 15 2
22 13 10 9 1 9 2 1 10 15 13 3 0 0 7 3 15 7 0 9 13 13 2
21 3 15 3 13 9 0 1 0 10 0 13 2 13 16 10 0 10 0 0 13 2
16 10 3 1 10 0 9 9 13 15 10 9 9 15 15 13 2
67 10 3 3 2 0 13 9 2 0 3 7 0 13 2 13 7 15 9 13 3 0 1 10 9 2 3 16 13 10 1 10 0 9 16 9 13 9 0 1 10 0 13 2 0 13 0 9 2 3 16 13 0 2 13 1 10 9 3 15 13 2 9 7 15 0 13 2
38 0 3 3 13 10 13 2 0 13 10 9 13 1 10 13 2 13 10 9 1 15 0 13 3 13 3 13 3 3 0 13 13 2 7 13 9 3 2
30 13 3 9 7 9 3 0 3 1 10 9 16 0 13 2 13 10 9 1 15 7 13 15 9 2 13 1 10 13 2
18 3 3 10 3 9 13 7 15 1 9 13 2 7 1 9 0 13 2
7 15 3 13 13 15 13 2
27 3 3 13 15 13 9 2 10 9 13 0 1 0 9 3 13 7 13 2 1 10 15 13 9 15 13 2
16 10 3 13 15 9 3 15 0 10 9 13 7 13 15 0 2
6 13 3 15 10 9 2
25 13 3 3 15 9 0 3 7 0 2 3 15 13 10 9 2 7 0 15 13 1 0 9 13 2
21 10 3 16 13 10 9 2 10 9 13 0 9 13 7 15 13 10 15 0 13 2
23 13 3 3 15 10 9 13 9 0 3 7 0 0 15 3 9 13 2 0 0 9 13 2
18 13 3 3 0 10 9 16 10 0 10 0 9 10 9 0 13 0 2
21 10 3 3 15 3 10 9 13 9 13 16 15 13 2 10 7 3 3 15 13 2
18 9 3 13 10 0 0 2 1 3 10 0 10 9 13 7 10 9 2
15 10 3 15 0 13 9 1 10 9 9 3 3 10 9 2
10 3 10 0 9 10 9 13 13 9 2
24 15 3 3 10 9 15 3 13 7 1 10 15 9 2 10 7 0 9 1 13 10 9 13 2
16 16 3 15 13 7 13 15 10 9 2 13 10 0 13 0 2
17 3 10 3 9 13 3 1 15 13 2 7 15 13 10 13 13 2
13 15 3 1 10 9 13 2 15 7 0 13 15 2
28 16 15 13 13 2 15 16 13 1 0 0 9 13 2 7 10 9 3 7 0 13 1 0 10 9 15 13 2
12 9 3 3 10 0 9 13 0 7 15 13 2
7 9 3 3 9 13 15 2
43 9 3 9 13 9 2 15 13 9 2 13 9 7 0 9 2 13 10 9 2 13 7 3 13 0 9 13 2 7 13 1 10 9 0 3 15 13 7 0 9 0 13 2
75 3 3 13 0 0 9 3 0 0 2 13 10 9 1 15 1 0 13 9 2 1 15 13 1 10 9 7 9 15 15 9 13 7 13 0 0 2 3 7 13 13 3 0 3 13 2 3 3 15 3 13 2 1 15 3 13 10 9 0 3 13 2 13 0 7 0 9 2 7 10 9 15 10 0 2
11 9 3 13 13 9 10 9 10 9 9 2
9 1 10 3 3 13 0 3 13 2
25 15 10 10 9 13 13 16 9 10 9 13 15 13 2 7 10 10 9 9 3 9 0 13 15 2
23 13 3 10 1 15 13 0 13 1 10 9 2 13 3 10 9 7 10 9 0 13 13 2
27 3 15 2 16 13 13 10 9 2 13 10 9 13 9 9 0 2 13 7 15 9 10 9 9 9 9 2
23 10 13 3 1 10 9 9 13 1 10 9 2 15 7 13 13 3 1 10 0 9 13 2
23 3 3 10 3 9 3 13 2 7 10 3 9 0 0 13 2 1 9 13 10 0 9 2
15 3 10 3 9 13 10 9 7 13 10 9 10 9 13 2
8 10 3 9 10 9 0 13 2
6 3 3 13 1 9 2
23 3 16 13 1 10 9 9 2 9 15 9 9 13 9 3 7 9 13 10 3 3 13 2
29 10 3 16 13 3 13 10 9 1 9 9 2 10 0 9 13 0 2 0 0 15 13 13 10 0 9 10 9 2
19 13 3 0 10 9 2 16 15 13 13 2 0 0 9 0 0 10 9 2
28 3 3 10 1 9 9 3 13 2 16 0 9 13 2 7 10 1 9 9 13 10 13 1 0 10 9 13 2
21 10 3 10 9 13 10 9 10 1 9 7 10 15 3 0 13 10 9 0 9 2
29 3 3 13 3 10 9 1 15 15 13 2 7 13 1 15 10 13 1 10 0 9 16 13 15 13 9 10 9 2
25 1 3 3 0 7 0 9 13 10 9 10 9 2 7 10 0 15 1 3 9 7 9 0 13 2
23 3 3 3 9 13 1 0 15 0 13 2 1 7 10 9 13 13 15 15 0 13 0 2
24 1 3 15 9 3 2 13 0 9 1 15 9 13 2 13 2 13 7 9 9 9 10 9 2
9 3 15 13 9 15 9 13 9 2
22 10 13 9 1 10 9 13 15 16 13 3 10 15 9 2 13 7 3 10 9 0 2
16 13 3 10 9 10 9 10 9 2 13 1 15 15 0 13 2
22 3 3 10 9 0 13 3 9 0 9 3 10 15 0 15 13 9 2 13 10 9 2
27 10 3 9 13 15 9 13 9 2 15 13 9 3 13 0 9 7 0 2 0 3 13 15 9 9 9 2
36 13 3 10 9 10 9 2 10 9 10 0 9 13 0 9 2 13 7 15 1 10 9 10 9 0 13 9 2 10 7 9 13 10 9 0 2
27 13 3 15 7 13 10 9 2 13 1 10 9 10 9 9 13 2 13 7 13 13 10 13 1 15 13 2
21 1 3 15 10 9 10 10 9 9 13 16 13 10 10 9 15 9 13 1 15 2
30 15 3 3 13 10 9 2 16 13 10 9 2 13 9 9 0 7 0 3 9 7 0 0 10 15 2 13 15 15 2
20 13 15 9 13 9 2 13 7 1 15 13 2 3 7 13 9 0 15 13 2
16 3 16 3 0 15 3 13 2 13 3 10 3 0 13 3 2
20 15 13 10 9 2 16 15 13 10 9 13 10 1 9 13 13 1 10 9 2
12 13 3 13 10 15 9 10 0 9 13 9 2
14 10 3 1 15 13 3 3 15 0 1 9 13 13 2
31 10 3 13 3 15 13 9 2 3 16 13 3 7 13 0 16 3 13 2 3 15 15 13 10 9 7 1 9 0 13 2
32 16 3 13 15 13 1 10 9 0 13 10 9 2 15 3 10 9 13 1 15 2 0 15 16 13 10 3 15 9 10 0 2
25 3 10 3 0 1 15 13 0 13 10 9 2 13 7 10 15 9 0 9 13 7 3 10 0 2
21 15 13 7 3 9 13 1 10 9 10 9 15 13 9 3 0 13 7 9 0 2
14 16 3 10 9 9 0 13 13 2 13 10 9 15 2
19 13 15 9 10 9 0 13 13 1 10 0 10 9 2 16 3 0 13 2
6 13 3 13 13 15 2
19 15 13 10 9 3 13 10 9 13 10 0 3 9 7 13 1 10 9 2
24 10 3 3 3 15 10 9 2 9 13 0 9 2 3 3 1 9 13 13 10 9 1 9 2
21 16 3 13 13 2 0 1 0 13 10 9 13 0 15 0 15 3 3 9 13 2
13 9 3 0 9 9 13 2 15 7 13 13 3 2
20 16 3 0 13 2 13 9 13 13 3 7 13 2 13 9 3 7 9 0 2
37 9 3 16 13 15 2 13 10 0 13 10 9 13 13 7 13 3 0 13 10 9 2 13 9 13 10 15 13 15 2 0 13 16 3 15 13 2
11 3 15 13 13 2 13 10 15 9 13 2
9 3 3 3 3 13 3 3 13 2
18 13 3 13 9 3 7 9 13 2 1 7 3 9 13 0 1 9 2
5 3 3 15 13 2
10 3 3 15 13 10 9 7 13 13 2
25 10 3 16 13 10 9 0 3 7 0 13 2 13 7 13 10 9 10 9 13 0 9 13 15 2
11 10 3 3 13 0 3 13 3 15 13 2
14 16 3 3 13 3 10 9 2 0 13 10 9 15 2
21 16 3 3 13 15 13 3 13 2 15 3 3 13 2 16 3 0 9 13 13 2
9 13 3 3 15 2 13 7 13 2
17 15 3 13 13 2 10 7 10 9 9 9 3 1 15 13 13 2
14 3 3 3 15 13 13 10 9 7 15 3 13 13 2
15 10 3 3 13 0 9 13 7 10 13 3 13 10 9 2
18 3 3 13 10 9 1 10 13 3 13 10 9 2 7 3 13 15 2
29 0 3 13 13 9 2 15 3 13 10 15 9 2 10 7 15 13 0 13 13 1 10 9 1 15 13 10 0 2
17 13 3 10 9 0 10 0 9 2 13 1 10 0 10 9 13 2
36 16 3 0 9 10 9 13 13 2 13 1 9 10 9 2 10 15 9 9 3 13 2 13 7 1 10 9 13 13 0 13 10 9 10 9 2
47 13 3 10 9 10 15 0 10 0 13 3 1 15 7 13 10 9 10 9 2 7 10 3 13 2 10 7 0 15 9 13 13 13 10 9 10 9 2 9 0 3 0 7 3 9 13 2
15 3 16 13 0 10 9 2 9 1 0 15 13 13 15 2
21 13 1 10 9 0 1 15 13 3 10 9 0 2 13 7 1 15 0 1 9 2
37 10 3 15 13 10 3 9 13 2 10 3 0 13 2 10 7 3 0 15 9 9 13 2 10 7 0 10 9 13 13 9 2 3 0 9 13 2
45 9 3 0 10 9 13 2 13 9 9 9 0 1 9 2 3 3 3 13 10 13 1 10 9 2 13 15 10 0 9 13 2 13 7 10 9 10 9 10 9 3 3 13 13 2
23 13 3 7 13 9 2 13 13 10 9 9 10 9 1 2 13 10 3 9 7 10 9 2
31 16 3 13 0 2 13 1 10 9 10 9 13 15 3 13 15 0 13 9 13 10 15 9 13 0 1 15 9 0 13 2
5 10 3 13 3 2
19 10 3 15 1 10 9 9 2 15 3 15 13 2 13 0 15 13 9 2
8 13 3 15 13 1 15 0 2
24 10 3 3 0 9 10 13 13 2 15 7 13 3 7 9 13 0 2 1 15 13 10 9 2
14 16 3 3 15 1 0 0 0 13 2 15 10 13 2
8 13 3 15 1 9 0 13 2
23 9 3 15 3 3 13 13 13 1 9 0 13 2 3 7 13 15 13 10 0 13 15 2
13 10 3 13 1 10 9 3 3 13 10 13 9 2
21 13 3 1 9 13 10 9 13 2 3 13 1 9 3 7 9 15 13 13 15 2
25 9 3 10 3 9 10 9 13 9 3 3 0 13 2 9 7 3 3 13 13 15 10 0 13 2
28 16 3 15 13 10 9 2 13 15 10 9 9 2 0 3 9 10 9 13 15 15 13 1 9 13 10 0 2
25 10 3 9 16 13 10 9 3 13 2 3 13 1 0 9 2 16 3 13 13 2 7 13 15 2
4 13 3 3 2
17 13 10 9 0 13 10 9 2 13 15 7 13 10 13 13 15 2
7 3 13 15 3 3 13 2
5 15 3 13 3 2
28 13 3 15 1 15 13 2 13 15 1 0 9 7 13 13 1 3 13 2 13 0 15 16 3 0 0 13 2
23 16 3 13 15 10 13 13 10 9 2 13 10 9 10 0 3 13 1 15 7 13 15 2
8 9 3 3 10 0 13 9 2
48 9 3 13 15 15 13 9 1 10 13 2 0 3 2 1 3 13 15 1 10 9 15 9 2 3 13 10 9 2 3 7 16 15 13 2 13 13 16 13 3 10 9 7 10 13 13 3 2
23 10 3 3 13 13 13 1 10 9 0 13 3 2 7 9 10 0 13 3 1 0 13 2
32 9 3 16 13 15 2 13 7 0 13 16 3 10 9 10 1 13 13 7 16 1 9 0 1 9 13 2 13 1 10 9 2
48 16 3 10 9 13 10 9 13 15 3 0 9 7 10 9 2 10 3 15 7 0 9 13 9 0 9 9 2 9 7 10 9 10 15 2 1 9 3 7 0 9 3 7 9 2 0 0 2
27 15 3 3 13 1 9 13 2 16 7 10 9 13 3 13 10 9 2 9 13 15 16 13 15 10 9 2
34 13 3 9 3 3 13 2 13 15 13 10 9 10 9 13 3 10 9 7 10 9 2 9 7 13 13 13 3 7 13 15 13 15 2
21 13 3 10 9 7 13 13 10 9 10 9 2 13 7 3 13 3 7 15 13 2
12 13 3 15 10 9 16 13 0 9 9 13 2
14 10 3 3 13 13 7 0 13 0 15 3 9 13 2
27 15 3 13 7 13 10 0 10 9 13 1 10 9 2 3 7 13 2 16 15 13 2 13 13 10 0 2
23 9 3 9 9 0 13 2 9 7 1 13 13 10 15 10 9 15 10 9 15 3 13 2
11 13 3 13 10 9 15 13 15 10 9 2
19 10 3 1 15 13 13 16 13 13 10 9 2 16 13 7 3 13 0 2
6 10 3 13 15 15 2
20 13 3 10 9 7 13 2 7 15 1 9 13 10 1 10 9 9 13 9 2
12 10 3 0 0 3 10 0 9 9 13 13 2
14 3 3 0 3 9 3 9 7 10 0 0 13 13 2
9 3 3 1 15 15 15 13 13 2
25 13 10 9 16 3 13 3 7 13 10 9 3 1 9 0 2 13 3 15 1 7 9 13 0 2
7 3 3 3 10 0 13 2
21 1 0 3 3 10 9 15 0 13 2 7 10 3 10 9 13 3 1 0 13 2
5 13 10 9 15 2
19 3 3 3 3 13 15 3 13 15 13 0 13 9 3 10 0 7 15 2
28 3 3 3 13 1 10 9 0 13 13 9 2 7 15 13 9 13 3 7 9 0 13 1 9 2 13 9 2
19 15 3 13 9 2 13 9 2 3 13 10 9 7 9 1 15 0 13 2
12 3 3 3 15 15 7 10 0 9 13 13 2
17 3 3 13 10 9 1 0 2 15 3 13 7 15 0 15 13 2
14 10 3 9 0 1 9 13 1 9 3 7 10 13 2
14 13 15 10 9 13 3 7 13 10 9 13 15 15 2
13 3 3 13 13 1 9 2 9 7 15 3 13 2
19 13 3 3 9 3 7 9 13 3 1 9 3 10 9 7 10 9 15 2
8 15 13 10 9 13 10 9 2
32 13 3 15 1 10 9 10 9 13 10 13 2 3 13 16 13 2 3 13 0 3 13 3 3 13 2 13 7 0 9 13 2
24 10 3 15 13 2 13 1 10 3 3 13 7 13 0 2 1 9 7 13 0 10 15 9 2
27 13 3 13 1 10 10 9 9 2 13 3 15 13 1 0 2 13 7 15 1 10 9 10 0 10 9 2
26 10 3 9 13 10 9 0 2 16 3 13 10 9 13 15 10 9 2 13 9 16 13 9 9 13 2
7 3 3 10 9 0 13 2
20 9 3 13 7 13 10 0 0 7 0 13 10 9 9 13 2 13 9 13 2
27 1 15 3 13 9 3 13 9 13 1 9 2 9 7 13 13 13 0 2 10 9 10 9 10 15 13 2
8 1 3 3 15 15 15 13 2
26 13 10 9 0 1 10 9 2 13 9 0 10 9 10 0 9 13 16 13 9 13 9 13 10 9 2
24 9 13 2 3 13 15 10 9 7 15 13 2 16 3 13 3 13 9 2 13 15 15 13 2
41 13 3 10 9 10 9 2 7 9 13 3 9 10 9 10 0 2 13 1 10 9 2 13 15 1 9 13 10 9 9 13 0 15 13 7 15 15 15 13 13 2
14 15 3 3 3 0 13 7 10 9 13 10 9 13 2
16 13 3 1 15 10 9 0 13 13 2 10 7 9 13 0 2
9 3 3 3 3 1 15 9 13 2
8 15 3 9 10 15 9 13 2
17 1 3 3 10 15 9 13 2 10 7 1 9 3 7 15 13 2
18 15 3 2 16 13 0 13 2 0 3 9 13 9 2 15 0 13 2
8 9 3 13 13 13 1 9 2
25 3 16 3 15 1 9 13 9 0 15 2 13 15 15 15 13 2 16 7 10 15 0 0 9 2
14 0 3 15 13 1 15 7 13 1 15 9 13 13 2
15 3 3 0 10 3 3 13 2 13 15 7 13 1 9 2
19 13 15 10 9 13 0 9 0 9 13 13 2 13 7 13 15 0 13 2
4 13 3 15 2
25 13 1 9 15 13 2 9 10 9 13 2 3 7 13 10 9 7 13 13 9 15 9 9 13 2
5 9 3 15 13 2
19 13 3 9 0 9 2 7 10 3 15 10 9 13 7 13 13 1 9 2
19 15 9 13 0 2 1 10 7 9 13 9 2 3 10 9 10 9 13 2
17 13 3 10 9 10 13 9 2 0 15 13 1 10 0 13 13 2
38 1 3 15 10 3 9 3 10 9 7 10 9 10 9 0 10 9 13 1 15 13 7 13 3 13 10 9 9 2 1 3 9 3 7 9 3 0 2
11 13 3 10 0 10 9 13 1 9 13 2
22 16 3 1 9 13 2 13 15 10 9 0 15 10 0 13 7 15 13 15 13 0 2
9 10 3 13 0 13 15 10 0 2
30 13 3 15 13 13 15 3 7 15 0 0 2 0 9 0 13 2 3 13 7 15 13 13 15 9 10 0 0 0 2
7 3 3 15 13 13 0 2
26 15 3 3 13 0 9 13 15 1 9 13 2 7 15 13 9 9 13 3 0 3 15 7 10 0 2
11 3 3 13 3 2 13 1 9 10 0 2
16 9 3 3 9 13 0 13 2 7 3 0 13 1 9 13 2
13 9 3 16 13 9 15 13 2 13 9 13 15 2
17 10 3 9 13 10 9 13 16 0 13 1 15 16 9 0 13 2
25 13 3 15 10 9 9 3 13 0 2 7 9 15 3 0 13 9 13 2 13 13 15 15 13 2
24 13 3 10 0 9 3 2 16 13 0 10 9 2 13 13 10 9 3 3 16 9 3 13 2
21 13 3 15 7 13 10 9 13 2 7 0 3 9 13 7 15 13 10 9 13 2
49 13 3 0 10 9 13 10 9 13 3 7 13 2 3 0 13 1 15 0 9 2 7 3 3 13 15 1 10 15 9 2 15 15 15 9 10 9 13 2 15 0 13 10 15 9 1 10 9 2
12 10 3 15 13 13 16 15 13 10 9 9 2
15 9 3 13 2 15 3 13 2 10 9 15 3 3 13 2
44 9 3 3 13 1 9 0 7 0 3 10 9 13 2 9 7 13 9 1 10 15 9 2 13 10 1 9 9 9 1 9 0 7 0 9 13 2 3 16 0 10 9 13 2
20 0 3 9 13 3 15 15 13 7 13 1 9 2 13 7 3 13 9 13 2
20 3 3 1 9 10 9 3 7 10 9 13 10 9 13 10 1 0 10 9 2
15 9 3 9 0 15 0 13 13 1 15 2 1 15 13 2
30 3 3 9 13 3 7 13 13 7 9 9 15 13 9 13 2 16 13 15 0 2 15 7 13 3 0 10 9 13 2
43 9 3 13 9 0 13 2 9 3 3 9 7 9 3 1 9 13 13 2 7 3 10 13 9 13 2 16 3 15 13 2 16 3 0 13 10 9 16 3 10 9 13 2
22 10 3 13 9 3 1 10 0 10 9 13 9 13 2 10 9 0 10 9 9 13 2
15 13 3 9 3 3 9 3 9 3 9 3 9 7 9 2
21 15 3 3 13 0 3 2 13 7 3 10 9 13 2 1 3 9 13 7 9 2
15 13 3 9 10 9 9 2 9 3 9 2 9 7 9 2
11 9 3 10 9 1 10 13 9 0 13 2
22 3 9 13 7 9 13 13 13 2 3 9 13 2 3 9 2 3 9 2 7 9 2
23 10 3 16 0 13 13 2 1 9 0 13 10 9 13 10 9 2 13 10 9 9 3 2
25 0 3 3 10 13 0 0 3 15 13 13 0 2 10 7 10 0 9 13 3 13 7 10 9 2
10 1 3 3 10 0 9 3 15 13 2
28 16 3 13 1 9 10 9 13 10 9 13 9 3 0 2 3 7 10 9 2 1 15 13 3 0 10 9 2
17 13 3 15 9 9 13 13 9 2 0 3 15 13 13 10 9 2
11 1 3 3 9 3 15 9 13 9 13 2
17 13 3 0 9 13 10 13 10 9 7 13 15 0 15 9 13 2
11 9 3 0 3 0 13 13 15 0 13 2
10 1 15 3 0 9 10 15 13 13 2
28 1 10 10 0 15 9 3 9 3 9 7 9 13 0 0 1 9 2 10 7 9 15 10 9 10 9 13 2
12 9 3 0 13 2 9 7 0 7 3 0 2
20 3 1 15 13 9 10 9 13 13 13 2 16 15 1 9 13 15 9 0 2
16 9 3 3 13 2 7 15 3 13 13 2 3 13 0 15 2
15 15 3 3 3 13 2 13 7 13 13 10 0 10 9 2
38 15 3 3 13 15 13 2 15 10 0 13 13 10 9 2 1 15 3 13 13 2 7 16 3 13 7 13 2 13 15 2 16 7 3 13 2 13 2
9 10 3 16 13 13 2 13 13 2
17 13 3 15 1 10 9 2 15 3 15 13 16 0 13 10 13 2
9 1 3 10 13 15 13 10 9 2
11 16 3 13 0 0 0 2 10 9 13 2
12 16 3 0 13 0 0 2 13 13 10 0 2
17 13 3 1 0 10 0 15 13 1 3 15 2 0 7 10 0 2
7 3 3 1 9 13 13 2
37 0 3 10 15 3 13 1 9 13 2 13 15 13 9 0 10 0 0 2 10 3 15 1 9 10 9 13 2 10 7 3 13 1 15 0 13 2
10 13 3 3 10 9 9 3 7 13 2
8 0 3 0 9 13 9 3 2
21 3 3 3 10 0 9 13 10 15 13 0 13 2 7 1 10 9 10 0 9 2
16 3 9 3 0 13 13 2 7 3 3 1 9 13 9 13 2
16 13 3 0 15 0 3 0 9 2 0 7 3 0 9 13 2
17 9 3 0 13 2 1 10 13 13 0 2 15 3 0 13 9 2
12 10 3 10 0 13 9 13 9 1 0 9 2
7 10 0 3 13 0 13 2
20 3 3 16 0 13 2 3 13 1 9 10 9 2 7 1 10 9 9 13 2
19 3 13 16 13 0 3 7 0 10 9 13 10 9 2 3 10 9 13 2
29 13 3 15 3 13 10 15 9 7 9 2 7 0 3 15 13 2 0 9 13 13 15 13 3 0 13 7 0 2
12 15 3 15 13 3 13 2 15 3 13 13 2
31 0 3 15 10 13 13 2 0 7 10 13 9 2 0 3 7 0 1 2 3 7 0 13 13 10 13 3 0 9 13 2
21 15 3 3 10 9 9 7 9 13 2 1 9 15 3 13 7 13 10 0 9 2
11 13 3 15 1 10 9 13 15 15 13 2
23 9 3 0 10 13 1 15 0 13 1 10 9 2 7 10 0 9 2 10 0 9 13 2
18 3 15 0 15 3 13 13 2 15 9 3 0 13 2 15 3 3 2
21 1 15 13 13 13 10 9 10 9 2 3 10 3 10 3 7 2 7 0 3 2
9 15 3 3 13 1 15 13 13 2
28 15 3 3 13 13 3 3 3 1 10 13 2 16 3 0 13 9 9 10 9 16 3 1 9 7 9 13 2
8 9 3 3 3 13 15 13 2
5 3 3 3 13 2
9 13 3 3 10 9 9 9 13 2
14 9 3 13 0 10 3 0 9 7 10 1 9 9 2
13 10 3 3 13 0 15 13 2 16 3 0 13 2
30 10 3 3 9 9 0 1 9 7 9 13 2 7 9 0 0 13 2 13 3 9 3 3 9 3 0 9 7 0 2
19 3 1 3 10 9 0 13 16 3 3 13 2 13 7 1 10 0 9 2
31 9 3 7 9 2 16 10 9 0 13 1 9 2 13 9 1 9 1 9 2 13 1 10 15 13 15 3 9 13 0 2
26 10 3 13 15 15 13 13 15 9 2 9 13 9 13 9 1 10 9 13 2 13 15 13 1 9 2
41 9 3 0 10 9 10 9 7 10 9 15 1 13 2 16 3 10 9 0 0 9 13 1 9 13 15 1 9 3 13 2 3 7 13 10 9 13 0 13 9 2
9 10 3 3 9 13 13 15 15 2
24 9 3 16 13 15 13 1 10 9 2 9 3 13 0 7 13 1 9 10 15 2 1 9 2
13 1 0 3 15 9 9 13 1 15 3 10 9 2
15 10 3 0 9 13 0 9 13 9 1 9 13 9 13 2
29 10 3 9 0 2 15 3 10 9 13 2 10 3 9 7 10 9 1 10 0 13 13 9 0 9 15 15 13 2
13 9 3 3 10 0 15 13 2 7 9 9 9 2
16 9 3 15 0 13 9 1 9 2 3 7 9 3 7 9 2
16 0 3 10 9 10 0 13 13 1 9 15 2 15 7 13 2
15 9 3 3 7 9 1 15 13 2 9 7 1 15 0 2
6 15 9 9 9 13 2
25 0 3 3 10 9 10 9 3 13 1 9 10 9 2 9 13 2 10 7 15 9 13 0 15 2
13 3 3 9 13 3 9 0 7 0 10 9 9 2
33 13 3 1 10 0 9 15 1 0 3 15 2 0 7 13 10 0 3 0 9 2 0 3 13 0 10 9 10 0 7 9 0 2
11 16 3 3 9 2 13 0 0 9 0 2
29 10 3 3 0 9 7 10 9 13 10 9 2 3 13 9 13 2 7 3 3 13 15 10 0 15 13 10 9 2
24 9 3 9 2 15 9 13 9 2 13 10 9 13 2 13 7 1 10 15 9 13 10 0 2
9 15 3 3 15 0 10 9 13 2
12 0 0 9 3 9 13 7 3 3 9 13 2
30 15 3 1 3 10 9 0 9 13 2 16 7 3 15 3 15 9 13 10 0 9 7 0 15 13 2 9 0 13 2
7 15 3 13 13 1 9 2
27 9 3 13 10 3 15 9 1 9 10 9 13 2 10 3 9 9 1 9 10 9 2 10 7 3 0 2
19 3 3 13 10 9 3 15 10 0 9 2 13 3 7 10 3 13 9 2
13 13 3 0 9 0 1 9 13 7 9 13 9 2
8 13 3 0 1 9 7 9 2
15 15 3 0 9 3 13 9 2 7 15 1 9 0 9 2
19 10 3 9 13 10 9 9 0 1 9 13 2 0 13 1 9 9 0 2
28 10 3 9 13 10 9 9 1 9 9 13 9 3 2 1 15 13 1 10 9 9 13 9 15 13 9 9 2
27 13 3 3 0 10 9 9 15 2 7 3 9 0 3 0 1 0 9 13 2 16 3 10 9 10 9 2
7 15 0 9 9 10 0 2
8 0 3 0 13 9 1 9 2
17 0 3 10 9 9 3 13 13 0 9 2 9 7 13 3 3 2
6 9 3 3 13 9 2
11 0 9 9 13 7 13 1 10 9 13 2
22 3 3 10 9 10 9 13 10 9 9 1 9 13 9 2 10 9 13 13 10 9 2
16 13 3 0 9 2 9 13 10 9 13 10 9 13 9 9 2
15 13 3 15 9 13 15 10 0 9 7 13 15 0 9 2
15 15 3 3 10 9 9 9 2 1 10 1 10 9 13 2
4 13 3 15 2
13 10 3 0 9 13 3 9 13 15 3 15 13 2
22 10 3 0 3 9 13 2 16 3 13 0 13 9 2 7 13 13 0 13 15 13 2
13 9 3 3 3 13 2 7 13 15 3 13 9 2
30 10 3 3 13 2 9 7 13 10 9 10 9 3 13 9 9 2 16 3 15 13 2 9 10 3 9 9 7 9 2
23 15 13 10 9 2 13 9 13 10 13 15 9 15 13 9 0 7 0 9 15 15 13 2
21 3 13 3 9 0 2 15 13 9 1 0 10 9 13 1 15 13 15 13 13 2
16 10 2 16 15 13 2 3 10 9 9 13 0 7 10 0 2
20 0 1 10 0 9 13 10 9 10 9 2 16 9 13 9 3 7 9 13 2
16 0 3 10 9 9 15 13 13 2 7 15 13 10 3 9 2
46 1 15 13 10 3 9 9 9 9 2 10 7 9 10 3 9 7 10 10 0 9 9 9 9 13 2 13 15 1 9 2 9 3 3 13 7 10 9 1 0 9 13 10 0 13 2
47 16 3 13 10 9 1 10 9 2 10 9 13 10 9 1 3 9 7 9 2 13 7 1 9 2 16 10 9 13 0 10 1 10 9 2 9 3 13 7 10 0 9 13 1 15 13 2
12 13 3 1 10 9 13 9 13 1 10 9 2
12 13 3 1 9 15 10 9 13 1 9 15 2
13 3 13 9 2 16 13 2 9 13 7 15 13 2
7 13 16 9 13 13 15 2
17 3 3 15 3 3 13 13 3 16 15 9 13 10 9 15 13 2
30 3 3 3 15 9 10 3 0 15 16 9 13 15 13 13 2 0 7 9 10 9 13 2 7 3 13 16 15 13 2
20 10 3 3 15 3 13 13 2 10 7 13 15 2 13 16 0 13 10 9 2
13 10 3 3 0 15 3 13 7 15 9 13 13 2
16 9 3 9 13 15 15 13 2 16 3 13 7 0 15 13 2
13 9 3 13 10 9 7 13 10 9 13 15 13 2
39 13 3 9 9 9 2 15 3 15 13 13 9 15 10 9 13 2 7 3 13 10 15 0 15 1 9 1 9 13 2 0 7 9 3 13 13 1 15 2
29 10 3 3 15 1 10 9 13 13 1 9 10 9 2 9 7 13 3 13 9 1 15 13 13 13 13 1 9 2
50 9 3 10 9 13 1 10 9 10 9 9 9 0 3 3 13 2 16 3 13 3 13 10 1 9 1 9 2 0 3 10 9 13 10 9 9 13 2 1 15 7 9 9 10 0 9 10 9 13 2
13 9 3 1 15 13 1 10 9 9 13 13 9 2
13 10 3 9 13 9 1 1 9 13 10 1 9 2
17 13 3 3 9 1 0 13 2 15 9 3 0 7 9 13 13 2
11 10 3 9 0 13 10 9 1 9 9 2
18 13 3 10 9 1 10 9 0 13 1 9 0 15 13 9 13 13 2
10 13 3 15 15 9 13 13 9 9 2
11 15 3 16 13 13 10 9 2 13 13 2
48 13 3 15 10 9 2 9 10 9 9 10 9 13 0 13 3 13 15 9 2 13 3 10 9 7 13 10 0 3 13 3 2 1 15 10 0 1 9 13 13 0 0 2 15 3 9 13 2
11 13 3 1 9 13 1 0 9 13 15 2
9 10 3 15 13 2 13 9 13 2
19 10 3 15 13 2 10 7 3 10 0 15 9 13 2 13 13 9 9 2
9 1 15 10 9 1 9 13 15 2
18 13 10 9 9 13 10 9 7 15 0 13 13 9 9 1 10 9 2
8 10 9 15 1 10 9 13 2
23 15 16 13 13 10 9 2 3 13 3 13 13 7 1 15 13 13 2 13 15 1 9 2
8 3 3 13 15 3 13 3 2
4 3 3 13 2
19 9 3 16 13 15 13 1 10 9 2 13 9 1 9 13 9 1 9 2
11 3 3 1 0 9 0 13 1 9 13 2
9 13 3 10 9 1 10 9 9 2
12 10 3 9 0 13 9 10 9 2 9 0 2
14 9 3 3 13 10 9 13 1 9 2 13 9 13 2
37 9 3 3 9 13 2 9 7 1 15 13 1 10 13 9 2 7 15 3 9 13 2 15 7 9 9 0 13 9 13 10 9 2 9 7 3 2
7 1 3 15 3 9 13 2
18 0 9 3 1 9 9 13 16 13 1 10 9 2 13 10 9 9 2
14 16 3 0 13 2 10 3 9 13 1 10 9 13 2
6 0 3 9 9 13 2
28 10 3 9 0 9 0 0 9 13 2 7 10 3 9 3 10 0 3 10 9 7 10 9 15 13 10 13 2
8 13 3 3 0 9 7 9 2
32 13 3 1 10 9 0 13 10 9 10 9 2 15 9 3 13 2 9 2 13 3 9 12 9 2 13 7 0 12 7 12 2
26 0 3 10 9 0 10 9 3 3 15 13 16 10 3 0 15 13 9 13 10 15 9 13 3 13 2
33 3 3 2 16 15 3 3 13 10 9 2 10 3 13 10 9 1 15 16 13 2 13 15 9 9 13 10 9 2 13 7 3 2
21 3 3 3 10 9 10 9 3 0 9 13 2 15 7 0 9 0 7 3 13 2
10 10 3 3 9 10 9 9 0 13 2
15 10 3 9 13 10 9 13 13 13 9 0 7 3 13 2
15 1 15 3 13 15 2 13 15 13 10 9 1 10 9 2
18 10 3 9 13 13 3 3 15 15 13 13 2 3 7 15 13 13 2
9 10 3 9 13 9 13 10 9 2
18 1 3 10 9 12 9 0 15 1 9 13 9 2 15 9 13 9 2
6 9 3 3 9 13 2
25 13 3 1 10 9 2 0 13 1 10 9 13 10 9 10 9 2 15 13 13 1 9 10 9 2
32 13 3 15 1 10 9 2 0 10 9 13 9 3 7 9 10 9 7 10 9 10 9 2 0 7 13 13 3 1 10 9 2
13 10 3 15 10 9 13 2 13 1 10 9 13 2
21 16 3 1 10 9 13 2 13 3 1 10 0 13 1 9 12 2 7 9 13 2
20 10 3 9 13 3 15 10 9 2 13 9 12 2 13 1 10 9 13 9 2
11 13 3 10 9 0 0 9 10 9 13 2
16 10 3 3 12 15 9 13 2 10 7 12 10 13 13 0 2
5 13 3 10 9 2
33 13 3 1 10 9 13 10 9 3 10 9 7 10 0 9 0 0 3 13 10 9 15 13 2 7 3 13 10 9 13 1 9 2
29 10 3 13 9 10 9 10 3 9 7 10 9 13 2 10 7 9 10 9 13 3 15 0 0 7 15 13 13 2
11 10 3 9 1 9 13 13 13 10 9 2
14 10 3 9 15 13 13 15 3 3 10 9 3 13 2
12 3 3 13 15 3 7 9 0 7 0 13 2
29 3 15 3 10 9 0 9 13 2 10 7 15 1 10 9 13 3 13 13 9 9 10 9 0 15 3 9 13 2
16 9 3 3 1 10 1 9 3 13 0 3 15 7 9 13 2
50 16 3 15 13 9 10 9 9 2 13 0 1 10 9 13 13 1 10 9 2 7 3 13 9 9 2 15 0 15 0 9 13 3 13 2 7 1 9 13 9 3 1 9 10 1 9 16 9 13 2
13 15 3 3 9 0 10 9 3 13 13 10 9 2
39 10 3 0 9 1 9 1 9 3 13 9 16 3 10 13 2 7 9 13 0 1 10 15 0 13 2 13 7 7 13 13 1 9 0 7 10 13 13 2
16 9 3 2 16 3 0 15 13 2 0 9 9 13 9 13 2
7 3 3 10 0 9 13 2
22 16 3 10 1 10 9 9 13 9 2 10 10 9 13 9 13 15 15 0 13 9 2
31 13 3 9 7 13 15 0 1 10 9 2 13 9 9 9 9 13 9 0 2 15 16 13 2 13 3 15 13 9 3 2
13 13 3 15 1 10 9 3 13 13 9 3 13 2
8 15 3 3 15 9 0 13 2
20 9 3 13 9 13 9 1 9 3 9 7 9 2 3 13 3 9 7 9 2
13 13 3 15 9 3 13 1 10 9 1 10 9 2
28 10 3 0 13 9 0 7 13 9 13 10 9 2 9 3 0 13 2 0 3 15 0 13 1 0 13 9 2
12 10 3 2 16 9 13 2 13 15 10 9 2
28 16 3 9 3 13 9 0 16 13 10 9 2 10 0 13 9 0 10 9 0 1 0 3 10 9 0 3 2
11 3 15 0 9 13 2 15 10 9 13 2
28 3 3 1 10 9 9 13 9 13 10 13 7 1 10 9 10 9 13 2 7 9 9 15 13 10 13 0 2
28 3 3 1 9 13 10 9 0 15 3 13 9 13 2 9 0 13 2 1 10 9 3 7 10 0 9 13 2
23 3 3 10 9 9 9 0 9 3 7 9 13 1 10 9 2 7 3 1 10 9 13 2
9 3 3 3 9 3 9 13 13 2
28 3 3 15 3 13 15 10 9 2 7 13 15 15 13 0 9 2 3 10 9 10 0 3 13 15 3 3 2
11 10 3 9 7 10 9 13 13 9 9 2
20 15 3 3 13 2 0 7 13 0 9 0 10 9 13 2 15 3 3 1 2
15 10 3 9 0 13 15 13 2 15 7 1 9 13 13 2
41 13 3 1 9 1 10 9 10 9 9 9 3 7 9 2 16 13 10 9 9 2 13 0 3 9 7 10 9 3 2 10 7 13 13 10 9 1 9 10 9 2
19 15 3 3 9 13 2 15 10 0 13 9 2 10 7 9 3 9 13 2
35 16 3 1 9 9 10 9 2 13 3 15 1 10 9 9 2 13 1 10 9 1 9 2 3 3 1 10 9 10 9 9 1 9 13 2
10 9 3 10 3 0 10 7 0 13 2
11 0 3 15 0 13 7 0 15 13 9 2
11 13 1 10 9 15 7 3 1 10 9 2
18 13 3 0 10 0 15 13 2 13 15 3 7 10 9 13 10 9 2
14 3 16 3 3 9 9 0 13 2 0 10 9 13 2
19 16 3 9 9 3 10 0 15 9 0 7 9 13 2 0 10 9 13 2
27 10 3 3 9 0 0 9 13 13 1 9 2 3 0 10 9 13 15 2 7 0 9 0 10 9 13 2
9 13 3 3 15 7 9 0 9 2
6 3 3 0 15 13 2
17 15 3 10 9 9 1 10 9 13 2 3 10 9 13 15 13 2
16 10 3 9 15 2 16 0 9 13 2 13 1 0 9 15 2
7 9 3 3 13 7 13 2
10 9 3 3 13 9 2 16 3 13 2
21 9 3 15 10 9 13 10 3 9 13 7 9 13 1 10 9 3 15 0 13 2
8 13 3 9 13 1 9 9 2
21 10 16 15 13 0 13 2 15 3 7 10 0 2 10 9 10 9 9 0 13 2
5 3 15 15 13 2
22 15 10 1 9 9 0 3 13 9 9 7 9 13 0 2 9 13 15 9 13 9 2
6 9 3 3 9 13 2
56 9 3 2 16 1 10 9 9 13 10 9 10 9 2 13 7 13 0 1 0 9 13 2 13 7 7 13 1 10 9 13 1 10 9 10 3 9 3 10 9 3 10 9 7 10 9 2 7 3 13 10 9 0 0 13 2
14 15 3 13 7 13 9 0 2 13 13 0 9 13 2
17 10 3 3 9 13 9 13 10 0 2 1 12 9 2 13 9 2
12 10 3 12 9 0 13 3 13 7 3 13 2
16 10 3 3 9 3 13 10 9 2 3 7 3 10 9 13 2
10 3 3 10 9 10 9 13 10 0 2
24 10 3 3 3 10 9 9 0 13 2 10 7 3 15 0 9 2 0 9 13 7 15 13 2
7 10 3 3 15 0 13 2
14 15 3 15 13 3 9 0 7 0 13 2 15 13 2
12 9 16 10 0 10 9 0 13 2 9 13 2
36 10 3 9 13 3 3 3 0 9 0 0 2 10 7 0 7 0 3 3 15 9 0 13 10 9 13 2 13 9 2 13 0 3 0 9 2
17 13 1 9 0 2 9 13 9 0 12 7 12 9 2 13 0 2
29 9 3 0 15 0 3 7 0 7 0 9 13 2 3 7 9 12 3 9 0 13 10 9 2 9 7 0 9 2
12 10 3 0 9 10 0 13 9 0 12 9 2
23 13 3 15 1 15 3 13 3 3 1 10 9 10 9 13 2 7 10 9 0 9 13 2
22 13 3 10 9 13 10 9 10 1 10 9 13 2 13 7 9 0 13 15 1 9 2
15 3 3 10 9 1 10 0 9 0 13 2 13 1 15 2
9 10 0 3 10 9 13 0 9 2
18 9 3 13 1 10 9 12 2 0 0 2 7 9 3 7 9 3 2
11 13 3 0 9 13 12 9 9 1 9 2
4 9 9 15 2
6 3 13 9 3 0 2
7 9 3 10 9 10 9 2
10 13 3 15 1 10 9 9 10 9 2
15 13 3 3 10 9 9 0 2 13 7 12 9 10 9 2
12 10 3 0 15 9 13 2 15 9 13 9 2
12 13 3 1 9 2 13 0 3 0 7 0 2
8 13 3 15 1 10 9 9 2
12 10 3 3 9 0 10 9 1 10 9 13 2
13 13 3 3 15 0 13 3 15 1 0 10 9 2
25 0 3 3 10 9 9 13 2 0 7 3 9 13 2 3 0 0 0 10 0 9 2 0 7 2
43 1 3 9 0 10 9 13 1 0 1 10 3 10 9 0 0 3 7 0 2 1 7 10 0 9 9 9 0 2 3 1 15 3 15 13 2 12 9 3 2 13 0 2
37 1 0 3 10 0 9 0 13 2 9 3 10 9 7 10 9 2 3 1 0 10 9 0 9 13 2 7 0 3 1 15 2 1 15 12 13 2
13 9 3 1 15 3 9 1 0 10 9 13 13 2
19 13 3 3 10 9 13 9 3 7 9 0 2 1 15 13 13 10 13 2
9 1 3 10 0 9 9 13 0 2
16 1 3 10 9 9 0 13 3 13 2 7 15 9 13 0 2
38 9 3 3 3 0 3 13 2 7 9 15 13 9 16 3 9 0 10 0 2 15 3 10 9 13 1 0 2 16 13 10 9 13 9 0 10 9 2
42 13 3 10 0 15 2 15 3 3 0 13 2 10 9 0 13 3 1 10 9 7 13 1 10 9 2 3 3 1 9 10 9 1 10 0 9 2 16 13 10 9 2
23 3 3 3 3 13 1 10 10 9 10 9 9 2 0 7 15 13 9 0 1 9 13 2
12 3 16 13 10 9 2 9 0 0 13 15 2
23 1 3 10 9 9 13 0 2 13 7 3 0 9 0 2 1 15 13 10 0 10 9 2
36 1 3 10 0 9 3 13 13 16 3 0 0 2 1 7 10 0 9 3 13 9 0 9 9 0 10 9 3 16 10 9 13 10 9 0 2
15 15 3 15 3 13 2 15 7 13 1 9 2 15 13 2
27 0 10 9 9 3 10 9 13 3 13 13 2 9 7 10 9 13 7 10 9 13 13 3 13 10 9 2
15 10 3 3 9 0 3 13 2 13 7 3 0 9 0 2
36 10 3 9 0 0 3 3 7 0 13 9 2 15 1 10 0 9 9 13 2 15 10 9 3 13 7 10 9 2 3 7 3 3 9 12 2
27 10 3 0 13 2 10 0 9 12 0 13 2 15 9 13 9 2 15 3 13 9 1 10 9 13 0 2
11 0 3 13 10 9 1 10 9 0 13 2
59 10 3 3 0 13 15 9 2 15 9 13 9 2 0 7 0 13 10 0 13 15 3 9 13 15 15 13 2 15 7 10 9 13 9 0 3 7 3 13 2 7 0 3 13 9 15 2 3 3 3 7 10 9 2 13 0 13 3 2
40 0 3 10 9 9 13 0 0 2 15 15 1 10 9 0 13 2 15 3 9 13 3 3 15 13 0 16 3 3 1 10 15 9 10 1 10 9 13 13 2
14 10 3 9 9 13 2 1 15 13 10 9 2 9 2
29 7 3 10 16 13 1 0 10 9 1 9 2 13 10 9 9 3 3 1 10 0 0 9 13 7 1 12 9 2
24 15 3 3 0 13 2 9 7 13 1 0 10 9 10 9 0 9 9 7 9 0 15 13 2
35 3 3 0 9 13 9 9 2 0 15 13 1 10 9 2 9 3 1 10 9 3 13 2 9 7 10 0 15 13 12 3 7 0 9 2
16 10 3 13 9 1 0 10 9 13 1 10 9 10 9 13 2
13 16 3 10 13 2 9 13 9 9 1 15 13 2
29 1 15 3 13 10 9 15 10 3 9 13 7 10 0 10 1 9 9 2 16 3 13 10 9 13 15 10 9 2
14 15 3 3 1 9 13 2 0 7 1 15 9 13 2
41 10 9 13 12 9 2 10 7 9 0 13 2 1 10 0 9 16 15 13 1 10 0 9 1 0 13 2 13 9 13 2 7 13 2 16 15 13 2 0 15 2
6 15 3 3 15 13 2
17 16 3 13 10 9 10 9 2 9 0 0 1 10 3 9 13 2
91 13 9 0 2 16 7 10 13 10 9 0 7 10 9 13 2 13 10 9 10 9 0 1 15 13 9 2 1 15 13 15 2 1 15 13 10 0 9 15 3 10 9 10 9 1 10 9 7 10 9 10 1 10 9 1 10 9 13 13 9 0 1 10 0 9 10 9 2 15 7 1 0 3 3 10 9 10 9 15 13 13 9 2 13 10 9 9 3 7 9 2
11 10 3 0 0 9 3 9 0 0 13 2
25 1 10 3 0 9 10 9 9 15 13 0 1 0 10 9 2 13 7 1 10 9 9 13 15 2
19 10 15 15 0 13 9 9 16 13 9 2 13 10 9 13 0 13 9 2
9 3 3 3 3 13 3 3 13 2
13 0 10 9 13 0 1 15 1 9 13 10 9 2
26 9 3 3 0 13 13 10 9 0 15 13 2 3 9 13 7 0 10 9 13 2 7 3 13 15 2
17 13 3 10 9 13 9 3 3 2 10 7 9 7 9 13 15 2
15 16 3 0 3 13 9 7 0 2 3 3 9 9 13 2
10 0 3 3 10 9 0 15 13 13 2
25 10 3 3 9 1 0 10 9 10 9 13 2 13 3 10 9 10 15 9 9 7 10 9 9 2
39 13 3 3 9 10 0 3 9 3 13 1 9 7 9 2 7 3 3 9 1 10 9 9 3 13 10 1 9 13 2 15 0 13 9 7 0 0 9 2
23 0 3 10 9 10 9 13 0 3 9 0 0 13 1 9 0 13 2 3 3 13 3 2
83 16 3 10 9 13 1 10 9 13 1 9 9 2 15 10 3 9 1 9 9 2 13 3 1 9 2 13 3 1 0 9 9 2 10 7 1 9 9 13 1 10 9 9 13 2 0 3 10 9 9 16 13 13 10 9 13 0 2 3 15 10 15 0 9 10 9 1 9 13 1 10 9 13 13 2 10 7 15 13 0 13 13 2
32 3 3 3 13 10 9 10 9 15 13 2 7 15 13 3 3 15 0 13 16 10 0 3 9 15 3 10 9 3 13 13 2
40 1 3 10 9 13 10 1 9 9 13 10 9 3 2 13 3 13 0 13 9 12 7 12 1 0 10 9 10 9 13 0 9 2 13 7 10 9 13 13 2
20 16 3 9 0 13 13 3 10 9 2 3 7 10 0 0 3 3 13 13 2
28 16 3 10 9 9 13 9 1 0 7 12 9 15 13 2 7 10 0 9 13 2 3 3 13 1 10 9 2
7 10 3 9 13 13 15 2
21 16 3 13 13 3 10 9 2 13 3 10 9 7 13 10 9 13 1 10 9 2
24 16 3 13 3 0 10 9 3 13 2 7 13 15 0 9 3 13 2 13 9 9 3 0 2
26 3 15 3 9 13 10 9 0 2 9 7 9 13 2 16 9 3 13 0 0 7 15 10 9 13 2
21 3 3 3 15 15 13 13 2 7 3 15 13 15 0 15 13 2 13 3 15 2
48 13 10 9 0 1 9 10 9 2 3 1 10 9 13 2 7 3 3 10 9 13 0 2 3 13 1 10 9 10 9 2 13 10 9 2 16 0 10 9 13 13 2 13 3 1 10 9 2
16 3 3 3 13 7 1 15 13 13 15 1 10 0 10 9 2
29 13 3 1 10 9 2 15 3 10 10 9 9 13 1 3 10 9 7 1 10 9 2 13 3 10 9 0 15 2
22 10 3 9 9 13 1 10 9 13 9 2 10 0 9 0 13 13 2 13 10 9 2
28 16 3 3 13 7 13 10 9 10 1 10 9 13 2 10 3 3 13 10 9 13 1 10 9 13 3 0 2
31 13 3 3 0 10 1 10 9 9 13 7 15 1 10 9 13 10 1 10 9 10 9 13 2 13 3 15 16 1 9 2
9 3 3 1 0 15 13 10 9 2
8 3 9 3 3 3 0 13 2
20 10 3 9 10 9 0 3 3 15 13 0 15 13 2 1 7 3 3 15 2
21 9 10 0 1 9 15 3 7 10 9 13 2 1 10 9 2 9 0 0 13 2
11 3 0 10 0 9 10 9 10 0 9 2
39 3 10 9 10 9 0 2 15 10 9 9 13 2 13 0 10 9 0 0 0 2 3 9 10 9 1 9 13 10 9 0 9 3 13 0 9 9 0 2
9 13 3 0 10 9 0 12 9 2
28 9 3 0 0 3 0 9 13 16 9 10 1 10 9 9 0 2 10 15 13 0 2 10 9 13 9 13 2
9 15 3 10 13 10 9 13 13 2
19 10 3 9 10 9 13 3 0 2 7 10 13 10 9 10 9 13 15 2
34 13 3 1 10 9 13 3 10 9 7 13 10 9 2 3 16 3 1 9 0 10 9 13 1 10 9 2 7 9 3 7 9 13 2
15 10 3 0 9 0 2 16 3 10 0 2 13 1 9 2
14 13 3 9 15 0 0 0 15 15 13 9 9 13 2
17 10 3 3 0 9 3 13 9 13 2 3 9 3 9 7 9 2
28 10 3 10 9 9 3 0 13 13 16 1 0 3 10 3 13 2 16 7 0 15 15 13 2 1 0 13 2
17 10 3 9 3 10 3 9 7 10 9 10 9 13 9 3 9 2
36 1 3 9 7 9 0 0 9 9 13 2 13 9 3 13 2 3 13 16 10 3 13 1 10 0 9 3 10 13 9 13 1 9 0 13 2
10 13 3 15 9 7 1 10 9 13 2
40 10 9 9 13 10 3 15 7 9 15 9 9 13 2 15 10 9 13 10 0 10 9 2 7 13 3 15 10 9 10 9 13 7 3 13 10 9 10 9 2
15 9 3 3 13 1 10 9 10 9 16 3 3 10 9 2
18 0 3 0 9 0 15 13 10 3 1 3 0 10 9 2 13 13 2
19 10 9 15 13 10 1 10 9 13 1 10 9 2 13 0 2 0 0 2
8 3 3 9 0 13 9 0 2
24 13 3 1 3 12 9 7 12 9 0 13 2 7 10 3 3 13 10 9 10 7 3 13 2
11 13 3 3 3 0 0 10 9 7 0 2
10 10 3 0 15 3 0 9 9 13 2
14 1 0 3 9 9 0 13 2 1 7 10 0 0 2
36 16 3 13 13 1 10 9 7 13 10 9 2 9 3 10 9 7 10 9 0 3 3 13 2 10 7 9 13 1 10 9 13 1 10 9 2
17 1 10 9 3 3 3 0 3 13 13 0 9 1 9 10 9 2
14 1 3 15 3 3 1 9 13 10 9 7 1 9 2
18 16 3 10 9 13 13 3 1 10 9 2 0 9 10 0 13 9 2
8 10 3 3 9 15 13 15 2
12 13 3 10 9 9 13 2 13 0 10 9 2
8 9 3 0 13 7 9 0 2
18 1 0 3 9 13 13 3 9 3 9 3 9 3 9 7 0 15 2
10 1 3 9 3 15 9 13 13 9 2
10 15 3 3 15 9 1 10 9 13 2
10 1 9 0 3 10 9 0 13 15 2
41 16 3 10 9 13 9 0 2 15 16 13 0 2 1 0 9 13 0 2 1 3 15 13 9 9 2 13 7 1 0 0 9 13 2 0 3 10 0 1 0 2
19 3 3 2 16 15 13 0 9 13 2 15 3 13 15 1 15 13 0 2
5 13 3 1 9 2
15 0 3 3 13 0 10 9 0 2 13 15 13 10 13 2
25 0 3 10 9 13 0 2 15 3 9 3 15 13 0 2 10 7 3 9 3 7 0 9 13 2
44 16 3 3 13 10 9 13 10 0 10 9 13 3 10 0 2 7 16 15 15 0 13 2 3 15 3 13 2 15 13 0 9 13 13 15 2 1 15 10 10 0 13 13 2
19 10 3 3 9 13 1 10 0 9 7 3 10 0 10 0 7 0 13 2
31 13 3 10 15 9 15 13 0 3 13 2 7 1 9 13 10 9 13 2 7 0 13 13 3 3 13 15 2 3 13 2
11 16 3 3 13 2 13 10 9 13 9 2
11 13 3 3 1 15 13 9 10 13 13 2
32 10 3 3 0 9 0 15 13 2 3 7 3 3 13 13 2 0 7 15 13 3 13 16 3 13 15 7 1 0 9 13 2
18 16 3 13 13 7 13 2 0 15 10 9 9 13 13 10 0 9 2
9 0 3 9 0 0 15 9 13 2
7 10 13 1 10 9 13 2
6 3 3 3 13 9 2
16 9 3 13 10 13 3 15 13 2 16 3 13 0 9 13 2
30 16 3 3 13 9 10 15 9 0 2 1 9 13 13 2 3 3 10 9 15 0 13 2 9 7 13 13 3 0 2
8 9 3 15 13 16 3 13 2
7 0 3 15 3 9 13 2
11 10 3 3 0 10 9 13 10 9 15 2
16 13 0 9 0 13 1 9 9 3 1 10 9 13 9 0 2
23 0 3 3 3 13 13 10 15 2 16 9 13 2 1 9 1 9 13 1 10 9 13 2
7 9 3 15 3 13 0 2
6 10 3 0 13 3 2
13 1 9 9 13 9 1 10 9 13 9 0 9 2
9 10 3 3 13 2 10 7 13 2
18 0 3 9 0 9 9 13 1 10 9 2 1 15 10 9 13 13 2
25 3 16 13 9 2 3 0 13 1 10 9 16 15 15 0 9 13 1 10 9 13 1 10 9 2
6 13 3 13 13 15 2
6 13 15 10 9 9 2
7 9 3 13 10 9 9 2
8 10 3 9 9 13 0 3 2
5 3 3 3 13 2
6 3 3 15 9 13 2
7 13 3 0 0 10 9 2
9 10 3 0 13 13 7 13 15 2
25 16 3 13 2 13 10 9 13 1 10 9 2 7 1 15 3 3 0 15 15 13 16 15 13 2
28 0 3 3 9 3 13 13 7 9 2 0 13 2 0 7 0 15 13 2 9 0 13 3 13 10 9 13 2
9 3 3 0 7 0 0 9 13 2
10 3 3 3 10 9 13 0 15 9 2
8 9 3 3 10 9 0 13 2
25 13 3 15 9 12 15 15 0 13 16 3 9 0 2 10 7 3 13 13 1 9 2 13 15 2
27 13 1 9 7 13 9 13 1 9 2 7 15 3 3 13 15 3 9 13 13 2 10 7 9 9 13 2
16 7 3 10 9 3 0 10 9 13 2 13 9 1 15 13 2
30 10 3 9 0 3 0 13 13 7 0 2 13 3 1 9 3 7 9 9 2 3 10 9 9 2 0 7 9 9 2
11 13 3 15 3 0 13 0 10 9 13 2
12 10 3 9 13 3 0 7 0 13 10 9 2
24 9 3 1 15 9 9 0 0 13 13 2 1 7 15 9 15 13 3 9 10 9 13 0 2
7 15 3 15 13 9 13 2
43 10 3 9 9 13 3 1 9 2 7 3 10 9 15 1 10 9 10 12 3 7 0 13 10 9 2 9 7 13 12 2 15 10 0 1 9 1 9 3 7 9 13 2
16 1 15 9 13 13 9 0 13 2 9 7 13 13 9 9 2
15 10 3 0 10 9 10 9 13 1 0 1 10 0 9 2
14 10 3 0 9 13 1 15 2 3 13 10 0 9 2
21 15 3 3 9 13 0 3 10 1 9 9 10 9 13 7 10 0 0 13 13 2
29 10 3 9 13 15 1 15 2 13 9 3 9 9 13 12 9 2 9 7 2 3 0 13 15 15 2 12 9 2
23 3 10 3 1 10 9 13 10 9 0 10 9 13 2 13 9 3 9 0 7 9 0 2
20 9 3 9 0 7 0 1 15 13 10 9 2 10 0 0 1 9 0 13 2
24 1 10 3 9 9 0 9 13 13 13 2 15 13 3 7 13 9 9 15 1 10 9 13 2
30 10 3 3 1 9 10 9 0 10 0 13 10 9 13 2 10 7 1 9 3 7 9 13 9 13 9 0 1 9 2
22 10 3 3 9 0 10 0 3 0 9 13 10 9 2 1 15 10 9 13 9 13 2
13 3 3 13 13 9 2 0 13 0 10 9 13 2
10 13 3 10 9 13 9 10 9 9 2
5 9 15 13 9 2
12 15 13 10 9 13 10 9 13 9 15 13 2
17 10 3 9 13 3 15 15 13 7 10 9 9 2 13 10 9 2
44 9 3 1 15 2 16 15 9 3 13 2 13 1 10 9 13 1 10 0 1 10 9 9 2 9 3 13 1 10 9 9 10 9 2 7 9 1 9 10 13 10 9 13 2
13 13 3 10 0 10 9 13 10 9 9 13 15 2
12 3 3 3 13 16 15 1 9 13 15 13 2
15 13 3 13 10 15 2 7 15 13 13 13 15 3 13 2
14 3 13 9 0 13 2 7 3 3 16 1 9 13 2
15 16 3 15 13 13 3 1 10 0 2 15 15 0 13 2
24 15 3 13 10 9 13 9 10 0 2 13 7 15 1 0 15 13 10 9 2 13 0 13 2
19 10 3 1 15 10 9 13 13 13 9 3 7 10 9 15 1 10 9 2
19 13 3 7 13 10 9 0 9 10 9 13 0 10 13 9 2 13 15 2
9 10 3 15 9 13 0 9 13 2
19 16 3 0 13 13 7 9 0 13 2 0 3 13 9 9 0 0 13 2
13 3 3 13 9 1 10 13 9 10 3 16 15 2
17 16 3 13 13 10 0 1 10 9 2 0 15 1 15 9 13 2
7 13 3 13 0 10 9 2
18 13 3 3 13 0 0 16 13 1 10 15 2 13 9 2 13 13 2
19 3 3 15 13 13 13 0 3 15 13 2 3 7 15 13 13 15 13 2
16 16 3 15 13 2 9 13 0 3 0 0 7 0 0 0 2
5 9 3 0 13 2
21 9 3 13 10 0 9 2 10 9 7 13 2 13 9 13 3 15 13 1 15 2
8 10 3 3 13 7 13 0 2
55 9 3 9 1 10 9 13 10 15 9 9 2 15 3 10 9 13 2 7 0 13 15 13 3 15 7 3 13 2 16 10 9 10 1 9 3 13 2 15 13 7 13 15 1 9 2 15 13 10 9 7 10 9 15 2
18 16 3 13 10 9 2 9 13 13 9 13 1 10 9 10 9 0 2
28 9 3 10 9 13 9 9 13 10 9 9 0 2 13 3 9 1 12 3 3 9 2 7 15 13 1 9 2
7 3 3 13 3 9 13 2
14 16 3 3 13 10 9 2 13 9 15 1 10 9 2
9 16 3 15 3 13 2 15 13 2
10 15 9 13 7 15 0 13 10 13 2
14 3 13 9 1 10 9 0 0 10 3 15 13 15 2
27 15 3 10 0 13 3 1 9 7 13 3 2 16 15 15 13 13 3 2 16 15 13 10 9 1 9 2
9 9 3 13 15 9 13 13 15 2
21 10 3 10 9 13 16 15 3 13 3 15 13 2 10 7 9 15 13 1 9 2
7 13 3 3 10 9 15 2
17 15 1 3 9 13 0 9 13 2 1 7 13 1 15 13 0 2
25 16 3 0 15 9 13 9 10 0 0 13 1 15 2 15 15 13 13 15 15 15 0 15 13 2
31 9 3 15 13 7 13 10 9 13 1 9 13 9 10 9 9 2 9 7 13 1 10 9 0 9 13 1 10 9 9 2
22 10 3 13 10 3 1 10 9 13 7 10 1 10 9 2 13 9 1 9 13 15 2
9 3 3 15 3 13 13 10 9 2
17 13 15 10 9 13 1 0 10 9 0 2 9 9 10 9 13 2
23 16 3 15 3 9 2 9 13 15 10 9 9 2 3 3 15 15 3 0 13 9 13 2
9 9 3 9 15 0 13 13 9 2
41 10 3 10 9 9 9 9 2 16 15 10 3 9 13 7 13 16 13 0 2 13 9 1 10 9 13 13 2 16 7 13 3 0 7 10 9 13 2 13 15 2
8 3 3 15 3 9 0 13 2
17 9 3 2 16 10 9 3 13 2 13 0 10 15 9 13 9 2
23 0 10 9 2 0 3 0 9 9 13 2 13 0 13 2 7 3 3 13 3 15 13 2
27 0 3 3 13 15 13 1 15 13 2 3 7 16 15 10 9 13 2 13 10 9 3 7 10 0 13 2
6 9 3 10 9 13 2
25 10 3 3 0 10 0 9 3 15 13 7 3 3 0 9 13 2 13 10 0 9 13 0 9 2
35 9 3 13 9 0 9 13 1 10 13 10 9 10 9 9 2 16 3 13 2 13 15 10 9 1 10 9 2 13 7 10 0 13 15 2
17 15 3 15 13 3 7 13 15 9 13 2 9 10 0 13 9 2
11 15 3 15 2 16 3 13 2 9 13 2
20 10 3 3 1 10 9 9 10 9 2 0 9 13 2 15 15 10 0 13 2
8 9 3 7 9 10 0 13 2
27 0 3 3 1 9 3 9 7 9 2 9 10 0 13 2 0 7 1 9 3 9 7 9 2 9 13 2
25 3 3 3 10 9 10 3 1 10 9 0 9 13 2 10 7 1 10 9 3 9 7 9 9 2
7 9 3 7 9 13 15 2
17 3 3 3 15 13 1 10 9 2 10 7 9 7 10 9 0 2
5 9 3 13 0 2
10 9 3 13 0 2 15 7 0 13 2
16 15 3 13 9 9 9 2 10 9 13 1 10 9 13 3 2
9 9 3 9 15 13 0 3 0 2
25 16 3 9 13 3 2 10 13 10 0 13 13 15 7 15 9 1 15 2 13 7 10 9 13 2
26 15 3 10 0 15 13 2 10 7 9 13 3 13 7 9 13 2 9 13 16 3 13 1 10 13 2
11 13 3 15 2 7 1 9 13 7 9 2
4 9 3 13 2
10 9 3 0 9 13 2 15 13 9 2
6 9 3 15 10 9 2
11 10 9 10 0 0 10 0 10 0 13 2
26 9 9 13 13 2 15 9 13 9 0 3 0 3 7 3 1 9 0 9 0 13 7 9 0 9 2
20 7 3 13 0 9 9 7 9 9 7 9 0 0 9 9 13 0 2 0 2
4 13 3 9 2
14 15 3 3 9 0 13 9 2 9 13 9 1 0 2
7 3 13 9 0 9 9 2
11 7 15 9 13 9 0 9 13 2 0 2
15 13 3 15 9 9 2 16 13 10 3 13 3 3 13 2
19 7 15 13 13 9 9 3 13 2 15 3 0 0 3 7 0 3 13 2
9 15 3 0 13 9 1 9 0 2
12 13 3 3 9 9 9 0 9 9 0 13 2
9 13 3 9 0 9 9 3 0 2
14 12 3 15 9 13 9 9 3 1 0 0 9 13 2
44 7 16 3 3 9 13 2 1 3 13 9 9 13 2 1 3 9 0 13 2 15 3 13 12 9 0 2 15 9 13 1 9 2 0 9 13 2 0 1 0 9 0 9 2
12 1 3 0 9 3 7 9 9 13 1 9 2
12 15 3 13 1 9 13 9 0 2 0 9 2
18 1 3 13 9 0 13 2 0 3 9 1 9 13 13 9 1 15 2
6 15 3 0 13 0 2
28 15 15 13 9 9 0 13 3 13 0 9 2 15 3 1 9 0 13 9 2 15 3 9 1 9 13 0 2
13 10 3 3 9 0 1 0 13 13 9 0 9 2
12 15 3 3 13 3 3 3 0 9 3 13 2
15 13 3 1 9 9 3 13 9 0 2 1 3 13 13 2
20 1 3 3 9 7 0 9 9 9 13 1 9 7 9 2 1 3 9 9 2
7 0 15 1 9 13 9 2
6 3 3 13 9 9 2
26 13 3 0 0 9 3 13 2 15 9 3 13 7 9 0 2 9 3 0 2 15 3 0 13 9 2
10 1 9 3 9 3 0 3 9 13 2
16 9 3 3 9 3 7 9 13 2 15 13 13 9 9 13 2
25 9 3 3 0 3 13 0 0 9 0 2 16 15 3 0 13 2 16 13 9 9 9 0 3 2
31 7 3 9 13 13 9 9 2 9 3 9 3 9 3 9 3 9 3 9 3 9 3 9 3 9 3 0 9 3 0 2
11 15 3 1 0 13 9 9 2 0 9 2
5 0 3 13 9 2
17 15 3 3 10 3 0 9 0 13 2 0 3 9 0 13 9 2
15 9 3 9 13 0 2 16 3 15 0 9 9 13 9 2
10 9 3 7 9 7 9 13 1 9 2
21 15 12 3 9 1 9 13 2 0 2 9 3 0 12 1 9 13 1 0 9 2
18 0 3 9 3 7 9 13 2 0 9 2 0 3 13 9 1 9 2
27 7 15 3 16 15 0 13 2 0 13 2 7 1 9 3 13 2 9 1 9 2 0 3 13 9 9 2
8 10 3 3 13 9 0 13 2
7 0 3 0 3 13 9 2
8 13 3 13 2 0 13 9 2
6 0 3 0 13 9 2
3 3 13 2
13 15 3 3 0 13 9 2 3 3 15 0 13 2
12 13 3 0 9 9 3 3 9 13 9 0 2
6 0 3 0 13 9 2
3 3 13 2
7 13 3 0 9 9 0 2
6 13 3 15 13 9 2
6 13 3 9 9 0 2
5 9 3 13 0 2
18 13 3 9 13 0 9 2 1 3 9 13 9 13 7 3 13 3 2
31 10 3 1 9 9 13 9 0 2 0 3 0 13 9 0 0 2 0 3 1 9 9 3 13 2 3 3 13 13 3 2
8 15 3 3 15 0 13 9 2
10 0 3 9 13 0 2 0 13 9 2
28 13 3 9 13 9 3 0 0 3 9 2 9 13 2 0 9 9 13 2 9 3 15 9 13 1 0 9 2
30 9 3 16 10 0 13 0 13 1 9 0 1 9 2 3 13 1 9 0 9 2 3 3 0 9 1 0 9 13 2
6 15 3 1 9 13 2
12 0 3 9 0 13 2 3 3 0 13 9 2
15 1 3 13 0 0 9 2 3 3 9 9 1 0 13 2
21 10 3 9 0 3 9 7 0 9 2 13 9 3 7 9 2 16 1 9 13 2
17 15 3 9 13 7 9 13 0 13 10 0 9 3 1 9 13 2
15 13 3 13 9 0 13 9 2 15 3 3 9 3 13 2
21 9 3 13 0 3 9 7 9 0 7 9 2 13 3 9 2 13 3 9 9 2
30 0 3 9 7 9 0 3 15 13 9 13 9 0 2 9 3 2 15 9 1 0 9 0 0 13 13 3 9 9 2
20 3 3 3 13 9 0 9 2 16 3 1 15 13 0 9 2 15 15 13 2
16 1 15 3 9 13 7 9 9 3 0 2 7 9 13 0 2
54 3 9 0 13 3 9 0 9 3 9 3 7 9 0 9 3 9 3 9 3 9 3 9 3 0 3 9 9 3 9 3 9 3 2 0 0 2 9 3 2 15 3 0 0 9 13 2 16 3 15 0 0 13 2
11 9 3 0 7 0 13 9 2 0 9 2
22 7 13 9 2 16 0 3 7 0 2 3 3 9 13 2 7 0 7 0 9 13 2
12 0 3 9 0 13 9 12 2 0 9 13 2
4 0 3 13 2
12 15 3 0 13 9 1 0 9 7 9 0 2
16 15 3 3 3 9 9 13 2 13 9 3 0 7 9 9 2
20 15 3 0 13 2 16 9 1 9 13 2 15 3 9 0 13 1 9 0 2
13 9 3 1 9 13 9 3 9 3 13 9 0 2
38 15 3 3 13 9 0 9 1 9 0 1 9 9 10 3 3 9 13 0 9 1 0 13 9 9 9 3 13 7 9 9 9 1 0 1 0 9 2
18 3 3 15 9 13 3 0 1 9 3 1 0 3 9 0 3 9 2
9 3 3 15 13 9 0 9 13 2
7 15 3 13 13 0 9 2
17 15 3 9 13 13 0 9 2 0 3 0 3 0 3 0 3 2
6 15 3 13 12 9 2
9 2 15 3 9 13 7 0 9 2
14 3 3 15 13 13 9 9 2 13 9 9 7 9 2
7 3 15 9 13 9 0 2
9 0 3 1 9 7 9 9 13 2
9 0 3 9 7 9 13 0 9 2
7 0 3 3 13 3 0 2
16 15 9 0 0 9 9 13 2 15 3 0 13 2 0 13 2
30 9 3 9 3 0 0 3 9 9 3 2 15 0 0 13 0 3 9 2 15 9 0 13 2 13 13 9 1 9 2
23 9 3 9 13 1 9 13 9 3 0 9 3 0 9 9 3 2 15 3 0 13 9 2
15 13 3 3 0 9 0 3 1 0 9 0 1 9 9 2
10 15 3 9 13 2 0 3 9 13 2
17 0 3 3 13 9 0 13 9 2 9 3 9 0 0 9 13 2
12 3 3 3 0 3 2 3 3 13 2 13 2
9 9 3 3 9 0 13 1 9 2
28 13 3 3 9 9 1 9 9 0 13 2 0 3 2 0 9 7 0 9 2 0 1 9 2 0 1 9 2
16 13 3 9 0 2 15 3 9 13 1 0 9 0 13 9 2
13 15 3 13 9 13 2 15 1 0 9 9 13 2
15 15 3 3 0 1 9 13 9 0 3 9 13 13 3 2
19 3 3 3 2 7 3 15 0 9 13 9 0 1 9 13 2 13 9 2
26 0 3 15 13 9 3 3 2 15 0 3 9 13 9 2 7 3 15 9 13 2 16 9 3 13 2
16 0 3 9 3 7 9 13 7 9 13 2 0 13 9 0 2
22 3 3 2 16 0 2 0 9 13 9 2 7 3 7 0 3 2 16 9 13 0 2
18 1 3 9 9 1 0 13 2 1 3 9 9 13 2 15 3 13 2
22 7 3 1 9 9 13 9 2 3 9 13 2 15 3 13 9 3 13 7 9 13 2
17 13 3 9 7 9 0 9 3 13 13 3 2 9 3 9 13 2
13 3 3 3 0 1 9 13 0 1 0 13 9 2
15 13 3 15 9 0 2 15 1 0 9 13 9 0 9 2
25 13 3 9 3 7 9 0 2 16 15 13 0 1 9 13 3 0 3 13 2 9 0 1 9 2
15 3 15 3 3 3 0 9 13 2 7 13 9 0 13 2
6 9 3 13 9 0 2
25 15 3 9 0 3 3 13 7 13 2 7 15 13 2 0 3 13 13 1 9 9 7 9 0 2
13 15 3 15 13 9 0 9 1 0 13 13 3 2
12 3 15 13 13 0 1 9 0 0 1 9 2
20 13 3 15 9 13 9 1 0 2 0 1 9 9 2 0 1 9 13 0 2
9 15 3 13 9 0 13 9 0 2
35 3 3 13 1 9 2 16 15 3 1 9 0 9 0 7 0 13 2 15 15 3 13 9 7 9 13 9 13 2 15 3 1 0 13 2
12 3 3 3 3 9 7 0 9 13 10 9 2
21 13 3 9 9 9 0 13 0 9 3 13 0 9 9 13 9 9 3 9 0 2
10 2 0 3 13 9 2 15 0 13 2
15 15 15 13 9 9 2 13 3 9 7 0 9 7 9 2
7 10 3 3 0 9 13 2
7 15 0 0 7 0 13 2
20 13 3 9 9 7 9 0 9 2 0 3 9 15 0 1 9 13 9 9 2
9 0 3 3 9 0 13 9 9 2
18 9 3 9 0 9 1 9 13 13 0 9 1 9 3 7 9 0 2
23 9 3 9 0 13 0 1 9 9 1 9 2 1 9 0 2 13 9 3 7 0 9 2
7 7 15 1 9 13 0 2
20 3 15 3 9 13 0 2 15 3 13 0 3 9 0 0 9 13 0 9 2
7 0 3 13 13 0 9 2
16 3 3 13 13 9 2 15 3 13 2 16 13 9 0 9 2
23 3 3 3 13 9 0 3 9 9 2 3 3 0 9 0 9 13 13 2 9 9 13 2
31 15 3 3 9 3 7 9 0 9 1 9 13 13 9 0 2 15 3 3 9 0 9 0 1 9 13 13 13 9 9 2
10 3 3 15 13 9 9 3 9 3 2
8 3 13 13 9 0 9 13 2
15 15 3 3 13 9 9 3 13 2 0 3 3 13 9 2
4 13 3 13 2
12 9 3 0 9 13 13 3 3 3 13 9 2
12 0 3 13 9 0 9 2 15 3 13 13 2
9 9 3 15 3 0 13 0 9 2
20 13 3 9 1 2 9 3 15 13 9 2 16 13 9 0 9 0 1 9 2
15 1 15 3 0 1 9 9 9 13 9 0 0 1 9 2
8 15 3 0 13 13 9 9 2
8 3 13 13 9 0 9 13 2
21 1 0 3 3 9 13 3 3 13 0 9 9 0 0 9 2 15 1 9 13 2
11 7 15 13 0 9 9 13 0 9 0 2
8 3 3 1 9 13 0 9 2
12 9 3 13 0 0 9 0 0 9 1 9 2
21 2 1 3 15 9 0 9 13 2 15 0 13 0 0 13 9 2 13 9 9 2
15 13 2 3 3 0 13 9 7 9 2 9 13 9 9 2
18 9 3 13 0 3 9 0 3 9 2 16 13 9 0 2 0 9 2
7 0 3 13 0 1 0 2
20 15 3 9 13 7 0 9 9 3 13 13 2 0 3 1 9 13 9 0 2
14 15 3 3 9 0 13 2 13 3 1 9 13 9 2
25 15 3 3 9 1 9 13 2 0 3 13 9 13 9 2 15 3 3 1 9 0 0 13 0 2
10 3 3 13 9 13 9 3 3 13 2
6 13 3 1 9 9 2
26 3 15 3 9 13 1 9 13 13 1 9 2 0 1 9 9 2 3 3 13 2 9 0 9 13 2
24 3 15 9 3 7 0 9 0 2 15 13 0 9 9 1 9 2 9 9 13 1 9 3 2
15 0 3 15 0 3 13 1 0 9 3 7 0 9 13 2
13 15 3 3 0 9 0 13 3 13 12 0 9 2
18 3 3 15 13 9 0 9 3 3 9 0 2 0 3 9 13 9 2
18 16 9 3 13 7 9 0 2 3 3 15 13 9 9 3 9 3 2
21 3 3 3 0 0 0 9 7 9 1 13 9 0 9 3 9 7 0 9 13 2
34 15 3 0 3 9 7 9 0 13 9 0 1 9 0 13 9 0 2 0 13 1 9 3 13 0 1 9 0 1 9 1 9 0 2
3 3 13 2
7 15 3 3 13 9 0 2
23 3 3 0 13 2 10 15 3 3 9 2 3 3 13 9 2 9 3 0 9 13 0 2
21 3 3 3 0 3 9 7 0 9 13 9 0 1 0 9 13 9 1 0 9 2
3 3 13 2
10 9 3 13 9 3 3 16 10 1 2
21 15 12 3 9 1 9 13 0 3 2 9 3 0 12 1 9 13 1 0 9 2
14 15 3 9 13 1 9 0 9 0 0 1 9 13 2
16 9 3 3 13 9 3 2 9 3 9 3 3 9 13 0 2
43 0 3 13 9 0 2 9 3 0 13 2 13 3 9 0 13 2 3 3 13 0 9 9 1 0 2 9 3 13 0 9 0 2 9 3 0 9 0 9 9 3 0 2
8 3 3 1 0 13 9 0 2
8 9 3 0 13 9 0 13 2
6 15 3 13 0 9 2
26 3 3 3 3 9 13 0 9 2 7 3 15 3 3 3 9 13 9 2 1 3 3 0 13 9 2
12 3 3 3 1 9 7 1 9 13 13 3 2
19 10 3 9 3 1 9 3 7 9 13 9 1 0 2 0 9 13 0 2
15 3 3 9 0 13 13 2 13 3 3 9 0 0 9 2
11 13 3 9 0 7 9 9 9 3 0 2
29 10 3 13 0 9 9 0 2 9 3 9 0 13 0 2 9 3 13 3 0 3 13 9 13 9 3 9 3 2
6 9 3 0 13 9 2
20 13 3 3 9 13 7 9 9 13 3 2 3 16 9 7 9 0 1 13 2
16 0 3 3 0 1 9 13 15 3 13 2 15 3 3 13 2
7 0 9 13 9 9 13 2
12 9 3 0 13 0 9 2 9 3 13 9 2
4 13 3 9 2
10 3 3 0 13 3 13 1 0 9 2
16 12 3 9 3 7 9 0 9 3 13 0 3 1 9 13 2
18 12 3 3 9 3 7 9 0 9 1 9 13 0 3 1 9 13 2
6 15 1 0 9 13 2
9 1 3 15 9 3 13 1 9 2
9 7 3 9 9 13 7 0 9 2
5 15 3 0 13 2
11 9 3 13 9 0 2 9 3 13 3 2
10 9 3 0 9 0 13 9 13 0 2
30 15 1 9 9 13 9 0 13 9 3 7 0 9 3 2 3 9 3 7 9 3 13 0 13 2 13 0 9 0 2
16 3 3 3 0 9 13 13 9 9 1 13 3 3 3 13 2
29 15 3 0 9 3 7 0 9 9 0 13 7 0 9 2 15 3 0 3 9 2 0 3 15 9 0 1 9 2
7 13 3 15 0 13 9 2
29 1 3 13 13 3 9 3 7 9 0 2 13 3 3 3 13 3 2 7 13 13 2 15 3 13 9 1 13 2
10 1 3 9 0 9 13 0 9 0 2
9 3 3 3 9 0 1 9 13 2
15 0 3 1 9 9 1 0 9 13 1 9 0 9 9 2
6 0 3 1 9 13 2
20 15 3 10 0 13 13 0 2 15 13 9 0 9 2 13 0 13 1 9 2
26 3 3 3 9 7 9 13 1 9 2 7 3 13 0 7 0 0 1 9 2 0 3 15 9 13 2
16 7 16 9 13 0 1 9 2 0 3 1 0 13 0 9 2
13 0 3 13 3 9 1 0 2 15 0 9 13 2
17 0 3 9 13 9 9 0 9 0 2 15 3 13 0 1 9 2
12 3 3 9 3 0 9 13 2 1 9 0 2
16 15 9 3 13 1 9 2 9 13 2 7 9 0 0 9 2
8 0 3 1 9 9 13 13 2
12 9 3 1 0 13 0 9 0 9 13 0 2
28 7 3 3 13 9 0 9 0 7 3 15 3 0 7 0 13 2 16 3 3 0 13 9 9 3 9 3 2
24 0 3 13 7 0 2 3 3 9 0 13 7 9 0 3 9 3 9 3 9 7 9 9 2
10 9 3 1 0 0 13 9 13 9 2
4 13 3 9 2
25 9 3 1 0 13 0 9 9 3 9 3 2 9 3 1 10 9 2 9 9 3 9 3 13 2
9 13 3 9 0 7 9 7 9 2
20 13 3 3 1 9 3 3 3 3 9 0 9 1 0 2 9 3 0 13 2
22 13 3 9 2 9 13 13 2 9 3 0 2 9 1 13 2 0 9 7 0 9 2
9 3 3 0 13 0 9 0 9 2
16 7 16 3 15 13 9 13 2 13 13 2 13 3 9 0 2
14 9 3 13 13 10 9 9 1 9 0 0 2 13 2
27 0 3 0 13 9 9 0 7 13 9 7 9 1 0 1 0 9 13 2 7 9 2 15 3 0 13 2
14 9 1 9 13 9 0 13 1 9 0 1 9 9 2
8 3 3 13 9 9 9 13 2
9 13 3 15 9 13 1 9 0 2
17 1 3 9 13 9 9 0 13 2 1 9 9 3 7 9 9 2
13 0 3 3 13 9 9 2 15 0 13 1 9 2
20 15 3 3 3 1 9 0 0 9 0 13 0 9 13 9 3 7 0 9 2
28 7 16 3 9 0 9 13 2 9 3 9 13 9 2 3 3 3 13 13 7 13 9 9 0 9 9 0 2
7 15 3 15 0 13 9 2
16 3 3 15 13 2 16 3 0 9 0 13 9 1 9 9 2
8 1 3 15 13 0 9 13 2
19 7 3 15 9 3 0 13 9 2 16 3 15 13 9 0 3 0 3 2
9 15 7 1 9 9 13 13 0 2
7 0 3 3 1 9 13 2
20 7 15 9 0 1 9 13 2 15 13 9 0 2 15 9 13 0 1 9 2
5 13 3 9 9 2
21 9 3 3 13 9 2 1 15 15 9 9 13 12 2 15 13 9 7 9 9 2
7 0 3 9 0 13 9 2
16 15 3 9 7 9 7 9 13 13 1 9 9 9 7 9 2
19 7 15 3 9 7 9 0 9 1 9 13 0 2 13 9 3 0 13 2
9 3 15 9 0 9 13 13 3 2
7 15 3 3 9 9 13 2
15 15 3 13 9 9 3 9 3 1 9 9 1 9 9 2
31 7 9 0 9 9 7 9 13 0 2 15 9 0 13 9 1 9 0 1 9 0 2 9 3 2 15 9 0 13 9 2
6 3 3 0 9 13 2
12 9 3 3 13 9 0 13 1 9 9 9 2
9 15 3 15 0 7 0 13 9 2
13 9 3 0 13 0 9 9 9 3 7 9 9 2
13 15 3 15 9 0 1 9 13 13 1 0 9 2
22 15 13 9 13 2 0 13 2 0 1 9 13 9 9 9 2 7 15 0 13 9 2
6 0 3 9 9 13 2
17 9 3 3 13 0 9 9 9 13 0 9 9 1 9 0 0 2
8 9 3 3 13 1 0 9 2
12 0 3 0 1 9 13 0 13 9 0 9 2
11 13 13 13 3 2 9 3 13 9 15 2
13 3 3 0 13 9 9 2 3 1 9 13 12 2
10 15 3 3 13 13 2 15 3 0 2
6 1 3 3 9 13 2
12 10 3 3 9 3 0 7 9 13 2 0 2
15 0 15 3 13 9 2 3 1 9 0 9 9 13 0 2
9 15 7 0 3 3 1 9 13 2
9 13 3 3 9 9 1 9 13 2
16 7 9 9 13 7 9 9 2 7 0 0 13 7 9 9 2
11 15 3 13 9 7 9 13 9 1 0 2
8 15 3 3 0 13 3 13 2
14 3 3 13 9 0 9 2 15 3 1 9 13 0 2
22 3 3 3 9 13 2 3 10 0 13 13 0 13 9 0 2 15 15 9 13 13 2
7 13 3 13 9 9 9 2
17 3 3 3 3 1 9 13 2 3 15 1 9 13 7 0 13 2
16 3 3 9 3 1 9 13 2 9 9 3 13 7 9 0 2
13 3 9 13 13 9 15 2 16 15 13 9 9 2
7 3 3 9 13 9 0 2
4 13 3 9 2
18 15 3 3 0 9 9 13 9 9 1 0 1 0 9 13 9 0 2
7 15 3 13 13 9 9 2
18 15 3 15 1 9 13 0 2 15 3 0 13 1 9 0 0 13 2
3 3 13 2
9 1 3 13 9 9 3 9 3 2
29 9 3 13 0 16 0 9 9 13 2 1 3 9 13 9 7 9 2 0 3 9 1 9 13 9 0 9 0 2
3 3 13 2
14 3 3 1 9 13 0 0 9 0 0 9 1 9 2
8 13 3 7 13 9 0 9 2
14 1 3 15 9 3 9 7 9 9 9 0 13 9 2
10 1 3 15 3 9 9 13 9 0 2
9 0 3 15 9 9 13 9 9 2
28 3 3 9 13 2 16 15 13 9 7 3 9 13 1 9 0 2 3 13 3 2 16 3 15 0 0 13 2
11 3 15 13 2 3 3 0 13 2 13 2
26 3 3 3 13 1 9 9 9 1 1 3 0 7 1 0 9 9 15 0 2 15 3 9 9 13 2
7 3 3 1 9 9 13 2
6 9 3 13 9 0 2
10 3 3 13 9 9 0 9 9 9 2
13 16 3 13 2 0 15 15 9 13 3 7 3 2
7 15 3 1 9 13 0 2
12 0 3 0 9 9 9 0 13 0 9 13 2
10 15 3 1 9 13 2 3 9 13 2
14 3 9 3 13 0 9 13 3 1 3 9 7 9 2
6 13 3 3 9 13 2
11 9 3 13 0 9 0 0 3 7 0 2
18 3 12 3 9 9 1 9 0 13 13 2 0 0 2 15 1 9 2
19 3 3 3 13 3 7 9 9 13 2 0 13 1 9 2 9 13 9 2
27 9 3 0 3 13 0 13 2 3 3 0 13 13 3 3 13 9 0 1 9 2 15 9 9 1 9 2
19 15 3 3 9 9 13 13 2 16 9 3 13 9 9 2 15 9 13 2
51 3 16 3 0 9 1 9 13 2 2 15 3 0 9 0 13 2 0 2 7 3 9 3 15 13 2 2 9 3 9 0 0 9 9 9 0 13 2 3 0 0 0 2 1 9 2 0 3 7 0 2
8 15 9 9 13 0 7 9 2
6 0 3 3 13 9 2
24 3 3 15 3 9 9 13 2 15 3 3 9 9 7 9 13 9 9 13 9 1 9 9 2
4 15 9 13 2
10 15 3 9 13 9 9 3 9 3 2
9 15 3 3 0 9 7 9 13 2
17 0 3 3 3 0 9 13 9 9 9 2 15 13 1 9 9 2
16 3 3 13 15 0 13 9 2 3 7 3 13 7 3 13 2
7 3 3 3 9 13 0 2
6 0 3 9 13 9 2
8 3 3 3 15 13 0 0 2
15 9 3 13 3 0 9 9 9 2 3 3 13 0 13 2
6 3 3 13 13 9 2
14 13 3 3 15 0 13 9 0 3 3 9 9 13 2
12 3 3 3 15 3 13 9 1 0 13 9 2
6 0 3 0 9 13 2
16 13 3 10 0 10 0 9 9 0 13 2 1 3 9 13 2
11 9 3 9 0 0 0 0 13 2 0 2
23 3 3 3 1 9 1 9 9 0 9 13 9 0 0 1 9 13 13 9 9 7 9 2
8 10 3 13 9 0 0 9 2
6 0 3 3 13 9 2
9 3 3 9 9 13 13 7 0 2
13 3 9 13 9 0 3 3 1 9 13 9 13 2
11 15 3 3 2 0 13 1 9 2 13 2
7 15 15 3 1 9 13 2
6 13 3 15 0 0 2
14 3 3 13 2 3 15 3 15 3 13 3 9 13 2
9 9 3 13 1 3 9 9 13 2
9 9 3 1 9 13 1 9 13 2
6 13 3 3 0 13 2
25 15 3 13 13 9 7 9 9 2 9 13 2 0 9 13 2 15 3 15 13 7 3 0 13 2
20 15 13 3 9 0 9 2 9 3 9 0 3 3 13 9 2 0 3 9 2
6 0 3 9 9 13 2
7 13 3 9 13 9 9 2
5 13 3 0 3 2
18 15 3 9 3 13 0 7 0 9 2 15 3 9 9 13 0 9 2
15 3 3 0 9 0 9 13 2 15 3 13 7 0 13 2
4 13 3 9 2
18 3 3 1 9 13 0 13 2 0 0 9 0 13 9 9 3 13 2
13 3 3 0 13 1 9 0 0 9 9 0 9 2
16 15 3 13 3 9 7 0 9 9 13 2 3 13 1 9 2
20 10 3 3 9 13 9 2 9 13 2 0 3 0 3 9 2 15 9 13 2
18 15 3 0 0 13 9 0 0 13 2 10 3 0 9 10 13 0 2
31 0 13 9 9 7 0 13 3 3 15 2 16 3 13 2 13 2 3 3 15 13 2 0 3 3 15 9 9 3 13 2
13 3 3 15 3 0 1 9 0 13 3 0 9 2
10 3 15 3 3 3 13 13 9 0 2
10 9 3 13 9 2 15 0 0 13 2
18 16 3 15 3 13 10 0 13 13 2 15 3 3 9 13 0 9 2
24 15 3 3 9 0 0 13 13 2 1 3 9 13 0 13 2 15 3 15 0 9 3 13 2
10 10 3 3 9 3 3 13 13 3 2
9 0 3 9 2 3 3 3 13 2
9 10 3 9 9 9 1 13 0 2
15 3 3 1 9 13 2 0 3 3 13 2 0 3 13 2
25 15 3 9 13 7 9 2 15 3 0 13 2 9 0 0 9 2 15 3 9 9 13 0 13 2
16 0 3 9 0 13 0 13 2 16 3 15 0 9 13 9 2
11 16 3 3 13 2 3 15 13 0 13 2
7 9 3 9 7 9 13 2
9 3 15 15 3 3 13 0 9 2
36 3 3 9 9 3 13 2 7 3 13 7 3 3 9 0 13 2 16 3 15 0 9 7 9 13 2 16 0 13 9 2 3 10 0 0 2
11 10 13 1 9 13 2 10 3 0 13 2
11 15 3 3 13 2 15 15 15 1 13 2
17 16 3 15 3 9 0 0 13 2 9 0 13 2 13 3 9 2
10 13 3 9 2 15 3 13 9 0 2
12 3 3 3 9 13 2 16 3 9 0 13 2
30 3 3 13 1 9 2 3 3 13 2 0 10 9 2 7 0 2 16 3 13 2 16 3 13 3 1 0 0 13 2
4 3 0 13 2
9 10 13 13 2 7 10 13 13 2
16 7 13 2 15 3 13 2 7 3 13 2 15 3 3 13 2
10 9 3 15 13 2 9 3 0 13 2
23 15 3 3 3 9 13 2 15 3 2 16 0 13 2 13 10 9 7 13 0 1 9 2
12 15 3 1 13 13 2 15 3 13 0 9 2
20 16 3 3 3 0 1 0 13 7 3 0 13 2 3 3 0 3 15 13 2
10 3 3 10 3 1 9 13 9 13 2
8 9 3 9 0 13 0 13 2
8 3 3 9 13 1 9 13 2
9 9 3 3 3 7 9 13 9 2
14 3 3 9 15 9 0 13 0 13 2 0 13 9 2
10 15 3 9 13 2 13 15 3 9 2
14 0 3 9 13 0 9 13 3 3 9 13 1 9 2
7 0 3 13 0 9 13 2
9 3 3 3 0 13 9 0 9 2
10 9 0 13 13 9 2 9 3 13 2
20 15 3 3 9 3 7 9 12 13 2 3 3 13 9 13 10 0 13 9 2
20 0 13 2 0 3 13 2 0 3 13 2 16 3 0 0 13 9 13 9 2
18 3 3 0 0 13 2 16 3 10 3 13 13 0 9 7 9 13 2
7 3 3 3 1 15 13 2
8 3 3 3 7 3 3 13 2
6 0 3 13 9 9 2
11 3 15 13 13 9 3 9 9 3 9 2
10 3 3 13 1 3 3 1 3 0 2
10 3 3 0 9 13 9 3 3 13 2
6 9 3 10 9 13 2
7 3 3 0 9 9 13 2
19 3 3 3 9 9 0 1 9 0 9 13 0 2 0 3 3 9 13 2
16 3 0 13 13 9 9 2 9 3 3 13 2 9 3 13 2
7 3 3 13 13 0 9 2
13 9 3 0 13 2 9 3 0 2 9 3 0 2
11 16 3 3 9 2 1 3 9 3 13 2
7 0 3 9 13 0 9 2
20 13 3 9 2 3 3 13 2 1 9 2 1 9 13 7 1 9 2 0 2
19 15 3 9 13 0 13 2 3 3 9 9 1 9 13 9 13 13 9 2
18 0 3 13 9 2 13 1 9 2 0 7 0 2 16 0 0 3 2
11 16 3 0 13 2 0 3 1 9 13 2
16 9 3 0 0 13 2 15 3 9 3 0 2 9 9 13 2
19 3 3 15 3 13 1 9 1 3 9 13 2 10 3 9 0 3 13 2
31 15 3 3 0 0 13 9 13 0 2 0 2 15 9 13 0 3 9 13 2 3 13 1 9 2 7 1 9 9 13 2
7 0 3 9 1 9 13 2
14 13 3 2 3 3 9 9 13 3 1 9 0 13 2
11 15 9 3 9 13 7 9 9 13 0 2
6 9 3 13 9 0 2
8 3 3 13 0 9 3 13 2
5 9 13 7 9 2
4 13 9 9 2
15 13 3 9 9 0 13 9 2 0 2 3 3 15 13 2
33 3 3 3 0 9 0 13 2 3 3 13 3 9 3 7 0 0 7 0 13 9 1 9 2 3 3 13 2 16 15 13 9 2
3 9 13 2
7 9 3 13 3 15 13 2
7 9 3 13 3 13 9 2
34 13 3 9 0 9 3 0 2 0 13 9 0 9 2 13 10 0 9 2 3 3 9 9 9 13 9 9 1 9 13 9 13 9 2
13 10 3 0 3 9 13 9 9 9 13 9 13 2
21 3 3 9 9 13 3 2 16 9 0 3 0 0 13 2 1 3 9 13 9 2
9 7 15 13 13 9 13 3 13 2
12 13 3 13 0 9 2 3 3 1 0 13 2
7 15 3 0 9 13 13 2
29 16 3 3 9 9 13 9 0 2 13 13 0 1 9 13 2 0 13 13 2 3 3 13 2 13 3 1 9 2
5 0 3 15 13 2
12 16 3 3 3 13 2 15 3 15 9 13 2
6 3 3 9 9 13 2
7 1 9 3 3 0 13 2
12 3 3 15 13 3 9 13 0 3 0 9 2
17 0 3 0 9 2 0 1 9 13 2 13 9 2 0 13 9 2
17 9 3 3 0 13 9 13 2 13 1 9 2 15 9 0 13 2
8 13 3 9 9 3 0 13 2
8 3 3 9 13 2 13 9 2
6 13 3 9 7 9 2
22 0 3 9 0 9 3 0 9 1 9 13 9 0 13 2 7 0 13 3 0 9 2
16 9 3 13 2 9 3 1 9 13 2 15 3 9 9 0 2
11 3 3 3 15 0 13 13 0 3 13 2
12 3 3 1 9 9 13 2 3 3 15 13 2
7 3 3 1 9 13 0 2
16 9 3 3 15 2 16 0 9 0 2 3 13 9 9 9 2
5 0 3 9 13 2
21 7 1 9 0 3 13 2 15 9 1 0 1 9 13 3 3 9 13 0 9 2
29 3 3 13 0 9 7 3 9 13 0 13 1 9 9 0 2 3 0 0 9 13 1 3 0 9 7 9 0 2
8 3 3 15 9 13 9 13 2
15 3 1 0 9 9 3 9 3 13 2 0 3 9 13 2
14 7 3 3 0 7 0 9 0 13 1 9 0 13 2
26 3 3 0 9 0 2 15 3 1 9 13 2 9 3 1 9 13 2 15 0 13 2 13 9 0 2
17 7 3 13 9 9 2 3 15 13 2 9 3 0 7 0 9 2
8 9 3 1 0 0 9 13 2
16 15 13 2 16 15 9 13 2 3 3 0 13 13 1 9 2
14 1 3 9 9 9 3 13 13 13 2 9 3 13 2
22 0 3 9 2 3 3 9 0 13 2 9 13 9 9 2 16 1 9 9 13 9 2
12 9 3 3 9 13 0 2 16 9 3 13 2
21 0 3 3 9 13 9 13 0 3 1 9 1 9 0 9 0 13 9 1 9 2
27 15 13 9 1 0 2 3 1 9 13 9 9 3 3 3 13 1 0 2 3 13 0 0 9 9 13 2
24 15 13 9 13 3 13 2 16 3 15 3 0 9 13 2 9 3 0 13 1 3 9 13 2
3 3 13 2
11 3 0 9 2 1 9 3 0 13 9 2
6 0 3 0 9 13 2
20 0 13 13 1 9 13 9 3 7 9 2 3 3 9 0 9 9 0 13 2
26 3 3 3 12 1 9 9 0 13 9 9 2 3 3 3 9 9 13 0 9 9 0 13 13 0 2
15 15 3 1 0 9 13 9 1 9 9 2 9 0 13 2
5 15 13 9 13 2
8 3 9 3 13 7 9 13 2
18 13 3 0 9 7 1 9 9 9 1 9 2 3 3 9 9 13 2
15 3 13 7 3 9 13 9 13 2 16 15 9 0 13 2
30 3 3 3 13 0 3 9 7 9 9 2 9 3 0 9 3 9 13 2 7 9 0 9 3 3 13 0 3 9 2
39 1 3 0 13 9 2 1 9 13 2 13 9 9 2 0 0 9 13 9 2 9 3 0 7 0 2 15 0 2 3 9 13 2 10 3 0 13 9 2
23 9 3 13 9 0 9 13 2 3 3 0 13 9 9 2 9 1 0 7 0 1 9 2
7 9 3 3 13 1 9 2
18 7 9 0 13 2 3 13 9 2 16 3 15 0 9 1 9 13 2
14 9 3 13 7 9 2 16 15 13 9 7 9 0 2
10 3 3 9 13 0 9 7 9 13 2
23 13 3 9 12 3 9 7 12 9 2 12 3 13 2 0 3 1 9 13 9 9 0 2
20 3 16 3 9 3 9 3 10 3 9 9 13 2 3 3 9 13 13 0 2
7 9 3 1 9 13 13 2
27 16 3 15 9 0 9 13 2 3 3 9 9 0 9 13 13 1 0 9 2 3 3 0 9 13 9 2
17 7 3 3 9 13 1 0 9 2 9 13 13 2 3 15 13 2
26 9 3 1 9 13 13 3 9 3 2 16 13 9 9 0 13 2 9 13 2 16 3 13 9 9 2
13 9 3 13 0 0 13 9 3 13 9 9 0 2
7 9 3 0 1 9 13 2
9 0 3 0 13 9 2 3 13 2
19 15 3 3 3 13 2 0 1 9 13 2 9 0 13 2 1 9 0 2
10 9 0 13 2 0 3 1 9 13 2
19 0 3 9 2 0 3 1 9 9 13 2 16 3 9 3 0 13 9 2
32 3 3 1 9 13 0 9 13 9 3 13 7 9 0 2 13 3 15 9 0 9 2 3 3 15 9 13 3 3 15 9 2
33 3 3 3 3 9 3 13 0 9 2 16 3 1 9 1 9 2 15 3 0 13 9 0 1 9 13 9 1 0 9 1 0 2
12 3 3 15 1 9 0 9 9 3 1 13 2
9 10 3 13 0 9 13 9 9 2
9 3 15 13 9 13 13 9 0 2
15 15 3 15 9 9 13 2 3 15 10 0 0 13 9 2
7 0 3 9 3 13 0 2
8 3 3 3 13 9 9 0 2
8 9 3 15 13 0 9 13 2
18 9 12 1 9 9 2 1 9 13 9 0 9 2 0 13 0 9 2
25 3 3 3 9 13 3 3 9 13 9 2 16 3 3 0 3 9 9 7 9 0 9 13 13 2
11 1 15 3 9 13 3 0 3 0 3 2
23 0 3 9 0 9 13 13 1 9 9 3 1 0 13 2 13 3 7 0 3 3 13 2
32 3 3 13 9 3 0 7 0 9 7 9 13 9 3 0 9 2 15 13 9 13 9 9 0 0 2 0 3 3 9 13 2
7 0 3 0 13 9 9 2
26 3 3 10 0 2 0 3 13 9 9 13 2 0 9 9 13 1 9 0 2 3 3 0 13 9 2
6 0 3 0 13 9 2
5 3 15 15 13 2
7 3 3 0 9 13 13 2
5 3 3 13 0 2
9 3 3 3 15 9 13 9 9 2
7 9 3 9 13 0 9 2
7 0 3 13 13 1 9 2
9 3 3 1 9 0 9 0 13 2
9 3 0 13 2 10 3 0 13 2
3 9 13 2
19 0 3 9 0 1 9 13 2 3 12 9 3 0 13 3 13 3 0 2
10 10 3 9 0 13 2 0 3 13 2
10 9 3 13 2 16 3 9 0 13 2
20 15 3 3 13 2 15 15 15 3 13 2 0 3 13 2 16 9 9 13 2
21 3 3 3 15 9 9 13 0 10 0 2 10 3 3 0 3 0 0 2 0 2
14 15 9 3 0 3 13 13 1 9 7 0 9 13 2
8 3 3 9 0 9 13 13 2
7 3 3 9 0 13 9 2
11 16 3 3 13 2 3 15 0 0 13 2
6 3 3 13 9 9 2
19 16 3 15 3 13 7 15 9 13 0 7 3 13 2 3 0 13 13 2
16 16 3 15 3 3 13 1 9 2 9 3 13 13 2 13 2
16 0 3 9 0 3 0 13 2 15 3 3 15 9 13 9 2
17 3 3 0 3 3 0 13 2 3 3 0 9 3 3 0 9 2
11 16 3 0 13 2 3 3 0 0 13 2
9 3 3 0 9 0 13 1 0 2
16 3 3 3 1 9 9 13 0 9 9 0 3 3 0 0 2
11 3 3 15 3 13 2 13 3 3 9 2
8 3 3 1 9 13 0 13 2
12 3 1 9 3 1 9 3 13 3 3 13 2
5 9 3 9 13 2
14 3 3 9 9 13 1 9 9 1 13 2 7 13 2
14 3 3 1 0 9 13 13 9 2 7 0 1 9 2
17 15 9 13 9 7 9 0 2 15 3 9 13 7 9 13 3 2
15 3 3 1 0 9 1 9 0 0 1 0 13 0 9 2
9 3 3 3 9 13 9 1 13 2
7 0 3 1 0 9 13 2
14 3 3 9 13 0 13 2 16 3 13 13 9 9 2
11 3 3 1 9 0 13 13 3 3 13 2
22 3 3 1 0 13 2 3 3 0 2 9 0 2 16 9 0 13 2 3 3 0 2
5 0 3 0 13 2
8 3 3 0 9 9 13 9 2
10 0 3 1 9 13 1 3 15 9 2
9 3 3 9 1 13 13 13 0 2
7 9 3 15 3 15 13 2
18 3 3 3 1 9 9 3 13 3 3 1 9 13 2 3 3 13 2
4 3 3 13 2
7 15 3 3 3 0 13 2
3 3 13 2
6 0 3 9 13 9 2
20 9 3 3 0 13 2 0 3 13 3 3 2 0 3 13 2 0 3 13 2
12 9 3 0 3 13 2 15 15 0 9 13 2
7 9 3 15 13 3 0 2
11 9 3 1 3 13 3 1 9 13 9 2
15 15 3 9 13 9 1 0 2 3 3 9 9 13 13 2
7 15 3 9 0 13 9 2
16 15 3 3 13 9 0 9 9 1 0 2 3 0 9 13 2
9 15 3 9 13 9 13 3 9 2
8 9 3 13 0 13 9 13 2
13 9 3 10 0 3 0 13 9 2 0 3 0 2
16 9 3 3 0 13 2 3 3 13 0 3 3 3 9 13 2
15 13 3 15 3 0 13 9 3 0 3 9 0 3 9 2
14 9 3 0 9 7 9 0 13 2 9 3 0 0 2
7 3 3 3 9 13 13 2
19 15 3 3 9 7 0 0 9 7 9 0 7 9 0 13 1 9 13 2
17 13 3 9 9 13 13 3 13 3 9 15 13 3 3 13 9 2
16 1 3 0 9 13 9 9 9 13 2 15 1 9 0 0 2
10 0 3 13 2 16 0 3 7 0 2
15 1 0 3 13 9 13 9 13 2 15 9 13 9 0 2
30 0 3 0 9 0 9 3 3 13 0 1 9 13 2 0 3 13 0 9 0 3 9 0 2 15 3 13 9 13 2
7 9 3 13 9 13 0 2
30 0 3 3 13 9 9 0 13 3 9 7 1 9 9 13 9 7 9 7 9 0 2 9 0 0 1 0 9 13 2
6 0 3 3 0 13 2
5 9 3 13 9 2
6 1 0 3 13 0 2
19 15 3 9 13 0 0 9 2 10 3 0 0 2 0 2 3 15 13 2
9 0 3 0 13 2 0 3 13 2
8 3 9 13 9 2 3 9 2
11 15 3 9 9 13 0 9 3 9 3 2
14 9 3 3 3 15 13 15 2 15 0 0 13 13 2
18 15 3 3 3 1 9 0 13 9 2 7 3 3 15 13 9 0 2
13 3 3 15 9 0 13 3 13 2 13 1 9 2
12 13 3 15 3 0 9 1 9 13 0 0 2
11 3 3 15 13 2 9 3 1 9 13 2
20 15 15 3 13 9 2 13 3 16 0 13 0 9 2 15 15 3 9 13 2
9 13 3 15 0 9 9 13 9 2
22 9 3 9 3 9 3 0 9 13 1 9 2 16 3 9 9 3 9 9 9 13 2
15 13 3 1 9 9 9 13 2 13 9 0 9 2 0 2
5 3 3 13 9 2
8 3 3 9 0 13 9 9 2
7 3 13 9 13 0 9 2
16 0 3 3 9 0 9 9 7 9 13 2 13 3 3 9 2
19 3 3 15 3 1 9 7 9 9 13 13 2 16 3 0 9 13 9 2
31 3 3 7 9 0 13 9 9 1 0 7 3 0 1 9 2 3 3 3 9 0 9 13 3 3 3 3 0 9 13 2
12 0 3 3 13 1 0 9 13 9 0 9 2
20 15 3 9 13 7 9 0 0 9 1 0 9 13 9 2 3 1 0 13 2
5 9 3 3 13 2
20 9 3 13 0 9 13 9 2 9 3 15 13 13 0 1 9 7 9 9 2
9 9 3 0 7 9 13 9 13 2
19 13 3 9 0 2 13 9 9 0 9 3 9 13 7 1 0 9 13 2
8 7 15 9 3 13 9 9 2
16 0 3 9 7 9 9 9 13 1 0 9 9 3 7 0 2
6 9 3 3 9 13 2
15 15 3 0 13 0 13 3 13 1 3 9 7 0 9 2
15 0 3 0 3 9 7 9 0 1 9 13 1 0 9 2
28 13 3 1 9 7 9 0 2 15 3 15 13 7 9 0 13 2 15 9 13 9 2 13 3 15 3 3 2
22 15 3 9 13 9 2 15 13 0 3 9 0 3 9 13 2 13 13 9 2 0 2
9 3 3 0 13 3 0 9 13 2
6 15 3 3 0 13 2
7 7 15 9 0 13 9 2
9 3 3 3 0 3 13 13 9 2
7 15 3 3 13 0 9 2
19 0 3 3 15 9 0 3 0 3 0 1 9 13 2 16 9 0 13 2
53 3 3 13 9 0 2 16 0 9 13 9 3 0 3 13 2 16 3 3 0 9 9 3 3 9 13 2 7 15 13 13 12 9 0 9 2 15 3 15 3 13 2 13 9 9 13 2 15 15 0 0 9 2
3 3 13 2
7 13 3 9 0 9 13 2
7 7 15 13 9 0 13 2
8 0 3 1 9 9 13 3 2
30 13 3 0 9 2 0 9 9 2 9 3 1 0 9 0 13 2 0 0 2 1 9 13 2 15 13 9 9 0 2
23 0 3 3 9 9 0 3 9 9 3 0 13 9 3 0 13 2 9 3 1 9 13 2
16 1 0 3 0 13 9 3 15 0 2 3 9 9 13 13 2
35 15 7 9 3 13 9 0 13 2 0 0 2 1 3 0 9 0 9 13 13 9 9 2 0 2 15 3 9 3 7 1 9 13 9 2
7 15 3 9 9 9 13 2
22 15 7 9 3 9 13 9 1 13 2 9 3 15 1 9 13 9 0 0 13 9 2
46 1 3 9 3 9 3 13 2 1 3 9 3 9 3 9 3 13 2 1 3 9 2 1 3 9 13 2 1 3 0 9 0 0 13 0 2 0 0 2 0 13 1 9 13 9 2
15 9 3 13 1 9 0 9 9 2 0 13 9 3 13 2
28 1 3 9 9 0 13 2 3 15 0 2 12 2 15 13 1 9 9 9 2 15 15 3 9 9 9 13 2
17 10 7 9 3 9 13 2 7 13 9 2 10 3 13 0 9 2
8 9 3 3 13 13 0 9 2
8 0 1 9 2 13 3 9 2
12 13 7 9 1 15 13 2 13 3 13 3 2
6 15 7 3 9 13 2
8 3 3 3 15 3 0 13 2
6 13 3 3 9 0 2
23 3 3 15 13 0 9 2 1 3 9 0 2 13 9 2 1 3 15 0 9 13 3 2
10 15 3 9 13 13 13 1 0 9 2
14 7 3 3 3 16 0 3 13 9 7 9 3 13 2
12 1 3 9 3 9 3 13 13 9 13 9 2
6 1 3 13 9 0 2
7 1 3 13 0 0 9 2
13 1 3 3 0 0 13 9 7 9 9 0 9 2
13 1 3 9 0 0 9 0 13 0 9 13 0 2
15 0 3 3 1 0 0 9 3 7 3 13 13 13 0 2
7 15 3 1 0 13 9 2
8 7 1 9 13 9 9 13 2
8 13 3 9 9 9 13 13 2
9 3 3 15 9 13 0 0 0 2
7 1 3 9 13 0 9 2
11 9 3 15 1 0 9 13 0 1 9 2
7 15 3 7 3 9 13 2
6 9 3 13 0 0 2
13 0 3 1 9 9 13 9 9 9 9 0 13 2
10 0 3 13 7 13 13 9 9 13 2
14 15 3 1 0 9 0 3 7 3 0 13 13 13 2
13 1 3 0 0 13 13 9 0 9 0 7 3 2
9 1 3 9 9 0 13 13 9 2
6 13 3 3 15 3 2
7 9 3 13 9 0 13 2
9 1 3 0 9 0 13 0 9 2
26 15 3 1 0 9 13 0 9 13 2 15 3 1 0 9 0 3 9 9 13 2 15 3 13 13 2
11 0 3 13 2 0 3 3 9 13 13 2
22 10 3 9 0 1 9 0 0 13 2 1 3 13 9 2 0 0 2 9 0 9 2
27 9 3 2 15 9 13 9 3 13 2 0 1 9 13 2 1 3 9 9 13 9 2 1 0 9 13 2
6 15 3 3 9 13 2
23 10 3 1 0 9 0 2 0 13 9 2 0 0 3 0 3 0 3 9 13 1 13 2
8 0 3 3 13 9 0 13 2
24 15 3 0 13 13 7 13 0 2 1 3 0 13 9 0 2 9 3 3 13 9 1 0 2
22 15 3 9 16 13 9 0 2 15 3 13 3 2 3 3 9 7 9 13 3 13 2
6 9 7 9 15 13 2
24 10 3 0 9 3 15 13 0 9 2 7 3 15 3 10 3 3 0 0 3 13 0 3 2
9 0 3 1 9 9 9 0 13 2
16 0 3 1 0 13 9 13 2 3 3 9 9 3 0 13 2
22 1 3 9 13 0 3 7 0 2 0 0 9 13 2 0 2 0 3 9 9 13 2
14 15 1 3 9 9 13 2 1 3 9 9 13 3 2
15 15 3 0 13 13 2 0 3 9 13 9 2 9 0 2
9 0 3 15 13 9 13 12 9 2
11 10 3 9 1 9 3 9 3 9 13 2
15 15 3 3 0 1 9 13 9 9 2 0 3 9 13 2
11 3 3 1 13 9 9 13 9 1 9 2
7 15 3 9 13 3 13 2
6 15 3 9 13 13 2
17 15 3 1 0 9 13 9 1 0 9 2 1 3 15 13 9 2
8 15 3 1 9 13 9 0 2
29 3 3 3 3 0 13 1 9 2 15 3 3 3 13 1 9 7 9 15 3 3 3 13 1 9 0 3 13 2
11 0 3 9 9 3 9 3 9 3 13 2
10 15 3 3 1 9 9 9 13 13 2
12 10 3 9 13 9 0 2 3 3 9 13 2
5 7 13 0 9 2
41 15 3 3 1 9 13 7 13 9 2 15 3 13 9 9 1 9 13 2 15 3 3 1 9 13 1 9 0 7 0 9 0 1 9 2 13 9 7 0 9 2
7 15 3 3 1 9 13 2
5 13 3 3 15 2
9 15 3 3 13 2 15 3 13 2
8 15 3 13 3 3 7 3 2
21 15 3 9 9 13 9 9 2 7 0 9 3 2 13 13 2 15 3 13 13 2
15 1 3 0 9 13 9 2 1 3 9 9 13 7 9 2
25 0 3 1 9 9 13 13 0 9 9 13 2 10 3 13 13 9 0 2 1 3 9 0 13 2
18 15 3 3 0 13 9 3 3 3 15 9 13 2 7 0 13 9 2
32 1 3 9 13 9 13 13 2 0 3 13 9 0 2 15 3 1 0 9 9 0 13 2 15 3 3 0 13 1 0 9 2
5 3 3 9 13 2
8 15 3 9 0 9 13 3 2
15 1 3 0 13 9 2 0 9 9 9 0 2 0 13 2
17 3 3 9 9 15 13 9 13 9 3 13 7 1 0 9 13 2
38 16 3 3 9 0 9 13 2 15 3 3 3 13 7 9 15 2 0 3 0 9 13 13 2 3 3 13 9 1 0 9 13 2 3 13 0 9 2
4 3 3 13 2
17 3 13 1 9 13 0 9 2 9 0 9 7 9 13 2 3 2
9 3 3 3 0 9 0 9 13 2
11 15 3 1 9 3 13 0 9 13 9 2
4 13 3 9 2
15 15 9 3 3 0 0 0 13 2 1 3 15 13 9 2
6 15 0 13 9 0 2
11 7 3 13 9 0 7 9 13 3 13 2
8 9 3 3 13 1 9 9 2
17 15 3 9 3 7 9 9 13 2 15 3 3 3 13 3 0 2
23 3 3 3 15 13 3 3 13 9 0 2 3 1 9 0 0 13 15 2 9 0 13 2
26 3 3 0 1 9 13 13 9 13 9 2 10 3 0 13 9 0 9 13 2 1 3 0 9 13 2
9 0 3 1 9 3 13 9 9 2
14 3 3 3 0 1 0 13 9 1 0 13 9 0 2
3 3 13 2
12 3 3 3 9 9 13 15 13 13 9 9 2
17 3 3 1 0 9 13 3 1 9 9 3 9 0 7 9 9 2
7 9 3 3 13 9 9 2
9 15 3 1 13 13 9 0 9 2
46 3 3 3 1 0 9 9 0 9 13 2 1 0 3 13 2 0 3 9 0 2 0 3 3 9 9 3 0 13 1 0 3 13 2 16 3 13 2 3 15 1 0 13 0 13 2
21 0 3 9 3 9 0 3 9 9 3 7 9 9 3 0 9 1 0 0 13 2
6 15 3 9 0 13 2
6 0 3 13 9 9 2
16 1 3 3 1 3 9 13 0 2 9 13 9 0 0 9 2
9 15 0 9 9 1 0 13 9 2
9 15 9 13 2 0 3 9 13 2
7 3 15 13 1 0 13 2
20 3 3 3 9 3 0 9 9 13 13 9 13 0 9 2 3 3 13 9 2
5 13 3 9 9 2
8 1 3 0 13 9 0 9 2
6 0 3 9 13 9 2
18 13 3 2 3 3 15 9 13 7 3 9 0 2 13 9 0 9 2
3 3 13 2
8 1 3 15 13 9 0 9 2
38 15 3 3 13 9 0 9 2 0 3 0 9 13 13 2 0 13 9 2 9 3 9 13 2 15 3 3 3 9 0 9 13 3 0 9 9 13 2
10 1 9 3 3 15 3 0 13 9 2
27 13 3 9 0 9 3 7 9 9 13 9 13 2 3 3 15 0 13 1 3 13 3 13 3 3 13 2
18 0 3 9 2 0 9 2 0 13 9 2 1 9 9 13 2 3 2
8 15 3 15 1 13 13 9 2
7 0 3 13 1 0 13 2
10 0 10 3 9 0 0 9 13 13 2
5 15 3 3 13 2
8 0 3 3 13 9 0 13 2
11 3 3 13 9 2 3 3 0 13 15 2
3 3 13 2
22 7 3 13 9 0 9 2 7 0 13 9 0 3 9 13 3 13 9 0 13 13 2
17 7 3 13 0 9 2 0 9 0 13 1 13 2 1 9 0 2
11 1 3 0 9 9 9 13 13 1 9 2
6 0 3 9 9 13 2
9 13 3 9 0 13 1 9 0 2
17 15 3 13 9 2 0 0 9 2 9 13 9 1 0 13 3 2
14 1 3 0 9 13 9 13 2 1 3 9 13 0 2
22 15 3 9 7 9 0 9 7 9 13 3 3 2 7 1 9 9 1 9 13 0 2
6 3 3 3 9 13 2
5 13 3 0 9 2
14 9 3 9 7 0 9 9 13 1 9 9 0 13 2
9 3 3 3 9 9 13 9 9 2
11 3 0 9 13 9 3 0 7 9 9 2
12 0 3 13 9 2 13 9 2 0 9 9 2
12 15 3 9 7 9 0 13 9 9 0 13 2
18 3 3 15 9 9 13 2 16 3 0 9 15 13 9 9 13 13 2
16 3 3 3 3 15 3 9 15 13 13 1 10 9 3 15 2
3 15 13 2
10 3 3 0 3 13 2 16 15 0 2
11 10 3 0 13 0 9 13 3 0 13 2
9 7 13 15 10 0 0 13 3 2
29 3 3 13 10 0 0 13 16 13 3 0 2 3 0 0 10 0 9 13 0 13 2 1 3 15 3 10 0 2
15 3 3 15 13 1 9 13 13 10 9 2 13 13 15 2
13 7 15 13 2 15 3 13 15 13 13 10 0 2
30 3 3 13 15 1 10 0 13 0 10 9 2 7 3 13 3 13 1 10 9 2 13 16 0 10 0 1 10 0 2
24 7 15 3 3 2 16 15 13 1 10 9 1 10 0 2 13 0 10 13 2 13 3 13 2
17 3 0 15 3 0 13 15 13 2 7 7 13 15 0 10 0 2
10 7 0 0 13 13 2 7 3 13 2
14 0 3 1 3 3 1 15 13 2 3 3 13 13 2
16 3 3 15 3 13 0 15 13 7 13 3 13 10 15 9 2
31 15 3 13 16 1 9 13 0 15 13 3 0 9 13 2 3 0 1 9 2 7 3 13 3 3 16 15 15 13 13 2
5 13 0 7 13 2
2 13 2
6 15 13 3 13 13 2
4 13 15 13 2
13 0 3 13 13 2 15 3 13 13 3 3 9 2
10 13 3 15 10 9 7 15 10 9 2
16 3 3 13 3 10 13 3 0 13 7 3 3 3 9 13 2
13 13 3 3 10 0 15 10 13 1 10 0 9 2
21 0 3 10 9 13 16 13 10 0 13 7 3 13 15 3 7 0 10 9 13 2
12 13 3 7 13 10 9 15 10 0 13 0 2
26 10 3 9 13 10 9 7 10 9 0 2 13 1 9 15 2 13 3 9 13 10 9 15 13 13 2
13 13 3 2 15 13 13 10 0 7 15 10 0 2
40 0 3 10 9 13 13 10 9 10 9 0 7 0 2 7 0 13 10 0 9 13 16 10 9 13 3 1 9 2 0 3 3 10 0 9 13 1 0 0 2
15 15 3 3 13 2 15 3 3 0 13 1 0 9 13 2
61 7 9 15 13 15 13 10 13 1 10 9 1 0 2 7 9 3 0 7 9 7 0 0 0 2 0 13 3 1 10 0 2 7 1 10 0 9 10 3 0 0 15 13 2 7 3 7 10 0 0 10 9 0 10 0 9 13 1 10 9 2
4 3 3 13 2
10 7 0 3 15 1 3 1 9 13 2
10 3 3 15 3 15 13 13 0 13 2
4 7 3 13 2
30 13 3 16 3 0 15 13 2 9 15 7 12 15 13 10 0 0 2 7 0 0 10 9 0 0 10 0 0 13 2
15 13 3 3 0 9 10 3 0 0 13 7 10 0 0 2
4 7 3 13 2
5 7 3 13 3 2
15 13 3 10 3 10 9 0 0 2 10 3 3 0 0 2
19 16 3 3 2 0 3 13 2 7 15 0 7 13 16 13 0 15 13 2
7 13 3 2 13 15 13 2
14 3 0 3 13 2 7 10 0 2 10 0 10 0 2
6 7 3 3 13 13 2
3 13 3 2
3 13 3 2
4 3 3 13 2
37 3 3 16 13 15 3 7 15 1 9 0 0 2 10 1 0 9 0 3 15 13 7 13 0 2 7 1 9 13 1 3 10 0 0 3 13 2
20 3 7 1 10 0 7 0 6 13 2 1 10 13 13 0 13 3 10 9 2
3 13 0 2
28 3 3 0 15 13 2 7 15 13 13 16 15 13 10 3 0 7 10 0 7 0 7 0 7 0 7 0 2
32 15 3 0 13 1 15 13 7 3 13 1 0 9 0 13 0 0 13 2 16 13 2 7 15 7 15 7 10 0 9 0 2
11 3 16 15 13 2 1 0 0 13 3 2
12 3 3 3 3 13 0 16 3 1 0 13 2
3 3 13 2
20 3 15 0 13 0 7 0 7 0 2 0 7 13 2 10 3 0 0 13 2
2 13 2
2 13 2
15 3 3 0 3 13 2 15 13 0 13 0 3 7 0 2
13 0 3 3 13 0 13 7 3 7 1 10 9 2
12 13 3 0 2 0 13 7 13 13 10 9 2
8 3 3 0 3 13 7 13 2
3 0 13 2
30 3 3 0 3 13 2 16 3 10 13 13 13 9 2 7 0 3 13 2 10 15 13 10 13 7 15 13 7 15 2
3 0 13 2
21 13 2 1 0 13 15 15 0 13 16 0 3 0 9 13 3 13 0 10 9 2
12 16 15 3 13 2 13 15 1 9 3 13 2
2 13 2
3 7 13 2
33 16 3 3 15 9 13 16 10 9 0 10 0 9 13 0 13 2 15 3 15 13 1 0 15 3 13 10 0 3 7 10 0 2
12 7 3 3 0 13 3 13 10 0 7 3 2
8 10 3 0 13 7 0 13 2
12 16 13 2 0 0 13 9 0 7 0 13 2
27 7 15 13 3 15 13 10 0 15 3 0 10 9 13 2 7 10 0 2 15 3 0 9 13 2 0 2
7 7 0 15 13 10 13 2
2 0 2
8 13 3 15 15 3 3 13 2
5 13 3 10 15 2
17 15 10 0 16 0 13 13 1 10 9 2 7 16 13 0 13 2
6 7 15 13 0 13 2
26 13 15 13 7 13 7 13 7 13 7 13 7 13 7 0 10 0 13 16 0 0 13 7 3 0 2
5 15 15 13 13 2
11 3 7 13 15 13 7 0 0 10 13 2
17 13 3 15 2 0 10 13 16 13 13 13 2 7 1 0 15 2
21 3 3 16 13 3 13 2 1 15 13 2 7 10 0 16 13 2 1 15 13 2
17 3 16 13 13 2 1 15 13 2 7 16 13 2 1 15 13 2
10 3 16 13 13 2 7 16 13 13 2
24 13 3 15 2 16 16 15 13 7 15 13 2 3 16 13 13 13 2 7 16 13 13 13 2
12 3 16 13 13 13 2 7 16 13 13 13 2
5 7 3 13 3 2
14 3 3 10 13 7 13 15 13 7 13 15 1 15 2
9 7 15 3 3 13 3 10 0 2
14 3 16 13 13 13 1 15 13 2 7 16 13 13 2
12 0 15 13 1 9 0 2 16 10 0 9 2
2 13 2
13 7 3 3 16 3 13 1 9 13 13 7 0 2
3 0 13 2
13 3 3 13 16 3 13 2 3 3 0 13 0 2
11 15 3 3 2 16 13 2 13 0 13 2
7 15 3 13 2 3 13 2
17 13 3 3 15 3 15 3 13 7 3 13 13 3 3 13 0 2
37 7 16 3 0 15 13 7 13 2 3 3 15 13 16 3 7 15 1 10 0 9 10 1 10 9 9 13 7 3 13 13 3 3 15 0 13 2
8 3 3 0 3 10 9 13 2
6 0 3 15 13 9 2
12 3 3 13 15 13 2 16 3 0 15 13 2
33 10 3 13 0 0 7 3 13 1 10 0 3 15 13 10 13 2 7 15 15 13 10 9 2 16 15 3 1 13 3 0 3 2
14 7 3 0 15 10 9 13 0 2 16 0 13 0 2
21 13 3 3 15 10 9 13 7 3 13 3 16 1 10 9 9 10 9 9 13 2
19 16 3 15 13 15 13 2 0 15 13 13 16 3 15 13 1 10 0 2
4 7 3 13 2
13 13 3 16 3 0 15 13 0 13 0 10 0 2
12 7 3 0 3 15 13 3 0 16 0 0 2
7 15 3 0 13 10 9 2
4 13 15 3 2
9 3 13 15 13 3 9 3 3 9
23 0 3 15 13 7 9 7 9 7 0 0 0 13 13 3 2 13 3 9 0 15 13 2
5 3 3 15 13 2
4 13 3 3 2
6 3 3 3 13 13 2
7 1 0 3 13 9 9 2
6 13 3 3 3 3 2
8 10 0 3 3 3 13 13 2
7 3 13 7 3 15 13 2
6 13 3 15 3 13 2
36 16 3 3 15 15 13 15 15 3 2 0 0 9 13 9 10 0 7 15 13 13 0 10 9 2 13 3 16 15 3 7 0 13 7 0 2
5 7 3 13 15 2
8 10 3 9 3 13 15 13 2
10 3 3 9 0 13 13 7 10 0 2
3 3 13 2
7 3 9 3 0 0 13 2
24 1 0 15 13 7 9 10 13 2 3 13 3 16 10 9 1 10 0 13 13 7 0 13 2
5 7 3 13 15 2
10 7 1 9 13 10 13 10 9 13 2
18 3 3 3 10 9 9 13 9 9 3 13 9 7 0 10 9 13 2
18 7 15 15 13 3 2 16 16 15 0 13 2 0 15 10 9 13 2
5 3 3 0 13 2
2 3 2
10 7 15 3 9 9 13 3 10 9 2
2 13 2
15 13 3 3 13 10 9 0 1 15 9 9 13 13 0 2
7 1 15 9 9 0 13 2
12 10 3 9 0 1 15 9 9 0 3 13 2
14 7 3 10 0 0 13 10 9 10 1 10 9 9 2
7 15 10 0 13 10 9 2
42 15 3 15 3 13 2 16 16 3 13 15 13 10 9 13 3 7 13 13 3 7 13 2 0 13 10 0 2 7 13 10 0 15 3 0 9 7 10 0 10 9 2
22 7 3 3 16 1 0 13 13 2 15 16 13 2 3 3 3 1 15 10 9 13 2
25 3 3 9 3 10 13 10 13 13 3 3 0 13 2 15 3 3 13 10 0 13 7 10 9 2
15 3 10 13 13 13 10 9 2 10 3 13 13 10 9 2
14 9 3 9 7 9 9 9 3 13 1 0 10 9 2
8 13 3 13 0 7 13 0 2
18 3 3 3 10 3 3 13 3 13 15 13 1 0 2 0 0 13 2
15 3 3 3 0 3 3 13 13 13 15 0 15 0 13 2
19 13 3 15 2 15 10 9 10 9 13 13 1 10 9 15 1 15 13 2
11 0 3 15 13 0 15 3 3 0 13 2
22 7 0 0 13 1 10 9 2 16 0 10 0 1 0 13 2 0 3 1 15 0 2
7 13 15 0 3 3 0 2
13 7 3 13 16 10 9 15 13 3 1 0 13 2
21 13 3 3 16 1 10 3 10 3 0 7 10 0 3 0 15 13 7 0 0 2
4 7 3 13 2
13 3 3 3 13 16 10 10 9 0 13 0 13 2
8 15 3 0 15 16 0 13 2
17 3 7 3 3 3 13 2 7 16 3 3 2 3 3 3 13 2
2 13 2
21 1 9 3 15 3 0 15 13 10 0 2 16 15 16 3 13 0 13 3 13 2
18 13 3 16 15 0 9 2 7 3 0 13 3 10 9 16 3 13 2
45 16 3 3 13 3 10 3 0 7 10 0 2 3 13 16 3 3 13 1 9 9 9 9 9 13 9 2 7 3 10 9 3 13 13 16 3 3 0 13 2 7 10 9 13 2
14 3 3 3 13 16 3 13 13 10 3 0 7 3 2
10 3 3 13 3 2 7 15 9 13 2
56 1 9 15 13 0 13 15 13 2 16 1 15 13 10 3 0 7 7 7 10 1 9 9 13 2 13 0 16 0 3 1 0 10 0 13 7 16 3 1 9 13 3 13 1 0 2 7 3 7 10 0 9 3 0 13 2
48 10 3 3 1 15 9 2 10 13 9 13 9 2 10 9 13 10 9 1 10 13 9 10 9 9 1 10 9 7 1 10 13 9 1 10 0 9 10 9 1 9 1 10 9 9 10 9 2
33 1 13 3 3 9 9 13 0 9 9 7 9 9 9 2 13 7 3 1 9 9 0 1 10 0 2 1 15 13 0 9 0 2
15 1 3 15 9 10 9 13 1 10 9 1 0 10 9 2
21 9 10 9 9 3 7 9 13 9 2 1 7 9 7 9 3 13 1 10 9 2
15 15 0 13 10 9 7 10 9 13 2 13 0 9 13 2
15 3 13 10 9 13 10 9 2 3 3 13 1 10 9 2
20 9 3 0 9 1 10 9 13 13 0 3 1 10 0 9 2 9 7 0 2
24 10 3 9 13 1 10 10 9 9 2 13 0 10 9 15 0 3 10 9 10 9 13 0 2
16 3 3 10 9 0 9 13 13 9 0 0 10 0 7 0 2
16 13 3 15 3 10 9 9 2 1 10 9 9 13 0 9 2
18 3 3 15 13 1 9 1 9 9 13 2 3 13 1 10 13 9 2
35 3 9 3 13 3 13 1 10 9 13 13 2 10 7 9 1 3 10 10 9 9 7 10 10 9 9 2 16 13 2 13 13 10 9 2
40 16 3 15 0 10 1 10 9 13 2 10 3 9 13 13 10 9 1 9 7 9 2 15 7 1 0 10 9 13 10 0 7 0 9 2 13 1 10 9 2
44 10 3 9 13 13 10 0 13 3 10 9 2 13 7 10 9 1 10 9 10 9 2 3 3 10 9 0 7 0 10 9 13 2 3 7 10 9 10 9 13 13 10 9 2
17 10 3 3 13 1 10 9 10 9 3 13 1 10 9 10 13 2
24 10 3 9 13 10 9 10 10 9 9 2 13 1 9 0 9 10 13 10 1 10 9 9 2
12 13 3 10 3 9 9 2 10 7 9 9 2
16 15 3 1 10 9 9 13 13 13 9 10 3 13 10 9 2
17 13 3 0 10 9 9 13 10 9 7 13 10 1 10 9 9 2
36 16 3 10 9 7 10 0 9 10 0 10 9 13 10 0 9 3 7 9 10 13 9 1 9 2 13 10 1 10 9 9 13 1 10 0 2
25 0 3 13 10 9 10 10 10 9 13 2 16 13 9 13 10 9 10 9 3 13 10 0 9 2
42 9 3 3 3 9 3 9 3 9 7 9 1 10 9 13 2 3 13 10 1 10 9 9 2 0 7 9 3 9 3 9 7 9 10 0 15 13 13 1 10 9 2
41 10 3 1 9 13 10 9 13 10 3 3 10 9 13 10 9 13 10 9 2 16 10 9 13 2 1 7 10 10 9 13 13 9 10 13 13 1 10 0 9 2
27 15 10 3 13 3 10 9 2 10 7 13 1 0 9 2 13 10 0 0 9 7 13 10 10 9 9 2
19 0 3 9 13 1 10 0 9 13 13 2 16 15 9 0 10 9 13 2
30 1 3 15 10 1 9 9 13 10 9 3 9 7 9 13 2 10 9 0 1 10 9 13 10 1 10 0 9 9 2
22 9 3 16 13 10 9 13 7 10 9 13 2 13 1 10 9 1 9 10 9 13 2
16 16 3 13 1 9 2 1 10 9 10 9 13 1 10 9 2
17 13 3 1 10 9 0 13 9 3 10 9 7 10 0 15 9 2
22 16 3 13 1 10 13 9 2 3 13 10 0 2 16 0 10 9 1 9 9 13 2
9 13 3 3 10 9 10 9 0 2
7 10 3 0 0 0 13 2
47 10 3 9 13 9 3 10 1 10 9 13 1 9 7 9 0 2 9 3 1 9 7 9 0 2 9 3 1 9 7 9 0 2 9 3 0 1 10 1 10 9 13 2 9 7 0 2
15 10 3 9 10 1 9 3 9 7 9 13 13 10 9 2
18 9 3 3 15 10 9 13 2 0 3 0 0 2 10 7 0 0 2
14 10 3 3 9 1 10 9 10 9 13 1 10 9 2
17 13 3 10 10 10 9 13 3 13 7 13 1 10 0 10 0 2
28 13 3 10 3 9 0 9 10 0 2 10 7 1 9 13 9 10 10 9 9 2 0 13 1 9 7 9 2
14 15 3 13 10 9 13 0 0 1 10 9 13 15 2
45 10 3 9 13 16 0 3 13 1 0 9 2 7 13 0 13 2 13 1 15 1 0 16 1 3 10 13 10 9 13 10 9 0 2 1 7 3 10 9 1 15 13 3 0 2
19 0 3 7 0 10 9 13 2 13 15 16 1 0 0 9 15 13 13 2
22 13 3 16 10 9 3 1 10 9 13 10 9 2 10 7 9 1 10 0 9 13 2
26 10 3 3 9 13 0 2 7 1 15 9 0 2 10 7 0 9 10 1 15 13 1 10 9 0 2
33 10 3 3 9 1 0 13 1 10 9 2 9 7 10 3 10 9 13 13 3 9 7 9 10 9 2 13 7 13 13 10 9 2
16 16 3 13 10 9 13 1 9 2 13 7 13 1 10 9 2
30 13 3 1 10 9 3 9 0 3 9 15 7 9 3 0 13 10 0 2 3 7 3 9 1 10 0 9 3 0 2
15 13 3 10 10 9 13 1 15 1 10 1 10 9 9 2
22 10 3 3 1 9 13 9 15 10 9 13 13 1 10 9 2 13 10 10 9 9 2
42 9 3 1 10 9 10 9 13 1 0 10 9 2 7 1 3 9 9 10 0 9 13 13 0 10 9 2 3 7 1 10 13 9 13 1 10 0 9 3 7 3 2
15 16 3 13 1 10 0 9 2 13 10 0 13 10 9 2
34 3 3 13 10 9 13 10 1 10 9 0 2 3 0 13 10 0 9 2 16 13 15 10 0 3 0 10 0 9 1 10 0 9 2
40 10 3 0 9 10 3 1 10 0 9 13 7 10 10 9 7 10 0 9 13 3 0 13 10 13 2 16 15 0 13 10 13 1 10 9 10 1 9 13 2
21 13 3 10 0 9 1 10 10 9 9 13 2 10 7 9 10 10 9 9 13 2
15 0 3 3 9 10 1 0 9 13 10 1 9 13 13 2
27 13 3 15 13 2 16 9 9 13 10 3 9 0 13 2 15 7 0 1 10 9 13 7 0 13 9 2
18 3 15 13 0 13 13 9 10 9 0 7 0 10 3 1 15 13 2
31 10 3 1 10 9 13 10 9 13 2 16 3 13 10 9 0 1 10 9 13 7 13 13 1 15 0 1 10 9 13 2
23 1 3 10 9 15 13 13 2 3 0 13 10 9 3 1 9 2 7 1 9 13 9 2
45 10 3 9 13 1 10 9 10 10 9 9 13 9 9 2 1 10 9 13 1 15 2 13 7 10 9 13 10 9 2 0 10 9 0 10 0 9 13 7 1 0 9 13 13 2
15 10 3 9 13 13 16 3 0 15 10 9 10 9 13 2
9 10 3 13 10 9 0 9 13 2
22 3 3 13 10 1 10 0 9 0 10 9 13 1 10 0 9 0 13 1 10 9 2
14 10 3 9 13 15 13 13 2 16 13 13 10 9 2
28 10 3 9 13 13 1 10 1 9 9 2 13 0 10 9 9 2 3 1 9 13 15 7 3 13 0 13 2
15 13 3 3 9 10 9 2 10 10 9 9 3 3 13 2
20 13 3 10 9 3 10 1 9 13 9 7 9 2 13 15 0 13 10 9 2
14 10 3 3 9 0 10 9 13 13 10 13 10 9 2
14 10 3 9 3 13 13 10 9 1 10 0 10 9 2
37 13 3 9 0 2 7 10 3 9 9 13 10 9 10 9 2 10 7 9 13 10 9 7 13 1 10 9 1 10 9 2 0 13 13 10 9 2
26 3 3 13 10 9 7 10 9 1 9 13 2 3 7 10 9 13 2 1 0 9 0 13 10 9 2
17 10 3 9 13 10 9 7 10 9 10 9 2 3 13 10 9 2
11 0 3 3 15 13 2 3 0 7 13 2
41 9 3 10 9 13 0 3 10 1 10 9 9 9 13 2 10 7 9 3 13 10 10 9 9 2 13 10 10 9 0 2 13 0 7 13 10 9 13 10 13 2
30 16 3 3 15 0 13 9 13 2 3 3 10 9 13 13 2 1 3 10 9 0 13 2 1 7 10 9 0 13 2
50 10 3 0 9 3 2 1 9 15 10 9 13 10 9 2 1 0 10 9 13 10 13 9 7 9 13 2 7 0 13 15 13 2 7 13 3 15 10 9 9 0 13 2 13 7 9 13 10 9 2
30 1 15 3 13 10 9 2 16 10 13 1 9 13 10 9 3 13 2 7 10 9 10 9 13 0 13 10 0 9 2
8 13 3 10 9 13 1 15 2
24 10 3 3 0 1 10 10 0 9 13 2 10 7 0 1 10 10 0 9 3 7 9 13 2
21 9 3 13 3 10 0 2 10 10 13 9 13 10 9 13 3 13 13 10 0 2
7 3 13 3 13 7 13 2
25 13 3 10 9 7 13 15 13 3 13 2 13 1 15 0 0 10 0 2 0 13 10 0 9 2
38 15 10 9 13 13 1 0 9 0 7 0 10 9 13 2 7 13 10 13 15 3 10 1 10 9 2 7 0 10 9 13 15 1 10 0 3 13 2
17 10 3 9 0 13 2 7 13 9 10 0 13 15 9 0 9 2
44 10 3 1 10 9 15 9 9 2 10 9 13 0 2 0 7 7 10 9 13 0 2 13 1 10 10 9 9 9 13 1 10 1 10 9 2 7 10 1 10 0 13 13 2
15 13 3 10 9 13 1 0 9 7 13 1 10 13 9 2
14 0 3 3 13 13 3 13 10 9 13 1 10 0 2
51 9 3 10 9 10 9 13 15 3 9 13 0 7 10 9 2 13 10 3 0 9 0 13 7 13 15 2 16 1 10 0 9 13 10 9 2 0 7 10 9 13 13 13 7 10 9 10 9 3 13 2
20 3 3 10 3 15 0 13 2 10 7 9 1 10 9 0 9 7 0 13 2
55 1 3 15 10 3 1 10 0 9 13 10 9 3 10 1 10 9 13 1 10 0 2 10 7 9 10 3 9 13 2 10 7 9 13 2 0 9 10 13 13 13 1 10 0 2 3 16 13 10 9 10 10 0 9 2
18 9 3 10 9 10 9 13 2 15 13 3 13 2 3 1 9 13 2
22 15 3 3 10 9 9 13 2 13 3 13 0 9 13 7 13 10 1 10 9 9 2
28 7 3 3 13 15 0 0 13 2 13 10 9 13 1 10 9 13 10 13 7 1 0 13 10 10 9 9 2
19 15 3 3 3 10 9 13 9 13 1 10 10 9 9 2 13 10 9 2
24 3 3 0 3 1 10 1 10 9 13 2 0 7 1 10 0 7 1 0 1 10 9 13 2
22 10 3 3 9 13 10 0 9 2 10 7 9 1 0 13 10 9 3 0 13 9 2
25 13 3 15 2 3 13 10 9 10 9 0 1 10 3 9 9 3 9 9 7 3 9 9 13 2
28 16 3 3 10 9 13 1 10 0 9 2 3 3 3 15 1 10 9 13 7 10 9 0 0 3 13 9 2
26 3 3 10 3 9 13 13 1 10 9 2 10 7 9 13 1 10 9 10 13 1 15 3 0 13 2
14 10 3 9 13 13 1 0 10 9 13 10 9 3 2
48 9 3 13 7 10 0 9 13 2 10 3 9 13 0 13 10 9 2 13 15 2 7 1 9 3 3 13 2 13 10 9 15 2 1 7 10 9 7 3 13 3 3 13 7 13 0 13 2
17 10 3 3 1 9 10 1 9 9 13 0 13 10 9 10 9 2
8 15 10 9 15 3 3 13 2
36 15 0 9 13 10 3 13 9 1 10 9 3 13 2 10 15 7 9 3 13 1 10 0 10 9 9 2 7 3 13 13 3 16 13 3 2
12 3 10 10 9 3 9 3 3 15 13 13 2
9 15 3 3 10 9 13 10 13 2
15 15 3 3 13 16 0 10 9 13 13 13 10 0 9 2
30 3 3 15 3 3 10 0 13 10 9 10 9 2 15 10 9 10 9 13 10 3 9 13 2 10 7 9 3 13 2
16 3 15 0 10 13 13 0 13 10 15 10 10 0 9 13 2
16 13 3 3 1 10 9 13 10 0 9 2 7 1 10 9 2
13 10 3 3 10 9 9 2 10 7 10 9 13 2
23 3 3 3 15 15 3 10 0 10 9 9 0 13 16 10 9 1 10 1 9 9 13 2
19 0 3 10 9 13 10 3 9 13 2 10 7 9 13 1 10 0 9 2
15 3 3 0 10 1 15 1 10 9 10 9 1 9 13 2
18 3 3 10 10 9 9 0 2 7 0 3 10 9 13 15 10 9 2
11 9 3 0 3 9 7 10 9 13 9 2
9 9 0 0 9 9 9 9 13 2
16 13 3 3 9 10 9 9 2 9 0 13 9 0 7 9 2
17 15 3 3 1 10 0 10 9 9 13 13 1 10 0 10 13 2
16 7 3 0 10 9 13 2 10 1 10 9 9 13 13 9 2
25 3 3 10 13 10 9 9 13 13 13 1 10 10 9 0 7 13 0 10 9 13 1 10 9 2
26 10 3 10 10 9 9 13 1 9 10 0 13 0 10 9 2 7 13 10 9 1 9 10 13 9 2
20 3 3 0 9 13 13 9 0 3 1 10 0 2 0 7 7 10 15 0 2
11 13 3 10 9 13 13 1 9 10 9 2
19 3 3 0 9 13 2 13 10 9 13 7 10 9 0 13 13 10 0 2
19 10 3 9 13 3 1 9 10 9 2 13 7 10 0 9 0 7 0 2
17 3 15 13 10 3 9 0 7 0 2 10 7 0 10 0 9 2
19 15 3 9 3 13 9 10 9 2 13 7 10 1 10 9 9 10 0 2
32 15 3 1 9 7 9 0 9 13 3 0 1 10 1 10 0 9 2 7 3 1 0 10 9 2 7 0 15 13 3 13 2
47 13 3 9 1 10 10 9 9 1 10 9 2 10 3 15 0 10 9 13 13 7 10 9 10 0 13 2 0 7 9 10 0 13 9 2 13 16 13 0 10 9 13 13 1 10 0 2
15 9 3 1 10 9 9 10 9 0 10 9 10 0 13 2
34 10 3 9 1 0 9 13 2 10 3 0 10 1 10 9 13 10 9 13 0 3 9 13 2 3 0 7 13 13 1 10 9 13 2
60 1 3 10 9 9 13 0 0 1 10 9 13 10 9 13 2 16 13 10 0 13 10 9 2 16 10 9 10 0 9 13 0 10 10 9 9 13 7 1 10 9 0 16 10 3 9 3 3 13 2 10 7 9 3 1 10 9 13 0 2
16 3 3 3 13 15 1 10 9 0 10 9 13 1 10 0 2
14 10 3 9 2 13 15 9 0 0 2 13 10 9 2
12 13 3 15 10 9 0 10 1 10 9 9 2
20 13 3 9 0 0 9 1 0 13 2 7 9 13 13 13 1 10 0 9 2
19 13 3 1 0 10 9 13 1 3 10 9 9 2 1 7 10 9 9 2
24 1 3 15 10 9 13 10 1 9 13 2 13 7 3 10 9 0 13 1 10 9 2 13 2
7 3 13 1 9 13 3 2
29 10 3 9 13 3 13 10 1 10 9 2 9 3 9 7 10 15 0 0 0 13 1 10 9 13 13 1 9 2
34 10 3 10 9 9 13 10 10 0 9 2 13 1 10 9 1 0 10 9 2 7 10 10 9 9 9 13 7 13 10 9 15 13 2
28 1 3 15 13 9 1 10 9 13 13 1 10 9 9 2 13 3 10 9 2 13 7 10 1 10 9 9 2
32 10 3 9 10 10 9 13 2 3 13 15 3 0 13 2 10 3 9 0 13 3 2 1 7 10 9 10 1 10 9 13 2
14 1 3 15 10 9 10 3 10 9 9 13 15 13 2
4 13 3 9 2
38 3 3 9 3 10 9 13 2 7 13 1 9 13 7 10 3 9 10 9 13 2 10 7 9 13 2 15 7 1 10 0 9 13 1 10 9 13 2
62 10 3 1 10 9 10 9 13 13 3 1 10 9 10 9 9 2 3 7 3 9 0 7 9 0 1 10 13 13 2 1 7 15 10 9 9 0 13 1 10 9 10 9 2 13 13 0 10 9 2 0 7 13 10 10 9 9 13 1 10 9 2
13 10 3 3 1 9 9 0 0 9 10 9 13 2
20 9 3 1 10 9 13 10 3 10 9 9 13 2 10 7 9 0 13 13 2
12 10 3 1 10 0 15 13 13 1 9 3 2
23 1 3 15 1 10 9 13 10 3 9 13 2 10 7 9 13 7 10 10 9 9 13 2
27 10 3 9 1 15 13 2 13 10 9 1 10 9 1 10 9 2 13 10 3 9 7 10 9 10 9 2
60 1 3 0 10 9 9 3 13 0 9 13 1 10 9 2 16 3 15 13 2 3 13 13 10 1 10 9 9 2 16 7 15 10 9 13 2 13 10 10 9 9 2 16 9 3 13 15 13 9 7 9 2 10 7 9 13 13 15 13 2
16 3 3 3 10 0 9 0 13 9 3 13 1 0 10 9 2
20 13 3 15 0 10 1 9 13 13 7 13 2 1 0 9 13 13 10 9 2
26 0 3 7 0 9 13 2 10 3 9 2 10 0 0 9 13 2 13 13 1 10 9 13 10 9 2
12 9 3 13 1 10 9 13 10 9 10 9 2
15 3 3 10 1 10 9 9 13 3 0 13 1 10 9 2
19 3 3 3 15 0 13 0 10 9 2 0 13 15 0 13 0 10 9 2
22 9 3 0 9 13 1 9 13 2 10 3 9 13 10 1 10 9 7 1 10 9 2
18 10 3 3 9 13 10 9 13 13 10 9 7 13 1 10 13 9 2
30 3 3 10 9 13 2 3 0 13 10 9 10 0 9 15 13 10 9 2 7 0 1 10 9 13 13 1 10 9 2
42 15 3 0 3 10 0 9 10 9 13 10 10 0 9 2 10 3 10 1 9 9 10 0 9 13 9 2 7 10 1 10 9 9 1 9 9 0 9 13 10 9 2
20 10 3 0 10 9 13 10 10 9 9 7 10 0 9 2 13 13 10 9 2
50 3 0 10 9 13 1 10 9 7 10 9 10 13 2 10 3 9 13 10 9 2 13 1 9 0 1 9 1 9 2 10 7 1 10 9 13 1 0 10 9 13 1 15 2 16 3 13 10 9 2
32 10 3 9 13 10 3 9 9 3 13 13 10 10 9 9 2 10 7 1 9 9 13 0 13 1 10 9 2 13 15 0 2
25 13 15 1 10 9 13 7 13 2 16 13 10 1 9 9 13 1 10 9 7 1 10 9 13 2
22 3 10 9 1 10 9 10 13 13 2 13 13 10 0 9 10 9 10 0 9 13 2
21 3 3 10 10 0 0 13 2 13 13 10 1 9 10 3 9 7 10 9 9 2
21 10 3 0 9 10 9 13 1 10 9 2 13 13 10 0 7 9 13 10 9 2
19 13 3 10 9 13 1 9 3 2 16 1 10 9 7 9 3 15 13 2
24 3 3 13 10 0 9 2 10 3 0 9 13 9 2 10 7 0 10 1 10 9 13 9 2
33 10 3 10 9 9 13 9 0 1 10 9 10 13 1 10 13 10 9 7 1 10 0 9 2 7 16 1 10 9 13 10 9 2
28 9 3 10 1 10 9 7 9 13 10 9 2 10 3 0 9 13 9 7 9 2 1 10 10 9 0 13 2
21 0 3 10 9 9 13 1 3 10 9 7 1 10 1 9 1 10 0 9 9 2
9 9 3 7 9 10 0 9 13 2
28 15 3 13 13 0 1 10 9 7 3 13 1 10 0 10 9 0 13 9 2 16 0 13 9 1 10 9 2
11 10 3 0 9 13 10 0 10 9 9 2
18 15 3 3 0 10 9 13 13 2 7 10 9 1 9 7 9 13 2
29 10 3 9 10 3 9 13 13 10 0 2 15 7 1 10 0 9 10 9 13 2 1 15 13 13 10 9 13 2
15 10 3 9 10 3 0 13 13 10 9 2 13 0 9 2
21 16 3 1 10 0 13 2 13 10 9 15 1 10 9 13 2 7 0 13 9 2
14 10 3 9 13 10 9 7 0 13 9 13 3 13 2
12 10 3 9 13 2 9 13 10 0 10 9 2
14 0 3 3 13 10 13 2 3 10 15 7 0 13 2
16 3 3 10 13 1 10 3 13 2 13 7 13 1 10 9 2
25 10 3 9 13 10 9 10 9 13 10 0 2 7 10 3 10 9 13 2 15 7 10 9 13 2
17 10 3 9 3 13 2 0 10 9 9 0 13 10 9 3 13 2
15 3 3 9 3 13 13 2 1 10 3 7 13 3 13 2
49 10 3 9 7 9 9 1 10 9 13 2 10 10 9 7 9 2 3 7 3 9 9 2 13 15 13 2 10 3 0 3 13 2 16 7 13 10 0 9 1 9 13 2 3 15 10 9 13 2
15 1 3 0 9 13 0 9 1 3 15 0 13 10 9 2
25 16 3 10 9 1 10 9 13 10 9 7 9 13 2 13 1 15 13 10 9 7 0 9 13 2
14 10 3 3 9 0 10 9 13 0 9 10 9 13 2
24 1 3 10 9 13 9 10 3 9 0 2 10 7 9 1 10 0 1 10 1 0 9 13 2
26 10 3 9 1 9 13 10 3 9 10 13 10 9 10 0 13 2 10 7 15 13 13 10 13 9 2
23 10 3 9 13 10 9 10 3 0 1 10 9 13 2 10 7 9 13 13 1 10 9 2
15 9 3 13 0 13 10 9 2 0 3 0 15 9 13 2
21 13 3 10 9 0 13 1 0 9 2 13 0 10 9 10 0 9 0 0 9 2
23 10 9 10 0 9 13 1 10 9 13 2 16 13 10 9 13 1 10 9 13 10 9 2
60 3 10 9 13 10 9 1 10 9 2 0 13 16 10 1 10 9 9 13 2 10 9 13 2 13 7 10 0 13 1 10 9 1 10 9 2 13 9 1 10 9 1 10 0 9 3 7 0 2 15 10 0 9 13 3 0 10 0 9 2
13 9 3 3 0 9 13 0 9 0 13 10 9 2
11 3 10 3 1 10 9 13 1 15 13 2
19 15 3 3 13 1 10 1 10 9 13 2 13 10 9 1 10 0 9 2
24 9 3 13 1 9 10 0 9 13 10 1 10 9 9 2 0 9 13 10 1 10 9 0 2
18 16 3 0 0 15 13 2 9 13 9 2 10 3 1 15 13 13 2
45 15 3 13 0 3 7 0 9 0 13 1 10 9 2 13 0 3 9 3 0 10 0 9 2 9 7 0 0 10 0 2 7 3 0 9 9 10 13 10 9 2 1 10 0 2
20 15 3 3 13 10 0 9 7 13 13 10 9 10 13 10 9 7 10 9 2
15 13 3 10 9 1 10 1 10 9 9 13 10 9 13 2
28 1 3 0 9 13 10 9 7 13 10 1 10 9 13 9 2 13 1 10 9 1 10 9 2 13 10 0 2
36 3 10 3 0 9 0 13 7 9 0 7 9 0 13 2 10 7 10 0 9 13 0 13 10 9 7 13 1 10 0 9 1 10 13 9 2
40 3 3 0 10 1 9 9 13 2 10 3 9 0 1 10 9 9 13 2 10 7 9 0 3 13 2 13 1 3 10 9 7 9 9 7 10 0 9 13 2
27 15 3 10 0 10 9 13 13 1 10 9 2 7 10 9 10 13 13 7 0 13 13 10 1 10 9 2
29 3 3 9 10 9 9 2 13 9 0 7 13 10 9 2 13 3 13 1 10 9 2 13 10 9 13 10 0 2
37 10 3 9 3 0 13 13 10 9 2 13 7 10 10 9 9 13 1 10 9 1 9 2 13 0 3 3 0 10 0 2 9 7 1 10 0 2
22 13 3 3 10 9 7 13 10 9 10 9 2 13 13 10 0 13 10 10 9 9 2
40 15 3 3 9 0 13 10 1 10 9 9 2 15 3 13 9 0 7 9 13 2 10 7 9 0 13 1 10 1 10 9 13 10 0 7 1 10 9 13 2
18 15 3 3 13 13 3 1 10 9 2 0 13 0 0 0 13 13 2
26 13 3 0 1 10 9 0 16 0 2 10 3 9 0 9 13 2 10 7 1 10 9 13 10 9 2
41 0 3 15 13 10 3 9 0 10 9 2 15 1 9 0 13 10 1 9 2 0 10 0 1 10 9 13 2 7 15 13 2 1 15 13 13 1 10 13 9 2
23 3 3 9 9 7 9 13 3 13 2 1 0 9 13 10 9 3 15 3 13 10 9 2
15 13 3 15 3 10 0 1 10 9 0 2 0 13 9 2
57 13 3 10 9 0 1 15 13 13 10 9 9 2 1 15 9 13 0 9 2 15 13 13 13 10 3 9 7 13 1 9 1 10 0 9 2 3 13 9 0 2 13 7 1 10 0 9 10 3 9 13 2 10 7 9 13 2
25 13 3 3 9 1 10 13 9 2 15 13 2 16 13 10 9 13 1 10 9 2 13 10 9 2
15 15 3 1 9 10 9 13 13 10 1 10 9 13 9 2
20 3 10 9 13 10 9 2 10 9 0 10 9 13 13 1 10 9 10 9 2
23 10 3 1 10 9 10 9 9 10 3 0 13 10 9 13 10 9 7 13 9 3 13 2
29 3 3 10 9 1 0 10 9 13 10 0 2 7 9 10 9 3 13 2 13 0 10 9 10 9 13 10 13 2
23 10 3 9 13 15 13 2 0 13 9 10 13 2 7 9 13 15 3 0 10 0 9 2
29 10 3 0 13 1 0 9 0 10 3 0 13 10 13 2 0 7 13 9 7 10 9 13 13 15 13 10 13 2
32 9 3 0 9 13 2 7 15 13 3 1 10 0 9 2 0 13 10 9 3 0 1 10 9 2 7 3 1 10 15 0 2
24 15 3 10 1 15 13 0 9 13 2 3 0 1 0 9 13 10 9 7 9 0 0 13 2
43 3 3 0 10 9 13 0 10 9 10 1 9 13 10 9 7 9 10 9 10 9 10 9 2 7 10 9 1 10 0 9 10 9 10 3 15 2 10 7 10 0 13 2
39 3 3 10 1 10 9 7 10 1 10 9 1 10 9 13 10 9 10 0 9 2 10 1 9 0 13 13 10 1 10 9 13 2 13 10 10 9 9 2
51 3 10 10 0 9 1 0 13 1 3 10 9 13 13 10 9 7 0 9 1 15 2 1 7 10 9 3 0 13 10 9 2 7 3 10 13 10 9 13 2 7 10 3 13 3 9 1 10 9 13 2
23 3 3 15 10 0 9 13 10 13 9 3 1 15 13 2 1 7 10 0 10 13 13 2
37 13 3 10 0 9 10 9 13 7 10 1 9 1 9 13 1 9 2 3 3 10 9 1 10 0 9 13 13 10 3 0 9 7 10 0 9 2
26 1 3 10 13 9 1 10 9 10 9 0 9 0 13 10 9 2 15 9 3 13 1 10 0 9 2
20 3 3 10 9 3 0 10 3 13 2 10 7 13 2 13 15 10 9 13 2
34 10 3 9 1 9 0 9 13 1 15 13 2 16 10 9 0 13 13 10 9 2 3 10 9 0 10 9 3 13 13 1 10 9 2
30 10 3 3 9 2 10 3 9 13 2 0 7 9 0 9 13 0 13 10 3 10 13 9 7 10 0 9 10 13 2
24 10 3 9 13 16 13 13 1 9 9 2 3 13 1 15 9 9 10 0 13 3 7 13 2
23 10 3 9 1 10 9 10 3 9 10 13 10 9 9 13 7 10 15 10 13 9 13 2
17 10 3 9 10 13 13 2 13 10 1 10 9 9 13 10 9 2
32 10 3 15 0 3 1 9 13 10 0 10 9 2 10 7 0 1 10 0 13 10 0 2 1 10 9 10 13 10 9 13 2
19 10 3 9 1 9 13 10 13 0 2 7 10 0 10 9 1 0 13 2
13 0 3 13 9 10 3 9 15 7 10 9 13 2
20 0 3 1 15 10 13 13 10 9 2 16 0 10 9 1 15 13 9 0 2
51 13 3 15 1 10 9 10 0 3 0 16 0 9 13 13 1 10 9 2 7 3 16 13 10 9 0 10 13 1 10 0 13 2 3 7 1 10 9 2 15 0 1 10 9 13 13 10 9 10 13 2
52 0 3 1 10 0 13 2 15 3 10 9 13 2 1 15 3 0 10 0 10 9 9 13 2 7 3 1 10 10 9 1 10 9 9 0 13 15 10 9 2 16 0 13 10 9 2 3 1 10 9 13 2
20 13 3 10 9 3 9 0 2 10 0 13 9 0 2 10 7 9 9 0 2
19 1 3 15 13 9 7 0 9 9 13 2 0 13 9 1 9 7 9 2
13 9 3 0 1 15 13 13 10 9 15 0 13 2
37 3 15 3 1 10 0 9 13 13 7 1 10 9 10 9 13 2 10 7 9 0 0 13 0 13 7 9 0 13 2 16 13 1 15 0 9 2
33 9 3 10 0 13 10 9 13 1 10 9 2 7 1 10 9 10 9 9 13 3 0 1 10 9 2 7 3 1 0 10 9 2
17 13 3 0 15 9 2 16 13 1 10 9 13 10 9 0 0 2
32 3 3 3 10 0 13 9 3 7 9 13 1 15 9 2 1 3 10 13 13 9 2 1 7 10 0 13 0 13 10 13 2
25 10 3 0 3 13 9 13 2 7 10 9 3 13 3 1 15 0 2 7 3 1 10 0 9 2
21 10 3 9 3 10 9 13 15 3 13 13 7 9 0 10 9 10 9 9 13 2
29 15 3 1 15 13 13 0 1 10 9 10 9 2 7 13 1 15 0 9 9 2 9 13 10 13 1 15 9 2
18 15 3 13 3 0 9 0 2 13 7 1 10 9 1 10 9 0 2
16 13 3 0 9 13 1 10 9 7 13 10 9 1 10 9 2
32 15 3 3 0 10 9 0 1 10 9 13 2 7 3 9 1 9 13 13 3 1 0 10 9 7 10 13 15 1 10 9 2
41 1 0 3 10 13 13 10 9 2 7 13 3 16 0 15 13 10 13 15 13 2 0 13 10 3 13 9 3 9 2 16 0 9 0 13 9 3 9 7 9 2
34 1 3 15 13 10 9 1 3 10 9 13 9 0 9 7 9 2 0 7 0 13 1 9 0 13 1 10 9 10 1 9 9 0 2
13 13 3 0 3 1 10 9 13 9 9 9 13 2
12 15 3 3 13 2 13 10 9 1 10 13 2
11 10 3 9 9 13 13 1 0 10 9 2
14 10 3 3 0 10 13 1 0 10 9 3 15 13 2
17 1 13 3 3 9 9 3 13 0 9 9 9 7 9 9 9 2
22 1 3 15 10 3 10 9 9 1 9 1 10 1 9 13 9 13 13 1 10 9 2
17 3 3 13 2 16 10 9 13 2 13 1 9 2 13 10 9 2
11 13 3 10 0 9 1 9 0 10 0 2
12 15 3 3 3 0 13 10 9 13 10 9 2
13 3 10 9 13 10 13 13 13 10 9 10 9 2
5 15 3 13 13 2
6 10 3 9 13 15 2
19 0 3 13 9 10 9 9 13 1 15 7 0 10 9 1 10 9 13 2
16 1 3 15 1 10 9 13 1 0 9 0 1 10 0 9 2
16 10 3 3 9 3 13 0 13 1 10 9 10 10 9 9 2
13 10 3 9 13 10 13 7 13 13 10 13 9 2
18 9 3 10 9 1 10 0 9 10 9 13 3 13 10 13 10 0 2
16 3 3 15 13 13 1 9 9 13 13 10 1 10 9 9 2
25 15 3 13 10 1 10 9 13 10 13 10 9 9 13 9 7 9 13 0 1 10 10 9 9 2
5 15 7 13 13 2
11 10 3 9 13 10 1 15 13 10 9 2
6 0 3 13 10 9 2
11 10 3 9 10 9 13 0 13 10 9 2
14 3 3 15 13 13 10 9 13 3 7 1 9 13 2
17 3 10 3 0 0 13 3 0 13 10 9 7 0 1 0 13 2
13 0 3 0 13 9 10 1 10 9 9 10 9 2
12 13 3 10 13 10 9 13 13 15 10 9 2
16 13 3 16 3 13 1 10 9 10 9 3 9 13 10 9 2
12 3 13 13 10 9 7 13 13 1 10 9 2
13 10 3 3 0 13 9 13 0 0 13 10 9 2
15 1 3 10 9 9 1 10 9 13 7 9 13 0 13 2
9 15 3 3 13 1 0 10 9 2
18 1 9 3 9 9 1 9 10 0 9 13 9 9 7 9 9 9 2
16 3 3 13 15 10 9 1 10 9 15 13 10 13 10 9 2
23 3 3 3 9 1 10 9 3 9 1 10 0 9 7 0 15 13 10 9 13 10 9 2
13 3 3 3 13 0 1 10 0 9 13 10 0 2
26 3 3 9 13 1 10 9 10 9 3 13 1 10 13 3 13 10 9 1 10 3 13 3 10 9 2
18 3 3 13 1 10 9 0 0 0 9 13 1 9 9 13 10 9 2
15 13 3 15 13 10 9 13 10 9 13 10 1 9 9 2
14 10 3 3 13 3 13 10 9 3 13 1 10 13 2
28 13 3 15 1 3 10 9 9 13 10 13 13 10 0 10 9 9 13 0 9 1 10 1 10 9 13 9 2
13 0 3 0 0 1 10 10 0 9 9 13 13 2
8 10 3 3 9 1 15 13 2
10 13 3 0 7 9 13 0 0 9 2
14 3 3 3 13 3 10 0 10 9 1 0 10 9 2
21 9 13 13 16 10 10 9 1 15 13 1 10 9 3 13 7 13 9 10 0 2
14 1 0 9 13 15 1 10 13 10 9 13 15 13 2
9 15 3 3 13 1 0 10 9 2
23 1 3 10 9 9 13 13 10 9 7 13 10 3 9 15 13 7 13 10 1 10 9 2
13 15 3 3 1 15 3 13 13 9 0 7 0 2
18 13 3 10 9 13 1 10 9 10 1 10 9 1 10 1 9 9 2
19 9 3 10 9 13 10 9 13 13 13 10 1 10 9 1 10 9 9 2
17 1 13 3 3 9 1 9 10 0 9 13 9 9 7 9 9 2
14 3 3 3 13 1 10 13 13 13 7 9 13 13 2
12 3 3 10 0 9 0 13 10 10 9 9 2
11 13 3 9 0 0 13 9 1 9 13 2
17 1 3 10 9 9 1 9 13 9 0 9 13 1 10 13 9 2
9 15 3 3 13 1 0 10 9 2
17 1 13 3 3 9 9 3 0 13 9 9 9 7 9 9 9 2
17 1 3 15 9 3 0 7 0 9 13 1 0 13 10 13 9 2
14 3 3 3 13 10 9 3 3 13 10 10 9 9 2
10 13 3 15 1 10 13 3 10 9 2
16 0 10 9 1 9 13 10 9 10 13 3 13 13 10 9 2
15 10 3 3 9 10 13 9 13 13 1 10 9 1 9 2
10 1 15 3 13 10 9 10 0 13 2
22 3 3 1 10 13 9 1 10 9 1 10 9 9 13 10 9 1 10 0 13 9 2
8 13 3 1 10 9 9 13 2
21 10 3 9 10 3 0 13 15 3 3 13 13 7 10 0 13 13 15 10 9 2
22 10 3 9 13 0 13 9 10 9 7 1 10 9 10 9 10 9 10 9 0 13 2
14 10 3 9 0 13 1 10 9 9 0 15 9 13 2
12 1 15 3 13 0 9 7 0 9 13 13 2
15 15 3 1 0 10 1 10 9 9 0 10 9 13 13 2
12 15 3 10 9 1 9 10 9 0 13 0 2
20 1 3 15 13 1 10 9 9 3 10 10 9 13 9 7 9 9 13 9 2
17 1 13 3 3 9 9 3 0 13 9 9 9 7 9 9 9 2
14 1 3 10 3 13 9 13 9 1 0 13 10 9 2
19 10 3 9 13 3 10 9 10 0 9 7 9 13 13 10 0 9 13 2
20 10 3 9 13 0 7 0 13 10 9 0 3 13 7 15 10 0 13 13 2
18 3 3 13 0 7 0 9 13 1 10 0 9 3 0 7 0 9 2
9 15 3 3 13 1 0 10 9 2
19 1 13 3 3 9 1 9 10 0 9 13 9 9 9 7 9 9 9 2
12 1 3 15 0 0 7 0 13 9 10 9 2
21 1 3 10 9 13 9 0 13 13 10 9 1 0 7 10 9 0 10 0 13 2
13 3 1 15 13 3 10 9 13 10 1 10 9 2
26 10 3 9 10 9 9 1 10 0 9 3 1 10 9 13 10 9 7 1 10 9 3 10 13 13 2
15 10 3 9 13 1 10 1 10 9 9 13 1 15 9 2
15 15 3 0 3 1 10 0 9 13 9 0 10 9 13 2
15 1 3 15 3 13 10 1 10 9 3 3 10 9 13 2
13 3 3 1 15 10 1 9 1 10 0 9 13 2
14 3 3 10 9 13 1 10 9 1 10 9 13 15 2
12 1 3 15 9 7 9 13 9 1 0 9 2
9 15 3 3 13 1 0 10 9 2
16 1 13 3 3 9 9 13 0 9 9 9 7 9 9 9 2
14 15 3 3 1 10 9 13 1 9 10 9 13 13 2
15 1 13 3 3 9 9 13 0 9 9 7 9 9 9 2
15 10 3 9 13 9 10 0 10 9 3 3 13 10 13 2
14 13 3 3 0 3 0 7 3 10 9 7 9 0 2
22 3 3 0 15 13 13 13 10 0 9 1 10 9 9 7 10 1 10 0 9 9 2
19 1 3 10 9 9 13 10 9 9 10 9 13 10 9 10 1 15 13 2
7 13 3 10 1 9 9 2
27 10 3 3 9 13 3 9 13 1 10 9 13 9 10 9 15 9 13 10 9 7 10 9 1 15 13 2
10 13 3 15 0 13 10 0 10 9 2
19 10 3 13 7 15 13 1 10 9 13 10 9 7 13 15 9 0 13 2
17 3 3 13 10 9 7 10 9 10 9 13 13 10 10 9 9 2
12 3 3 3 9 13 9 13 10 9 13 13 2
15 1 13 3 3 9 9 13 0 9 9 7 9 9 9 2
14 10 3 3 9 1 0 9 1 10 10 9 9 13 2
13 3 10 3 1 10 9 7 10 9 1 15 13 2
14 1 3 15 3 1 9 7 9 13 1 0 0 9 2
9 10 3 9 0 10 0 9 13 2
5 15 3 13 13 2
18 3 3 10 1 10 9 9 10 13 3 13 7 0 10 0 13 13 2
10 3 10 3 1 10 9 1 15 13 2
17 15 3 13 9 9 3 7 0 1 10 0 9 13 13 10 9 2
25 10 3 9 3 9 13 7 3 13 10 1 9 13 13 10 1 10 9 9 10 9 0 9 13 2
15 1 13 3 3 9 9 13 0 9 9 7 9 9 9 2
17 10 3 1 10 9 9 10 1 10 9 13 1 10 9 9 13 2
9 15 3 13 9 3 9 7 9 2
16 3 3 15 3 9 1 9 10 9 9 13 13 13 10 9 2
11 1 3 15 9 3 9 13 1 9 13 2
14 13 3 3 10 9 10 0 9 13 1 9 10 9 2
15 10 3 3 0 10 9 15 13 13 7 1 0 9 13 2
16 1 3 15 9 3 9 10 9 13 13 10 9 1 10 9 2
13 9 3 13 10 1 10 9 13 10 9 1 9 2
5 15 3 13 13 2
17 13 3 10 9 0 15 13 10 1 10 3 9 13 9 10 9 2
33 10 3 3 1 9 13 9 3 10 1 9 1 9 9 7 10 0 10 0 10 9 9 13 15 13 10 9 15 13 9 10 9 2
18 13 3 10 9 1 10 10 0 9 7 10 0 9 15 13 10 15 2
14 1 3 15 1 10 9 13 13 1 9 10 13 9 2
17 9 3 3 1 0 9 0 9 13 0 13 10 9 1 10 9 2
9 15 3 3 13 1 0 10 9 2
20 10 3 9 13 15 13 1 10 9 10 0 10 13 10 9 7 10 9 0 2
13 0 3 13 3 13 3 7 1 10 9 13 13 2
9 3 3 13 13 10 9 1 9 2
17 1 13 3 3 9 9 3 0 13 9 9 9 7 9 9 9 2
17 1 13 3 3 9 9 3 13 0 9 9 9 7 9 9 9 2
17 13 3 9 0 13 0 1 0 13 7 10 9 3 13 10 9 2
9 3 3 10 0 13 1 10 9 2
17 13 3 1 10 9 10 13 1 15 13 7 10 13 10 9 13 2
15 0 3 10 9 13 13 10 9 10 0 13 1 10 9 2
17 1 13 3 3 9 1 9 13 0 9 9 9 7 9 9 9 2
17 1 3 15 9 10 10 9 9 13 1 9 13 10 10 9 9 2
13 1 3 15 13 1 9 0 10 9 13 10 9 2
23 1 3 15 13 9 10 0 9 1 10 9 13 0 0 9 15 7 10 10 9 9 13 2
24 9 3 3 13 10 13 9 16 13 0 2 3 3 0 10 9 13 1 10 15 13 13 15 2
18 0 3 13 9 10 10 0 9 16 13 1 0 0 9 13 10 13 2
12 15 3 10 9 13 10 1 10 9 9 13 2
11 3 15 13 10 13 10 9 9 0 13 2
14 3 3 10 10 9 9 10 13 1 10 9 0 13 2
18 13 3 3 10 9 1 9 0 13 7 9 7 10 0 9 3 13 2
20 13 3 10 9 0 1 10 10 9 9 7 1 10 9 10 9 0 13 9 2
11 1 15 10 1 9 13 1 10 0 9 2
10 3 10 3 1 10 9 1 15 13 2
9 0 3 13 9 0 10 9 13 2
12 13 3 10 9 9 0 3 13 1 10 9 2
12 1 15 10 1 9 13 13 1 10 13 9 2
14 1 13 3 3 9 9 13 0 9 9 7 9 9 2
14 15 3 13 1 10 9 13 10 9 13 1 10 9 2
19 0 3 3 10 13 13 13 13 16 0 7 1 10 13 10 13 13 9 2
13 10 3 9 16 0 0 9 13 3 13 10 9 2
14 9 3 9 13 3 9 0 0 13 1 9 0 9 2
20 0 3 9 9 0 2 3 9 9 0 1 0 13 2 1 9 0 13 3 2
31 3 3 9 0 2 9 9 3 0 3 9 0 9 13 2 13 2 3 3 9 2 15 9 13 2 13 9 15 0 13 2
11 9 3 13 0 9 3 2 9 3 13 2
29 15 13 2 3 1 0 9 0 9 10 3 9 13 2 15 3 3 13 0 9 0 2 15 3 0 3 13 13 2
7 13 3 9 15 1 9 2
18 9 7 0 13 13 1 9 2 9 3 3 13 2 13 3 0 9 2
6 3 3 13 3 3 2
6 9 9 3 0 13 2
11 3 3 13 1 9 0 1 9 9 9 2
10 0 3 9 0 3 13 9 13 0 2
13 13 3 9 1 0 0 9 2 9 3 0 13 2
11 13 15 9 3 3 13 3 9 1 0 2
9 3 3 13 1 9 0 0 9 2
5 3 15 9 13 2
9 3 3 13 1 9 0 0 9 2
15 9 3 3 0 3 9 9 13 9 0 15 13 1 9 2
4 3 3 13 2
10 9 3 1 9 9 15 9 0 13 2
6 13 3 9 9 0 2
7 0 3 1 9 13 9 2
6 3 3 3 13 13 2
12 7 1 9 3 9 13 13 13 0 9 13 2
5 9 3 13 0 2
13 9 3 9 7 0 13 2 1 9 0 3 9 2
12 3 3 1 15 15 9 9 9 13 9 13 2
21 9 3 13 0 3 10 7 0 2 10 7 0 3 1 0 13 9 9 1 0 2
10 7 7 0 3 3 0 1 9 13 2
4 13 3 13 2
5 0 13 9 9 2
7 13 3 3 13 10 0 2
8 13 3 15 13 15 0 9 2
5 9 3 9 13 2
6 13 3 0 1 9 2
8 13 3 3 15 3 9 13 2
9 7 3 13 2 9 3 13 9 2
6 0 13 3 13 15 2
7 7 9 9 15 3 13 2
7 13 3 9 15 13 9 2
6 13 3 7 13 0 2
7 15 3 13 15 9 3 2
6 13 9 15 9 9 2
9 3 3 3 13 3 3 13 9 2
5 0 3 0 13 2
7 0 3 9 15 9 13 2
7 9 9 3 3 13 13 2
11 3 3 3 13 0 0 1 0 13 3 2
14 3 13 9 2 3 9 2 9 0 1 13 0 9 2
15 13 2 13 15 10 9 2 16 3 15 9 3 13 15 2
14 9 3 3 3 1 9 9 13 1 15 1 9 0 2
7 0 15 9 9 13 9 2
16 7 0 0 3 13 0 13 2 16 7 13 9 13 10 13 2
6 13 1 9 0 9 2
17 15 3 1 15 0 3 9 13 2 7 9 0 2 7 9 9 2
8 1 0 13 7 13 0 15 2
11 15 3 9 3 0 9 9 15 13 9 2
17 7 0 9 2 15 7 0 13 9 2 10 1 13 9 2 13 2
6 13 3 9 0 9 2
5 15 1 15 13 2
12 0 3 9 0 9 15 3 13 9 9 9 2
17 0 9 0 7 0 13 3 9 0 9 9 3 0 13 1 9 2
14 13 3 3 1 15 9 9 3 3 13 7 13 3 2
9 0 3 3 3 9 3 13 9 2
7 7 0 0 0 13 9 2
9 0 3 3 0 9 13 3 0 2
19 7 9 3 13 0 0 2 0 9 3 1 0 9 13 13 9 1 9 2
16 7 10 0 0 3 9 2 16 0 13 2 3 3 13 15 2
9 13 3 3 2 7 9 0 13 2
7 3 3 13 9 9 15 2
7 9 10 9 13 0 9 2
7 3 13 9 1 0 9 2
7 13 2 9 0 9 9 2
7 10 0 13 9 13 9 2
5 0 9 0 13 2
7 15 3 13 0 0 0 2
7 9 13 0 15 9 3 2
8 3 15 1 9 13 0 9 2
7 7 0 13 0 3 15 2
7 7 3 9 1 9 13 2
8 7 9 3 9 9 13 9 2
8 15 3 10 9 9 13 9 2
8 15 3 3 0 15 9 13 2
8 10 0 3 9 0 15 13 2
7 7 15 13 9 0 9 2
12 9 3 0 0 9 13 3 16 0 13 9 2
8 13 3 15 15 13 9 0 2
7 3 3 0 9 13 13 2
4 0 13 9 2
8 9 3 13 3 0 0 9 2
12 15 13 13 15 0 9 2 0 13 0 9 2
10 0 1 9 2 7 15 7 9 13 2
8 15 3 3 0 13 10 13 2
7 9 3 3 0 13 9 2
8 3 3 1 15 0 15 13 2
7 3 10 9 3 0 13 2
6 13 13 15 9 0 2
10 13 9 0 0 13 9 15 0 9 2
7 13 3 0 9 0 0 2
9 3 3 1 0 0 9 9 13 2
6 15 3 3 13 9 2
9 13 3 0 9 0 9 9 0 2
6 3 13 9 0 0 2
13 10 0 3 16 13 9 2 0 13 9 13 9 2
15 15 3 3 3 13 9 3 2 9 3 0 15 13 1 2
22 9 0 13 2 13 9 2 0 9 2 0 9 15 2 0 3 1 9 9 0 13 2
3 9 13 2
15 9 3 13 10 0 0 2 15 3 13 3 13 9 1 2
9 13 3 9 0 9 0 13 9 2
20 16 3 13 9 9 15 9 9 2 13 3 9 13 2 15 3 15 13 13 2
17 13 3 15 13 1 9 10 3 2 16 3 13 9 0 1 15 2
9 7 15 3 3 13 0 9 9 2
9 0 3 3 9 13 9 0 9 2
10 0 3 13 9 13 9 10 1 9 2
5 7 15 13 0 2
17 0 0 15 13 9 0 2 13 3 0 3 0 2 0 3 0 2
7 3 3 13 13 9 0 2
7 13 7 13 3 0 9 2
8 13 3 9 9 7 13 9 2
20 7 15 13 10 9 13 1 9 9 9 13 3 9 2 0 9 3 9 0 2
3 13 3 2
15 9 15 7 9 2 0 3 13 2 13 3 13 0 9 2
6 15 13 0 3 9 2
4 7 3 13 2
4 3 3 13 2
19 7 15 7 15 9 13 0 0 13 9 2 7 13 9 9 0 3 13 2
15 3 3 9 15 1 13 13 3 9 3 16 0 0 13 2
7 13 3 3 1 9 0 2
6 0 13 9 0 9 2
6 13 2 7 13 3 2
4 3 15 13 2
7 3 3 9 0 0 13 2
7 13 0 9 15 13 13 2
6 15 15 13 9 9 2
4 3 3 13 2
5 13 9 9 9 2
2 13 2
4 13 3 0 2
13 7 3 3 0 9 2 0 3 9 9 3 13 2
14 9 3 0 9 3 3 0 15 13 2 3 9 0 2
14 16 3 3 15 7 15 13 9 2 9 13 3 0 2
21 7 3 3 3 15 13 13 15 9 3 13 9 9 2 15 3 3 13 9 0 2
8 10 0 3 0 15 9 13 2
27 9 3 9 3 0 13 2 16 3 10 0 9 9 0 7 2 0 9 13 2 9 3 13 1 9 13 2
8 9 3 3 0 9 9 13 2
6 13 7 9 13 9 2
8 7 3 0 15 13 9 1 2
6 3 3 10 9 13 2
8 0 3 13 2 7 13 13 2
5 15 3 3 13 2
5 3 9 13 15 2
9 7 3 15 13 9 7 9 15 2
7 0 1 9 3 13 15 2
8 7 3 0 9 3 13 15 2
6 3 0 9 15 13 2
5 0 13 9 13 2
7 3 3 0 13 13 0 2
7 3 0 0 9 13 9 2
14 15 3 9 13 0 13 2 10 0 16 3 0 13 2
8 7 0 13 9 0 13 13 2
14 1 0 13 7 9 0 9 13 15 15 9 13 13 2
6 15 3 0 13 13 2
7 9 3 13 7 9 0 2
8 9 3 13 0 10 0 9 2
10 0 3 9 13 13 9 1 15 0 2
9 13 3 0 1 9 0 9 3 2
4 9 3 13 2
10 13 3 9 0 0 9 13 9 0 2
13 3 0 13 9 2 2 0 9 15 9 13 3 2
12 9 15 9 7 15 3 9 13 1 9 13 2
9 15 3 9 0 13 3 1 9 2
11 1 9 3 3 15 13 10 0 0 13 2
6 0 3 13 13 9 2
12 13 3 9 3 9 13 15 15 0 13 9 2
5 9 13 0 9 2
12 13 0 3 3 2 3 3 13 15 0 9 2
10 9 3 9 0 13 9 15 13 9 2
12 0 13 9 0 9 13 1 9 16 13 15 2
8 0 3 13 0 9 9 9 2
4 9 3 13 9
4 0 3 13 2
7 13 3 9 9 9 0 2
9 3 3 0 9 9 13 9 9 2
19 3 9 3 13 0 0 13 2 10 0 3 3 2 15 0 9 9 13 2
19 3 3 15 9 9 13 15 9 13 2 0 9 0 9 9 3 0 13 2
9 9 3 9 1 9 13 9 0 2
9 0 3 3 9 13 9 9 0 2
7 0 3 9 9 0 13 2
7 10 0 3 1 9 13 2
8 0 3 1 9 9 13 9 2
13 9 3 0 2 3 13 9 2 9 1 9 13 2
14 9 3 2 15 9 13 3 13 0 0 0 0 9 2
12 10 3 13 9 0 15 1 0 9 13 0 2
12 15 3 7 13 13 9 0 15 7 0 9 2
9 0 3 15 1 9 13 10 9 2
6 0 3 3 15 13 2
10 0 3 9 1 9 13 9 3 13 2
13 3 3 13 7 13 1 9 13 15 7 13 9 2
8 15 3 0 9 3 13 13 2
14 3 3 3 9 15 7 9 13 2 13 13 9 9 2
5 3 0 13 15 2
4 7 13 15 2
2 13 2
13 9 3 9 3 1 9 9 13 15 9 13 9 2
12 0 15 13 9 3 0 9 9 16 15 15 2
9 0 13 0 9 9 9 3 0 2
5 7 13 1 13 2
14 0 3 13 9 9 13 3 0 9 0 0 1 9 2
11 0 3 3 13 1 9 13 9 3 13 2
5 0 3 7 13 2
4 3 13 9 2
9 3 13 9 10 9 0 9 13 2
7 9 3 9 3 13 9 2
38 3 0 0 9 9 2 3 3 9 2 3 13 9 0 1 9 13 2 3 3 1 9 13 9 9 3 2 3 3 7 13 0 9 1 9 13 9 2
7 13 9 13 9 9 0 2
15 3 13 3 3 3 3 9 9 0 2 3 9 9 13 2
12 9 3 3 13 9 9 2 13 3 0 9 2
12 3 13 0 9 2 0 16 15 9 13 3 2
7 0 13 9 9 13 9 2
12 10 0 3 0 0 0 3 9 1 9 13 2
7 0 3 3 3 13 0 2
6 9 3 13 15 9 2
6 9 9 3 15 13 2
3 13 9 2
16 13 3 3 0 9 13 1 9 2 3 9 0 15 13 9 2
6 1 13 3 9 13 2
11 9 3 3 9 0 9 9 3 13 13 2
8 9 0 3 9 13 9 9 2
17 9 3 0 9 0 0 1 15 9 13 9 9 0 0 13 13 2
8 15 3 1 15 0 0 13 2
5 13 9 1 9 2
14 7 1 0 0 9 0 1 9 2 0 3 9 13 2
7 13 9 2 13 1 9 2
5 0 9 3 13 2
13 3 3 13 0 9 2 3 13 0 9 9 13 2
16 15 3 1 9 9 13 3 0 0 2 9 9 3 0 0 2
16 6 3 3 13 7 0 9 2 1 0 9 0 13 0 9 2
7 13 7 13 7 13 9 2
6 0 3 9 3 13 2
9 13 7 13 2 13 0 9 9 2
8 13 13 9 1 0 0 0 2
5 3 3 15 13 2
7 9 3 3 9 0 13 2
6 3 13 9 3 3 2
6 3 13 9 10 3 2
10 3 3 15 13 2 3 3 13 9 2
5 13 3 9 9 2
9 9 3 3 15 15 9 13 13 2
15 16 7 15 1 9 13 13 15 2 9 9 9 3 13 2
2 13 2
6 13 2 3 13 9 2
14 13 13 15 13 9 2 16 3 13 0 10 0 9 2
9 1 0 9 9 9 15 13 9 2
8 3 3 9 1 9 13 13 2
7 0 13 3 9 13 3 2
7 7 0 13 0 13 9 2
8 15 3 13 15 15 9 1 2
7 0 3 13 0 3 13 2
5 0 13 13 13 2
7 9 13 10 9 0 13 2
6 10 1 9 9 13 2
11 13 3 2 16 13 2 3 3 1 0 2
6 13 9 3 3 0 2
7 3 3 13 10 9 9 2
7 13 3 13 9 9 15 2
7 3 13 0 9 1 9 2
9 3 0 13 3 9 9 9 9 2
6 15 15 13 13 9 2
11 1 9 13 13 15 3 0 10 9 15 2
15 0 3 0 3 1 9 9 13 3 2 16 0 13 9 2
10 15 13 3 9 3 2 16 13 3 2
19 0 3 9 13 13 3 3 1 9 9 13 2 0 3 13 1 0 9 2
7 13 3 3 0 1 9 2
6 13 3 9 13 0 2
8 13 3 9 7 9 10 9 2
13 3 9 3 15 9 9 13 3 13 1 9 9 2
10 3 15 13 0 13 9 0 1 0 2
12 16 3 15 0 9 2 13 13 7 0 9 2
5 15 15 0 13 2
5 13 3 10 0 2
16 0 3 1 9 9 0 13 0 2 10 3 13 0 9 3 2
13 0 3 13 7 13 15 2 9 13 15 0 9 2
9 9 3 13 7 9 2 15 3 2
25 1 0 7 13 15 0 9 0 3 9 7 13 9 2 3 3 9 15 2 9 3 0 0 13 2
19 9 3 7 0 1 15 3 9 2 15 3 7 9 13 2 13 9 1 2
13 0 13 15 9 9 2 10 13 13 10 9 0 2
6 0 13 1 9 0 2
15 16 3 15 7 9 13 0 2 9 10 3 3 13 9 2
15 13 3 9 9 9 13 0 3 7 15 9 9 13 0 2
15 9 3 9 15 9 13 2 3 3 3 9 9 13 9 2
15 13 3 9 0 9 13 2 3 3 1 9 9 13 9 2
5 0 13 15 9 2
8 13 3 9 9 9 1 9 2
14 0 3 0 9 13 9 15 3 0 0 13 9 9 2
10 13 3 9 9 9 0 9 3 9 2
11 9 3 9 0 3 9 9 3 0 13 2
7 15 1 9 13 0 9 2
10 15 15 3 0 13 2 15 13 3 2
8 9 3 0 13 0 9 0 2
10 1 0 3 9 15 9 0 13 9 2
8 10 0 9 13 9 0 15 2
6 15 3 3 0 13 2
6 15 3 13 3 0 2
8 15 3 3 3 13 10 13 2
5 0 3 9 13 2
5 0 9 15 13 2
31 15 3 9 10 13 9 1 9 9 13 2 7 10 0 7 0 9 9 2 1 9 15 0 9 9 9 0 13 9 13 2
15 1 3 9 10 0 7 0 9 3 9 3 13 9 3 2
23 0 3 9 0 13 2 0 3 9 13 2 3 15 9 3 3 15 9 9 10 9 13 2
9 0 3 10 0 7 0 9 13 2
17 9 3 10 0 0 9 13 3 2 9 3 0 7 0 9 0 2
13 10 0 3 9 1 0 9 13 0 9 1 9 2
26 15 9 9 9 13 9 2 15 1 0 9 0 13 9 13 0 2 9 3 9 3 3 13 9 13 2
16 0 3 13 9 1 9 9 2 3 3 13 1 15 0 13 2
7 9 3 9 9 13 9 2
12 0 9 9 10 13 2 7 0 9 9 13 2
2 13 2
20 9 3 9 9 2 9 3 7 9 13 2 16 15 7 9 0 3 13 9 2
14 0 3 13 13 0 9 7 10 9 3 0 0 9 2
5 15 9 13 9 2
11 13 3 9 3 0 2 1 3 9 9 2
7 9 3 9 13 9 9 2
10 0 3 10 0 1 15 13 15 9 2
8 0 3 13 15 15 9 13 2
19 0 3 3 0 9 13 2 1 15 9 0 13 9 9 9 13 13 13 2
11 3 3 3 15 0 13 3 10 1 9 2
4 13 3 15 2
18 9 3 0 13 13 13 2 9 3 1 13 0 7 9 1 9 13 2
31 15 3 15 13 9 1 9 3 13 0 9 2 15 3 13 2 7 9 9 9 13 7 13 9 1 9 7 9 13 0 2
12 13 3 0 9 2 7 9 13 9 13 15 2
25 16 3 13 7 9 0 13 9 2 1 0 9 9 13 2 0 9 13 13 9 2 15 9 15 2
8 13 3 13 9 1 9 9 2
12 0 3 9 13 9 9 13 7 9 9 13 2
29 3 3 13 2 9 0 13 3 3 0 3 13 9 2 3 3 13 2 3 0 9 2 13 3 3 15 13 9 2
31 9 3 9 13 2 16 15 0 13 2 13 15 9 13 2 10 3 0 0 13 15 3 7 9 15 7 9 0 3 0 2
10 0 3 13 9 9 3 7 0 13 2
7 0 0 13 15 3 13 2
9 3 3 3 13 15 15 13 1 2
17 3 3 0 3 10 0 15 0 9 9 7 9 0 15 13 9 2
5 13 3 10 0 2
21 0 3 2 3 13 2 0 13 9 10 3 1 9 0 2 16 3 1 9 13 2
9 3 3 13 0 9 15 13 9 2
8 0 3 13 3 9 9 0 2
7 3 15 13 0 9 9 2
8 0 9 13 9 3 3 0 2
8 3 3 3 13 9 0 9 2
8 0 3 13 13 10 13 13 2
9 3 15 13 3 13 0 0 9 2
18 15 3 9 9 0 13 13 2 7 13 0 15 9 0 7 0 13 2
6 9 3 0 13 0 2
7 0 3 3 0 13 9 2
14 3 0 15 3 15 9 13 0 2 13 15 9 0 2
11 13 0 3 13 9 9 0 3 0 9 2
12 0 3 13 9 2 0 3 13 9 13 0 9
12 13 0 9 0 9 0 2 16 0 3 13 2
12 13 3 1 7 0 9 3 13 9 7 0 2
6 13 3 0 13 0 2
11 13 3 15 9 15 3 13 0 13 9 2
12 0 3 13 9 13 13 2 16 13 0 7 2
20 15 3 13 2 15 3 7 13 10 0 2 15 1 9 13 0 9 13 13 2
9 9 3 0 13 3 7 13 9 2
13 0 3 13 9 9 0 7 0 9 9 1 0 2
11 10 9 9 9 9 9 0 1 9 13 2
15 7 9 0 2 9 3 0 2 0 9 9 2 3 13 2
6 15 9 3 13 1 2
7 0 13 3 0 13 0 2
7 3 13 15 0 13 3 2
16 0 3 9 13 9 9 2 3 13 0 9 9 13 0 9 2
10 9 3 3 3 13 3 0 9 13 2
4 3 13 9 2
7 7 15 13 3 13 13 2
13 3 3 9 15 13 9 2 9 13 3 0 9 2
6 9 9 13 9 9 2
7 3 3 9 13 0 9 2
7 9 3 13 9 13 0 2
9 9 3 9 9 0 13 2 13 2
16 15 13 2 0 9 2 9 2 7 9 0 2 9 13 9 2
19 7 16 9 13 9 0 2 9 3 9 13 15 2 9 13 9 13 13 2
7 0 13 3 1 0 9 2
8 3 3 10 13 1 9 13 2
21 15 3 3 3 2 3 0 9 9 3 13 2 9 3 9 13 9 9 1 0 2
21 16 3 9 9 13 7 9 13 2 0 9 9 9 1 9 13 0 3 9 9 2
7 9 3 9 13 9 0 2
18 13 3 3 0 13 13 2 7 0 3 0 13 9 9 0 0 9 2
13 7 9 13 2 3 3 9 9 0 9 0 13 2
28 16 3 3 0 9 0 13 9 0 13 2 0 3 9 9 9 1 3 13 2 0 3 3 13 9 9 9 2
8 9 3 0 0 13 9 13 2
17 3 3 7 9 9 13 0 9 3 2 3 1 9 13 0 9 2
7 9 3 9 0 0 13 2
18 3 3 9 9 9 13 9 0 1 9 2 3 3 0 13 0 13 2
14 7 3 1 15 9 9 9 13 2 3 13 13 9 2
19 13 3 9 0 9 2 13 0 9 9 9 2 1 0 3 0 13 9 2
9 10 0 3 3 9 0 9 13 2
19 9 3 0 9 3 13 2 9 3 0 0 9 13 2 0 13 0 9 2
14 9 3 3 9 13 0 9 2 16 0 9 9 13 2
17 0 3 9 2 3 3 3 16 12 9 13 2 3 3 13 15 2
13 15 1 0 13 9 9 16 15 7 3 13 9 2
9 7 0 13 3 15 3 0 9 2
14 13 0 3 13 15 9 9 13 0 13 1 10 0 2
25 9 0 13 0 9 2 9 3 0 9 0 2 0 3 9 9 1 0 3 2 13 3 0 9 2
7 0 9 3 15 13 13 2
22 9 15 13 3 9 9 2 0 2 0 9 2 15 10 0 9 13 2 0 9 1 2
29 3 13 15 2 16 2 16 9 13 0 9 13 2 13 0 9 9 2 0 3 13 0 9 2 3 10 13 13 2
17 16 3 9 9 13 9 9 9 2 3 13 0 9 9 9 13 2
11 1 3 13 0 9 2 3 13 3 13 2
16 0 3 3 1 9 9 13 2 0 3 1 9 9 13 13 2
17 9 3 13 1 9 9 13 2 13 0 9 2 16 0 13 9 2
7 9 3 13 0 13 9 2
16 13 3 9 13 0 2 0 13 3 9 2 13 0 1 9 2
9 15 15 1 15 1 9 1 13 2
17 0 3 9 0 9 0 9 13 2 3 13 15 3 9 0 13 2
11 15 9 9 0 13 13 15 9 9 13 2
13 15 3 13 2 9 15 13 9 2 3 15 13 2
4 13 13 3 2
13 9 3 9 10 13 3 1 9 3 0 13 9 2
12 3 15 9 9 9 7 0 9 13 0 13 2
5 0 3 13 15 2
16 9 3 1 0 9 9 0 13 2 13 3 0 9 0 9 2
16 9 3 15 10 3 13 3 3 13 9 2 9 9 3 13 2
12 16 3 0 13 13 9 2 13 9 1 9 2
12 15 3 15 3 13 9 9 13 2 13 13 2
13 13 3 9 0 9 9 0 9 13 2 13 9 2
5 13 3 1 0 2
9 13 3 3 15 0 9 13 9 2
23 0 3 0 13 9 2 9 13 3 0 9 2 13 13 2 3 0 15 2 1 0 9 2
4 0 13 0 2
10 0 3 13 13 0 15 9 13 9 2
7 15 3 3 0 3 13 2
15 7 3 2 16 3 13 9 15 2 9 3 0 13 13 2
25 7 9 2 16 3 3 15 3 13 2 13 2 7 13 1 9 2 16 7 15 1 0 13 0 2
14 0 3 0 9 9 13 0 9 9 13 2 9 13 2
9 15 3 9 10 13 13 3 0 2
10 3 3 3 0 3 13 9 9 13 2
13 0 3 13 9 0 13 9 1 0 0 3 9 2
7 13 3 0 9 0 9 2
23 15 3 1 9 9 3 3 13 2 3 3 3 13 0 9 2 3 3 1 9 13 13 2
5 0 3 13 9 2
11 13 3 9 0 13 2 16 13 9 9 2
10 13 3 9 9 0 9 13 10 9 2
21 15 3 3 0 3 9 0 1 9 0 13 9 2 13 3 1 9 9 3 9 2
6 0 0 9 13 9 2
14 16 3 15 0 9 13 0 2 0 3 0 9 13 2
5 1 3 13 15 2
9 13 3 3 0 3 9 9 13 2
5 0 3 13 13 2
16 13 1 9 9 9 2 0 9 9 13 2 0 9 0 13 2
7 0 3 15 1 9 13 2
7 9 3 3 1 0 13 2
9 0 9 15 13 0 9 0 0 2
8 13 2 13 2 7 13 9 2
14 13 3 9 10 0 9 3 13 2 9 3 0 13 2
7 7 3 0 13 15 13 2
7 13 3 16 0 13 9 2
7 15 13 9 0 0 0 2
13 13 3 13 2 13 3 9 13 15 0 1 9 2
13 13 3 13 2 13 3 9 13 2 13 0 0 2
9 0 3 3 3 9 3 13 9 2
9 13 10 9 9 2 16 13 9 2
8 9 15 13 9 7 9 9 2
7 3 1 9 0 13 9 2
7 15 3 0 3 9 13 2
2 13 2
9 0 7 9 3 9 15 13 0 2
6 0 9 13 12 9 2
9 3 3 7 9 15 0 13 13 2
9 9 13 9 9 2 3 13 9 2
9 7 15 13 2 3 9 13 0 2
3 3 13 2
7 9 3 3 15 9 13 2
8 7 15 3 13 0 3 13 2
7 0 9 13 0 13 9 2
8 3 3 3 9 0 13 9 2
11 0 3 13 0 9 2 3 3 15 9 2
9 0 3 9 0 13 3 0 13 2
11 15 3 3 1 0 9 15 13 13 9 2
10 3 16 13 15 0 2 10 9 13 2
8 3 0 13 9 0 13 0 2
10 9 3 0 15 3 13 13 0 9 2
9 3 15 3 9 9 13 9 0 2
12 13 16 0 9 9 0 9 13 15 13 9 2
9 0 3 0 13 9 13 0 9 2
25 13 3 16 15 3 0 9 9 13 1 9 2 15 3 9 1 3 13 2 0 3 9 0 13 2
15 15 1 9 9 3 13 0 15 13 9 7 9 1 9 2
8 9 3 13 10 0 9 9 2
8 0 3 0 9 15 9 13 2
6 9 3 0 9 13 2
13 0 3 9 7 9 13 2 9 3 0 13 9 2
9 9 3 3 13 2 16 0 13 2
7 9 3 9 0 13 9 2
19 15 3 1 9 9 13 0 1 9 2 1 9 0 2 15 15 13 9 2
7 3 3 0 15 13 9 2
11 3 3 1 0 3 13 7 0 0 9 2
8 0 3 10 9 0 0 13 2
9 3 0 13 2 15 9 3 13 2
7 3 0 3 0 13 9 2
14 3 3 3 10 13 3 1 9 9 9 13 0 9 2
3 3 13 2
12 3 3 0 9 0 13 10 9 9 9 1 2
10 13 3 3 15 3 2 15 3 3 2
12 16 15 13 2 9 0 9 13 0 9 13 2
14 15 9 13 9 3 9 9 13 13 3 3 13 9 2
12 9 3 0 2 9 3 9 0 3 13 9 2
12 0 3 13 9 0 1 9 9 9 9 1 2
18 9 0 3 7 0 9 0 13 9 9 16 3 3 0 13 13 13 2
12 9 3 13 13 9 9 2 3 0 13 9 2
22 0 13 15 9 13 9 9 3 2 3 3 15 13 10 13 9 0 13 9 13 0 2
16 1 0 0 2 13 13 2 13 0 9 2 13 13 0 9 2
12 0 3 0 1 9 9 1 9 13 0 9 2
8 15 3 13 9 1 9 3 2
12 3 0 7 13 7 13 3 13 13 0 9 2
13 3 13 2 7 13 9 1 9 13 9 15 13 2
8 3 3 10 0 1 0 13 2
12 7 10 0 1 9 0 0 9 13 0 9 2
10 0 3 13 9 9 9 0 3 9 2
14 3 3 3 3 0 15 3 13 9 13 3 9 0 2
10 13 3 15 9 9 15 9 13 9 2
12 9 3 13 10 0 9 9 13 9 9 9 2
7 13 0 7 0 0 9 2
17 13 3 15 0 2 0 9 3 13 0 3 9 2 9 9 9 2
6 13 13 3 9 0 2
15 9 3 13 2 9 0 9 0 0 9 13 0 3 9 2
14 0 13 0 1 9 13 1 9 0 0 13 1 9 2
4 15 15 13 2
29 3 7 10 9 3 10 0 0 0 9 0 0 9 9 9 9 10 9 10 9 2 9 3 0 3 9 13 13 2
6 9 0 0 0 13 2
7 13 13 15 9 3 9 2
10 13 13 2 3 1 9 0 3 13 2
6 13 3 15 9 9 2
2 13 2
5 13 3 15 9 2
8 13 10 0 15 10 0 9 2
3 13 13 2
5 15 15 13 13 2
3 13 0 2
5 13 0 13 9 2
7 9 3 13 1 9 0 2
12 0 3 13 7 0 2 0 2 9 3 0 2
4 13 13 9 2
5 1 9 3 13 2
5 13 3 0 15 2
5 13 9 3 13 2
7 13 13 7 13 0 9 2
4 13 0 13 2
5 13 3 0 15 2
4 13 3 9 2
7 7 9 13 13 10 0 2
7 7 15 9 13 0 9 2
4 13 3 0 2
4 7 15 13 2
7 9 3 13 9 13 9 2
7 7 13 9 7 13 9 2
4 13 3 9 2
3 13 3 2
5 13 3 0 15 2
5 0 1 9 13 2
6 13 3 15 0 9 2
22 15 3 9 15 13 9 13 9 2 16 3 13 10 9 9 13 2 0 3 13 9 2
12 15 3 0 13 0 9 13 9 9 1 0 2
16 0 3 15 10 0 9 13 9 2 9 3 0 9 13 3 2
9 3 3 10 13 9 0 13 15 2
7 10 13 3 3 13 3 2
6 0 13 10 0 9 2
12 9 9 3 3 13 9 9 9 13 1 9 2
14 1 15 0 15 13 9 3 2 0 2 3 13 9 2
8 0 3 9 7 9 0 13 2
15 15 10 9 0 3 13 9 2 15 10 0 0 13 9 2
2 13 2
5 3 0 13 0 2
4 15 15 13 2
7 3 15 0 0 13 13 2
7 0 3 0 13 1 9 2
6 13 15 0 13 13 2
13 3 13 15 9 13 2 16 7 15 13 13 9 2
7 7 3 0 9 13 1 2
13 13 15 1 9 0 9 9 13 2 13 1 9 2
7 13 3 3 13 9 15 2
8 13 3 2 13 2 3 13 2
6 13 15 3 9 3 2
13 7 15 3 13 3 2 16 13 9 13 9 0 2
8 1 15 3 0 3 13 15 2
10 0 3 9 0 9 9 3 13 3 2
11 15 3 3 13 10 9 3 0 1 13 2
5 13 9 0 9 2
6 13 13 15 10 0 2
6 3 1 9 9 13 2
7 3 3 13 13 3 1 2
8 13 3 2 9 3 13 9 2
8 7 3 13 9 3 0 9 2
6 3 3 13 0 9 2
6 0 9 9 15 13 2
7 13 2 16 9 9 13 2
10 3 3 13 7 9 9 13 0 13 2
6 3 15 9 9 13 2
12 0 3 15 13 9 2 15 9 15 13 9 2
28 6 0 9 7 0 9 2 9 3 9 2 0 3 9 0 9 2 9 3 9 2 7 10 9 9 9 13 2
9 13 0 9 13 10 0 9 13 2
11 15 10 0 9 9 13 1 15 9 0 2
4 3 15 13 2
14 0 13 3 15 13 2 3 3 15 0 9 0 13 2
18 10 13 3 13 9 13 3 0 2 13 16 10 10 9 13 0 9 2
15 3 3 3 13 3 3 7 13 9 0 3 15 15 13 2
9 0 3 9 13 9 15 13 0 2
17 0 3 13 9 9 0 2 15 9 9 0 9 13 7 0 9 2
8 15 9 9 13 0 9 13 2
13 13 0 1 9 9 0 9 2 7 15 3 13 2
8 9 9 11 11 9 11 9 11
4 11 13 10 11
5 11 3 13 10 11
9 11 3 13 10 11 7 10 9 15
11 11 3 13 10 11 7 10 11 1 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
8 11 3 13 10 11 1 10 11
8 11 3 13 10 11 1 10 11
5 11 3 13 10 11
7 11 3 13 10 11 10 9
9 11 3 13 10 11 1 10 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
13 11 3 13 10 11 7 10 9 15 1 10 9 11
9 1 3 10 9 11 11 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
29 15 3 10 9 1 11 1 11 9 12 7 1 11 1 10 9 11 9 12 7 1 10 9 11 1 10 11 9 12
8 10 3 11 11 10 9 3 13
18 13 10 9 15 11 10 11 16 3 13 15 13 1 9 13 1 9 0
16 11 3 10 9 15 0 13 7 3 13 15 13 13 3 13 15
10 11 9 11 3 13 13 11 10 9 15
9 10 3 1 15 13 1 9 13 0
19 13 3 9 7 13 10 9 15 11 15 3 13 10 9 15 1 10 9 15
14 0 3 0 13 16 13 10 13 1 9 1 10 9 13
18 13 3 11 1 10 9 13 3 13 15 10 9 9 7 13 10 9 15
8 7 3 13 15 16 15 13 9
6 7 13 10 9 15 11
7 3 13 10 13 9 10 0
12 13 3 15 10 9 1 10 9 7 13 13 15
27 13 3 10 9 11 13 7 15 11 1 15 7 13 15 10 9 7 9 10 9 13 1 15 3 10 11 13
4 15 3 13 15
4 1 11 10 11
12 7 15 11 9 11 3 0 13 1 10 9 11
12 1 15 3 13 13 15 13 10 9 15 10 11
6 13 13 3 1 10 9
11 16 3 13 13 15 16 3 15 13 13 15
25 15 3 13 10 9 13 7 6 10 9 15 13 1 10 9 13 15 16 13 13 1 3 13 10 9
8 13 3 10 9 13 9 0 3
30 7 13 1 10 9 13 10 9 1 11 10 9 15 7 13 13 15 7 13 10 9 15 13 15 9 9 7 9 7 9
16 7 13 1 9 3 13 1 11 1 0 9 13 1 10 9 15
19 13 13 10 9 7 10 9 15 7 13 1 11 7 13 3 16 3 13 15
32 15 3 13 13 10 9 7 10 9 15 9 7 13 1 11 7 13 3 1 10 9 11 16 13 10 13 1 9 1 10 9 13
6 1 11 13 10 9 15
37 3 11 13 16 13 1 10 9 13 3 7 13 13 15 10 9 10 1 11 7 1 15 10 9 15 1 0 7 3 1 10 9 15 13 1 10 9
9 3 13 10 13 1 11 10 9 13
8 9 1 11 13 9 7 9 0
12 11 13 10 9 15 7 3 13 13 16 3 13
15 13 3 10 11 6 9 9 13 1 9 10 11 1 11 13
15 13 3 16 11 13 10 11 1 10 9 15 11 13 3 13
10 13 3 1 9 13 1 10 9 10 11
17 7 13 13 1 9 13 11 16 13 10 13 1 10 9 16 0 13
16 1 3 10 9 0 13 11 10 9 13 1 10 0 10 11 13
1 13
6 13 3 10 9 10 9
10 0 3 13 10 13 1 11 10 9 13
5 9 13 1 10 0
5 0 13 10 9 15
18 0 3 10 11 13 10 9 15 1 9 9 7 9 0 1 10 9 15
9 10 3 9 13 15 9 7 9 0
27 3 13 1 15 11 7 15 10 11 7 15 10 9 10 11 7 13 1 10 11 9 1 15 13 10 9 15
13 13 3 0 10 9 7 9 13 1 10 9 13 15
10 9 9 15 13 15 13 1 10 13 9
6 13 3 9 0 10 9
6 7 3 13 13 1 15
10 3 3 10 9 1 10 9 10 9 13
12 15 3 9 3 13 9 0 13 7 1 9 13
8 15 3 15 13 1 9 1 9
15 10 3 1 15 13 0 15 13 15 3 13 0 10 9 13
8 0 15 13 1 9 0 7 9
20 15 10 9 1 10 9 15 7 13 10 9 15 7 13 10 9 15 1 10 9
6 10 3 9 13 9 0
5 15 3 13 15 13
7 13 3 10 11 13 1 15
2 13 3
8 3 3 13 13 15 13 15 9
3 3 13 15
9 13 3 10 11 3 13 1 10 9
15 7 6 13 10 9 7 13 9 9 13 3 9 13 1 15
10 0 13 10 9 15 10 0 1 15 13
14 3 10 11 13 1 10 9 1 10 9 13 1 10 9
6 7 13 10 13 13 15
12 16 9 13 10 9 13 16 10 9 0 9 13
4 15 3 13 13
1 13
15 3 1 9 0 13 10 9 7 1 15 9 13 1 9 9
8 16 9 13 10 9 13 15 3
3 13 3 16
18 10 9 15 13 1 15 7 1 9 13 15 16 13 1 9 10 9 15
2 3 13
6 3 13 9 10 9 15
24 3 13 15 10 9 1 9 0 3 7 13 15 15 10 9 10 9 7 10 9 15 7 13 15
8 0 15 15 13 16 13 13 15
2 13 11
2 13 3
9 9 10 9 15 13 7 15 0 13
12 3 13 15 10 9 7 6 9 13 7 13 15
24 7 13 10 11 13 13 1 11 10 0 1 9 11 7 11 16 13 10 13 1 11 10 9 13
33 9 11 7 9 11 9 9 1 10 11 11 10 9 10 9 10 13 1 9 9 13 0 7 10 13 1 9 7 9 9 9 13 15
8 1 3 13 10 11 13 7 13
6 13 3 10 9 10 9
24 13 3 1 10 9 10 11 13 12 9 11 10 13 11 7 11 10 9 15 13 9 1 10 9
3 13 3 9
3 7 13 15
8 6 1 15 7 13 15 9 9
28 7 13 3 13 0 12 9 11 10 10 11 7 11 10 9 15 1 10 9 1 11 10 9 15 13 10 9 15
3 7 13 15
27 7 13 1 0 10 11 13 1 10 9 15 7 13 10 9 10 9 7 13 15 9 7 15 9 1 10 9
9 7 13 10 9 15 1 0 10 11
21 7 13 15 15 10 3 13 0 9 7 9 13 7 13 7 13 7 0 7 13 15
18 7 13 15 9 0 1 10 11 7 11 7 11 7 11 7 1 10 11
8 13 3 10 9 13 1 10 9
8 7 13 15 13 15 10 9 15
12 0 10 0 10 9 16 15 13 10 9 10 9
6 0 10 13 16 15 13
10 0 10 13 7 13 10 9 16 15 13
6 0 10 0 16 15 13
10 0 10 0 10 9 16 15 10 9 13
7 0 10 0 16 9 9 13
12 0 10 13 1 9 16 15 13 10 9 10 9
16 0 13 3 13 15 7 13 7 13 15 0 1 15 13 1 15
6 15 13 10 9 10 9
8 16 3 10 9 13 1 15 13
12 1 15 13 3 3 3 13 3 13 1 10 9
6 15 13 10 9 10 9
7 3 13 9 13 1 9 13
20 7 13 9 7 13 15 1 10 9 7 1 10 9 7 13 15 10 1 10 9
23 3 13 10 9 15 1 10 9 16 13 15 10 0 9 7 13 10 9 15 10 1 10 9
10 3 13 16 13 13 10 9 7 10 9
4 6 3 13 15
23 16 3 13 10 9 7 10 9 9 12 7 12 9 3 3 13 1 10 9 16 3 15 13
22 15 16 3 13 12 10 9 0 10 0 7 13 3 10 9 0 13 1 10 9 10 9
14 15 3 3 13 7 13 0 0 13 1 10 9 10 9
23 13 3 15 16 16 3 13 15 10 9 0 10 9 7 9 3 3 13 1 10 9 10 9
5 13 16 13 10 0
2 3 13
8 15 3 3 13 0 13 10 9
12 15 3 3 13 0 0 13 1 10 11 10 9
42 16 3 13 10 9 15 1 10 9 7 3 13 16 10 9 15 13 15 1 15 13 3 10 9 15 1 10 9 7 13 0 13 10 9 15 7 3 13 13 10 9 15
30 13 13 10 9 15 0 16 15 13 1 15 1 10 9 16 15 13 10 9 10 9 7 10 9 10 9 7 1 9 13
3 6 13 15
10 3 3 13 3 16 3 13 10 0 9
3 13 16 13
2 3 13
15 16 3 10 9 15 10 0 13 15 13 15 7 13 1 15
14 7 16 10 0 15 9 13 15 13 15 7 13 1 15
18 13 3 15 16 13 12 10 9 15 7 3 0 10 9 15 1 11 13
2 13 3
9 15 3 13 10 9 15 13 15 9
23 15 3 13 15 16 15 10 13 10 9 15 1 9 9 13 15 13 7 15 3 13 13 13
6 3 13 16 13 10 0
7 13 3 10 9 10 9 15
7 15 3 13 15 3 13 3
10 7 1 10 9 16 9 13 10 9 15
9 7 1 11 16 9 13 10 0 9
15 7 1 10 9 15 13 16 3 13 12 9 0 13 7 0
9 13 3 10 9 15 6 6 3 3
8 10 3 0 0 1 10 0 13
7 9 1 9 7 9 1 9
8 15 3 13 15 3 13 10 0
13 7 15 15 13 1 10 0 9 13 15 3 10 0
10 7 15 15 13 9 12 13 1 15 12
12 10 13 15 13 7 10 13 1 15 13 3 13
3 13 16 13
9 13 10 3 15 7 13 10 0 15
34 13 10 0 15 7 13 1 10 13 15 16 13 9 10 9 15 10 1 9 16 10 9 15 13 1 0 7 0 7 13 1 0 7 0
9 16 3 13 10 13 15 15 9 13
7 3 3 10 9 10 15 13
10 7 16 13 10 9 15 0 15 0 13
12 13 3 15 0 3 10 9 15 10 0 0 13
14 13 3 10 9 15 3 13 1 10 9 1 10 13 15
13 16 3 3 9 3 13 1 10 9 15 10 1 9
3 6 13 15
4 13 10 9 15
33 15 3 13 9 3 13 10 0 15 15 13 10 0 15 16 10 15 9 13 1 10 0 7 10 9 15 10 13 1 10 0 13 15
8 7 3 13 3 13 3 10 9
17 3 13 1 10 9 7 1 10 9 10 9 13 13 16 13 10 9
4 13 10 9 15
22 15 3 3 13 13 1 10 9 15 7 13 10 9 15 13 10 9 15 10 1 10 0
7 13 3 3 13 3 10 0
8 13 3 16 1 10 9 15 13
4 3 3 13 15
13 13 3 10 9 15 15 9 13 1 10 15 13 15
4 3 3 13 15
10 9 15 10 1 10 9 13 10 9 15
10 13 10 9 15 3 1 9 3 1 9
13 7 13 15 10 9 15 3 7 15 13 10 9 15
12 7 3 13 15 1 9 7 13 15 1 10 0
16 16 3 13 10 9 10 9 15 13 7 15 10 9 15 10 0
14 16 3 3 13 10 9 3 10 9 15 13 10 9 15
9 3 3 13 3 13 3 10 9 0
10 13 3 10 9 15 16 13 10 9 13
3 6 13 15
11 7 10 9 15 10 13 1 10 0 13 15
18 3 13 15 9 1 10 9 3 9 7 9 13 7 3 9 13 7 13
19 13 3 15 9 1 9 3 7 9 7 9 13 7 3 9 3 13 7 13
12 3 3 13 10 9 15 3 13 3 10 9 15
7 10 9 10 9 13 10 9
12 16 13 10 9 15 0 0 10 9 15 0 13
13 16 3 10 9 15 0 13 0 10 9 15 0 13
12 16 3 10 9 10 1 15 9 13 10 9 15
16 7 3 10 12 13 7 10 0 13 7 12 13 7 10 0 13
6 3 13 9 13 7 9
4 1 0 13 15
13 3 13 10 9 15 15 13 7 10 9 15 15 13
12 3 10 9 0 13 10 9 7 10 9 10 9
23 13 1 10 9 10 9 16 3 13 7 13 7 13 1 9 7 10 9 15 10 0 13 15
5 3 15 3 13 15
13 15 3 1 15 13 13 13 1 10 9 15 9 12
2 3 13
2 7 13
15 13 3 15 16 3 11 1 15 10 9 15 13 3 12 0
22 16 3 10 9 10 9 3 13 7 3 1 9 13 10 9 3 13 3 0 3 15 0
12 3 3 13 13 15 13 7 15 13 7 15 13
6 15 3 0 10 9 13
11 13 3 10 9 15 10 0 16 13 0 0
6 3 3 13 1 10 3
6 0 10 9 10 9 15
5 3 13 16 3 13
13 1 15 3 9 13 13 7 1 15 9 13 13 15
12 15 3 13 10 9 10 1 10 9 10 9 15
9 10 3 1 10 15 9 9 3 13
6 7 3 13 10 9 15
7 13 10 9 1 10 9 15
8 7 6 10 9 1 10 9 15
25 3 13 10 0 10 9 7 13 10 9 15 1 10 9 16 13 15 1 10 9 15 7 13 13 15
4 13 7 13 15
3 13 7 13
4 13 7 13 15
13 15 3 10 13 13 7 10 13 13 7 10 13 13
4 7 7 9 13
4 3 9 13 15
26 16 3 15 0 13 13 9 0 13 10 9 15 15 3 10 9 15 10 1 10 9 13 0 10 13 15
8 0 3 13 10 9 7 10 9
5 13 1 10 0 9
18 3 0 7 0 10 9 10 13 1 10 9 7 0 13 10 13 1 15
17 3 0 7 13 10 9 10 13 1 10 9 7 0 13 10 13 15
5 3 3 13 9 0
6 1 10 9 15 13 15
9 3 13 1 9 9 7 1 9 9
7 3 15 9 0 9 0 13
13 3 13 9 0 9 0 13 7 9 0 9 0 13
11 15 9 3 13 9 0 13 7 1 9 13
7 3 1 10 9 15 13 15
7 0 13 15 1 0 10 9
20 9 9 3 10 15 9 13 7 10 15 9 9 13 7 10 15 9 9 0 13
5 7 3 13 15 16
3 3 13 15
7 13 1 15 10 13 10 9
20 7 13 10 9 7 13 10 9 7 13 10 9 7 13 10 9 0 7 3 13
5 13 3 1 10 9
25 7 13 10 9 7 13 10 9 7 13 10 9 7 13 10 9 0 7 13 7 13 10 9 15 0
16 7 13 16 13 10 11 10 9 0 13 10 9 1 10 9 15
13 13 3 13 15 3 9 13 7 3 3 10 9 15
10 13 3 15 1 10 9 13 15 9 0
7 7 6 0 13 13 15 13
6 9 16 13 13 15 13
1 13
6 7 3 13 15 10 9
5 7 13 15 10 11
19 13 15 13 7 13 15 13 10 9 7 13 10 9 15 13 11 1 9 15
12 13 3 15 1 11 13 15 9 13 15 7 13
11 9 10 9 15 13 1 10 9 0 3 13
2 13 15
4 15 13 13 15
9 7 0 13 9 7 13 10 9 15
11 3 3 15 9 13 1 9 13 1 15 9
6 7 13 0 13 7 13
5 7 0 13 7 13
8 7 10 9 15 13 0 7 13
9 13 3 10 11 13 7 13 10 13
3 6 13 15
7 3 1 10 11 0 9 13
11 10 3 9 10 9 13 1 10 9 10 0
9 3 13 10 9 7 10 9 10 9
6 7 13 10 11 10 9
1 13
4 3 13 13 15
8 7 13 10 9 1 10 9 0
15 7 13 10 11 1 10 9 11 13 10 9 15 13 7 13
10 7 13 10 9 15 7 13 15 10 9
20 7 13 10 9 9 7 15 10 3 13 13 16 13 10 13 1 11 10 9 13
9 0 10 9 15 13 7 10 9 13
13 13 3 10 11 0 9 1 15 13 13 1 10 3
6 7 13 12 9 13 15
6 9 13 15 3 3 13
5 7 13 15 10 11
10 10 9 9 13 7 10 9 10 9 9
6 0 3 10 9 13 15
4 15 3 13 15
10 13 15 7 13 10 0 13 10 15 0
11 7 13 15 1 10 9 13 15 10 9 15
15 7 6 9 0 13 1 10 9 16 10 9 13 1 10 9
3 15 3 13
5 7 13 13 15 13
1 13
3 7 13 15
12 3 13 13 10 9 7 10 9 7 13 9 0
5 10 3 9 13 13
12 15 13 0 16 3 10 9 7 10 9 15 13
30 7 13 15 1 10 3 1 10 9 10 0 13 15 12 13 1 10 9 13 0 3 16 3 13 15 13 1 10 9 0
4 7 6 13 13
6 13 3 1 9 13 15
9 13 3 3 1 15 9 9 0 13
6 10 3 9 13 15 13
3 7 13 15
1 13
7 15 3 13 13 1 10 9
17 7 6 13 15 10 9 1 10 9 1 10 9 7 13 1 10 9
20 7 6 15 10 9 13 1 9 10 11 7 13 15 13 16 13 1 10 9 15
11 7 13 1 9 13 7 13 1 10 0 9
8 7 6 13 15 0 1 9 13
10 7 13 10 11 10 9 15 13 10 0
4 13 15 10 9
8 7 6 15 10 9 13 1 15
2 0 13
7 3 13 0 1 10 9 15
11 15 3 13 0 13 13 15 10 9 7 13
3 13 7 13
15 16 3 13 16 9 13 10 9 10 9 1 10 9 13 9
4 3 13 10 0
7 7 13 13 1 10 9 15
15 13 3 10 9 13 7 13 10 9 10 13 9 0 10 9
2 13 15
4 7 13 13 15
7 7 13 15 13 1 10 9
13 6 0 9 7 0 13 13 10 11 7 10 9 15
8 7 13 10 9 13 10 9 15
11 1 15 1 10 9 7 0 13 10 9 15
10 3 9 13 10 13 9 7 10 3 13
5 9 13 7 3 9
7 3 3 13 13 0 7 0
7 3 13 15 10 9 11 13
13 1 15 15 7 10 9 13 10 3 9 15 3 13
5 7 13 15 10 11
14 3 13 10 9 10 9 13 1 15 1 15 13 10 9
12 13 3 9 3 13 1 15 10 9 7 3 13
7 7 13 9 0 1 9 0
14 16 3 3 13 10 9 7 10 9 13 7 10 9 13
10 7 13 9 0 1 9 0 7 0 13
10 0 15 13 15 6 9 13 13 15 13
15 10 9 15 3 13 7 13 13 10 9 15 1 15 7 13
10 7 13 10 11 13 15 7 10 9 15
14 7 6 9 13 12 9 13 3 13 10 9 10 9 15
4 13 3 1 15
7 15 3 13 7 13 15 13
1 13
6 9 10 9 15 13 15
8 7 13 10 9 1 10 9 0
18 7 13 10 11 1 10 9 10 9 7 13 10 9 7 10 9 13 13
1 13
7 3 3 13 10 9 7 13
3 7 13 15
12 7 13 3 10 11 13 15 12 0 13 7 13
4 13 15 9 11
14 13 3 1 10 9 13 15 10 0 7 13 15 10 11
5 13 16 13 0 13
2 13 15
2 6 9
6 3 13 10 9 15 13
5 7 13 15 10 9
3 13 15 13
10 15 3 13 13 15 1 0 10 9 0
9 15 3 13 6 13 15 9 0 13
7 7 13 10 9 13 10 0
5 7 13 10 9 13
6 3 13 3 1 10 11
8 1 10 9 10 9 13 10 9
28 7 13 10 11 10 9 15 7 10 9 13 1 10 9 15 7 13 10 9 10 9 7 13 15 9 7 15 9
5 3 13 10 9 15
4 10 3 9 0
4 10 3 9 0
13 13 3 10 9 10 9 16 13 9 1 10 9 15
21 7 13 10 12 9 15 13 15 9 9 0 16 13 15 7 13 15 9 7 15 9
45 0 11 10 13 11 7 11 10 9 15 7 11 10 10 11 7 11 10 9 15 11 7 11 11 7 11 10 9 11 10 10 11 7 11 11 10 0 7 11 10 11 10 3 13 15
9 0 10 12 13 10 11 13 15 13
11 1 9 9 3 13 7 1 9 9 3 13
10 13 3 13 13 16 13 10 9 10 9
2 13 13
2 0 13
2 0 13
2 3 13
2 3 13
22 3 13 9 7 9 7 9 1 10 9 15 3 9 1 9 7 12 9 7 9 7 9
7 0 3 10 9 10 9 15
6 7 3 13 16 3 13
7 13 3 1 10 9 13 15
13 7 16 3 13 10 9 0 13 10 9 15 1 15
26 7 15 3 3 13 15 7 13 10 9 15 13 1 10 9 7 10 9 0 13 10 9 1 10 9 15
3 6 13 15
13 0 13 9 11 7 11 1 9 9 3 10 9 0
9 6 15 13 15 3 9 1 0 9
11 13 3 0 3 10 9 7 0 3 10 9
12 13 3 15 1 9 7 1 10 9 15 13 15
15 7 1 9 3 7 9 13 1 15 1 9 15 7 10 9
9 13 3 15 1 0 10 9 15 13
16 3 3 15 13 10 13 7 10 9 10 9 15 10 13 1 15
17 13 3 9 9 1 9 7 9 9 7 13 9 1 9 7 13 15
9 7 13 13 1 15 1 10 9 15
7 10 3 13 1 9 0 13
12 3 3 13 15 1 10 9 0 13 1 10 0
13 3 3 13 10 9 10 11 16 13 10 9 10 9
16 0 10 9 16 13 3 10 9 15 7 10 9 3 10 9 15
10 16 10 9 11 13 15 3 10 9 15
4 3 3 13 15
12 15 3 13 13 15 3 13 7 0 15 3 13
10 15 13 15 1 10 9 13 1 10 9
10 7 15 1 10 9 13 13 1 10 9
14 7 3 13 1 10 13 10 9 10 3 9 3 13 13
13 7 12 1 15 3 13 1 10 9 1 10 9 15
10 15 3 3 10 9 10 9 15 13 13
3 3 3 13
4 0 9 13 15
21 15 3 15 13 1 15 1 10 9 13 7 15 1 15 1 10 9 15 10 1 9
19 15 3 3 13 15 1 10 9 13 7 15 15 1 10 9 15 10 1 9
9 3 13 16 13 13 9 1 10 9
6 3 13 13 9 7 9
7 7 0 10 9 10 9 15
38 10 13 9 7 9 1 15 3 13 15 0 7 10 13 9 7 9 1 15 3 13 15 0 7 15 3 13 10 9 15 7 13 1 15 3 13 15 0
17 10 13 10 9 15 13 15 7 10 13 10 9 15 1 15 13 15
13 10 13 15 15 13 7 10 15 13 13 10 13 15
19 10 13 9 1 9 9 9 9 13 7 10 13 0 1 9 0 9 0 13
23 7 15 3 13 12 10 0 0 9 0 0 1 9 9 6 13 15 3 3 13 10 9 15
11 7 13 16 13 10 11 13 10 12 9 15
10 13 3 10 13 7 13 1 10 9 15
3 7 0 13
6 7 13 10 11 13 15
7 13 13 11 15 13 7 13
16 0 13 7 0 13 0 13 7 0 13 7 0 13 7 0 13
9 7 0 13 15 3 3 13 1 15
11 0 3 13 13 10 11 13 10 9 1 11
6 15 13 1 10 0 13
4 7 15 13 13
10 6 10 10 0 13 1 10 9 10 9
3 7 15 13
2 9 13
3 6 13 15
3 7 0 9
5 0 13 1 15 13
3 6 13 15
9 3 13 1 0 9 0 11 10 9
18 1 3 10 9 11 10 9 1 3 10 9 10 9 13 7 9 13 15
20 15 3 10 9 7 10 9 1 11 13 7 16 13 13 0 13 11 10 13 13
4 10 13 9 13
6 15 3 13 10 9 0
12 0 13 9 13 1 10 9 15 13 10 0 13
4 13 7 3 13
9 13 3 11 7 13 7 13 7 13
2 9 13
9 6 9 9 7 9 9 9 7 0
8 7 13 10 9 1 10 9 15
15 3 13 13 10 9 1 15 13 10 0 9 15 16 3 13
3 6 15 11
20 3 16 1 11 7 11 13 10 9 10 13 1 15 3 3 1 9 7 9 13
3 3 13 15
10 11 7 11 0 13 1 9 9 3 15
7 7 15 11 3 1 9 13
13 3 13 15 16 9 11 0 13 1 9 9 3 15
8 1 0 10 9 13 10 11 13
20 13 15 9 9 10 9 7 10 9 16 13 0 1 0 7 0 7 13 15 0
32 15 15 13 1 10 9 15 7 15 13 10 9 3 3 10 9 7 10 9 15 13 3 3 10 9 7 15 3 13 10 9 13
12 6 1 15 15 10 13 7 13 7 15 13 15
23 13 10 9 15 1 15 7 13 1 15 16 0 13 7 0 10 9 7 13 9 10 9 15
11 10 3 9 15 0 7 10 9 15 0 13
12 1 0 10 9 13 10 11 10 9 1 10 0
6 10 3 9 13 13 15
11 6 10 9 15 13 15 3 13 13 1 9
11 3 13 15 13 11 16 13 7 10 1 15
28 3 13 1 10 9 10 9 7 10 9 10 9 13 15 3 13 13 15 13 7 10 1 15 3 3 10 9 0
20 7 3 13 1 10 9 16 10 9 10 9 1 10 9 10 9 13 7 0 13
9 13 3 15 16 10 9 0 13 3
15 16 3 13 15 13 9 13 7 3 9 3 3 13 10 0
9 9 3 13 10 9 10 9 10 9
6 7 6 9 9 13 0
4 15 3 13 15
22 15 13 1 15 9 15 13 9 12 7 16 13 0 10 9 1 9 3 13 15 7 13
5 15 3 13 9 9
6 3 13 10 9 3 13
4 3 13 10 9
4 13 15 10 9
8 7 13 7 13 0 3 10 0
16 7 13 15 0 7 13 15 15 7 13 15 16 3 0 15 13
9 16 13 10 13 1 11 10 9 13
15 6 10 9 15 15 13 10 0 15 1 15 13 10 9 15
11 13 10 9 15 1 15 7 9 10 9 13
13 3 13 7 13 7 13 15 1 10 9 10 9 15
16 9 13 3 13 7 9 13 3 13 16 3 13 1 9 10 9
6 7 10 9 15 9 13
7 3 13 15 13 0 7 0
7 7 13 15 10 9 7 13
6 3 0 13 10 9 11
5 10 3 9 13 13
13 0 3 13 10 9 3 3 1 10 11 9 10 9
7 13 3 10 9 15 13 15
16 15 9 13 1 15 13 7 15 9 7 9 13 1 15 3 13
10 7 16 10 11 10 11 13 1 15 13
6 3 3 13 10 9 15
17 16 3 1 9 9 15 13 10 9 3 13 1 15 10 9 10 9
27 7 3 13 15 13 1 10 9 10 0 7 10 9 15 13 16 3 0 13 10 0 7 3 10 9 15 13
15 10 3 13 1 15 1 15 13 7 10 3 13 1 15 13
4 1 0 13 15
7 15 9 7 9 13 10 9
7 10 3 10 9 9 3 13
12 7 15 3 13 9 1 10 9 10 9 13 15
20 7 13 10 9 0 7 10 9 15 0 7 13 10 9 0 7 10 9 15 0
8 9 9 3 13 0 13 0 13
9 1 3 10 9 10 9 10 9 13
20 10 0 9 1 10 0 9 13 10 0 7 10 0 9 1 10 0 9 13 0
18 13 3 15 16 15 9 0 15 13 10 9 13 1 15 9 1 9 9
12 1 3 10 9 15 13 7 1 10 9 15 13
9 3 13 15 15 10 9 7 9 13
5 15 3 13 13 15
18 9 0 7 9 9 13 7 9 3 13 15 3 3 10 9 11 10 9
19 9 9 13 1 10 9 1 10 9 0 7 13 15 16 13 1 10 9 11
5 7 6 0 11 3
24 9 9 13 1 10 9 1 10 9 0 7 13 15 16 13 1 10 9 10 9 13 10 9 11
5 7 6 0 11 3
18 3 3 10 0 9 13 1 10 9 13 1 0 9 13 9 7 3 13
7 1 10 9 15 13 3 13
8 7 13 13 13 7 13 7 13
25 3 13 7 13 1 15 12 0 9 0 15 7 13 13 3 7 13 10 0 10 9 0 0 10 0
17 3 15 13 10 9 6 10 9 7 10 9 15 13 3 13 15 13
4 13 3 15 15
13 6 10 9 15 7 10 9 15 3 13 13 15 13
7 15 3 13 13 10 13 15
9 7 13 10 9 1 10 9 15 13
8 6 10 9 15 7 10 9 15
20 15 3 3 13 10 9 10 9 15 10 1 9 15 15 9 7 9 7 9 13
14 1 10 9 0 13 10 11 1 10 9 13 1 10 9
7 7 13 15 0 1 9 13
6 6 13 10 13 10 13
18 7 1 10 13 15 15 3 13 1 10 9 7 13 10 9 7 13 15
11 9 3 13 13 7 1 10 3 13 9 13
13 0 3 13 1 10 9 7 13 10 9 7 13 15
20 0 3 13 1 10 9 10 0 7 13 9 15 3 12 15 3 12 15 3 12
4 10 13 9 13
6 7 13 10 9 13 15
4 15 3 13 13
10 3 15 13 13 10 9 10 9 10 9
7 15 3 13 13 15 7 13
10 15 3 3 13 3 15 13 13 1 15
16 1 0 1 9 15 13 16 13 3 13 7 13 3 13 7 13
8 7 13 15 10 9 11 10 13
13 9 13 7 3 3 13 7 13 13 7 3 3 13
34 13 3 10 9 10 9 0 7 10 9 3 13 7 10 9 15 13 16 13 10 9 7 10 9 13 7 10 9 13 7 13 7 13 15
22 6 13 15 16 0 9 7 0 13 13 15 13 7 3 13 7 13 15 13 7 3 13
20 15 13 10 9 10 9 7 3 13 13 10 0 7 13 10 13 1 10 9 15
7 0 13 10 1 10 9 13
18 10 3 1 10 0 13 0 13 10 10 9 13 7 3 1 9 13 15
19 3 13 3 9 1 15 7 0 13 13 3 9 7 9 1 10 9 3 13
28 10 3 1 10 9 13 0 13 10 10 9 13 7 10 9 10 9 7 10 9 10 9 13 10 9 7 0 13
29 10 3 1 10 0 9 13 0 13 10 10 9 13 7 13 15 3 13 7 13 15 3 12 15 3 12 15 3 12
5 0 9 13 15 13
13 16 3 13 10 9 7 9 13 3 13 3 10 9
8 13 3 10 9 10 9 13 15
9 9 3 0 9 13 1 10 15 9
4 3 3 13 9
4 15 3 13 15
4 0 9 0 13
5 10 3 9 13 15
5 13 3 13 13 15
10 3 3 13 10 9 13 1 15 10 9
14 13 13 0 1 10 9 7 1 9 10 9 13 10 9
13 13 0 10 9 7 13 15 1 9 1 10 13 15
8 10 3 9 13 1 10 9 15
5 0 9 13 15 13
16 0 13 10 9 10 9 9 9 15 13 9 13 1 10 9 15
7 15 0 3 13 15 10 9
22 3 3 13 0 10 9 13 7 13 9 16 13 10 9 10 9 7 13 1 10 9 15
24 0 15 13 10 11 1 9 10 9 7 1 9 15 13 15 16 13 10 13 1 10 9 11 13
6 13 1 9 10 9 15
4 13 13 1 9
8 3 13 10 9 13 1 10 9
7 7 13 15 10 9 15 13
8 13 15 10 9 10 9 10 9
4 15 3 13 13
6 10 3 9 13 10 9
8 10 3 9 13 10 9 10 0
9 10 3 0 10 13 15 13 10 9
6 10 3 9 9 9 13
5 10 3 9 9 13
15 3 3 13 10 9 7 9 13 3 13 1 10 9 10 9
30 13 10 9 10 9 10 9 15 7 13 1 10 9 15 15 10 9 7 10 13 10 9 7 13 15 1 10 9 10 9
13 3 10 0 13 3 10 9 1 10 9 10 9 15
4 10 13 9 13
16 7 1 10 9 15 13 7 13 15 15 13 7 13 10 9 0
12 3 0 13 10 9 10 9 9 9 13 0 9
13 13 3 12 0 9 13 13 15 15 13 7 13 15
17 3 0 13 10 9 10 9 9 13 1 10 9 7 1 15 9 13
14 15 16 13 13 1 10 9 7 13 13 10 0 1 9
7 3 13 1 10 9 10 9
19 13 10 9 7 13 10 0 1 0 10 0 7 13 15 1 10 9 10 9
9 3 13 10 9 7 10 9 10 9
2 13 15
1 6
4 15 3 13 15
22 1 0 15 9 13 10 9 10 9 0 13 9 9 15 13 1 10 9 15 0 7 0
17 7 13 1 10 9 15 13 15 1 10 9 15 16 13 15 7 13
8 3 0 10 9 0 7 10 9
7 3 0 13 10 10 9 9
17 3 10 9 15 13 11 7 10 9 15 11 7 11 7 11 7 11
5 3 3 0 0 15
4 7 13 1 15
5 10 3 11 13 15
10 7 3 13 3 9 0 1 10 9 15
16 1 0 10 9 13 11 10 9 10 9 11 7 13 10 9 15
5 0 13 11 10 9
13 15 13 1 10 0 7 1 0 10 9 13 1 15
18 10 3 11 13 10 11 13 7 1 9 13 1 11 10 9 10 9 15
5 3 13 15 13 15
12 7 13 15 13 13 10 9 16 3 9 15 13
18 15 3 13 1 10 9 15 13 15 13 3 1 9 10 9 11 10 9
19 7 13 10 9 1 10 9 7 10 13 13 13 7 13 13 11 1 10 9
16 7 13 10 9 15 1 9 7 13 10 9 7 13 10 9 15
16 7 13 10 9 15 13 10 9 7 13 15 7 13 13 10 11
13 13 3 10 11 13 3 1 9 1 0 9 1 0
10 7 13 10 9 13 15 0 1 10 9
8 0 3 13 13 15 10 9 13
12 13 3 10 9 16 13 1 10 9 13 15 9
4 15 3 13 15
4 3 9 13 13
4 13 15 15 13
4 15 3 13 15
10 3 13 3 3 3 12 9 7 12 9
3 15 3 13
14 7 13 15 7 13 7 13 10 13 10 9 12 9 0
11 10 3 13 13 9 3 12 1 9 7 9
19 7 13 10 9 13 1 10 9 7 13 15 1 10 3 16 15 13 10 9
11 7 13 10 9 13 1 10 9 1 0 13
6 0 3 13 0 13 3
12 10 3 9 3 0 10 9 13 13 1 10 9
5 13 3 0 10 9
12 0 3 9 10 9 13 1 15 13 1 10 9
5 3 3 13 15 13
1 13
2 15 13
2 3 13
6 13 3 15 10 11 13
12 9 16 15 13 13 15 13 1 15 1 10 9
3 15 3 13
1 13
3 9 13 15
12 3 3 10 11 13 10 9 13 15 7 13 15
4 0 1 15 13
9 7 13 15 1 10 9 13 10 9
8 10 3 1 10 9 13 15 13
4 3 9 9 13
8 7 13 13 1 10 9 1 11
4 7 15 13 13
10 1 15 10 9 15 13 10 9 10 0
8 3 3 13 10 9 3 9 13
5 15 3 13 13 15
13 1 15 3 15 13 10 9 10 9 1 10 9 15
5 10 3 9 13 13
14 13 10 9 7 10 9 7 10 13 9 7 9 9 13
24 15 3 13 10 9 7 10 9 9 15 3 1 15 13 3 3 13 10 9 15 7 10 9 15
10 7 13 10 9 10 9 1 10 9 15
7 10 9 0 10 9 15 13
8 10 3 9 15 3 13 1 15
8 3 3 13 15 13 9 9 9
6 7 13 10 9 13 15
3 13 7 13
6 3 13 10 9 13 15
8 13 16 10 9 13 10 9 13
4 15 3 13 13
2 13 15
4 9 13 0 0
9 0 3 0 16 13 0 1 9 13
6 13 3 10 11 13 15
3 15 3 13
5 3 3 15 0 13
17 3 13 16 15 10 13 1 10 9 1 10 9 13 7 1 9 13
15 10 3 13 1 10 9 1 10 9 13 7 0 13 10 9
6 0 13 10 13 10 9
9 10 3 0 9 13 3 13 10 9
12 7 13 3 10 11 13 1 10 9 11 7 11
5 13 15 9 9 11
5 10 9 15 3 13
6 15 3 3 13 15 9
8 7 13 10 9 15 13 15 13
6 13 15 16 13 1 15
11 3 13 3 3 1 10 9 10 13 9 11
6 15 3 13 13 15 13
4 15 3 13 13
11 3 13 13 10 9 10 9 7 13 10 9
3 15 3 13
2 6 9
16 3 3 10 9 13 1 10 9 10 13 1 10 9 10 9 15
6 3 13 10 11 13 15
4 13 15 3 13
18 7 13 3 10 11 13 1 10 9 10 11 7 13 1 10 9 13 3
22 7 13 15 9 0 13 1 15 0 0 0 0 7 0 0 7 13 15 1 10 9 15
18 7 13 15 16 10 9 13 13 0 13 0 0 7 0 13 7 0 13
5 7 13 10 9 11
8 10 3 11 13 10 9 15 13
15 13 1 10 9 16 3 9 12 13 15 7 3 13 15 13
11 7 13 15 0 3 13 16 13 1 10 9
5 7 13 15 10 11
3 15 9 13
3 15 3 13
4 12 7 0 9
27 7 13 10 9 13 1 10 9 13 10 12 9 7 10 9 7 13 13 7 13 10 9 10 3 9 10 9
14 7 13 15 7 13 7 10 13 10 9 13 12 9 0
10 10 3 13 13 12 9 1 9 7 9
14 7 13 10 9 13 1 10 9 7 13 1 10 9 11
5 15 3 13 13 15
3 0 13 13
1 9
4 13 3 10 9
2 7 3
2 3 9
5 13 3 13 10 9
14 10 3 9 10 9 13 13 10 3 9 10 9 3 13
10 7 13 10 9 1 10 3 13 9 13
5 10 3 11 13 15
10 13 7 13 1 10 9 10 9 7 9
7 15 3 13 1 15 13 16
3 9 3 13
5 13 3 10 11 13
9 15 13 1 15 0 16 9 3 13
11 7 13 10 12 9 10 12 7 15 9 13
9 3 3 13 16 3 1 9 13 15
9 13 3 1 10 9 10 9 7 9
21 3 13 16 3 13 13 1 10 9 10 9 7 9 7 1 10 9 10 9 7 9
15 13 3 10 11 1 10 9 11 10 11 13 10 9 15 13
9 15 13 10 9 13 10 9 10 9
3 15 3 13
3 0 3 11
7 0 3 11 7 12 10 9
6 15 3 15 15 13 13
5 13 3 11 11 13
10 15 13 10 11 10 9 10 9 10 13
6 13 3 10 11 13 15
19 0 13 11 11 16 9 7 9 3 13 15 7 10 9 15 10 1 10 9
32 13 15 10 9 10 9 10 9 7 15 3 13 1 10 9 13 13 1 10 9 7 15 3 13 1 10 9 13 13 1 10 9
12 3 13 10 9 16 15 13 16 15 13 10 11
32 1 3 13 10 11 13 10 9 15 16 13 15 1 11 13 7 0 13 1 10 0 7 9 7 9 7 13 7 10 0 9 13
3 0 15 9
5 3 3 13 15 0
6 15 3 13 13 10 11
4 13 1 15 11
7 3 10 11 13 10 9 15
16 16 15 13 1 15 13 13 15 7 13 10 9 15 7 13 15
10 15 3 3 13 10 9 15 13 13 15
11 15 3 3 13 10 9 15 1 15 13 15
8 7 15 13 9 9 10 9 15
25 13 3 10 9 10 9 13 1 10 9 10 9 15 1 10 9 15 7 3 13 15 1 10 9 15
26 6 13 15 16 13 15 10 3 13 15 3 3 13 9 16 3 13 10 9 10 9 13 1 10 9 15
12 7 13 1 15 7 13 10 9 15 3 10 9
9 10 3 9 15 13 0 3 10 9
10 7 6 13 15 11 7 11 13 1 15
7 13 3 10 11 13 10 11
6 9 0 13 15 3 13
15 3 15 13 6 9 0 13 15 7 6 9 1 10 9 13
10 0 13 10 9 15 10 0 1 15 13
11 7 13 10 9 13 1 9 15 7 13 3
8 7 13 10 11 7 13 15 13
4 13 7 3 13
12 13 3 10 9 15 15 13 3 3 10 11 0
11 7 13 15 1 10 9 13 15 10 11 13
13 15 13 10 9 16 15 10 9 10 9 1 0 13
10 15 3 10 9 13 16 11 13 13 0
6 11 3 13 7 13 15
17 13 3 15 16 11 3 13 7 3 13 15 7 13 1 15 15 13
10 3 3 10 9 10 9 13 13 1 15
11 3 13 10 9 16 1 11 10 9 13 15
12 7 13 1 10 9 13 15 9 13 15 7 13
10 9 13 15 10 9 16 13 7 3 13
11 3 3 13 1 10 9 7 3 1 10 9
10 6 9 0 7 13 1 3 1 15 13
4 1 3 13 15
4 13 15 15 3
19 7 13 15 10 11 7 13 1 15 10 9 7 13 10 9 1 10 9 0
9 3 13 10 9 10 11 1 0 13
7 1 15 15 3 13 13 15
4 15 3 13 15
4 1 10 9 15
10 16 13 9 3 9 9 13 10 9 0
3 13 3 3
6 7 13 7 15 13 15
10 13 3 15 1 10 11 13 15 10 11
17 13 10 9 10 9 13 1 9 9 7 13 15 7 10 0 9 13
3 7 13 3
14 13 3 15 1 11 13 10 10 9 13 10 11 7 13
6 10 9 15 3 13 9
10 7 13 1 10 9 13 15 10 11 13
4 15 15 13 11
10 10 9 10 9 1 15 13 9 7 9
8 1 10 9 15 7 1 10 0
9 13 3 1 10 0 13 15 10 11
5 3 0 13 10 9
23 16 3 3 13 15 13 1 9 13 9 7 10 13 0 9 13 7 13 10 9 15 13 9
10 1 0 10 9 13 10 9 10 11 13
10 7 13 9 13 15 1 0 15 7 13
3 6 13 15
16 16 3 13 7 13 3 10 9 3 3 13 1 10 9 10 9
17 15 3 13 15 3 10 9 0 0 13 10 0 1 10 9 10 9
13 7 15 3 13 12 9 0 1 10 9 15 15 13
29 15 3 3 13 12 10 0 0 10 13 1 15 13 15 16 13 9 0 1 10 9 15 7 13 1 10 9 10 9
6 9 3 13 13 10 9
9 3 6 10 9 1 15 10 9 13
23 0 15 13 13 1 10 9 0 7 0 3 12 9 7 12 9 13 13 1 10 9 10 0
13 7 16 10 9 15 13 15 13 15 7 13 1 15
18 0 15 13 0 1 10 9 13 3 12 9 13 13 1 10 11 10 9
7 13 3 13 12 10 0 0
20 13 3 15 16 10 9 15 1 9 1 15 13 10 9 10 9 15 10 1 9
22 16 13 15 9 12 9 7 13 12 1 15 3 13 10 12 1 10 9 13 13 10 13
20 7 16 13 13 15 6 13 15 16 13 1 15 3 3 1 10 12 10 3 13
17 3 3 13 9 1 10 9 15 10 1 9 16 13 12 10 0 0
7 16 15 13 13 10 9 15
21 16 3 3 13 13 1 15 3 12 7 12 16 1 9 12 9 7 12 13 15 9
7 16 3 13 15 13 10 9
14 16 3 3 10 9 13 13 15 3 10 0 7 10 9
21 15 3 13 1 10 9 13 13 1 9 7 15 3 13 1 10 9 13 13 1 9
27 3 13 15 16 16 12 13 1 15 1 10 9 1 15 9 15 3 13 13 15 1 10 9 15 10 1 9
16 3 3 13 12 7 12 13 1 10 15 9 3 13 1 0 15
6 3 13 10 11 13 15
2 1 3
4 13 15 10 11
9 3 13 15 1 3 7 1 3 12
10 13 3 15 13 13 12 15 9 12 9
22 3 13 3 15 13 13 15 10 9 13 7 10 9 7 10 9 7 15 15 13 7 13
8 13 3 10 9 0 13 15 13
7 13 1 15 7 15 13 15
14 13 3 10 9 10 9 0 13 15 7 10 9 13 15
4 13 16 15 13
8 13 3 10 9 15 13 15 13
14 15 3 3 13 7 13 13 15 1 9 16 13 10 13
18 13 3 10 9 15 10 13 13 3 7 13 13 10 9 15 15 10 13
8 3 13 15 10 9 15 13 15
11 9 0 15 10 9 0 13 15 16 13 15
13 3 13 3 15 13 10 9 15 3 3 15 15 13
16 7 13 10 9 15 13 15 10 9 16 15 13 15 10 13 15
23 7 13 16 13 10 11 10 9 0 13 1 10 11 7 13 1 10 9 10 11 1 10 11
9 7 13 15 10 9 13 15 7 13
9 3 13 13 10 9 15 1 15 9
4 15 3 13 13
12 3 13 16 10 13 1 9 0 7 0 13 15
2 7 13
21 1 0 13 9 10 9 7 10 9 7 13 10 9 15 7 13 10 12 1 9 12
7 3 3 13 12 7 9 12
9 15 3 11 13 13 9 9 7 13
3 13 15 16
11 11 1 10 9 15 13 15 13 10 9 15
6 1 9 3 3 13 3
17 13 3 15 16 15 3 13 10 9 15 3 1 9 7 13 0 13
4 13 15 10 9
13 16 3 13 10 9 10 9 1 10 9 3 13 13
4 15 3 13 15
28 13 3 9 15 1 9 9 13 3 7 13 9 15 13 1 10 9 7 13 9 15 13 15 1 10 9 10 9
4 10 13 13 13
11 3 13 15 9 16 10 9 13 15 7 13
5 10 3 9 13 15
5 10 3 11 13 15
10 13 10 9 7 3 13 15 13 1 15
8 10 3 0 13 10 9 10 9
7 7 13 10 9 15 13 3
4 15 3 13 15
6 15 15 13 1 10 0
4 12 13 10 0
10 16 3 13 1 10 9 13 13 10 9
1 15
1 13
4 10 3 11 13
4 13 15 10 9
3 15 3 13
4 13 15 10 11
21 16 13 0 13 13 13 15 10 13 7 13 0 7 13 9 1 9 7 6 13 15
6 13 3 10 9 13 13
5 13 3 13 9 0
7 10 3 11 13 10 9 15
19 3 3 13 15 16 0 13 9 1 9 9 13 3 0 1 10 9 10 9
7 13 3 10 9 13 3 13
6 13 3 10 11 13 15
10 1 9 0 0 13 1 3 9 0 15
6 3 13 10 11 13 15
7 6 15 13 15 7 13 15
4 15 3 13 15
33 6 13 15 16 15 10 13 15 1 10 9 3 13 10 9 10 9 1 9 9 15 13 3 0 1 12 9 13 10 12 9 10 11
27 7 15 15 13 9 7 9 7 9 7 9 7 9 7 9 7 9 1 10 15 9 0 13 7 9 0 13
8 0 3 13 0 0 7 0 0
15 13 3 1 10 9 1 9 10 9 13 15 1 10 9 15
15 7 13 1 0 9 13 0 13 1 10 9 0 7 0 13
13 13 3 15 1 10 9 7 15 3 13 0 13 15
3 15 3 13
11 1 3 10 0 13 13 0 13 7 13 15
7 15 3 13 0 10 9 0
2 13 15
4 16 15 15 13
6 13 3 15 1 10 9
11 0 3 13 13 10 9 10 9 10 9 15
14 13 10 9 7 13 10 9 13 1 10 0 1 10 0
8 13 3 10 0 13 16 0 13
7 7 13 10 1 9 3 15
7 13 3 13 1 10 9 13
20 0 10 0 12 9 13 7 0 15 15 13 10 13 10 9 10 9 7 10 9
6 15 3 13 12 15 13
4 3 9 13 15
5 13 10 15 7 13
10 7 3 13 15 15 13 13 1 10 15
10 7 10 9 15 0 13 16 15 0 13
9 3 13 10 0 0 7 10 0 0
17 7 13 10 11 1 11 13 10 12 1 0 7 1 10 9 13 15
19 6 13 1 11 7 10 9 10 9 13 10 9 7 9 7 13 15 1 9
17 7 13 15 10 9 1 10 13 7 13 7 13 7 10 0 9 13
4 15 3 13 15
2 13 15
20 13 16 13 0 10 12 9 15 12 1 0 7 12 1 0 15 1 10 9 15
5 13 3 10 11 13
4 3 13 15 13
8 13 13 10 9 15 15 13 13
2 13 15
1 13
21 10 3 13 1 0 15 7 1 0 3 13 15 0 13 7 15 13 1 10 9 15
9 13 3 10 12 13 1 10 12 9
6 10 3 11 13 15 13
13 13 16 10 9 10 9 13 15 7 10 0 13 15
5 3 3 13 1 15
22 7 15 3 13 1 15 0 13 13 15 9 7 15 3 13 1 15 13 0 13 15 9
18 3 10 9 10 9 3 13 13 7 13 7 13 10 9 15 9 1 0
9 7 13 15 1 11 13 15 9 0
4 13 15 9 11
7 10 3 9 13 15 16 13
5 15 3 0 13 13
5 9 13 15 9 11
8 7 13 10 11 13 15 7 13
4 15 13 13 15
2 13 15
6 9 16 13 10 9 15
16 13 1 10 9 10 1 15 7 3 13 9 13 7 9 1 15
3 13 13 15
13 7 16 15 15 13 15 13 16 10 9 15 9 13
4 3 3 13 15
11 0 3 13 16 13 10 13 1 10 9 13
4 13 10 9 11
16 6 10 9 15 13 15 0 7 13 1 9 7 1 9 9 9
11 10 3 0 9 13 15 10 9 1 10 9
11 10 3 9 10 13 15 7 10 13 13 13
14 6 10 9 11 13 10 13 1 9 9 6 1 10 0
10 7 13 15 1 11 13 15 10 9 13
3 15 13 0
4 10 3 9 13
10 0 13 10 9 11 10 1 11 10 11
1 13
6 10 9 15 9 9 13
12 7 13 15 0 7 0 1 10 9 7 13 15
29 13 3 10 9 7 10 9 10 0 15 13 7 10 9 10 13 1 10 9 7 13 6 10 9 11 13 7 13 15
4 13 15 0 13
5 10 3 11 13 15
1 6
12 7 13 15 13 1 10 9 1 11 7 13 3
7 3 3 13 1 10 9 13
22 7 13 9 12 1 10 9 13 1 15 7 15 13 1 15 3 3 9 0 7 13 15
5 7 13 3 10 9
6 7 13 10 9 13 13
5 3 3 13 10 9
6 13 3 10 11 13 15
26 16 13 9 7 3 13 3 0 10 10 9 13 7 3 16 10 9 0 13 13 7 13 1 10 9 13
10 7 15 15 3 13 1 10 9 13 13
17 7 13 15 1 10 9 13 15 13 10 9 7 10 0 10 9 13
5 1 15 9 0 13
6 13 3 10 11 13 15
19 13 15 3 15 9 12 15 16 13 15 3 15 15 13 1 15 9 0 13
11 10 9 10 11 3 13 1 9 7 1 9
6 16 13 1 9 13 15
6 1 15 3 3 13 15
8 16 3 13 1 9 13 10 9
7 15 3 3 9 13 10 11
5 7 13 10 11 13
4 13 15 7 15
9 3 15 13 15 1 15 9 0 13
4 9 13 9 12
4 13 10 0 13
7 9 13 3 13 1 10 9
4 15 3 13 13
2 3 13
3 0 13 13
4 15 3 13 13
3 7 3 13
9 15 1 10 12 13 10 9 10 9
1 13
2 10 0
4 13 15 10 11
16 6 13 15 16 10 9 7 10 9 13 15 1 10 9 10 9
12 13 3 11 1 15 1 9 9 7 3 13 15
3 0 9 13
24 9 13 9 15 13 9 7 9 15 13 7 13 1 15 9 7 13 9 7 13 15 9 7 13
18 16 3 13 10 9 10 9 13 10 9 15 1 10 9 13 10 9 15
16 7 13 10 9 10 9 15 15 3 13 15 3 13 15 3 13
11 3 13 0 9 0 10 0 7 13 15 3
9 0 3 13 1 15 10 9 15 13
4 13 10 9 15
9 10 3 9 13 10 9 13 1 15
8 6 13 15 7 13 10 9 15
9 7 13 15 13 1 10 9 7 13
12 3 3 13 10 9 10 9 15 13 10 9 0
2 13 15
19 0 3 13 15 7 10 9 13 0 9 15 13 15 10 9 1 10 9 15
4 13 15 10 11
5 3 13 1 10 9
10 9 15 13 10 13 0 13 1 9 9
15 13 3 10 9 7 10 9 10 9 15 13 16 1 15 13
12 7 13 15 13 13 10 9 16 1 9 15 13
10 7 13 10 11 3 13 1 9 15 13
13 13 10 9 10 9 9 9 15 13 9 10 9 15
15 7 13 10 9 15 13 10 13 1 10 9 7 3 13 13
5 3 13 0 9 13
3 13 10 13
10 10 9 15 7 10 0 13 7 15 0
16 15 3 13 13 15 3 1 10 0 9 15 3 1 10 9 15
10 10 3 0 13 10 9 15 13 7 13
18 10 3 9 13 7 13 10 9 15 13 10 9 0 7 10 9 15 13
5 3 13 10 9 15
5 10 3 9 0 13
6 10 3 13 3 13 0
21 7 13 10 9 0 1 10 9 13 15 15 13 0 7 7 0 7 13 10 9 13
14 13 3 10 9 13 10 13 13 3 9 3 13 9 9
8 9 3 13 3 3 13 9 9
3 15 3 13
6 3 10 9 13 10 9
12 13 15 9 7 9 13 15 1 10 9 10 0
9 3 13 10 9 7 10 9 10 9
11 3 13 10 9 9 13 16 15 13 1 9
10 7 13 15 10 9 15 1 10 9 13
19 9 13 16 0 13 7 10 9 10 9 1 9 13 7 3 13 15 1 15
6 13 3 15 15 15 13
6 13 13 9 9 7 3
8 13 3 10 11 10 9 15 13
4 15 15 13 9
5 15 3 13 15 9
5 7 13 15 10 11
7 15 10 9 0 7 10 9
1 13
3 3 13 15
11 13 3 10 9 9 7 10 10 9 10 9
7 7 13 13 7 13 15 13
3 9 11 13
19 16 15 13 3 13 9 13 10 9 15 10 9 15 7 13 9 10 9 15
22 13 3 1 15 12 9 7 10 0 13 13 7 3 13 9 13 10 9 15 10 9 15
10 3 7 10 0 7 10 0 1 10 12
6 0 3 15 13 10 9
4 15 3 13 15
6 13 3 10 11 13 15
16 1 3 10 9 7 13 7 13 7 3 9 9 1 10 9 13
15 1 3 10 9 10 0 3 13 10 13 15 1 10 9 13
13 15 13 10 9 11 7 10 9 11 7 10 9 11
6 3 13 9 0 7 13
9 7 13 10 9 13 1 10 9 15
20 10 3 9 13 16 13 10 9 13 1 10 15 7 13 12 1 15 0 13 15
4 15 3 13 15
7 0 13 10 0 7 0 9
3 0 0 15
6 13 10 3 15 3 15
12 1 0 10 12 9 0 10 9 13 7 10 9
9 13 3 10 9 13 15 10 11 13
6 15 15 13 1 10 11
3 15 9 13
2 13 15
9 3 3 11 1 9 13 9 15 13
5 13 9 10 9 15
14 13 1 0 15 16 3 13 10 0 15 1 10 9 15
10 16 3 11 13 15 9 3 9 15 13
16 7 15 13 13 15 9 7 13 15 1 0 10 9 13 15 3
11 3 10 11 13 10 9 7 10 9 15 13
10 1 10 11 9 13 10 9 7 10 9
5 13 3 7 3 13
11 13 3 9 0 7 13 1 10 9 10 9
9 0 3 10 9 15 3 13 13 15
11 15 3 10 9 15 13 1 10 13 10 9
9 13 3 10 9 15 7 13 10 9
25 13 3 10 9 1 10 9 7 10 9 1 10 9 7 10 9 1 10 9 7 13 1 10 9 9
5 15 3 3 13 9
6 12 3 13 15 10 9
8 12 3 13 15 10 9 10 0
10 7 13 9 16 9 15 13 12 10 11
7 10 3 0 15 13 15 9
10 15 3 13 15 13 7 15 13 15 13
16 6 3 15 9 7 9 9 16 13 10 9 10 9 1 10 9
9 15 3 3 13 7 10 13 13 13
25 6 15 9 7 9 9 16 13 10 9 7 10 0 13 12 9 7 3 13 13 15 9 11 0 15
8 15 3 13 1 10 9 15 13
16 0 7 0 15 3 0 13 10 9 7 10 9 10 13 10 9
1 7
8 15 3 13 1 10 9 15 13
11 15 3 3 13 1 10 9 10 1 15 13
13 0 15 3 0 10 9 7 10 9 10 13 10 9
15 10 3 13 1 10 9 13 1 15 7 1 15 10 1 15
18 7 10 13 1 10 9 13 1 10 9 10 9 7 1 10 13 1 15
30 6 15 9 7 9 9 16 13 10 9 7 10 9 7 10 9 7 13 10 0 10 9 10 9 7 10 9 7 10 9
10 9 0 10 13 10 9 10 3 9 13
22 6 15 9 7 9 9 16 13 10 1 10 9 7 10 9 3 3 13 1 9 7 9
15 9 0 13 0 10 1 10 9 16 13 3 10 1 15 0
23 6 15 9 7 9 9 16 13 9 13 15 3 3 13 0 3 3 13 9 0 7 15 9
9 3 3 15 3 3 13 10 9 0
20 6 15 9 7 9 9 16 13 10 9 10 9 7 13 10 9 10 0 7 13
18 16 13 1 10 9 10 9 15 3 3 13 9 15 1 10 9 10 9
10 3 13 15 16 9 13 10 13 10 9
10 9 9 9 3 13 1 10 9 10 11
12 1 0 6 15 13 1 15 9 7 0 7 9
19 1 15 13 7 13 7 1 15 13 1 10 9 15 7 13 1 9 1 9
31 3 13 1 15 15 9 0 13 1 10 9 1 10 9 11 10 0 1 10 9 11 9 11 15 13 1 10 9 7 10 9
7 13 0 15 1 10 9 0
31 11 11 10 13 10 9 7 13 10 13 1 15 3 13 13 10 9 15 15 9 9 13 10 9 15 1 10 9 7 3 13
7 6 13 15 10 9 15 0
3 13 3 15
6 13 10 13 1 9 9
19 7 13 10 11 1 10 9 13 7 13 10 9 15 13 15 10 9 10 9
5 15 3 13 13 15
3 6 13 15
10 3 3 13 3 9 1 9 15 3 13
15 13 3 15 1 10 9 10 9 13 15 10 9 1 0 13
2 13 15
14 3 0 13 7 15 10 9 10 15 9 7 9 10 9
5 13 3 15 15 13
8 0 3 13 1 10 9 15 13
3 7 0 13
7 13 3 13 9 7 9 9
1 13
2 3 13
8 13 3 13 7 3 13 10 9
16 13 3 9 1 9 7 9 1 9 7 13 9 7 9 1 9
19 3 13 15 1 9 7 13 15 7 13 13 1 15 10 9 1 10 9 15
7 7 0 9 13 7 13 0
11 7 1 10 13 10 9 13 10 9 10 0
7 10 3 13 1 9 0 13
21 7 13 0 10 9 10 9 1 0 10 9 1 9 15 10 9 7 3 13 10 9
53 3 3 13 10 9 10 9 10 13 1 11 10 9 13 1 9 0 10 13 13 3 10 1 10 11 13 1 10 9 10 1 10 9 3 13 13 10 1 10 9 15 7 10 1 10 9 3 13 3 13 10 9 15
13 6 3 10 1 9 13 7 10 13 1 0 10 9
11 13 3 16 3 13 10 9 15 9 7 9
8 1 3 10 0 13 10 9 0
13 3 16 15 15 13 6 3 10 11 7 3 3 13
18 13 3 9 7 9 7 13 9 0 7 9 16 13 16 0 3 10 0
3 6 13 15
11 16 3 13 15 6 1 10 0 13 3 13
4 6 1 10 9
2 3 13
19 3 3 10 9 13 1 9 7 13 1 9 3 13 10 9 10 9 10 9
32 3 3 1 10 9 10 9 0 10 9 13 7 10 9 3 13 10 9 15 7 10 9 13 1 10 9 7 10 9 10 9 13
35 7 3 13 10 9 10 9 10 9 1 9 7 13 15 10 9 10 9 7 13 10 9 10 9 13 1 10 9 10 9 1 9 7 9 0
23 7 13 10 9 15 1 9 0 7 13 10 0 15 1 10 12 9 1 9 9 1 9 15
7 1 3 10 9 13 10 9
16 3 3 10 9 15 13 0 7 10 9 13 13 16 3 10 9
13 3 3 15 3 13 0 15 13 16 3 13 1 9
3 6 13 15
11 3 3 13 10 9 0 16 3 15 0 13
22 1 3 10 9 0 7 9 15 13 7 10 9 10 9 7 10 9 3 3 10 9 0
14 3 3 10 9 10 11 3 13 10 9 10 9 10 9
43 3 3 13 1 10 9 10 1 10 9 13 7 13 13 7 13 1 15 9 13 11 1 10 9 7 3 13 16 13 10 9 7 13 0 3 13 7 10 9 10 9 10 9
6 3 13 12 1 10 9
5 12 13 7 12 13
5 12 13 1 10 9
5 12 13 7 12 13
23 0 3 13 16 16 13 10 9 15 9 10 9 13 13 3 7 3 3 13 13 10 9 15
23 15 3 13 10 0 9 7 0 15 13 10 9 1 10 9 15 10 13 15 10 9 1 9
12 0 10 9 0 15 13 10 9 15 13 3 13
11 6 13 15 16 1 15 10 13 15 13 15
55 16 3 13 10 0 9 1 10 9 15 13 15 10 9 7 13 13 10 9 15 13 3 7 13 1 10 13 13 10 9 10 9 0 1 9 15 3 13 7 1 9 15 3 13 7 13 15 7 10 9 15 1 10 9 13
9 3 13 10 9 7 10 9 10 9
18 3 13 10 9 10 9 12 9 15 13 10 9 15 13 1 9 10 9
11 10 3 0 13 10 9 3 13 1 15 9
12 10 3 0 13 9 1 10 9 1 10 9 15
5 0 3 9 9 13
3 6 10 9
3 13 1 9
11 3 13 15 10 9 0 7 13 10 9 15
6 10 3 0 10 0 13
5 13 3 10 0 13
6 3 3 13 15 7 15
8 13 3 1 10 13 7 13 15
8 0 3 13 3 10 0 9 13
4 9 9 13 15
4 15 3 13 13
3 6 13 15
10 13 3 16 3 13 10 9 7 10 9
33 3 3 9 13 13 10 0 9 7 13 15 10 13 15 7 15 3 13 12 9 15 3 12 15 3 12 0 1 10 0 9 7 13
15 3 13 10 10 12 9 13 13 1 15 7 13 0 12 9
7 3 10 10 12 13 0 12
15 1 3 0 9 13 10 9 10 9 0 7 13 9 1 15
12 7 13 10 10 12 9 13 13 0 12 9 13
5 9 12 9 15 13
4 0 12 9 13
5 13 15 10 9 15
9 3 9 0 7 0 1 0 13 0
4 1 0 15 13
7 13 1 10 9 10 9 15
5 9 12 9 15 13
1 13
5 13 15 10 9 15
9 3 9 0 7 0 1 0 13 0
4 1 0 15 13
7 13 1 10 9 10 9 15
9 13 3 3 10 10 12 9 13 13
16 9 13 15 16 0 13 9 13 3 3 13 7 13 3 3 13
1 13
7 13 3 10 9 15 13 15
15 0 9 7 0 13 16 13 3 3 13 7 13 3 3 13
18 13 15 3 13 10 9 15 10 9 7 13 15 13 3 10 15 1 9
13 13 3 1 15 10 9 7 13 10 13 10 12 9
7 10 3 13 15 13 7 13
10 10 3 3 13 3 15 13 13 1 15
10 7 10 0 9 13 1 10 9 10 0
34 7 13 1 15 15 10 9 7 13 15 1 15 3 10 9 13 10 9 1 10 9 7 13 10 3 9 1 0 15 10 3 9 1 0
8 3 13 10 9 10 1 0 15
1 6
13 10 13 10 9 15 13 10 13 15 9 1 9 9
6 13 3 7 13 15 13
4 13 7 13 15
5 0 13 7 13 15
4 0 7 13 15
7 1 9 13 7 13 1 15
6 3 13 15 10 0 13
7 9 3 15 13 13 7 13
4 7 13 7 13
7 3 3 15 13 0 7 13
4 7 0 7 13
12 3 3 15 13 13 7 1 9 7 13 1 15
6 7 13 10 9 13 15
6 3 13 7 10 1 0
17 13 1 15 13 1 10 9 10 0 10 13 10 9 7 10 9 15
7 13 3 7 3 13 15 13
5 13 7 3 13 15
6 0 13 7 3 13 15
5 0 7 3 13 15
8 0 7 1 9 7 3 13 15
20 9 3 15 13 13 7 13 7 0 7 0 7 0 7 1 9 7 3 13 15
3 6 13 15
11 1 15 3 13 12 0 10 0 3 15 13
12 7 13 0 1 9 0 10 3 0 1 9 0
14 7 13 16 13 10 11 15 10 9 0 13 10 9 15
17 13 16 1 12 9 10 9 13 7 10 9 10 9 13 1 10 13
17 3 13 10 9 7 10 0 10 9 1 10 9 10 9 10 13 11
2 13 3
11 3 1 10 9 16 3 9 13 1 10 9
6 13 3 10 9 13 13
5 1 15 10 9 0
8 13 3 0 13 0 7 13 0
6 13 3 10 11 13 15
5 15 9 13 10 9
7 3 3 10 0 13 1 15
5 15 3 3 3 13
15 13 3 0 10 9 0 1 10 9 15 1 10 13 15 13
18 3 3 13 10 9 0 1 0 10 9 13 3 15 13 0 1 9 15
13 3 13 12 10 12 10 13 11 11 1 10 9 13
9 15 13 15 13 7 15 15 13 15
6 15 3 13 15 12 9
11 10 3 0 10 0 13 10 9 10 11 13
7 3 13 13 15 13 10 9
3 15 3 13
7 13 1 10 9 1 10 0
3 10 9 13
5 10 9 15 3 13
9 1 15 13 10 9 1 10 9 15
4 7 13 10 9
8 0 3 13 13 1 10 12 9
4 7 13 15 13
9 6 13 15 16 12 1 15 13 15
8 7 13 3 13 13 15 12 0
4 15 3 13 13
12 10 13 1 15 10 9 1 10 9 0 15 13
12 6 3 10 9 0 1 15 10 9 10 9 13
9 0 13 15 16 3 13 10 9 0
7 13 3 11 10 13 15 13
4 3 15 13 9
2 13 15
2 15 13
5 7 13 10 9 13
1 13
5 0 13 10 9 15
8 7 13 9 7 13 13 15 13
4 13 1 15 15
15 0 3 13 10 9 15 10 9 10 1 0 13 1 9 9
3 13 3 15
27 3 3 13 1 3 1 0 10 9 10 9 1 10 9 0 3 15 13 1 15 0 1 10 9 10 9 15
9 15 15 13 1 15 1 10 9 0
2 13 3
9 13 10 9 7 13 10 9 10 9
10 1 3 10 13 15 13 15 1 10 11
6 13 3 10 11 13 15
8 16 15 13 1 15 15 3 13
4 13 15 10 11
14 6 13 15 16 1 0 10 9 16 9 13 3 13 15
11 3 16 13 15 1 15 13 3 3 15 13
6 3 7 15 10 9 13
14 3 13 1 15 10 11 1 9 13 11 7 13 10 9
7 13 3 1 15 13 3 13
13 7 13 10 11 7 10 12 9 11 13 13 7 13
3 3 13 15
7 0 13 10 9 15 1 9
6 13 3 7 13 1 15
8 3 3 3 15 13 7 3 15
13 7 13 1 10 9 7 13 15 13 7 13 10 11
8 3 3 13 12 9 13 1 15
8 13 7 13 16 3 13 1 9
4 10 3 9 0
4 10 3 9 0
6 3 1 0 13 13 13
6 7 13 3 13 15 13
13 7 13 15 3 13 13 1 0 10 15 9 13 3
8 3 13 1 10 9 7 13 15
5 13 10 0 7 13
13 6 13 10 9 7 10 9 10 9 13 1 9 0
1 13
1 13
26 7 3 15 13 6 11 12 10 12 13 7 1 15 9 0 1 9 7 9 1 10 9 7 0 10 9
8 10 3 13 15 13 15 9 13
2 13 15
6 7 3 13 10 11 13
2 13 9
3 7 13 15
5 10 3 11 13 15
11 3 13 13 10 9 1 10 11 7 13 15
23 7 6 12 10 1 11 13 10 9 13 10 9 15 7 13 10 9 10 9 13 15 10 9
5 3 13 15 10 11
8 15 3 10 13 9 1 9 13
17 7 13 16 3 13 13 10 9 15 7 13 15 3 0 12 9 9
9 3 3 13 10 9 16 3 13 13
9 1 0 10 9 13 10 11 10 9
11 1 9 1 10 9 13 13 7 3 13 15
10 0 3 0 13 16 13 10 9 10 9
7 3 10 9 15 13 15 13
17 15 3 13 10 11 13 1 11 10 9 3 10 9 7 10 0 13
21 10 3 9 7 10 9 0 13 9 1 10 11 16 15 13 7 3 13 0 13 9
5 0 3 13 12 13
2 0 13
6 7 13 10 9 13 15
2 15 13
4 15 0 15 13
4 10 3 11 13
6 7 13 10 9 13 15
4 13 15 10 11
2 15 13
19 1 3 13 10 9 10 9 13 1 0 10 9 7 13 1 10 9 10 9
8 3 10 9 13 10 9 15 13
1 13
5 15 3 9 13 9
5 13 3 13 10 9
3 15 15 13
3 0 9 13
4 15 3 13 13
2 13 15
6 11 15 13 10 13 15
8 10 3 11 13 3 1 10 9
6 7 13 15 12 9 13
7 3 15 13 1 11 10 0
6 15 3 13 1 15 13
6 0 13 1 11 10 0
6 7 3 13 1 9 16
4 3 13 10 9
9 1 0 3 13 10 13 13 10 11
6 3 3 15 1 15 13
8 7 3 10 9 15 0 15 13
6 3 13 13 7 13 16
4 3 13 10 9
9 7 13 10 11 10 9 11 13 16
6 16 9 13 3 13 15
5 7 13 3 13 3
19 9 3 13 9 13 15 10 9 7 10 0 10 9 1 10 11 16 13 15
9 7 13 15 13 7 13 11 10 9
18 3 13 11 10 13 15 16 13 13 13 10 12 9 10 9 7 0 13
4 13 13 9 0
3 15 3 13
11 7 13 10 9 1 10 9 13 7 13 13
7 10 3 9 13 10 9 13
11 3 13 13 15 1 10 9 16 9 9 13
14 9 3 13 13 1 15 10 9 10 9 1 9 10 0
10 3 13 10 9 0 9 9 1 10 3
9 3 13 10 13 1 11 10 9 13
26 7 13 10 12 9 10 9 10 13 15 13 1 9 11 7 13 15 1 10 9 10 9 3 13 15 9
6 7 13 15 10 9 13
4 10 3 11 13
2 15 13
12 7 1 10 13 15 1 10 9 7 0 15 13
5 3 13 15 10 11
5 3 13 15 15 13
13 7 3 13 15 1 3 12 9 16 13 10 9 3
7 13 3 3 9 0 13 11
7 13 3 15 13 15 10 11
7 13 3 16 1 9 13 15
13 13 3 15 1 10 9 13 1 15 10 9 15 13
6 15 15 7 10 0 0
8 0 3 13 3 1 9 1 15
6 13 3 10 9 13 15
3 15 3 13
2 10 11
4 13 15 10 11
2 13 15
1 13
3 15 3 13
4 15 3 0 13
1 13
20 13 3 10 11 16 15 13 7 3 9 13 13 9 13 10 9 1 10 9 13
6 0 13 1 10 9 0
2 15 13
10 10 9 15 1 15 7 1 10 9 15
5 3 13 15 10 11
7 10 3 11 13 13 16 13
30 7 13 15 9 0 13 15 7 13 9 1 9 13 1 10 9 15 7 9 1 10 0 15 7 13 1 15 13 15 13
5 13 10 9 10 0
13 7 13 1 15 13 10 9 7 13 1 10 9 15
19 7 16 13 15 13 15 10 9 13 15 10 9 15 7 13 15 1 10 13
7 13 3 13 9 0 9 11
18 7 13 1 9 13 11 15 13 9 9 13 13 15 13 9 1 9 13
5 7 13 3 13 13
10 7 13 1 10 9 15 10 9 15 13
7 0 13 11 10 9 10 0
13 3 13 1 15 12 9 12 1 0 7 12 1 0
11 10 3 13 13 15 13 10 9 15 7 13
21 10 13 10 9 7 1 12 9 13 13 15 16 9 13 10 9 7 13 1 10 9
10 3 10 9 13 1 10 9 7 0 13
4 15 3 13 13
9 13 3 1 10 9 7 13 1 15
4 13 1 10 9
5 13 3 16 13 15
3 13 3 16
3 9 13 9
12 10 3 15 7 10 9 10 13 1 15 13 15
13 1 3 0 9 9 13 1 15 10 9 1 9 0
2 0 13
7 9 15 9 15 3 15 13
8 15 3 10 3 13 13 13 16
3 11 13 0
17 7 3 13 12 1 15 7 13 9 13 7 9 7 13 9 13 15
4 10 3 0 13
1 13
6 13 16 13 11 13 15
31 7 6 10 9 10 9 13 3 1 3 1 12 7 10 9 13 7 10 9 13 7 10 9 13 7 0 9 10 13 0 13
17 7 13 1 10 9 1 10 9 15 13 1 10 0 9 7 13 0
19 10 3 9 7 10 1 15 13 10 11 13 10 9 7 10 13 13 3 13
5 3 9 9 13 0
17 13 3 3 9 0 1 3 13 15 13 10 11 1 10 11 13 15
20 1 15 13 11 10 9 7 11 10 10 11 7 11 9 7 10 9 10 9 11
17 0 3 13 13 9 0 1 11 10 9 11 15 3 0 13 10 11
9 0 13 10 11 13 10 9 10 11
14 13 3 3 11 10 9 7 10 0 11 13 1 10 9
17 10 3 3 15 13 1 10 9 13 10 9 7 10 9 1 11 13
9 9 13 16 0 10 0 13 3 13
4 1 12 9 13
19 13 3 13 10 9 1 10 0 9 16 13 10 9 13 15 7 13 10 9
4 13 1 10 0
8 7 13 10 0 9 0 10 0
2 13 9
3 13 3 13
12 15 3 13 13 10 9 13 10 9 1 10 9
19 3 3 9 10 13 1 12 9 13 11 10 9 7 10 0 11 13 10 9
5 7 6 9 13 0
15 9 3 9 13 1 9 7 13 13 10 9 7 13 1 15
14 13 3 10 9 15 3 9 7 10 9 15 0 3 9
7 13 3 10 9 13 10 9
3 3 13 15
3 3 13 3
4 13 3 3 13
6 6 13 10 9 3 13
8 7 0 13 13 10 9 15 16
11 13 1 10 0 7 6 13 15 1 10 11
3 6 13 15
16 7 13 0 1 10 9 1 9 7 9 0 13 13 10 9 15
6 7 6 11 13 15 13
10 15 3 13 13 15 10 9 7 13 15
5 3 13 15 10 11
2 3 13
1 13
17 13 3 15 6 15 10 9 13 1 10 9 13 10 9 0 10 13
14 7 13 1 10 0 9 7 13 9 0 13 10 9 13
11 13 16 10 9 15 9 13 13 15 15 13
13 7 16 13 0 1 10 9 15 13 7 15 0 13
10 7 13 10 9 0 1 0 1 10 3
20 10 3 12 9 13 1 10 11 1 10 9 3 13 15 10 11 7 13 15 13
3 15 3 13
9 13 15 15 9 1 9 7 1 9
26 13 13 15 10 9 13 15 1 10 9 10 9 7 10 9 7 10 0 9 13 15 13 15 15 13 15
14 7 6 15 1 15 13 15 10 9 1 10 9 10 9
12 9 10 9 11 11 3 13 1 10 11 10 9
14 6 15 13 10 9 15 1 9 15 15 13 10 9 15
4 13 10 9 9
5 0 13 10 9 15
24 7 13 1 15 15 10 0 9 7 10 9 15 7 13 1 15 1 10 11 9 13 10 9 15
20 7 13 10 11 13 9 9 7 9 0 1 10 9 15 7 13 9 7 9 0
3 7 13 13
17 13 10 0 15 1 15 15 3 13 0 13 13 10 9 10 9 15
4 15 13 15 9
7 0 3 13 15 1 9 0
18 7 3 13 1 10 9 13 13 10 9 7 10 9 3 9 13 1 15
7 15 13 10 9 15 10 0
3 1 15 13
9 7 3 10 9 15 13 1 10 9
21 7 13 1 10 9 12 9 13 1 10 11 7 13 1 10 9 7 10 9 13 15
27 1 3 10 13 10 11 13 10 11 1 10 11 13 10 9 10 9 16 13 10 9 7 13 10 9 10 9
6 13 7 13 1 10 9
18 7 13 1 10 9 10 11 13 11 7 11 10 9 11 13 1 10 9
9 6 1 15 7 13 15 13 9 9
7 7 3 13 10 9 13 15
25 7 13 0 13 11 10 10 11 7 11 10 9 15 7 15 1 10 9 13 10 9 7 3 13 15
15 7 13 10 9 15 11 1 10 9 1 10 9 13 1 15
4 7 13 1 11
8 7 3 10 9 13 1 10 9
6 7 13 1 10 9 15
12 13 3 13 15 3 9 13 7 3 3 10 9
6 15 15 7 15 11 9
3 13 13 15
4 13 15 15 13
4 10 0 10 9
5 7 13 15 10 11
5 13 7 13 1 15
14 7 13 15 10 9 10 0 7 13 9 0 13 1 15
7 7 13 0 16 13 15 13
9 3 10 9 10 0 13 7 13 15
13 7 13 10 9 15 3 3 1 0 10 9 10 11
17 7 3 1 10 9 13 13 1 10 9 11 7 11 1 11 7 11
12 10 3 9 11 13 13 7 3 13 15 1 15
7 7 13 13 15 13 10 9
8 7 13 15 10 9 7 13 15
17 0 3 13 16 13 10 9 13 1 15 15 10 3 13 7 10 13
20 7 13 0 3 13 0 9 7 9 0 13 7 3 13 13 10 9 16 13 15
15 7 13 15 11 7 10 1 15 7 13 15 7 13 15 16
3 15 13 15
3 7 13 15
10 13 3 1 10 13 9 16 3 3 13
4 1 0 3 13
15 7 13 13 1 10 9 15 1 0 10 11 7 10 9 13
5 16 13 13 15 13
9 7 13 13 10 9 15 13 7 13
1 13
9 7 3 13 1 15 10 9 7 13
9 7 13 15 3 13 15 7 13 15
22 13 15 15 13 7 13 15 13 10 9 7 13 1 10 9 15 15 13 11 1 9 15
29 15 3 13 13 13 0 7 13 10 9 16 3 15 13 1 9 3 13 7 3 1 0 9 13 7 13 1 15 3
16 7 13 0 16 3 13 7 10 1 10 9 7 13 15 10 9
9 7 13 13 1 15 0 13 1 12
22 7 3 13 13 15 1 10 9 13 10 9 3 13 7 13 13 10 9 3 10 0 13
5 9 13 15 10 9
13 13 3 15 10 9 3 13 7 13 1 10 9 15
4 15 0 3 13
1 13
15 7 3 13 10 11 10 9 15 16 3 13 1 15 13 15
7 15 0 13 1 10 9 15
20 15 13 0 13 10 0 13 15 10 9 7 13 13 7 13 10 9 15 7 13
18 16 3 13 16 9 13 10 9 10 9 1 10 9 13 9 13 10 0
1 13
10 13 10 9 15 7 13 1 10 9 15
19 7 13 7 3 13 10 9 13 1 15 16 13 15 7 13 10 9 13 16
6 7 13 3 1 10 9
10 7 15 10 9 13 1 15 7 13 15
14 7 13 13 11 10 10 11 13 1 10 9 7 13 15
2 13 15
4 7 13 13 15
10 13 3 0 7 13 15 3 9 10 9
13 7 13 16 13 1 10 9 7 0 13 10 9 15
6 7 13 10 11 13 15
10 3 9 13 10 13 9 7 10 3 13
6 3 13 13 0 7 9
9 7 13 10 9 11 7 10 9 13
5 7 13 7 13 15
17 1 15 10 9 11 7 10 9 10 9 13 10 3 15 9 3 13
14 3 13 10 9 10 9 1 15 10 9 1 15 13 13
16 13 3 9 3 13 1 15 10 9 7 3 13 1 0 10 9
8 15 9 9 0 13 1 9 0
16 16 3 3 13 10 9 1 15 10 0 10 0 7 0 9 13
8 7 15 13 9 0 1 9 0
15 16 3 3 13 10 9 10 9 7 10 9 13 7 10 9
20 7 13 15 1 10 9 13 1 10 0 7 10 9 15 13 9 13 13 10 9
5 7 10 9 13 15
3 7 13 15
15 3 13 15 13 11 16 9 13 7 13 15 7 10 1 15
31 3 13 1 10 9 10 9 1 11 9 7 10 9 10 9 13 15 3 13 13 3 3 10 9 7 13 3 10 1 15 13
3 7 13 15
13 10 9 1 10 9 13 7 3 10 9 1 10 9
10 3 9 13 10 9 10 9 3 10 9
13 7 13 3 1 9 7 13 3 9 13 13 10 9
12 7 13 15 16 1 10 9 13 15 16 13 15
4 13 1 10 0
3 7 13 15
11 13 10 9 0 13 7 13 9 13 7 13
3 15 3 13
15 7 13 15 1 9 13 1 10 9 10 9 15 13 10 9
3 13 10 9
7 7 13 7 13 10 9 15
15 7 13 10 9 3 1 10 9 9 13 1 15 16 15 13
12 0 3 13 16 13 15 16 15 13 15 13 9
14 7 10 9 10 0 3 15 13 13 15 7 13 13 16
6 15 13 10 9 10 9
9 7 0 13 15 16 3 15 0 13
14 7 13 1 10 9 7 13 15 13 15 7 13 1 15
18 7 13 12 16 13 1 15 7 16 13 15 13 7 13 9 13 10 9
10 7 13 10 12 7 13 9 10 11 11
28 7 11 7 11 7 11 7 11 7 11 7 11 10 10 11 7 11 7 11 10 0 7 11 11 15 3 13 15
11 7 13 3 9 16 3 13 15 3 9 13
8 7 13 10 1 15 13 13 15
4 13 3 16 13
21 7 10 9 10 1 11 13 13 16 11 13 7 16 1 10 9 10 9 13 10 9
7 7 13 15 1 9 13 15
5 3 13 11 11 13
12 7 16 9 1 15 13 3 13 10 9 0 13
15 7 16 10 11 13 1 15 13 7 3 13 13 7 9 13
18 6 13 15 16 15 13 10 9 10 9 10 9 7 10 9 15 3 13
20 15 3 3 13 1 10 9 10 0 3 13 9 1 10 9 7 0 13 0 9
2 3 13
3 9 0 13
17 7 13 10 9 15 7 10 9 15 7 3 13 13 1 15 13 15
15 6 10 9 15 7 10 9 15 7 10 9 15 3 13 15
4 7 13 15 13
9 15 13 10 9 15 7 10 9 15
1 13
7 10 9 15 7 10 9 15
15 15 3 13 10 9 10 9 0 9 15 7 9 7 9 13
7 7 3 13 13 1 10 9
13 7 13 15 1 9 0 7 13 15 1 10 9 15
1 13
5 6 13 10 13 13
18 7 13 1 10 13 15 3 13 1 10 9 7 13 10 9 7 13 15
13 7 16 13 10 9 13 7 1 10 3 13 9 13
17 7 15 13 1 10 9 7 13 10 9 7 13 15 7 9 3 13
24 7 15 13 1 10 9 10 0 7 13 9 13 7 13 7 13 1 12 7 1 12 7 1 12
5 15 13 9 13 13
15 7 16 13 1 0 13 15 10 1 15 1 10 12 10 9
3 7 13 15
8 15 10 9 13 10 9 10 9
25 0 3 10 3 1 9 15 13 16 13 13 7 3 13 7 13 13 7 3 13 16 13 7 13 15
11 3 13 10 9 0 7 3 15 10 9 13
5 10 13 10 9 13
38 7 0 3 13 10 1 10 0 13 15 3 13 10 9 3 1 9 13 15 7 3 13 9 1 15 7 0 13 3 13 9 7 9 1 10 9 3 13
8 7 15 13 10 1 10 9 13
29 0 13 10 10 9 13 7 10 9 10 9 7 10 9 10 9 7 10 1 10 0 9 13 13 10 9 7 0 13
26 7 0 13 10 1 10 9 10 0 13 15 13 10 9 7 13 7 13 12 12 7 12 12 7 12 12
17 7 13 15 16 3 13 10 9 16 1 10 9 13 7 1 10 9
6 3 16 1 10 9 13
6 16 15 13 9 13 13
3 13 15 13
9 1 15 9 13 13 15 7 13 15
5 15 3 13 13 15
10 7 15 3 13 3 15 13 13 1 15
2 7 13
31 3 13 10 9 10 9 3 9 13 10 9 1 10 9 7 13 7 13 9 7 9 7 10 9 13 7 13 3 3 13 15
14 0 10 9 13 0 9 3 9 3 0 9 1 10 9
12 3 13 10 9 10 9 7 1 15 15 9 13
43 3 9 9 15 3 13 1 10 9 0 13 15 10 9 10 1 10 9 7 3 13 13 7 13 0 15 10 9 7 13 9 0 16 13 1 10 9 15 10 9 10 9 13
11 7 0 9 0 13 15 10 9 3 13 13
6 1 3 9 3 13 15
8 1 0 3 10 0 9 13 15
9 7 13 15 1 0 10 9 0 13
4 13 1 10 3
17 7 13 10 9 13 15 3 13 1 10 9 7 15 9 13 1 15
10 7 13 15 1 10 9 1 10 9 13
6 7 13 15 7 13 15
6 9 3 13 15 16 13
9 7 13 13 10 9 7 13 10 9
1 13
1 13
8 7 13 10 9 7 13 9 0
3 7 13 15
8 7 13 9 0 7 13 1 15
13 15 3 0 13 16 7 10 9 7 10 9 15 13
12 7 13 1 10 3 10 9 1 10 9 10 0
72 7 13 15 1 10 9 3 13 15 1 10 9 9 1 9 0 15 10 9 13 1 10 9 7 7 9 3 15 13 15 13 1 10 15 3 9 7 9 13 7 13 1 15 10 9 7 10 9 13 7 15 13 15 13 7 3 9 7 9 1 10 9 7 1 10 9 13 13 7 13 15 9
15 7 13 10 11 1 3 13 7 13 15 7 13 9 0 13
10 15 15 7 15 11 9 10 9 10 0
4 13 15 10 9
3 13 3 15
3 7 13 15
3 15 9 15
3 7 13 15
6 9 9 15 16 0 13
11 7 13 15 0 16 3 15 13 1 10 9
10 13 3 3 1 10 9 9 9 0 13
9 13 15 1 10 9 16 1 15 13
3 7 13 15
14 7 10 13 15 13 7 13 1 10 9 7 1 10 9
7 7 13 13 15 13 10 13
19 7 13 1 10 11 7 13 10 13 13 13 7 13 10 13 10 9 7 13
13 7 13 15 10 13 3 13 10 13 7 1 10 9
9 7 13 13 15 13 1 10 9 15
7 7 3 13 15 7 13 15
19 13 1 10 9 15 1 10 15 7 13 15 15 10 9 15 13 7 13 15
16 7 13 7 13 13 1 10 11 15 13 15 10 11 7 15 13
36 7 13 12 10 9 9 11 7 13 15 13 1 10 9 15 7 13 15 0 13 16 10 9 15 3 13 16 13 13 10 9 15 16 13 7 13
12 7 13 1 15 7 13 15 9 0 7 13 15
43 7 9 13 1 9 9 12 9 7 0 13 1 0 9 7 13 10 1 15 15 7 15 13 7 3 1 10 0 13 13 10 1 10 11 13 1 10 9 3 13 10 9 15
3 13 3 16
17 7 3 13 10 9 10 9 15 7 13 10 9 16 13 1 10 9
17 7 3 10 11 13 1 15 10 1 15 9 13 13 1 10 9 13
5 15 15 13 10 9
6 7 13 15 10 9 15
3 15 15 13
6 7 13 13 10 0 13
20 10 3 9 13 7 13 13 15 13 15 13 7 13 15 7 13 15 15 10 9
6 9 10 9 15 13 15
10 13 1 9 7 13 0 1 10 9 15
9 3 15 13 13 1 10 9 13 16
4 10 9 15 13
5 15 3 13 10 9
2 3 13
2 0 13
19 7 13 1 10 9 10 9 7 13 9 7 13 7 13 0 7 13 13 15
4 15 13 7 13
6 10 9 3 13 7 13
3 7 13 15
22 15 3 13 15 13 10 9 10 9 7 10 9 7 10 1 15 7 13 3 13 10 9
8 7 13 10 9 10 9 13 15
4 10 9 15 13
7 7 3 13 10 9 7 13
4 13 3 9 12
5 7 13 3 9 0
13 7 13 15 0 16 15 13 0 7 13 13 15 13
15 7 13 3 7 13 1 10 9 15 7 13 15 10 9 15
8 7 13 9 13 13 1 10 9
6 7 10 0 13 13 13
18 3 0 13 10 9 10 9 10 11 7 9 11 7 11 7 11 7 11
9 7 3 13 10 9 15 3 1 15
4 7 13 1 15
26 7 13 15 10 11 16 3 13 9 0 3 3 1 10 9 15 7 1 10 0 15 7 1 10 9 15
15 7 3 13 3 13 15 9 16 3 0 0 13 10 9 13
6 7 13 1 10 9 15
6 7 13 10 9 3 13
47 7 13 10 12 7 13 15 13 12 12 7 13 15 9 10 9 10 0 7 13 15 16 15 13 1 9 3 3 9 0 3 9 3 9 3 1 10 9 9 7 13 9 7 3 13 12 9
11 3 3 13 1 9 3 13 16 3 13 3
23 7 15 3 9 3 13 15 7 13 15 13 3 13 10 9 10 1 10 9 15 1 9 15
16 7 13 13 16 13 7 9 0 13 7 13 9 0 0 7 13
28 7 13 10 9 11 0 3 13 10 9 15 7 13 16 11 10 13 13 1 0 7 1 0 13 10 9 1 15
6 15 3 13 16 11 13
9 15 3 13 16 9 3 12 10 9
5 13 3 10 11 13
6 15 15 13 11 0 13
9 3 13 15 13 10 9 10 9 15
12 10 3 11 13 15 7 13 15 13 7 3 13
24 10 3 11 13 10 11 13 15 9 0 7 0 7 13 15 7 13 15 0 13 7 3 15 13
37 7 13 9 0 16 11 10 9 15 9 13 10 9 15 7 10 9 7 10 0 10 11 7 13 10 9 15 10 11 7 13 13 10 11 7 10 13
6 10 3 9 13 10 9
8 13 15 15 3 13 7 13 15
4 7 13 15 16
6 7 13 13 10 9 15
3 15 3 13
5 10 9 11 10 13
10 7 13 3 1 9 1 10 9 13 13
12 13 16 3 13 15 1 9 10 9 11 10 9
15 7 0 13 10 9 1 10 9 7 10 13 3 13 13 15
11 7 3 13 10 9 9 13 13 10 9 15
16 7 13 10 9 15 13 7 13 10 9 15 7 13 15 1 9
15 7 13 10 9 1 10 11 7 13 15 15 15 13 7 13
11 6 15 0 1 0 1 0 9 7 13 0
12 13 3 10 13 7 10 13 0 7 7 13 13
9 7 13 1 0 9 10 9 1 0
19 7 13 15 13 7 13 15 0 7 3 1 15 10 9 13 3 7 13 15
21 7 13 13 0 9 7 13 1 15 16 13 3 9 3 13 9 7 13 13 15 0
14 13 15 16 13 1 10 3 9 7 9 13 15 15 13
5 15 3 13 13 15
4 13 15 15 13
9 13 13 9 12 9 7 13 15 13
4 15 3 13 15
3 15 9 13
1 13
3 7 13 13
4 12 7 12 9
11 7 13 15 13 15 9 9 1 10 0 9
9 7 13 9 9 1 12 7 1 12
5 7 13 15 7 13
10 7 13 9 12 9 9 7 1 10 9
8 7 13 10 13 10 9 12 9
8 7 13 15 13 1 10 9 13
16 7 0 13 13 10 9 1 0 10 9 7 0 0 1 10 9
25 7 13 15 13 1 10 13 13 3 10 9 0 15 1 0 9 10 9 13 1 15 13 1 10 9
4 7 13 13 15
14 15 3 13 15 1 10 9 13 13 16 9 13 7 13
9 15 3 3 13 1 15 7 13 15
1 13
2 3 13
11 7 13 1 15 1 10 9 7 13 10 9
7 7 3 1 0 1 15 13
12 3 3 13 1 10 9 7 13 15 10 9 13
10 7 13 1 10 9 13 1 11 7 13
27 7 13 15 1 10 9 3 13 15 13 0 10 9 0 7 13 1 10 9 10 3 13 13 3 13 16 13
6 7 15 3 13 15 13
64 7 13 15 10 9 15 16 0 9 0 13 0 13 10 9 10 3 9 7 15 10 0 16 3 0 13 10 9 3 13 13 10 9 10 0 7 1 9 16 3 13 3 13 7 15 0 13 15 13 13 9 9 7 9 7 9 7 13 15 10 9 7 10 9
18 1 15 3 13 10 9 15 1 10 9 10 0 7 0 9 13 10 9
4 15 3 13 15
25 3 13 11 1 15 10 9 3 13 16 0 10 9 10 9 15 13 10 3 9 15 3 13 1 15
8 3 3 13 15 13 9 9 9
10 13 10 9 10 9 13 10 9 10 9
3 7 13 15
16 13 10 9 15 7 10 9 15 7 10 13 9 7 9 9 13
3 15 3 13
37 16 13 9 10 9 7 10 9 8 15 13 9 15 3 1 15 13 3 13 15 15 13 10 9 7 10 9 13 10 9 10 9 10 9 15 15 13
5 7 0 0 0 13
7 7 13 3 10 9 13 15
5 13 15 15 7 13
12 15 13 1 10 9 13 1 15 15 13 13 15
11 7 10 1 10 9 13 13 10 13 10 9
3 7 13 15
5 3 3 15 0 13
34 3 13 16 15 10 3 13 1 10 9 3 13 15 13 16 3 13 15 1 10 9 7 1 10 9 7 1 10 9 13 13 15 10 9
12 13 3 16 10 1 10 9 13 0 13 10 9
25 3 3 1 10 9 10 9 10 9 10 0 13 9 9 9 9 9 9 9 9 9 0 9 9 9
10 15 0 10 0 3 13 7 13 10 9
8 3 3 13 13 1 10 9 11
11 7 13 1 9 15 13 13 7 3 13 13
11 7 13 15 16 10 9 13 1 10 9 15
3 7 13 15
5 13 0 13 10 9
13 3 3 13 0 13 10 9 10 9 7 10 9 13
6 15 3 13 7 13 15
2 6 9
12 7 10 9 1 10 9 13 1 10 9 10 9
12 1 0 10 9 13 13 1 10 9 15 10 9
20 7 3 13 1 10 9 11 13 1 11 1 10 9 10 11 1 0 10 9 11
14 7 13 15 0 7 0 7 13 15 16 13 15 10 9
30 7 13 15 1 10 9 1 0 13 10 9 1 10 9 15 7 13 13 10 9 15 7 13 1 10 9 13 7 13 15
4 8 15 13 13
16 7 13 15 10 9 7 3 13 10 9 10 9 15 7 13 3
6 7 13 15 16 15 13
4 7 3 13 13
11 3 15 13 7 10 0 13 13 7 0 13
15 13 1 10 9 16 3 9 12 13 15 7 3 13 15 13
12 7 16 13 15 0 1 9 15 13 1 10 9
6 7 15 15 1 3 13
7 7 13 15 10 9 15 16
9 3 0 13 15 3 13 9 1 9
3 15 13 9
3 15 3 13
1 12
14 7 13 10 12 9 13 13 7 13 10 9 15 16 13
4 7 13 10 9
4 7 13 9 0
4 7 13 15 13
4 13 3 3 12
3 7 13 15
15 7 3 13 1 10 9 1 10 9 15 13 1 10 9 11
17 7 13 10 9 7 13 13 15 13 1 15 9 1 10 9 13 15
6 15 10 9 0 13 9
9 6 13 15 16 13 10 9 0 9
9 7 13 15 3 13 13 1 10 3
4 7 13 15 13
1 13
10 13 1 10 9 10 9 7 10 9 11
5 7 13 1 15 16
3 9 3 13
6 15 13 16 9 3 13
2 3 13
6 3 13 13 10 9 15
26 9 13 3 13 7 9 13 3 13 7 3 13 16 10 12 9 13 1 10 12 7 15 9 9 0 13
2 13 15
1 12
12 16 3 10 12 1 10 12 15 9 9 9 13
2 7 13
3 7 13 15
4 7 13 1 11
10 7 13 15 0 7 13 15 16 15 13
26 7 13 10 9 10 0 13 15 1 10 9 7 13 1 10 9 15 13 10 9 15 13 15 16 15 13
3 7 13 13
8 13 10 9 16 3 9 13 13
17 3 3 13 10 9 1 10 9 15 7 13 7 13 7 13 3 0
7 7 13 15 1 9 15 13
10 7 1 10 9 13 10 9 15 13 15
6 15 15 13 10 9 13
18 15 3 13 15 13 16 11 10 9 7 15 11 15 3 16 12 10 9
4 7 0 13 15
6 15 3 15 15 13 13
5 13 10 11 13 15
4 15 13 10 11
8 7 13 15 16 15 13 1 15
5 7 9 10 9 13
8 7 13 10 11 15 13 13 15
12 15 3 13 7 13 10 9 15 13 11 7 13
14 13 1 15 11 16 3 13 10 10 9 7 10 10 9
10 7 13 10 9 1 10 9 15 13 15
15 15 13 1 15 13 13 15 7 13 10 9 15 7 13 15
10 15 3 3 13 10 9 15 13 13 15
14 15 3 3 13 10 15 9 1 15 7 10 9 13 15
37 15 3 16 13 15 7 10 15 9 1 10 9 0 10 9 7 0 7 10 9 10 9 13 15 3 13 1 10 9 10 9 15 1 10 9 10 0
3 7 13 15
24 6 13 15 16 13 15 3 10 13 15 3 3 13 9 16 3 13 10 9 10 9 13 1 9
45 7 1 9 12 13 10 11 10 11 7 10 11 7 10 11 7 13 15 1 9 0 1 0 0 7 13 1 15 7 10 9 15 13 13 0 3 15 9 1 10 9 3 13 3 13
11 7 13 15 11 1 11 7 13 13 10 11
7 7 13 10 11 13 10 11
18 9 0 13 15 3 13 7 13 12 9 15 12 7 11 12 7 11 12
3 0 3 13
7 0 13 10 9 15 10 0
2 13 15
12 7 3 13 3 15 13 7 10 11 0 1 15
23 7 13 15 1 10 9 13 15 16 15 15 13 13 3 3 3 10 9 10 9 1 0 13
13 7 10 9 13 1 15 13 15 13 10 1 0 13
4 7 13 15 13
4 15 3 13 15
5 11 13 0 13 15
5 16 0 13 7 13
16 7 13 15 16 7 11 13 7 13 15 15 13 3 13 1 15
15 7 13 1 10 9 13 9 0 1 15 7 9 13 1 15
12 7 3 15 10 9 13 15 13 7 13 13 15
3 7 13 15
7 7 13 15 12 1 10 9
24 9 13 10 9 15 1 15 13 9 0 7 3 3 15 13 13 7 13 7 13 10 9 7 13
11 7 13 10 9 15 16 15 13 7 3 13
8 6 9 0 1 3 1 15 13
4 1 3 13 15
4 13 15 1 15
5 7 13 15 1 15
5 7 13 10 9 15
7 15 9 13 3 0 13 15
3 15 3 13
2 1 3
9 7 16 15 13 13 15 13 1 15
8 10 3 11 13 15 10 16 13
4 15 0 10 13
1 13
4 13 15 10 9
15 13 3 10 11 16 13 10 9 13 10 9 10 0 13 15
8 10 0 7 0 9 15 13 15
8 13 1 15 7 3 13 1 15
10 7 13 3 0 16 10 0 13 16 13
11 10 3 11 13 10 9 15 13 15 7 13
6 3 15 3 13 13 15
3 7 13 15
11 0 10 9 1 15 13 13 3 3 1 9
13 7 3 13 13 1 10 11 7 3 13 16 15 13
26 13 3 10 9 15 7 13 15 16 10 9 10 9 13 1 9 9 7 13 15 7 13 1 12 9 13
9 15 3 13 10 9 7 13 15 13
7 7 1 10 9 13 13 15
3 15 3 13
9 1 15 3 13 1 10 9 15 0
8 7 13 13 10 12 7 13 15
11 16 15 13 0 13 13 15 0 7 15 9
13 7 13 9 13 15 1 0 15 7 13 15 13 15
13 15 3 12 10 9 0 13 1 10 9 15 15 13
12 7 15 3 15 13 3 15 13 7 10 13 15
4 10 3 11 13
3 3 13 15
15 15 3 13 15 13 9 1 10 9 15 7 13 0 13 15
9 15 3 3 13 1 15 1 15 13
23 15 3 3 13 15 9 9 1 9 15 16 11 13 6 13 15 16 3 3 13 10 9 15
27 7 15 3 13 12 10 0 0 10 13 0 13 15 3 16 13 9 0 1 10 9 15 7 13 1 10 9
9 7 16 13 15 10 9 15 13 15
22 0 13 15 0 13 1 10 9 3 10 12 9 13 13 1 10 11 1 10 9 10 0
17 0 13 15 13 1 10 9 0 3 10 12 9 13 13 1 10 11
9 7 16 10 9 15 13 15 13 15
29 0 15 13 0 13 1 10 9 10 9 3 12 9 13 13 1 10 11 3 10 9 15 3 13 7 10 9 3 13
4 15 3 9 13
3 0 10 9
10 16 3 10 9 0 13 1 15 15 13
8 13 1 15 9 7 13 1 15
25 7 3 13 13 1 10 9 10 11 7 1 10 11 7 13 3 9 1 15 7 3 13 3 13 15
4 15 15 13 11
3 15 3 13
7 13 11 9 9 13 7 13
5 10 3 11 13 15
9 1 10 9 15 13 15 10 9 0
9 1 3 9 9 0 7 0 13 15
25 1 0 13 9 10 9 15 7 10 9 15 7 13 10 12 1 9 12 16 3 13 12 7 12 9
11 7 1 10 9 3 10 9 1 0 13 15
12 15 3 13 10 9 15 7 13 15 13 1 15
10 7 16 15 13 10 9 15 13 15 13
7 7 13 15 9 16 13 15
6 10 3 9 13 10 13
8 13 3 10 11 13 7 13 15
6 13 10 9 13 1 15
8 10 3 0 13 10 9 10 9
3 6 13 15
9 7 13 15 13 13 10 9 1 15
12 7 13 15 1 9 13 12 7 13 15 13 15
8 9 0 15 13 16 9 0 13
5 10 3 11 13 15
4 15 15 13 0
3 10 9 13
2 3 13
2 3 13
2 3 13
2 3 13
8 13 10 9 15 7 10 9 15
4 15 3 13 15
10 10 3 11 13 15 13 15 7 13 15
3 12 15 13
1 13
16 15 13 13 7 13 10 0 7 13 9 1 9 7 6 13 15
5 13 3 13 9 0
8 7 13 10 11 13 10 9 15
12 3 3 10 10 9 13 1 10 9 10 9 13
7 10 3 11 3 13 13 15
10 9 3 0 13 1 10 9 10 9 13
17 0 13 9 1 10 9 10 9 13 3 0 1 10 9 10 9 13
7 15 3 3 13 13 1 15
4 7 15 13 13
7 1 9 0 7 3 1 9
6 15 3 0 1 10 9
7 6 15 13 15 7 13 15
3 13 10 11
3 6 13 15
53 15 13 15 13 9 7 9 7 9 7 9 7 9 7 9 7 9 1 15 7 1 10 9 16 3 13 0 3 1 10 9 0 9 7 9 7 9 7 9 7 9 7 9 1 9 7 1 10 9 10 13 9 0
9 0 3 13 0 0 7 10 0 0
20 13 3 1 10 9 13 1 11 7 13 13 15 10 11 7 13 10 3 13 13
40 6 13 1 11 7 10 9 10 9 13 10 9 7 10 9 7 13 15 9 7 13 15 10 9 7 13 15 7 13 15 7 13 15 7 13 7 1 12 9 13
9 9 13 16 15 3 13 15 13 15
4 15 3 13 15
5 15 13 15 13 15
4 15 3 13 15
17 13 15 16 12 15 1 0 7 12 15 1 0 13 1 10 9 15
5 10 3 11 13 15
4 3 13 15 13
1 13
5 10 3 11 13 15
13 10 9 15 15 13 13 7 10 9 15 15 13 13
16 10 3 13 1 0 15 3 1 0 3 13 15 13 7 15 13
10 7 13 10 12 13 13 1 11 7 11
7 7 13 15 10 11 13 15
15 13 16 10 13 13 10 9 13 15 7 10 0 15 13 15
6 3 3 3 13 1 15
19 7 3 10 9 10 9 3 13 13 7 13 7 13 10 9 15 9 1 0
4 7 13 1 11
22 7 13 15 1 11 7 10 9 15 7 9 0 10 9 11 11 0 9 13 1 10 9
11 7 13 16 11 10 9 13 13 13 7 13
5 9 11 11 13 15
6 7 13 15 0 16 13
5 15 3 0 3 13
4 9 11 13 15
6 7 13 10 0 13 15
1 13
1 13
2 13 15
11 15 3 13 10 9 15 13 13 1 10 11
6 7 13 15 10 11 13
4 15 15 13 13
3 9 16 13
1 13
5 10 9 15 13 15
9 7 3 13 7 13 15 1 10 9
21 7 16 13 1 11 7 1 11 1 10 9 10 9 13 12 10 9 15 7 13 15
21 13 1 10 9 10 1 15 7 3 13 1 15 13 9 13 1 15 15 9 3 13
4 13 15 7 13
11 10 9 15 9 13 7 3 15 13 3 3
17 7 13 7 13 10 9 13 1 10 9 3 1 10 9 7 13 15
5 15 13 13 10 9
8 15 3 13 15 3 13 10 11
3 7 13 15
17 7 13 10 9 1 10 11 7 13 15 10 9 15 7 13 1 15
16 7 0 10 9 15 13 1 10 9 15 3 9 13 1 10 9
7 6 13 10 13 1 9 9
12 13 10 13 9 10 9 15 11 6 1 10 0
7 7 13 1 11 1 10 9
8 7 10 3 13 15 1 11 13
23 7 13 9 1 3 13 9 13 16 3 15 13 1 15 7 13 1 15 15 13 3 3 9
6 10 3 9 3 13 9
4 7 13 13 15
5 7 13 10 9 15
4 7 13 1 11
43 7 13 1 10 9 13 13 10 13 7 10 13 1 10 9 7 10 9 10 9 7 10 9 10 13 10 9 13 7 3 13 16 15 13 9 1 10 9 7 13 7 13 15
12 3 13 16 10 9 15 9 9 13 15 10 9
12 7 13 10 9 7 10 9 7 13 3 15 13
3 13 3 15
9 15 3 10 9 13 1 10 9 15
9 7 13 3 13 10 9 13 1 9
6 7 13 10 11 13 15
2 9 13
5 10 9 15 13 13
6 7 13 10 11 13 15
31 6 13 15 16 15 3 13 10 9 0 13 7 13 1 10 9 7 3 13 1 10 9 15 7 13 16 15 13 13 13 15
4 1 0 13 15
24 7 3 13 13 13 16 15 13 1 15 16 3 10 9 15 10 1 10 9 13 15 10 9 15
5 7 13 3 1 11
20 7 1 10 9 13 15 13 1 15 10 9 7 10 9 7 10 0 7 13 15
5 1 15 9 0 13
10 7 15 15 10 9 0 13 16 0 13
5 10 3 11 13 15
10 10 9 10 11 1 9 13 7 1 9
5 7 13 1 15 13
5 16 13 1 9 13
6 1 15 3 3 13 15
2 7 13
2 1 9
3 13 10 9
9 0 3 13 10 11 3 16 9 13
5 7 10 11 13 15
9 3 15 13 15 1 15 9 0 13
6 7 13 15 1 9 13
18 9 9 13 7 13 9 7 13 9 7 13 9 7 13 15 9 7 13
18 7 13 1 10 9 10 9 9 16 1 10 9 13 1 10 9 10 9
7 7 13 15 13 7 13 0
7 7 3 13 1 15 15 9
5 3 0 13 7 13
12 7 0 13 7 0 15 15 3 13 15 3 13
5 3 12 13 9 0
7 13 15 0 1 15 13 16
4 13 10 9 15
8 0 3 10 9 1 15 13 16
4 0 13 10 9
8 6 13 15 7 15 13 10 9
10 7 13 13 15 7 13 15 1 10 9
5 7 10 9 0 13
10 9 15 13 10 13 0 13 1 9 9
10 1 9 13 0 7 13 0 1 9 15
8 7 13 15 13 7 13 10 9
8 13 3 16 1 15 10 9 13
4 7 13 15 13
14 7 13 1 15 15 10 9 7 10 9 16 15 13 9
11 9 13 16 0 13 7 3 13 15 1 15
6 13 9 9 13 7 3
4 13 7 3 13
8 15 3 13 15 10 9 13 15
3 15 15 13
5 13 15 9 16 13
3 15 3 13
7 15 10 9 0 7 10 9
4 15 3 13 15
5 10 3 11 13 15
10 10 9 13 9 7 10 10 9 10 9
4 7 13 1 15
14 7 13 9 1 15 15 13 9 3 13 7 13 15 13
29 9 11 13 15 16 16 15 9 13 7 13 9 7 3 13 9 3 13 10 9 15 10 9 7 13 9 10 9 15
10 7 10 0 13 9 7 13 3 13 9
10 7 10 0 13 15 7 13 3 13 9
4 7 10 0 3
6 0 15 3 10 9 13
9 1 10 9 3 13 15 15 13 9
6 10 3 12 13 15 9
4 13 15 10 11
16 3 3 1 0 13 7 13 7 13 7 13 3 9 1 10 9
21 1 3 10 0 16 13 3 13 1 10 9 11 1 10 9 3 13 15 10 9 13
12 15 10 9 11 7 10 9 11 7 10 9 11
6 3 13 9 0 7 13
15 7 13 12 10 9 13 15 13 13 16 3 13 15 13 15
5 15 13 9 0 15
6 13 10 11 16 0 13
7 9 10 9 15 9 1 13
29 7 13 9 10 9 15 1 0 10 9 15 7 1 0 10 9 15 7 1 0 10 9 15 7 1 0 10 9 15
2 0 0
6 13 10 3 15 3 15
6 0 0 15 9 3 13
14 3 9 1 9 13 16 12 13 7 3 13 15 1 15
33 7 10 13 15 1 0 10 9 7 1 0 10 9 7 1 0 10 9 7 10 13 10 3 3 15 0 13 15 10 9 7 10 9
8 3 3 13 1 10 9 10 9
6 7 15 3 13 15 13
9 7 13 10 11 13 13 1 10 9
10 3 13 10 9 16 10 11 9 11 13
8 0 11 13 1 10 9 10 0
6 13 10 9 10 9 15
10 0 11 13 15 9 7 3 15 13 9
6 7 1 10 9 15 13
24 13 1 10 9 10 13 1 9 13 7 9 1 10 9 7 9 1 10 9 7 9 1 10 9
14 10 13 10 9 10 9 7 9 0 13 0 13 0 9
14 7 13 1 10 9 13 3 10 9 13 9 1 10 9
16 7 0 0 13 0 7 13 12 9 0 13 9 12 15 13 9
7 7 13 10 9 15 13 15
17 6 13 15 16 10 9 0 10 0 0 15 13 10 13 1 10 9
12 7 13 15 1 10 9 13 15 12 10 9 15
2 9 13
5 15 9 7 15 9
5 7 10 11 13 15
5 13 0 10 0 9
10 3 3 13 9 1 9 15 3 3 13
23 7 13 15 1 10 9 10 9 1 10 9 13 15 1 0 10 11 7 11 7 11 7 11
14 13 15 3 0 13 7 15 10 9 3 13 0 13 15
5 13 3 15 15 13
13 0 13 1 10 9 15 13 16 15 13 7 0 13
9 3 3 13 9 7 9 9 3 13
6 13 13 7 3 10 9
9 13 3 9 1 9 7 9 1 9
4 13 9 1 9
2 13 9
3 9 9 0
10 7 1 15 10 9 0 13 13 10 9
20 7 3 13 15 13 3 13 15 13 7 0 3 13 15 1 0 10 9 0 13
11 3 3 13 15 10 13 7 10 9 10 0
17 7 13 9 9 1 9 7 9 9 7 13 9 1 9 7 13 15
9 7 13 13 1 15 1 10 9 15
7 10 3 13 1 9 0 13
23 3 3 13 10 9 10 9 13 3 3 13 10 13 13 3 10 1 10 11 13 1 10 9
13 6 3 10 1 9 13 7 10 13 1 0 10 9
24 13 3 10 9 0 9 15 3 13 0 1 9 9 15 13 10 9 1 10 3 7 3 3 13
12 7 16 3 13 9 10 9 3 3 13 15 9
9 7 1 10 0 15 13 13 10 9
14 7 3 16 15 15 13 13 3 10 11 13 3 3 13
17 13 3 9 7 9 7 13 9 7 9 1 10 13 16 0 10 0
3 15 3 13
36 7 1 0 10 9 1 10 9 0 10 9 13 7 10 9 3 13 10 9 15 7 10 9 13 1 10 9 13 7 10 9 10 1 10 9 13
15 7 3 13 10 9 10 9 13 1 9 1 9 0 7 9
7 1 3 10 9 13 10 9
17 3 15 3 10 9 0 13 7 13 10 9 13 16 3 10 9 13
13 3 3 15 3 13 0 13 13 16 3 13 1 9
15 6 13 15 16 3 3 13 10 9 0 16 15 0 15 13
6 10 9 7 10 9 13
22 1 3 10 9 0 7 10 9 15 13 7 10 9 1 9 7 10 9 3 3 10 9
1 13
1 13
24 3 9 0 13 10 9 15 7 13 10 9 15 10 9 15 10 9 15 7 10 9 13 16 13
2 13 3
17 3 13 3 3 10 9 10 9 13 7 3 7 9 7 9 7 3
6 3 13 3 13 15 13
23 13 3 10 9 7 10 0 1 12 9 7 13 10 9 7 10 9 3 15 1 9 13 13
2 13 3
4 3 1 10 9
5 3 13 9 10 9
7 13 10 9 13 15 10 9
6 13 3 15 13 1 15
8 1 15 10 9 0 10 9 13
3 7 13 15
4 10 3 11 13
2 13 15
4 15 15 9 13
5 0 9 13 1 15
5 15 3 3 3 13
3 15 13 13
21 6 3 13 15 3 3 13 10 9 1 0 10 9 7 15 13 0 13 1 9 15
15 7 11 11 10 12 10 12 13 1 10 9 16 15 13 15
9 15 3 13 13 7 13 15 9 13
6 7 13 3 15 3 13
15 7 10 0 9 10 0 16 10 9 13 13 15 10 9 15
8 3 13 13 13 16 13 10 9
11 13 1 10 9 7 13 15 9 9 9 13
13 3 13 10 9 15 3 10 9 1 10 9 15 13
12 7 15 15 13 9 0 13 0 7 3 13 15
18 7 13 10 9 7 13 1 10 9 7 13 3 13 15 7 13 10 9
7 7 0 13 13 1 10 12
8 7 13 15 7 13 10 11 13
13 6 13 15 16 12 1 15 13 15 10 13 1 15
8 13 13 7 13 15 12 1 12
10 12 10 12 10 13 1 15 1 10 9
11 3 10 3 9 10 9 13 3 13 1 15
12 6 3 10 9 0 1 15 10 9 10 9 13
8 0 15 16 3 13 10 9 0
12 7 13 15 13 9 13 13 7 13 15 7 13
1 13
5 0 13 10 9 15
11 7 13 9 13 13 15 7 13 1 15 15
11 0 13 10 9 15 10 9 10 13 1 0
26 6 13 15 16 3 3 3 13 1 10 9 10 9 1 10 9 0 3 15 13 0 1 10 9 10 9
8 7 13 13 1 10 9 10 9
6 7 13 15 10 11 16
4 15 13 16 13
7 13 10 9 7 10 9 13
10 7 1 10 13 15 13 15 1 10 11
5 10 3 11 13 15
17 6 13 15 16 15 3 0 10 9 16 3 3 9 13 3 15 13
4 15 3 3 13
9 16 15 13 13 15 3 3 15 13
5 3 3 7 15 13
13 7 13 1 9 15 10 9 11 7 13 10 9 15
4 13 3 16 13
18 7 13 10 11 7 11 7 11 1 15 7 13 13 7 13 7 13 15
4 13 3 7 13
6 9 10 9 15 0 15
6 13 10 9 0 1 15
8 7 3 15 15 13 7 15 15
10 7 13 7 13 15 13 7 13 10 11
2 11 13
5 3 13 12 9 13
8 10 3 9 0 10 3 9 0
8 7 3 13 13 10 15 9 13
12 13 3 15 10 9 13 7 3 13 15 13 15
7 7 13 10 0 7 13 15
5 13 10 0 7 13
1 13
3 13 10 9
1 13
1 13
5 6 10 13 15 13
8 13 3 10 13 15 9 15 13
5 15 3 13 0 13
5 13 15 7 13 3
10 7 13 3 13 15 13 9 7 13 15
18 12 3 15 10 13 13 10 9 13 10 9 10 9 7 13 15 10 9
6 7 13 10 11 13 15
10 3 1 9 13 1 9 7 9 13 15
13 1 9 13 1 15 1 10 9 13 7 3 13 15
5 7 13 15 13 15
13 7 12 15 9 13 15 13 9 1 0 7 13 15
7 15 3 13 10 9 0 13
25 7 10 11 1 3 13 15 1 3 1 10 9 10 9 7 13 13 1 10 9 7 13 1 10 9
19 10 3 9 7 0 10 9 13 1 10 11 9 1 10 13 15 7 3 13
11 0 3 13 1 15 7 0 10 9 3 13
8 7 15 13 13 1 15 13 16
5 15 13 15 13 16
8 7 3 3 0 13 10 9 15
10 7 13 10 9 1 0 13 10 11 13
4 15 0 15 13
7 15 3 13 7 3 13 15
8 3 10 9 13 15 7 13 15
8 15 13 10 11 10 9 10 0
4 10 3 11 13
20 15 13 7 13 10 9 10 9 1 0 13 10 9 7 13 1 10 9 10 9
5 15 3 9 13 9
3 15 15 13
8 10 3 15 13 15 0 13 9
16 7 13 15 13 15 7 13 15 10 9 7 13 15 7 13 15
1 13
6 7 10 9 9 15 13
22 7 13 10 11 3 1 10 9 13 12 10 9 10 9 7 13 10 11 13 13 15 13
8 3 15 1 10 9 13 10 11
9 7 13 3 1 10 9 7 9 13
11 7 10 9 13 15 13 3 13 10 13 16
4 0 1 15 13
4 15 3 3 13
9 7 1 0 3 10 13 13 10 11
4 3 1 15 13
4 7 3 0 13
7 15 3 13 13 7 13 16
6 7 3 1 0 9 13
12 7 13 10 11 10 9 3 13 15 10 11 16
7 16 9 13 3 3 15 13
3 7 13 13
24 7 3 3 9 13 10 9 1 10 0 7 10 9 7 0 10 9 13 10 11 13 7 13 11
5 7 13 15 10 11
6 15 13 10 9 10 0
5 15 3 13 15 13
6 10 3 11 3 13 15
3 3 13 15
4 13 15 15 13
10 10 3 11 3 15 13 16 13 10 11
9 1 3 9 13 15 12 9 15 13
15 13 3 10 13 11 1 10 9 13 15 1 10 9 9 13
9 7 13 10 9 13 13 3 13 15
7 13 13 15 10 9 10 0
12 10 3 9 13 10 9 16 3 10 11 13 15
7 10 3 11 3 13 13 15
10 15 3 13 13 15 13 10 9 10 0
4 15 3 3 13
2 13 15
5 10 3 11 13 15
4 15 3 3 13
2 13 15
16 10 3 9 13 15 3 10 9 15 13 9 7 13 0 10 9
10 7 13 15 9 7 13 15 13 0 9
4 7 13 13 15
4 13 9 10 0
15 7 13 15 10 9 9 7 13 15 7 13 10 9 13 15
5 7 13 15 16 13
19 7 13 13 15 11 0 13 1 9 10 9 11 7 11 16 13 10 9 15
12 7 13 15 1 10 11 9 15 13 13 9 9
4 15 3 3 13
15 7 13 15 7 13 10 9 15 13 9 1 15 15 15 13
7 13 3 9 0 7 13 15
8 7 13 10 9 10 9 15 13
14 7 1 15 13 12 9 12 1 0 7 12 1 0 15
11 7 10 13 13 15 13 10 9 15 7 13
15 6 10 13 10 9 7 13 12 9 13 15 13 1 10 9
11 3 3 10 9 13 1 15 1 10 9 13
4 15 3 13 13
14 10 11 10 9 11 13 3 1 10 9 16 13 7 13
7 7 10 13 1 15 13 15
9 7 10 0 9 13 10 11 9 0
4 8 8 8 8
3 15 13 13
10 10 9 15 10 9 15 1 15 13 15
6 7 15 10 13 13 13
2 11 13
12 13 3 15 7 13 9 9 13 9 13 15 13
6 13 16 13 11 13 15
7 10 3 11 13 9 0 13
12 7 10 9 10 9 13 1 12 1 3 1 3
13 13 3 10 9 10 13 1 0 15 16 3 13 13
7 3 0 10 9 9 13 9
43 13 3 3 9 1 3 13 1 15 7 11 10 9 7 11 10 11 10 0 7 11 9 7 11 15 16 13 1 10 11 13 15 7 13 15 7 15 0 10 13 15 1 11
16 10 3 11 13 16 3 13 7 13 10 9 13 15 16 3 13
26 7 13 9 13 15 13 10 9 7 13 15 1 9 15 13 13 1 9 7 13 9 1 10 9 10 9
12 10 3 11 10 9 7 11 10 11 13 3 13
19 7 13 10 9 11 10 9 7 11 10 11 7 11 13 9 16 13 13 15
14 7 3 3 10 12 10 9 13 1 10 9 13 10 9
4 7 13 1 15
10 15 13 15 10 9 1 10 9 10 9
7 7 13 13 16 13 10 9
4 15 3 13 15
2 3 13
6 11 13 10 9 10 13
1 13
3 3 13 3
1 13
5 10 9 3 13 15
2 7 13
6 3 15 13 3 13 15
6 7 13 13 1 10 9
10 13 3 15 9 7 9 7 15 15 13
2 13 3
15 13 3 3 0 9 13 0 11 10 9 1 15 13 12 9
10 0 13 13 10 1 15 13 13 7 13
10 7 0 13 16 13 7 13 1 15 13
14 1 3 0 12 1 15 13 13 1 0 9 13 1 9
20 0 13 15 10 12 13 7 13 10 9 15 7 9 16 10 13 15 13 3 13
3 7 13 15
11 13 1 10 9 0 13 10 9 15 10 9
5 10 13 7 13 13
4 10 3 13 13
6 9 3 10 13 0 13
6 1 10 9 15 9 13
11 9 13 7 16 0 15 13 3 3 15 13
18 10 3 3 9 1 10 13 15 13 1 10 9 7 13 1 0 10 9
16 0 3 13 13 3 10 9 13 7 10 9 13 1 10 13 9
43 16 0 13 13 9 1 10 13 1 15 9 3 13 15 10 1 9 9 7 9 13 10 9 13 3 15 13 3 15 3 3 15 13 0 11 16 13 1 15 13 9 10 9
27 13 1 10 9 11 9 10 11 9 15 9 11 1 9 11 7 9 15 1 10 9 11 7 10 9 15 11
17 13 3 0 0 1 10 9 13 1 15 10 9 7 9 10 9 0
18 7 3 13 15 9 16 13 10 11 9 7 0 13 1 10 9 15 13
12 13 3 15 9 9 13 1 0 10 9 10 9
4 7 13 11 13
6 13 3 1 15 10 9
22 3 13 11 16 13 10 9 15 7 10 9 15 11 13 9 15 7 13 10 9 15 11
13 7 13 9 15 7 9 7 0 1 10 9 15 13
32 13 3 0 1 9 7 9 7 9 3 3 13 7 9 0 13 3 1 9 9 15 7 0 10 9 11 13 1 9 10 9 15
24 7 15 13 1 15 1 9 7 9 11 13 9 9 1 9 7 0 1 9 0 13 9 9 13
4 1 15 13 0
13 15 3 13 9 7 10 9 15 13 1 10 9 15
6 7 13 10 9 13 15
26 7 6 13 13 7 3 13 13 1 15 9 13 0 16 15 3 13 10 9 15 15 13 1 10 9 15
16 7 13 10 9 13 10 11 7 13 1 10 13 15 1 10 9
14 13 3 3 13 13 15 7 13 16 9 13 1 10 9
8 7 15 13 13 15 7 13 0
10 1 3 0 10 9 13 11 10 9 15
7 7 13 15 9 12 13 16
13 3 15 13 9 1 9 15 13 13 9 15 1 9
36 1 3 10 9 10 0 13 10 9 11 1 10 9 1 9 10 11 15 9 11 1 9 13 9 15 9 11 1 9 11 7 10 9 10 9 11
1 13
5 13 10 9 1 15
13 15 3 1 10 9 13 7 13 15 13 10 9 0
3 3 13 11
6 13 3 9 1 10 9
14 7 6 13 1 9 7 13 9 7 13 10 9 15 11
35 0 13 0 7 9 0 13 7 13 15 9 10 9 10 9 11 10 9 15 7 13 1 10 9 11 1 10 9 7 10 9 15 3 13 9
6 13 3 11 1 10 9
6 7 13 10 9 13 15
10 9 0 13 1 15 7 9 0 13 15
30 7 6 11 10 9 15 3 15 13 9 1 9 15 7 0 9 0 13 15 10 13 9 16 3 13 1 10 9 15 9
3 13 3 11
4 6 10 9 9
6 13 15 1 10 9 15
6 7 13 1 15 10 9
26 13 3 11 1 10 9 0 13 1 10 0 1 9 1 9 11 7 13 1 10 9 11 7 13 10 11
12 7 13 9 0 10 11 7 13 9 0 7 13
13 7 3 15 0 16 13 10 9 10 9 15 1 15
22 6 3 16 13 10 9 10 9 15 1 10 9 15 13 1 9 10 9 1 10 9 15
12 7 0 10 13 16 13 9 10 13 15 1 9
3 7 13 11
25 13 10 9 15 10 9 7 13 10 9 15 1 10 9 10 9 15 16 13 1 10 9 10 9 15
16 6 3 1 10 3 13 15 15 10 9 16 13 15 0 10 0
16 7 0 10 9 15 7 10 9 15 1 9 7 9 10 13 15
7 13 9 1 9 7 13 0
7 13 13 0 7 13 13 0
21 13 11 9 15 13 9 3 13 1 10 9 15 10 11 7 10 9 15 1 10 9
14 13 3 11 1 15 3 9 12 7 13 1 10 9 15
12 10 3 11 13 10 9 10 13 15 7 13 9
19 7 13 10 0 7 10 0 15 16 13 9 10 9 15 1 15 7 13 15
21 7 13 1 10 9 10 0 13 13 10 9 7 13 15 1 10 9 10 9 15 11
6 7 13 10 9 15 13
5 7 13 1 15 16
11 15 13 1 10 9 15 15 13 10 9 0
11 13 3 10 9 15 10 15 3 13 13 15
5 7 13 9 13 13
5 11 13 10 9 15
3 7 13 15
15 13 3 10 9 15 3 7 10 9 15 7 13 13 10 9
30 7 13 1 15 9 10 13 15 7 1 0 10 0 10 11 13 15 10 9 0 7 13 15 10 13 1 10 9 15 13
11 7 11 10 9 15 13 9 0 7 13 13
45 0 9 10 9 10 11 16 13 7 13 9 10 9 15 7 13 9 9 15 1 9 11 9 15 3 13 1 9 10 0 1 9 9 15 9 1 0 15 7 1 9 15 10 13 15
39 13 9 1 10 9 15 7 13 9 0 15 9 15 13 1 11 10 9 15 10 13 15 3 1 9 0 13 13 15 1 9 7 9 1 15 15 10 9 15
7 3 15 3 9 9 0 13
47 13 3 1 9 9 13 9 15 10 13 9 9 10 9 15 1 9 9 15 1 9 9 9 15 1 15 13 15 9 1 9 13 10 1 9 7 9 9 13 10 13 10 9 15 1 9 9
19 10 3 9 13 7 13 9 7 13 1 10 0 1 9 9 15 1 10 11
15 13 3 1 10 9 0 13 9 1 9 11 13 15 10 9
9 7 13 15 13 0 1 10 15 9
36 13 3 1 10 13 15 3 13 10 9 10 13 15 7 13 10 9 15 10 0 7 13 15 7 13 15 1 9 16 3 13 15 9 1 10 9
18 7 9 13 1 10 9 10 15 13 7 13 9 10 9 1 10 9 15
14 7 9 9 13 15 7 9 9 13 15 7 13 9 0
5 7 13 15 10 9
2 3 13
23 6 3 13 15 9 0 15 13 15 10 9 16 13 15 3 9 15 13 11 9 1 9 11
5 13 9 13 1 9
14 7 3 13 1 10 9 9 9 0 13 10 9 7 13
16 7 13 3 13 1 15 1 10 9 10 9 10 9 13 1 15
16 13 3 1 11 7 13 10 9 0 10 13 15 10 9 13 15
18 7 13 13 7 13 10 7 11 7 10 11 7 10 9 13 1 10 9
13 13 3 13 1 10 9 10 13 15 1 10 9 0
13 7 15 10 13 13 1 10 13 1 10 9 1 15
19 7 13 10 9 13 7 13 10 9 1 15 15 13 7 13 3 13 1 15
26 7 16 13 9 12 10 13 15 7 13 10 9 15 11 10 13 1 10 9 1 10 13 15 1 10 9
44 7 16 13 10 9 10 9 15 1 10 9 11 13 15 1 11 13 10 9 3 13 1 9 9 16 15 0 13 9 0 10 9 13 7 10 13 9 1 10 13 1 10 9 9
26 7 6 9 13 1 11 15 9 11 7 10 9 0 0 7 0 13 9 10 11 7 9 13 0 1 15
19 7 13 15 13 1 10 9 10 0 3 13 9 16 3 3 13 10 11 9
8 7 13 1 10 9 1 10 9
32 7 1 10 13 10 9 10 9 11 10 13 15 1 10 13 10 9 1 15 7 15 13 15 1 10 9 7 13 10 9 7 13
15 7 13 10 9 15 7 10 9 15 13 1 10 13 1 15
11 7 13 15 11 7 13 1 11 10 9 15
15 6 0 13 1 9 7 9 0 1 10 11 7 1 9 13
15 3 15 3 15 10 9 13 9 16 3 13 1 0 9 9
32 0 13 1 9 0 13 1 9 9 12 1 10 9 15 7 15 9 1 9 12 15 3 13 10 9 9 7 9 13 9 7 9
17 7 15 10 9 13 13 10 9 7 13 1 15 15 10 13 9 11
16 7 16 13 15 1 10 9 9 13 1 10 11 1 9 15 11
13 7 13 10 9 15 1 9 1 11 10 9 10 9
32 7 16 13 9 12 13 15 1 10 9 10 9 7 13 10 9 1 10 13 15 13 11 10 9 1 11 7 3 13 10 9 15
27 13 3 15 13 1 10 9 13 9 9 7 13 15 1 10 0 7 10 0 7 3 13 13 1 11 13 15
21 7 13 1 9 12 13 15 1 10 9 13 1 0 10 9 7 13 15 7 13 15
13 13 3 15 10 13 15 1 10 9 7 10 9 15
5 9 15 13 15 3
9 6 10 9 15 7 15 13 13 15
4 15 16 13 15
11 3 13 16 1 10 10 9 15 13 13 15
9 7 15 3 13 10 9 15 13 15
12 7 13 1 15 7 13 1 11 7 13 13 15
12 7 10 9 15 13 15 10 9 1 10 9 15
14 7 11 13 1 10 9 7 9 7 9 1 9 7 9
22 7 13 1 15 10 9 10 11 13 9 9 1 9 9 3 13 1 9 9 11 10 9
4 13 10 9 9
5 0 13 10 9 15
21 15 9 13 7 15 9 7 9 13 7 13 10 0 1 0 7 10 0 1 9 0
8 7 13 15 9 10 9 10 9
8 13 3 10 13 9 13 1 15
10 9 9 15 13 15 13 1 10 13 9
6 13 3 9 0 10 9
15 13 3 15 16 13 10 9 1 10 9 0 13 9 10 11
11 3 3 7 10 9 1 10 9 10 9 13
12 15 3 9 3 13 9 0 13 7 1 9 13
6 7 13 15 10 9 13
3 15 3 13
4 13 3 13 15
14 10 13 12 9 13 10 3 13 7 10 13 9 3 13
9 13 3 3 9 13 7 13 1 15
5 15 3 13 1 15
7 15 0 1 10 13 15 13
6 13 3 15 3 13 13
4 15 13 3 15
4 7 13 1 15
9 15 13 15 13 7 13 10 9 15
24 13 3 10 9 7 13 15 1 10 9 15 1 10 11 16 15 13 10 11 13 13 15 10 11
5 15 3 9 13 15
19 15 10 9 1 10 9 15 13 10 9 15 7 13 10 9 1 10 9 15
6 10 3 9 13 9 0
9 0 3 3 3 0 13 13 10 9
33 10 3 11 10 9 13 1 15 1 11 10 9 10 9 15 7 1 15 15 13 0 10 11 13 3 0 1 15 13 10 11 1 9
33 13 3 1 10 13 0 10 9 3 11 13 7 13 13 10 9 7 13 10 9 10 0 0 9 3 9 1 15 7 9 1 9 13
7 15 13 10 9 15 10 0
3 1 15 13
23 11 3 0 9 0 13 1 10 11 7 13 1 10 9 1 10 9 9 12 13 1 10 9
5 13 3 15 10 9
12 16 9 13 10 9 13 10 9 0 16 13 9
6 7 13 1 15 10 11
9 13 16 3 1 9 0 13 10 9
13 7 13 15 13 15 15 10 9 10 9 1 9 9
5 7 13 15 10 9
9 15 3 16 13 1 15 13 15 15
6 7 13 10 11 13 15
9 13 9 10 9 15 7 15 0 13
15 13 3 15 1 11 7 13 1 10 9 10 9 7 13 15
9 16 9 13 10 9 13 15 3 3
25 13 3 16 10 9 15 13 1 15 10 13 15 7 16 1 9 13 15 16 13 1 9 10 9 15
8 7 13 13 15 10 11 16 13
11 7 13 15 9 10 9 13 1 15 1 9
12 7 13 10 11 1 10 9 10 9 1 10 11
9 7 9 13 1 0 10 9 1 15
24 7 13 1 11 3 13 13 7 13 1 10 13 15 1 10 9 10 9 1 10 9 7 13 13
16 7 13 15 9 10 9 11 7 13 10 9 13 9 3 13 13
10 9 9 1 15 15 1 13 15 13 0
16 13 15 13 0 9 7 0 9 13 13 1 9 13 9 9 0
6 13 3 13 1 15 16
9 3 13 10 9 0 1 10 13 15
19 7 15 13 15 7 13 1 10 9 10 9 10 13 1 10 9 15 7 13
5 3 9 13 11 0
6 3 13 15 10 9 0
3 9 13 15
13 15 13 13 1 10 11 13 3 3 1 10 9 15
12 6 13 15 16 15 9 0 13 1 10 9 15
49 1 9 3 13 15 16 0 9 13 1 10 9 11 1 10 11 16 13 10 9 1 9 12 7 9 12 16 13 9 0 1 15 10 9 7 1 15 15 13 11 3 3 1 11 10 11 1 9 9
20 7 0 0 13 1 10 11 1 11 10 9 7 15 15 13 3 3 11 10 9
32 7 13 15 9 1 10 9 13 0 7 13 13 15 1 10 9 7 13 15 1 9 10 9 1 15 10 9 13 15 16 13 15
7 15 3 13 1 0 15 13
13 7 13 1 10 9 15 16 1 9 13 10 9 15
14 7 1 10 9 13 9 13 9 9 0 7 13 9 0
3 13 13 15
4 13 15 15 13
4 10 0 10 9
6 7 13 15 10 11 13
5 13 7 13 1 15
14 7 13 15 10 9 1 10 0 13 1 15 15 13 15
15 15 10 9 0 16 1 9 7 9 13 10 0 9 7 13
10 13 3 1 10 9 13 1 10 9 11
13 9 3 10 11 13 13 9 0 7 13 15 1 15
10 7 13 1 15 13 10 9 7 13 15
5 3 3 13 13 15
14 13 3 10 9 15 15 13 13 9 0 13 15 1 15
10 15 3 12 0 15 10 9 13 13 15
10 13 3 3 9 1 0 13 7 13 16
13 13 3 9 13 13 1 0 9 7 10 9 13 15
12 7 13 1 15 7 13 15 10 3 13 1 15
6 15 3 13 1 15 16
15 3 10 0 9 13 15 13 10 9 10 9 16 1 0 13
8 7 13 13 1 10 9 10 11
30 13 3 1 10 10 9 13 15 7 13 10 9 10 9 7 15 13 13 1 10 9 11 7 13 12 9 13 1 10 9
9 10 3 9 1 15 13 13 10 9
16 13 3 1 12 10 9 15 13 11 13 15 1 10 9 13 0
8 16 3 13 13 13 1 10 11
11 13 1 10 9 7 13 10 9 15 1 9
4 7 13 11 13
7 9 1 0 9 13 15 13
8 1 3 10 9 15 13 10 9
7 7 0 13 13 9 9 0
5 13 3 10 9 15
12 7 13 10 0 1 10 0 9 10 13 13 15
8 13 1 15 16 9 0 13 9
29 9 3 13 15 7 15 10 1 15 1 10 9 10 9 15 13 3 3 7 11 7 11 9 11 15 13 9 10 11
7 7 13 1 10 11 10 11
2 3 13
6 1 10 3 9 13 13
11 7 13 10 9 1 10 9 13 15 13 15
15 7 13 1 10 13 15 1 12 10 9 7 6 9 0 9
6 9 16 13 13 15 13
1 13
1 13
7 7 3 10 9 13 1 15
6 7 15 13 15 15 13
18 7 13 13 15 10 9 7 13 1 10 9 15 3 13 11 1 9 15
18 13 3 3 10 9 1 15 7 13 9 0 13 7 13 1 10 9 15
28 7 13 1 12 10 9 7 15 13 13 7 13 13 9 7 9 15 13 13 1 15 9 10 11 7 11 7 11
8 7 9 9 13 1 10 13 15
27 7 3 13 15 13 15 1 10 9 13 1 10 9 1 10 9 13 15 1 10 9 1 10 0 1 10 11
6 7 13 10 9 15 13
6 9 13 15 10 9 15
9 7 13 13 10 9 7 10 9 13
6 15 13 0 15 13 9
11 13 3 10 11 10 9 15 13 13 1 15
6 15 13 1 10 9 15
14 15 13 0 13 13 15 10 9 15 3 13 13 7 13
3 13 10 13
2 15 13
11 13 7 13 10 9 15 13 1 10 9 15
17 7 3 13 1 15 13 1 15 13 13 1 10 9 15 13 10 9
3 13 0 3
16 7 1 0 13 7 13 9 9 11 13 1 10 9 7 13 15
2 13 15
6 7 13 15 13 13 15
12 7 13 9 0 9 7 0 15 13 1 15 13
13 7 13 10 9 7 10 9 15 1 10 9 15 13
10 1 15 1 10 9 7 0 13 7 13
10 3 9 13 10 13 9 7 10 3 13
8 3 13 13 0 7 0 1 9
5 15 3 13 1 15
19 10 9 11 13 0 7 9 13 3 3 10 10 9 10 3 15 13 7 13
6 10 3 11 13 1 15
16 13 3 9 7 3 13 1 15 10 9 3 13 1 0 10 9
7 13 3 3 9 1 15 16
18 16 3 3 7 10 0 13 7 10 0 3 13 10 9 10 1 10 0
8 7 15 13 9 0 1 9 0
17 16 3 3 13 10 9 10 0 10 9 7 0 13 7 10 9 13
7 7 9 0 1 9 0 13
6 7 15 13 0 13 0
2 13 3
21 13 3 1 9 0 13 15 1 0 7 13 10 9 15 10 9 7 13 13 10 9
8 15 13 15 3 13 13 10 9
7 7 13 10 11 1 15 13
14 3 0 13 15 13 11 16 13 15 7 10 1 15 13
30 3 13 1 10 9 10 9 7 10 9 10 9 13 7 13 7 13 3 10 1 15 15 3 13 13 3 3 0 10 9
13 7 13 15 16 9 13 10 9 10 9 3 10 9
12 13 3 1 0 9 13 15 1 10 9 7 13
12 7 13 9 3 7 10 9 15 10 0 13 0
9 13 3 10 9 10 0 13 10 9
6 13 7 13 1 10 0
3 7 13 13
6 13 3 10 11 1 15
13 13 15 16 13 10 9 13 7 13 9 13 7 13
6 7 13 15 15 13 15
4 13 10 9 15
8 15 3 13 7 13 10 9 15
20 13 3 1 10 9 0 13 15 1 10 9 13 7 13 13 1 10 9 10 9
56 7 16 13 9 13 10 9 15 7 13 1 15 12 15 3 9 13 11 15 7 13 11 7 11 10 9 15 7 11 7 11 7 11 7 11 7 11 7 11 7 11 11 7 11 10 13 9 7 11 11 7 11 11 15 13 9
47 7 13 1 15 13 1 9 0 7 9 0 9 15 7 9 0 10 9 1 15 10 11 7 11 7 10 0 11 7 11 15 13 13 15 7 13 1 10 9 15 7 10 13 1 9 0 13
15 7 15 10 9 13 13 15 16 9 1 15 13 7 13 15
11 7 15 13 10 9 15 1 10 9 15 13
10 0 10 0 16 15 13 10 9 10 9
6 0 10 13 3 16 13
6 0 10 13 3 16 13
9 6 3 10 9 15 0 1 10 9
10 1 10 15 3 13 10 9 10 9 15
10 3 6 15 10 0 16 13 10 9 15
7 6 15 10 13 3 16 13
8 6 10 13 3 16 13 7 13
8 6 3 3 13 15 15 10 9
10 1 10 15 3 13 10 9 10 9 15
4 13 10 0 15
4 13 10 13 15
5 13 1 10 13 15
22 10 13 15 1 10 9 13 3 10 0 7 1 10 13 15 10 9 3 10 9 3 13
12 15 13 15 13 7 1 10 13 10 15 3 13
13 7 3 13 16 13 15 10 9 3 15 13 15 3
10 7 16 13 10 13 15 15 15 9 13
11 7 3 16 13 10 13 15 15 15 9 13
6 3 10 0 10 15 13
8 3 0 0 13 16 13 10 0
11 3 13 10 0 15 7 13 7 13 15 13
19 7 13 10 9 15 0 7 13 9 0 16 15 0 13 1 10 0 7 0
8 13 0 3 10 9 15 0 13
7 7 3 13 7 3 3 13
3 13 7 13
4 13 7 13 15
10 9 0 13 13 13 13 1 10 9 15
5 13 3 3 9 15
5 3 13 0 0 13
5 3 0 1 9 13
6 3 13 9 1 10 9
12 15 3 13 10 9 10 1 10 9 10 9 15
10 10 3 9 10 1 10 0 9 3 13
25 3 13 13 10 9 15 9 13 13 10 9 10 1 10 9 15 0 10 1 10 9 15 9 3 13
22 9 13 0 10 9 1 10 9 15 7 3 13 10 9 10 1 10 9 10 9 15 13
8 0 3 9 1 10 0 9 13
11 3 3 1 9 13 9 7 1 9 9 13
21 10 0 9 1 10 0 9 10 9 13 10 0 7 10 0 1 10 0 13 10 0
11 15 3 15 13 9 9 7 3 13 15 13
18 15 10 13 1 15 7 13 15 10 9 7 13 15 13 15 15 13 0
15 0 13 9 13 9 15 13 7 13 7 13 9 1 10 9
19 9 3 13 13 10 9 10 9 0 7 3 13 13 15 1 10 3 13 15
20 10 3 13 7 3 13 0 13 9 13 9 1 10 9 1 9 15 13 10 9
8 7 13 10 9 10 9 0 0
14 16 13 15 10 9 15 1 10 9 10 9 13 1 11
19 13 3 1 10 11 13 1 15 0 10 0 13 15 16 13 13 10 9 15
16 15 3 13 1 10 11 13 15 3 13 16 0 13 15 13 0
11 13 3 10 9 15 7 10 9 15 13 15
6 10 3 11 13 1 15
13 3 3 15 3 3 13 10 9 13 9 10 9 13
3 9 3 13
7 3 7 15 13 1 15 13
12 3 3 15 9 13 1 9 13 13 1 15 9
6 7 13 0 13 7 13
5 7 0 13 7 13
8 7 10 9 15 13 0 7 13
14 13 3 0 10 11 13 15 7 13 10 13 15 9 13
2 13 15
7 3 1 10 11 0 9 13
28 16 3 13 10 9 10 9 7 6 13 13 0 9 10 9 15 7 15 13 9 7 9 10 9 0 13 1 15
11 7 13 15 10 9 13 1 15 7 13 15
2 3 13
5 7 13 13 10 9
6 10 3 13 13 7 13
3 9 15 13
1 13
13 7 13 10 0 7 13 13 7 13 15 10 9 15
15 7 13 10 9 0 1 0 10 11 1 15 7 15 10 9
9 7 13 11 10 9 15 1 15 0
14 7 13 12 15 10 9 15 10 11 13 1 10 9 13
7 15 13 10 13 7 0 13
7 13 3 1 15 10 9 13
8 11 10 9 13 15 1 15 13
7 15 13 10 13 7 0 13
18 1 0 10 9 13 0 1 9 7 9 7 9 0 7 0 0 13 13
9 7 0 13 15 3 3 13 1 15
12 13 3 10 9 11 13 13 1 10 9 1 11
6 15 13 1 10 0 13
4 9 1 9 13
4 7 15 13 13
5 9 1 0 9 13
12 6 10 1 9 0 7 9 13 1 10 0 13
1 9
3 3 0 9
5 0 13 1 15 13
15 6 13 10 9 15 1 9 15 15 13 10 9 15 1 15
2 13 15
8 0 1 0 9 9 11 15 13
11 10 3 0 1 10 9 10 9 0 15 13
17 10 3 9 7 10 0 10 9 10 9 13 1 15 3 13 1 15
12 15 3 13 10 9 10 9 0 7 15 13 0
5 13 15 7 3 13
4 13 7 3 13
13 13 3 11 10 9 3 13 9 7 13 9 7 13
2 9 13
10 13 10 9 10 9 13 7 13 7 13
9 7 13 10 9 1 10 9 15 15
10 13 3 15 15 10 9 16 13 1 15
8 7 13 1 10 9 10 9 13
11 13 3 10 9 10 13 15 13 1 15 13
17 0 16 13 9 13 3 15 7 15 10 9 15 13 15 16 0 13
7 7 13 10 11 13 1 15
5 11 13 15 15 13
5 12 9 13 9 15
9 10 12 13 9 12 10 3 0 12
6 3 13 15 13 0 13
6 15 3 15 0 13 15
6 13 16 15 10 0 13
4 15 3 13 15
2 3 13
4 13 0 10 9
5 13 15 1 10 9
7 9 15 1 10 9 3 13
13 0 3 10 9 13 15 10 9 7 10 9 15 13
4 9 15 3 13
6 9 10 9 15 3 13
7 0 3 9 13 15 10 9
9 13 15 10 9 10 0 16 13 0
6 15 3 0 13 0 13
3 13 3 15
4 13 15 10 9
7 7 13 10 13 13 1 15
7 15 0 13 15 3 9 13
5 10 9 15 13 15
5 7 13 1 10 3
57 7 15 13 1 9 7 9 13 7 13 10 9 10 9 7 10 12 1 15 7 9 15 15 13 13 1 9 0 7 9 11 10 13 9 1 15 9 12 13 7 11 9 11 9 11 7 11 7 0 0 15 13 15 1 10 13 15
14 13 3 9 0 7 10 1 9 13 1 15 13 1 9
8 13 10 13 10 13 10 9 15
20 7 1 10 13 15 15 3 13 1 10 9 7 13 7 10 9 10 9 13 15
14 7 0 13 1 10 9 7 13 13 1 10 3 13 9
13 7 0 13 1 0 10 9 7 13 10 9 13 15
5 10 13 9 13 13
11 13 3 15 10 9 15 15 0 13 10 9
3 15 3 13
22 15 13 13 10 9 10 9 10 9 10 3 0 1 9 16 13 3 13 7 13 3 13
5 13 3 0 10 9
7 10 9 13 10 9 10 9
8 10 3 1 10 9 13 10 13
16 3 13 10 9 7 13 10 9 1 10 9 15 16 3 13 13
14 7 0 9 3 13 15 1 9 13 7 1 9 9 13
24 10 3 1 10 9 13 0 13 10 13 7 1 9 7 9 7 9 10 9 13 13 7 3 13
22 10 3 1 10 0 9 0 13 15 1 9 0 7 0 13 10 9 13 7 13 1 9
21 15 3 9 13 13 15 9 7 1 9 13 7 1 9 13 16 10 13 13 10 9
18 3 3 13 0 15 3 0 13 7 0 15 3 3 13 7 1 0 13
4 13 3 3 13
18 15 3 3 13 13 15 7 15 3 3 13 3 15 13 13 13 1 15
19 13 3 1 15 10 9 15 7 10 9 15 7 3 13 13 15 1 10 9
6 15 3 13 13 1 15
15 9 15 7 9 15 0 13 10 10 9 10 9 13 7 13
6 13 3 1 12 10 9
13 7 15 13 1 9 7 10 9 15 7 13 1 15
6 13 1 10 3 10 9
2 7 13
4 13 3 15 13
5 13 3 13 15 13
11 15 3 13 13 10 9 7 10 9 10 9
5 7 13 7 13 9
3 13 3 15
4 3 10 9 15
6 13 3 13 13 1 15
15 15 3 0 13 16 7 10 9 13 7 10 9 7 13 15
29 13 3 15 1 10 9 13 9 15 1 10 9 13 9 7 9 0 3 13 9 7 1 9 3 13 7 1 10 9
11 13 3 10 11 13 13 15 7 9 0 13
2 13 15
3 3 15 13
10 13 3 10 9 10 0 13 1 10 9
22 0 3 9 13 15 7 13 9 7 9 13 7 13 10 9 13 1 10 9 1 10 0
6 13 3 15 10 11 13
10 15 3 13 9 16 13 9 0 1 15
11 7 13 15 16 3 13 15 1 10 9 13
19 13 3 3 9 9 0 13 1 10 9 7 13 15 16 13 15 1 0 13
23 13 3 10 9 1 10 9 13 1 10 9 7 13 10 9 1 10 9 1 10 9 7 13
16 13 3 10 13 10 13 13 7 13 1 10 9 7 1 10 9
30 13 3 13 10 13 7 13 1 10 11 7 13 13 10 9 1 15 10 9 13 13 7 13 1 10 9 10 11 7 13
9 13 3 15 10 13 3 13 10 13
6 15 3 13 1 9 13
13 13 3 15 10 9 1 15 13 10 9 13 1 15
4 13 3 15 13
12 13 1 10 9 15 7 13 15 15 13 10 9
11 13 3 1 10 13 10 11 13 15 10 9
5 13 3 15 13 15
13 7 6 13 9 15 9 11 7 15 9 10 9 13
9 1 3 10 13 15 10 9 13 15
36 7 9 13 1 9 9 1 9 12 15 9 13 0 10 9 3 13 1 15 13 13 1 13 10 9 10 9 15 7 3 13 10 9 10 9 15
4 7 13 10 11
4 15 10 13 15
10 13 3 15 13 10 11 7 10 1 15
4 10 3 11 13
3 13 15 15
26 13 3 10 9 16 3 13 13 13 7 13 15 1 15 9 13 15 13 1 15 10 9 7 3 13 3
4 15 3 13 15
6 9 10 9 15 13 15
3 13 1 9
10 3 15 13 13 15 1 10 9 13 16
4 13 10 9 15
6 10 3 11 13 13 15
4 0 13 7 13
26 13 3 1 10 9 3 13 13 15 1 15 3 3 11 7 11 7 11 7 10 9 10 9 7 10 9
6 13 3 15 7 13 15
3 15 3 13
2 3 13
4 3 13 7 13
6 7 13 15 13 16 13
13 7 13 10 9 15 7 13 3 7 13 15 13 13
5 7 13 10 9 15
8 15 3 13 15 15 13 10 13
30 13 3 10 12 13 15 9 7 9 1 15 10 9 7 9 13 7 13 15 13 10 9 10 9 7 13 7 13 1 15
13 15 13 1 10 9 7 9 7 9 7 9 7 9
5 7 1 12 9 13
11 7 1 15 3 9 13 3 13 7 3 13
23 7 15 3 3 13 15 13 1 10 9 0 3 10 9 1 10 9 15 13 1 9 1 15
34 13 3 11 10 9 10 13 15 7 13 1 10 13 1 15 16 11 13 1 0 1 15 3 16 11 13 0 3 16 9 15 10 0 13
3 13 3 11
3 11 15 13
8 15 3 13 0 1 15 13 0
4 7 13 13 15
8 7 13 10 9 13 15 15 13
10 7 13 15 13 1 0 1 9 13 11
22 10 3 9 13 13 15 7 13 15 13 15 1 10 9 10 9 7 10 9 13 9 13
21 13 10 9 16 13 1 10 3 9 7 9 13 7 13 9 16 3 1 0 9 13
4 13 3 1 15
4 13 15 13 15
3 15 3 13
21 3 13 15 0 3 9 12 7 9 12 16 3 13 15 13 1 15 10 9 0 9
5 13 3 3 9 12
6 13 3 1 10 9 15
6 7 13 3 7 13 0
13 7 13 7 13 15 7 13 10 13 15 9 9 12
17 7 13 1 10 13 15 13 1 0 13 15 10 9 7 13 15 13
6 15 15 10 9 13 13
4 15 3 13 13
14 11 10 9 15 3 11 15 3 16 9 15 10 0 13
3 13 3 15
4 11 3 13 13
4 10 11 10 9
4 13 3 1 15
18 16 15 13 1 15 13 13 15 7 13 10 9 15 1 9 7 13 15
10 15 3 3 13 10 9 15 13 13 15
12 15 3 3 13 10 9 15 1 15 0 13 15
13 15 3 13 9 13 10 9 0 15 3 13 7 13
4 13 3 15 3
17 13 15 10 3 13 15 3 3 13 9 16 3 13 10 9 10 9
9 13 3 1 10 9 0 3 9 12
18 7 13 1 10 13 15 10 9 10 9 15 0 7 10 9 15 0 13
24 7 6 9 12 13 15 15 13 11 7 11 15 13 1 9 13 10 9 15 15 13 13 1 11
10 10 3 11 7 10 1 15 13 13 9
13 13 3 13 10 9 15 7 10 12 9 10 13 15
9 0 3 15 13 13 9 7 13 15
9 13 3 1 10 13 15 1 10 9
7 7 9 13 1 10 9 13
7 0 13 10 9 15 10 13
9 7 1 10 13 10 9 13 11 0
13 7 15 13 7 15 13 1 0 10 9 15 15 13
14 13 3 10 3 9 13 15 1 10 9 13 15 9 0
12 9 13 15 13 1 10 9 15 16 0 15 13
20 7 6 9 13 15 7 3 13 7 13 15 1 9 7 3 13 1 15 13 15
11 7 13 10 9 15 16 13 15 7 3 13
5 13 3 10 11 13
13 6 9 0 7 13 1 3 13 1 15 7 13 15
10 3 3 13 15 13 15 10 9 7 13
18 13 3 10 11 10 9 10 0 7 13 10 9 7 13 15 10 9 15
12 15 3 13 1 15 15 13 13 1 10 9 15
9 13 15 1 10 9 15 10 9 0
10 10 3 9 10 9 13 13 1 9 9
23 15 3 13 10 9 0 7 13 13 1 15 16 3 13 15 7 13 13 15 1 10 9 0
11 13 3 9 1 15 10 15 3 13 0 15
18 10 3 11 13 10 9 10 9 15 13 9 13 15 1 15 7 13 15
9 7 15 3 15 13 13 10 13 15
5 13 3 10 11 13
17 9 13 15 1 10 9 15 13 9 7 13 15 16 3 13 1 15
5 13 3 1 15 11
2 3 13
9 15 3 3 13 1 15 1 15 13
26 13 3 1 10 13 10 9 10 9 15 7 15 10 9 15 13 10 13 1 11 7 13 9 1 9 15
9 7 13 13 1 9 9 16 13 15
11 9 13 13 9 13 1 10 9 7 13 15
4 13 3 13 15
5 7 13 1 0 9
10 7 13 15 1 10 9 13 15 1 15
5 13 15 3 3 13
5 7 13 15 10 11
10 10 9 9 13 7 10 9 10 9 9
11 10 3 9 10 9 3 13 3 10 9 13
2 13 15
3 15 3 13
8 13 15 0 13 13 10 9 15
3 13 3 15
7 13 10 0 13 10 15 0
8 15 3 13 13 10 9 10 9
4 13 3 7 0
3 13 15 9
18 15 13 10 9 15 1 9 7 13 1 10 3 0 13 10 9 10 9
26 1 3 0 13 10 9 3 0 12 7 13 15 1 12 1 9 15 1 15 9 7 9 3 13 0 13
4 13 3 1 15
4 10 3 9 0
4 10 3 9 0
13 13 3 10 9 10 9 16 9 13 1 10 9 15
1 13
7 3 13 9 3 9 3 9
8 1 15 3 3 13 9 0 13
4 9 10 9 0
12 7 16 13 3 9 9 13 1 15 10 9 15
6 16 3 3 1 15 13
12 1 15 3 10 9 13 13 7 13 10 1 15
7 0 3 10 9 10 9 15
22 7 1 15 3 9 13 7 13 15 13 10 13 15 7 13 10 1 15 0 7 13 15
7 13 1 15 10 9 10 9
15 3 10 9 10 13 15 1 10 9 15 1 10 9 13 15
9 3 0 13 16 13 10 9 10 9
15 13 3 15 16 11 1 10 9 0 0 13 3 10 9 0
6 6 15 11 6 15 11
21 3 16 1 11 7 11 13 10 9 10 13 1 15 3 3 1 9 7 9 13 13
7 7 15 11 3 1 9 13
3 1 11 13
11 10 13 15 15 13 7 10 13 15 15 13
7 13 3 10 12 1 9 13
10 9 3 10 9 13 15 1 10 9 15
3 13 3 15
9 13 10 11 3 9 1 10 9 13
10 3 1 0 3 13 16 10 9 15 13
10 13 3 16 10 9 15 13 1 10 9
12 1 15 10 9 13 1 10 9 10 0 7 13
20 13 15 9 9 10 9 7 10 9 16 13 0 1 0 7 0 7 13 15 0
6 7 13 1 10 9 13
34 15 15 13 1 10 9 15 7 15 13 15 13 10 9 3 3 10 9 7 15 13 10 9 3 3 10 9 7 15 3 13 10 9 13
8 7 13 1 10 9 1 0 13
23 13 3 15 16 0 9 7 9 13 13 15 15 13 7 3 13 7 13 15 13 7 3 13
8 7 6 0 15 13 13 15 13
6 9 15 13 9 0 13
5 15 3 13 1 15
5 1 10 9 15 13
4 15 3 13 13
34 13 9 10 9 15 1 0 10 9 15 7 1 0 10 9 15 7 1 0 10 9 15 7 1 0 10 9 15 7 10 3 15 3 15
2 3 13
4 0 13 7 13
9 15 3 13 13 15 13 1 10 11
5 7 15 13 15 3
4 13 10 11 13
20 9 15 13 1 11 1 11 7 9 13 15 7 13 15 7 9 13 13 13 0
12 3 3 3 9 13 1 10 9 13 7 13 13
12 7 1 10 3 13 12 9 13 10 9 7 13
13 13 15 7 15 3 13 15 1 10 13 15 13 15
13 15 0 10 12 3 13 15 13 10 13 1 10 9
3 15 3 13
6 10 13 10 9 1 15
5 13 3 15 10 11
5 13 7 15 13 3
18 7 0 13 9 13 11 15 3 13 1 10 9 10 9 13 10 9 15
7 10 3 11 13 1 0 9
3 13 3 13
12 9 3 13 15 16 10 9 15 0 15 13 13
6 13 3 15 16 15 13
6 13 3 13 15 10 9
7 11 11 13 7 13 1 0
4 12 3 13 9
19 7 13 1 10 13 15 1 9 15 13 16 13 13 15 10 9 15 1 15
11 9 13 15 13 3 3 11 13 10 9 15
3 13 3 15
3 3 13 13
5 9 13 10 9 15
4 13 10 9 15
10 10 9 15 10 0 13 15 10 1 9
6 7 13 15 10 9 15
4 7 13 1 15
13 15 1 15 13 9 7 13 1 15 9 7 13 15
19 9 13 15 12 9 16 9 15 13 1 9 1 15 7 3 13 15 13 15
5 7 0 3 13 13
4 3 15 9 13
14 3 10 9 13 7 10 9 15 1 15 1 10 9 13
5 3 13 13 13 15
21 16 3 3 13 15 13 1 10 13 9 15 1 3 10 9 15 13 13 15 15 13
4 13 7 13 15
3 13 7 13
4 13 7 13 15
13 15 3 10 13 13 7 10 13 13 7 10 13 13
14 15 3 1 15 10 9 13 10 9 9 3 9 13 15
9 7 7 9 3 1 9 9 15 13
25 16 3 15 0 13 13 9 0 13 10 9 15 15 3 10 9 10 1 9 13 9 0 10 13 15
8 7 13 13 9 7 15 13 0
4 7 13 10 9
5 15 3 1 15 13
9 1 11 10 9 10 9 13 10 9
9 0 3 13 9 1 9 13 1 15
8 15 3 13 15 10 9 13 15
13 16 3 3 10 11 1 15 13 3 13 10 9 15
8 3 13 1 11 13 15 10 9
14 16 3 15 1 11 13 10 9 10 9 15 1 15 13
16 16 3 1 9 9 13 10 9 3 13 1 15 10 9 10 9
14 3 10 0 13 13 10 15 9 1 9 13 10 13 15
19 16 3 0 15 13 13 15 10 9 15 13 1 15 13 7 10 9 15 13
15 10 3 13 1 15 1 15 13 7 10 3 13 1 15 13
7 13 1 10 9 15 3 13
6 7 13 13 13 7 13
23 3 13 7 13 0 9 0 15 12 7 13 13 3 7 13 10 0 10 9 0 0 10 0
16 13 3 1 10 13 15 0 13 15 9 9 1 10 9 13 15
3 15 3 13
10 3 0 10 13 10 9 10 9 7 13
6 10 3 9 13 13 13
12 9 13 7 9 3 13 15 3 3 10 9 11
17 3 3 13 11 10 9 9 3 13 7 10 9 10 9 10 9 0
15 9 9 13 1 10 9 1 10 9 10 9 0 7 13 15
16 3 13 1 10 9 10 9 13 10 9 11 7 6 0 11 3
13 9 9 13 1 10 9 1 10 9 0 7 13 15
20 15 9 13 1 9 13 7 1 10 9 7 1 10 9 16 10 13 10 9 13
8 10 9 10 9 13 10 9 15
9 16 3 0 13 3 10 9 15 0
10 13 3 3 10 9 10 1 15 9 13
23 16 3 10 9 15 0 0 3 13 15 9 0 13 0 0 3 3 10 9 10 9 13 15
11 1 3 10 13 13 15 9 16 13 1 15
3 13 3 13
12 10 3 9 13 13 16 3 0 13 1 10 9
12 3 15 10 9 10 1 10 9 7 10 9 13
10 0 3 10 13 10 3 3 10 3 13
11 3 10 13 13 9 7 6 15 0 15 13
24 7 6 15 10 9 16 13 10 9 7 10 9 7 15 9 7 13 10 9 7 10 9 10 9
7 0 13 13 7 0 3 13
17 6 15 10 9 16 13 10 9 1 10 9 7 10 9 1 10 9
17 6 15 16 13 3 10 9 10 0 7 10 9 10 13 1 3 13
7 13 3 15 10 0 13 15
21 3 15 10 0 6 16 13 10 9 9 0 7 0 12 10 9 15 3 13 10 9
14 6 15 16 13 10 9 10 9 7 10 9 15 13 15
18 3 9 13 7 13 10 9 10 9 15 16 15 3 13 15 15 3 13
8 1 0 7 10 9 10 9 13
42 13 1 15 9 7 9 7 1 15 13 7 13 16 13 10 9 15 10 9 10 13 1 9 9 1 10 9 0 1 9 11 1 9 11 10 13 1 10 9 7 10 9
3 6 13 15
5 13 1 10 9 0
10 6 15 10 0 16 13 10 9 10 9
24 7 3 13 15 13 10 9 7 10 9 3 13 7 13 15 1 0 13 13 15 1 10 9 15
17 1 15 13 10 9 10 9 16 13 15 13 13 1 10 9 15 0
10 13 15 1 10 9 10 9 15 13 9
12 15 3 13 13 15 3 13 7 0 15 3 13
24 1 15 15 1 10 9 13 1 10 9 13 7 15 1 10 9 13 1 10 9 13 1 10 9
6 13 3 15 10 9 15
15 3 13 1 10 13 10 9 7 1 0 3 13 0 15 13
5 13 3 15 15 13
2 0 13
6 3 12 9 13 9 12
10 7 12 1 15 3 13 13 1 10 9
9 7 3 10 9 10 9 15 15 13
2 3 13
3 0 9 13
3 13 3 15
13 10 3 13 15 1 10 9 13 1 10 9 10 9
9 10 3 1 10 0 9 13 3 13
22 3 3 13 15 1 10 9 7 10 9 7 10 9 3 13 3 7 15 13 7 15 13
13 10 3 0 9 13 15 1 15 10 9 15 13 13
7 13 3 15 1 10 9 15
10 9 13 10 9 15 13 1 15 10 9
4 15 3 13 15
4 13 3 1 15
20 13 7 13 1 15 9 16 3 1 10 13 15 10 9 15 13 1 10 13 15
6 9 15 0 13 10 9
5 7 13 1 15 13
10 15 13 16 3 13 3 13 10 9 15
2 7 13
2 0 13
8 9 13 0 0 13 1 9 0
1 13
1 13
1 13
5 13 3 15 10 9
10 0 0 10 9 10 9 15 13 1 15
5 15 3 13 15 13
6 13 3 1 10 9 15
4 1 0 15 13
11 3 13 10 9 15 13 7 10 9 15 13
11 10 9 0 13 10 9 7 10 9 10 9
5 7 10 9 13 15
6 15 3 15 13 10 9
12 15 3 1 15 13 13 13 1 10 9 15 9
8 13 10 9 3 7 13 7 13
3 13 3 15
11 3 11 1 15 10 9 15 13 3 12 0
21 16 3 1 9 10 9 13 3 7 3 1 9 13 10 9 3 13 15 3 15 0
12 7 15 3 13 15 13 7 15 13 7 3 13
8 15 3 10 9 13 16 13 0
9 3 13 10 9 15 7 0 13 15
9 3 13 10 9 15 13 15 10 9
7 13 10 13 15 7 13 9
17 13 15 9 3 13 9 0 1 10 9 3 9 3 13 7 9 13
12 3 3 13 10 9 15 3 3 10 9 15 13
9 13 15 10 9 13 7 10 9 13
20 7 15 0 9 13 10 9 15 3 13 1 10 9 16 13 7 13 3 13 15
12 6 13 15 16 13 7 13 15 7 13 13 15
14 3 15 13 0 16 15 9 3 13 10 9 10 9 13
5 13 3 15 10 11
11 9 1 15 10 9 0 13 7 3 1 15
4 7 13 10 9
22 15 3 13 10 0 9 10 0 15 13 10 9 1 10 9 15 10 13 1 9 10 9
12 0 10 9 0 15 13 10 9 15 13 13 3
11 3 13 15 16 1 15 10 13 15 13 15
10 10 3 3 13 13 3 0 9 13 0
16 15 3 15 13 0 0 13 1 15 7 15 13 0 0 13 15
12 9 13 13 1 10 9 7 15 13 16 3 13
10 9 3 13 13 7 3 13 16 15 13
8 13 16 9 13 13 1 10 9
3 3 13 15
3 7 7 9
17 13 3 1 10 3 12 1 12 9 13 12 1 12 7 12 1 12
5 13 3 3 10 9
14 3 13 9 13 1 9 3 13 16 9 13 7 13 3
10 7 3 9 13 13 16 9 13 7 13
10 9 10 9 10 9 7 10 9 13 13
7 10 3 9 0 3 3 13
9 15 3 7 1 15 3 13 10 0
37 16 3 13 1 10 9 15 1 9 1 10 9 13 9 13 1 15 16 13 15 1 10 9 7 10 9 15 13 10 9 7 10 9 15 13 1 9
2 13 15
4 7 13 13 15
14 13 16 10 0 0 0 1 15 10 0 13 16 0 13
3 3 13 15
7 7 16 3 13 15 3 13
28 7 0 10 12 1 15 13 10 9 1 10 11 7 13 15 13 16 15 9 13 1 15 10 9 10 13 1 11
3 3 13 15
7 7 16 3 13 15 3 13
17 9 13 15 13 1 10 9 15 7 13 13 9 1 15 7 3 13
15 6 12 9 16 15 13 13 9 1 10 9 0 7 3 13
2 13 15
5 3 3 10 9 13
5 15 3 13 13 15
15 9 13 15 3 0 10 9 16 15 13 1 15 7 13 9
8 7 16 3 13 9 1 10 13
10 13 3 13 1 12 10 9 1 10 9
18 7 6 9 9 13 9 9 12 7 13 13 7 3 13 13 1 10 0
6 9 13 1 10 9 15
5 7 13 15 10 9
7 7 3 13 7 13 10 9
22 13 3 10 9 13 16 10 9 13 10 11 13 10 9 16 12 9 13 1 15 13 13
11 1 15 3 13 13 7 3 10 9 10 9
19 9 0 15 10 9 3 13 10 9 15 7 10 9 1 10 9 7 13 13
25 0 3 9 11 13 15 13 10 11 6 12 7 12 9 3 13 13 1 10 9 0 10 9 10 9
22 7 0 13 15 13 15 10 13 15 7 15 10 9 13 1 15 10 0 10 13 1 15
11 15 0 13 10 9 10 9 7 15 13 15
11 0 13 9 9 15 13 9 13 1 9 15
16 7 13 7 13 1 9 7 10 9 10 9 13 1 10 9 15
3 7 3 13
15 0 13 9 15 13 9 13 1 9 9 12 16 15 13 0
12 7 13 1 9 7 9 13 7 9 13 1 11
4 13 3 15 15
5 9 3 0 10 13
15 13 13 1 10 0 9 16 0 13 15 13 13 7 3 13
19 16 15 3 13 10 9 7 13 10 9 7 13 3 13 7 13 10 9 13
3 9 13 15
5 3 13 15 3 13
3 3 13 13
11 13 1 15 7 13 7 1 10 9 15 13
2 7 13
2 13 15
6 13 1 15 15 9 9
29 3 13 10 9 7 10 9 10 9 3 13 11 7 11 7 11 7 15 10 9 1 10 9 10 9 15 3 13 3
13 7 6 13 0 15 13 0 7 13 0 15 13 0
9 1 15 10 9 13 15 9 13 15
9 13 7 13 3 16 11 13 15 13
3 7 13 15
5 13 13 10 9 0
13 6 13 9 7 9 13 3 7 3 7 10 0 13
30 11 11 10 13 10 9 7 13 10 13 1 15 3 13 13 10 9 15 15 9 9 10 15 9 1 10 9 7 3 13
11 13 15 16 3 3 13 15 16 13 3 13
6 13 10 13 1 9 9
21 7 13 1 10 13 15 1 9 15 10 9 10 9 9 13 9 7 15 13 13 15
8 7 6 9 15 13 0 1 15
11 7 13 10 11 13 1 10 0 7 9 13
6 13 10 9 13 7 3
3 15 3 13
17 15 15 9 7 9 1 9 13 7 3 3 13 15 1 9 10 9
6 7 3 13 13 1 0
14 13 3 1 10 13 9 13 3 10 9 13 13 1 15
27 3 13 1 15 1 9 3 13 1 10 9 16 0 15 13 13 1 15 7 13 10 15 7 15 13 13 15
3 13 0 9
9 7 3 13 1 9 10 0 9 13
17 7 3 13 13 13 1 10 0 9 16 3 13 10 13 15 13 15
3 9 13 0
11 3 15 10 13 15 13 7 10 13 15 13
6 13 3 7 10 13 15
30 3 13 9 7 9 3 13 10 9 15 7 10 9 15 7 10 0 15 7 9 0 16 3 15 13 15 7 13 9 15
17 7 3 13 9 13 0 0 0 0 7 0 13 16 3 13 13 15
8 13 3 15 1 10 9 10 0
8 13 3 15 10 13 0 13 15
9 0 15 13 9 1 10 9 10 9
4 15 3 13 15
6 7 13 1 12 15 13
4 10 0 13 15
8 9 13 7 13 9 13 13 15
2 13 15
3 13 15 13
3 7 0 13
8 9 9 13 12 7 13 13 15
3 13 15 13
8 9 13 7 1 0 3 13 13
9 7 13 10 9 13 10 9 15 0
8 3 13 10 9 13 10 9 15
20 13 3 1 10 9 7 9 10 9 7 10 0 7 0 7 0 7 0 13 3
4 7 13 10 9
8 9 13 15 13 7 3 9 13
14 13 1 10 9 7 9 7 13 13 16 13 15 10 9
14 13 3 15 16 15 10 9 0 10 13 13 15 10 9
37 16 15 13 1 15 7 3 13 10 9 15 7 10 9 7 10 9 7 10 9 7 10 9 7 10 9 3 3 7 10 15 9 3 13 13 15 9
15 15 3 13 10 9 15 7 13 1 15 3 13 13 15 9
17 15 3 1 15 13 9 13 3 0 13 13 10 9 16 13 1 9
17 16 3 13 15 9 7 3 13 13 15 10 13 13 15 13 13 16
9 0 10 9 13 13 7 3 13 13
13 16 3 3 3 15 3 13 9 13 13 10 1 9
17 3 3 15 1 15 15 3 13 15 10 15 13 3 13 13 15 9
4 0 3 10 9
8 7 1 9 7 1 9 0 13
3 3 13 15
4 10 13 9 13
12 13 3 15 13 15 10 9 7 10 0 13 15
8 13 3 1 15 10 9 0 13
27 15 9 1 15 13 12 9 7 13 1 15 12 3 13 10 12 1 10 9 7 13 1 10 13 16 13 15
21 7 13 13 1 10 9 15 13 7 13 1 10 9 13 10 9 7 10 9 13 15
9 13 15 16 13 10 9 15 10 13
23 7 15 9 9 13 12 16 13 9 12 3 13 9 7 13 10 9 7 13 3 16 15 13
8 7 13 13 10 9 7 9 13
8 13 15 16 13 10 9 15 13
2 13 3
5 9 15 13 12 9
7 7 13 10 0 15 10 9
8 9 13 15 10 13 9 10 9
5 7 13 15 10 9
15 13 3 15 15 13 9 0 1 10 9 0 7 15 13 13
18 7 13 13 12 10 9 10 9 0 7 13 15 1 10 9 15 13 9
5 1 15 3 13 13
7 15 0 10 9 15 13 9
5 15 3 9 3 13
9 13 13 1 10 9 15 7 13 15
8 9 13 1 10 9 7 1 15
6 3 13 0 13 9 15
7 7 13 13 1 10 9 15
5 13 3 15 10 9
8 9 13 1 10 9 7 1 15
6 3 13 0 13 9 15
8 13 3 10 9 1 10 9 15
25 13 9 10 0 7 13 15 7 13 9 1 10 9 15 7 9 1 10 9 7 13 10 9 10 0
3 7 13 13
9 13 3 10 9 15 10 0 1 9
17 10 9 15 13 7 13 10 9 15 10 9 10 0 16 13 15 13
6 13 3 7 3 13 13
7 10 3 9 15 13 13 15
6 15 3 13 13 10 9
21 6 0 9 13 15 7 3 9 15 13 7 15 3 13 9 16 1 10 9 15 13
19 16 3 10 9 15 0 10 13 15 10 9 1 9 13 13 15 10 0 9
4 15 3 13 15
12 9 15 3 1 15 13 7 15 10 15 15 13
6 13 3 7 1 10 9
16 9 15 13 0 15 13 9 7 0 13 15 3 13 10 13 15
5 7 13 15 13 15
5 15 0 13 1 15
6 13 10 9 10 9 15
5 3 3 13 3 13
6 13 3 1 15 10 9
11 15 13 16 10 9 15 13 10 9 1 15
15 13 15 13 16 3 13 1 10 9 13 15 1 10 9 15
12 7 13 12 0 10 9 10 9 15 13 10 0
5 15 13 10 9 15
3 15 3 13
3 12 9 9
4 15 3 13 15
9 13 15 10 9 7 13 3 13 12
4 15 3 15 13
3 12 9 9
2 13 15
7 13 15 10 9 7 13 12
11 7 13 10 9 10 9 10 9 16 3 13
18 3 10 9 10 9 0 0 1 10 9 10 9 1 10 9 10 15 13
4 7 15 15 13
19 10 0 1 0 3 1 0 0 13 7 10 1 0 0 3 1 0 0 13
14 16 3 1 10 0 9 0 3 13 10 0 15 15 13
6 15 9 13 12 9 13
16 7 3 10 12 13 7 10 0 13 7 12 13 7 10 0 13
6 3 13 9 13 7 9
11 13 3 0 15 10 9 0 13 7 13 15
3 7 13 15
7 10 3 9 13 10 9 15
9 3 10 1 9 0 9 1 10 9
7 10 9 7 10 9 1 11
15 0 3 13 10 9 7 10 9 13 3 10 9 12 9 13
17 15 10 13 10 9 15 7 13 0 13 7 10 13 1 9 13 13
14 9 3 15 13 0 7 13 9 7 9 13 1 9 3
22 0 3 15 9 11 13 1 10 9 15 13 7 13 13 1 10 13 1 10 9 10 0
15 13 3 13 10 0 7 13 15 1 10 9 1 10 9 11
7 13 3 3 10 0 7 13
21 7 1 10 11 13 10 9 15 13 1 9 13 11 1 3 7 11 1 10 9 15
4 7 15 13 13
3 13 3 11
16 9 13 16 13 10 0 15 1 10 9 15 7 11 3 10 0
4 3 3 3 13
26 7 1 15 0 1 15 7 15 9 0 13 16 10 13 13 3 1 15 3 13 7 10 3 1 15 13
2 13 3
31 13 3 15 9 16 13 15 1 10 9 10 9 15 13 3 12 9 16 13 15 16 3 3 15 13 1 10 9 0 10 9
4 13 3 15 11
5 13 11 7 10 9
3 15 3 13
12 3 9 11 7 16 15 1 0 13 1 15 13
14 16 11 7 10 9 3 13 3 16 15 1 0 13 13
6 13 3 1 10 9 15
12 0 13 10 10 9 3 13 6 3 1 15 13
22 13 15 16 9 0 13 1 10 9 15 7 13 1 10 9 3 16 13 10 0 10 12
2 13 15
12 16 13 10 9 15 13 15 7 16 13 13 15
6 7 13 10 9 10 9
4 13 3 10 9
11 16 13 9 3 9 9 13 3 10 0 0
6 13 7 13 1 10 9
4 7 13 3 15
16 15 3 1 15 9 13 13 7 13 15 13 1 10 9 13 15
3 3 13 13
4 7 3 13 15
11 3 3 15 3 13 15 10 13 15 13 16
3 9 0 13
4 15 13 13 13
15 7 13 1 10 13 1 11 7 15 13 1 0 11 7 11
19 7 13 15 1 15 9 13 15 12 0 9 15 13 3 7 15 13 9 13
4 11 9 13 15
4 7 13 13 15
5 13 13 15 10 9
24 12 3 1 15 13 16 13 13 1 9 0 13 10 9 7 13 1 9 1 10 9 15 13 15
4 7 15 13 9
5 13 3 10 11 13
4 3 10 12 13
3 10 12 3
12 3 13 13 13 9 10 9 3 3 10 0 0
3 7 13 15
2 13 13
14 3 13 10 9 10 9 1 9 7 13 6 3 7 3
9 6 3 10 9 10 9 1 15 13
5 13 3 1 10 9
15 13 9 3 13 12 10 9 10 9 10 9 13 7 3 13
3 7 13 15
2 6 3
2 6 3
25 3 3 10 9 13 1 10 1 10 9 1 10 1 9 13 3 13 10 9 10 9 1 10 9 15
17 7 3 13 1 10 9 11 3 13 7 1 10 9 10 9 10 9
19 13 13 13 13 1 15 9 13 11 1 10 9 7 13 10 9 7 13 0
7 3 3 13 1 10 9 11
1 13
1 13
1 13
1 13
1 13
11 1 10 15 13 15 9 10 9 10 9 13
30 1 0 10 9 15 13 1 10 9 7 10 9 15 1 10 9 3 13 13 15 7 10 1 9 3 3 13 1 10 3
4 13 10 9 11
15 15 3 13 10 9 15 13 13 15 7 15 3 13 13 15
2 13 15
6 12 13 7 10 0 13
6 13 12 13 1 10 15
3 10 12 13
4 7 13 13 15
2 3 9
4 15 3 13 15
8 3 10 9 3 7 10 9 13
14 9 15 13 1 15 9 10 9 3 13 7 9 3 13
12 9 3 13 1 10 9 0 7 13 1 15 13
6 13 15 1 10 9 15
5 7 3 13 1 9
27 16 3 10 9 3 13 7 9 13 1 3 10 13 15 9 10 9 0 13 15 16 3 1 9 13 13 15
4 13 3 10 9
7 13 15 10 9 10 9 13
9 13 15 16 13 10 9 15 1 9
13 3 10 9 10 9 13 3 13 10 9 1 10 9
19 13 3 7 1 15 10 13 1 15 16 13 0 7 13 10 0 10 9 0
7 9 12 13 1 10 9 13
7 10 12 9 7 10 0 9
21 10 9 13 15 16 3 13 3 10 0 10 9 0 0 9 7 3 3 0 10 9
4 13 3 10 9
20 10 3 9 3 13 3 13 3 10 9 13 1 10 9 7 13 10 9 15 13
6 10 9 13 15 10 0
2 13 15
10 13 0 13 1 10 9 15 3 3 0
11 3 15 10 13 15 13 10 3 13 15 13
9 13 3 15 3 10 9 16 15 13
6 10 3 11 13 15 13
8 10 3 0 13 10 9 10 9
3 6 13 15
15 15 3 3 13 10 9 10 9 3 9 3 3 13 1 15
6 7 13 15 15 9 13
7 9 0 15 13 9 0 13
5 13 3 15 10 11
4 15 15 13 0
2 3 13
2 3 13
2 3 13
2 3 13
8 13 10 9 15 7 10 9 15
3 15 3 13
5 0 15 13 1 9
6 13 3 10 11 13 15
16 15 15 13 13 7 13 0 7 13 9 1 9 7 6 13 15
6 15 3 13 0 0 13
4 13 3 0 3
6 13 3 15 10 11 13
12 3 3 10 10 9 13 1 10 9 10 9 13
16 0 3 13 9 1 9 9 13 3 0 1 10 9 10 9 13
4 13 3 10 13
4 7 15 13 13
3 13 3 11
7 6 15 13 10 0 13 15
4 15 3 13 15
3 6 13 15
35 15 13 15 13 9 7 9 7 9 7 9 7 9 1 10 9 10 9 15 3 3 13 0 1 10 9 0 7 1 10 9 10 13 9 0
7 13 3 10 12 13 1 15
16 6 13 1 11 7 13 15 10 13 1 10 9 10 9 10 9
18 7 15 15 0 13 7 13 10 9 0 13 1 15 7 3 13 10 13
8 13 3 9 13 13 15 13 0
8 13 3 15 16 11 10 0 13
3 7 13 13
5 11 9 11 13 15
7 7 10 13 13 15 16 13
5 15 3 0 3 13
9 13 3 10 11 13 15 13 1 15
5 13 3 15 13 15
3 15 3 13
3 9 16 13
5 7 10 11 13 15
1 13
5 10 9 15 13 15
9 7 15 10 9 13 13 9 10 9
5 7 13 13 10 11
6 7 6 9 9 13 11
18 7 13 13 10 11 15 13 7 3 13 1 10 9 16 10 9 0 13
15 7 13 1 10 3 13 1 9 16 13 15 16 0 13 13
12 7 16 13 1 10 9 13 10 11 13 1 15
3 11 13 13
7 7 13 13 7 13 15 13
11 7 13 15 13 13 16 1 0 9 13 13
7 13 3 11 13 1 10 9
17 6 10 0 15 10 13 9 10 0 13 7 16 15 15 13 13 9
11 3 9 10 9 0 13 16 3 15 9 11
11 13 3 10 9 10 9 13 7 13 10 13
24 13 3 15 0 13 13 9 1 10 3 13 11 15 7 13 15 16 3 13 10 9 10 9 13
12 9 15 0 13 1 9 3 13 15 9 7 13
13 13 3 12 9 15 13 15 12 9 7 13 1 15
4 13 1 15 13
12 10 3 9 15 13 15 7 13 9 1 15 13
6 3 13 0 13 1 15
5 13 3 10 0 13
7 9 10 9 15 12 13 9
14 3 0 9 16 1 0 0 13 13 9 13 1 12 9
5 7 13 10 0 13
7 10 9 15 9 13 12 9
4 13 3 3 0
6 3 15 1 13 12 9
5 7 10 0 13 13
7 13 3 15 16 9 0 13
2 13 15
8 1 10 9 15 13 15 0 9
15 13 16 15 9 0 13 13 15 3 13 7 13 15 3 13
10 7 1 15 3 13 15 10 9 1 9
8 7 15 13 1 9 3 15 13
4 7 10 13 13
12 13 1 15 10 9 7 13 10 10 12 9 13
7 13 15 16 15 10 13 13
9 1 3 10 3 13 7 15 13 13
19 3 10 0 15 0 10 3 13 15 13 1 15 13 3 7 13 15 1 15
8 7 13 0 13 3 13 1 11
19 7 13 16 13 1 11 7 11 1 10 9 10 13 9 13 12 10 9 13
21 13 1 10 1 9 1 15 13 13 9 13 1 15 15 3 9 13 7 13 15 13
10 7 16 15 15 13 1 15 13 3 13
6 16 10 9 15 9 13
11 13 3 15 10 9 13 10 9 15 1 15
4 15 13 10 9
3 15 3 13
6 16 10 9 15 9 13
17 7 13 15 1 10 11 7 13 15 10 9 1 10 9 13 10 11
10 13 3 15 13 10 9 15 1 10 9
29 13 3 15 3 1 10 9 10 9 10 9 13 0 10 9 10 9 13 13 10 9 9 0 1 15 15 13 9 13
6 13 10 9 1 9 9
5 9 13 10 9 15
3 7 13 13
9 13 15 16 16 0 13 10 9 13
11 7 16 13 13 10 9 13 1 15 13 16
14 3 13 3 15 3 1 10 9 15 0 10 1 9 15
6 3 3 13 1 9 15
45 3 13 9 1 15 7 13 10 0 15 9 15 7 13 15 7 13 15 3 7 13 15 7 10 9 15 1 15 7 3 13 9 1 9 1 15 16 15 3 13 10 9 10 9 15
1 13
6 15 3 15 13 9 9
9 7 13 13 10 1 9 1 10 9
20 10 3 9 7 10 9 13 15 13 7 10 0 10 9 7 3 13 10 15 13
7 10 9 3 0 13 15 13
29 7 13 1 12 10 9 13 15 10 9 1 10 9 7 13 13 10 9 7 10 9 1 10 0 7 13 13 1 15
16 13 15 1 15 9 0 13 7 15 13 10 13 15 10 9 0
8 13 15 3 15 9 7 13 15
10 10 9 10 11 1 9 13 7 1 9
5 16 13 1 9 13
5 1 15 3 13 15
10 16 3 13 1 9 10 9 0 13 15
6 13 3 13 11 9 13
5 7 13 3 13 3
9 3 15 13 15 1 15 9 0 13
9 13 3 1 10 9 13 10 9 0
11 9 13 9 7 13 15 9 7 13 9 0
7 10 3 9 13 15 13 0
5 7 13 0 13 9
9 15 3 7 0 13 7 13 13 0
4 7 13 0 13
6 13 3 10 9 10 9
2 15 13
6 13 10 9 15 10 0
3 3 0 13
4 0 13 10 9
7 13 15 16 15 13 10 9
7 7 13 15 1 10 9 13
11 13 7 13 10 9 0 7 13 10 9 0
3 13 3 13
2 3 13
5 15 3 13 15 13
6 15 3 13 10 13 0
8 15 10 13 1 0 10 9 13
7 1 15 3 3 13 13 15
9 13 3 16 1 15 13 10 9 0
22 7 13 13 0 13 15 0 13 16 13 15 9 16 13 15 10 9 7 10 9 10 9
4 7 13 15 13
19 9 13 16 3 13 7 13 7 3 13 9 7 1 9 10 9 10 9 13
7 13 15 9 9 13 7 3
8 13 3 15 10 9 13 1 15
5 15 13 9 7 9
1 9
5 15 3 13 1 15
11 3 13 10 9 9 7 10 10 9 10 9
16 7 3 13 13 15 9 1 10 9 7 13 1 10 9 15 13
13 13 3 15 10 9 10 13 9 3 13 13 15 13
27 9 11 13 15 16 15 9 13 13 9 7 0 0 13 16 13 10 9 15 10 9 7 13 9 10 9 15
4 12 3 9 13
10 3 3 3 10 12 3 13 9 7 13
5 0 3 10 9 13
10 10 9 3 1 10 9 15 15 13 9
6 10 3 12 13 15 9
5 7 13 15 10 11
8 10 9 10 9 0 13 7 13
17 10 3 13 10 9 0 13 7 10 9 10 1 0 7 13 7 13
5 7 3 13 3 13
23 16 3 13 10 0 3 11 13 1 10 9 16 13 9 10 9 11 7 9 11 7 9 11
7 9 3 3 13 0 7 13
4 15 3 15 13
6 13 3 15 10 9 13
3 9 3 13
6 3 3 13 13 15 15
4 13 3 1 15
7 3 13 10 11 13 11 9
14 13 1 0 15 16 3 13 10 0 15 9 10 9 15
10 11 3 9 15 13 7 3 15 9 13
8 13 3 15 10 9 13 10 9
35 13 1 10 9 10 13 13 1 9 7 13 9 1 10 9 7 9 1 10 9 7 9 1 10 9 15 13 10 9 10 9 7 9 0 13
4 0 13 0 9
12 13 3 13 10 13 1 10 9 10 9 15 0
11 13 3 15 9 0 13 3 12 9 7 13
11 0 3 0 1 10 13 15 13 1 10 9
13 7 15 13 1 10 9 16 9 0 7 9 13 13
15 0 15 13 13 9 1 15 3 13 9 1 9 15 3 13
4 13 3 15 13
5 9 3 3 0 13
8 7 15 10 9 3 13 0 13
3 15 3 13
8 0 3 13 1 10 9 15 13
6 15 13 7 10 9 13
8 3 3 13 9 7 9 3 13
10 13 3 0 13 0 7 3 3 10 9
3 3 13 15
8 13 9 1 9 7 9 1 9
10 9 7 0 7 1 9 9 7 9 13
27 1 3 0 15 13 1 15 10 9 15 7 13 13 1 10 9 7 9 13 1 9 7 9 1 10 9 15
4 13 15 1 9
9 13 3 1 10 9 15 3 13 13
24 13 3 7 1 9 7 9 7 0 7 9 7 13 1 15 7 13 13 1 15 1 10 9 15
9 7 9 1 10 9 15 3 3 13
8 1 10 9 15 13 10 9 15
14 3 3 13 13 1 9 11 3 13 16 13 10 9 15
12 6 10 1 9 13 7 10 13 1 0 10 9
33 13 3 9 0 1 10 9 7 9 10 9 0 7 13 9 9 7 13 1 10 9 15 7 11 13 13 1 9 16 15 13 9 9
31 7 13 9 1 9 7 9 7 9 7 1 10 9 9 9 1 9 9 9 7 9 13 9 1 9 7 9 10 13 10 9
6 10 3 9 10 9 13
15 13 3 0 13 13 7 13 10 9 15 16 13 10 9 15
4 7 13 9 15
7 13 10 9 7 15 10 9
15 3 3 15 3 13 0 13 13 16 3 13 10 9 10 9
14 6 13 15 16 3 3 13 10 9 0 16 3 15 13
6 10 9 7 10 9 13
7 10 3 9 15 3 3 13
25 13 3 15 16 13 15 10 9 1 9 7 9 7 9 0 7 13 1 15 0 10 9 0 3 9
21 13 3 1 15 9 13 16 13 13 0 15 10 13 13 7 13 1 10 9 10 9
8 13 3 10 9 1 10 9 13
12 7 15 10 9 13 1 15 1 10 9 13 15
20 13 3 10 9 10 0 10 13 9 7 13 10 9 7 10 9 10 3 13 15
4 13 3 10 9
14 13 3 11 1 11 10 13 11 13 1 10 9 10 12
12 7 13 13 10 9 7 9 10 3 15 13 15
7 7 13 7 13 15 9 13
18 13 3 10 9 10 0 1 15 13 13 10 9 7 13 11 7 11 13
4 15 3 13 15
3 3 13 13
4 15 3 13 15
12 6 13 15 1 10 9 13 15 9 9 9 13
8 13 15 1 10 9 1 15 13
6 7 13 10 9 10 9
4 13 15 10 9
2 3 13
10 13 3 13 3 13 15 7 13 10 9
11 7 16 13 10 9 13 7 10 9 1 15
4 7 13 1 15
12 9 13 0 10 9 13 1 15 1 10 15 13
17 13 3 15 16 3 3 3 13 15 16 15 13 1 10 9 10 9
5 7 13 9 13 13
6 13 0 7 13 1 15
9 7 13 9 13 13 7 13 15 13
9 0 13 10 9 15 10 1 15 13
5 0 13 1 15 9
8 7 10 9 3 1 10 13 13
14 0 10 9 10 0 9 1 10 9 15 10 1 15 13
12 3 6 10 9 10 13 15 1 15 1 10 9
18 3 10 9 3 10 9 1 10 13 13 3 6 10 9 0 1 15 13
16 7 15 13 13 1 15 10 15 3 13 1 15 10 0 13 13
12 10 9 10 9 13 15 7 10 13 15 9 13
4 15 3 3 3
15 7 10 0 1 15 13 3 10 0 7 10 13 3 10 13
8 15 3 0 10 13 7 10 13
3 3 10 13
9 15 3 1 0 15 13 3 10 13
11 15 3 13 10 13 1 15 1 10 9 15
12 11 11 6 10 11 13 15 10 13 3 10 9
8 7 15 3 13 13 10 9 15
4 15 3 13 15
12 9 1 15 0 13 7 1 9 7 1 9 13
3 15 3 13
2 13 15
11 11 3 13 3 9 16 3 13 3 13 15
12 16 13 15 1 9 7 9 7 9 3 15 13
3 15 3 13
4 15 3 13 15
20 7 3 10 13 9 13 3 7 9 7 10 3 13 13 10 9 15 7 13 9
12 13 3 15 16 0 10 13 13 13 1 15 0
4 7 1 0 13
7 7 3 10 1 15 9 13
5 9 6 9 3 12
4 15 3 13 15
2 0 13
6 13 3 15 3 10 9
7 13 3 1 10 9 13 15
5 13 3 13 1 9
14 7 15 13 1 15 3 9 9 7 13 10 9 13 13
9 3 3 10 9 15 7 10 15 13
8 13 3 15 9 1 9 13 15
6 7 13 1 9 3 13
12 7 13 10 9 15 3 9 9 13 1 10 9
2 15 13
7 13 13 16 3 13 1 9
20 3 15 13 6 9 7 10 13 11 12 10 12 13 15 7 13 10 11 13 15
7 11 9 10 9 10 9 13
8 13 3 10 1 15 10 13 13
5 9 3 13 1 9
17 7 13 12 15 1 15 10 9 10 9 7 13 10 9 15 10 0
5 13 3 10 11 13
6 7 13 10 9 13 15
15 13 3 11 1 10 13 1 15 9 7 9 10 9 7 0
15 1 9 13 15 1 15 1 10 9 3 13 10 9 1 15
11 7 0 13 15 10 9 7 10 9 10 9
11 13 3 15 13 7 13 1 10 9 10 9
5 10 3 11 13 3
14 13 3 9 1 0 10 9 7 13 13 10 11 0 15
13 13 3 15 9 15 13 1 10 9 7 13 15 13
5 15 3 13 15 13
7 7 1 0 0 13 15 13
5 3 15 1 15 13
4 15 3 11 13
3 9 3 13
9 7 13 3 9 12 0 15 13 13
7 1 9 3 0 1 15 13
4 7 3 0 13
26 7 3 3 13 15 13 9 7 13 10 9 13 10 11 7 13 10 11 10 9 10 9 3 13 15 16
7 16 9 13 3 13 15 3
5 7 13 3 13 3
14 7 10 9 10 13 15 13 15 13 7 13 15 13 13
6 13 15 13 10 13 15
7 7 0 0 13 13 1 15
21 7 16 13 9 13 10 9 10 9 9 7 7 9 7 13 15 1 10 9 15 13
7 16 15 13 10 11 13 15
6 16 15 13 3 3 13
6 16 3 13 3 3 13
16 1 10 3 3 13 10 9 10 9 13 1 0 10 9 10 9
3 13 3 15
7 15 3 13 10 9 10 9
5 15 3 1 15 13
5 15 13 16 15 13
3 15 3 13
11 7 13 0 10 9 15 13 15 1 10 11
5 13 3 13 15 13
17 0 13 13 10 9 15 7 13 9 9 13 7 13 15 11 9 13
6 10 3 11 13 15 13
6 15 13 10 9 10 0
5 15 3 13 15 13
2 15 13
7 15 13 0 1 10 9 0
30 11 3 13 13 16 10 9 0 13 7 13 16 1 10 9 11 13 13 15 1 11 13 3 15 1 11 1 0 10 9
8 10 3 11 13 10 11 13 3
21 13 3 1 0 9 13 13 15 1 10 13 1 15 7 13 15 9 13 1 15 13
6 13 3 15 1 9 0
5 15 3 15 13 15
10 13 3 10 9 7 10 9 3 13 15
15 13 3 9 10 7 11 7 10 11 1 15 10 9 1 15
7 13 3 1 9 13 1 15
26 13 15 10 9 0 3 13 10 9 7 6 15 1 15 13 15 13 1 10 9 0 0 15 13 1 15
3 7 7 11
5 13 3 15 1 15
8 7 6 15 0 9 13 13 15
4 13 3 15 13
2 13 0
5 13 3 15 10 11
15 15 13 1 9 15 13 1 10 9 7 9 13 1 10 9
4 15 3 13 13
1 13
2 13 15
6 15 3 0 13 1 15
6 15 0 9 13 1 15
4 13 3 15 13
13 15 3 13 9 0 13 15 13 7 13 10 9 15
7 7 11 13 13 10 9 15
7 10 3 11 13 10 9 15
19 7 16 13 15 13 11 15 0 13 1 9 13 15 10 9 13 1 10 11
14 13 3 15 0 9 10 9 7 9 15 13 7 13 15
6 9 11 3 13 1 15
16 3 1 15 13 7 1 10 9 15 16 6 13 9 1 15 13
14 0 10 9 7 10 9 15 3 13 7 9 15 3 13
5 3 13 13 10 9
3 13 1 15
2 13 15
13 3 16 1 10 0 9 0 13 1 10 0 15 13
22 7 16 13 1 10 9 10 13 9 3 13 15 7 10 0 15 3 1 0 15 3 0
4 10 3 11 13
3 9 13 15
5 3 3 13 15 13
7 13 3 10 9 15 13 9
5 7 13 10 9 13
2 15 13
12 13 3 15 7 10 9 13 9 13 15 7 13
9 16 15 13 10 9 10 0 13 15
6 13 3 7 9 1 15
5 10 9 10 0 0
7 12 3 10 13 0 13 15
5 3 15 13 10 11
4 13 15 7 15
4 7 15 3 3
5 0 3 15 13 13
5 0 3 15 0 13
2 7 13
9 11 13 15 3 13 1 10 9 15
3 7 13 15
3 6 15 13
7 3 1 15 13 1 10 9
7 13 3 10 9 10 9 0
7 7 13 9 0 10 11 13
8 9 1 9 15 13 10 9 15
4 0 3 13 13
10 13 3 10 9 10 13 13 10 9 13
6 3 10 9 0 0 13
16 7 15 10 13 9 1 10 9 0 13 10 13 13 10 9 13
18 13 3 15 10 0 15 1 3 7 9 10 13 15 1 10 11 13 0
7 7 9 13 9 7 9 13
19 13 3 9 15 13 13 1 10 11 15 13 10 9 7 3 13 10 9 15
6 13 3 13 9 7 9
8 7 10 3 9 13 1 10 9
15 10 3 12 10 9 9 0 1 10 9 13 13 15 13 9
8 13 3 10 9 13 1 10 9
9 13 3 3 13 10 9 10 9 11
9 7 6 9 12 13 15 1 9 13
7 15 13 10 13 1 10 0
5 3 13 3 7 13
28 13 3 13 15 3 13 1 10 11 13 10 9 10 9 16 13 13 1 9 9 0 7 13 7 10 0 9 13
19 7 13 10 9 15 7 13 1 10 9 13 15 0 10 12 7 15 10 0
16 13 3 10 9 11 7 11 7 11 10 11 7 10 0 1 15
5 13 1 10 9 0
31 7 6 12 1 15 1 15 10 9 13 13 1 9 13 9 12 1 11 15 9 11 7 15 13 1 15 1 15 10 13 0
14 7 13 1 10 13 15 7 13 7 0 11 13 13 15
4 13 3 1 15
9 15 10 9 0 15 13 1 15 13
3 7 13 0
9 13 3 12 15 9 11 13 1 15
15 15 0 13 11 7 3 13 10 13 1 15 1 10 9 0
1 15
4 15 3 13 15
37 10 1 11 10 9 15 13 9 9 0 1 9 7 9 1 10 9 7 15 10 9 3 7 13 15 10 9 7 10 9 15 1 9 9 7 13 15
14 7 3 7 1 15 0 0 0 9 13 16 15 0 13
8 7 7 9 15 1 15 13 15
21 13 0 1 10 9 7 3 13 10 9 15 13 13 3 9 9 13 15 13 15 13
17 7 13 15 10 1 15 1 10 9 7 13 3 3 7 10 9 13
5 7 15 13 1 15
14 6 0 7 0 10 9 10 13 1 15 15 13 10 9
12 3 0 13 13 10 11 7 13 1 10 9 15
18 7 13 1 11 7 1 15 10 9 13 15 1 15 10 9 10 1 15
4 7 13 15 13
12 13 1 15 16 1 9 13 7 13 3 10 9
6 7 13 10 13 1 15
8 15 3 13 10 9 7 13 15
6 7 15 0 13 1 15
4 7 13 1 15
19 3 10 9 15 13 13 1 15 16 13 15 1 10 9 16 13 15 10 9
26 7 13 15 10 9 13 1 11 7 13 13 10 12 7 10 1 15 13 16 3 13 10 9 7 13 11
9 0 3 15 13 0 13 1 0 15
8 13 3 7 0 13 13 9 13
12 15 13 13 7 1 15 9 13 1 10 9 15
12 13 10 9 15 7 10 9 15 16 15 13 0
15 13 15 7 13 16 9 9 7 9 3 13 3 15 13 13
11 3 3 13 15 1 10 9 7 13 13 15
4 13 15 0 3
7 15 3 13 15 9 0 9
4 13 3 1 15
9 3 13 15 10 9 10 13 10 9
33 7 13 15 16 3 13 13 10 11 7 13 1 0 10 0 9 7 13 1 10 9 15 9 1 9 9 1 15 10 9 13 1 11
3 15 9 0
10 7 15 13 10 9 10 9 15 1 15
12 15 3 13 1 10 9 16 15 13 1 9 9
13 13 3 15 1 1 11 7 13 10 9 15 13 15
27 7 13 1 10 13 15 15 13 1 15 7 15 13 1 11 1 9 0 7 13 3 1 10 9 13 10 9
12 15 1 15 13 7 1 15 13 3 12 15 13
12 1 15 9 13 7 10 9 13 10 9 10 9
13 7 10 9 1 10 9 13 7 10 9 15 3 13
5 13 9 13 1 9
3 9 15 11
14 0 13 1 9 16 13 1 10 9 16 15 13 1 15
11 3 13 0 10 9 7 16 13 1 10 9
13 13 10 9 10 0 15 13 15 9 13 1 10 9
10 1 10 0 13 7 10 0 15 3 13
32 15 3 13 15 13 15 9 9 9 13 10 13 1 10 9 15 15 3 1 9 7 1 9 9 7 1 9 9 7 1 9 13
23 7 10 9 9 13 7 13 1 15 7 13 10 9 15 9 3 0 1 9 0 9 7 9
7 11 13 1 15 7 13 13
4 0 13 15 13
11 10 1 15 13 1 15 13 16 0 15 13
12 3 1 10 9 15 15 15 13 7 9 1 9
6 3 10 9 1 11 13
12 10 0 9 10 13 1 10 9 10 9 0 13
19 7 0 13 10 9 10 11 16 13 10 0 1 11 9 7 9 16 13 15
3 15 15 13
8 7 13 7 3 13 7 13 16
5 15 3 13 10 11
3 7 13 15
2 15 3
1 13
4 10 9 13 15
2 7 13
1 3
3 13 3 15
2 15 13
6 16 9 13 10 13 15
1 13
6 15 9 13 1 10 0
6 7 13 13 1 10 9
6 7 13 15 7 13 15
14 15 3 13 16 15 3 13 10 11 7 11 7 10 9
5 13 15 10 11 13
4 15 13 1 9
16 10 1 15 13 15 3 13 15 0 16 13 15 10 9 10 9
12 0 1 11 13 1 10 11 3 13 10 11 13
10 10 3 13 10 11 13 1 15 7 13
6 0 13 1 15 15 13
12 1 15 13 9 15 1 15 13 16 0 15 13
17 7 15 3 13 15 7 16 13 10 11 1 0 13 15 1 9 13
5 7 13 11 13 16
15 7 15 3 13 15 7 10 13 15 13 1 9 0 15 13
18 1 15 3 13 10 9 13 7 13 1 15 0 13 10 13 1 9 0
12 7 15 13 7 13 16 0 13 10 9 10 9
18 10 3 3 13 10 11 7 1 10 9 15 12 7 13 10 11 13 13
10 13 10 12 9 15 13 7 13 10 11
9 13 10 11 7 13 15 13 13 15
2 15 13
7 9 15 13 13 9 3 13
2 13 15
3 13 7 13
13 13 3 7 13 3 13 7 1 15 13 10 9 0
4 9 13 3 0
11 13 0 0 10 9 10 0 11 7 13 15
7 13 10 11 15 13 13 11
5 13 15 10 11 13
6 15 13 11 10 9 11
6 15 13 11 15 13 11
10 10 3 13 13 1 10 11 7 13 11
5 7 13 15 10 11
2 13 15
7 13 11 10 11 7 13 15
3 13 15 11
6 1 11 13 15 0 13
3 13 15 11
3 13 7 13
11 13 11 10 11 13 1 15 7 13 1 15
8 13 3 9 1 15 9 3 13
3 13 15 11
11 1 10 15 11 13 13 1 10 9 13 15
3 13 15 11
7 9 15 13 10 9 10 9
5 15 9 13 10 11
5 13 11 7 13 15
10 16 13 15 16 13 15 1 10 9 13
3 0 0 13
3 7 13 15
17 13 10 9 13 7 10 9 10 9 13 7 13 1 10 9 10 9
18 7 10 9 10 0 9 13 1 11 10 11 7 13 10 9 10 11 3
12 13 3 7 10 11 7 10 9 15 1 10 9
10 7 9 3 13 16 13 10 9 10 9
8 3 13 10 9 10 11 1 15
3 9 3 13
4 13 15 10 11
5 15 15 7 15 9
5 15 3 13 15 13
18 13 3 3 0 9 12 1 10 9 10 0 13 13 1 9 12 7 12
4 13 15 10 11
4 13 10 9 9
5 7 13 15 1 3
3 7 13 15
6 13 3 7 13 10 9
30 16 3 13 10 9 10 9 9 13 7 3 13 3 13 10 3 9 13 10 13 10 9 13 10 9 10 9 7 13 15
7 15 13 10 0 9 1 3
23 0 13 9 10 9 10 11 1 11 10 11 7 13 10 9 15 7 13 1 15 10 9 15
24 1 0 13 1 11 15 7 10 9 15 7 10 9 15 7 10 9 15 7 3 13 3 0 9
13 7 3 13 10 9 10 0 7 13 1 11 10 11
48 7 13 1 10 9 10 13 9 7 9 7 9 7 10 9 13 7 13 9 1 9 15 13 1 10 9 10 7 9 7 10 9 7 10 9 13 10 9 7 10 9 13 7 10 10 9 13 13
3 13 0 3
7 13 10 9 15 16 13 13
7 10 9 10 9 15 13 15
7 15 9 13 15 16 0 13
5 13 11 7 13 15
10 13 10 9 0 7 1 12 9 13 15
4 13 3 10 0
15 12 7 12 9 13 10 9 0 7 15 1 12 9 13 15
23 16 3 13 1 0 13 10 9 15 16 0 13 7 13 10 9 7 10 9 15 13 10 11
24 16 3 13 1 10 11 1 10 9 1 10 9 0 13 1 10 9 15 13 15 10 9 15 13
23 0 3 11 3 13 15 15 1 10 15 13 15 7 16 3 9 13 16 15 13 1 10 9
12 13 3 9 1 10 9 11 9 15 9 10 0
8 0 13 1 15 9 7 13 15
7 9 13 16 1 9 13 9
17 15 3 13 0 10 9 13 15 15 13 16 3 13 10 9 1 15
4 6 6 13 15
12 16 3 15 13 3 3 13 13 10 9 10 9
5 13 1 15 10 11
6 3 13 9 13 9 13
2 13 11
4 6 6 13 15
16 16 3 15 13 1 9 7 9 3 13 13 1 10 9 10 9
5 3 13 16 13 15
4 13 15 13 3
18 10 9 3 13 13 7 10 9 15 13 7 3 13 3 13 7 3 13
8 3 13 15 10 13 1 10 9
5 13 11 7 13 15
5 13 11 7 13 15
10 15 13 10 9 10 11 7 0 3 13
15 16 10 0 13 15 7 3 13 3 16 13 15 10 0 13
22 7 15 13 1 10 9 3 3 10 1 10 9 13 10 9 10 9 10 13 1 10 9
25 7 3 11 13 10 9 1 10 0 3 13 13 10 9 10 9 16 15 10 13 1 15 13 9 0
25 3 3 13 10 9 10 9 16 10 9 10 0 13 16 15 10 13 1 15 3 13 7 13 9 0
21 3 3 13 10 9 10 9 1 10 9 16 13 10 9 7 16 13 10 9 1 15
6 10 13 1 15 3 13
22 0 3 13 10 9 16 10 9 13 1 10 9 7 13 10 9 3 10 9 3 10 9
20 15 3 10 0 13 13 10 9 7 3 13 1 10 9 16 3 13 10 9 15
19 10 3 13 10 9 13 1 10 9 16 13 15 10 9 16 1 9 13 13
20 1 0 13 10 11 7 10 9 15 1 10 0 9 7 3 13 1 15 7 13
19 13 3 7 11 13 1 11 3 10 11 16 9 0 13 3 7 13 7 13
8 3 3 13 13 1 10 9 11
11 13 3 9 1 10 9 11 1 0 1 9
8 7 13 1 10 11 7 13 15
13 3 13 9 13 15 16 3 13 13 15 1 10 9
6 0 15 15 13 16 13
11 3 13 15 10 11 7 16 13 13 1 0
6 10 13 10 9 9 13
17 10 3 9 10 9 10 13 7 13 15 9 13 1 10 9 10 9
7 0 3 10 9 10 15 13
6 0 13 13 15 3 13
6 10 3 13 1 15 13
16 10 1 10 9 13 15 13 7 13 13 7 10 9 15 15 13
11 10 13 15 10 9 13 16 10 9 0 13
10 15 3 13 10 9 10 9 10 9 13
7 3 3 1 9 13 10 9
12 10 9 13 10 9 7 15 13 1 10 9 15
8 10 13 1 10 9 13 9 0
15 10 13 10 9 3 13 9 7 10 9 10 9 13 1 15
36 16 3 13 10 11 16 13 10 9 16 11 0 9 13 7 13 3 11 3 11 0 3 13 7 10 9 15 13 10 11 7 13 3 1 10 11
6 13 3 3 9 10 11
12 10 3 11 13 1 10 9 13 3 1 10 9
4 9 13 3 0
7 13 9 1 10 11 13 9
4 13 15 10 11
3 13 15 13
11 10 3 9 15 13 1 10 9 16 9 13
11 3 15 0 13 1 15 13 13 9 9 13
25 16 13 10 9 10 9 7 15 13 10 13 15 13 15 13 15 3 13 15 7 13 3 15 9 13
4 13 15 10 9
9 9 7 9 13 7 10 9 13 0
6 3 13 10 9 10 13
26 3 15 0 13 10 9 15 11 15 13 15 10 9 7 0 1 15 13 7 10 9 15 7 10 9 15
5 13 11 7 13 15
33 15 3 3 13 1 10 9 15 15 13 15 3 3 13 1 10 9 7 10 9 15 15 13 15 13 1 15 9 9 13 1 9 0
5 13 1 15 10 9
2 13 15
8 13 13 10 9 15 7 13 3
5 13 10 9 7 13
3 9 3 13
4 13 15 10 11
3 9 3 13
12 12 3 9 13 7 3 15 13 3 13 15 9
3 0 0 13
6 9 13 16 9 13 15
8 10 9 15 1 10 9 0 13
12 7 15 13 16 1 11 13 10 9 3 13 13
4 13 15 10 11
5 15 13 15 3 13
11 15 13 15 13 16 10 9 1 10 0 13
17 7 13 9 7 3 13 3 10 0 9 13 10 9 1 9 7 9
9 7 3 10 9 0 13 10 13 15
4 13 15 10 9
7 13 16 11 13 10 13 11
6 3 13 0 13 15 0
5 15 13 10 13 15
13 7 1 0 13 10 9 15 7 13 16 1 9 13
6 15 3 13 15 13 7
4 15 13 1 15
16 13 3 10 9 15 10 9 7 13 1 10 9 7 13 10 9
5 3 0 13 10 11
8 13 1 10 9 7 13 1 15
2 9 13
4 15 3 13 15
8 15 9 13 13 15 15 3 13
6 13 3 10 9 1 15
5 3 15 13 15 13
4 13 15 10 11
11 3 15 13 16 3 0 13 7 10 9 13
13 13 10 9 15 7 13 10 9 16 0 13 1 9
20 3 10 13 9 13 7 13 9 1 9 0 16 3 10 13 3 13 7 10 13
16 1 3 0 10 9 13 0 16 0 13 10 13 7 0 10 13
8 15 13 15 13 15 3 15 13
9 15 13 7 15 1 10 9 15 13
18 1 3 10 9 0 0 13 1 15 10 9 1 10 9 10 9 13 16
5 13 15 15 15 13
8 7 0 0 13 1 10 9 15
5 10 7 9 13 16
6 3 1 10 15 9 13
13 0 3 13 7 13 16 0 13 3 10 9 10 9
10 1 3 10 12 9 13 3 1 10 11
13 0 3 11 13 16 9 1 10 0 9 9 3 13
19 16 3 13 1 10 11 13 15 10 0 15 13 15 13 1 11 1 10 9
7 3 15 3 13 1 10 9
9 13 3 0 15 10 9 13 1 11
23 0 13 16 11 13 1 10 11 1 10 11 13 1 15 7 13 16 13 7 13 15 10 9
3 13 3 13
6 13 3 10 11 1 15
9 16 3 9 7 9 13 3 3 13
5 13 1 15 10 0
7 9 13 16 13 10 9 15
4 13 15 10 11
12 13 10 9 10 9 15 13 15 10 11 7 13
15 3 3 15 13 10 9 13 15 7 13 16 10 9 15 13
10 13 3 10 9 1 15 1 15 3 13
11 13 3 15 16 3 9 0 13 15 10 9
14 13 3 10 9 16 0 10 9 1 15 13 15 10 11
4 10 9 15 13
8 7 13 15 7 10 9 15 0
12 1 0 13 10 9 10 0 7 13 11 1 11
9 1 0 13 9 10 13 0 0 0
14 13 3 15 9 3 12 7 12 9 13 1 10 9 15
14 0 13 10 11 13 7 13 16 0 3 9 13 13 15
3 13 0 13
4 13 15 10 13
14 9 9 3 13 16 3 13 10 9 13 15 1 10 9
4 13 15 10 11
1 13
12 7 13 0 10 9 7 13 10 9 15 7 13
7 13 3 9 1 0 10 9
6 13 3 10 0 10 13
9 9 13 7 3 13 15 13 10 9
2 13 15
6 13 10 9 15 7 13
2 13 15
7 15 13 10 9 10 13 15
7 10 3 13 3 13 15 13
9 10 3 11 13 9 13 1 10 9
12 1 0 13 15 10 11 1 10 9 7 13 15
3 13 0 13
14 13 10 9 7 13 10 0 16 11 13 10 13 15 0
13 7 1 0 13 10 0 10 11 16 0 13 1 9
4 15 3 13 15
9 10 9 15 1 3 13 7 15 13
7 13 3 10 11 7 13 15
4 6 6 13 15
15 3 13 10 9 13 1 15 15 16 3 15 13 10 9 13
22 10 3 9 13 10 9 7 15 13 15 15 15 13 7 0 0 13 15 9 16 15 13
16 3 3 10 9 13 10 0 7 13 3 3 10 9 15 13 13
22 7 3 10 9 13 15 7 10 9 15 13 10 9 16 15 13 10 9 3 13 10 9
12 10 3 13 10 9 3 13 10 9 10 13 15
31 6 6 13 15 16 10 10 9 15 13 7 13 10 13 15 13 9 0 7 1 9 3 13 7 13 1 10 9 1 10 9
17 3 3 10 9 13 9 1 15 3 7 10 9 13 9 13 1 15
10 7 9 13 15 9 13 16 9 9 13
30 16 13 9 1 15 15 10 1 10 9 13 10 9 15 7 13 10 10 0 13 1 9 9 10 10 0 13 1 9 9
7 3 13 15 13 1 15 15
23 3 13 13 7 10 9 10 15 0 13 16 3 13 10 9 10 15 7 10 9 10 13 15
11 16 15 13 1 15 10 9 15 3 13 0
17 0 13 10 13 1 15 7 13 16 0 13 10 9 15 13 1 15
8 15 13 1 11 7 13 10 9
8 0 13 10 9 10 13 7 13
8 15 3 13 10 9 0 10 11
24 10 3 9 15 13 15 10 9 16 13 15 0 10 9 15 13 13 1 15 16 10 9 15 13
9 7 10 13 15 9 0 13 1 15
26 7 9 15 3 13 7 9 15 13 7 10 9 15 3 13 1 15 13 16 15 13 0 0 15 3 13
11 13 10 9 16 15 13 1 15 9 0 13
7 7 0 13 10 13 1 15
9 7 3 13 13 1 15 16 9 13
10 16 0 13 1 10 9 10 0 0 13
18 3 13 15 13 9 1 15 13 7 10 9 10 1 10 0 9 3 13
9 3 13 16 15 13 15 1 10 9
9 13 10 13 15 11 1 15 15 13
7 16 3 13 11 13 3 15
5 1 3 15 0 13
12 16 3 10 0 9 3 13 3 10 15 9 13
12 1 0 13 10 11 1 10 9 10 11 10 11
13 13 3 1 10 9 11 7 3 13 1 10 9 15
9 13 3 3 10 9 10 9 10 0
17 13 3 10 9 10 11 7 13 16 0 9 13 1 15 13 1 11
6 3 13 9 16 13 0
5 0 3 13 13 15
6 0 3 13 15 13 13
4 13 15 10 11
11 12 9 9 3 13 15 16 0 0 15 13
6 7 0 15 13 1 0
3 13 10 11
4 13 10 9 13
7 13 3 9 0 1 10 9
8 13 3 10 9 10 9 3 12
19 13 3 10 9 10 11 7 13 7 13 10 13 3 7 1 10 9 15 13
7 16 3 13 13 10 9 15
17 13 3 7 13 12 9 9 1 10 12 9 10 0 15 13 10 13
10 0 13 3 10 9 10 1 10 9 13
19 11 3 13 16 13 13 7 13 15 16 13 9 13 3 1 10 9 15 0
21 16 3 0 13 13 10 9 15 1 10 9 7 13 1 9 13 1 10 9 1 11
11 13 3 15 10 9 7 3 13 11 1 15
7 10 7 9 9 0 13 13
21 13 3 3 9 12 7 12 13 10 11 13 1 10 9 7 1 10 9 13 7 13
2 15 13
2 3 13
37 10 3 10 9 10 13 1 10 9 13 16 9 15 3 13 3 3 3 12 7 16 3 13 10 9 15 10 11 1 10 9 7 0 10 9 15 13
15 15 13 9 1 11 1 10 9 3 13 10 9 13 10 9
26 16 3 13 10 9 16 11 3 13 3 7 10 9 15 13 15 1 10 9 7 13 1 11 13 10 11
8 7 13 15 1 10 9 13 15
4 9 3 3 13
4 6 6 13 15
14 13 15 3 16 13 9 7 16 13 1 10 9 7 13
21 13 3 10 9 10 13 7 10 9 10 13 1 9 0 15 10 9 10 9 13 15
4 13 3 1 15
8 15 13 16 13 10 9 10 9
5 13 11 7 13 15
12 0 13 10 9 10 9 16 13 1 15 13 0
10 15 3 13 15 9 16 13 7 13 15
2 15 13
12 10 9 15 10 9 13 1 10 0 3 13 13
7 9 1 10 9 13 15 13
4 6 6 13 15
22 3 11 13 15 10 9 1 10 9 7 10 9 15 13 15 10 9 1 10 9 10 0
16 10 3 9 10 9 13 10 13 1 10 9 7 9 13 10 9
7 9 3 13 15 10 9 0
5 13 3 15 10 11
6 15 13 10 9 10 9
16 10 13 1 15 3 3 13 7 10 13 1 15 3 3 13 3
9 7 13 15 16 7 13 7 3 13
24 0 3 13 10 9 10 13 15 16 15 15 13 15 3 13 1 15 7 13 15 1 10 0 9
29 0 3 13 10 9 10 9 15 16 15 10 13 10 9 7 13 1 15 13 9 0 7 13 15 15 1 10 0 9
9 15 13 10 9 10 13 1 10 9
2 7 13
15 3 0 13 11 10 9 11 15 15 13 10 9 7 10 9
9 3 3 13 0 16 1 10 9 13
5 13 11 7 13 15
4 3 13 1 15
5 13 13 1 10 9
11 15 10 13 1 10 9 7 13 13 1 15
13 3 3 10 9 13 15 3 3 10 13 1 10 9
4 0 13 10 9
4 6 6 13 15
5 10 13 13 9 0
6 15 13 10 9 10 9
11 10 9 15 13 1 10 0 10 9 7 13
11 16 15 13 1 10 15 9 13 1 10 9
16 7 10 9 3 15 15 13 1 10 10 9 9 10 9 15 13
7 13 3 1 15 10 0 13
8 3 13 15 0 13 10 9 13
5 13 3 15 10 11
4 6 6 13 15
19 16 3 13 10 9 10 9 10 9 7 13 15 10 9 3 13 9 1 15
20 10 13 15 10 9 7 13 15 10 9 13 9 0 7 15 13 15 10 0 9
17 10 13 15 10 9 7 13 15 10 9 1 15 13 7 15 1 15
21 3 13 15 10 13 9 7 15 13 1 10 9 3 10 13 15 3 0 13 1 15
15 0 13 10 9 10 1 9 13 3 3 13 10 9 7 13
9 10 13 0 10 9 13 1 10 9
7 0 13 1 9 13 1 11
8 0 3 13 1 10 9 15 13
5 0 13 10 9 0
4 15 13 15 13
12 16 3 13 10 9 10 9 13 3 13 10 0
5 10 9 13 10 13
5 10 9 3 13 15
11 10 9 15 15 13 15 9 13 7 9 13
8 7 13 1 15 15 15 3 13
17 13 3 1 9 10 11 15 13 10 3 13 7 15 13 10 13 15
2 7 13
16 1 0 3 0 10 9 15 13 1 10 3 7 3 1 15 13
5 3 3 15 13 13
4 13 15 11 11
4 9 1 15 13
4 9 9 0 13
12 7 15 13 7 13 16 15 13 10 0 10 9
2 13 15
6 7 1 15 12 9 13
6 13 3 10 11 11 11
8 1 0 13 10 11 1 10 11
13 3 3 13 1 10 11 13 16 13 15 10 0 13
9 13 3 3 10 9 10 0 10 9
7 13 3 1 15 10 9 15
18 13 3 7 13 1 10 11 16 3 10 9 15 13 10 9 15 15 13
7 16 0 13 13 15 10 9
8 3 3 10 9 15 13 1 15
4 13 15 10 11
8 10 3 9 10 15 3 13 0
6 3 13 10 9 13 15
14 15 3 13 16 15 13 1 15 16 10 9 15 0 13
5 15 13 1 10 9
7 0 13 15 13 1 10 11
18 16 3 13 10 9 15 1 10 9 3 3 0 13 3 3 7 1 0
10 10 3 0 13 15 1 10 9 7 13
3 3 13 0
6 15 3 13 16 0 13
2 15 13
5 3 7 13 10 9
12 3 3 10 9 13 13 11 1 10 9 7 13
5 13 3 10 0 13
6 3 0 9 13 3 13
6 13 3 15 11 7 13
10 10 15 9 3 13 15 7 10 13 15
9 10 1 15 13 10 9 10 0 13
17 10 3 13 10 9 10 13 15 0 0 13 7 9 1 15 3 13
7 7 15 1 15 13 10 9
4 15 15 13 13
3 13 10 9
2 9 13
4 15 15 13 13
5 13 11 7 13 15
21 10 11 13 15 10 9 3 16 1 10 9 13 7 1 10 9 7 1 9 13 9
9 3 13 1 9 7 10 0 9 13
6 13 3 15 1 10 9
6 3 0 13 15 13 13
2 7 13
6 9 13 7 15 15 13
10 3 3 13 10 9 16 0 13 10 11
5 7 0 13 3 13
7 7 15 13 7 13 3 13
15 7 1 15 3 13 7 13 0 10 13 15 15 15 3 13
11 15 13 15 16 1 15 13 7 0 15 13
17 13 3 15 13 7 15 13 1 15 10 9 16 3 13 10 9 15
10 0 3 13 1 10 9 1 15 7 13
11 10 11 3 13 3 0 9 13 15 0 13
20 13 10 9 10 9 13 1 15 0 7 13 9 10 9 7 10 9 16 13 15
4 13 3 10 11
13 13 15 7 3 13 7 3 13 15 15 3 13 13
6 13 3 10 0 1 15
8 3 13 0 13 16 3 13 15
12 3 1 10 9 10 9 13 13 7 13 10 9
7 15 13 10 9 0 15 13
13 13 15 7 3 13 7 3 13 15 15 3 13 13
15 1 3 10 0 9 10 0 10 9 13 10 11 7 13 13
6 16 15 13 13 7 13
8 3 3 13 9 16 11 3 13
9 1 10 9 3 13 10 9 0 13
5 0 13 3 10 9
2 15 13
4 0 13 10 11
2 15 13
8 3 3 1 10 11 10 11 13
8 9 3 13 1 10 9 1 15
13 13 3 10 9 1 10 9 7 9 7 13 15 0
5 1 15 3 13 15
3 13 10 9
9 3 13 3 9 3 0 13 10 9
4 13 15 10 9
4 3 3 15 13
11 7 10 9 0 10 3 13 10 9 0 13
8 13 11 1 15 12 13 1 15
4 13 7 13 15
7 3 3 15 1 10 11 13
10 13 7 13 16 9 1 10 11 3 13
7 7 13 0 1 10 9 15
8 11 3 13 1 10 9 10 9
20 13 3 10 9 7 10 9 1 15 9 1 9 13 7 13 15 1 0 13 15
7 9 0 10 9 13 3 13
10 1 3 10 9 11 15 13 10 0 13
9 0 3 13 13 15 16 13 13 15
11 10 3 11 3 13 10 9 13 1 10 9
9 16 3 13 13 15 13 13 1 15
9 10 0 15 0 10 9 1 15 13
30 15 3 13 7 1 10 9 13 13 12 1 12 13 1 10 0 1 10 0 7 13 0 10 11 7 10 9 1 0 13
12 13 3 10 11 7 15 13 1 10 9 13 15
8 10 9 3 13 0 10 9 15
3 15 15 13
2 15 9
5 13 3 15 10 11
4 3 15 15 13
7 3 3 15 13 10 11 13
6 15 13 10 9 10 9
15 10 13 15 3 3 13 1 10 9 7 13 10 9 10 9
5 13 3 15 10 9
4 15 1 15 13
5 13 11 7 13 15
18 3 16 15 13 1 15 0 13 10 9 15 16 13 3 13 7 3 13
5 15 1 10 9 13
4 15 3 13 15
21 3 16 13 3 15 10 9 10 15 0 13 16 0 3 13 7 15 7 10 13 15
16 7 1 10 9 3 10 15 13 13 16 12 9 10 9 0 13
14 15 13 10 13 1 15 7 13 1 15 10 13 15 9
3 13 3 15
2 13 11
9 16 15 13 3 10 9 15 3 13
11 0 10 9 13 1 10 9 13 1 10 9
10 7 15 13 15 16 3 13 10 9 15
4 13 3 3 15
11 15 13 7 13 15 7 1 10 9 15 13
7 3 15 13 15 3 13 13
4 13 3 10 0
3 7 13 15
5 15 1 10 3 13
5 15 1 10 3 13
6 15 1 10 9 0 13
7 15 3 13 1 10 9 0
9 13 3 15 16 13 1 10 9 15
12 16 3 3 13 16 15 13 13 1 10 9 15
3 13 3 15
4 13 15 10 11
6 10 9 15 7 13 15
7 0 13 1 15 13 7 13
17 7 10 13 15 0 13 7 15 15 13 1 15 0 13 1 10 9
7 3 13 16 10 9 15 13
4 13 3 10 11
24 3 13 10 9 10 9 3 13 16 15 13 7 1 15 13 15 7 3 13 15 10 9 0 13
7 7 10 13 15 1 15 13
9 13 3 10 11 1 10 13 15 0
21 16 15 13 1 10 9 10 15 3 9 15 13 7 13 10 9 7 10 9 13 15
3 13 1 15
7 9 11 13 7 15 13 3
4 3 15 13 16
2 0 13
4 13 15 10 11
11 10 3 9 3 13 1 10 9 1 10 9
9 16 3 10 9 15 13 3 0 13
5 13 16 9 11 13
13 7 13 15 13 16 10 9 10 15 3 13 1 15
7 15 15 13 1 10 9 13
9 7 15 3 15 13 1 10 9 13
4 13 7 13 15
4 13 15 10 11
10 16 9 10 11 13 10 9 10 11 13
4 0 11 3 13
7 15 13 10 9 10 9 15
2 13 15
5 15 1 9 3 13
5 12 9 13 10 9
9 16 10 9 9 15 13 13 3 15
8 15 3 1 10 9 13 7 13
9 3 3 1 15 13 7 0 15 13
8 16 3 13 13 10 9 10 15
15 15 1 10 9 10 9 13 7 10 9 10 9 15 13 13
17 0 0 13 1 9 7 1 10 9 3 13 16 3 13 9 1 15
15 3 13 10 9 1 10 0 13 16 9 13 7 10 9 15
7 15 1 15 13 15 1 9
9 16 9 13 1 15 15 3 13 15
10 10 13 1 10 9 10 9 10 9 13
11 1 0 15 3 13 16 1 10 9 3 13
11 3 3 13 15 16 9 13 15 7 9 13
2 13 11
13 15 9 3 13 7 13 10 9 15 7 15 13 15
5 13 10 13 7 13
4 6 6 13 15
13 16 15 10 15 9 13 9 3 3 13 1 10 9
4 13 15 10 0
5 3 13 16 9 13
13 16 15 10 9 15 13 3 3 13 9 1 10 9
10 3 15 0 13 10 9 15 11 15 13
3 15 15 13
2 13 11
9 16 15 13 15 10 9 15 15 13
11 13 10 9 15 10 13 15 15 15 13 16
3 9 15 13
4 7 3 13 15
11 7 16 13 16 3 13 15 13 0 15 9
15 11 10 9 15 13 16 13 10 9 10 15 7 13 7 13
6 13 3 10 0 1 15
7 12 9 3 13 7 11 13
3 13 15 11
4 6 6 13 15
5 16 11 13 15 13
7 13 3 9 16 13 1 15
7 7 13 15 10 9 15 13
11 9 15 13 0 7 10 9 15 16 0 13
2 13 11
16 7 0 13 7 10 9 15 7 16 13 10 9 10 9 1 15
11 15 13 13 10 9 10 13 15 16 9 13
6 13 9 3 15 13 13
9 3 1 10 9 13 9 13 10 9
21 0 13 13 3 7 13 9 1 10 9 7 13 15 10 9 1 10 9 7 13 15
7 13 3 7 13 7 13 13
13 10 3 9 7 10 13 15 10 0 16 9 13 13
7 3 0 13 10 13 7 13
5 15 13 16 0 13
2 15 13
5 3 7 0 15 13
3 0 13 16
2 15 13
2 13 0
16 10 9 10 13 11 9 13 7 13 15 10 9 7 13 15 16
6 13 1 10 11 7 13
5 13 3 7 13 13
2 13 15
3 3 13 0
1 13
8 13 15 1 10 9 10 3 0
9 3 3 13 15 7 10 9 3 13
4 15 3 13 15
10 9 13 15 1 10 9 7 13 7 13
6 13 3 1 10 9 15
12 3 13 0 1 9 10 9 16 10 9 3 13
2 15 13
5 7 9 13 1 15
5 13 3 10 0 3
6 15 3 13 16 9 13
24 3 13 3 10 0 1 15 16 13 0 7 13 16 15 13 10 9 15 10 13 7 13 15 13
11 0 13 10 9 15 15 15 13 16 0 13
4 3 3 13 3
7 13 3 10 9 15 7 13
15 3 3 3 13 3 13 7 15 13 15 10 9 15 3 13
2 15 13
2 9 13
9 0 13 10 9 15 16 13 10 0
13 3 3 13 10 0 16 16 15 15 13 11 0 13
7 1 0 10 9 15 13 16
2 9 13
12 13 3 10 9 1 0 15 13 0 7 13 15
4 13 9 10 9
8 15 13 16 10 9 0 0 13
3 13 3 0
7 12 13 16 0 13 3 13
3 13 3 15
3 15 13 15
2 13 15
6 13 15 3 7 3 13
4 15 3 13 13
7 3 3 15 13 15 9 13
4 13 15 7 13
6 15 3 10 11 13 9
7 15 13 16 11 13 10 9
6 13 10 9 7 13 15
17 1 0 3 10 0 13 16 15 3 13 3 13 7 13 15 10 9
19 13 16 0 10 9 3 13 7 16 15 0 13 7 10 9 15 13 0 13
11 1 10 9 3 13 16 13 15 9 0 13
10 16 3 13 0 1 9 3 13 13 15
4 13 7 13 15
4 7 13 15 3
7 15 13 1 10 9 10 9
4 13 0 7 13
8 7 15 13 9 16 13 1 15
4 13 15 10 11
10 7 13 15 7 10 13 1 15 0 13
3 15 3 13
2 13 9
18 1 9 15 1 10 9 0 13 16 10 3 13 13 7 10 13 0 13
11 13 1 10 9 10 1 15 13 7 13 15
5 3 3 15 0 13
4 13 15 10 11
7 16 0 13 3 3 13 9
4 3 3 13 16
1 13
4 10 9 15 13
19 10 3 13 1 10 9 1 10 9 10 9 7 13 3 0 9 13 7 9
10 10 3 13 1 10 9 9 13 10 9
21 0 10 9 13 7 10 9 10 9 15 13 7 10 0 9 13 1 9 7 13 15
18 3 10 0 15 13 1 15 13 7 10 9 15 13 16 13 10 9 15
16 0 3 3 3 13 7 13 1 15 16 3 13 10 0 10 9
7 0 10 9 13 15 10 11
9 0 3 3 13 15 13 15 13 15
4 13 3 10 11
4 15 13 10 9
13 1 15 16 15 13 13 7 13 7 13 7 9 13
12 10 9 3 13 3 3 16 13 7 13 7 13
8 15 13 16 9 13 7 0 13
6 15 13 10 9 10 0
11 10 9 10 0 10 9 15 13 1 10 9
29 10 9 7 3 13 9 15 3 13 10 9 0 13 10 9 13 7 13 10 9 7 13 7 10 9 13 15 7 13
33 15 13 10 9 10 0 7 13 10 15 7 13 15 10 15 3 13 15 10 9 7 15 13 10 9 7 10 9 15 13 1 10 9
16 3 0 13 15 13 7 10 9 15 13 7 13 12 9 12 9
16 1 0 15 10 9 13 16 15 13 10 9 15 16 3 13 15
11 15 13 15 1 15 7 15 13 15 1 15
10 9 13 13 15 7 9 13 3 13 15
8 0 10 9 13 1 10 9 15
10 9 3 13 1 10 0 1 10 9 0
4 9 13 7 13
3 15 15 13
6 0 10 9 3 13 13
6 3 9 13 0 9 13
7 13 3 10 9 1 10 11
2 9 13
11 7 13 10 11 1 10 9 1 10 9 11
6 1 3 10 9 15 13
8 16 15 13 10 11 13 15 9
3 13 10 11
15 10 9 15 15 13 1 10 9 10 9 15 0 13 1 15
12 7 15 3 13 16 3 13 1 10 9 10 15
37 10 9 10 15 10 9 15 13 7 15 13 15 7 13 15 7 15 13 15 9 0 7 3 3 13 1 10 9 7 3 13 15 15 1 10 9 15
17 10 9 15 13 15 15 0 13 7 15 13 13 1 10 9 10 9
8 13 3 9 10 0 16 13 15
4 13 15 10 11
8 0 9 0 13 15 1 10 9
6 1 15 15 9 15 13
17 1 0 9 3 13 15 7 1 9 7 16 15 9 13 13 15 9
4 13 15 10 11
10 3 13 13 1 10 9 15 16 15 13
32 16 0 13 9 1 15 10 9 13 10 9 7 3 13 13 10 9 15 10 9 13 7 13 1 10 9 15 13 16 13 16 13
3 9 9 13
11 16 3 13 10 9 10 9 15 3 13 15
25 16 3 13 3 16 15 3 13 10 9 13 16 13 7 13 16 1 15 10 9 7 15 1 10 9
10 13 3 15 13 7 13 1 10 9 15
8 7 0 13 1 15 7 13 16
14 11 3 9 13 15 15 3 15 13 11 1 0 0 13
17 13 3 15 13 11 1 11 1 10 9 10 11 7 11 10 9 15
21 13 3 11 10 13 10 9 9 7 13 10 9 15 10 9 15 15 10 9 11 13
7 13 3 10 9 1 15 13
5 9 13 15 13 13
5 13 3 10 11 13
21 0 10 9 3 13 1 9 7 1 10 9 10 9 16 13 10 9 10 9 1 15
14 16 3 13 16 13 3 3 13 1 15 13 9 12 9
5 13 1 10 11 3
4 13 15 10 9
11 9 3 13 15 13 10 0 7 3 13 3
2 13 11
6 3 12 9 13 10 9
15 16 15 13 1 10 9 3 13 16 10 9 10 9 0 13
15 16 3 15 13 1 10 9 13 16 10 9 3 13 1 15
5 7 13 16 13 15
5 13 3 15 10 9
4 9 16 13 13
8 13 3 10 11 1 10 9 15
10 0 3 13 16 1 10 9 10 9 13
7 3 3 13 15 10 11 9
12 11 13 7 13 1 15 16 13 16 3 13 3
4 7 13 1 15
7 13 3 15 16 13 1 15
12 13 3 10 11 13 15 12 9 13 1 10 9
10 13 3 11 3 10 11 3 1 9 12
18 0 3 1 10 0 13 1 10 1 11 7 11 16 13 15 1 10 9
10 10 3 11 16 13 16 11 13 13 15
6 11 3 1 10 9 13
6 13 3 10 11 1 11
10 9 16 13 3 3 3 13 10 9 15
4 13 10 9 15
4 13 15 10 11
10 13 16 13 1 10 9 1 10 0 9
4 13 15 10 11
7 15 13 10 9 7 10 9
22 10 13 1 15 3 16 13 13 7 15 10 13 7 13 1 15 3 3 13 1 10 9
2 13 0
2 6 9
12 7 0 13 13 7 13 11 10 9 15 3 13
6 10 9 13 7 13 15
9 0 16 13 13 0 7 13 1 15
18 3 3 13 10 11 1 10 9 7 13 1 10 9 3 13 15 10 11
32 10 3 0 10 13 1 15 1 10 9 7 13 15 13 10 11 16 3 13 7 13 13 15 13 16 13 1 10 9 16 13 3
17 10 3 11 16 13 3 13 11 13 15 13 15 1 10 9 13 15
20 11 3 16 13 15 13 7 10 13 15 0 13 13 10 9 7 13 15 7 13
3 3 13 15
4 9 13 7 13
3 13 10 11
4 13 3 10 0
4 13 3 13 15
5 15 3 1 15 13
10 11 3 3 13 1 15 13 1 10 9
8 13 3 9 7 9 13 1 15
3 13 10 11
7 13 15 10 9 10 13 11
3 9 3 13
3 0 3 13
4 13 15 10 11
4 13 3 10 9
9 10 3 11 13 10 9 3 7 13
6 9 13 15 16 13 15
7 15 3 13 16 3 15 13
6 7 0 13 9 0 13
3 11 6 3
16 13 10 13 13 10 9 7 10 9 9 7 10 9 15 9 13
6 13 15 7 13 15 13
17 0 3 1 10 0 10 13 1 10 11 7 13 15 13 13 1 15
14 15 3 1 15 13 1 10 9 7 13 15 15 13 11
10 13 3 10 9 7 10 9 9 7 13
9 15 13 16 0 10 9 0 13 9
13 12 3 15 1 15 11 9 13 10 9 0 13 15
22 15 3 13 15 7 13 16 13 15 16 12 9 13 1 10 9 7 3 0 10 9 13
9 1 0 3 10 9 13 16 13 15
27 11 3 3 9 13 1 10 0 7 13 3 1 10 9 1 10 0 1 11 13 9 7 3 13 1 10 9
21 13 3 3 10 9 10 0 7 13 0 1 11 1 10 9 1 10 9 16 13 15
12 13 3 10 11 7 13 1 15 1 10 9 13
10 15 13 15 16 3 3 13 1 10 9
18 13 3 10 9 7 10 9 9 16 16 15 13 3 13 13 16 13 15
9 13 3 15 9 3 7 10 11 13
22 10 3 11 13 9 9 9 0 0 13 10 9 10 11 7 13 10 9 15 10 9 15
9 10 3 9 13 1 10 9 10 9
14 13 3 11 10 11 12 1 10 9 15 10 13 15 13
12 1 15 0 10 9 3 13 12 9 7 13 0
21 13 3 0 3 16 1 10 0 13 15 7 16 9 13 7 10 9 13 10 13 13
4 13 3 10 11
11 13 15 16 1 10 9 10 9 15 13 15
28 13 3 10 9 0 1 10 0 16 3 13 7 13 3 1 10 11 0 7 16 3 10 11 13 15 13 1 0
21 13 3 10 9 16 3 10 11 13 16 0 1 15 13 10 0 7 13 1 10 11
27 10 3 9 0 10 13 1 10 9 13 16 13 11 1 11 13 10 9 10 9 7 13 1 9 15 7 13
1 6
11 13 10 13 1 9 9 7 10 9 10 11
11 13 3 10 11 9 13 1 15 3 13 13
4 3 13 9 11
9 6 10 9 15 13 13 1 9 9
20 13 3 10 9 10 13 1 15 16 10 11 13 1 10 9 7 13 15 1 0
14 1 0 3 13 15 10 9 16 13 0 15 13 10 9
6 10 3 9 13 1 15
5 13 16 3 13 15
6 13 10 9 1 15 13
12 13 3 9 15 1 10 13 16 13 1 10 9
13 0 3 13 11 10 1 11 10 11 7 13 15 13
5 9 13 10 11 13
6 10 3 11 13 15 13
9 13 10 9 16 13 10 9 10 9
4 6 6 13 15
14 16 3 10 9 10 9 13 1 10 9 13 15 0 13
6 16 3 13 0 9 13
22 10 13 10 9 15 13 15 7 10 13 10 9 15 1 10 9 0 1 9 0 13 15
17 16 15 15 13 15 13 7 3 13 15 3 7 10 9 10 15 13
8 3 10 9 15 13 7 15 13
8 7 1 0 13 1 10 9 0
5 9 13 15 10 9
6 13 3 9 1 10 9
5 7 13 7 3 13
9 10 3 9 10 13 13 13 9 13
2 15 13
4 13 11 7 13
10 3 1 15 10 9 0 13 7 1 15
19 3 10 9 10 9 0 13 3 7 15 16 13 1 10 9 15 13 1 15
8 0 3 13 13 15 9 13 13
5 13 3 15 10 9
23 15 13 1 10 9 16 10 11 13 1 10 9 7 3 13 15 16 13 13 10 9 10 9
7 15 13 0 10 9 10 9
8 3 0 9 10 9 1 15 13
10 13 16 10 9 13 16 3 9 15 13
10 7 10 13 1 10 9 3 13 3 13
8 0 13 11 7 13 13 1 15
20 0 3 15 9 13 1 15 3 13 1 15 16 10 9 11 10 9 13 15 13
6 9 15 13 10 9 15
6 7 10 9 9 15 13
23 13 15 10 9 7 13 15 10 9 16 3 13 10 9 7 13 10 9 7 13 7 13 15
12 0 13 11 16 13 10 9 15 7 13 1 15
20 3 3 3 1 10 9 0 13 1 15 7 1 10 9 3 13 16 3 0 13
12 13 3 10 9 10 9 3 3 10 9 10 9
21 10 13 1 15 3 13 1 15 7 1 10 13 15 7 10 13 15 13 10 13 15
17 15 9 1 10 9 13 16 15 10 13 1 15 1 10 9 3 13
14 7 16 15 15 13 10 9 7 3 13 15 3 13 15
13 10 13 15 7 3 13 10 9 15 13 10 13 15
10 10 9 15 13 0 13 15 10 0 9
20 3 15 1 15 3 13 7 10 13 15 9 15 15 9 13 15 13 7 15 13
9 7 13 16 10 9 15 9 0 13
11 15 3 15 13 3 13 15 10 9 3 13
49 7 9 13 10 9 3 13 1 10 9 16 13 15 11 11 11 13 16 15 13 15 10 9 1 10 9 7 16 1 9 13 7 1 10 9 13 13 1 10 9 7 13 10 9 7 13 9 13 15
20 3 13 9 1 10 9 7 13 13 10 9 10 9 7 13 10 9 15 13 13
2 13 15
6 9 15 15 13 10 9
5 13 11 7 13 15
7 15 15 13 15 3 13 3
4 13 3 1 0
3 13 15 11
3 13 11 15
4 13 15 11 11
13 9 3 10 9 15 0 7 3 10 9 7 10 9
3 13 15 11
10 10 13 3 13 9 13 7 13 0 0
7 7 15 0 13 7 3 15
5 13 3 10 13 15
4 1 0 13 16
4 13 15 13 15
3 15 13 15
5 10 9 7 10 9
3 7 3 13
2 13 3
19 16 3 15 13 15 10 9 10 9 7 10 9 3 15 13 15 13 10 9
12 9 3 13 15 16 3 15 13 15 3 15 13
4 6 6 13 15
8 16 0 13 0 13 16 13 15
5 3 1 15 15 13
4 15 13 15 13
5 7 16 10 9 13
12 10 13 1 15 10 9 13 1 15 10 9 15
13 3 13 15 1 10 13 16 13 3 13 16 15 13
4 6 6 13 15
7 10 13 3 15 13 15 13
10 6 6 13 15 16 12 1 15 13 15
9 13 1 15 10 9 13 1 15 13
16 13 13 12 1 10 9 15 1 10 9 10 11 15 13 10 11
8 13 3 0 11 11 7 13 15
6 13 15 13 1 15 13
11 13 3 0 3 1 10 9 10 11 13 15
3 9 15 13
10 0 13 15 15 13 10 9 7 13 15
10 7 1 10 9 3 13 1 0 10 11
4 13 3 15 11
4 15 13 13 3
10 0 3 15 13 10 13 1 15 13 15
25 15 3 13 16 10 9 13 11 16 13 15 11 13 15 9 13 1 10 9 7 10 0 16 15 13
7 13 3 10 9 0 13 3
5 16 3 13 13 11
12 3 13 10 9 10 9 7 10 9 13 1 15
6 9 3 0 1 15 13
19 13 15 7 3 13 10 0 16 3 15 13 15 3 13 13 3 15 13 3
7 9 0 13 15 16 13 15
8 3 13 15 16 3 15 13 15
13 1 0 13 15 16 15 9 13 16 9 13 1 15
3 9 3 13
2 13 11
8 3 15 13 3 13 15 3 13
3 13 15 11
8 9 1 15 3 13 15 13 3
6 10 9 15 1 15 13
2 13 11
4 6 6 13 15
9 3 3 9 13 16 15 13 15 3
5 3 13 15 10 9
8 13 1 10 9 7 1 15 13
11 16 3 3 13 3 15 16 13 13 9 15
21 7 16 13 7 13 9 15 3 13 7 13 15 1 15 16 3 13 15 3 15 13
7 7 3 15 13 13 10 9
10 9 3 13 3 13 7 3 13 10 9
3 13 15 11
10 15 13 10 9 7 10 9 7 10 9
9 15 13 1 10 9 3 3 1 15
8 16 13 15 3 10 9 15 13
3 13 15 11
8 9 13 15 10 9 7 13 15
10 0 9 1 15 13 7 3 13 15 11
6 10 13 15 13 10 9
3 3 15 13
4 13 15 10 9
13 3 13 16 15 1 10 9 7 10 9 1 15 13
10 10 9 15 15 13 15 1 15 3 13
12 13 15 16 15 1 10 9 7 10 9 1 15
4 6 6 13 15
16 10 13 1 15 10 9 15 15 13 3 0 13 7 0 0 13
6 3 15 1 10 9 13
17 7 15 3 13 1 10 9 15 0 13 16 13 10 9 1 10 9
10 16 15 13 15 1 10 9 15 15 13
8 16 13 15 10 9 10 15 13
34 7 15 13 10 9 7 0 9 13 15 16 1 15 13 1 10 9 10 9 10 9 15 10 9 3 13 13 16 3 13 15 7 13 15
3 13 1 15
8 3 0 7 10 9 15 3 13
10 15 3 13 15 16 15 13 7 15 13
20 1 0 10 9 13 15 16 15 1 10 9 15 7 15 1 15 7 15 1 15
13 10 13 10 9 15 7 13 15 0 13 10 13 15
17 10 3 13 15 13 1 10 9 15 7 15 13 15 7 13 15 15
6 13 15 11 3 10 11
13 9 7 15 13 16 15 13 13 15 7 3 10 9
23 16 15 13 15 10 9 15 13 7 10 9 15 13 15 7 1 15 13 7 9 1 15 13
9 10 3 13 15 10 9 15 3 13
13 7 10 9 15 13 3 13 15 7 10 13 15 9
6 0 13 15 1 15 13
26 10 3 9 10 9 10 0 15 13 10 9 1 10 9 15 0 15 13 15 7 13 15 15 15 13 15
3 9 13 15
5 9 10 15 13 15
8 3 3 10 9 13 15 13 15
5 13 7 13 1 15
16 16 13 15 13 3 16 13 1 10 9 16 10 9 0 15 13
10 7 3 13 15 16 13 16 3 13 13
5 3 0 13 1 15
12 13 3 10 10 9 9 7 1 15 3 13 15
17 7 3 13 10 9 16 13 10 9 7 3 13 15 10 9 3 13
1 13
13 15 13 10 9 10 0 7 10 9 15 10 9 13
10 3 15 0 13 1 10 9 15 13 15
7 13 1 15 7 15 1 15
23 3 10 9 3 13 9 13 1 15 16 3 13 1 10 9 3 3 15 16 3 1 15 13
4 15 13 10 9
3 15 10 9
19 10 13 1 15 7 15 1 15 0 13 9 0 16 1 15 3 13 13 15
18 16 13 1 15 7 10 9 15 1 15 13 15 3 13 13 7 13 15
14 1 0 13 10 9 15 16 9 0 13 7 13 15 9
6 13 1 10 9 10 15
25 16 10 9 15 13 13 1 10 9 15 3 3 15 10 9 15 10 9 13 7 13 15 1 10 9
16 0 13 15 16 10 9 10 15 1 15 13 7 10 9 15 13
12 0 13 10 9 10 15 16 13 15 3 13 15
14 0 0 9 15 13 16 10 9 15 13 1 10 9 15
14 3 13 15 9 16 10 9 3 13 15 13 15 10 9
14 15 3 13 9 16 15 15 13 1 10 9 15 13 15
34 3 15 15 13 7 15 13 15 7 13 15 16 15 13 7 9 13 7 10 9 15 13 16 15 3 13 10 9 1 10 9 15 13 15
10 16 10 9 15 13 13 16 15 0 13
11 16 1 10 9 13 10 9 3 10 0 13
20 16 3 1 10 9 3 13 7 15 13 15 1 10 9 1 0 13 15 10 9
7 13 10 9 15 15 13 15
6 16 15 13 3 15 13
9 16 10 9 15 13 7 10 15 13
16 7 0 15 13 1 15 1 10 9 15 16 3 13 10 13 15
9 16 3 13 7 13 15 9 3 13
8 10 15 13 3 10 9 15 13
14 16 10 9 3 13 1 15 15 15 0 13 9 3 13
12 3 3 7 13 7 13 7 15 7 10 9 15
3 13 15 3
24 3 13 10 9 15 15 13 15 1 10 9 10 9 10 9 15 1 10 9 13 0 13 1 15
10 3 15 3 13 16 1 9 1 15 13
6 0 13 15 16 3 13
3 0 13 15
10 7 0 13 16 3 13 10 9 7 15
15 7 0 13 15 16 3 13 10 9 13 15 16 15 13 15
13 3 3 13 1 10 13 15 7 15 1 15 13 15
2 3 13
11 7 16 0 13 15 10 9 13 15 10 9
6 7 15 10 9 13 15
5 13 15 16 15 13
10 16 3 3 13 10 9 3 13 1 15
44 7 13 0 13 10 9 1 9 7 1 9 7 1 9 1 9 3 16 3 13 1 15 1 9 3 16 1 10 9 13 7 3 13 15 1 3 9 16 10 9 10 9 0 13
14 3 3 13 0 10 9 10 9 13 15 1 10 9 15
14 3 3 13 1 15 7 15 13 13 7 10 13 13 15
11 0 15 13 16 1 10 15 13 7 13 15
7 15 15 13 10 9 15 13
11 1 0 13 16 1 10 15 13 7 13 15
11 0 7 3 13 15 7 3 0 7 13 15
8 13 3 1 10 9 15 1 15
2 13 3
7 0 15 13 15 13 10 0
4 3 13 15 13
9 13 11 16 13 15 13 7 13 15
7 1 0 13 1 15 16 13
11 0 7 3 13 15 7 3 0 7 13 15
9 6 6 13 15 16 13 7 13 15
4 10 3 9 13
11 10 9 3 13 9 13 16 13 10 9 15
18 3 3 13 10 9 3 13 10 9 1 10 9 16 13 9 1 10 9
7 3 15 3 3 3 9 13
17 3 3 13 15 7 13 15 10 9 7 10 9 15 15 13 1 15
9 7 1 0 10 9 15 3 13 15
4 6 6 13 15
11 16 15 13 10 9 13 15 1 10 9 15
9 1 3 3 13 15 1 10 9 15
15 13 9 3 3 1 9 13 15 7 9 1 10 9 13 15
20 1 0 10 9 1 10 9 15 13 7 3 13 15 16 15 13 10 9 1 15
18 0 3 10 9 13 15 16 15 15 13 7 13 16 15 1 10 9 13
9 13 1 10 9 7 13 1 10 9
9 3 13 10 9 7 13 1 10 9
4 13 10 9 15
9 13 3 1 9 13 7 9 15 13
7 1 0 13 16 1 9 13
2 3 13
15 6 13 9 7 13 16 13 0 1 10 0 7 15 0 13
10 7 3 13 0 16 10 9 1 15 13
8 0 13 15 16 1 15 9 13
5 1 10 9 9 13
2 7 13
12 0 13 11 7 13 10 9 15 1 10 9 13
4 9 13 10 9
18 0 3 13 10 0 9 16 13 15 10 0 0 9 7 15 13 11 11
14 15 15 13 1 10 9 10 9 13 15 13 15 16 13
19 7 3 13 15 15 9 1 15 10 9 15 13 1 10 10 9 13 1 15
12 13 15 10 9 10 9 15 13 15 1 10 9
11 15 13 7 15 15 13 7 10 9 15 13
24 3 10 9 15 13 15 13 15 7 15 13 7 13 3 16 1 15 13 7 13 16 15 15 13
4 15 1 15 13
13 3 1 10 9 13 7 1 15 13 15 16 15 13
17 7 3 13 1 10 9 7 15 1 10 9 13 7 15 1 15 13
16 9 0 13 15 1 10 9 15 15 13 15 16 13 12 3 15
31 16 13 1 15 15 13 15 1 10 9 15 15 13 15 7 13 7 15 1 15 13 3 3 10 9 10 9 16 10 9 13
20 3 3 1 15 13 7 0 13 1 10 9 16 13 10 9 10 15 13 1 15
15 3 13 16 13 15 1 10 9 7 16 13 15 1 10 0
12 1 10 9 3 13 3 15 3 13 1 10 9
5 13 15 1 10 9
6 10 9 10 15 9 13
12 7 1 15 13 15 16 13 3 15 13 1 9
44 3 1 0 3 13 0 7 3 1 10 13 1 10 9 15 1 15 16 15 12 13 3 15 9 1 15 7 15 1 15 16 3 15 1 15 13 16 10 9 13 16 15 15 13
15 7 15 10 9 15 13 15 13 15 16 13 12 3 15 12
29 9 15 13 15 13 16 3 13 15 3 0 13 1 15 16 13 10 9 10 15 15 13 15 16 13 15 1 9 9
8 9 0 7 10 9 15 3 13
11 15 3 15 13 7 0 13 16 15 15 13
21 7 13 15 10 9 15 7 13 16 10 9 15 13 15 1 15 13 7 15 1 15
24 0 13 11 13 1 10 9 15 1 10 9 10 11 3 13 9 1 15 13 15 7 10 9 15
23 10 3 11 13 10 9 7 1 10 9 7 1 10 9 9 13 3 1 9 7 9 7 9
12 11 3 13 15 10 13 1 15 13 7 13 15
2 13 15
3 11 10 0
3 13 15 11
2 15 13
9 13 3 3 11 10 13 15 1 15
13 16 3 13 15 15 13 13 1 10 3 7 13 3
2 15 13
3 11 10 0
2 13 11
5 13 15 16 15 13
7 16 3 15 13 13 0 13
7 16 13 10 9 15 13 16
8 15 13 15 3 13 1 15 15
20 11 3 11 13 9 13 15 7 13 10 10 9 9 7 13 15 10 9 10 0
6 13 10 9 1 10 9
11 10 9 15 13 15 10 9 3 3 13 15
22 10 3 9 7 10 9 7 10 9 10 0 13 10 11 7 13 15 7 13 1 11 0
11 13 3 9 10 11 15 13 9 10 9 0
15 13 3 11 10 13 10 0 16 13 12 9 13 1 10 9
9 13 3 10 11 11 11 7 0 9
17 10 3 9 0 13 0 10 9 7 13 10 11 1 10 9 10 9
8 10 3 11 13 1 10 9 3
8 13 3 10 11 10 9 10 9
10 3 3 15 1 10 9 13 10 9 0
2 13 0
2 3 13
14 13 3 10 9 7 10 9 9 13 16 9 13 7 13
10 13 3 3 10 11 1 15 13 7 13
15 10 3 9 13 10 11 1 10 9 15 7 1 10 9 15
3 13 15 11
3 15 15 13
6 13 10 13 15 13 15
6 13 0 13 15 13 15
13 0 3 15 13 12 13 10 9 13 9 10 11 13
4 3 13 10 9
3 13 15 11
7 16 3 13 13 1 10 0
10 13 3 15 10 11 13 1 11 10 9
3 13 3 15
8 3 3 15 1 10 9 15 13
4 13 0 7 13
2 3 13
14 13 12 1 10 9 10 9 0 13 15 13 11 10 9
9 3 15 15 13 1 10 9 1 15
4 7 3 9 13
10 13 3 10 11 1 10 11 1 10 9
14 7 0 3 13 1 10 9 16 3 13 7 13 10 9
9 13 3 10 11 3 1 15 7 13
6 15 9 13 10 9 0
4 13 7 13 15
11 16 3 13 0 0 13 3 3 15 13 15
9 13 15 15 7 1 10 9 15 13
5 13 3 15 10 0
5 15 3 13 13 15
15 13 3 1 10 9 3 10 11 7 13 10 11 7 13 15
6 15 13 10 9 10 0
2 13 11
11 1 15 15 0 13 7 15 15 13 1 15
4 3 15 0 13
10 10 9 10 15 7 10 9 13 15 15
2 15 13
2 13 11
21 16 1 10 9 0 13 10 9 10 15 10 9 3 10 15 13 16 3 13 10 0
9 3 3 10 9 10 15 3 13 3
5 13 3 15 10 11
3 13 10 11
5 15 13 16 9 13
15 15 1 0 13 7 1 0 13 1 10 9 16 13 10 9
10 15 10 13 1 10 9 13 15 10 9
4 13 15 10 11
11 7 0 13 3 13 1 10 0 7 13 15
6 15 15 13 1 15 9
8 13 3 13 15 10 9 10 0
4 13 3 3 13
5 3 0 7 10 11
5 13 3 10 11 9
9 3 3 13 10 11 10 11 7 13
22 7 10 9 13 9 1 9 13 15 10 9 7 9 0 13 15 7 13 1 15 7 13
4 7 13 15 9
11 13 13 15 15 3 16 13 16 9 3 13
13 13 3 10 11 3 13 10 0 9 7 10 0 9
3 7 13 15
3 6 10 9
10 16 3 13 15 10 9 7 10 9 13
1 13
1 13
7 15 3 3 13 1 15 9
3 13 10 0
14 15 9 13 7 1 10 9 13 13 16 9 9 15 13
20 16 3 13 10 11 0 10 9 3 13 7 13 1 10 9 3 7 13 10 11
3 3 13 15
7 10 3 11 9 3 13 15
4 13 15 10 11
3 15 3 13
2 13 11
12 3 13 9 1 15 15 16 3 13 13 15 3
9 1 0 10 13 15 15 0 9 13
7 1 0 10 11 13 13 15
5 10 3 0 13 13
8 16 0 13 3 13 9 10 9
8 15 10 9 15 13 13 10 9
22 10 3 11 13 10 9 0 13 3 10 11 7 13 1 9 1 9 13 0 3 3 11
4 7 13 10 0
4 13 10 9 15
3 13 3 0
1 13
1 13
2 13 15
4 13 15 10 11
3 13 10 9
7 3 3 13 15 15 16 13
34 13 3 10 11 7 13 15 10 9 13 1 10 13 9 9 15 13 3 11 3 15 13 7 1 15 15 12 3 7 3 0 3 10 11
11 13 3 7 9 10 11 7 13 1 10 9
3 13 3 13
7 11 10 0 10 9 10 0
19 0 3 10 9 0 13 10 0 16 3 13 10 9 10 9 3 13 10 11
8 13 3 10 11 10 9 10 0
10 3 13 10 9 10 0 7 16 0 13
3 13 10 11
3 15 13 13
21 10 3 9 16 13 10 11 13 10 9 15 7 13 12 9 15 9 9 7 10 9
11 13 3 10 9 0 1 10 3 0 1 0
4 13 3 1 15
4 16 10 9 13
12 13 10 9 15 15 7 1 10 9 15 13 9
6 10 3 3 9 0 13
14 11 3 13 10 9 7 10 9 13 15 13 13 10 9
5 9 13 10 9 15
4 3 13 10 9
4 13 10 9 15
14 1 0 13 10 11 16 3 15 13 16 13 10 9 13
1 13
4 9 13 9 0
10 9 3 0 9 9 13 13 15 10 9
1 13
7 7 13 10 9 13 10 9
35 10 3 0 16 9 13 16 3 13 1 10 9 10 9 1 10 9 13 3 0 10 9 0 10 9 13 10 11 16 13 15 10 9 7 13
30 1 3 10 11 13 16 13 3 15 13 3 13 15 10 9 7 12 10 9 9 15 10 9 13 7 13 3 9 7 9
20 7 10 13 13 7 0 15 13 10 9 7 0 13 16 0 13 16 7 15 13
7 13 3 0 16 10 9 13
4 9 3 13 15
5 7 3 0 9 13
27 1 3 0 13 10 11 11 10 1 11 13 9 10 11 13 3 1 10 9 10 0 16 13 10 9 10 11
4 7 13 10 11
19 13 3 7 11 10 13 1 15 9 10 0 13 9 9 7 9 3 9 12
19 13 3 10 9 10 11 7 13 15 9 1 10 9 3 9 13 10 0 13
19 13 3 1 10 9 3 13 9 7 1 10 9 9 0 1 15 3 15 13
15 3 3 1 10 9 10 0 16 3 13 10 9 13 10 11
24 10 3 12 10 9 11 10 9 13 3 9 3 13 1 10 9 7 13 10 9 13 1 10 9
19 13 3 7 13 1 11 11 7 1 10 0 9 15 13 10 11 7 13 15
13 13 3 10 11 7 10 0 9 7 13 1 10 9
20 7 10 0 9 13 3 10 11 7 13 0 1 10 9 7 13 13 13 10 9
3 3 3 13
36 13 3 11 11 13 15 7 13 1 10 9 7 13 10 9 13 7 10 9 15 13 1 10 9 15 3 1 10 9 13 7 3 13 1 12 9
17 3 3 13 3 10 0 9 10 13 0 1 10 9 7 13 7 13
11 3 3 13 10 9 16 13 15 1 0 13
7 13 3 3 1 15 10 9
8 11 3 13 1 10 9 3 13
3 9 15 13
3 13 15 16
10 13 10 9 15 7 3 13 3 13 15
17 0 13 13 1 10 3 7 13 10 11 13 7 3 13 16 11 13
3 13 15 11
3 9 15 13
2 15 13
8 0 13 16 10 9 13 13 15
3 13 15 11
1 11
5 13 0 13 15 3
1 9
3 15 13 9
3 13 15 11
3 3 15 13
6 3 3 13 1 10 9
15 13 11 10 9 13 10 9 16 13 10 9 7 0 13 15
33 13 3 0 10 9 0 10 12 9 7 10 9 13 3 13 10 9 1 10 9 10 0 13 10 11 7 13 1 10 0 7 13 15
2 9 15
10 7 0 13 13 10 9 7 10 9 15
7 13 3 10 9 13 10 9
4 13 3 15 3
2 9 15
7 7 0 13 13 7 13 15
7 16 15 13 10 9 13 15
4 16 15 13 13
16 11 3 12 1 10 12 10 13 11 3 13 1 15 16 13 11
6 13 3 15 10 0 9
3 13 10 9
4 15 3 13 15
14 7 1 9 12 3 13 3 10 9 15 7 11 1 15
13 13 10 11 10 9 13 7 13 1 10 0 7 13
4 3 13 10 11
27 13 10 9 15 3 7 13 10 9 15 7 13 10 9 15 7 13 1 10 9 15 7 3 13 0 7 0
5 13 11 7 13 15
7 10 9 15 7 10 9 15
4 13 15 10 11
6 0 10 3 13 7 13
20 0 3 3 7 0 9 13 10 11 1 10 9 15 3 13 13 1 10 9 0
23 0 3 13 16 13 16 11 13 10 11 10 9 10 9 7 16 13 9 13 1 10 9 15
3 13 3 3
27 13 3 11 11 7 11 10 13 11 7 11 10 1 11 10 11 7 10 10 11 7 15 1 10 9 15 12
4 13 15 11 11
2 13 13
5 13 3 15 1 15
13 13 7 13 1 10 9 7 1 0 10 9 13 15
9 9 3 3 13 13 11 1 10 9
8 3 3 13 10 9 16 11 13
5 9 3 15 9 13
2 13 15
1 3
11 13 1 10 0 9 10 9 10 9 7 13
12 13 3 7 3 15 13 13 1 10 9 10 9
11 13 3 10 9 0 15 13 10 11 10 11
3 10 9 13
20 11 3 11 13 16 10 9 13 10 9 13 13 3 0 7 13 15 1 10 9
17 3 3 13 3 1 10 9 7 3 1 9 12 13 10 9 10 9
14 16 3 13 1 10 9 13 9 13 7 9 13 7 9
7 13 1 10 9 15 13 3
14 13 11 11 7 13 10 9 1 10 9 0 9 0 12
7 3 0 13 3 13 10 9
4 13 15 10 11
2 6 13
15 15 3 13 10 9 13 15 15 15 13 13 16 10 9 13
10 0 3 0 13 11 10 9 13 1 0
6 11 11 13 15 0 0
2 13 15
7 6 9 15 13 16 13 15
2 13 15
4 13 10 9 15
4 13 15 3 0
4 11 11 13 15
2 13 15
4 13 10 9 15
4 13 15 10 0
4 11 11 13 15
8 13 10 11 16 13 15 10 0
2 13 15
3 7 13 15
4 9 15 15 13
2 13 15
4 13 10 9 15
4 6 6 13 15
9 16 13 0 13 15 7 13 3 13
16 3 3 13 13 10 9 15 7 15 15 13 7 13 3 3 13
9 0 3 13 13 15 9 13 10 9
5 7 0 13 13 15
2 13 15
8 0 3 13 10 11 13 10 11
4 9 0 3 15
4 13 15 10 11
9 16 15 13 13 16 13 15 1 15
3 15 15 13
14 13 3 0 10 9 1 10 9 16 10 9 0 3 13
10 7 3 13 15 10 11 16 3 13 7
19 0 13 10 9 10 13 1 0 7 13 0 7 13 16 0 15 10 9 13
25 15 7 13 15 13 1 10 13 15 1 0 9 1 9 12 13 15 7 13 10 1 10 9 10 9
17 7 13 13 15 1 11 3 13 7 13 10 9 10 9 15 13 15
5 3 11 3 13 9
11 15 3 1 9 13 0 3 1 0 0 9
7 15 3 3 13 13 15 13
11 9 3 1 10 9 0 13 10 9 10 11
43 3 15 13 13 9 7 9 15 10 9 13 1 10 0 9 7 13 9 13 10 0 9 1 15 7 13 15 9 1 7 11 7 1 15 10 11 7 11 7 1 0 10 9
14 7 0 13 13 15 13 7 9 13 15 1 10 9 15
8 9 0 15 13 13 1 10 9
20 0 10 11 10 13 1 15 1 10 9 3 13 15 9 13 15 13 1 10 9
16 3 13 1 11 1 9 10 13 9 15 13 1 11 9 13 9
34 7 16 13 1 10 9 13 3 13 13 10 7 11 7 11 7 11 7 11 11 7 11 11 7 11 11 11 7 11 10 9 7 11 11
19 0 15 13 13 3 10 9 1 9 7 11 10 9 10 11 7 10 9 15
9 13 7 9 9 1 10 15 3 12
23 9 9 13 13 10 9 15 13 10 9 10 0 1 9 11 1 11 10 13 9 10 13 11
12 3 13 13 1 15 7 13 10 9 10 9 0
22 15 7 0 13 15 10 13 11 16 13 10 9 0 10 0 9 15 11 0 13 9 9
5 13 3 1 9 9
18 13 10 9 15 0 7 3 13 10 13 1 15 7 10 9 15 13 0
39 13 3 10 13 15 9 1 15 9 15 13 7 13 1 15 10 9 11 13 1 10 9 11 1 10 9 15 13 1 15 9 10 9 15 1 15 13 12 0
3 7 13 13
30 15 9 9 15 13 15 13 1 0 10 12 12 13 10 9 10 9 0 7 9 1 15 13 11 13 1 10 9 10 0
16 7 13 9 15 7 13 10 9 1 11 7 13 1 10 12 9
14 7 1 10 13 10 9 10 9 13 15 3 1 10 15
29 7 13 15 13 9 3 9 7 13 1 12 15 15 7 13 15 9 0 7 13 13 0 9 3 10 9 13 13 15
15 13 3 1 11 13 0 9 0 1 15 9 10 1 10 9
19 13 3 10 9 0 13 10 9 7 13 16 13 12 15 10 0 9 13 15
8 3 6 0 0 13 10 13 0
12 7 3 15 13 15 10 0 9 15 1 15 13
52 9 7 9 7 9 7 10 13 10 11 11 7 7 11 11 7 10 11 11 7 7 11 11 7 10 9 10 11 10 1 11 7 10 13 0 0 7 7 9 9 7 9 13 13 15 10 15 9 10 0 10 9
9 13 3 15 7 13 0 1 0 13
4 15 13 0 13
14 13 3 10 9 1 10 12 13 10 9 15 7 13 15
16 9 0 7 10 13 11 15 0 15 0 13 7 13 10 9 15
6 7 13 1 10 0 9
3 13 10 9
29 13 1 10 9 15 1 15 9 7 13 10 9 15 7 10 9 15 7 10 9 15 9 13 7 10 0 15 9 13
21 3 1 10 9 15 7 1 10 9 15 1 10 9 0 13 1 10 9 15 7 13
19 7 13 9 1 10 9 3 7 9 1 10 9 3 9 7 9 7 9 9
10 10 9 13 1 9 7 10 9 1 9
2 7 13
6 9 9 13 10 9 0
58 11 10 0 9 13 1 10 9 1 15 9 7 9 7 9 15 13 1 15 10 9 1 0 15 3 0 13 0 10 13 9 7 9 10 9 0 1 9 0 13 13 15 10 9 13 13 10 9 10 9 16 3 13 0 13 15 1 15
5 11 3 13 1 15
15 13 10 9 15 1 15 3 16 1 0 15 13 16 3 13
20 1 0 13 15 10 9 7 13 10 9 15 3 3 3 10 9 15 13 1 9
15 3 3 13 10 9 15 1 11 7 13 10 0 15 13 9
4 13 15 9 9
39 9 3 13 7 13 16 9 13 15 10 9 1 9 10 9 15 13 1 10 9 15 13 13 1 10 9 10 11 16 7 13 1 11 7 10 9 15 13 9
11 0 10 11 13 10 9 15 15 15 13 9
25 10 0 3 10 9 13 10 7 9 10 9 10 0 13 1 10 9 13 0 0 15 7 13 7 13
7 3 3 11 13 1 10 9
3 13 3 15
5 13 9 10 9 15
14 13 1 0 15 16 3 13 10 0 15 9 10 9 15
21 3 3 13 15 9 11 16 7 9 15 7 11 13 10 9 0 10 11 15 15 13
4 15 13 9 9
27 9 3 1 15 13 13 7 13 0 15 1 10 9 11 11 1 9 10 9 15 7 13 10 9 10 0 9
21 15 3 13 10 9 7 10 9 15 7 15 10 1 3 15 3 13 9 10 9 15
9 0 3 9 0 13 7 13 15 13
7 13 1 10 9 10 0 0
17 10 3 3 13 10 9 15 13 7 13 1 10 9 0 9 3 12
17 13 3 13 10 9 10 9 7 10 9 10 9 10 9 7 10 9
5 13 3 15 9 9
30 1 9 7 13 3 1 10 9 13 7 1 9 9 13 9 1 9 7 9 9 13 10 9 7 13 9 1 0 10 9
11 10 3 9 13 10 13 1 9 1 10 15
15 11 3 7 11 13 1 10 9 1 10 9 10 9 10 0
31 3 15 9 0 1 9 9 15 13 13 15 13 1 9 1 10 9 10 9 10 13 0 10 13 9 1 10 13 1 10 9
13 15 13 11 7 11 13 13 1 10 9 13 9 13
9 13 3 11 1 15 1 10 11 13
3 13 1 15
3 13 3 11
6 15 3 13 0 15 13
8 1 10 9 11 11 10 0 13
8 3 13 15 10 0 9 13 15
28 3 3 13 10 9 15 7 10 9 7 13 13 7 13 7 13 1 15 1 10 9 13 7 13 7 13 10 9
37 3 13 15 10 9 15 13 7 13 10 9 13 3 15 16 15 13 10 1 10 9 13 1 10 0 9 10 9 7 13 9 7 9 1 10 13 15
21 13 3 15 10 11 7 10 11 13 15 10 9 1 15 1 10 9 10 13 11 0
19 9 9 15 13 1 0 7 15 15 13 3 0 9 7 9 13 10 13 15
33 10 9 11 7 10 9 11 7 10 9 11 10 9 10 9 15 13 10 9 15 11 15 15 3 13 7 13 1 9 11 13 0 13
30 3 1 10 9 10 9 15 0 15 13 7 13 13 10 9 15 7 10 9 10 1 15 13 15 10 9 0 1 15 15
13 3 3 9 13 16 1 9 13 3 3 10 13 15
16 10 3 9 15 13 1 9 15 10 9 13 10 11 15 13 3
47 13 3 7 13 1 10 13 15 10 9 16 3 13 9 9 1 9 10 9 7 13 10 13 15 11 11 15 13 9 3 13 1 9 9 15 15 13 10 9 1 9 10 0 1 9 15 9
4 9 3 13 16
9 15 13 1 15 15 3 13 1 15
2 13 3
13 15 9 15 3 3 13 10 9 0 13 1 10 9
20 15 13 10 9 10 9 7 10 9 15 13 10 9 1 10 9 15 13 1 11
11 7 1 10 9 15 13 15 10 9 10 9
20 15 0 13 10 9 10 9 15 13 15 13 15 1 10 13 15 1 10 9 15
47 13 3 15 1 10 9 13 15 10 9 7 10 9 10 9 7 10 9 13 1 10 13 15 10 9 7 13 1 10 11 10 9 10 1 0 7 13 15 10 9 7 13 1 9 1 10 3
14 0 3 10 13 10 9 13 7 13 9 10 9 9 12
40 13 3 1 10 3 13 15 10 9 7 10 0 7 10 9 1 11 7 11 10 9 7 11 7 11 7 11 7 15 13 1 9 0 7 13 15 1 10 0 13
10 1 15 9 7 1 15 9 0 13 15
8 3 9 13 9 0 13 1 15
15 0 13 10 9 10 13 1 15 10 9 10 13 1 9 9
25 3 3 13 1 15 15 10 9 7 3 9 13 0 1 10 9 10 13 1 9 1 15 13 13 15
25 13 3 10 10 11 9 7 11 7 13 16 9 0 13 7 9 13 13 7 15 16 1 10 11 13
11 13 3 15 1 10 9 13 13 1 15 13
5 15 13 10 9 0
17 3 3 3 0 9 13 1 15 15 10 13 11 0 7 3 13 13
19 7 16 3 1 0 13 1 10 9 13 15 3 13 1 10 9 0 15 9
14 7 13 15 13 3 3 13 7 13 1 10 9 10 11
13 16 0 13 1 10 9 15 13 3 3 10 9 13
10 3 13 3 15 15 13 7 13 3 13
15 9 3 13 0 12 10 9 1 15 13 10 9 0 10 9
17 13 3 13 1 10 0 7 13 15 1 15 10 9 7 10 0 13
11 15 3 13 3 13 9 1 10 9 7 13
29 9 15 10 13 10 9 7 10 9 7 10 9 7 15 10 1 15 10 10 9 15 1 9 0 9 11 9 15 13
7 3 13 9 7 9 13 0
20 13 10 9 10 9 7 10 9 13 1 10 15 1 10 9 7 1 10 11 15
43 7 10 3 9 13 1 10 9 15 7 13 10 9 15 1 9 15 13 10 9 15 1 10 10 9 15 13 15 1 9 7 9 7 9 13 1 10 9 10 0 9 15 11
25 10 3 9 10 13 13 9 7 9 12 7 7 12 15 10 13 15 13 0 13 7 13 15 0 0
21 7 9 0 13 10 9 10 9 10 9 11 11 10 9 9 7 0 13 1 15 15
7 3 3 0 15 13 1 15
20 15 3 9 9 7 9 13 13 13 10 9 10 13 7 13 1 10 9 10 9
8 13 3 15 3 3 15 9 13
31 11 3 10 13 11 1 10 9 15 13 13 9 9 9 0 10 9 13 15 9 13 13 10 9 7 13 1 10 9 10 9
31 9 3 15 11 9 1 11 10 9 15 13 9 7 13 1 10 9 13 7 10 9 7 13 9 15 1 10 9 10 9 13
11 3 13 15 13 7 13 1 10 15 9 13
10 15 16 13 1 10 9 15 10 9 0
6 3 13 9 7 10 9
9 13 3 10 11 10 9 0 13 13
8 7 13 9 0 1 15 10 13
9 13 3 10 0 13 15 7 13 13
15 13 3 3 9 12 9 7 10 9 15 3 13 10 13 13
5 13 3 1 15 11
3 15 3 13
2 6 0
5 10 3 11 1 15
8 15 16 13 15 13 10 9 9
14 6 10 9 10 13 10 9 15 1 10 9 7 13 15
9 13 3 3 1 10 9 15 7 13
14 13 3 10 9 13 15 0 7 13 13 1 10 9 15
14 7 13 9 0 1 0 10 9 7 1 15 10 13 0
12 10 3 0 15 13 13 15 7 13 15 10 9
35 3 3 13 13 10 9 9 9 7 7 9 16 3 1 10 9 13 10 0 7 13 1 9 7 9 16 13 11 3 3 10 9 13 15 15
19 13 3 3 10 9 10 3 9 11 13 0 7 13 1 9 0 15 13 0
29 13 3 10 9 7 15 10 1 15 10 13 9 10 9 13 9 7 13 10 9 1 10 9 7 13 15 1 9 0
14 9 3 9 1 9 13 10 9 10 9 13 7 15 13
15 13 7 13 13 1 10 9 10 9 15 10 9 10 9 0
11 13 3 13 1 10 9 1 10 9 7 13
10 10 3 13 9 3 13 15 1 10 9
14 10 9 13 13 1 15 9 7 10 9 13 1 10 9
5 13 3 3 15 13
21 16 3 13 10 9 0 10 7 9 10 9 7 10 9 13 1 15 15 3 13 0
6 13 3 15 13 15 16
17 6 10 9 15 13 1 10 9 13 1 10 9 13 7 13 10 9
12 3 13 10 9 1 10 9 13 15 3 1 9
7 13 3 15 13 1 10 9
6 7 13 15 10 9 13
18 7 6 13 10 11 10 9 15 7 13 13 1 15 10 9 10 9 0
7 13 3 11 7 10 9 13
6 13 13 9 3 3 9
13 10 9 10 9 15 13 11 15 15 13 13 1 9
18 0 10 9 9 7 9 13 10 0 15 10 13 9 10 11 7 9 9
8 15 3 13 13 7 13 13 15
20 13 3 15 1 10 9 9 9 11 9 0 15 10 9 13 3 0 10 9 13
4 13 7 1 15
17 1 3 0 10 9 13 11 13 13 15 15 15 13 9 9 3 12
12 15 13 7 15 15 13 15 13 7 13 1 15
16 1 0 13 11 10 0 1 10 9 10 9 7 13 9 1 15
9 3 0 13 7 15 15 13 15 13
8 13 1 10 9 0 7 13 15
13 3 16 13 1 9 10 9 0 7 10 9 0 13
13 16 3 1 9 13 3 13 13 15 16 3 0 13
18 13 3 15 7 13 10 9 13 13 3 13 1 10 9 10 11 7 13
17 15 7 9 1 10 9 7 1 9 3 13 13 7 13 10 11 11
25 1 3 10 9 0 13 10 9 13 9 10 9 1 10 0 16 13 1 10 9 10 0 10 9 15
9 13 3 10 12 10 9 10 9 13
18 13 3 9 9 1 15 13 12 0 9 7 9 15 13 1 10 9 0
10 15 3 10 9 7 10 9 10 9 13
42 7 13 10 9 1 15 10 9 7 13 11 9 0 9 7 9 0 7 11 7 11 7 11 7 11 7 11 7 11 9 9 15 13 1 10 9 7 13 13 15 10 9
15 7 10 9 10 9 13 7 13 10 9 10 9 1 11 3
8 0 7 9 10 9 13 10 9
34 13 3 15 10 1 10 9 10 13 9 7 0 7 9 7 10 1 11 7 11 13 10 11 7 3 13 13 10 9 7 10 9 15 13
5 3 13 9 13 16
19 13 7 10 9 7 10 0 7 10 9 7 13 13 15 7 13 1 10 9
5 13 7 9 0 13
15 10 9 0 3 13 13 9 1 10 9 10 0 7 10 9
21 13 3 15 13 16 11 10 0 0 13 10 9 0 7 13 10 9 15 13 15 11
17 7 13 1 15 15 10 13 1 10 9 13 10 9 15 3 9 9
4 13 3 10 9
3 15 3 13
23 10 9 10 9 13 10 9 15 11 13 1 10 11 16 3 13 15 1 11 7 13 1 15
10 13 1 10 9 15 7 1 10 9 15
9 7 6 1 10 9 15 3 15 13
8 3 13 1 9 0 13 1 11
46 7 3 1 10 13 10 9 15 13 15 1 10 9 0 1 15 15 3 13 7 3 13 15 9 1 15 3 9 9 7 13 13 15 1 9 15 7 10 9 15 1 15 3 13 15 9
21 13 3 3 10 9 16 13 10 9 15 0 1 9 0 7 13 15 7 13 9 12
22 7 10 9 15 3 13 13 15 10 9 13 7 1 0 13 7 13 15 1 10 9 0
9 7 10 9 13 10 11 13 1 11
36 7 13 10 9 1 15 7 13 15 1 15 10 9 15 7 13 15 9 7 9 1 11 9 11 7 13 15 13 1 11 7 1 0 10 9 15
19 13 3 9 1 0 10 11 7 11 7 9 0 7 3 13 9 10 9 15
12 13 3 11 13 9 1 11 13 10 9 15 0
17 7 1 10 0 13 11 10 9 15 7 0 13 10 11 10 9 15
20 13 3 11 13 11 10 9 15 7 15 10 9 1 9 12 7 13 11 1 11
27 7 13 15 7 10 9 15 7 13 1 11 7 13 1 10 9 15 13 11 9 9 1 10 9 11 1 11
32 3 3 13 10 9 10 9 15 13 10 9 10 11 13 10 9 7 13 1 11 16 15 13 9 0 1 11 15 3 13 10 11
10 1 15 9 13 11 7 13 0 10 9
9 15 13 9 12 1 10 9 10 9
14 13 3 15 13 15 10 9 11 7 13 15 15 1 9
7 7 13 11 1 15 9 0
8 13 3 0 1 9 7 9 15
18 16 3 13 15 0 9 13 1 10 9 15 13 10 9 15 10 9 11
13 7 13 15 13 13 7 13 9 10 13 13 10 0
14 13 3 13 10 9 16 10 9 1 9 15 13 9 15
3 9 9 13
3 3 13 15
8 10 3 13 10 3 13 15 13
8 15 15 13 9 7 9 1 15
11 3 13 15 15 13 15 9 13 3 10 0
17 13 3 11 1 10 9 0 7 13 0 1 9 9 3 13 9 12
17 7 13 9 12 13 15 1 10 0 10 9 11 9 1 9 9 9
7 13 3 15 13 13 9 9
7 0 3 13 11 3 13 13
5 13 3 15 10 9
6 13 10 9 10 9 15
9 10 3 9 1 15 13 9 0 13
19 13 13 10 9 10 9 15 10 1 11 7 10 9 15 13 7 13 13 15
7 7 3 6 13 15 1 11
20 0 13 15 13 9 7 9 1 9 11 7 1 0 9 7 1 10 0 9 12
9 0 13 10 11 10 13 10 9 11
51 0 13 10 13 1 10 9 1 10 0 1 10 9 10 13 15 1 10 9 11 7 10 9 15 15 13 9 13 13 15 15 3 13 0 13 10 9 15 7 13 7 13 1 10 9 15 1 11 13 10 11
6 13 15 9 15 13 15
15 10 3 11 0 15 13 15 1 9 11 3 13 15 13 15
19 7 13 1 10 9 0 7 13 9 10 9 7 13 1 10 9 10 9 15
12 13 3 10 9 7 13 15 13 10 9 10 9
13 3 9 7 9 13 15 9 12 1 10 0 9 11
18 7 13 10 9 10 11 7 10 9 10 9 11 10 9 15 13 13 15
5 7 13 15 3 11
5 11 3 13 15 9
7 7 3 10 0 1 0 13
4 3 10 9 13
4 10 9 15 9
12 15 9 13 15 13 9 7 15 9 10 9 15
7 3 10 9 15 13 0 15
14 0 7 0 9 7 10 9 15 3 10 9 10 0 13
6 3 10 9 15 3 15
26 7 13 10 13 1 10 9 10 0 15 3 15 9 7 9 13 15 13 10 9 1 9 9 7 3 13
13 13 3 0 13 10 9 15 7 13 10 9 1 15
21 13 3 0 9 0 13 1 10 9 13 9 9 7 11 13 1 0 10 9 7 13
19 13 3 9 0 13 10 9 15 7 13 3 1 15 7 13 1 10 9 13
13 7 10 9 13 10 9 15 1 10 9 9 13 11
7 7 13 10 11 13 7 13
6 9 11 13 10 9 15
7 13 3 10 9 13 9 0
4 7 0 13 13
7 11 3 13 13 10 9 15
12 15 13 1 10 9 10 11 7 11 1 10 9
12 13 3 10 11 9 0 7 13 9 0 1 15
9 11 3 13 10 9 1 10 9 13
8 13 7 9 7 9 13 1 9
8 10 3 3 13 13 13 10 9
12 11 3 13 1 10 9 10 11 13 15 10 11
10 0 3 10 13 9 0 13 9 0 13
8 13 3 0 9 1 10 9 0
29 9 3 15 9 11 13 1 10 9 13 7 13 10 9 10 11 13 13 15 15 0 15 13 15 1 0 1 0 13
9 0 13 10 9 10 9 10 13 0
11 13 3 15 1 10 0 9 10 9 13 15
21 16 3 13 10 11 13 1 10 9 10 9 7 10 9 11 11 13 9 7 7 9
9 10 3 11 3 0 13 7 13 13
11 13 10 11 13 7 9 7 9 0 13 13
10 0 3 13 13 1 10 9 10 9 11
10 3 13 10 9 1 15 7 13 9 0
19 13 3 10 11 16 1 10 9 10 9 10 9 13 10 9 13 15 9 13
15 13 3 15 10 9 0 16 15 3 13 10 9 13 9 0
5 11 3 13 1 15
17 10 9 15 1 15 13 1 9 16 10 9 10 9 13 1 9 13
10 3 13 15 9 7 9 1 10 9 0
10 10 3 9 15 3 13 0 1 10 9
10 1 3 9 9 7 9 9 13 15 13
5 13 3 10 11 13
14 13 15 1 15 1 10 9 16 15 13 1 15 15 13
13 15 3 3 13 7 13 10 9 10 9 13 1 11
6 0 7 9 10 9 13
7 9 3 9 13 1 11 13
14 13 7 13 1 9 1 10 9 10 13 1 11 1 11
3 0 13 0
13 13 7 13 7 13 1 10 9 15 13 10 9 11
6 13 3 10 9 10 11
6 13 7 13 10 9 0
12 13 3 10 11 13 15 13 11 10 9 7 13
5 3 3 13 15 13
3 15 3 13
9 3 3 3 13 16 3 15 13 15
9 10 3 9 10 9 15 13 13 0
7 1 10 9 10 9 15 13
5 10 9 15 15 13
8 3 13 1 10 9 10 9 15
7 13 3 10 9 10 11 13
2 13 15
12 1 15 10 9 13 0 1 15 7 1 0 15
14 16 3 13 1 10 9 13 1 15 9 7 13 10 9
2 6 9
20 7 13 13 10 9 7 13 0 1 10 9 10 7 11 7 10 9 7 13 15
18 16 3 13 1 10 9 9 9 13 10 11 7 3 13 15 3 10 9
6 13 3 10 9 15 13
17 11 3 13 1 11 7 13 13 10 9 15 1 10 13 15 1 11
40 10 3 11 3 13 9 7 9 1 10 9 10 9 13 10 9 13 1 15 9 1 11 1 10 9 16 16 15 13 13 10 9 9 7 7 9 13 13 1 11
17 3 7 15 13 9 1 10 9 7 13 1 10 9 13 9 13 15
5 11 11 15 15 13
2 13 3
2 15 3
6 15 13 11 15 15 13
14 7 13 7 13 1 10 9 7 13 15 15 15 13 13
15 10 3 9 10 13 15 13 0 13 3 10 9 15 3 13
7 13 3 10 9 15 15 13
6 13 3 15 13 1 11
11 7 13 9 12 3 13 7 3 13 7 13
16 13 3 15 9 1 11 9 11 7 13 1 15 1 9 10 9
3 15 3 13
3 6 15 9
5 10 3 9 1 15
15 6 3 13 7 13 9 11 9 13 7 13 15 9 16 13
3 13 3 11
16 9 13 1 0 1 10 9 0 15 0 10 0 15 13 1 11
14 7 3 13 9 1 10 9 13 15 10 13 10 9 15
6 13 3 1 15 10 9
12 15 3 13 15 15 13 15 1 10 9 15 13
15 13 3 11 7 13 1 10 9 7 13 1 15 10 9 13
9 7 3 13 15 1 10 9 3 9
9 13 7 7 13 13 7 13 9 13
24 13 3 1 10 1 11 9 9 15 7 3 1 10 9 13 10 11 16 0 13 10 9 10 9
7 13 3 15 10 13 7 13
24 3 0 13 10 13 1 11 10 13 10 9 0 7 3 1 0 13 16 13 15 13 1 10 9
17 11 3 3 13 7 13 0 10 13 1 11 13 16 0 13 10 11
7 13 3 10 11 10 9 15
14 13 3 10 9 15 9 1 10 9 13 15 13 1 9
8 13 3 1 11 13 13 10 9
9 7 15 13 15 3 13 16 13 9
31 11 3 13 15 13 1 10 9 7 13 15 3 1 10 9 13 10 9 7 16 13 15 7 3 1 11 13 1 10 9 11
15 7 13 1 15 13 7 13 1 11 13 1 10 9 10 9
7 13 7 7 13 1 10 9
5 15 3 13 13 15
14 13 3 11 13 1 15 13 3 1 10 0 10 13 11
16 13 3 3 9 15 9 11 1 9 12 13 1 9 15 13 13
5 7 13 15 10 11
5 11 13 15 11 11
4 13 7 13 15
3 7 3 13
15 7 13 15 15 10 13 11 7 10 11 15 13 1 10 9
12 1 11 3 15 13 9 9 11 15 13 13 11
9 13 3 1 10 9 0 13 15 13
6 13 3 13 15 1 9
20 1 3 13 11 10 11 10 9 13 16 11 13 1 15 13 12 9 1 15 13
5 3 13 13 1 15
5 13 3 11 13 15
25 15 13 13 1 10 9 7 13 15 15 10 9 13 7 13 9 7 9 15 13 1 15 13 10 11
17 13 3 3 15 10 11 7 13 10 9 13 7 13 1 10 9 13
2 11 13
10 13 3 10 0 7 10 9 13 15 13
13 0 3 13 1 0 10 11 7 13 0 1 10 9
11 13 3 9 0 13 1 11 1 15 11 9
52 9 3 15 1 11 9 11 9 1 9 10 13 0 0 7 13 10 9 1 15 10 9 15 13 9 0 10 9 7 13 10 9 3 13 1 9 3 3 1 9 0 10 9 9 10 9 13 1 15 7 13 15
1 11
8 15 3 13 15 7 0 13 13
3 15 13 9
13 10 9 15 7 10 9 15 13 1 9 1 10 9
11 0 13 1 15 11 9 15 13 9 1 9
27 16 3 13 10 9 10 13 15 13 12 10 9 7 9 0 10 13 15 7 13 0 15 13 15 1 10 11
18 10 3 3 13 15 7 10 9 13 13 11 1 10 9 13 1 9 0
6 13 3 0 7 13 13
39 13 3 15 13 1 15 9 7 13 10 9 13 7 13 9 15 3 9 0 12 9 13 1 10 9 1 15 13 15 10 9 7 9 10 9 7 9 10 9
5 7 13 9 1 15
4 10 3 11 13
9 3 9 16 3 13 15 0 7 0
7 15 10 9 13 15 3 13
13 0 3 13 1 3 7 3 13 10 9 1 10 9
41 16 3 1 15 13 10 11 15 3 13 10 9 15 13 6 10 9 10 13 1 10 11 13 10 9 10 11 13 1 10 9 7 13 13 16 11 10 13 11 3 13
11 10 3 11 13 1 10 9 13 10 9 15
4 6 9 13 15
7 13 3 11 1 10 9 13
5 6 15 13 15 13
6 15 10 9 1 15 13
31 11 9 9 0 7 13 10 9 13 7 1 0 10 9 10 0 13 1 9 0 13 15 1 10 9 15 7 13 9 1 15
4 13 3 15 13
16 10 3 3 13 13 1 15 7 15 10 9 10 1 11 13 15
7 10 3 3 13 1 10 11
16 16 3 13 10 13 10 11 13 15 10 11 13 1 10 9 13
6 10 3 11 13 15 13
1 13
5 3 15 0 9 13
4 13 7 1 15
11 15 13 16 0 13 9 0 13 7 13 0
11 7 15 13 10 9 15 0 7 0 13 9
2 13 3
4 15 9 13 15
4 7 10 11 13
26 1 0 9 1 0 10 9 13 10 0 13 1 10 9 15 7 6 9 13 1 15 1 9 0 7 13
13 11 13 15 10 9 7 10 9 15 13 1 10 9
8 0 13 1 9 11 9 1 9
5 3 3 13 1 15
16 3 3 15 15 1 10 9 13 13 15 10 13 15 1 10 9
6 13 3 11 10 9 13
22 1 9 13 16 3 13 9 10 9 7 1 15 9 10 13 15 7 13 9 0 15 13
12 10 9 15 13 10 9 11 13 9 1 11 11
4 0 13 15 9
19 15 13 10 13 9 1 0 10 11 13 1 10 11 1 10 9 15 13 11
15 7 15 9 15 15 13 1 7 10 9 10 0 7 1 11
36 0 10 9 13 1 10 0 9 7 13 15 0 13 3 15 10 9 7 9 10 13 1 10 9 15 15 13 7 13 15 1 10 13 15 1 0
20 7 13 15 13 10 9 7 13 16 15 13 10 13 1 10 9 9 13 7 0
17 0 15 10 9 13 9 9 13 1 10 9 15 15 10 13 1 15
18 3 13 10 11 10 9 0 13 10 9 10 0 1 15 10 13 10 9
21 7 13 10 1 9 0 15 13 10 11 16 3 1 10 9 10 9 10 0 9 13
9 13 3 15 13 9 7 13 10 9
3 3 13 11
6 3 13 15 13 9 15
21 13 3 10 9 7 10 9 10 13 1 10 11 16 3 10 9 13 10 9 10 9
14 16 3 13 11 1 11 13 1 15 10 1 9 13 16
8 13 1 9 9 13 7 13 15
7 13 3 11 13 15 3 13
27 15 13 1 9 11 13 7 13 1 9 9 13 9 15 3 9 0 12 9 13 1 10 9 7 13 1 15
21 1 15 13 13 7 13 10 9 10 9 7 10 9 7 10 9 7 10 9 10 9
6 13 3 3 9 13 15
2 13 3
12 3 9 16 0 7 0 3 13 1 10 9 15
8 13 3 9 1 0 1 10 9
7 15 10 9 13 15 3 13
12 0 3 13 1 3 7 13 3 0 1 10 9
17 7 6 3 12 9 13 1 10 9 1 15 13 13 1 11 1 15
9 13 3 10 9 15 13 15 15 13
16 13 3 1 15 3 10 12 9 0 7 13 1 10 9 10 9
19 1 3 10 13 15 13 13 10 9 10 0 1 15 3 3 1 15 1 9
8 13 3 10 9 10 9 16 13
4 11 3 13 9
6 15 3 13 1 9 0
25 16 3 10 0 9 13 15 10 9 3 3 15 13 1 10 9 11 11 15 15 13 0 13 10 9
9 13 3 0 13 7 13 10 9 13
11 3 3 10 9 10 9 10 9 1 9 13
22 13 3 15 1 15 9 0 7 0 15 13 1 11 13 3 1 10 9 13 10 9 11
9 0 7 9 10 13 13 1 10 9
20 13 3 10 9 1 10 9 10 9 10 13 1 11 1 15 7 13 11 1 11
30 15 13 7 13 10 9 10 10 9 13 7 13 15 10 9 10 9 13 10 9 16 13 9 0 7 0 9 0 7 9
6 7 13 9 0 10 9
11 13 3 1 11 13 11 7 13 13 1 11
14 13 3 15 3 9 0 13 1 10 9 7 13 9 0
11 1 0 3 10 9 13 1 11 9 1 11
19 13 3 12 1 15 9 11 13 1 10 9 9 0 13 13 1 0 10 9
18 10 3 9 3 13 15 13 15 15 1 9 13 10 13 1 10 11 9
12 15 7 13 13 1 10 0 1 9 11 7 11
17 1 0 3 10 9 13 10 9 11 10 9 13 15 10 1 10 9
7 13 3 11 10 9 11 9
36 13 3 16 0 13 10 0 13 13 7 11 13 3 9 10 0 15 3 13 13 1 9 13 12 9 9 13 15 13 1 10 9 13 15 10 9
13 9 3 13 3 13 1 10 9 1 10 9 1 15
20 16 3 13 13 15 10 11 10 9 0 13 10 11 13 1 12 9 13 9 12
8 9 7 1 10 9 13 10 9
9 13 3 10 9 10 11 13 15 13
3 13 1 9
8 7 13 15 10 9 1 10 9
6 13 7 10 9 1 15
3 13 3 3
3 7 13 15
7 13 10 9 15 7 13 15
14 7 13 13 7 3 13 16 0 13 10 13 1 10 9
33 13 3 0 9 7 0 13 1 10 9 10 0 10 13 1 10 9 15 0 13 15 7 13 13 9 12 7 3 13 10 9 1 15
7 7 10 11 1 15 13 13
23 3 13 3 16 13 9 10 9 15 7 13 15 1 9 11 7 15 10 9 10 9 10 0
12 13 3 15 10 9 10 9 13 9 13 9 11
13 7 13 10 9 10 11 1 10 9 3 13 10 9
9 13 3 13 13 10 11 1 10 9
5 15 3 1 15 13
1 13
3 15 3 13
4 10 9 13 15
6 13 3 13 15 7 13
15 13 3 15 10 9 13 13 3 10 9 15 13 1 10 9
2 13 7
6 13 11 7 10 9 0
6 7 13 13 1 0 9
15 13 3 9 13 9 3 0 1 10 9 15 3 10 11 13
6 13 3 13 0 7 0
15 0 3 9 10 11 13 9 0 13 1 10 9 13 1 15
4 10 3 9 13
5 9 9 7 3 9
18 3 3 13 15 9 9 16 15 3 13 10 9 10 9 7 13 0 13
8 10 3 9 10 9 13 7 13
15 11 3 7 11 13 1 11 13 10 9 13 11 10 13 11
31 13 3 1 11 1 10 13 9 9 7 9 10 7 11 7 11 10 13 11 7 11 10 0 11 7 11 10 9 0 7 11
10 3 13 7 13 7 13 10 9 15 13
30 15 3 3 13 1 10 0 9 13 1 11 3 7 13 1 11 7 13 1 11 13 10 9 10 9 1 10 9 10 0
5 13 3 3 11 9
25 13 3 0 10 9 1 11 13 9 15 9 9 0 15 9 11 15 13 1 10 9 11 11 9 0
11 0 13 11 7 11 13 13 10 9 10 9
19 13 3 15 11 10 9 3 3 13 10 9 15 13 13 10 9 1 10 9
12 11 3 10 3 11 13 9 0 13 1 15 13
20 6 0 15 9 7 15 9 9 9 0 15 9 3 13 13 10 9 9 10 0
12 3 7 13 1 15 9 7 9 7 13 13 9
13 3 13 10 9 10 13 13 13 1 10 9 10 9
13 13 3 1 10 11 10 1 11 13 1 11 10 11
8 11 3 13 1 15 13 1 11
21 0 3 13 1 10 11 13 1 11 10 0 7 13 1 10 9 10 9 10 9 13
15 1 3 10 9 10 9 7 10 9 13 10 9 1 15 13
13 9 9 16 15 13 1 15 9 9 1 10 9 13
8 13 3 11 7 13 10 9 13
8 7 1 0 13 9 1 11 9
19 7 3 13 9 7 13 15 10 9 10 11 9 11 9 1 9 11 9 12
13 7 13 15 13 10 11 15 1 9 15 3 13 13
16 13 11 10 10 11 9 1 10 9 15 15 13 15 10 9 15
26 0 10 9 1 10 9 1 9 13 10 11 9 11 13 11 1 9 10 9 15 9 9 15 10 9 11
8 16 3 13 10 11 10 9 13
7 15 15 13 13 3 13 15
19 9 9 9 9 11 7 10 1 15 13 10 9 15 10 9 10 9 0 13
15 16 3 13 15 10 1 15 13 13 1 10 9 13 1 9
7 10 3 9 13 15 1 0
21 15 13 1 9 0 10 13 15 1 10 11 1 11 15 3 13 9 15 1 10 9
20 7 15 15 13 10 1 10 9 9 13 16 0 10 9 13 10 9 15 13 11
7 3 3 1 10 0 9 13
4 9 15 13 15
14 16 3 13 15 1 0 3 13 13 1 9 3 13 16
7 13 15 10 0 11 10 0
7 3 13 10 0 15 13 9
20 11 3 3 0 9 13 10 10 9 9 13 7 13 1 10 9 15 7 13 9
8 15 3 10 9 13 3 13 9
13 0 3 13 15 9 9 16 1 0 15 9 9 13
15 1 15 15 3 13 1 9 11 13 1 0 15 10 13 13
24 13 10 9 7 13 7 13 16 9 13 15 1 10 9 15 9 15 3 3 13 16 15 13 15
13 13 3 15 13 1 10 3 9 13 15 10 9 0
27 13 3 10 9 13 0 10 0 7 10 13 9 10 11 7 10 11 15 13 15 13 15 13 10 9 10 9
17 13 3 10 0 10 9 13 9 7 13 10 1 11 13 13 7 13
8 13 7 10 11 7 10 11 13
9 15 13 0 0 13 10 9 10 9
16 16 13 15 7 3 0 13 15 10 0 9 6 13 1 10 9
14 13 15 1 9 9 10 13 15 1 9 1 0 10 9
19 13 3 10 9 13 7 13 10 9 10 9 7 13 15 13 13 1 9 0
10 13 3 10 9 10 9 1 0 10 9
29 10 3 0 13 10 13 9 10 0 7 10 0 10 9 7 13 9 1 10 11 7 11 7 13 15 1 10 9 15
8 10 3 9 13 9 7 9 0
25 13 3 1 11 1 10 15 13 15 1 10 9 10 0 7 13 3 16 13 0 7 7 9 0 9
14 10 3 13 0 13 7 13 10 9 10 9 1 10 9
6 13 3 10 9 10 9
7 7 15 3 13 1 10 0
5 15 3 1 10 9
34 16 3 13 9 10 9 7 7 0 1 10 9 15 13 7 13 15 13 13 1 10 9 10 11 11 7 11 7 10 9 7 3 13 13
17 3 15 9 1 11 0 10 9 13 0 1 9 9 15 15 3 13
6 13 1 10 9 15 0
4 3 13 7 13
7 10 9 13 9 13 1 15
16 13 7 10 11 11 10 3 11 11 16 15 13 10 13 10 9
22 10 7 9 10 11 10 13 1 10 9 9 7 9 1 10 9 13 1 10 9 13 13
18 13 3 10 9 11 7 11 13 10 9 15 13 1 10 9 13 7 13
4 9 15 0 13
31 3 15 0 13 15 9 13 15 1 0 10 0 13 1 9 13 15 13 10 9 7 10 9 7 10 9 7 15 10 1 15
20 3 3 0 15 13 13 3 15 9 13 7 9 0 13 9 7 9 10 9 15
22 13 3 1 11 7 11 0 7 13 10 9 7 13 10 11 13 1 10 9 13 15 13
10 13 3 10 9 15 13 13 1 10 9
9 3 10 3 13 1 10 11 1 11
29 13 7 10 9 0 7 13 0 13 1 10 11 7 1 11 7 1 11 13 10 9 10 9 13 13 10 9 7 16
11 1 0 9 13 15 13 1 10 9 10 9
16 13 3 15 1 9 0 13 1 9 13 15 10 9 1 15 13
18 7 13 10 11 13 1 10 11 7 13 1 10 11 10 9 13 1 11
8 13 3 9 3 0 1 10 9
10 7 15 13 1 10 11 13 10 9 16
10 16 3 13 10 9 10 11 3 13 13
35 13 3 9 7 9 3 0 10 11 7 10 11 1 15 13 13 11 7 11 7 15 15 1 15 1 10 9 7 0 1 11 1 10 9 0
25 15 3 3 13 1 10 9 13 10 7 11 7 11 13 10 9 10 9 7 13 9 0 15 10 9
14 13 3 1 11 13 1 10 9 7 10 9 7 10 0
8 13 7 15 10 9 13 1 15
12 13 3 15 10 1 10 9 10 9 13 13 16
12 13 3 10 9 7 10 0 13 1 10 9 0
9 0 3 9 13 13 11 13 1 15
26 9 9 15 13 16 1 9 0 1 15 13 10 9 1 10 9 15 13 10 9 10 9 10 9 7 13
28 7 10 9 9 13 15 13 10 9 10 0 3 3 15 7 15 13 1 15 7 7 15 10 9 13 10 9 15
22 3 3 15 13 10 9 13 9 1 10 9 10 9 15 7 10 9 15 7 15 13 13
14 7 1 10 9 10 9 11 13 13 1 15 9 3 0
23 13 3 15 10 9 7 13 11 7 11 13 15 13 10 9 9 7 9 1 10 9 1 15
8 1 3 10 13 15 13 11 13
7 7 0 13 10 9 10 9
2 3 13
39 1 0 13 7 13 10 9 11 10 13 7 10 13 15 13 7 13 15 16 3 13 10 0 10 9 10 9 7 15 10 9 1 15 13 10 9 15 1 15
7 13 9 13 0 0 1 9
31 3 15 13 3 13 10 1 10 9 13 1 10 9 7 13 15 10 13 10 9 10 9 7 10 9 7 10 0 7 10 9
18 11 3 1 9 0 1 9 10 13 15 13 1 10 9 1 15 9 13
34 3 13 10 9 7 10 0 1 0 10 9 13 9 1 15 13 1 11 1 10 11 7 11 11 10 13 11 7 11 9 13 1 10 9
19 10 9 7 10 0 9 10 1 10 11 7 11 7 11 9 10 1 9 13
12 13 3 11 7 11 3 0 1 9 13 10 15
25 13 3 10 9 10 0 7 15 15 0 13 15 9 1 0 10 3 13 0 7 9 7 0 7 9
6 1 15 13 15 3 13
1 13
14 15 3 3 13 13 1 11 7 13 10 9 13 10 9
6 13 3 13 1 10 9
13 13 3 9 13 1 9 1 10 9 1 10 13 15
18 11 3 7 11 13 1 11 13 7 13 1 3 0 0 10 9 10 9
17 13 3 13 10 9 1 9 15 1 15 13 10 9 10 9 3 13
10 11 3 13 13 3 10 11 10 13 11
19 11 3 13 10 13 1 15 1 11 7 3 13 15 1 10 9 3 13 0
17 13 3 9 16 13 15 1 15 10 7 11 13 10 11 13 1 11
13 11 3 13 11 13 13 10 9 10 9 1 10 9
7 13 3 1 11 7 1 11
24 7 6 9 15 13 3 9 11 9 9 0 0 9 3 9 15 13 1 10 1 11 7 11 9
20 0 13 10 11 1 15 13 7 13 13 15 1 10 0 10 13 1 10 9 0
20 16 3 13 10 9 13 15 13 10 9 10 13 1 10 9 7 0 10 1 11
13 10 3 3 9 13 10 9 7 13 10 9 1 9
18 13 3 10 11 7 0 9 13 1 10 0 9 13 10 9 1 10 11
17 13 3 1 10 11 13 1 10 11 13 7 3 13 15 10 9 11
7 7 9 1 9 10 11 13
10 9 9 15 13 13 7 13 15 7 13
5 13 1 11 13 15
18 16 3 10 9 13 3 13 13 1 11 13 16 13 15 10 9 13 15
9 13 3 1 0 10 9 13 9 15
21 10 7 9 10 9 13 1 10 9 1 9 3 13 9 13 7 13 13 10 13 9
23 7 15 9 9 11 9 9 11 13 10 9 13 15 10 9 13 10 9 13 10 13 1 11
13 16 13 15 0 10 9 13 13 1 10 9 15 13
3 7 13 15
22 13 3 13 15 1 10 9 9 15 13 9 9 13 15 15 9 0 13 10 9 15 13
8 0 13 10 11 7 15 13 13
14 0 10 9 9 10 9 10 0 13 15 13 15 9 9
8 13 3 11 7 13 10 9 13
9 13 15 1 9 11 11 13 1 15
31 13 3 10 9 15 16 13 10 9 10 9 15 13 10 11 7 10 11 13 1 10 9 1 10 9 7 13 15 10 9 13
21 0 10 9 13 15 10 9 0 13 7 13 9 15 3 13 15 13 7 13 0 13
29 7 13 10 9 1 15 7 10 9 13 15 10 9 13 13 0 7 13 15 9 13 1 9 13 10 9 3 13 15
18 15 9 0 13 13 15 1 10 0 9 7 10 9 13 15 1 10 9
11 1 3 10 9 11 7 11 13 13 10 9
5 13 3 15 10 9
11 13 3 3 10 9 15 7 15 10 9 13
6 13 3 9 0 11 13
4 15 13 15 0
4 0 3 13 3
18 13 3 9 13 7 0 13 13 10 11 7 10 11 7 13 15 3 13
7 9 15 15 13 13 16 13
3 15 3 13
12 13 1 10 9 11 7 13 15 7 10 9 15
14 13 7 15 1 10 9 13 9 7 13 3 13 10 9
9 9 3 13 13 10 9 10 9 13
4 13 10 9 0
11 13 3 10 9 10 9 0 1 10 11 16
5 13 10 9 16 13
6 3 3 13 13 1 9
6 10 3 11 13 1 15
10 13 15 3 0 9 0 13 13 1 9
7 3 3 7 13 0 15 13
9 13 7 10 9 10 9 10 9 0
17 13 3 13 16 0 13 7 13 13 15 7 13 13 13 1 10 9
16 13 3 1 10 9 13 1 10 11 7 13 13 10 9 7 13
15 13 3 10 11 7 10 11 13 1 11 3 13 9 10 0
32 1 3 10 13 10 11 13 1 15 7 1 9 12 13 15 1 10 9 13 7 13 16 10 11 13 13 7 13 1 0 7 16
8 0 13 11 11 15 15 13 15
24 7 15 1 15 13 7 13 10 11 7 10 11 10 7 13 9 9 0 9 7 10 0 3 0
11 10 10 9 13 0 3 3 13 15 13 11
13 7 0 15 1 10 9 9 13 9 0 13 13 11
21 13 3 10 9 7 10 9 13 0 7 13 10 0 1 10 11 7 10 0 13 15
23 10 3 9 3 1 9 13 10 7 11 7 10 11 1 11 15 13 1 10 9 10 0 13
23 0 3 13 0 10 1 11 15 13 10 9 1 15 9 1 9 13 10 9 16 13 0 3
16 0 3 3 1 15 13 7 10 0 9 10 0 7 9 3 0
29 16 3 13 10 1 10 11 0 16 3 1 10 11 13 1 10 11 10 9 10 9 13 3 3 13 7 13 10 9
9 13 7 10 7 11 7 10 11 3
19 1 3 10 11 13 15 10 11 13 10 9 15 1 15 13 0 13 10 9
21 13 3 3 1 10 9 10 0 7 10 13 7 1 10 9 1 15 9 1 10 13
13 15 3 7 10 9 7 0 9 13 15 7 15 13
7 15 3 13 10 0 0 13
2 15 3
5 0 9 13 9 13
9 13 7 15 1 10 0 9 13 13
11 13 13 15 10 0 0 10 1 15 13 9
7 13 3 13 15 13 0 13
18 0 3 15 7 10 13 0 1 15 0 13 3 13 15 7 13 15 0
9 13 3 11 1 0 10 0 9 13
8 9 0 1 15 3 0 15 13
13 13 3 7 13 10 9 15 13 3 9 1 15 13
8 15 3 13 13 0 15 13 15
38 10 9 10 13 10 9 7 15 10 1 15 0 9 7 9 13 9 3 1 0 9 13 7 1 9 0 13 13 15 0 13 15 9 7 9 7 10 15
39 13 7 1 12 15 9 9 13 1 15 9 10 9 13 13 9 7 10 9 10 9 15 13 10 9 16 3 13 15 7 13 3 3 3 1 12 0 15 13
8 3 3 15 10 1 15 9 13
5 15 3 3 9 13
22 9 3 13 10 9 3 13 13 9 7 9 7 9 9 9 7 9 9 10 0 13 0
39 10 3 3 9 10 9 13 10 9 10 3 13 10 9 15 3 13 16 13 9 1 15 13 13 10 9 1 9 1 9 15 13 9 13 15 13 15 1 0
3 15 3 13
6 13 15 1 0 3 3
7 3 10 11 13 1 0 15
20 15 3 9 13 15 13 1 15 7 11 10 9 7 9 9 11 7 0 1 15
41 7 13 15 0 9 11 0 10 9 3 13 1 10 11 7 11 9 15 1 10 13 11 13 15 10 0 1 10 11 13 15 7 1 10 0 13 13 1 15 7 13
5 13 3 9 10 9
8 13 3 1 10 9 1 15 9
24 16 3 13 1 10 11 10 7 11 7 10 11 13 10 9 10 11 13 10 0 13 10 11 11
11 13 3 15 7 13 13 10 9 13 1 15
7 10 9 15 1 10 9 15
2 0 15
7 1 10 3 1 10 9 13
20 11 3 10 9 13 10 9 1 0 10 9 15 7 0 10 0 13 13 7 13
10 13 3 10 9 1 9 1 9 10 11
13 13 3 9 7 9 12 13 1 15 10 9 10 9
30 11 3 9 13 10 11 13 3 10 0 10 11 7 13 15 1 10 9 13 16 1 10 9 13 0 10 9 13 10 9
13 13 3 10 11 13 10 9 13 10 11 1 10 0
15 16 3 13 9 15 3 9 0 6 0 1 9 3 13 15
15 16 3 9 13 1 9 7 9 7 9 10 1 15 13 0
6 9 15 0 3 13 13
10 13 3 15 11 10 9 13 1 10 9
25 10 3 11 3 13 9 0 10 9 13 13 1 10 11 7 1 15 11 7 11 13 1 11 10 9
3 13 3 9
8 13 3 1 11 7 0 13 3
9 15 3 13 1 10 9 13 10 0
24 13 3 15 1 0 9 13 3 13 7 13 7 13 3 13 1 15 10 9 13 13 1 10 11
28 7 13 1 11 13 7 13 10 9 13 1 11 7 13 9 15 13 13 3 10 0 9 7 11 13 15 10 9
18 0 3 15 11 9 9 10 9 9 0 13 1 11 0 13 1 10 9
16 13 3 15 11 7 11 13 15 7 3 15 13 10 9 10 9
15 13 3 15 13 1 10 11 13 10 9 13 10 9 13 15
9 15 13 13 0 10 13 1 10 9
14 3 3 10 0 13 3 13 1 10 9 13 10 11 11
21 13 3 1 10 10 11 13 1 11 11 13 10 0 9 13 1 11 7 13 15 9
4 13 7 1 15
5 3 9 0 13 13
4 15 3 1 15
3 15 3 13
4 1 15 3 13
3 15 3 13
4 1 10 11 9
3 13 3 11
19 11 13 9 9 10 9 13 1 10 13 1 15 16 13 0 13 1 10 11
22 13 3 13 1 10 9 10 9 11 7 13 15 10 11 9 13 10 9 10 0 1 15
5 13 7 9 7 13
25 16 3 15 13 7 13 13 10 9 1 10 9 13 1 15 13 10 9 1 9 13 1 10 9 11
21 0 3 13 1 9 12 16 15 10 13 10 11 13 10 9 10 9 0 7 7 9
37 9 7 3 10 13 10 9 13 1 10 9 11 16 3 1 10 13 13 1 10 9 15 9 7 9 7 13 1 15 10 9 10 7 9 10 0 13
22 13 3 15 3 10 13 0 9 13 1 10 13 10 9 10 0 10 9 10 9 11 13
7 13 15 10 11 15 11 13
10 13 3 15 11 0 9 12 9 0 13
8 13 3 10 9 10 0 13 15
4 15 3 15 13
37 0 3 13 0 15 0 7 7 9 10 13 10 11 7 13 9 1 15 15 7 13 10 9 10 9 11 0 7 10 13 13 13 7 13 10 9 15
12 0 3 10 10 0 13 13 10 9 13 1 15
10 7 13 10 9 15 7 13 9 9 12
10 3 1 9 10 9 10 9 13 7 13
20 16 3 13 0 13 10 11 1 10 9 13 10 11 7 11 13 1 11 13 16
10 1 10 13 15 3 13 15 3 11 13
12 13 3 1 10 9 0 9 3 0 1 10 9
24 11 3 15 9 9 13 9 0 11 13 10 9 3 0 9 15 13 7 10 1 10 0 9 13
37 3 0 3 0 13 15 10 9 1 9 13 7 3 10 10 0 9 9 11 1 15 13 13 7 3 13 10 9 15 15 0 10 11 7 10 9 13
8 13 3 7 13 0 9 13 13
4 0 10 11 0
6 7 13 10 9 10 9
13 13 7 3 1 10 9 13 11 7 11 9 9 11
18 15 3 3 10 9 13 15 9 13 1 15 13 3 13 15 1 10 9
6 15 3 3 15 15 13
13 13 3 10 9 13 7 10 0 3 13 15 1 13
10 10 3 11 13 10 9 13 13 10 9
15 13 3 16 0 13 9 13 12 1 15 3 1 9 12 13
4 0 10 11 0
7 13 3 10 9 10 9 13
13 0 3 13 0 13 13 15 13 13 7 15 0 13
12 13 3 10 9 0 7 0 7 13 10 9 15
18 16 3 3 11 7 10 1 15 9 13 1 15 9 0 13 7 9 13
2 13 15
20 3 3 13 13 9 1 10 3 15 0 13 1 15 3 13 13 9 10 9 0
6 7 0 13 13 10 9
18 1 3 10 13 10 9 13 10 11 10 9 7 13 13 13 13 1 11
21 13 7 9 12 13 9 15 1 10 0 13 13 1 10 11 13 9 10 13 1 11
21 13 3 15 11 11 0 9 3 11 7 11 7 11 0 7 11 9 3 11 7 11
7 0 3 13 13 15 1 11
24 15 3 13 1 10 9 10 0 1 11 7 13 1 15 1 10 11 1 9 12 3 13 9 12
18 1 3 10 12 10 9 13 15 13 9 10 11 13 15 13 13 10 3
10 13 3 9 0 1 10 9 3 13 13
29 13 3 15 9 9 11 1 10 9 13 9 0 13 10 11 1 0 13 1 10 9 13 1 10 9 3 7 13 0
2 3 13
7 10 3 9 15 1 15 13
16 13 3 7 13 10 9 7 13 1 0 7 13 1 9 3 13
9 13 3 10 9 13 7 13 3 3
15 15 3 13 1 10 9 13 1 10 11 3 13 13 10 11
7 3 3 13 13 13 0 13
8 7 3 13 10 13 13 1 11
6 10 3 13 13 1 11
15 13 3 10 11 13 10 11 16 3 13 15 13 1 10 11
13 13 3 16 0 13 15 10 9 10 9 13 1 11
12 1 3 10 11 13 1 11 13 10 0 10 9
7 16 3 13 1 15 13 15
36 15 13 1 0 9 1 15 13 1 10 11 3 1 15 10 15 9 13 13 10 9 1 15 9 7 9 7 9 10 13 15 1 10 9 10 0
33 16 15 13 10 13 10 3 13 15 7 13 15 3 7 1 9 13 0 7 7 9 10 1 9 9 7 9 1 10 9 15 11 11
19 7 3 6 15 13 16 3 13 10 9 15 15 15 1 15 13 13 10 9
14 3 13 15 1 10 3 9 16 0 13 1 10 9 15
12 3 3 13 10 3 13 15 10 9 10 9 15
27 13 15 7 15 10 9 1 15 15 10 9 10 0 13 9 13 10 9 10 9 15 13 1 10 9 10 0
30 15 13 16 13 1 10 9 15 9 0 1 15 3 13 10 9 7 1 15 0 13 9 13 13 10 13 10 9 1 15
15 3 13 13 16 9 9 7 9 3 13 1 9 13 12 0
24 7 10 3 13 15 10 9 7 10 9 10 9 15 10 13 13 7 13 10 9 1 10 13 15
7 9 7 9 7 9 15 13
20 15 13 15 16 3 13 13 13 10 13 13 7 10 9 10 9 11 16 15 13
6 0 13 3 13 3 13
11 7 0 13 13 10 9 15 1 15 15 13
28 0 3 9 13 15 7 13 1 10 9 10 11 13 15 13 3 1 10 9 15 13 16 3 13 10 9 15 13
6 13 3 15 1 10 9
23 16 3 13 13 15 13 1 15 13 13 1 10 11 10 3 3 1 10 11 7 3 1 11
8 7 13 9 13 1 11 13 13
15 13 3 10 11 7 13 15 0 13 1 11 7 13 1 11
35 16 3 13 15 13 10 9 13 13 13 15 15 1 9 7 9 1 1 10 9 7 13 10 9 1 10 9 13 13 15 7 13 1 10 9
6 0 3 13 1 10 0
19 15 3 10 9 13 1 11 13 1 11 7 13 10 9 13 9 12 1 15
22 10 3 3 13 13 1 11 7 13 1 10 9 11 10 9 13 1 10 12 13 1 15
7 0 3 13 9 12 9 13
30 13 3 9 0 13 15 1 10 11 9 9 11 7 13 1 15 7 13 10 9 10 11 13 15 10 9 7 10 9 13
6 0 13 10 9 10 0
16 16 3 13 0 13 15 7 7 10 0 10 3 13 15 1 11
8 15 13 13 7 13 15 10 9
18 15 3 3 0 13 7 3 13 1 11 3 13 1 10 9 10 9 11
6 3 13 3 15 13 13
5 10 9 10 9 13
9 1 3 10 9 0 13 13 1 11
18 13 3 3 10 9 1 11 1 15 13 1 15 13 11 15 0 0 9
15 10 7 13 13 10 11 1 15 1 11 15 7 13 10 0
18 7 13 15 13 1 12 0 15 13 10 9 1 10 9 1 10 9 15
3 13 7 15
13 13 9 15 9 13 10 13 7 15 9 10 9 13
25 13 3 1 15 16 9 13 1 11 10 1 10 9 15 0 13 3 13 15 10 9 7 10 9 13
3 15 3 13
4 3 13 13 9
6 0 3 13 15 15 13
8 13 15 9 12 9 13 1 15
30 0 13 13 1 15 7 13 1 15 16 13 10 9 7 13 15 16 15 13 1 15 15 13 7 13 3 0 13 10 9
32 3 10 11 13 10 9 10 13 9 1 15 13 13 1 10 9 13 10 9 10 9 10 9 16 15 13 1 12 0 15 10 9
28 16 3 13 10 12 9 13 10 1 10 11 0 13 15 1 10 9 13 15 10 9 7 13 1 15 10 9 13
3 9 9 13
18 0 13 10 9 10 1 10 9 7 10 9 7 10 9 0 15 3 13
20 13 3 13 11 10 0 1 10 9 1 15 15 13 16 1 10 9 13 10 11
24 13 7 10 9 0 7 13 9 10 9 7 13 10 11 13 15 1 10 9 7 3 13 10 9
23 13 7 15 13 13 9 10 9 10 9 16 0 13 11 15 3 13 9 7 9 13 1 15
12 15 3 13 10 9 7 10 9 13 13 10 11
8 15 3 0 15 13 1 10 9
16 3 13 3 15 13 10 0 1 10 9 13 13 15 1 10 9
17 16 3 13 1 10 9 13 13 15 1 10 9 1 10 9 10 9
2 13 15
11 13 7 13 1 10 9 10 11 13 10 9
7 3 13 15 13 15 1 15
3 15 3 13
2 3 13
4 13 3 10 11
12 15 9 3 13 0 9 10 11 3 0 9 9
6 13 15 13 1 10 9
14 13 3 15 10 11 13 1 10 9 13 10 9 10 9
9 0 3 9 13 13 10 0 9 13
11 9 9 7 9 13 15 10 1 15 3 9
11 13 3 16 10 0 9 13 15 3 13 9
2 7 13
26 15 0 10 9 13 1 9 13 7 13 1 9 9 7 7 9 3 3 10 9 13 15 7 15 10 9
19 13 3 15 13 7 13 10 11 1 9 3 1 10 9 13 9 0 1 15
10 13 7 1 10 9 7 13 9 13 15
5 11 11 15 15 13
3 15 3 13
3 15 13 9
4 13 7 1 15
8 15 13 11 10 0 15 15 13
2 13 3
3 15 13 9
6 10 3 9 13 1 15
14 13 13 1 11 7 3 15 13 1 15 15 13 15 13
18 16 3 3 13 1 10 9 10 9 0 13 1 10 13 15 13 1 11
21 11 3 15 9 0 1 10 9 13 1 15 10 13 0 13 1 15 7 13 13 15
3 11 9 13
8 7 15 0 10 9 13 1 15
33 10 9 10 9 15 13 15 13 10 9 15 7 13 10 0 7 13 9 1 10 9 15 16 13 9 15 1 15 9 15 13 7 13
4 7 3 15 13
11 13 13 7 13 10 9 15 13 10 9 15
21 13 3 15 13 1 11 7 13 15 1 10 9 13 15 1 9 7 13 15 13 15
14 13 7 13 1 9 1 11 16 3 13 15 9 1 15
3 7 15 13
16 9 0 13 16 15 13 13 7 13 1 10 9 10 13 1 15
22 7 16 13 10 9 11 10 9 15 3 0 13 13 7 13 7 13 10 9 10 13 15
13 13 3 15 1 0 10 9 7 13 10 9 15 13
6 13 1 10 9 10 0
5 3 3 13 15 13
33 13 3 15 7 13 10 9 7 9 13 1 10 9 13 10 9 13 15 1 10 9 13 9 13 15 16 13 1 15 9 3 13 15
13 16 3 13 15 10 9 13 1 10 13 9 10 11
8 3 9 0 7 0 13 15 13
9 13 3 10 9 13 10 9 13 13
6 10 3 9 0 0 13
2 13 15
3 15 0 13
4 15 3 13 6
4 13 3 10 9
7 15 0 9 10 9 0 13
4 10 3 11 13
9 3 3 13 1 15 10 13 15 13
14 7 10 9 3 13 13 16 0 13 7 16 15 13 13
7 13 3 10 9 10 11 13
13 9 9 15 15 9 0 13 10 9 1 0 10 9
12 10 3 9 11 13 10 13 15 13 15 10 9
6 3 10 11 1 15 13
7 13 15 13 10 9 9 13
4 10 3 13 13
5 10 9 10 9 13
4 13 7 10 11
10 13 3 16 9 10 9 15 3 13 3
18 13 3 10 11 16 10 12 9 13 9 10 3 0 9 13 1 10 9
7 9 9 15 9 13 9 9
7 1 9 7 9 0 15 13
11 9 3 3 13 3 13 9 7 9 7 9
5 9 3 13 10 0
15 13 3 9 0 7 13 15 10 9 10 9 10 9 13 13
7 15 0 13 1 10 9 0
27 0 3 13 9 13 10 9 16 13 10 11 1 15 13 10 9 13 13 15 1 0 15 13 7 1 10 9
9 10 3 13 9 13 15 10 9 13
1 13
19 13 3 9 13 9 10 0 13 15 13 7 13 7 13 16 15 13 10 11
9 13 3 0 12 10 0 10 9 13
8 15 13 10 9 7 10 0 13
10 9 13 15 15 13 16 15 13 10 11
21 3 3 15 13 10 9 1 10 9 16 13 15 1 15 3 13 13 3 10 1 15
18 13 3 10 9 10 9 11 10 9 13 7 13 1 10 9 13 10 11
8 13 3 10 11 12 10 9 13
5 13 3 15 13 15
11 15 3 3 13 15 13 1 10 9 7 13
16 10 9 11 13 15 13 0 10 9 13 1 15 13 15 13 15
12 13 3 10 9 15 10 9 7 13 1 0 13
6 15 13 15 13 13 15
24 13 3 16 10 0 13 10 13 15 16 3 10 11 13 1 10 9 3 13 15 3 13 1 15
28 13 3 15 1 15 9 0 12 15 13 15 7 13 7 13 16 15 13 15 7 3 13 0 13 10 1 15 9
7 7 13 15 12 10 9 13
18 13 9 12 16 13 1 11 7 9 12 7 9 12 1 0 9 10 9
18 9 7 13 16 13 10 11 13 1 11 10 9 13 9 13 10 9 0
7 11 11 10 0 9 11 13
21 10 9 0 13 1 10 0 7 13 13 1 15 13 1 10 9 13 13 16 0 13
14 13 7 13 10 9 1 15 13 15 13 1 10 9 15
16 15 13 13 1 9 10 9 15 15 3 0 9 7 9 13 9
16 15 13 1 10 11 7 13 10 9 10 9 13 3 10 11 15
22 1 3 12 9 13 10 9 11 1 0 15 7 9 11 15 15 13 10 9 1 10 11
8 13 3 15 13 13 10 11 13
25 0 9 13 1 15 7 9 13 10 9 0 1 10 15 9 3 7 7 3 13 0 11 1 15 9
15 16 3 3 1 0 15 13 13 13 15 15 3 10 15 9
9 13 3 3 10 0 13 0 3 13
9 13 7 10 11 13 15 10 9 13
62 1 0 9 13 15 9 10 9 0 13 3 10 1 15 13 13 15 13 16 3 0 13 15 9 12 1 15 13 13 1 11 7 7 1 10 9 13 15 1 15 13 7 9 13 9 7 1 10 9 7 1 10 9 7 13 13 15 1 15 3 13 15
15 1 0 7 0 13 0 9 13 1 10 9 7 10 9 3
27 1 9 3 0 9 13 1 10 9 15 13 7 9 1 15 13 15 13 1 10 9 3 1 9 7 1 9
18 15 3 1 10 11 0 15 13 1 15 13 7 13 16 15 13 1 15
31 7 0 0 13 15 13 9 13 15 1 10 9 3 1 12 0 9 15 13 1 15 13 16 1 9 0 15 13 3 1 15
26 1 3 9 15 13 10 11 1 11 10 0 9 13 0 13 10 11 7 13 15 1 10 1 11 11 9
17 13 3 15 1 9 7 9 7 10 9 10 13 0 13 10 11 13
4 10 3 13 13
5 9 3 13 13 15
9 9 3 13 13 9 10 11 11 11
12 13 7 9 13 10 0 10 11 13 10 11 13
13 11 3 13 10 0 1 12 9 13 1 11 1 11
32 13 7 15 10 9 7 10 0 10 0 1 10 11 7 13 15 13 9 1 15 16 13 15 1 11 9 13 13 15 1 10 9
16 10 3 3 11 13 13 10 11 1 11 15 3 13 1 9 13
16 10 3 1 15 13 0 13 16 15 13 1 10 9 0 13 15
23 13 3 1 15 9 3 0 12 7 12 13 1 11 10 3 13 1 10 9 13 10 11 13
15 7 1 10 9 10 0 7 1 10 9 7 1 9 15 13
10 13 1 11 13 3 1 0 13 1 15
4 13 3 10 11
8 0 15 13 3 3 15 3 13
13 16 3 3 13 7 0 9 13 15 3 13 10 13
13 16 3 15 13 15 0 13 15 15 15 13 15 13
2 9 13
2 9 13
3 1 9 13
16 16 3 0 9 13 3 10 11 10 9 13 10 1 10 11 13
25 9 15 13 13 1 11 9 1 15 13 15 1 11 13 10 9 7 10 0 10 0 13 1 15 9
27 1 15 13 16 3 13 9 0 13 15 9 16 3 10 13 1 9 13 10 9 9 7 9 13 1 10 9
16 13 3 3 9 15 13 10 3 13 1 10 9 13 13 10 9
12 1 15 13 10 9 15 9 13 15 15 13 0
18 13 3 15 10 1 0 9 13 16 13 13 1 11 7 3 13 1 0
20 10 3 11 13 13 15 1 10 10 11 9 13 13 15 16 15 13 15 1 9
5 11 3 1 10 11
4 3 13 13 15
34 10 3 3 13 10 11 7 10 11 1 0 9 7 13 1 10 9 1 7 9 7 9 10 1 9 10 9 7 13 10 11 13 10 11
4 7 13 10 11
30 11 9 7 15 10 13 15 9 13 0 1 15 0 10 9 10 0 13 15 1 7 11 7 3 13 3 13 15 13 3
8 0 3 0 13 10 11 13 13
9 1 15 0 15 13 10 9 3 13
18 3 13 15 1 15 7 3 1 15 9 11 16 10 9 13 13 15 13
13 0 3 15 13 13 9 3 3 10 1 15 9 13
5 13 15 1 15 13
7 3 10 11 13 10 9 13
28 1 15 15 13 1 0 9 11 13 15 0 1 15 13 3 13 3 9 15 13 15 10 1 0 9 7 7 9
39 10 3 3 9 15 10 1 9 10 1 9 13 1 10 9 15 1 7 11 13 15 10 0 13 15 3 16 13 13 16 1 10 0 9 10 15 9 13 9
29 7 3 1 9 10 1 10 9 15 9 13 1 10 9 13 13 1 15 10 9 15 1 9 9 7 9 13 13 13
7 1 15 9 13 1 0 9
10 15 0 13 1 15 16 10 9 0 13
15 15 3 3 13 15 1 10 9 11 10 0 13 0 0 13
15 7 0 7 10 0 15 1 9 13 10 1 10 9 9 13
15 13 7 15 13 9 7 1 15 10 9 3 13 15 13 13
34 1 15 13 1 10 11 1 9 7 9 10 10 9 9 0 1 10 9 13 9 3 1 10 9 10 9 13 15 9 7 10 1 15 13
15 15 7 13 15 1 10 9 13 9 13 1 15 10 0 9
5 11 11 15 15 13
5 0 15 1 9 13
3 15 3 13
3 15 13 9
6 15 13 11 15 15 13
62 1 0 3 13 15 13 15 9 7 9 15 7 13 15 7 13 15 13 15 1 10 9 7 1 10 9 1 15 15 13 15 13 9 15 10 13 1 9 1 9 7 10 9 10 11 1 10 9 10 13 15 9 9 7 9 1 10 13 9 10 1 15
38 3 9 11 3 13 0 10 0 9 7 10 1 11 0 7 7 11 15 7 10 9 10 11 7 10 9 13 13 7 13 1 10 9 0 10 9 9 13
11 1 0 15 0 13 13 1 10 9 13 13
47 9 3 13 10 1 10 9 1 10 9 0 13 13 0 7 7 0 15 1 13 15 7 10 9 13 13 13 7 11 16 0 10 11 16 0 1 9 0 9 13 13 10 7 9 7 10 9
10 0 3 15 13 10 11 0 10 9 13
2 13 11
7 10 0 15 9 1 9 13
11 13 3 1 0 10 9 1 15 3 13 13
7 13 3 15 0 3 13 15
7 3 3 13 1 9 13 0
5 13 9 11 10 9
3 13 16 13
6 10 3 11 1 10 11
6 1 0 15 13 9 13
3 10 3 11
31 13 7 10 9 7 10 9 10 7 11 7 10 13 15 7 13 13 1 15 13 16 15 9 7 9 0 15 13 10 9 0
5 11 3 10 11 13
9 13 13 10 9 0 16 3 13 9
22 16 3 13 10 13 15 1 10 11 13 10 7 11 7 15 0 9 9 9 11 9 0
19 13 3 9 0 13 13 1 10 1 10 11 9 13 13 1 15 11 9 9
6 10 7 0 13 1 11
14 3 7 10 11 10 11 13 13 1 10 9 13 9 13
12 7 3 13 13 10 11 1 10 10 9 13 0
21 1 0 3 9 13 7 3 13 1 10 11 3 13 15 10 9 13 10 11 1 11
16 3 7 13 15 13 1 9 15 13 0 9 15 1 9 13 11
22 0 3 9 13 7 13 3 0 10 9 1 10 3 10 9 3 13 13 10 11 13 15
24 9 13 16 1 9 7 0 9 3 0 10 9 7 10 9 7 3 10 9 15 13 13 10 9
15 10 3 9 10 9 7 10 9 3 13 3 10 1 11 13
28 0 3 10 9 13 1 9 10 0 13 9 13 3 16 13 13 1 11 13 9 10 11 13 1 9 7 1 9
12 13 3 9 13 10 9 13 13 3 13 10 11
12 13 3 10 9 7 3 13 13 10 9 13 13
12 13 7 16 1 10 11 13 13 10 9 3 13
17 3 3 13 15 10 3 9 13 7 10 0 0 10 9 10 9 13
21 7 3 9 7 9 13 1 0 9 9 7 3 0 13 0 13 9 15 10 13 15
12 0 7 9 13 3 13 10 11 1 0 15 13
19 13 3 6 9 13 15 3 13 1 10 11 13 7 10 9 0 7 10 9
6 7 10 3 13 15 13
16 13 3 15 0 10 9 10 9 15 13 15 15 7 13 9 13
3 3 13 11
3 3 13 9
12 13 3 10 9 16 3 13 1 15 9 13 15
7 1 9 3 15 13 15 13
21 16 3 0 9 13 13 15 1 10 11 1 0 10 9 13 10 9 13 15 15 9
5 7 13 13 9 12
16 13 7 16 3 1 0 9 13 1 9 13 9 12 13 9 13
30 10 3 9 13 13 1 10 9 7 13 10 9 1 10 9 9 3 1 9 9 13 13 13 10 11 10 9 7 10 9
11 16 3 0 13 1 10 9 15 13 3 13
13 16 3 15 9 13 13 13 10 11 0 13 9 13
8 0 3 9 13 0 13 15 13
5 3 13 15 13 9
7 0 3 1 10 15 9 13
15 13 3 0 7 13 9 13 10 9 1 15 7 13 13 13
8 0 3 13 15 3 0 13 9
9 13 3 10 15 9 1 10 9 12
12 13 3 9 13 10 9 13 10 9 1 10 9
14 9 3 15 13 13 9 1 15 13 16 13 13 10 9
24 7 10 9 13 13 1 10 9 3 13 10 9 10 9 7 13 10 9 10 13 13 1 10 9
15 13 3 1 9 0 13 10 9 7 10 3 9 13 13 0
13 10 3 9 9 13 16 10 9 13 16 15 13 13
11 10 3 9 13 13 10 11 13 15 10 9
26 13 7 10 13 13 13 0 1 10 9 13 7 10 0 15 3 1 9 15 3 1 15 10 1 10 9
8 7 3 13 15 13 1 10 9
9 7 13 3 13 16 11 10 9 13
15 13 3 9 13 15 15 1 10 9 10 13 7 1 10 9
21 13 3 10 11 9 15 9 7 13 1 10 9 9 1 10 9 13 13 10 9 15
16 3 9 13 10 9 0 15 13 1 10 9 10 9 13 3 13
12 15 3 3 13 10 9 1 10 9 13 15 0
10 15 3 13 15 13 13 7 13 3 0
17 1 0 3 15 13 7 13 15 0 1 15 13 13 13 15 13 9
22 1 3 10 1 10 9 0 13 9 10 0 10 9 9 11 15 13 15 12 9 3 13
24 13 3 10 9 10 11 9 7 9 13 13 1 15 10 11 13 7 13 13 10 9 15 13 15
14 1 3 12 9 13 1 9 13 1 10 9 0 0 9
19 7 1 12 9 13 9 0 13 1 11 3 13 9 13 1 15 13 9 12
6 7 3 1 10 11 13
17 16 3 13 1 10 11 13 10 11 13 1 15 1 10 13 15 9
12 13 3 1 9 12 13 15 10 13 10 0 0
6 13 3 15 13 1 15
35 15 9 9 15 0 13 10 9 7 10 9 10 0 9 1 11 13 1 10 9 10 0 15 13 15 13 13 1 10 15 9 9 13 1 15
15 13 3 10 0 13 13 9 3 3 10 9 15 13 15 13
5 15 3 1 15 13
21 15 7 9 1 15 13 1 10 11 7 13 15 10 9 13 7 13 15 1 15 0
7 13 3 1 15 13 15 13
12 1 3 3 10 9 0 0 15 13 16 3 13
36 13 3 15 9 13 1 15 1 10 9 0 15 13 13 10 9 10 9 13 7 15 1 10 11 1 7 10 9 11 7 10 9 1 3 1 9
6 7 15 3 13 10 13
3 15 3 13
27 0 7 13 1 15 13 13 10 11 9 12 16 3 10 9 10 0 13 1 11 10 9 1 10 9 15 13
13 9 13 7 3 3 13 7 13 13 7 3 3 13
17 13 3 10 9 10 9 0 7 10 9 3 13 7 10 9 15 13
17 16 13 10 9 7 10 9 13 7 10 9 13 7 13 7 13 15
13 0 3 13 15 16 10 9 13 0 10 9 10 9
3 15 3 13
30 13 3 9 0 1 0 9 7 13 15 10 13 1 15 13 10 9 10 9 7 13 10 1 10 9 11 1 15 9 3
81 11 9 11 11 0 9 13 1 9 9 15 13 1 10 9 15 1 9 0 1 10 9 15 10 13 1 9 11 1 9 10 13 9 9 1 9 1 9 9 1 9 0 11 11 10 9 15 1 15 13 9 7 9 1 9 9 1 15 10 9 1 10 9 15 1 15 13 3 15 0 11 11 15 10 13 1 11 0 9 0 0
12 9 15 7 9 1 9 9 15 7 9 11 11
29 13 3 13 15 16 15 13 9 15 0 1 10 13 15 0 3 13 13 1 15 1 10 1 15 9 15 7 7 15
30 3 13 3 15 13 9 16 3 13 13 1 15 7 13 1 10 3 16 15 9 13 3 1 15 3 3 1 10 0 9
10 9 7 7 0 0 7 7 0 9 13
11 3 10 1 15 0 3 15 10 1 11 13
5 3 3 13 10 9
14 9 3 9 13 1 9 15 10 13 0 7 0 7 9
10 9 3 9 1 15 13 1 9 1 9
6 10 3 0 1 9 13
5 10 9 3 15 13
23 10 3 0 15 1 9 9 10 9 13 13 15 7 0 15 9 7 9 1 10 13 15 0
22 3 13 10 9 3 3 9 13 7 13 7 13 1 10 9 15 7 13 10 0 15 9
22 13 13 0 13 7 13 10 9 10 0 9 1 9 9 0 9 7 9 7 9 7 9
44 3 13 15 10 9 1 10 9 10 9 15 1 9 10 13 10 9 15 1 15 15 13 10 9 10 9 1 10 9 7 13 7 13 10 9 1 10 13 15 13 0 1 10 9
1 6
48 10 7 3 0 15 13 10 0 9 1 10 1 9 3 7 7 10 0 13 10 0 9 10 0 13 1 10 9 15 1 15 0 1 0 10 9 13 7 10 9 15 13 10 9 15 1 15 13
46 7 3 3 13 10 9 13 1 9 13 15 10 9 1 0 9 13 10 3 13 13 15 9 9 9 9 0 9 9 9 9 9 9 9 0 9 0 9 9 0 9 0 0 0 0 0
8 3 0 13 6 9 15 10 13
8 1 15 3 13 10 0 15 13
6 10 3 15 13 10 13
15 13 3 16 10 9 10 9 13 1 9 1 10 10 0 13
21 13 3 0 6 9 10 13 10 10 0 13 7 13 15 16 15 13 10 9 10 9
26 1 3 10 9 15 7 0 9 13 15 9 1 9 9 7 9 9 10 9 15 13 15 1 10 9 15
14 10 3 1 9 9 0 9 7 9 7 9 13 9 0
15 10 3 1 9 7 13 10 9 13 3 10 9 9 7 9
16 9 3 7 9 7 9 15 10 13 10 0 0 7 0 7 9
7 3 3 13 9 1 10 9
7 15 3 3 13 3 3 13
8 7 15 1 9 13 1 9 13
19 3 3 9 10 3 9 13 9 10 10 9 13 0 9 3 13 15 13 9
24 15 13 10 9 10 9 0 1 10 9 15 13 15 10 9 7 1 15 10 9 13 3 3 13
17 1 9 3 13 10 9 10 0 10 9 1 10 9 15 1 11 11
56 16 3 15 0 13 7 13 9 7 13 1 9 7 13 10 9 7 13 10 13 13 1 10 9 13 7 15 9 13 0 9 10 1 9 9 0 9 0 13 10 9 10 9 7 10 9 1 10 9 10 3 13 0 15 3 13
5 10 13 3 13 13
5 10 13 10 9 13
12 15 1 9 13 1 10 9 10 9 10 9 13
7 9 3 3 13 16 9 13
10 16 3 9 9 13 10 9 15 9 13
16 16 3 10 9 10 9 10 9 13 3 10 9 15 1 9 13
17 7 13 10 1 9 9 10 9 13 15 10 1 9 7 9 9 9
16 3 3 10 1 10 0 0 13 7 10 1 10 0 1 9 9
12 15 3 10 0 10 0 7 15 10 9 10 9
4 0 1 15 9
5 15 3 16 13 15
9 3 10 9 15 10 9 10 9 13
2 3 13
5 13 3 10 9 0
4 15 3 9 9
2 3 13
10 16 3 10 9 15 9 9 13 15 13
3 1 9 13
2 3 13
7 3 3 13 10 9 10 9
22 16 3 10 9 10 9 1 10 15 9 13 1 10 9 15 15 3 3 15 3 0 13
11 7 3 3 13 7 3 13 15 15 13 16
7 13 10 0 16 13 10 0
5 15 10 9 0 13
2 3 3
10 13 3 0 7 7 9 15 1 9 13
3 3 13 16
5 3 13 0 3 12
4 3 13 10 13
6 3 13 10 13 10 9
2 15 13
2 3 13
4 3 13 1 12
5 9 13 10 9 15
4 10 9 15 13
6 9 9 1 10 9 15
7 15 10 9 9 7 9 13
6 0 10 9 15 13 9
7 9 7 9 1 10 9 15
5 7 9 9 3 13
10 3 1 9 9 3 13 15 9 1 15
5 1 3 9 9 9
14 3 3 1 9 9 9 13 13 1 10 9 7 10 9
11 9 3 9 1 9 11 11 1 15 10 13
4 3 3 13 9
21 15 3 13 7 13 10 9 10 9 13 3 10 15 9 1 10 9 10 1 11 11
48 15 13 10 9 9 1 9 1 10 15 9 1 9 10 9 15 1 10 9 10 13 9 1 10 9 10 9 1 10 9 10 9 15 1 10 3 9 1 10 13 15 0 7 13 10 1 9 11
1 13
2 10 9
5 3 7 1 9 9
8 13 3 13 9 9 1 9 9
5 7 0 10 9 0
3 3 3 9
17 6 3 9 16 12 10 9 15 13 9 1 9 7 9 1 10 9
5 3 13 7 9 13
10 15 3 13 13 11 10 9 15 1 9
4 7 3 1 9
5 15 3 10 9 13
10 13 3 11 10 9 7 13 15 1 9
12 10 3 13 10 9 3 13 1 9 7 1 9
32 10 3 3 13 13 3 1 10 13 10 0 13 10 9 15 1 9 3 3 11 13 10 9 10 9 15 10 9 13 9 1 9
8 0 9 15 3 3 13 9 9
12 10 9 3 0 1 10 9 7 3 1 10 9
9 13 3 13 10 11 10 9 1 9
6 1 9 13 7 1 9
6 3 1 9 7 1 9
50 7 9 13 9 9 10 9 10 9 10 1 10 9 1 10 13 15 9 15 10 13 1 9 1 10 13 15 9 7 9 9 10 3 1 9 0 7 3 10 13 10 9 10 1 9 9 10 9 15 11
21 3 3 1 9 10 9 10 11 7 10 9 15 10 9 15 13 9 7 1 9 9
5 10 3 9 9 13
7 3 3 3 13 9 3 9
33 1 0 1 9 16 1 9 1 10 13 0 10 9 15 10 9 3 10 1 10 9 0 7 3 10 1 9 11 15 13 9 15 15
3 3 13 16
15 1 15 13 9 10 13 10 0 7 13 10 3 13 3 13
16 15 1 9 1 9 13 1 10 13 15 9 0 9 1 10 13
5 3 13 10 9 15
27 1 3 10 9 10 9 3 13 10 9 7 13 10 9 13 9 10 9 7 13 16 15 13 0 13 3 13
6 3 3 13 15 1 9
39 3 13 3 1 15 0 16 13 15 7 3 1 15 15 13 13 10 13 1 10 13 11 10 9 15 1 0 15 13 1 10 9 15 7 13 1 10 9 15
38 13 3 1 9 9 13 1 10 9 1 10 9 15 11 11 1 15 3 10 9 13 10 9 1 10 9 0 1 15 13 7 13 1 9 10 9 10 9
23 3 0 3 7 3 13 1 10 9 13 16 10 9 9 13 10 3 9 9 10 3 9 9
12 3 3 11 13 15 0 3 1 9 1 0 13
6 3 3 1 0 15 13
18 13 3 10 15 9 1 15 10 9 16 3 0 13 15 11 1 15 13
15 0 3 3 13 3 1 10 9 15 13 1 15 1 10 9
21 16 3 0 13 13 10 9 1 10 9 10 9 15 0 3 13 13 1 10 9 15
21 3 0 3 7 3 13 1 10 9 1 10 9 15 11 11 1 15 3 10 9 13
30 1 0 3 1 12 9 10 9 1 10 9 13 7 1 10 9 10 9 3 3 1 15 9 10 9 13 1 15 15 13
7 1 3 9 9 13 1 9
24 7 13 10 9 1 11 1 11 3 1 10 3 13 1 10 9 10 9 11 15 13 9 10 13
30 16 3 10 10 12 9 10 0 13 0 3 10 9 10 9 7 10 9 1 9 10 10 12 9 11 11 1 10 0 13
8 7 3 3 1 12 13 10 9
8 10 3 3 9 1 12 1 9
8 10 3 9 1 0 9 1 9
33 16 3 10 10 12 9 10 9 13 1 10 12 0 3 10 10 9 10 9 7 10 9 10 9 13 1 9 13 1 10 12 11 11
22 3 3 3 1 12 9 1 15 9 1 9 3 3 1 12 9 1 15 9 1 9 9
23 3 3 1 10 9 10 12 9 0 13 10 0 3 3 1 10 9 10 12 0 13 10 0
3 15 3 13
7 13 10 9 16 10 9 13
2 3 13
9 15 13 10 9 3 3 13 1 15
13 7 13 16 15 13 1 11 11 1 10 9 15 13
27 13 3 15 1 10 9 1 10 9 16 3 13 11 1 0 1 10 9 10 9 3 3 15 1 9 9 13
34 16 3 0 13 10 9 10 9 15 7 3 10 9 13 0 13 16 10 0 15 9 13 16 13 10 9 10 9 10 3 13 15 10 9
7 10 3 13 13 1 10 9
7 15 3 13 10 9 13 3
6 15 3 13 13 10 9
17 3 3 15 13 15 13 0 3 10 9 13 3 10 9 1 11 11
42 3 3 13 10 9 1 10 0 15 9 1 10 13 10 9 15 7 13 10 9 15 9 9 10 9 7 13 15 10 9 3 1 0 13 7 10 9 15 9 9 10 9
5 9 3 15 3 13
8 3 3 13 1 9 7 1 9
2 15 3
9 13 16 3 13 1 9 7 1 9
26 9 3 10 9 16 13 9 10 9 13 3 1 9 1 15 13 9 9 13 3 1 10 9 13 10 9
8 0 13 1 10 9 10 9 15
26 3 3 13 10 9 15 0 10 9 7 10 9 1 10 9 3 3 13 10 9 15 0 10 9 1 9
10 16 3 9 13 10 9 0 13 10 9
9 15 3 9 13 3 1 15 3 13
5 10 3 9 0 9
16 3 3 13 1 10 9 13 3 10 9 13 10 9 15 1 9
6 10 3 9 10 9 9
17 7 13 9 13 3 9 13 16 10 9 13 10 9 1 15 9 13
9 10 3 0 9 10 13 9 13 9
11 16 3 13 10 9 13 1 10 9 10 9
11 3 3 13 10 9 9 13 16 13 9 0
18 16 3 13 10 9 0 13 1 10 9 10 3 13 15 9 13 9 0
26 3 9 15 3 15 13 10 9 1 10 9 10 11 1 10 13 15 0 10 1 0 13 16 13 10 9
20 3 3 13 1 10 9 13 1 15 13 16 13 15 1 9 9 7 3 9 9
3 15 3 13
2 3 13
20 7 10 9 3 13 3 3 1 9 10 7 3 9 3 13 16 3 10 9 13
2 3 13
13 9 3 13 10 9 1 10 9 13 1 15 15 9
5 1 3 9 9 0
21 13 3 10 9 10 9 13 15 3 13 7 13 15 10 9 10 1 9 0 1 9
14 10 3 9 9 13 1 10 9 13 15 7 1 15 13
13 3 10 3 9 0 7 10 9 0 7 0 7 0
2 3 13
22 7 10 9 16 13 9 1 10 0 15 13 9 16 13 1 9 0 10 9 1 10 9
7 13 3 16 10 9 0 13
8 15 3 0 13 13 1 10 9
11 3 3 15 13 0 13 7 15 13 0 13
12 16 3 15 3 13 0 13 13 10 9 16 0
12 3 3 3 15 13 15 7 10 13 1 15 9
14 13 3 16 3 13 1 15 0 13 1 10 9 15 0
13 3 3 15 13 13 0 7 15 3 13 0 0 13
18 16 3 15 3 13 15 0 13 3 15 13 15 7 10 13 1 15 9
15 13 3 10 9 10 13 15 13 10 0 16 15 10 0 13
28 13 3 0 9 1 10 9 15 13 10 9 10 9 15 7 13 15 1 10 9 10 9 10 13 1 10 9 15
3 0 15 9
9 15 15 13 1 10 9 10 9 0
10 9 3 10 9 1 11 11 10 9 15
14 3 3 0 15 10 9 13 9 9 10 3 9 9 9
20 10 3 9 10 9 10 9 1 11 11 13 15 1 10 9 10 9 7 10 9
46 10 3 0 10 9 1 15 13 1 10 9 10 9 10 15 9 13 1 9 9 9 7 1 9 13 10 9 1 10 9 16 10 9 10 9 13 1 15 10 3 1 9 13 7 1 9
7 10 3 1 9 10 10 9
6 10 3 9 10 9 9
8 10 3 9 10 9 9 7 9
8 3 10 9 10 9 9 1 9
10 10 3 9 10 9 3 13 7 3 13
9 10 3 1 9 13 9 13 3 13
11 16 3 15 9 11 3 13 0 3 13 15
32 16 3 10 9 10 13 10 11 1 0 13 1 15 10 13 1 0 11 11 13 3 10 0 9 15 1 10 13 15 9 1 15
12 3 3 9 9 13 3 10 9 10 1 9 13
7 16 3 1 9 13 13 13
9 16 3 9 10 9 10 9 13 13
9 15 3 9 9 13 0 9 13 9
15 3 3 13 9 9 3 1 9 7 13 9 9 1 15 13
3 9 10 9
17 13 3 16 3 0 10 9 10 3 9 1 10 13 9 13 1 15
12 10 3 9 10 9 10 9 10 9 10 9 13
14 10 3 9 10 9 13 3 0 7 1 10 13 1 9
20 3 3 0 10 9 13 1 10 9 10 9 1 10 9 10 9 10 9 10 9
12 13 3 16 15 10 9 13 7 13 1 10 3
24 3 0 3 7 3 0 10 9 10 9 13 15 3 15 1 15 13 9 13 10 9 10 9 15
4 10 3 9 13
6 9 3 13 3 13 9
9 16 3 15 3 13 13 1 9 13
9 3 3 3 10 9 13 10 9 15
15 10 3 15 13 3 13 3 13 7 0 10 9 13 9 0
17 10 3 13 10 9 13 15 10 9 10 9 16 1 9 13 1 0
16 13 3 16 10 13 10 9 15 13 1 0 10 1 9 0 13
19 3 15 13 3 13 0 10 9 10 9 15 1 10 13 15 0 1 0 9
6 15 3 13 0 3 13
6 7 15 13 0 3 13
8 16 10 9 1 15 15 1 15
22 15 3 10 0 9 3 13 7 1 15 15 13 15 3 3 3 1 15 10 15 15 13
5 15 13 1 0 9
3 9 10 13
3 15 10 13
18 11 11 10 13 3 3 13 15 13 1 0 10 9 15 3 13 1 15
21 15 15 13 1 10 9 10 11 9 7 9 7 9 7 9 7 9 7 9 7 9
6 1 15 13 0 10 9
9 7 1 0 15 13 1 10 13 15
40 13 3 16 7 9 7 9 7 9 7 9 7 13 7 13 7 9 7 9 7 9 7 15 9 0 13 15 13 1 10 9 10 9 10 1 11 11 10 9 15
25 9 13 1 11 3 13 13 15 10 9 15 1 9 0 16 9 15 13 0 7 0 9 10 9 15
50 13 3 9 13 0 15 1 10 11 1 10 9 15 10 0 15 1 9 15 13 9 15 10 9 7 10 9 7 10 9 7 10 9 7 10 9 7 10 9 15 10 9 7 1 15 10 11 10 1 9
10 10 13 1 15 9 0 1 10 9 6
9 3 15 3 16 13 10 9 10 9
13 3 16 13 9 11 15 9 7 1 11 13 15 9
19 0 13 3 10 9 10 9 0 9 10 9 7 10 9 10 9 13 1 9
10 1 10 9 0 13 7 13 10 11 9
14 3 0 3 7 3 9 1 12 9 13 11 10 9 15
32 3 3 13 7 13 15 0 7 0 16 10 1 9 9 10 9 13 3 1 9 7 1 10 13 13 15 16 10 0 13 10 0
2 3 13
3 10 11 13
3 15 3 13
5 3 9 1 10 9
2 3 13
9 13 15 3 13 7 13 15 3 13
12 3 3 3 10 13 7 10 13 7 10 13 9
7 13 3 10 9 10 11 16
22 1 15 0 13 15 16 13 1 15 10 9 15 7 16 13 10 9 15 1 15 10 9
4 15 3 13 13
3 13 15 3
3 15 3 13
6 10 3 9 15 15 13
6 3 13 10 9 10 13
4 15 15 13 3
22 7 3 13 9 10 9 10 9 1 10 15 9 13 15 3 1 9 9 15 3 1 9
6 3 7 1 10 11 13
12 13 10 3 9 15 9 15 7 10 3 13 13
8 7 13 1 10 9 3 13 15
4 3 9 15 15
5 3 13 9 9 13
15 16 13 10 9 10 9 11 3 10 9 10 9 10 9 13
10 9 3 13 7 13 13 9 1 10 9
16 16 3 9 8 13 15 9 3 11 3 13 7 3 11 3 13
3 15 3 13
13 16 9 10 3 13 9 13 9 9 3 10 1 9
9 11 3 13 9 9 1 9 3 13
2 1 15
8 16 3 1 9 7 3 1 9
2 3 13
17 9 10 3 9 10 15 9 7 10 9 1 10 9 1 15 1 9
11 13 3 15 16 9 9 13 7 3 1 9
18 13 3 10 10 9 9 7 10 0 9 13 13 10 9 10 9 3 13
9 9 3 9 11 1 9 15 10 13
15 11 3 13 16 10 9 10 1 9 10 13 9 13 1 15
7 10 3 1 9 9 3 13
6 3 13 1 10 9 15
1 7
5 15 13 1 10 9
6 0 13 11 1 0 13
3 7 15 13
14 1 15 10 9 13 1 10 9 15 7 1 10 9 15
8 0 13 10 9 10 9 15 13
5 9 3 13 1 9
5 9 3 13 1 9
7 15 10 13 1 15 3 13
8 3 3 13 9 0 7 7 9
11 10 3 0 9 15 13 1 15 10 13 15
9 15 3 15 3 13 10 9 9 13
7 3 3 13 1 15 3 13
6 3 3 13 15 3 13
5 3 3 13 1 13
6 3 3 13 16 3 13
6 7 3 15 13 10 9
3 11 3 13
6 9 15 13 10 9 15
5 3 10 9 1 9
6 10 3 9 1 9 11
2 7 13
3 3 3 13
2 7 13
3 0 11 13
6 15 13 15 1 3 9
5 1 9 0 13 15
5 11 3 13 7 13
5 13 10 15 3 13
6 0 13 10 15 3 13
12 0 10 9 13 10 9 15 1 9 13 7 13
2 13 3
2 3 13
10 3 3 15 9 13 1 9 11 9 11
9 3 13 10 9 10 9 15 15 13
9 7 3 13 1 11 15 13 10 9
7 3 13 10 9 1 10 11
6 7 15 13 15 10 9
10 13 15 12 9 15 3 13 9 10 11
12 3 3 3 1 10 3 9 9 1 9 9 13
2 15 3
6 15 13 11 0 3 13
4 10 3 9 13
4 10 3 0 13
19 13 15 10 9 9 9 9 10 3 13 7 9 10 3 13 1 10 3 9
3 7 11 13
29 13 10 9 15 1 9 7 1 9 7 1 9 7 1 9 15 13 10 9 15 10 3 13 7 10 9 15 3 13
2 13 3
2 3 13
12 7 10 15 9 10 9 10 9 1 10 13 15
18 16 3 10 9 15 9 9 7 10 9 15 9 9 15 3 10 9 15
22 1 15 3 3 13 15 9 9 10 9 15 13 16 13 15 10 9 7 13 15 1 15
15 16 3 10 9 15 9 9 15 10 9 3 3 9 1 0
8 16 3 10 9 0 3 10 9
8 7 16 10 9 0 3 10 9
26 16 3 15 10 9 13 15 3 9 13 13 1 15 7 9 10 9 10 9 10 9 13 3 13 10 9
2 13 3
5 13 9 16 15 13
3 10 9 13
5 15 3 10 9 13
5 3 0 13 7 13
13 16 3 10 9 10 1 9 9 3 13 3 15 13
6 13 3 9 7 9 9
5 1 3 10 13 9
4 3 3 15 13
8 0 3 13 10 9 3 13 15
25 16 3 15 1 10 1 9 13 9 7 1 9 13 1 9 15 3 0 10 1 9 13 10 0 9
34 3 3 13 15 13 9 10 9 0 16 3 13 1 15 0 16 9 1 9 10 11 13 16 3 10 9 10 9 13 7 3 15 11 13
2 3 13
5 13 1 11 10 13
4 13 9 1 11
12 7 0 15 10 1 15 9 3 13 10 9 15
9 0 3 10 9 7 10 9 10 9
26 3 3 15 3 13 10 9 3 3 13 10 0 9 3 3 0 3 13 10 15 9 16 3 0 3 13
12 13 3 10 9 10 15 1 9 16 10 15 13
8 6 9 9 7 9 7 9 9
10 3 0 10 9 15 7 0 10 9 15
5 15 3 13 9 9
5 7 15 9 15 13
7 7 15 13 15 7 13 15
6 15 10 9 1 10 9
1 6
23 13 3 15 9 1 10 9 10 9 13 10 9 15 9 13 0 10 9 0 10 0 9 15
27 7 3 13 10 9 0 7 13 10 9 10 9 1 10 13 15 15 10 9 10 9 10 0 7 0 7 0
31 13 3 1 10 9 10 13 15 15 10 13 1 15 3 13 1 15 13 13 7 13 1 10 13 0 3 10 9 13 9 9
31 3 3 1 12 9 0 9 13 10 3 9 15 3 10 15 13 9 3 10 0 12 9 13 1 11 10 3 1 12 15 9
10 13 3 9 1 10 9 10 13 15 0
7 16 9 1 10 9 10 9
6 16 10 13 1 10 9
4 10 13 1 9
4 10 13 1 9
4 10 13 1 9
3 10 9 0
6 13 10 0 13 10 0
5 10 9 1 15 0
4 10 9 3 0
3 10 9 13
3 10 9 13
3 10 9 13
3 10 9 13
5 10 9 10 0 13
3 10 9 13
4 13 7 3 13
3 13 1 13
5 10 15 1 15 13
8 3 10 0 13 7 10 0 13
5 3 13 0 1 15
5 15 0 1 0 13
5 13 0 1 15 9
9 3 15 13 0 7 13 9 10 9
2 13 3
2 15 9
2 13 9
8 7 16 13 10 0 15 13 15
4 16 13 13 15
10 0 3 13 9 9 13 1 10 9 15
5 15 9 9 13 13
8 3 3 13 9 3 3 1 9
7 10 3 13 1 9 13 13
10 3 10 13 10 9 10 10 9 9 13
12 10 3 9 3 13 9 10 0 9 7 10 0
6 13 3 3 13 10 9
8 10 0 13 7 13 9 1 15
6 16 3 10 0 13 13
6 3 3 3 10 9 13
4 9 3 9 13
7 9 1 9 10 10 0 13
13 3 9 13 3 0 1 10 9 7 3 1 10 9
8 9 3 9 13 1 15 0 13
4 13 15 10 9
5 10 10 9 10 9
5 10 10 9 10 9
5 10 10 9 10 9
8 15 15 13 3 3 10 15 13
7 10 3 13 10 0 9 13
28 10 3 3 13 3 13 3 13 3 13 7 3 15 0 9 1 10 9 0 13 1 10 13 10 3 15 3 15
5 9 3 9 10 9
9 3 3 3 15 10 9 3 16 13
3 10 9 13
4 10 3 9 13
6 13 3 10 9 10 9
6 13 3 10 9 10 9
17 3 1 9 3 13 3 9 7 9 3 9 7 9 3 9 7 9
14 7 13 10 9 11 11 7 10 9 9 3 13 1 9
5 10 3 13 9 13
7 10 13 10 3 13 3 13
8 10 3 3 13 10 13 3 13
5 10 9 3 15 13
7 15 15 13 10 13 0 9
6 10 0 9 13 7 13
2 13 3
6 13 3 10 9 13 15
5 15 3 13 15 9
6 0 1 10 0 9 13
6 10 13 10 9 9 13
5 7 10 13 9 13
4 13 3 10 9
11 7 10 3 13 9 3 13 7 13 10 9
9 15 3 15 15 13 7 15 15 13
7 16 7 3 13 10 9 13
13 1 0 3 11 13 7 13 16 7 0 7 13 13
7 15 3 15 13 10 9 15
8 7 3 15 15 13 10 9 15
7 15 3 13 10 9 10 9
2 13 3
2 13 15
3 13 9 16
10 3 3 0 15 1 15 9 13 10 9
12 7 0 13 3 10 3 13 9 10 9 7 9
11 13 7 13 1 9 11 16 15 0 1 15
9 3 3 10 13 15 0 13 0 0
12 16 3 1 9 10 9 15 13 3 1 9 13
10 3 10 9 15 0 13 1 15 11 13
6 3 13 3 15 10 0
14 10 3 1 0 13 10 11 0 10 9 7 0 10 9
13 3 3 10 10 9 13 7 10 10 9 10 1 15
11 15 3 0 7 0 10 9 10 1 9 13
15 0 10 3 13 9 7 13 9 7 1 15 10 9 15 13
10 15 9 15 13 1 15 13 1 10 9
8 0 10 3 13 15 1 15 13
10 10 3 13 16 13 13 16 3 1 9
14 13 3 15 10 0 10 9 10 0 13 7 3 15 13
10 0 15 10 3 13 1 10 0 1 9
7 3 3 10 11 3 15 13
8 10 9 10 13 15 13 1 15
21 15 3 13 1 10 15 9 13 16 1 10 9 7 1 10 9 10 9 10 9 13
33 10 3 9 10 9 7 10 9 13 15 10 15 13 1 15 1 11 11 16 3 1 12 9 13 10 9 7 9 10 9 15 11 11
13 3 13 15 3 3 10 11 13 15 1 9 10 9
2 3 13
11 1 0 13 15 1 9 7 10 9 15 13
3 7 3 13
6 13 9 1 10 9 15
12 13 15 10 9 10 9 7 13 15 15 10 9
4 7 3 9 13
10 13 10 9 10 11 7 10 13 13 9
25 10 3 9 10 9 13 15 15 9 7 9 1 10 13 1 10 13 15 1 10 9 1 9 9 0
23 13 3 9 15 3 0 15 1 15 16 7 0 0 13 9 13 15 10 9 13 3 15 13
44 3 3 13 15 1 9 3 13 15 1 10 9 10 13 15 1 10 9 1 10 13 15 9 11 11 1 10 9 13 10 9 10 9 16 13 10 9 10 9 0 13 1 9 0
11 13 3 10 9 1 11 11 10 1 10 9
40 3 3 13 15 13 15 3 13 11 1 15 1 9 9 9 7 9 1 9 9 7 9 1 9 9 9 16 15 1 11 7 3 1 10 11 13 10 9 10 11
3 7 3 13
11 15 3 13 1 15 13 7 15 3 13 13
41 3 3 3 9 13 1 10 9 0 9 3 13 10 13 1 15 1 0 9 16 3 13 1 10 9 13 3 13 13 15 7 1 15 13 3 16 15 0 1 9 13
8 3 3 13 1 11 13 10 0
16 13 3 11 7 9 9 15 13 1 10 0 10 0 10 1 11
6 13 3 7 9 13 15
15 16 3 10 0 15 13 10 9 13 3 1 10 0 13 15
14 0 3 13 7 13 15 10 9 0 13 1 15 1 9
56 13 3 15 9 1 10 9 15 11 11 7 1 10 9 10 9 13 15 1 10 9 1 15 1 10 9 16 13 1 10 13 1 10 11 7 10 9 15 10 1 11 0 10 0 13 16 13 1 9 1 15 1 9 9 13 15
1 6
31 13 3 15 9 10 9 15 13 9 10 9 10 1 9 16 15 13 1 9 3 10 0 7 13 15 1 15 3 15 13 9
9 3 3 15 9 0 13 7 15 0
37 13 9 7 9 10 0 15 1 11 11 15 1 10 9 15 10 15 9 13 15 3 15 0 13 7 3 15 10 9 10 9 7 10 1 9 15 9
12 13 9 10 0 15 15 13 9 10 9 1 11
7 13 11 15 0 13 1 15
23 13 9 7 9 10 0 15 7 0 15 15 13 0 1 10 9 15 7 1 15 13 1 11
6 13 9 10 0 1 11
5 13 10 1 10 9
5 13 9 10 0 15
9 13 10 1 10 9 10 13 1 9
8 13 9 7 9 10 13 1 9
9 13 9 10 0 15 0 13 1 9
12 13 9 10 0 1 9 7 10 9 15 7 15
11 13 9 9 9 9 9 7 10 1 15 9
5 13 15 1 9 0
7 13 15 10 9 15 10 11
22 13 3 15 9 13 10 10 9 7 10 9 1 10 9 13 15 13 13 7 13 1 15
24 10 3 0 10 9 15 11 3 13 7 10 15 9 7 1 10 9 7 9 13 10 9 10 0
7 10 3 15 9 1 15 13
4 1 15 3 13
13 13 3 15 0 13 1 10 0 0 3 1 10 0
14 10 3 9 10 9 13 10 9 1 10 9 15 1 9
10 13 15 15 11 10 13 10 9 1 9
10 13 15 11 10 0 15 7 0 10 9
11 13 15 9 10 9 10 9 7 9 10 9
54 10 3 13 15 13 1 10 9 15 7 10 9 11 11 1 9 9 9 0 13 13 3 3 1 7 9 0 1 9 10 0 9 1 9 9 1 15 10 9 13 0 0 9 1 11 11 15 10 9 1 10 9 10 9
1 6
43 11 0 9 11 11 1 9 9 7 11 10 9 10 9 10 9 10 13 1 11 13 1 11 11 0 0 1 15 10 13 10 9 10 9 15 11 11 1 15 9 15 7 15
12 9 15 7 9 1 9 9 15 7 9 11 11
15 15 3 13 15 1 9 0 1 10 9 10 9 15 11 11
35 13 3 15 9 1 10 9 10 9 15 11 11 16 10 15 13 15 7 3 13 1 15 9 13 3 13 1 10 0 9 7 1 10 0 9
15 13 3 15 1 15 9 15 1 10 11 16 9 1 15 13
7 13 3 0 16 0 15 13
4 15 3 13 11
3 15 3 11
3 15 3 11
3 13 10 11
11 3 11 13 1 15 7 1 10 9 11 13
6 13 3 3 10 11 9
7 0 3 13 16 15 0 13
19 3 3 13 15 11 13 7 13 3 1 9 9 16 3 13 10 9 10 11
11 10 9 3 10 10 9 10 3 13 9 13
7 10 3 13 15 9 9 13
11 13 10 9 10 0 7 10 9 10 0 13
2 3 0
2 3 9
8 3 13 10 9 10 9 10 9
27 16 3 1 10 9 10 9 3 13 10 9 1 10 9 10 9 13 10 9 1 10 9 10 9 13 10 13
34 16 3 0 9 13 7 9 9 13 15 3 13 11 13 0 3 9 9 3 9 15 3 10 0 0 7 7 9 11 9 9 7 9 9
17 3 10 0 10 9 0 10 9 13 7 10 0 10 9 0 10 9
50 7 10 0 10 9 13 10 9 16 13 10 0 7 10 0 10 9 13 10 9 16 13 10 0 7 10 0 10 9 7 10 13 13 10 9 10 3 13 16 10 13 13 16 3 13 15 9 1 10 9
28 1 15 3 15 13 1 11 11 15 13 9 15 1 9 9 7 7 9 7 9 16 3 13 10 13 1 9 13
19 3 15 13 1 15 9 13 3 1 9 9 7 9 13 15 10 9 10 9
14 3 3 13 13 15 1 15 3 3 11 11 3 0 13
6 9 3 13 1 10 0
14 9 3 3 10 9 0 7 10 9 10 9 0 10 13
18 7 13 9 9 1 9 10 13 15 13 10 9 1 10 9 1 9 15
10 16 3 13 3 3 10 9 10 9 13
3 7 3 13
21 15 9 3 13 7 9 3 13 7 1 9 9 3 13 15 13 10 9 10 13 15
8 15 3 13 10 9 1 10 9
10 10 3 9 15 13 3 10 9 10 9
13 3 3 10 10 9 15 13 3 3 10 9 10 9
23 15 3 3 10 9 10 9 13 7 10 9 10 1 10 9 16 13 10 1 10 9 13 15
10 0 3 9 3 13 10 10 9 10 9
11 9 3 15 13 7 3 13 13 16 3 13
5 10 3 0 13 15
5 0 3 1 15 13
8 15 3 13 9 9 15 13 15
5 15 3 9 11 13
5 9 15 13 3 9
5 7 3 3 3 13
4 3 3 0 13
14 3 3 1 15 9 7 9 3 0 13 7 1 9 13
15 3 3 13 15 15 3 13 11 0 3 15 11 3 9 13
4 15 3 13 11
4 15 3 13 11
10 9 1 15 13 3 0 3 10 9 13
13 3 7 10 13 13 15 7 10 13 7 10 13 9
8 10 13 3 7 10 13 12 13
10 0 3 10 0 9 13 1 10 0 9
4 9 3 13 0
5 9 9 9 9 13
13 1 10 9 10 9 10 13 15 3 0 9 9 13
3 0 3 13
5 0 3 13 3 13
19 16 3 15 13 1 10 9 9 9 9 0 9 9 9 0 10 9 0 13
4 10 3 9 13
14 3 1 9 13 7 0 10 9 15 13 10 9 15 13
9 16 15 10 9 13 15 13 9 13
6 16 15 10 9 13 13
8 15 3 13 3 3 3 1 9
14 3 13 16 9 9 13 7 10 9 10 9 13 1 15
11 16 15 10 9 10 9 13 13 0 10 9
16 16 15 13 0 13 1 15 1 10 9 0 0 13 16 13 0
11 10 3 9 10 9 0 9 1 10 9 13
2 13 3
8 10 13 10 0 1 10 9 15
2 7 3
9 9 13 10 9 10 0 16 13 0
5 3 15 13 1 9
2 15 15
3 11 3 9
11 3 15 13 9 3 9 11 7 9 9 9
10 3 0 13 1 10 9 16 0 15 13
13 15 3 1 0 13 16 1 15 13 7 1 0 9
4 7 7 15 13
9 15 3 15 13 7 3 1 0 13
24 3 3 1 9 15 13 16 3 13 10 9 15 7 13 10 0 10 9 7 13 10 9 10 9
9 7 3 10 9 13 0 1 10 9
4 15 3 15 13
6 15 3 13 15 3 13
9 16 3 7 13 15 13 3 3 13
3 3 13 13
2 3 13
9 7 6 3 13 16 3 15 15 13
2 13 3
18 10 9 15 10 9 0 13 3 0 16 9 13 10 9 7 9 7 9
5 15 3 0 1 11
2 15 0
3 15 3 0
2 15 0
20 1 10 3 9 7 13 7 13 7 13 7 13 7 13 7 13 13 10 0 9
2 13 13
2 13 13
2 13 13
11 3 13 15 13 0 7 3 9 15 0 13
11 16 3 12 9 13 1 11 7 3 0 9
10 1 3 11 11 1 10 9 15 15 13
3 9 15 13
31 1 0 0 13 15 11 15 13 15 9 0 7 0 1 9 15 15 13 10 9 15 10 1 11 11 3 3 1 15 9 13
9 3 3 13 3 15 1 15 13 15
19 13 3 3 1 15 16 10 9 13 7 13 3 10 9 10 13 7 10 9
11 3 3 1 9 10 9 10 9 7 1 9
11 1 9 13 1 15 7 1 9 9 7 9
19 3 13 1 15 9 7 0 9 15 3 1 10 9 16 9 15 10 9 13
56 15 3 3 13 10 9 13 3 10 9 3 13 3 13 10 3 0 13 1 10 9 10 9 11 13 15 7 10 15 9 1 10 9 10 9 15 11 13 10 0 10 11 1 9 10 9 16 10 9 13 1 10 9 10 9 11
5 3 0 10 9 15
9 3 13 16 0 9 0 10 9 13
11 13 10 0 9 16 13 0 9 3 13 0
7 3 3 10 9 15 13 11
18 3 13 3 1 9 0 7 1 9 9 7 9 7 1 0 9 7 9
14 3 3 10 9 10 9 0 7 10 9 7 9 7 9
26 3 3 13 15 3 13 16 15 9 13 13 9 7 9 7 9 7 0 7 9 7 0 10 0 7 13
6 15 3 15 10 3 13
5 3 10 3 15 13
6 10 3 3 10 9 13
6 13 10 0 1 15 0
17 13 15 15 9 13 1 10 0 13 1 10 0 7 3 1 10 0
9 7 3 13 16 10 0 10 9 13
2 3 0
13 0 3 3 9 16 13 10 13 1 10 9 0 13
4 1 9 15 13
15 3 3 13 1 15 15 0 15 13 13 1 0 10 9 15
9 7 9 1 9 13 7 0 1 0
11 3 3 3 9 15 13 16 9 13 1 15
5 1 15 3 3 13
5 1 15 3 3 13
9 7 3 13 16 0 9 9 3 13
2 3 13
23 7 9 7 9 7 9 7 0 7 9 7 9 7 9 3 9 3 0 3 0 9 9 13
4 7 0 15 13
2 7 13
2 7 13
16 7 13 1 10 9 10 9 11 11 7 1 10 9 10 9 15
7 15 15 13 7 3 15 13
8 10 3 9 7 0 7 0 13
14 10 3 9 3 10 9 7 10 9 7 10 9 10 9
14 10 3 9 7 10 9 13 7 15 13 1 10 9 15
9 3 13 16 10 9 15 9 11 13
9 13 3 10 9 10 11 13 9 9
2 3 13
11 7 3 13 16 10 13 10 9 12 9 13
8 10 3 13 10 9 12 9 13
10 15 9 15 3 13 9 1 10 9 13
8 10 3 13 1 10 0 9 13
22 7 3 13 16 10 9 15 9 10 1 15 0 9 13 15 13 1 9 7 3 13 15
3 13 3 9
8 13 3 10 9 1 10 9 15
4 1 3 15 13
15 1 3 10 9 0 10 15 9 13 7 0 10 0 9 13
7 10 9 10 9 10 9 13
10 10 9 10 0 9 3 13 7 10 9
13 3 3 3 10 9 10 0 9 3 13 7 10 9
30 3 13 15 3 3 3 1 0 1 9 16 13 10 9 7 3 1 10 15 13 16 3 13 15 10 11 1 10 9 15
8 0 3 13 1 9 3 1 9
8 13 3 15 9 13 3 7 15
7 13 3 10 0 7 10 9
7 0 15 16 13 3 3 15
5 16 3 3 13 13
29 10 3 13 13 3 15 7 10 9 9 1 9 3 13 16 3 3 13 13 0 7 10 9 13 7 9 9 3 13
8 10 3 0 13 15 3 10 9
15 16 15 9 9 13 0 7 0 13 13 1 15 3 13 15
17 7 9 16 15 13 9 0 7 0 13 13 1 15 3 13 10 9
7 3 3 10 9 15 0 13
4 3 3 0 13
6 16 3 10 0 13 13
10 3 13 10 9 7 10 9 1 10 0
8 15 3 13 9 16 10 9 13
8 7 15 13 9 16 10 9 13
7 7 3 1 10 9 15 13
2 3 13
4 1 9 13 15
2 3 13
13 10 9 15 13 7 10 9 15 13 7 9 9 9
9 0 1 10 9 15 13 1 0 13
3 3 15 13
8 7 16 3 13 0 13 3 13
7 3 10 0 13 9 13 11
2 9 13
4 3 13 9 9
10 0 1 15 13 9 1 0 13 1 9
8 1 3 10 9 9 9 3 13
9 9 3 13 3 13 1 9 0 13
2 13 9
3 13 1 9
3 3 13 9
6 16 3 3 13 3 13
7 7 16 13 10 9 3 13
7 9 3 10 9 13 10 0
4 15 3 15 13
3 0 3 13
7 13 3 10 9 10 9 0
5 13 3 15 0 13
10 10 0 13 10 10 9 3 13 10 9
13 10 3 13 13 10 10 9 3 13 10 9 7 13
6 7 10 9 7 10 9
15 10 0 13 10 10 9 16 13 0 7 10 9 7 10 9
11 10 3 13 13 10 10 9 3 13 10 9
22 0 3 1 10 15 0 0 13 3 16 9 15 13 7 1 10 0 7 0 10 9 3
2 3 13
1 13
31 15 3 13 1 10 9 15 0 3 13 9 9 3 13 1 10 0 9 7 0 13 1 10 0 9 13 10 15 9 3 13
15 3 7 10 13 10 15 9 3 13 7 10 3 13 0 13
9 9 13 1 15 9 13 10 9 15
13 16 3 13 10 9 0 13 15 13 13 0 1 9
10 0 3 13 16 3 13 1 10 15 9
7 13 3 3 15 9 9 13
4 10 3 9 13
10 16 15 13 13 15 3 13 3 13 13
10 16 3 15 13 10 9 0 13 1 15
19 1 10 9 3 10 0 13 16 15 9 1 9 7 16 15 9 3 3 12
46 7 3 16 13 13 9 7 1 9 7 1 9 3 13 9 0 7 9 0 7 15 12 9 10 9 1 15 10 15 7 15 1 15 7 12 9 11 11 1 15 10 15 7 15 1 15
6 7 3 1 15 10 9
18 15 3 10 9 1 3 10 9 3 0 13 7 10 9 15 0 13 13
9 7 16 13 13 7 16 3 13 13
23 16 3 15 13 15 10 13 9 1 9 13 3 10 9 15 0 13 13 1 10 10 0 13
14 13 3 10 13 1 10 15 9 10 9 1 15 11 13
15 3 3 13 1 10 9 7 13 15 10 9 13 1 11 13
20 3 16 9 13 10 9 15 3 3 13 9 1 10 9 16 3 10 9 15 13
3 3 13 0
3 3 13 9
8 3 10 9 15 15 13 1 9
9 16 0 3 13 9 7 3 15 13
8 10 15 9 10 15 13 13 0
7 3 3 13 9 13 7 13
19 3 3 13 9 9 9 13 3 3 10 0 9 7 10 9 10 9 7 11
10 7 0 15 7 11 3 13 9 3 13
5 15 13 0 9 3
12 7 15 13 9 7 1 10 9 10 9 3 13
12 3 1 9 0 13 7 3 10 9 0 3 13
6 1 3 10 11 9 13
6 3 10 9 13 10 9
5 7 1 15 3 13
18 1 15 3 13 16 13 1 9 10 13 13 7 10 13 1 9 10 13
13 16 15 15 10 0 13 0 16 15 15 10 0 13
18 7 3 13 10 9 0 7 15 13 16 3 15 9 13 10 9 10 11
19 3 13 16 10 10 0 13 10 1 10 9 13 10 10 9 13 10 9 13
13 3 7 10 9 13 10 10 9 13 1 10 9 13
6 15 3 3 13 15 0
6 0 3 15 3 13 3
5 10 9 15 15 13
7 16 3 13 3 13 15 9
7 6 3 15 13 16 3 13
7 16 3 0 0 13 9 13
5 16 3 0 9 13
6 15 3 15 13 10 9
16 16 13 0 13 10 9 1 10 3 13 10 9 15 1 10 9
9 7 13 10 0 3 0 16 0 13
16 10 1 9 3 1 9 3 13 0 1 9 16 10 1 9 13
8 13 10 0 0 16 10 0 13
8 10 15 13 15 16 3 15 13
10 15 3 13 1 10 9 16 9 15 13
15 3 13 16 10 1 9 13 15 3 13 12 3 13 10 9
4 3 13 16 13
16 15 3 10 13 15 13 0 3 3 16 0 9 13 15 3 0
6 3 13 3 3 9 13
48 3 13 3 15 13 9 16 10 9 15 15 1 10 9 13 7 15 1 10 9 13 7 15 1 10 11 13 1 10 9 7 1 10 9 7 15 10 0 0 9 13 7 15 10 0 0 13 9
6 13 3 1 0 13 9
6 10 9 3 13 10 11
9 7 3 1 10 0 15 13 10 9
5 13 3 1 10 0
16 0 3 9 15 13 1 10 3 13 15 9 0 3 3 0 13
6 7 9 13 3 15 15
12 7 13 3 15 15 13 7 13 12 9 12 9
13 7 13 10 9 3 15 15 13 7 1 10 9 13
11 7 13 3 15 15 13 7 13 1 10 9
5 0 3 3 13 0
12 13 3 1 9 15 1 15 10 9 10 9 13
7 3 10 13 13 13 3 13
7 9 15 3 13 3 3 0
23 0 3 10 9 15 3 13 15 13 1 15 13 7 13 1 10 9 3 10 9 10 13 13
3 3 0 13
4 13 15 15 13
13 10 9 10 9 15 13 3 9 10 9 10 11 13
11 10 9 15 13 3 9 10 9 10 11 13
8 3 12 9 12 9 10 0 13
8 10 3 15 1 10 12 9 13
5 13 10 11 1 9
9 3 10 13 10 9 9 10 9 13
5 7 16 9 15 13
9 7 16 15 13 9 7 3 9 13
8 3 13 3 15 9 10 9 13
8 3 13 9 9 13 7 9 9
8 3 13 9 9 13 7 9 9
4 7 13 10 9
4 3 0 15 13
6 15 13 7 3 15 13
11 15 10 1 9 13 13 15 13 1 10 9
9 10 9 3 10 9 7 10 9 15
19 16 15 13 15 10 0 7 13 13 15 10 13 15 13 15 13 1 10 9
17 16 3 15 15 13 0 0 13 3 13 1 0 10 13 7 10 9
10 9 3 13 3 10 15 7 0 10 0
9 3 3 10 9 15 13 1 0 9
13 7 3 13 7 13 7 15 13 15 1 9 9 13
28 0 7 0 13 7 9 7 10 9 10 9 3 3 15 15 15 13 3 13 10 15 0 7 10 10 0 16 13
14 13 3 15 16 15 15 13 7 3 13 15 10 9 13
12 13 3 15 13 16 15 9 10 9 10 11 13
5 9 3 9 10 9
6 9 3 10 11 10 9
12 15 9 13 7 13 1 9 13 13 10 9 15
8 12 3 13 7 10 0 10 13
7 16 3 3 13 9 3 13
9 16 3 0 9 10 13 7 13 13
6 10 9 3 9 9 13
10 3 3 13 9 1 9 7 9 1 9
13 7 3 3 13 9 1 10 9 7 9 1 10 9
13 1 0 13 10 9 9 13 1 10 9 1 10 9
14 3 3 10 9 1 10 9 3 3 10 9 1 10 9
6 10 3 15 1 10 9
4 1 15 15 13
7 13 13 9 0 10 9 13
7 3 10 9 1 9 13 15
16 16 3 15 13 0 13 15 0 9 3 13 7 10 9 10 9
15 0 3 13 3 13 16 3 1 10 0 7 1 10 0 13
14 13 3 3 9 1 15 13 16 10 0 0 13 1 15
11 13 3 15 1 10 15 3 13 0 9 13
16 0 3 10 0 9 13 1 10 13 7 15 3 13 15 3 13
10 3 3 9 3 13 1 10 13 7 13
11 7 10 9 10 9 13 7 13 10 3 13
2 13 15
4 1 0 3 13
8 0 15 13 10 9 10 1 15
6 0 13 1 10 15 9
8 3 3 10 9 1 10 13 13
11 0 10 9 10 0 9 13 1 10 15 9
9 0 13 3 3 13 1 10 15 9
19 3 3 3 13 10 9 0 7 10 9 13 10 9 10 9 13 16 15 13
15 13 3 9 15 7 3 1 10 9 13 7 1 10 9 13
11 1 0 1 15 0 0 7 0 7 13 0
7 16 3 15 13 3 3 13
12 13 3 1 10 9 13 16 3 1 10 9 13
9 3 9 15 13 1 10 13 15 13
11 16 15 13 1 9 13 16 3 1 9 13
7 10 3 0 16 3 13 13
9 1 3 10 0 9 3 13 15 13
4 9 3 9 13
4 10 3 0 9
8 7 9 9 13 7 10 0 9
4 7 9 9 13
10 10 3 0 9 10 13 10 15 1 15
10 0 3 13 10 9 10 9 1 10 13
9 15 3 3 1 10 9 13 9 9
8 0 3 9 9 1 10 0 9
8 0 3 9 9 1 10 12 9
4 0 3 9 9
3 0 3 9
4 0 3 9 9
3 0 9 9
4 0 3 9 9
15 15 3 0 13 10 12 7 10 0 9 13 0 0 3 13
25 3 3 10 9 12 13 7 9 0 13 15 3 10 9 10 9 0 13 12 13 9 3 3 10 11
21 16 13 10 9 16 3 13 9 3 13 1 10 9 3 1 0 3 13 1 10 9
22 7 16 13 10 9 16 3 13 9 3 13 1 10 9 3 1 0 3 13 1 10 9
8 16 0 10 9 9 3 10 9
6 16 0 9 3 10 9
15 3 3 10 9 13 10 9 12 0 15 1 10 9 3 13
10 16 3 13 10 15 12 9 3 10 9
5 3 3 0 3 9
22 3 13 3 10 9 13 10 9 9 15 3 13 7 3 10 9 10 9 9 15 3 13
7 10 3 0 15 3 9 13
26 7 10 9 13 10 9 10 13 0 13 9 16 3 13 9 1 10 9 7 10 15 1 15 13 10 9
9 7 16 13 12 9 13 15 10 9
7 16 13 9 13 15 10 9
9 15 3 13 9 11 7 9 1 9
24 7 15 3 13 10 9 1 10 9 0 9 0 9 0 9 3 9 3 9 9 9 9 9 9
3 3 15 9
3 3 15 9
5 3 15 9 13 9
4 3 15 9 13
3 3 15 13
6 13 3 10 9 10 0
7 7 3 1 9 9 15 13
28 7 16 13 9 7 13 10 9 15 7 15 10 9 7 16 13 15 10 9 16 9 13 9 3 3 13 15 13
21 7 16 13 15 10 13 15 7 16 13 10 9 15 16 13 9 3 3 13 15 13
3 10 9 13
2 3 13
4 10 9 3 13
2 3 13
2 3 13
2 3 13
4 3 13 10 0
5 3 13 1 10 9
4 13 3 10 9
2 15 13
2 15 13
2 15 13
4 16 3 9 13
3 16 9 13
3 16 9 13
8 1 9 3 13 7 1 9 13
9 3 3 13 10 0 10 1 9 13
3 13 3 0
3 13 3 0
7 13 3 3 1 9 1 9
5 3 3 9 1 9
4 3 13 1 9
6 3 3 13 3 3 13
9 3 3 13 9 9 9 10 12 0
5 0 3 0 10 9
8 13 3 10 0 3 3 16 13
3 15 3 13
4 9 3 13 9
10 10 3 13 9 13 9 7 9 7 9
5 10 13 9 15 13
5 10 3 13 9 13
10 13 3 15 15 13 9 3 3 16 13
17 0 3 10 13 3 10 13 9 3 16 3 13 16 10 9 9 13
11 7 3 16 0 9 9 13 15 13 1 9
15 3 3 15 1 10 9 16 3 0 9 13 3 13 10 13
5 13 3 1 9 13
11 0 16 13 9 9 13 1 9 7 15 0
18 16 3 3 13 10 9 10 9 13 10 13 0 7 10 13 1 15 0
15 3 3 15 16 9 13 9 1 10 9 10 9 13 16 13
7 3 10 13 9 13 16 13
8 16 3 13 9 10 9 15 13
3 15 3 13
3 13 10 9
5 13 3 3 10 9
3 13 10 9
5 13 3 3 10 9
23 3 16 13 9 10 13 10 9 10 9 3 13 10 6 1 10 15 9 16 15 13 3 13
10 15 3 3 3 13 7 10 0 3 13
3 13 10 9
10 9 3 9 13 10 9 7 10 9 13
5 10 3 9 0 13
22 1 10 9 13 16 1 0 7 1 9 0 13 10 9 0 7 3 3 13 15 13 9
12 3 10 9 1 9 13 3 10 13 7 10 0
9 10 3 9 3 10 0 7 10 13
22 16 3 13 10 9 0 1 10 15 7 15 13 9 13 3 9 7 0 3 13 16 13
13 16 3 15 13 13 3 15 0 3 9 13 1 15
22 10 0 10 9 15 0 13 7 3 13 1 9 13 10 9 13 16 3 9 1 15 13
5 3 13 0 9 13
2 9 13
2 9 13
2 9 13
2 9 13
4 15 1 9 13
8 16 3 3 13 9 13 1 9
6 15 3 13 7 10 9
8 16 3 0 13 13 10 0 13
17 13 3 1 12 15 13 16 15 13 7 15 13 7 9 9 9 13
8 3 3 13 9 10 9 7 9
13 3 1 15 10 9 10 0 10 9 1 10 9 13
5 3 3 13 15 13
11 16 3 15 13 13 1 9 10 0 9 13
7 0 3 13 9 13 1 9
13 7 1 15 10 9 10 9 13 7 1 15 0 13
5 16 3 15 13 13
12 3 9 15 13 10 13 7 10 13 3 13 9
7 15 3 3 7 1 9 13
31 13 3 15 9 10 9 15 13 15 15 7 13 1 15 7 13 1 15 7 13 15 9 13 15 16 13 3 16 3 3 13
16 3 13 1 12 9 3 1 15 10 0 13 1 3 15 3 13
3 3 13 11
4 3 10 9 15
9 0 3 15 3 10 9 13 3 15
31 9 3 9 13 15 13 7 10 9 15 10 1 15 3 0 13 7 0 15 15 13 3 15 3 7 10 9 10 9 1 15
10 7 3 15 7 0 3 13 7 3 13
18 16 3 11 13 16 13 1 0 3 13 1 15 15 16 9 0 3 13
16 16 3 11 3 13 0 3 7 10 9 15 0 7 10 9 15
23 13 3 7 9 10 9 16 13 1 10 9 16 13 10 11 15 3 13 16 3 0 3 13
8 16 3 0 3 13 3 11 13
9 16 3 11 3 13 0 10 9 15
6 3 13 1 10 9 15
14 16 1 10 9 0 1 11 13 13 0 0 15 9 13
9 3 3 11 13 1 0 9 10 13
14 3 3 1 10 11 15 13 3 3 1 10 11 15 13
6 0 3 1 10 0 9
2 9 11
8 3 15 10 11 1 10 9 15
20 3 10 9 3 13 10 9 10 9 7 9 3 13 15 9 7 15 9 7 9
14 13 3 15 13 16 15 13 15 10 0 1 10 9 15
7 15 3 13 1 10 9 15
25 3 3 13 15 10 15 3 3 0 10 9 13 10 13 15 10 15 16 13 10 9 10 15 1 15
8 3 15 13 10 13 1 10 0
10 16 3 0 3 13 15 3 13 1 15
6 15 3 15 13 15 9
16 1 9 13 3 10 15 9 9 15 13 1 11 11 10 9 15
10 16 1 9 13 1 11 15 15 10 9
7 16 0 3 13 13 7 13
5 13 9 0 9 0
5 13 3 7 3 13
5 9 3 9 15 13
4 1 9 15 13
3 7 13 15
4 3 13 10 0
4 15 3 9 13
9 0 15 15 13 3 13 16 3 13
14 10 3 9 13 15 9 3 13 7 0 10 9 0 9
21 3 15 9 10 0 9 7 0 3 9 0 3 9 9 0 3 9 0 0 3 9
6 7 9 0 7 9 0
7 7 0 3 10 10 0 9
5 0 3 10 10 0
11 0 9 9 7 0 9 9 7 0 9 9
6 9 3 9 13 1 9
6 3 3 10 9 10 0
3 13 1 9
3 13 1 9
3 13 1 9
3 13 1 9
3 13 9 0
3 13 9 0
7 16 13 9 0 13 3 0
8 13 10 0 9 11 1 9 13
8 7 3 0 10 0 7 10 0
3 3 10 0
6 10 0 9 1 9 0
5 10 0 9 1 9
15 15 10 0 0 3 10 0 7 15 10 0 0 3 10 0
13 7 3 13 10 9 10 0 13 3 10 9 10 0
4 6 9 15 13
3 15 3 13
10 13 3 7 10 0 13 0 7 15 13
13 13 3 10 0 0 13 9 7 10 0 0 13 9
19 3 3 10 0 0 13 9 7 10 0 0 13 9 3 13 10 9 10 13
5 13 10 9 1 9
5 3 15 9 10 9
7 10 3 9 10 9 10 9
7 10 3 9 10 9 10 9
15 10 3 9 9 10 13 15 10 9 1 10 9 15 11 11
18 1 3 10 9 10 1 10 0 3 13 10 9 10 11 3 3 15 13
20 1 12 9 0 15 1 15 13 13 15 15 3 13 16 3 3 13 3 9 13
16 3 3 13 15 3 13 1 9 0 13 13 10 9 15 1 11
11 16 3 13 0 10 3 15 13 1 15 13
3 11 3 13
15 1 15 3 13 13 7 3 13 16 15 15 13 3 3 13
8 3 13 3 15 3 1 9 13
11 13 3 9 15 13 1 15 16 10 9 13
10 9 3 15 13 0 7 0 7 13 0
10 16 3 13 11 13 16 3 13 1 15
8 10 3 9 9 13 3 3 15
9 13 3 15 1 9 16 13 1 15
6 13 3 15 1 10 9
15 1 3 11 10 9 0 13 15 16 13 1 15 1 10 9
8 7 3 3 13 9 16 3 13
4 13 3 3 13
4 13 1 10 9
1 13
5 15 15 1 9 13
32 13 3 15 9 13 10 9 11 16 13 9 10 11 7 1 9 10 0 13 15 16 3 15 13 10 0 7 15 10 13 7 13
16 13 3 1 10 9 11 7 11 7 11 16 10 15 9 0 13
8 13 3 10 15 9 7 10 15
4 13 3 10 0
6 13 15 10 9 10 11
5 13 15 10 9 15
6 10 9 10 15 9 11
8 16 15 3 13 10 9 13 9
2 8 8
7 10 9 10 9 11 1 15
9 10 9 15 1 15 15 1 11 11
29 11 9 11 11 1 9 9 7 11 10 9 10 9 10 9 10 13 1 11 1 10 0 15 10 13 1 0 10 11
12 9 15 7 9 1 9 9 15 7 9 11 11
9 16 3 13 1 10 15 9 7 9
17 16 13 1 10 15 9 10 13 1 9 10 0 9 15 3 15 13
18 7 10 9 15 0 1 15 13 16 3 9 13 10 9 3 3 10 9
27 3 3 13 15 13 9 1 10 9 15 10 13 1 10 11 16 1 9 1 9 13 16 13 15 3 10 13
23 7 0 1 15 10 9 10 9 13 16 3 13 13 1 15 7 1 10 9 10 13 10 0
35 15 1 0 9 13 15 7 13 1 15 13 16 3 3 13 13 3 15 1 15 10 9 16 1 0 9 10 1 15 9 1 0 13 1 15
34 10 3 9 15 0 13 10 9 10 9 15 16 1 9 7 9 10 9 3 1 9 0 7 1 9 9 13 1 10 9 3 3 1 15
12 3 3 0 13 15 7 7 15 13 7 3 13
33 7 0 10 9 13 0 1 15 13 16 0 9 13 7 1 15 13 1 11 7 3 1 11 13 1 15 7 1 15 13 1 10 11
8 0 3 13 3 3 10 9 13
17 7 15 13 1 9 13 16 13 1 15 10 6 6 7 10 3 3
16 0 3 10 9 16 10 9 15 10 1 15 3 13 6 7 3
29 10 10 9 3 9 11 11 10 1 15 1 15 13 1 15 7 11 7 11 3 13 6 7 3 7 6 1 15 13
8 15 3 9 9 1 15 10 6
12 3 7 1 15 10 6 10 9 1 9 1 15
26 10 3 13 15 1 15 1 11 7 13 15 9 10 3 13 15 7 13 10 9 10 9 1 10 9 15
4 10 3 9 13
12 13 3 15 0 10 3 3 1 9 1 15 13
16 16 3 15 13 15 3 15 10 13 15 3 3 10 13 1 15
25 7 13 0 15 16 3 13 9 13 1 15 13 15 13 13 1 15 15 16 10 15 9 15 15 13
25 1 3 0 9 7 9 9 13 15 1 0 9 3 16 13 7 10 9 16 13 15 13 3 1 15
15 16 3 15 13 3 15 13 7 1 9 16 3 13 15 15
25 0 10 0 10 9 0 10 1 10 0 16 10 3 3 15 13 7 13 16 10 0 9 13 10 0
15 1 0 3 3 13 16 13 10 9 15 16 1 15 0 13
19 7 3 15 15 13 16 15 13 1 15 1 9 11 16 3 13 1 10 11
6 3 3 15 10 9 13
36 13 3 1 10 11 1 10 9 10 11 3 9 15 13 1 9 3 13 9 10 9 15 10 3 13 15 11 10 9 15 7 13 15 13 1 11
23 10 3 9 9 10 3 13 15 1 10 11 7 10 9 10 9 15 13 1 15 1 15 9
13 3 11 9 13 10 9 1 10 13 7 1 10 13
7 15 3 9 1 9 1 9
5 7 1 0 15 0
15 3 3 13 3 10 0 13 10 9 10 9 7 3 1 9
4 13 3 15 13
12 7 3 13 3 15 0 9 1 15 7 1 15
16 10 9 15 15 13 13 1 10 9 15 13 7 13 1 15 9
24 13 16 13 9 11 13 1 15 13 3 9 7 9 9 13 3 1 9 0 7 1 9 9 0
10 9 3 0 13 1 10 11 1 10 9
4 10 3 9 13
4 10 3 9 13
42 16 3 10 9 10 9 1 9 13 9 13 1 9 16 3 13 13 10 9 11 1 10 9 11 1 10 9 10 9 15 10 13 3 3 3 10 9 10 9 13 1 9
14 7 3 3 13 10 13 1 0 10 9 1 10 13 9
12 16 3 10 13 1 9 0 3 10 13 1 9
29 13 3 0 9 0 9 13 7 3 3 11 13 9 1 10 9 15 1 10 3 13 10 9 11 1 10 9 10 13
5 7 13 10 9 15
13 7 1 3 16 3 13 11 9 1 10 9 15 13
9 16 3 3 13 1 9 13 10 9
6 10 3 9 10 9 13
6 3 3 10 9 9 9
40 1 0 13 10 9 0 3 13 3 13 7 13 10 0 10 9 3 13 1 9 7 13 10 9 10 9 7 10 9 10 9 13 15 1 15 9 9 1 10 9
42 16 3 3 13 13 10 9 15 1 10 13 13 13 1 15 10 9 10 9 0 13 10 9 10 0 1 10 3 13 10 9 10 9 10 9 10 11 15 13 9 10 9
8 3 3 15 13 7 11 11 9
26 3 10 9 10 13 1 9 9 13 15 13 1 10 9 15 1 9 10 9 10 9 10 9 1 9 11
20 13 3 10 9 0 1 0 9 16 10 9 10 9 13 10 9 7 3 1 15
38 1 15 13 7 3 13 13 7 3 13 13 7 3 13 13 7 3 13 3 10 9 10 11 1 10 9 13 16 3 10 9 10 11 1 10 9 15 13
22 3 3 15 10 13 1 9 13 1 11 16 3 10 9 10 11 13 1 10 0 9 15
6 3 10 9 1 15 13
36 13 3 10 0 9 10 9 1 10 13 13 3 7 13 3 15 13 3 7 13 13 16 10 13 10 9 11 3 15 1 11 13 7 13 1 15
20 10 3 15 1 15 16 10 9 13 1 10 0 10 9 13 1 10 9 10 9
25 10 3 3 0 10 9 15 1 9 1 9 0 9 9 13 15 3 13 15 10 13 7 10 3 13
4 10 3 13 0
5 10 3 3 13 0
21 13 3 16 16 10 0 15 9 10 9 13 9 1 9 13 9 0 0 1 10 9
20 7 3 1 0 13 10 9 15 10 1 9 13 13 16 3 7 13 3 0 13
23 7 3 10 13 1 10 9 13 13 1 15 3 13 13 7 13 16 13 10 0 1 10 9
14 13 3 3 7 13 16 13 1 10 9 13 1 10 9
14 13 3 7 13 3 13 1 10 9 7 13 1 10 9
10 3 7 13 7 13 7 13 0 15 13
25 10 3 15 15 13 13 1 10 9 10 11 16 13 0 10 1 10 9 1 15 13 7 0 7 0
8 13 3 10 9 10 9 9 13
3 9 3 13
8 13 3 3 1 10 9 15 13
24 3 3 3 15 13 15 7 9 13 15 9 1 15 16 13 1 10 1 9 13 7 3 1 9
14 10 3 9 10 11 13 15 13 0 16 12 1 15 13
4 3 10 15 13
17 7 1 15 13 16 10 13 3 15 13 7 10 1 15 13 7 13
9 3 15 1 10 3 15 13 1 9
10 16 3 13 1 9 11 7 3 3 13
7 3 16 15 1 11 0 9
3 10 0 13
3 6 13 0
10 1 11 3 13 3 10 9 13 1 15
3 13 1 11
3 13 10 9
15 10 3 13 9 1 15 9 13 16 15 13 9 9 1 15
13 13 3 3 13 3 1 0 10 9 10 9 13 15
2 13 3
10 9 0 13 15 7 1 9 9 13 15
4 6 3 9 0
17 1 10 9 10 9 10 0 7 0 1 9 7 9 1 9 7 9
34 3 0 7 0 3 13 7 13 3 13 7 6 13 3 13 7 3 13 3 13 3 3 13 3 0 0 3 13 3 15 13 7 15 13
6 10 9 15 13 1 15
5 0 10 9 15 13
4 3 13 1 15
6 13 3 1 10 9 15
10 10 3 0 9 3 9 13 13 3 15
6 15 3 9 9 7 9
12 15 3 9 11 1 11 7 15 9 0 1 0
7 15 3 9 9 9 1 9
6 15 3 9 9 13 13
5 3 13 10 9 16
14 13 1 15 7 13 7 13 15 9 7 15 13 15 9
13 3 13 1 0 15 7 13 13 9 7 0 3 13
3 13 9 9
19 0 3 13 10 9 0 13 15 1 15 9 9 7 9 13 9 1 9 9
2 15 13
2 15 13
2 15 13
4 1 9 3 13
13 13 3 16 1 10 9 15 13 1 10 13 7 13
5 0 15 9 1 15
3 13 10 9
8 13 10 9 1 15 10 9 15
2 3 9
2 3 9
13 7 10 13 10 0 13 15 10 9 1 10 9 11
33 3 0 3 1 10 9 15 7 3 1 10 9 15 13 1 15 13 15 10 15 9 10 15 9 10 15 9 1 15 16 15 3 13
10 13 3 1 9 16 1 15 13 1 15
10 10 3 1 9 9 9 1 9 0 13
7 10 3 10 9 9 9 13
24 6 3 15 0 10 1 9 13 15 13 15 9 7 9 7 9 7 9 7 9 7 9 7 9
28 3 16 3 13 15 3 1 10 13 7 1 10 13 7 1 10 13 10 9 15 10 1 15 1 15 1 10 9
3 1 0 13
20 1 3 10 9 15 3 3 13 1 10 9 11 16 13 10 9 15 1 15 15
20 7 10 9 15 3 1 15 13 13 10 15 15 9 16 1 9 7 9 13 15
7 13 16 1 15 13 1 15
38 13 3 15 9 10 9 10 9 10 13 1 10 9 10 11 16 1 0 9 9 10 9 10 9 15 7 10 1 9 9 15 13 1 10 9 10 9 15
24 3 1 9 13 7 1 9 0 1 0 9 13 15 10 9 7 10 9 10 9 10 1 10 0
32 7 3 3 13 7 15 13 0 10 9 7 15 1 9 9 1 10 13 15 11 16 3 13 3 3 13 1 15 3 10 9 0
16 3 1 9 13 7 1 10 0 9 7 10 10 15 9 0 13
21 13 3 10 9 10 9 15 11 11 16 1 15 13 0 13 16 15 10 0 9 13
16 0 3 15 13 15 3 0 10 13 7 3 10 13 13 1 3
19 3 3 3 10 13 13 16 3 10 9 10 13 3 3 10 13 1 10 13
13 16 3 10 9 13 3 3 13 0 3 3 3 13
10 3 3 16 0 9 15 9 7 1 9
24 1 10 3 9 10 15 9 1 10 0 9 16 3 10 0 9 13 1 10 15 9 16 13 9
2 3 13
27 9 3 10 9 10 13 10 0 9 1 15 1 10 9 11 16 10 3 9 13 0 3 13 0 13 1 15
42 3 0 3 7 7 13 1 10 9 9 15 1 10 9 0 10 13 1 15 1 10 0 10 9 9 7 9 15 13 0 3 15 15 13 1 10 9 0 10 13 1 15
11 13 3 0 3 0 1 9 7 3 1 9
22 13 3 15 10 9 15 15 13 1 0 3 0 13 3 3 0 0 9 0 10 1 15
9 7 1 11 9 15 7 1 15 0
7 7 9 15 9 9 9 11
18 10 3 9 10 9 15 7 15 9 1 15 1 15 13 1 9 10 9
15 1 3 3 10 9 10 1 10 0 0 15 13 10 13 15
25 0 3 13 13 10 9 16 13 1 15 7 13 10 13 9 15 0 0 13 3 3 9 3 3 9
2 0 3
15 10 13 3 3 3 13 7 10 13 1 9 1 9 3 13
11 0 3 13 10 9 3 1 9 7 1 9
6 0 3 9 13 10 9
21 13 3 10 9 15 9 13 1 15 16 1 15 3 15 9 13 13 1 15 9 0
2 3 13
1 13
7 10 9 15 13 1 10 9
23 10 3 13 9 10 13 7 9 1 9 13 7 13 10 9 15 7 13 10 9 10 9 15
13 1 15 13 1 15 9 15 13 1 15 9 10 9
22 3 10 9 10 9 0 3 0 13 13 10 9 10 0 7 3 13 1 0 9 10 9
44 1 10 9 10 9 0 13 10 9 1 10 9 10 9 15 1 10 9 10 11 7 9 10 9 1 15 7 1 15 7 15 9 1 15 13 15 1 10 13 9 10 9 1 15
8 9 10 9 1 10 0 15 9
25 0 3 15 11 13 15 1 10 9 7 9 10 11 15 1 9 3 0 1 15 13 3 13 1 15
20 13 3 10 3 13 13 10 9 15 13 13 1 15 10 13 15 3 1 9 13
18 16 15 13 15 11 13 0 13 3 1 15 16 3 15 11 3 3 15
33 16 7 3 0 15 13 1 10 9 15 15 13 10 9 1 9 7 3 1 9 15 3 13 16 3 13 3 3 13 15 1 10 9
8 3 10 9 3 13 0 7 0
10 10 3 9 10 9 0 7 10 9 13
17 0 13 10 0 16 15 13 10 9 1 9 13 0 3 13 10 9
11 3 3 13 13 7 13 15 15 10 15 13
12 7 15 1 15 15 13 7 13 15 15 3 13
9 3 3 3 3 13 1 15 13 15
37 3 1 10 0 13 1 0 9 9 3 13 13 10 9 15 1 15 13 1 10 9 15 1 9 1 10 1 15 13 3 1 0 9 1 10 0 13
6 10 3 13 1 9 13
13 3 3 10 15 13 0 13 0 7 15 10 9 13
6 6 13 15 0 15 9
4 7 3 13 15
5 13 3 15 9 9
22 13 3 16 3 10 9 13 11 1 10 9 15 13 10 9 15 1 10 9 10 1 11
26 16 3 3 10 13 0 11 13 15 3 13 7 9 0 13 15 3 13 7 9 0 15 3 13 3 13
18 16 3 3 9 10 9 7 3 10 9 7 1 15 13 1 15 1 15
16 7 9 13 15 13 16 15 13 16 3 10 10 9 9 13 15
18 0 9 13 13 9 1 10 15 9 7 13 1 15 7 13 3 13 15
10 10 3 9 15 13 10 9 13 1 11
9 7 1 15 0 15 15 13 7 13
2 1 15
4 16 3 13 15
3 10 9 13
10 10 3 0 9 9 0 13 1 9 11
3 7 3 9
8 0 3 10 11 13 1 9 9
12 3 0 3 16 3 10 9 15 13 3 9 9
2 3 13
6 3 15 15 13 0 13
15 16 3 3 3 3 3 0 13 15 16 3 15 0 15 13
16 15 13 3 1 9 13 7 3 1 9 1 0 10 9 10 9
7 3 3 13 10 0 0 13
21 13 3 16 15 15 13 16 15 13 16 15 13 16 15 13 16 15 1 9 15 13
7 1 9 13 3 16 15 13
2 0 13
2 3 15
2 9 13
2 3 15
3 9 11 13
3 9 11 13
2 13 13
12 1 9 3 1 9 3 1 9 3 1 9 3
7 1 0 3 12 1 12 13
2 3 13
2 3 13
2 3 13
5 9 1 10 9 13
14 1 10 3 10 9 15 10 1 9 10 9 15 10 9
6 15 13 7 3 15 13
8 16 13 13 10 10 9 15 13
17 10 9 7 9 10 9 11 13 10 13 0 1 10 9 16 3 13
27 1 11 10 9 11 10 9 13 10 9 0 13 15 7 1 9 1 9 13 1 10 9 7 13 10 9 15
2 13 13
3 3 13 3
7 13 3 1 9 7 9 9
4 1 10 0 13
11 1 3 15 3 13 3 3 1 10 9 15
7 16 3 13 13 3 13 0
3 9 3 13
15 13 3 3 15 1 15 13 1 15 13 15 7 13 1 15
21 7 10 9 10 9 16 3 13 13 15 9 10 9 9 11 16 15 13 16 3 13
10 1 0 3 10 9 13 16 13 1 15
3 7 13 15
6 10 3 9 1 9 13
16 3 3 3 13 1 10 9 15 16 13 1 15 10 9 10 11
14 3 13 1 9 1 9 1 9 1 9 7 9 1 11
6 3 3 13 3 0 13
2 13 0
3 15 15 13
6 15 3 13 1 15 13
10 15 3 13 10 3 9 16 3 15 13
5 13 15 10 9 0
11 6 0 0 3 13 13 1 15 7 3 13
7 3 3 13 10 15 7 15
13 3 3 13 10 9 10 9 13 7 10 9 10 9
10 15 3 3 13 7 13 1 10 9 15
6 16 3 15 13 0 13
2 13 3
6 7 13 9 9 15 13
6 13 11 7 13 10 9
4 3 13 15 11
5 3 10 0 9 13
4 3 10 0 9
5 3 13 16 15 13
5 1 9 1 11 13
28 3 3 13 15 13 15 10 9 15 1 15 7 13 0 10 13 7 3 13 1 10 9 7 9 7 9 15 13
5 0 0 13 1 15
32 13 7 13 3 13 10 0 3 13 3 10 13 7 10 0 15 16 16 13 1 10 3 3 13 16 9 13 10 1 15 13 11
9 15 1 15 3 13 7 13 1 15
10 7 3 13 1 9 7 13 1 9 9
15 3 3 15 13 1 15 7 13 1 15 1 9 9 1 15
7 15 13 16 13 1 10 9
9 7 3 13 15 16 11 11 1 15
4 16 3 0 13
9 13 3 16 13 16 15 3 13 0
11 3 3 13 15 1 10 9 7 1 10 9
9 13 3 3 15 13 15 3 0 13
6 0 7 13 10 15 9
24 1 0 0 13 13 16 13 3 3 13 1 10 9 15 10 9 13 15 1 9 7 3 1 9
1 13
1 13
3 10 15 13
1 13
5 13 15 1 0 9
5 13 15 10 0 15
20 10 9 10 9 11 11 7 10 9 10 9 7 10 9 10 0 9 1 15 15
44 9 15 7 9 1 9 9 7 9 15 11 11 10 13 15 1 10 9 15 16 13 15 1 10 9 10 13 0 1 10 9 10 9 7 9 15 15 10 9 1 10 9 10 9
1 6
33 13 16 3 3 13 1 10 13 15 1 9 11 1 0 9 15 3 13 0 16 3 15 13 10 13 15 7 13 13 10 9 10 11
15 7 3 16 15 7 9 1 9 13 1 15 13 15 9 13
6 3 13 3 3 3 13
7 3 3 9 13 7 10 9
4 7 13 9 13
15 13 3 15 9 10 9 10 13 1 15 16 3 13 1 9
14 7 3 15 1 9 13 15 7 13 7 1 9 11 11
39 13 3 10 15 9 3 1 10 9 16 1 9 13 10 9 10 9 7 13 15 7 13 1 10 9 1 0 9 1 10 9 15 3 9 13 10 0 15 9
52 16 3 13 10 13 15 1 9 9 15 7 13 1 10 9 15 13 10 9 15 1 15 16 13 15 1 10 9 3 3 13 9 7 9 7 13 1 11 1 10 1 15 9 7 13 1 11 7 3 13 1 11
15 3 1 12 9 13 1 11 13 11 7 13 1 15 9 12
13 0 3 10 9 3 13 3 3 11 10 9 10 9
10 3 13 1 10 9 10 11 7 10 11
5 0 3 13 13 16
11 10 13 15 3 3 13 10 9 15 3 13
6 7 13 1 15 10 9
13 3 1 12 9 3 13 1 11 1 11 13 3 11
4 13 3 1 9
10 7 13 15 10 9 15 13 1 10 9
11 1 0 3 10 13 16 1 0 13 7 13
15 15 3 1 9 13 10 9 16 10 9 10 9 13 1 15
12 1 3 10 13 13 15 15 3 13 15 15 13
6 9 10 9 9 3 13
66 15 3 10 13 15 13 7 10 3 13 16 13 10 9 10 9 3 11 10 9 10 3 13 11 1 9 10 9 13 7 15 1 10 9 7 13 10 9 10 13 15 11 7 11 7 11 10 13 9 13 0 13 15 7 11 9 16 15 1 10 9 15 3 1 10 9
11 0 10 0 16 13 15 3 13 0 0 13
13 16 3 13 11 1 11 1 9 15 13 16 13 13
11 1 10 3 13 15 1 11 1 10 9 13
11 16 3 13 13 7 13 15 13 10 1 9
16 7 16 13 16 3 13 1 10 9 10 9 13 10 11 1 15
14 16 15 0 13 3 7 3 3 13 3 10 9 13 13
8 15 9 0 7 3 1 9 0
39 13 3 16 3 13 9 1 9 9 3 3 1 9 11 11 7 15 1 11 11 13 16 13 1 9 11 7 3 1 9 9 16 1 9 9 3 13 15 9
14 16 3 13 13 1 11 13 3 0 0 3 11 9 9
2 3 13
10 16 3 15 13 0 3 13 9 15 13
9 15 3 1 9 9 13 16 9 13
5 13 3 1 15 11
22 15 3 3 13 1 9 1 9 13 10 10 9 10 9 10 13 15 7 13 15 1 15
6 3 13 10 9 10 9
9 16 3 1 9 9 3 11 3 13
13 6 0 9 15 15 13 15 1 9 11 11 13 13
6 0 0 13 13 1 15
10 1 9 9 10 9 13 7 1 9 9
5 13 9 3 9 13
4 16 3 3 3
18 10 3 13 15 10 9 7 13 9 1 15 1 9 9 7 1 9 9
10 3 11 13 10 9 7 13 15 1 9
10 13 3 16 10 1 9 0 9 13 11
16 13 3 10 9 16 1 9 13 10 9 10 9 13 10 11 16
6 13 1 15 15 10 9
9 15 3 1 9 9 13 1 9 13
19 13 3 16 0 15 15 3 13 15 10 13 1 10 9 10 9 10 13 15
14 10 3 9 3 13 1 9 7 10 13 15 13 1 15
41 11 15 13 1 10 9 10 9 13 1 15 9 16 13 0 15 10 13 1 9 16 1 10 9 10 9 10 11 13 1 11 11 16 10 9 10 9 13 1 10 9
4 9 1 9 13
8 3 9 13 9 15 13 7 13
10 10 3 11 13 10 9 7 10 9 15
3 0 3 13
20 9 13 1 10 9 10 1 12 7 12 9 13 9 3 13 1 10 13 10 9
9 16 3 1 9 10 9 3 1 9
4 15 3 10 9
17 10 9 1 13 16 15 13 10 9 15 13 13 1 9 1 9 9
6 10 3 9 12 3 13
5 10 3 9 12 13
2 3 13
14 16 3 13 9 10 13 13 3 1 9 13 3 10 9
18 7 13 10 9 10 15 1 9 16 10 9 1 9 11 11 13 10 13
15 1 10 3 13 10 9 1 9 13 13 1 10 13 9 13
8 13 3 10 9 3 1 9 13
11 15 3 9 9 13 1 10 9 1 11 11
7 15 3 1 11 13 11 13
5 3 13 9 7 0
5 3 13 0 7 0
8 0 3 15 12 13 1 11 11
12 16 3 15 11 3 10 11 9 13 1 9 9
2 13 3
13 3 3 15 16 13 0 1 10 9 10 9 13 13
28 16 3 13 10 9 10 9 13 10 9 10 9 15 13 1 9 13 1 9 16 10 1 9 13 16 10 9 13
3 9 10 9
6 3 3 13 9 7 9
7 16 3 9 3 9 1 9
12 7 3 3 3 13 9 13 10 9 3 13 9
23 3 3 13 9 3 3 13 1 9 3 13 3 1 10 0 7 0 9 15 3 3 13 13
8 9 13 7 9 7 9 7 9
8 13 3 15 16 3 15 3 15
3 15 15 13
32 13 3 16 1 9 10 9 13 15 10 0 7 10 9 15 1 10 9 15 3 13 7 13 7 3 9 9 13 15 3 11 11
5 3 3 10 9 15
12 13 3 15 16 16 0 10 9 15 13 13 15
6 3 0 15 13 13 15
11 13 15 3 3 7 13 15 13 16 15 13
15 0 3 13 1 0 3 7 3 0 1 10 13 15 1 15
4 10 9 3 13
16 13 3 16 11 12 9 13 12 1 10 9 7 12 1 10 0
17 7 10 3 1 10 9 1 9 13 10 3 1 10 0 1 10 9
3 15 13 13
16 0 3 13 12 9 12 3 1 9 11 1 9 13 15 13 11
8 10 3 11 9 13 1 10 11
5 13 3 10 3 11
6 13 3 1 10 9 15
2 13 3
5 13 9 10 3 13
6 13 7 13 10 3 13
12 3 0 10 9 10 0 3 3 10 13 10 9
8 15 3 9 1 11 9 9 13
14 7 3 3 10 1 9 13 13 10 1 9 3 3 3
5 7 15 13 10 9
7 13 10 9 7 10 9 15
5 10 9 15 11 13
8 13 3 7 3 3 9 9 13
1 13
11 15 11 13 15 16 16 13 11 15 15 13
13 13 3 3 15 9 13 16 9 13 0 10 9 13
7 13 1 11 15 1 9 13
3 10 9 13
15 1 3 11 11 7 9 15 13 7 9 7 9 1 9 13
6 15 15 13 9 3 13
7 10 9 3 1 10 13 15
6 0 9 0 10 9 13
10 15 13 1 15 1 9 16 15 0 13
10 10 3 13 15 13 10 9 15 3 13
10 15 3 9 16 9 3 13 15 3 13
6 6 3 13 10 13 15
6 15 3 1 9 13 9
16 10 3 15 9 1 12 9 13 1 10 13 10 3 15 3 15
11 16 3 15 13 7 13 13 3 1 15 13
2 13 3
8 9 13 7 9 9 3 3 13
7 10 3 9 13 1 10 9
11 0 3 15 13 16 3 15 3 13 0 13
8 16 3 9 13 3 13 1 9
42 0 3 13 10 9 10 9 15 13 9 9 9 9 9 9 9 9 9 9 9 9 9 9 9 7 10 0 0 15 13 15 3 13 16 10 10 0 13 9 9 3 13
6 1 10 0 3 13 9
14 10 3 10 11 11 10 9 13 1 10 9 7 10 9
6 16 13 9 9 3 13
7 3 13 0 15 13 15 13
11 15 10 9 13 7 3 13 10 9 10 11
10 16 3 13 15 13 15 15 13 13 15
19 10 3 9 15 13 0 7 3 1 15 0 10 9 13 7 3 1 10 0
6 0 3 10 0 9 13
2 3 13
3 9 3 13
8 15 3 3 13 9 0 3 13
12 10 3 13 1 10 9 1 10 9 13 9 0
6 10 3 0 13 3 13
6 9 3 0 13 3 13
17 3 3 16 9 13 13 10 0 1 15 3 3 1 10 0 10 9
8 13 0 15 9 13 10 15 9
17 3 3 10 13 0 9 13 7 13 15 13 16 1 10 15 9 13
10 7 3 9 15 13 7 9 7 0 9
6 10 0 9 15 15 13
11 15 3 10 9 10 11 1 10 9 15 13
12 10 9 10 9 15 11 11 1 10 9 15 9
1 6
16 11 9 11 11 1 9 9 10 0 10 13 7 0 1 11 11
12 9 15 7 9 1 9 9 15 7 9 11 11
32 1 15 1 15 3 13 13 1 9 10 10 15 13 1 10 9 10 9 15 1 10 13 15 1 9 9 15 10 13 1 10 11
26 1 15 3 13 13 10 9 10 9 10 0 15 13 9 10 9 15 1 9 10 9 1 9 10 9 15
143 1 0 3 15 13 10 1 15 9 1 10 9 11 7 10 9 10 1 15 10 0 3 13 13 1 15 9 13 1 10 9 15 16 10 9 10 9 15 11 11 10 9 10 9 13 15 9 9 7 9 1 9 15 13 10 9 10 9 15 1 10 13 15 15 13 10 9 10 9 15 15 10 9 10 9 10 9 15 1 10 0 7 15 10 13 9 10 9 15 1 15 10 13 1 10 9 10 9 10 9 15 15 13 1 10 11 13 15 1 0 7 13 15 1 0 15 1 10 0 1 15 9 7 9 7 9 7 9 7 15 9 13 3 0 1 10 9 0 7 7 1 10 13
28 7 15 13 1 10 9 15 7 15 13 9 1 15 10 9 15 13 10 9 15 10 9 10 10 15 1 15 13
37 7 15 13 0 10 9 7 10 9 15 1 15 3 13 1 10 9 10 9 0 1 10 9 10 9 10 9 10 9 10 3 13 1 10 9 10 9
30 1 15 3 15 15 13 3 1 10 9 10 9 15 13 10 9 10 9 7 10 9 7 13 9 9 9 3 3 10 0
57 10 3 9 0 13 1 9 1 10 0 9 15 15 13 15 7 13 15 0 10 9 13 10 11 9 13 13 7 13 7 13 1 10 0 1 11 11 16 13 1 10 9 10 13 10 13 9 10 9 15 1 9 1 15 1 11 11
7 10 3 9 13 13 1 9
7 3 1 9 16 3 15 13
19 15 3 13 9 13 1 11 11 1 9 0 15 13 10 9 16 1 15 13
45 3 13 16 3 15 10 9 1 9 10 13 9 1 10 13 9 1 9 0 16 13 10 9 0 1 11 13 10 9 10 11 7 0 10 9 10 9 9 3 13 7 0 1 10 9
17 3 3 1 11 11 15 10 3 13 3 13 3 1 10 9 10 11
59 15 3 13 10 9 15 10 13 10 0 12 7 10 9 10 9 13 10 9 1 10 9 15 10 9 10 9 1 9 13 16 10 12 13 1 15 1 12 0 9 13 9 7 13 10 0 1 12 9 10 9 1 10 9 13 10 9 1 15
25 7 13 13 9 15 10 3 7 9 10 3 16 1 15 13 10 9 10 0 1 12 9 1 10 9
51 3 3 3 13 0 7 0 7 13 9 10 0 7 0 10 9 13 1 10 9 10 9 7 9 13 0 15 11 11 1 15 15 9 13 13 1 9 0 1 9 1 15 3 15 13 1 9 10 9 1 9
105 0 1 15 11 10 9 10 11 1 15 10 9 16 3 13 10 9 10 9 10 9 10 13 15 1 15 16 1 9 13 15 10 9 3 13 1 0 1 15 13 13 13 10 9 15 1 10 9 10 11 15 0 9 3 13 10 9 10 9 3 3 13 10 0 9 15 7 9 1 9 13 10 9 0 7 0 7 0 10 9 1 11 11 1 10 9 15 13 9 1 10 9 10 9 10 9 10 13 15 1 10 9 10 9 15
14 3 13 3 13 1 10 9 15 1 15 15 13 9 15
86 0 1 13 10 9 15 1 10 9 1 15 15 9 1 9 7 1 9 13 16 13 15 1 10 9 10 9 15 9 13 1 10 9 15 1 10 3 9 13 10 11 1 10 9 1 10 9 15 1 9 13 7 13 16 13 13 1 15 10 0 15 10 9 7 9 7 9 7 9 13 7 10 13 10 9 9 10 11 16 13 1 15 10 9 10 9
36 10 3 13 1 15 13 3 15 13 3 13 1 10 9 10 13 1 15 15 10 9 1 10 9 7 1 11 11 1 15 10 9 10 9 10 9
1 6
36 13 3 15 15 10 9 1 9 3 13 10 9 15 13 1 15 9 7 9 1 9 13 15 1 9 13 13 10 9 10 9 1 10 9 10 9
14 12 9 7 12 9 3 3 13 1 12 9 10 9 15
6 12 9 12 9 12 9
14 12 9 7 9 15 10 1 15 7 1 15 7 1 15
5 13 1 9 13 9
4 13 9 10 9
15 10 3 13 15 13 3 3 16 3 13 1 10 0 10 9
15 10 13 0 13 3 10 13 1 15 10 9 16 13 10 15
124 7 15 13 15 3 9 15 3 9 15 3 9 15 3 9 7 9 1 10 9 10 0 1 9 9 1 9 10 9 10 11 16 13 10 15 1 10 9 10 9 7 10 9 10 9 10 9 1 9 0 1 9 9 10 9 10 11 16 3 13 0 13 7 13 15 9 10 9 1 10 9 10 9 1 9 1 10 9 10 9 13 3 1 9 13 1 15 10 15 15 13 10 9 11 1 15 15 10 9 13 7 13 1 15 9 10 9 1 9 1 9 12 0 9 10 9 10 9 13 1 9 15 1 9
54 0 3 13 7 13 1 9 3 15 13 3 3 10 9 13 1 9 10 9 15 13 10 9 13 13 10 9 10 9 1 10 9 10 13 1 15 1 10 9 10 9 15 15 13 15 13 10 9 1 9 9 15 1 9
59 15 3 3 3 13 10 11 16 3 15 13 7 1 15 13 3 13 9 1 10 11 13 15 1 10 0 9 10 0 9 10 13 1 10 9 10 9 13 3 10 9 10 9 15 7 13 10 0 9 10 1 9 13 1 9 7 9 10 9
4 13 7 3 13
5 7 13 9 10 9
4 10 13 3 13
15 3 3 13 13 10 0 9 10 0 16 13 13 10 9 13
22 15 9 0 1 10 9 15 3 13 7 3 15 0 1 9 10 9 16 13 9 10 13
15 7 3 13 10 9 10 0 10 9 1 15 13 1 9 9
16 15 9 7 9 7 9 7 9 7 9 13 1 15 1 15 9
31 13 3 9 10 9 3 9 0 7 13 1 9 3 3 10 11 13 15 7 13 15 1 15 9 7 9 10 9 1 9 9
26 9 3 7 9 15 7 9 7 13 1 15 3 13 0 7 9 7 9 7 9 15 3 13 7 3 9
5 15 15 13 0 9
13 1 0 3 13 10 9 10 9 1 10 9 10 9
5 3 3 13 0 15
4 13 3 3 9
5 3 3 9 1 9
9 7 3 13 10 9 10 0 10 9
4 3 3 3 13
10 10 3 3 13 1 15 0 13 3 13
6 15 3 10 13 9 13
2 3 13
13 13 10 13 7 13 1 10 0 7 13 15 10 11
19 13 3 3 3 13 3 3 0 7 3 0 13 10 9 16 10 9 0 13
48 7 3 13 9 1 15 13 9 7 13 1 9 13 15 9 7 9 7 9 0 13 7 13 10 9 15 10 9 13 3 1 15 1 9 10 9 15 11 11 10 9 7 9 13 15 1 9 11
25 10 9 10 0 9 3 10 9 16 9 13 9 10 9 3 3 10 11 9 10 9 15 9 10 9
15 7 3 10 9 13 10 11 3 3 10 9 10 9 1 15
49 10 9 13 10 9 3 3 10 11 13 10 9 7 15 13 1 15 16 15 13 13 10 9 10 9 1 9 16 13 15 15 0 10 9 3 13 9 7 9 7 15 10 0 7 16 13 0 7 0
7 10 13 10 15 9 15 13
24 15 3 3 10 15 9 13 7 13 7 13 15 3 3 10 11 10 9 16 9 13 10 9 15
20 1 0 13 9 10 9 7 10 9 7 13 10 9 7 13 10 12 1 9 12
9 15 3 13 1 11 7 1 10 9
14 3 3 15 10 1 12 0 10 15 9 3 13 3 15
7 10 3 9 16 13 10 9
8 10 9 13 10 9 15 1 9
4 0 3 13 0
16 7 10 9 3 13 10 9 15 7 13 15 1 9 7 9 9
58 10 9 13 10 1 9 9 1 9 7 9 1 9 9 15 3 10 11 3 1 9 3 0 7 3 9 11 13 10 9 10 9 1 9 1 9 13 3 10 9 7 3 9 13 16 0 16 15 13 0 0 13 1 9 7 9 7 0
12 10 0 13 1 9 7 1 10 9 10 9 15
15 13 10 9 10 9 1 10 13 15 13 1 10 9 10 9
31 3 3 13 15 10 9 1 9 7 9 7 1 10 9 1 10 9 1 10 9 10 9 0 1 10 0 10 9 1 10 0
19 1 0 13 10 9 10 9 16 13 13 1 10 9 10 0 7 0 13 13
42 13 3 13 10 9 15 1 9 7 13 10 9 10 9 7 13 10 9 1 9 10 9 10 9 1 15 13 10 9 10 9 1 15 13 15 10 9 10 0 10 13 13
71 7 10 9 10 0 13 7 10 9 10 9 15 13 9 9 1 15 9 7 9 13 1 15 9 1 9 7 1 15 13 1 15 9 7 9 1 15 10 0 7 1 15 16 15 13 9 1 9 10 9 15 1 9 13 10 9 10 9 1 15 13 1 9 16 1 15 13 3 13 15 13
14 9 10 9 7 9 1 9 1 9 9 7 9 11 11
20 11 7 11 9 11 11 15 10 0 1 11 11 10 13 1 11 1 9 7 9
12 9 15 7 9 1 9 9 15 7 9 11 11
50 13 10 9 15 1 15 10 9 15 3 1 15 9 15 1 15 15 1 9 10 9 13 1 10 9 15 1 10 9 1 0 9 1 10 3 13 15 0 16 10 13 1 15 9 0 13 1 9 11 11
37 3 13 0 15 0 13 1 15 15 1 10 13 15 1 10 9 15 1 7 10 9 15 7 1 10 9 7 9 10 9 9 15 10 9 15 15 13
13 9 3 15 10 9 16 13 15 15 1 9 11 11
43 7 0 13 16 10 9 15 3 3 7 3 13 1 9 7 15 9 1 10 13 15 10 13 16 13 0 7 0 1 9 11 13 9 9 10 1 11 11 1 9 7 9 9
50 13 3 15 13 9 16 10 1 15 3 1 9 10 9 13 16 10 9 15 0 1 11 13 1 0 10 9 7 10 0 15 7 10 0 10 9 1 9 13 10 9 15 3 13 3 10 9 10 9 13
11 15 3 1 9 13 16 1 9 10 9 13
15 15 3 1 9 10 11 13 3 3 13 9 13 10 9 15
2 15 3
14 3 16 15 9 7 9 7 9 11 13 7 1 0 13
3 7 3 13
48 13 3 16 0 15 13 1 9 1 10 15 9 7 9 10 9 11 11 1 10 9 7 9 15 16 1 15 13 7 1 15 9 3 3 3 3 13 11 1 10 9 15 7 1 9 7 1 9
9 15 3 10 13 11 7 10 13 9
10 16 3 10 13 1 9 0 15 9 9
15 13 3 1 10 12 10 9 13 1 10 13 7 1 11 13
4 0 3 3 0
8 10 3 13 10 9 0 1 15
35 7 0 13 13 16 13 7 13 15 15 1 10 15 9 7 9 10 9 16 10 9 15 13 1 11 11 1 15 1 10 15 9 3 1 15
51 0 3 10 9 10 11 13 16 7 13 7 13 15 7 13 13 10 1 15 16 13 1 12 9 12 9 13 10 9 10 9 7 3 13 1 15 1 10 13 15 13 15 9 9 15 3 9 7 0 1 9
31 3 15 13 10 1 11 3 0 10 1 15 13 7 3 10 1 15 13 10 0 9 13 15 13 1 15 7 3 13 1 15
58 16 15 3 9 1 11 16 15 9 9 16 15 9 9 16 15 9 7 9 13 15 10 9 16 10 15 13 10 0 9 13 0 10 12 13 15 1 9 7 1 9 7 10 9 15 13 13 15 3 10 15 0 13 7 3 10 0 0
31 0 13 1 15 15 3 1 11 11 15 1 9 9 13 3 9 13 10 13 0 9 7 15 13 9 9 13 1 9 9 13
29 3 0 15 3 3 13 3 3 1 10 9 15 0 7 3 0 3 1 10 9 15 1 9 7 9 10 15 9 13
16 9 3 13 10 13 1 15 7 10 13 7 10 13 1 10 9
44 15 13 1 9 7 9 16 13 0 7 0 9 9 0 0 9 0 7 13 1 15 13 3 9 1 9 9 9 13 1 9 15 1 9 11 16 3 1 0 13 7 1 0 13
17 7 16 3 13 1 10 9 7 9 10 9 15 13 7 13 15 15
9 10 3 15 3 15 13 7 13 15
17 13 3 1 9 11 11 3 13 15 16 3 15 13 13 10 1 15
10 15 3 13 0 15 3 10 1 15 13
15 10 3 9 15 13 16 3 9 9 1 15 13 1 10 9
9 13 3 1 9 16 3 0 3 13
33 0 3 13 11 10 9 7 0 7 9 15 15 3 9 7 9 10 9 15 13 1 15 16 13 13 15 15 7 13 16 13 16 13
5 3 3 13 0 9
5 7 10 9 13 15
13 3 15 3 0 7 3 15 16 3 9 1 9 13
13 3 3 13 15 16 13 15 3 13 7 15 0 13
7 10 0 9 15 13 1 9
11 10 15 13 15 15 3 3 0 15 3 0
4 13 10 0 9
3 13 10 9
9 16 15 13 0 13 1 9 15 3
10 15 13 15 9 0 13 1 10 11 9
76 7 3 7 13 15 9 13 1 10 13 10 9 11 11 10 9 15 1 15 10 15 13 7 13 9 16 11 13 7 13 1 15 3 13 15 9 10 1 9 7 10 1 9 11 10 1 9 9 1 10 9 10 13 15 7 10 9 10 9 15 7 9 9 15 13 10 9 15 16 13 1 10 9 10 1 0
11 13 3 16 13 1 15 3 13 1 11 11
6 9 15 15 3 13 13
2 12 3
5 15 3 0 0 13
11 7 16 15 3 13 3 0 10 9 15 13
7 3 1 15 13 10 15 13
13 9 15 13 9 7 13 10 3 13 3 13 9 15
39 15 3 10 9 1 9 13 1 3 3 9 13 9 11 11 15 13 10 9 10 9 15 0 10 9 10 9 15 1 10 9 10 13 15 7 13 15 10 15
15 3 9 15 0 7 0 9 7 9 15 3 13 1 9 0
10 11 13 7 11 13 10 15 13 1 9
4 6 13 3 15
4 13 1 9 3
2 3 13
1 13
3 10 9 3
19 15 13 7 1 15 10 9 7 10 9 1 9 10 9 15 13 1 10 9
20 7 10 9 10 9 10 13 15 9 13 10 9 15 7 10 9 15 1 11 11
25 10 0 9 15 13 0 15 0 15 0 15 0 15 0 15 0 16 15 9 7 16 15 9 0 13
13 15 7 13 7 13 7 13 7 13 1 15 0 13
19 13 3 1 9 3 16 3 3 13 10 1 15 13 1 15 3 13 13 3
5 3 16 1 9 13
3 13 3 13
3 13 3 13
14 1 15 7 1 15 13 7 13 7 13 7 13 7 13
6 15 13 1 10 13 15
7 3 3 13 13 15 10 9
27 13 3 3 15 9 16 1 9 10 9 16 13 1 11 15 15 9 13 1 9 9 7 9 3 3 15 0
14 3 16 13 10 9 7 13 10 9 10 13 1 9 15
14 13 13 1 11 10 1 15 9 9 9 0 0 10 9
17 10 3 9 15 13 15 9 15 1 10 9 15 1 9 1 11 11
13 10 3 9 7 9 15 10 9 1 10 9 10 9
1 6
6 13 15 0 1 11 11
6 13 15 10 1 15 9
5 13 15 15 10 0
20 11 9 11 11 1 9 9 7 11 10 9 10 1 11 0 7 0 9 1 11
8 9 15 7 9 1 9 9 15
78 13 10 9 7 9 10 9 15 11 11 3 1 15 13 13 10 9 15 1 11 11 7 10 9 15 13 1 15 10 0 1 10 9 10 13 15 1 10 9 15 13 1 10 9 10 9 10 9 10 13 1 15 3 3 1 15 10 9 13 13 7 13 3 3 1 15 1 15 9 13 7 13 10 9 10 9 1 9
25 3 13 1 11 10 0 9 15 15 13 0 1 15 9 10 11 10 3 13 15 10 15 9 1 9
79 1 0 7 15 1 15 9 13 3 13 1 15 13 7 13 16 13 10 9 10 9 15 1 15 9 7 9 0 13 3 10 9 1 15 9 1 15 9 0 13 7 13 10 9 10 9 1 15 9 13 1 10 9 10 9 15 1 15 9 7 9 1 9 13 10 9 10 13 15 1 10 9 10 9 10 0 1 10 9
27 15 13 15 1 10 9 10 9 7 13 1 10 9 10 9 10 9 15 1 15 13 10 9 10 9 10 9
36 15 13 9 10 9 10 0 0 15 9 16 1 15 13 10 15 1 10 9 7 1 10 9 10 0 7 10 0 7 9 7 9 7 9 7 9
19 10 15 1 15 7 1 15 13 7 15 13 1 15 7 10 15 1 15 13
13 15 13 9 0 1 10 0 16 13 1 15 15 13
35 3 1 15 13 15 10 9 13 7 1 15 13 10 15 1 15 13 1 10 9 10 9 15 1 15 7 10 1 10 9 7 10 1 10 9
67 7 15 3 13 13 7 0 10 9 1 10 9 10 0 3 3 13 1 10 9 10 9 15 1 10 9 13 15 0 7 0 7 0 1 15 16 3 13 10 9 13 7 0 7 3 13 1 10 9 10 9 15 13 10 13 1 15 9 10 1 10 9 15 13 15 11 9
57 3 13 1 10 9 1 15 7 13 10 9 10 9 10 11 1 10 9 15 1 10 9 15 15 13 10 9 15 13 15 9 1 10 9 10 9 10 13 15 1 15 13 10 9 10 9 10 9 10 13 1 10 9 7 1 10 9
51 3 3 13 10 0 15 15 13 10 9 13 15 10 9 10 9 10 9 0 1 10 9 15 13 11 1 15 10 9 10 9 15 15 13 13 15 9 7 13 15 9 1 15 9 16 13 15 9 0 1 11
15 1 15 3 13 13 1 10 9 15 10 13 1 15 1 9
56 13 3 15 13 0 9 13 1 15 7 10 1 11 7 15 3 13 10 9 15 1 9 16 13 10 9 15 13 1 9 7 1 15 9 10 9 10 9 1 9 10 9 10 9 11 1 15 13 15 10 9 10 9 7 9 0
8 0 13 16 15 15 13 1 9
89 13 3 15 15 13 10 13 1 10 9 7 0 9 1 10 9 10 9 1 10 9 10 9 7 3 1 11 16 1 15 13 15 10 9 10 9 3 7 13 1 15 13 15 13 10 9 15 9 7 9 1 15 7 13 9 0 1 10 9 10 9 10 9 1 10 9 10 11 13 15 1 10 9 1 15 3 13 1 10 9 10 9 10 9 10 13 15 1 0
42 7 15 0 13 10 9 7 10 9 10 9 15 13 15 1 15 13 15 15 10 9 13 10 1 15 9 10 9 15 13 0 15 7 15 13 1 10 0 13 15 10 9
13 13 10 9 7 10 9 13 1 9 13 15 1 15
23 3 3 15 15 13 1 9 7 1 9 7 1 9 9 7 9 7 9 15 13 9 10 13
5 10 3 9 10 11
44 15 15 13 13 1 9 7 9 10 9 15 13 13 3 13 1 10 9 10 9 15 7 3 13 10 9 1 15 15 10 9 1 10 9 7 9 13 7 13 13 10 9 10 9
15 16 13 1 11 1 10 9 10 9 15 3 13 1 9 13
14 15 13 15 1 9 10 9 1 10 9 7 9 10 9
17 16 3 13 10 11 10 3 13 3 10 11 13 1 0 10 9 13
8 10 3 13 3 10 1 10 9
13 13 3 7 10 9 15 13 1 10 11 1 10 9
15 3 10 11 13 10 9 15 3 3 15 1 15 13 1 9
26 13 3 10 9 10 1 10 9 9 9 9 9 0 7 10 9 15 13 9 1 15 13 10 9 10 9
10 1 15 3 15 13 3 16 13 1 0
45 3 13 1 15 13 10 0 9 1 10 9 15 7 13 10 0 10 13 1 9 1 9 10 13 15 3 3 13 9 7 0 9 7 9 0 9 9 0 7 10 15 7 1 15 11
26 13 3 3 0 10 9 0 7 13 9 9 9 9 9 9 13 15 7 13 15 16 15 1 15 13 9
11 1 15 3 0 10 9 15 13 9 10 9
17 7 10 9 10 11 13 1 10 9 15 1 15 3 13 1 12 9
3 7 0 13
8 10 9 10 11 13 1 15 3
11 1 15 9 13 7 13 15 9 9 9 0
22 7 15 15 15 3 13 1 9 7 1 9 15 1 9 9 11 13 10 9 9 1 15
9 10 9 13 10 9 3 13 1 9
10 10 9 13 10 9 7 3 13 1 15
6 0 3 0 13 1 9
10 10 9 3 13 10 9 15 16 3 13
21 10 9 13 1 15 10 1 9 9 3 1 9 3 0 7 1 9 9 13 10 9
21 15 3 13 1 9 13 3 10 9 7 3 9 13 16 1 9 13 10 9 10 9
10 10 3 13 13 15 13 7 3 13 9
18 10 9 10 0 7 10 9 10 9 13 13 16 3 15 13 9 1 9
37 10 9 13 13 1 15 1 9 13 3 3 1 15 16 10 9 13 15 9 10 9 13 10 9 10 11 1 15 3 13 16 13 15 3 13 15 13
9 1 9 13 1 10 3 10 9 13
45 10 1 15 15 13 15 11 10 0 9 7 0 9 7 9 1 9 15 13 1 15 1 15 0 16 13 10 1 15 7 13 10 9 15 1 11 10 0 7 0 9 15 13 1 15
5 15 15 13 10 3
30 13 15 11 10 0 15 7 11 10 9 11 1 15 13 9 16 13 1 15 13 15 7 11 10 13 11 10 13 1 9
26 13 15 11 10 1 15 9 11 11 3 13 1 15 1 10 9 16 13 0 7 13 1 15 9 10 9
17 13 3 15 16 13 0 9 1 15 7 10 1 11 7 10 1 11
9 13 15 11 10 9 10 0 7 11
13 13 10 1 11 9 7 11 7 10 1 9 15 9
23 7 3 13 1 15 10 9 13 16 3 1 10 9 9 13 7 10 1 11 16 3 15 13
10 13 10 9 15 13 1 9 16 15 13
6 10 9 10 15 9 11
4 10 9 1 15
15 11 7 11 7 11 10 9 9 1 9 9 7 9 11 11
4 9 15 7 9
80 13 10 9 3 1 15 15 9 13 1 10 9 15 3 13 15 10 9 10 9 7 10 9 10 9 7 10 9 10 9 10 9 15 11 11 1 10 9 7 9 15 13 9 13 1 10 9 10 9 15 16 10 9 15 3 13 1 15 1 9 0 7 3 1 9 7 1 9 0 7 9 0 3 13 15 13 1 15 1 15
32 7 15 9 15 13 7 10 9 13 10 9 1 9 0 1 9 9 0 16 13 15 9 15 10 13 1 10 11 7 1 10 11
36 1 15 3 13 10 9 10 9 3 0 1 10 11 7 1 10 11 7 1 15 9 10 9 15 10 1 10 9 13 16 3 9 13 15 13 15
37 0 3 13 9 10 9 15 10 1 15 16 3 0 13 7 13 7 13 3 13 1 11 13 1 10 9 15 13 1 15 10 9 10 9 1 0 9
33 7 3 3 1 9 9 13 3 13 7 1 9 9 9 9 7 13 1 9 9 7 1 15 7 1 0 13 1 9 13 3 11 9
13 7 13 0 1 0 15 3 16 9 13 10 15 9
21 3 13 15 13 13 15 3 0 10 9 10 9 7 3 10 15 9 16 0 15 13
9 13 3 9 10 9 15 7 10 9
17 9 7 9 13 1 10 3 13 15 15 13 1 15 10 9 10 9
47 15 9 7 10 9 3 3 7 3 7 3 15 10 13 13 3 13 3 12 0 15 3 9 9 15 13 15 7 13 7 13 1 10 13 15 3 10 9 10 13 15 1 10 15 9 7 9
34 7 1 0 3 15 13 10 9 3 16 13 9 9 1 15 10 9 13 3 9 9 7 3 13 3 9 9 15 3 13 1 15 10 13
21 15 3 9 13 1 15 1 9 9 9 3 9 3 13 10 9 15 13 1 0 9
17 3 13 13 1 15 15 3 11 7 3 7 3 7 13 15 10 11
22 15 3 15 9 7 9 7 9 9 3 3 3 15 1 10 9 15 11 1 10 15 9
9 15 3 13 10 9 15 7 10 9
40 3 3 13 13 13 1 11 0 7 13 11 10 9 15 7 9 10 9 1 10 9 10 11 1 10 13 15 7 13 1 10 9 15 10 15 13 1 10 9 0
7 0 3 13 16 1 0 13
16 7 3 16 1 15 13 13 15 16 13 13 3 3 13 7 13
25 1 0 7 15 3 13 13 1 10 13 10 9 15 16 13 15 10 13 7 1 0 13 10 9 15
39 15 3 9 13 10 9 13 1 15 1 15 10 9 15 13 1 15 1 10 9 15 9 7 9 3 13 1 10 13 15 10 9 7 13 10 9 10 9 15
18 0 3 10 9 7 9 15 7 10 9 15 11 13 10 9 15 1 15
46 15 3 10 9 13 7 13 10 9 1 15 7 1 15 3 3 15 1 15 1 10 13 15 10 9 0 1 9 1 10 9 7 9 15 1 10 9 10 9 15 11 1 15 10 0 15
1 6
29 0 3 9 13 15 7 13 1 9 11 16 3 13 1 15 10 3 13 15 13 7 13 9 3 7 13 16 13 3
10 13 3 15 9 13 15 1 10 9 11
61 0 3 13 9 10 9 10 9 15 13 15 1 10 9 13 0 15 10 15 9 13 1 9 7 9 3 1 9 9 3 3 10 9 10 3 13 10 9 10 3 13 7 13 1 10 9 10 9 15 16 0 9 1 15 0 3 3 13 15 7 13
11 3 3 13 15 10 9 1 9 7 1 9
9 0 3 15 0 13 1 10 13 15
12 7 3 13 15 1 15 10 9 1 0 10 11
31 13 3 15 9 13 3 7 13 13 7 13 10 0 7 13 10 9 15 3 15 13 16 13 3 1 10 3 7 15 9 13
20 3 13 3 15 13 9 1 10 13 16 3 13 3 3 10 0 10 3 13 9
20 16 3 13 16 11 13 7 13 3 3 10 9 10 13 1 10 11 13 1 15
23 0 3 15 13 1 9 9 16 15 10 13 10 13 1 10 9 10 9 3 3 13 10 13
23 3 0 10 9 1 9 1 9 9 7 1 9 9 13 1 9 7 10 0 1 11 13 0
6 7 3 3 1 9 13
13 1 3 10 9 7 10 9 9 3 9 13 15 13
13 0 3 3 13 16 9 9 3 9 1 9 3 13
21 3 13 9 7 9 3 0 15 13 9 3 10 9 10 1 9 13 7 3 3 13
14 15 3 9 3 13 1 9 16 10 9 15 3 9 13
9 15 3 15 9 9 13 7 9 9
5 3 13 9 7 9
10 10 3 13 9 13 7 10 13 9 13
14 15 3 9 13 13 13 9 9 7 9 7 9 9 9
11 3 13 15 7 13 12 10 12 3 3 13
27 13 3 15 9 13 10 13 1 15 7 13 15 1 9 7 13 15 7 13 15 3 1 9 1 10 9 15
3 13 1 0
3 13 3 15
4 9 13 10 0
3 13 10 0
3 13 1 15
18 13 3 15 0 1 0 15 13 7 3 10 0 13 1 15 7 1 15
2 3 13
3 1 15 13
9 0 3 9 9 1 11 11 1 15
4 10 9 3 13
3 15 3 13
3 10 0 13
5 1 15 9 0 13
30 0 3 10 9 10 9 13 15 0 7 0 15 10 9 7 10 9 7 10 9 3 1 10 9 10 9 15 11 11 13
4 9 13 1 15
7 13 10 9 15 1 9 0
10 13 15 10 9 13 10 9 15 10 9
16 11 7 11 7 11 10 9 9 1 9 9 15 7 9 11 11
12 9 15 7 9 1 9 9 15 7 9 11 11
53 13 13 10 9 3 1 15 9 3 0 13 16 13 10 9 15 7 13 10 9 12 0 15 15 1 15 16 0 15 1 15 13 1 10 9 10 9 1 10 9 15 7 9 1 15 10 9 15 7 10 9 15 13
105 9 10 0 9 10 9 1 10 13 15 10 9 10 9 1 15 7 13 16 0 1 9 13 10 13 15 9 7 15 10 13 9 1 15 1 10 9 10 9 11 1 9 1 9 9 15 1 9 9 13 9 10 3 13 9 7 10 3 13 10 9 10 9 15 11 15 9 13 9 0 1 9 10 9 7 1 10 9 10 9 15 3 13 13 1 10 0 15 7 13 1 15 10 13 16 13 10 9 15 1 15 1 10 9 0
49 1 15 7 13 3 1 15 16 15 13 10 9 10 9 15 7 13 15 9 9 7 9 9 1 9 16 13 10 9 10 9 15 11 1 15 7 15 1 15 1 10 9 10 9 15 7 9 11 11
7 3 15 15 13 1 15 9
40 3 16 3 13 10 9 0 7 13 10 9 10 9 10 9 10 9 10 13 7 13 1 15 13 9 7 9 16 15 1 10 9 10 9 13 13 15 16 13 9
13 7 3 10 13 13 1 10 13 15 1 10 15 9
7 10 3 9 3 13 10 9
8 0 10 13 3 16 1 0 13
57 7 3 13 10 0 15 10 9 11 13 10 9 10 9 15 7 13 10 9 10 9 15 15 13 10 9 1 9 10 11 1 15 9 7 9 7 9 9 7 1 15 9 9 10 13 16 15 10 9 10 9 3 13 1 10 13 15
27 7 1 0 13 15 10 9 9 9 1 10 13 15 10 9 16 13 0 10 3 13 10 9 7 13 10 9
45 15 3 13 13 10 9 3 1 15 9 13 1 9 16 13 15 10 9 1 9 1 9 1 9 9 7 9 9 1 15 7 13 15 1 10 9 15 1 9 9 10 9 15 11 11
37 0 3 10 9 15 11 11 7 10 9 10 9 15 10 13 15 7 13 9 0 7 9 0 1 9 13 15 10 9 7 13 1 15 9 7 9 0
5 3 3 15 10 9
13 0 3 13 10 9 15 13 15 7 13 1 10 0
12 13 3 1 9 1 15 16 15 13 13 7 13
18 10 3 9 13 15 10 9 1 10 9 10 9 7 1 10 9 10 11
27 13 3 15 9 1 9 10 9 15 11 11 13 15 1 15 9 3 13 7 3 1 10 9 15 13 1 15
33 0 3 13 3 13 13 15 16 3 13 1 15 7 3 9 13 1 15 7 1 9 7 9 9 7 9 13 1 10 3 13 15 15
15 3 16 3 13 9 7 16 15 9 13 15 1 10 13 15
18 10 3 0 13 7 13 1 9 11 11 16 1 9 13 10 15 9 13
6 15 3 9 3 13 13
13 16 3 15 3 13 10 9 15 1 10 9 0 13
5 3 13 15 16 13
9 7 3 3 0 13 7 13 3 9
14 0 3 10 9 10 9 13 15 10 9 3 1 15 9
5 10 9 1 15 15
12 10 9 10 15 9 11 15 13 9 1 15 9
10 10 9 10 9 15 11 11 1 15 15
20 11 9 11 11 1 9 9 9 15 7 11 11 10 9 15 11 0 9 1 9
12 9 9 9 1 9 9 7 11 11 10 9 15
30 3 13 15 13 1 11 13 1 11 16 13 15 3 13 7 13 9 7 9 0 15 9 13 3 3 9 9 10 1 9
34 10 3 9 10 9 13 9 1 0 9 7 9 0 7 9 0 15 15 13 13 1 9 13 13 9 3 13 7 15 13 7 1 15 13
56 13 3 16 0 10 9 16 15 15 3 13 13 0 16 0 9 3 13 0 3 7 0 0 7 0 0 7 0 9 7 9 9 9 9 9 9 0 7 16 15 0 10 13 9 13 1 10 9 10 9 10 0 9 15 13 15
25 9 13 10 13 15 11 11 10 9 15 16 0 15 13 13 1 9 10 0 13 0 7 9 7 9
7 7 13 16 13 13 1 9
24 7 1 0 13 16 1 15 0 13 11 11 10 0 9 1 9 10 13 13 1 15 1 9 0
17 10 3 9 10 9 0 0 0 9 9 7 9 1 10 9 10 9
1 6
32 0 10 9 13 15 9 11 1 10 13 1 15 9 16 13 1 15 10 0 9 13 9 7 0 9 15 15 13 1 10 9 13
13 15 13 11 7 11 15 13 10 11 16 13 3 13
12 13 3 0 15 13 9 9 9 9 1 15 9
19 1 9 7 15 10 1 9 13 16 0 7 0 9 13 1 15 9 7 9
22 12 3 9 12 7 9 9 7 9 9 11 11 10 13 15 9 1 15 10 9 9 0
15 13 3 13 10 9 1 15 9 13 0 9 1 9 7 9
31 3 3 9 1 9 0 1 9 7 9 13 15 3 1 9 7 9 7 9 7 9 0 7 15 13 9 13 9 1 9 0
7 9 1 9 13 1 15 9
12 13 3 9 3 13 7 13 9 7 13 1 9
4 11 3 0 13
2 3 11
7 10 3 9 13 1 9 13
15 13 3 1 10 9 16 13 1 9 7 9 7 9 1 9
7 16 15 9 13 0 9 13
34 13 3 10 9 0 13 12 9 9 0 0 0 0 0 3 0 3 9 7 0 0 0 10 0 9 3 13 9 13 1 9 1 15 9
13 16 3 15 10 0 9 13 3 13 3 9 9 13
10 3 0 16 3 13 1 9 13 10 9
18 13 3 7 9 0 13 1 10 3 16 3 1 9 13 7 9 10 9
5 3 0 3 13 0
4 3 13 0 13
9 9 3 0 3 0 0 0 1 15
17 10 3 3 13 9 15 0 13 7 0 9 1 9 10 1 11 11
8 0 15 13 13 13 1 15 3
21 16 3 13 16 13 3 13 1 9 9 13 15 13 9 9 13 9 7 9 10 9
8 7 3 0 13 10 10 9 9
44 10 3 9 3 13 16 1 0 9 13 15 10 9 13 9 0 7 9 9 1 9 0 13 10 0 9 13 13 13 9 15 10 9 13 1 9 1 9 10 0 7 13 10 9
11 3 15 9 9 0 7 15 0 1 9 13
7 13 3 1 9 9 7 9
20 0 13 10 9 0 13 9 11 11 13 10 9 10 9 7 10 0 9 15 13
5 13 3 15 1 9
8 10 3 0 9 1 0 13 0
15 10 3 9 1 15 0 13 9 13 9 10 3 7 10 13
18 1 0 3 13 7 13 16 13 1 9 13 15 13 9 15 9 3 0
4 13 0 7 13
20 15 15 10 9 13 7 9 13 10 0 1 9 1 9 1 9 1 9 1 9
9 16 13 13 10 9 10 9 10 9
17 3 13 10 1 15 9 15 13 15 1 9 1 9 10 9 10 9
10 1 0 13 16 15 10 9 0 13 15
5 13 15 7 10 9
10 0 3 13 7 15 13 7 10 13 15
19 0 3 13 7 13 3 9 0 3 9 0 3 9 0 3 9 1 15 9
5 9 13 10 3 9
19 16 3 15 9 9 7 0 13 13 0 10 0 9 13 7 9 13 10 9
7 0 3 13 0 1 10 9
19 10 3 3 9 7 13 13 1 9 7 13 10 9 7 10 9 9 7 9
6 7 0 13 16 0 13
30 9 13 3 0 9 12 13 12 9 9 1 9 0 13 16 13 16 13 16 0 9 13 16 13 13 16 15 9 0 13
4 0 3 9 13
14 3 3 13 10 11 13 13 13 9 16 10 0 9 13
21 3 3 3 0 13 13 10 9 3 0 3 0 7 3 0 7 0 13 10 3 13
13 13 3 0 13 13 13 15 9 13 10 13 9 1
7 3 3 15 13 1 10 11
17 16 15 0 13 9 13 15 7 3 13 10 9 16 10 3 9 13
13 1 0 9 3 13 3 3 3 1 12 7 12 9
11 10 13 1 15 13 16 3 10 0 9 13
20 13 1 10 9 7 11 11 7 10 0 9 16 0 13 1 9 15 13 1 9
8 9 3 15 13 7 13 9 0
3 15 0 13
14 3 13 7 9 0 13 1 10 9 7 10 0 15 9
9 15 9 10 9 0 13 13 1 9
4 15 3 3 13
22 15 13 1 9 9 10 0 9 15 9 0 13 16 3 10 9 10 9 7 10 9 13
10 10 3 0 13 9 3 13 16 9 13
12 7 3 13 16 0 13 7 0 10 10 9 13
4 0 13 7 13
50 16 15 13 7 3 13 13 9 10 10 9 15 11 11 7 10 1 9 9 13 15 13 7 13 1 9 7 9 1 15 13 9 9 9 9 0 9 13 9 10 9 7 13 10 9 13 9 13 10 9
8 13 3 9 0 10 9 1 9
11 15 3 13 1 10 9 16 3 13 15 13
7 13 3 9 7 9 0 13
7 15 3 6 9 9 0 13
8 13 3 9 9 9 9 9 9
6 13 10 0 9 10 9
15 13 10 0 9 1 15 13 7 13 10 0 9 1 0 9
63 13 1 9 10 13 10 15 7 11 11 10 13 1 11 11 10 0 9 13 15 10 9 0 0 1 10 9 10 9 15 11 11 15 9 0 13 10 0 7 0 9 10 9 10 13 7 9 10 13 10 0 13 9 9 13 0 15 13 15 9 7 13 13
5 15 9 7 9 0
1 6
21 6 11 10 9 13 13 10 0 9 7 9 10 0 9 15 15 13 1 10 9 13
17 11 9 11 11 1 9 9 1 9 9 10 1 11 11 11 0 9
12 9 9 9 1 9 9 7 11 11 10 9 15
61 9 13 10 9 15 13 1 9 1 0 9 16 0 13 10 1 15 9 1 10 9 15 9 7 9 13 15 13 13 15 10 9 16 9 13 9 13 10 1 15 0 9 15 13 0 1 10 9 15 11 7 10 9 15 11 13 3 16 3 1 15
20 1 15 9 13 15 13 10 9 10 9 15 13 1 15 1 10 9 10 9 15
14 3 3 13 15 10 9 9 9 7 9 7 9 7 9
79 3 3 13 10 9 10 9 15 7 15 10 9 15 7 13 10 9 1 9 9 10 13 15 7 13 9 0 3 1 10 9 15 7 1 0 9 7 9 10 13 15 1 11 11 1 9 0 13 3 3 1 10 9 10 9 15 11 11 13 3 10 9 13 3 9 7 9 1 10 9 1 15 13 15 9 7 9 7 9
17 13 3 15 13 7 13 16 0 13 10 9 15 13 1 0 10 9
16 9 13 13 9 15 1 15 13 1 9 7 9 10 1 11 11
15 13 0 16 13 15 15 10 1 10 11 15 13 11 7 11
26 13 9 10 9 10 11 9 16 3 15 13 7 10 9 15 3 13 7 13 1 11 3 13 15 7 13
12 13 15 10 9 13 9 1 9 1 0 10 9
8 7 15 1 11 13 0 15 13
30 15 3 9 15 13 1 10 9 10 1 11 11 7 15 13 1 15 1 0 9 0 13 0 9 15 0 13 3 0 13
11 15 13 13 10 10 9 9 16 10 13 13
11 16 3 7 13 15 3 13 16 3 3 13
8 10 13 9 13 0 10 9 13
8 13 3 15 10 9 9 1 15
13 13 11 11 13 1 0 1 9 11 1 10 9 15
14 1 15 13 1 9 3 0 7 10 9 10 9 3 13
19 1 0 15 13 1 10 0 16 3 15 9 13 10 1 11 11 1 9 0
5 16 3 13 3 13
4 16 13 3 13
6 16 13 3 0 13 15
5 16 13 0 0 13
15 0 13 13 1 10 9 3 13 1 15 0 1 9 10 13
13 13 15 0 13 10 9 9 0 13 10 9 10 9
5 10 3 0 9 13
19 15 13 11 7 11 15 1 10 9 13 13 9 3 13 7 13 10 15 9
26 10 3 0 9 10 9 13 13 10 9 0 13 9 10 13 15 7 13 1 9 15 10 13 10 9 9
16 1 0 3 9 3 13 0 9 0 7 0 7 3 0 7 0
5 7 15 3 1 9
4 15 3 1 9
5 10 3 0 9 13
14 13 3 9 9 9 9 1 10 13 10 9 1 0 9
41 9 3 9 3 13 13 7 0 13 1 15 0 0 1 9 13 10 13 16 13 15 10 9 9 1 9 9 7 13 1 10 10 9 9 13 1 15 1 10 0 9
10 0 3 13 16 1 0 9 13 9 0
34 13 3 10 9 0 0 9 0 0 9 0 0 0 0 0 0 0 0 0 9 0 13 0 3 3 0 13 9 9 10 3 9 15 13
3 7 0 13
26 1 0 3 13 10 13 1 10 9 7 13 9 13 9 13 9 0 3 13 7 3 1 9 9 13 13
22 15 9 3 11 7 11 13 11 3 3 0 13 10 9 9 13 10 9 0 1 10 9
12 10 3 9 15 0 13 15 3 3 10 0 13
10 15 9 13 7 1 15 15 13 10 9
11 7 15 3 10 13 13 3 1 11 11 13
12 0 3 9 7 9 13 1 10 0 13 7 13
31 15 3 13 1 15 13 7 13 13 1 15 13 7 16 1 9 0 9 13 10 13 15 13 1 9 1 9 10 1 11 11
28 15 9 0 7 0 1 9 1 9 1 9 1 9 10 1 9 16 0 13 10 10 9 9 1 15 9 0 13
21 13 1 10 9 7 11 11 10 13 13 13 7 0 7 10 9 15 7 10 9 15
3 13 10 9
1 13
6 13 1 15 9 7 9
33 13 3 9 3 10 13 9 3 13 7 1 10 0 9 15 13 9 13 10 9 7 1 3 10 9 10 9 13 1 3 10 9 13
5 15 3 13 1 15
1 13
3 9 13 9
4 10 9 15 13
11 15 3 3 13 7 10 9 10 9 15 13
3 10 9 13
3 10 9 13
31 0 13 15 10 10 9 9 15 13 15 10 9 1 0 10 9 10 0 9 3 0 3 15 7 3 15 10 13 10 9 15
5 13 13 1 15 3
12 11 3 15 13 13 10 3 9 7 13 1 11
3 11 1 11
3 11 1 11
5 11 13 0 1 15
5 11 3 13 1 11
16 10 9 15 13 1 11 1 11 13 13 7 10 9 3 10 9
7 11 10 9 0 15 0 13
8 13 15 10 9 1 10 9 15
4 15 3 15 13
6 3 3 13 10 15 9
12 1 10 0 15 9 15 15 13 7 15 15 13
24 10 3 9 15 13 7 13 15 16 1 15 10 9 13 7 13 15 10 9 7 13 1 9 9
1 6
8 13 11 7 11 7 10 11 9
4 11 13 1 11
6 11 3 13 1 11 13
4 13 1 9 13
13 13 15 11 7 11 7 11 7 11 7 10 9 15
4 10 9 1 15
53 11 9 9 9 3 11 11 1 9 0 9 7 9 9 10 1 9 1 9 9 0 15 13 10 0 9 1 9 0 13 3 9 0 10 9 15 1 9 15 13 15 1 9 10 9 15 9 11 0 9 1 0 9
35 0 1 13 15 1 9 16 10 13 13 7 13 1 9 0 3 15 15 13 16 15 13 0 12 9 9 9 13 0 3 1 9 9 7 0
47 13 3 10 9 0 13 3 9 9 3 0 3 0 3 0 3 9 3 0 7 0 0 0 0 0 0 13 10 1 10 9 0 9 16 0 13 7 13 1 10 9 10 13 7 10 13 13
26 13 3 0 0 0 7 9 3 10 1 10 9 15 13 13 15 0 9 13 13 15 3 13 0 9 1
7 13 15 1 15 0 15 9
7 9 3 9 0 9 9 0
21 1 15 9 13 15 3 16 13 1 10 9 3 13 0 9 7 9 9 13 10 9
4 15 0 10 0
16 10 3 13 7 0 15 0 7 13 15 7 10 9 7 10 9
14 10 3 9 13 0 13 7 0 7 1 15 9 0 0
8 15 3 13 15 13 10 13 9
12 9 0 13 0 0 13 10 9 10 9 10 9
34 9 3 1 9 0 3 0 3 9 0 13 0 16 13 10 0 0 13 0 0 0 0 0 13 10 0 9 16 3 10 9 10 9 13
19 1 10 9 9 9 9 0 0 16 10 1 0 13 15 13 13 1 15 0
28 9 0 9 13 1 15 0 13 3 13 3 13 7 15 9 13 0 16 10 9 10 10 9 15 9 13 1 15
64 13 3 10 9 10 9 0 15 9 13 15 16 13 10 9 7 10 0 9 3 7 3 7 3 13 1 10 3 9 13 10 0 9 7 9 10 9 10 0 9 7 9 15 11 11 15 13 15 1 15 16 13 15 1 15 9 7 13 15 9 0 9 0 9
9 0 13 7 13 7 13 1 15 9
23 13 15 9 9 13 13 1 15 9 0 0 13 15 13 0 13 0 15 13 9 1 15 9
21 13 3 3 3 15 0 0 13 13 9 7 9 0 1 9 7 9 13 0 13 15
57 16 3 10 9 7 10 9 13 10 9 15 9 3 1 9 10 1 9 15 13 15 7 1 10 15 9 13 15 1 9 9 7 9 9 0 15 13 1 15 3 1 11 11 10 9 15 16 13 10 0 9 9 13 1 9 9 0
7 0 13 0 7 0 10 9
11 0 3 9 7 9 7 9 7 9 0 13
5 13 3 0 7 0
17 0 9 1 12 7 0 9 13 13 16 13 10 0 7 13 13 0
13 3 13 11 1 15 7 11 13 13 1 15 1 11
11 9 10 0 7 9 3 13 16 15 15 13
16 13 3 3 10 15 0 9 13 1 10 0 9 16 3 13 0
6 13 10 13 15 1 9
5 10 9 1 15 15
29 9 9 11 11 7 9 10 9 9 10 0 7 0 15 7 9 10 9 7 9 10 9 15 7 10 1 9 15 9
12 9 15 7 9 1 9 9 15 7 9 11 11
47 13 10 9 15 3 9 15 13 1 10 9 15 13 15 10 9 7 10 9 15 13 1 10 9 11 7 1 15 10 0 16 10 9 10 9 15 0 13 1 9 15 0 10 1 15 1 11
19 9 3 0 13 7 9 1 10 9 15 16 10 9 10 0 13 1 15 9
32 13 15 1 10 15 9 15 13 1 10 9 9 10 3 15 0 3 3 7 15 7 15 0 15 13 15 15 0 13 10 15 9
20 1 3 10 15 9 15 13 13 16 3 3 1 9 10 0 15 13 7 1 0
32 3 3 1 0 13 1 9 16 0 15 13 3 3 3 9 7 1 9 9 0 3 15 15 3 3 15 7 1 9 7 1 9
9 16 3 15 13 9 13 15 3 15
10 16 3 15 13 15 7 13 0 15 13
6 15 9 13 10 15 9
2 15 13
9 16 3 13 15 16 3 15 15 13
13 13 10 9 15 13 15 13 16 3 1 15 13 13
6 3 3 7 13 15 9
9 13 3 16 1 10 9 15 13 15
16 13 15 11 10 0 15 1 11 11 9 9 9 9 10 0 15
10 10 9 10 9 11 11 1 10 9 15
31 3 7 3 3 10 9 13 10 9 1 10 9 1 0 10 9 0 13 15 1 9 15 13 9 15 1 15 7 13 10 9
41 15 13 9 10 9 7 9 10 9 15 13 7 10 15 10 9 10 9 15 9 10 9 13 13 1 0 10 9 1 0 0 0 13 10 9 15 0 1 15 13 9
6 15 3 13 3 10 9
4 15 3 13 15
2 7 3
11 15 13 15 1 9 7 15 13 15 1 9
10 3 3 3 13 10 0 1 10 9 13
6 7 13 15 15 9 9
6 7 1 3 10 9 13
12 10 13 10 9 15 9 7 10 9 15 9 9
4 1 3 10 9
15 1 0 13 15 10 9 10 9 15 9 9 1 10 0 15
16 7 15 1 9 9 10 9 13 7 9 10 9 15 13 10 9
5 15 13 15 3 13
12 7 15 3 9 13 7 3 9 13 15 7 13
11 15 3 10 0 13 7 10 9 15 3 13
7 1 15 3 10 9 13 3
14 13 1 0 15 16 3 13 10 0 15 9 10 9 15
10 1 0 13 3 13 15 10 13 16 13
31 15 9 13 13 1 10 9 1 10 13 1 15 13 13 10 9 9 7 7 9 7 0 9 7 9 0 9 1 10 15 9
11 3 3 9 13 10 9 10 13 1 15 13
5 13 3 3 15 13
12 15 13 9 16 13 15 7 9 9 16 13 15
6 13 15 0 15 1 9
5 9 7 9 13 15
11 1 10 3 13 15 10 15 15 13 15 0
8 3 3 3 13 15 10 15 13
25 13 3 15 1 15 10 15 7 1 15 10 15 0 9 1 9 13 10 9 10 9 15 1 9 13
10 10 7 3 13 7 10 13 1 12 15
9 1 15 9 3 13 9 15 13 13
7 13 10 9 15 10 9 15
5 1 0 9 13 15
12 3 3 6 15 7 10 9 15 15 13 10 9
42 16 3 10 9 13 9 7 9 3 0 3 13 10 15 16 1 10 9 13 10 10 9 13 10 9 0 13 10 9 7 13 0 15 9 9 1 15 10 13 0 13 9
9 3 3 3 9 13 7 9 11 13
10 1 15 3 13 0 13 13 10 13 13
28 3 9 0 9 0 0 13 10 9 7 9 10 9 15 11 0 13 10 13 15 3 3 11 1 0 10 9 15
17 0 3 0 9 1 11 13 16 15 0 9 13 10 9 10 13 0
6 15 3 9 13 1 15
15 7 11 3 0 1 0 10 9 15 3 9 1 9 10 13
24 11 3 3 9 1 10 9 15 15 9 13 15 16 10 9 7 10 9 10 9 1 9 0 13
7 3 3 13 10 9 10 0
37 3 16 10 9 15 13 3 13 10 9 15 3 1 10 9 1 10 9 10 9 1 10 0 3 13 10 9 15 1 9 7 13 10 9 15 12 9
4 3 13 10 9
7 15 3 3 13 10 9 15
12 3 13 1 10 9 15 16 13 1 10 9 15
20 7 13 15 1 0 9 16 15 10 3 13 16 3 13 15 1 15 11 10 9
14 0 3 10 11 13 16 10 9 10 9 1 9 0 13
3 1 10 13
15 3 16 10 9 15 13 3 13 10 9 15 3 1 10 9
4 15 3 13 13
5 15 3 13 12 9
10 3 10 13 15 10 9 13 1 10 9
8 7 13 16 3 13 13 1 9
15 13 3 16 13 9 13 1 10 9 15 13 15 1 15 13
7 3 3 13 13 3 3 0
14 7 3 13 10 9 10 9 0 3 13 10 9 10 13
9 13 3 1 10 9 10 13 3 13
19 3 13 1 10 9 15 16 13 1 10 9 15 3 10 9 1 9 9 13
14 7 13 10 9 1 10 9 10 0 1 15 10 9 15
6 16 13 1 10 9 15
23 16 3 13 15 13 1 15 7 10 0 13 3 13 1 9 3 15 13 9 3 1 11 13
16 1 0 9 3 13 3 16 10 9 15 13 3 13 10 9 15
13 16 3 15 11 13 3 3 1 0 13 1 0 9
7 3 13 9 10 9 10 9
20 10 3 13 1 10 9 15 7 0 13 1 10 9 15 3 1 10 0 10 9
17 13 3 13 1 0 10 9 16 3 1 10 0 15 9 13 10 9
8 15 3 0 7 13 10 9 15
5 1 15 15 10 9
15 13 3 9 0 13 10 9 11 10 9 10 9 13 10 9
18 3 3 13 9 3 13 13 10 9 15 13 3 1 15 1 9 1 9
17 13 3 1 9 10 9 10 9 16 13 9 7 9 13 1 0 9
32 15 3 9 1 9 13 1 9 13 10 1 10 9 16 13 9 7 7 9 1 9 13 13 10 13 7 13 16 3 15 13 9
15 7 1 15 13 3 1 10 9 3 3 1 15 13 1 9
15 7 3 15 15 13 10 9 7 13 1 10 9 3 3 11
4 15 3 13 15
5 3 3 1 0 13
9 15 9 1 10 9 1 10 9 11
19 7 13 13 15 10 13 15 0 9 0 13 1 10 9 9 1 10 9 11
14 1 15 0 15 10 9 7 0 13 16 0 13 10 9
31 7 3 13 13 9 1 10 9 3 9 13 10 13 15 15 10 9 10 9 10 9 10 9 7 13 9 13 9 3 0 9
8 15 3 10 13 9 0 9 0
3 0 3 13
7 7 0 13 16 13 10 9
39 0 3 10 3 13 13 7 10 9 10 0 7 0 13 9 0 7 0 13 9 9 9 7 13 9 7 13 3 13 1 9 13 15 10 9 10 9 7 13
24 9 3 10 13 10 1 15 13 3 9 7 13 9 0 0 1 15 3 13 13 9 1 10 9
14 13 3 1 15 0 10 0 7 13 9 16 3 3 13
23 3 3 0 10 9 13 10 9 15 7 10 9 15 13 1 10 9 15 13 10 0 7 13
29 13 3 0 15 10 0 13 9 1 10 9 10 9 1 9 16 3 0 13 9 3 10 1 9 7 9 13 10 9
16 10 3 11 13 10 9 16 1 15 13 0 13 13 1 15 13
6 7 3 13 13 10 9
38 1 15 0 13 10 9 13 10 9 10 9 10 0 10 9 15 13 9 16 1 12 9 0 1 15 0 13 10 9 0 9 13 10 13 13 10 13 9
65 0 3 10 11 9 11 9 10 9 10 0 10 13 11 13 1 10 9 10 9 7 13 15 15 3 0 1 15 13 11 0 3 13 9 9 3 3 3 9 11 15 13 9 9 0 0 0 7 9 9 7 9 9 13 13 3 10 9 10 9 13 9 1 10 0
29 7 10 3 1 10 9 11 10 9 13 9 13 13 10 9 1 10 9 0 13 10 9 15 3 13 1 10 9 11
14 15 3 3 13 1 15 13 11 7 10 13 10 9 13
10 1 3 15 9 10 0 1 10 0 13
12 7 3 9 13 1 11 3 11 10 12 13 13
32 16 3 3 9 1 10 0 9 13 10 9 3 1 15 13 15 3 9 1 10 9 11 0 13 9 7 3 1 10 9 11 13
10 13 3 10 9 1 9 3 9 9 13
3 13 3 16
9 15 9 1 10 9 1 10 9 11
26 9 3 3 13 13 9 1 10 15 0 7 0 15 3 13 10 9 9 3 0 9 1 15 13 10 9
12 7 10 3 0 13 13 9 1 10 9 13 13
13 15 3 1 10 13 15 1 10 9 0 13 10 9
6 0 3 13 3 15 13
22 10 9 3 9 13 9 13 9 10 9 3 10 9 10 1 10 9 9 1 10 9 13
5 9 3 1 10 13
11 15 3 9 1 10 13 9 7 7 9 13
8 3 0 13 15 3 0 15 13
17 16 3 3 13 1 9 3 3 13 9 13 10 13 1 9 10 9
14 15 9 7 9 13 10 0 3 13 11 13 13 10 9
16 3 3 0 13 9 15 3 0 13 9 9 15 1 0 9 13
12 16 3 10 0 0 13 0 3 3 0 13 9
4 13 3 15 13
3 6 9 13
46 7 13 1 10 9 11 7 1 10 9 11 9 0 3 1 10 9 15 13 10 9 15 1 9 13 15 10 9 15 13 15 1 9 11 16 15 3 13 1 10 9 15 7 15 13 15
2 13 9
2 13 9
3 13 10 9
9 3 15 13 15 1 0 1 0 15
14 3 0 13 10 0 15 7 10 9 15 3 3 13 3
7 1 10 13 0 13 10 0
7 10 3 13 7 13 1 9
21 9 3 13 10 0 1 15 10 7 9 7 10 9 7 10 9 10 9 15 13 0
39 1 3 10 0 9 9 10 13 0 0 0 13 9 7 10 9 10 9 13 3 9 1 15 9 0 13 10 9 7 10 9 11 10 13 7 10 9 10 9
8 1 15 3 13 3 13 1 9
91 0 3 3 13 1 3 10 0 9 3 13 10 9 10 9 13 1 3 10 0 3 10 9 0 10 9 3 1 9 15 13 1 15 7 10 10 9 9 0 13 10 9 10 0 3 13 10 10 0 9 3 10 0 9 13 9 15 9 1 10 9 10 13 1 15 9 7 7 9 13 3 13 1 9 13 10 13 0 1 9 7 9 7 0 9 9 9 1 9 9 13
40 11 3 13 9 10 13 0 1 10 0 7 0 9 3 0 0 13 3 0 10 9 7 1 9 9 7 9 1 3 10 0 9 13 3 1 10 0 0 9 13
46 16 3 10 9 9 7 9 7 9 9 13 10 13 13 1 10 10 9 9 15 3 10 9 10 11 15 1 9 0 15 13 0 10 9 13 10 9 15 1 0 9 1 10 13 9 13
26 7 1 0 9 0 9 13 16 9 13 1 9 10 1 10 0 9 9 10 9 13 10 13 10 0 9
8 3 3 9 9 9 13 10 13
7 3 3 10 0 1 9 13
11 0 10 9 10 9 15 13 1 15 10 9
14 7 10 9 3 7 15 10 9 10 9 10 9 3 13
19 9 3 10 3 9 10 1 10 9 0 13 0 3 10 0 0 9 1 0
23 3 3 1 0 13 0 11 0 10 0 7 1 0 10 9 3 13 10 9 10 9 1 15
25 7 16 3 13 15 3 10 9 13 1 10 0 1 9 1 9 0 16 13 15 3 13 1 9 9
15 3 3 3 1 9 10 9 1 9 9 1 10 9 15 13
33 7 1 15 13 10 9 3 13 1 3 0 9 3 3 10 11 3 13 1 10 0 13 9 1 0 1 9 13 10 15 13 1 9
7 7 1 15 9 9 1 9
8 0 3 9 9 7 9 13 9
6 3 13 1 10 9 13
5 9 7 9 3 13
4 9 3 13 15
6 9 7 1 9 3 13
2 3 13
15 6 13 1 9 9 13 1 15 10 13 10 9 10 9 15
7 13 10 0 16 10 0 13
13 1 15 9 13 13 1 10 9 10 9 11 11 3
19 7 15 3 9 13 1 9 13 7 10 0 3 13 9 15 3 13 13 9
27 0 3 12 1 9 13 9 1 10 0 13 1 0 10 9 10 0 13 16 13 10 0 15 9 10 9 15
9 12 3 9 13 1 10 0 10 13
8 13 3 15 3 10 9 10 0
4 1 3 10 13
11 0 10 9 15 13 1 15 1 10 9 0
37 13 10 9 10 9 0 0 3 10 13 7 13 15 1 9 9 7 0 9 3 13 10 9 15 3 9 15 7 13 3 0 3 15 13 13 10 9
28 3 3 13 15 1 10 13 10 9 10 9 3 1 9 13 9 0 3 15 9 9 7 9 9 13 13 10 0
12 13 15 9 11 1 9 1 12 7 12 9 13
27 15 13 0 13 9 10 10 9 10 9 13 7 10 9 10 9 0 13 1 15 13 7 10 9 10 9 13
4 13 3 10 13
2 15 9
2 15 13
5 13 9 10 9 15
21 3 3 10 9 13 7 10 9 10 13 15 1 9 13 13 13 15 0 9 7 13
10 3 13 3 10 9 15 15 13 0 9
13 9 3 13 9 16 10 9 10 9 13 13 10 9
11 3 3 0 15 15 10 13 13 7 3 13
17 10 3 0 15 1 9 13 7 16 13 3 13 10 9 15 1 15
12 15 3 3 13 9 1 9 7 9 1 9 9
6 1 0 3 13 10 0
15 9 13 13 10 9 9 9 1 10 3 1 13 10 13 13
15 9 11 13 10 3 13 9 7 3 13 16 13 15 10 9
8 1 3 10 9 13 13 10 9
5 1 3 9 0 13
14 13 3 13 10 13 9 16 13 7 10 13 15 9 13
27 9 13 11 1 10 3 13 13 13 9 1 9 10 9 15 1 15 13 10 9 7 10 1 9 9 13 9
21 9 13 1 9 10 9 3 0 1 9 13 1 11 7 11 10 0 10 9 10 0
13 13 3 10 10 9 13 9 15 9 7 9 10 9
18 9 3 0 11 9 1 9 9 13 3 1 9 9 16 0 13 10 13
25 1 9 13 0 15 3 13 10 9 7 3 15 13 7 13 7 13 16 0 7 0 13 1 10 9
8 10 3 0 13 13 16 9 13
12 7 16 3 0 13 1 15 13 13 3 9 13
7 3 3 0 13 0 13 0
4 13 3 15 9
32 9 13 11 10 11 13 7 10 0 13 10 10 9 13 1 15 13 16 1 11 13 15 9 13 16 3 1 0 13 0 10 9
6 3 15 3 1 9 13
10 9 1 13 13 11 10 11 7 10 11
16 9 11 13 1 10 9 10 9 11 13 7 1 10 9 15 13
21 9 11 13 13 0 1 10 9 15 16 13 0 10 9 7 3 13 10 9 10 9
31 9 11 0 13 13 13 9 9 11 3 13 13 10 9 10 9 3 0 13 9 9 0 9 13 10 11 9 10 9 10 11
9 9 13 11 3 13 10 9 10 9
6 10 3 0 3 13 13
17 9 13 10 9 7 10 9 10 9 16 3 10 13 10 0 13 15
9 9 10 9 11 13 13 1 12 9
13 9 11 10 9 3 13 10 13 13 10 9 1 9
18 13 15 3 13 10 9 1 11 11 11 11 11 7 7 11 7 10 9
5 15 1 9 13 9
2 13 9
3 13 9 9
3 13 9 9
3 13 9 9
3 13 1 9
3 9 13 0
11 15 3 13 3 13 10 9 16 0 9 13
1 13
1 13
1 13
4 1 9 9 13
23 7 0 15 13 1 10 9 3 13 10 9 10 9 1 15 0 15 13 16 3 1 15 13
50 3 7 15 0 13 13 15 9 9 9 13 15 7 10 0 9 1 9 13 10 13 15 9 13 1 10 10 9 9 7 9 11 15 1 10 13 15 9 13 9 9 13 1 0 7 10 9 10 9 13
18 13 3 10 0 13 1 10 0 1 15 9 16 3 13 10 9 15 13
5 15 3 13 9 13
6 13 3 15 9 15 13
3 1 9 13
6 3 9 15 13 10 9
7 15 3 9 15 3 13 9
15 16 3 1 13 9 15 0 13 15 3 9 7 3 9 13
11 3 10 3 10 9 15 9 13 9 7 13
10 3 0 3 13 10 9 10 9 7 13
13 15 3 9 1 3 10 13 3 13 9 13 7 9
10 0 3 9 0 10 1 15 13 13 9
24 3 10 13 9 7 10 13 9 13 7 9 0 13 10 9 15 16 3 10 0 13 13 3 3
50 9 13 1 15 7 10 9 15 1 15 13 10 9 13 16 15 13 1 10 9 10 9 16 15 9 9 3 13 13 7 1 0 13 10 0 16 15 9 7 0 3 11 15 1 9 12 13 10 9 15
10 13 3 16 3 3 13 13 10 9 13
10 9 3 9 3 13 3 1 9 13 15
27 3 3 13 13 7 13 9 7 9 7 9 7 9 7 9 9 7 9 9 15 10 13 13 3 13 15 9
4 0 13 7 0
18 16 3 0 3 13 1 9 13 10 13 0 3 15 10 0 1 9 13
7 15 10 9 10 9 13 3
4 3 3 13 13
12 3 3 15 13 3 0 10 9 7 3 10 9
16 10 3 3 3 13 10 10 13 9 3 13 16 13 10 3 13
15 11 9 7 9 11 11 9 10 12 9 10 1 10 9 13
18 15 9 13 9 15 3 9 13 0 13 16 10 9 15 10 9 13 9
19 16 3 15 15 13 9 13 1 10 13 9 15 3 7 3 13 7 13 15
9 10 3 13 13 9 9 13 7 13
12 3 3 13 10 9 0 16 13 15 1 10 9
8 9 0 0 1 15 10 9 15
23 13 3 10 9 1 10 9 7 13 10 9 7 10 9 15 13 7 10 9 10 9 15 13
9 3 3 10 0 1 10 9 15 13
18 0 9 15 13 9 16 0 13 13 10 9 10 9 15 13 10 13 15
3 1 9 13
6 10 3 9 0 13 0
10 0 3 13 1 10 0 9 13 7 13
6 3 10 9 13 13 9
6 10 3 9 13 13 9
5 3 13 9 15 0
23 15 9 0 7 15 9 0 3 13 13 1 10 9 10 9 1 15 3 13 9 7 9 9
15 13 3 15 9 0 1 10 13 0 1 10 13 0 1 9
7 9 3 9 9 9 3 13
19 3 13 15 9 7 9 9 1 9 13 10 0 9 10 13 13 10 9 15
20 3 16 15 9 9 13 7 3 9 0 13 9 13 10 9 10 9 15 1 9
10 13 3 15 7 13 7 3 13 15 13
25 10 3 13 1 9 0 10 10 9 7 13 3 9 9 13 7 9 9 0 0 1 10 9 15 13
17 16 15 13 0 13 3 13 9 15 7 13 9 15 0 0 10 9
15 9 15 3 1 9 13 10 9 10 9 15 11 11 10 9
55 16 3 13 1 9 15 9 0 1 9 0 13 3 3 0 1 0 9 7 13 1 10 13 10 9 10 0 7 13 15 13 3 3 7 10 9 13 15 13 3 7 13 1 10 9 15 3 13 1 15 7 13 9 9 0
4 13 9 15 0
20 3 10 9 13 10 0 10 9 0 1 9 7 9 10 9 15 13 10 13 15
11 3 10 0 13 15 7 0 13 15 1 9
10 3 15 13 10 0 9 10 13 1 15
16 16 3 9 13 0 1 10 9 13 10 0 15 3 15 3 13
13 15 3 0 10 9 13 13 3 1 12 13 15 0
7 10 3 13 3 13 13 3
2 3 13
9 16 3 3 13 13 3 13 9 9
11 3 13 7 3 13 3 1 9 9 13 13
3 13 9 9
14 15 10 9 9 15 16 9 13 15 13 9 3 3 13
34 16 9 7 9 0 13 7 13 10 0 9 13 3 15 15 1 15 13 1 9 13 7 13 3 13 3 15 10 0 10 9 15 10 9
12 3 3 10 9 16 3 13 9 0 13 1 15
3 7 13 15
7 15 9 13 7 15 9 13
18 13 15 10 9 15 1 10 9 7 15 15 13 1 10 9 15 10 9
7 15 13 16 12 13 10 9
6 3 10 9 13 7 13
16 11 10 9 15 3 1 9 13 13 11 10 9 15 1 10 9
21 13 16 10 9 13 10 9 15 7 1 10 9 10 9 13 7 13 10 9 10 13
10 13 3 11 10 9 7 13 15 1 9
4 7 9 9 13
11 13 16 1 9 13 9 7 3 1 9 0
17 3 3 3 11 10 9 3 1 9 13 13 10 9 7 0 9 13
16 3 3 10 9 1 9 0 13 3 3 10 9 1 9 0 13
15 16 15 1 9 3 13 0 0 9 0 13 3 0 10 9
21 6 3 10 9 0 13 7 1 9 0 13 13 1 0 9 3 10 9 10 13 13
10 3 3 10 9 0 9 13 7 0 13
6 6 0 9 0 9 13
23 10 9 13 1 10 9 15 10 13 0 10 9 7 13 10 9 10 9 7 13 1 10 11
18 15 3 9 9 7 7 9 9 7 7 0 13 7 13 10 9 10 0
7 10 3 9 15 13 9 13
2 0 0
18 1 15 13 10 9 7 9 7 1 15 13 10 9 10 1 9 9 13
8 1 10 0 9 13 9 7 9
7 3 13 9 15 0 3 13
13 3 10 9 1 10 0 9 13 10 0 7 10 0
10 3 13 9 15 9 9 13 7 9 9
5 3 0 0 13 9
6 15 0 7 0 1 15
11 13 1 10 0 9 10 9 15 1 9 9
11 3 3 9 7 9 3 9 7 15 0 9
19 10 3 3 9 0 3 0 13 3 0 0 0 0 9 7 9 0 0 0
9 9 3 9 1 9 13 10 13 9
7 3 9 7 3 9 1 15
12 3 3 1 10 9 15 10 13 1 10 9 15
4 13 7 3 13
7 13 7 13 7 3 13 13
8 7 3 13 1 10 3 13 15
12 9 3 13 16 10 9 10 9 9 13 10 9
12 15 16 3 13 9 13 10 9 0 10 9 13
7 7 13 16 3 10 9 13
9 1 9 13 10 9 15 13 1 15
4 0 3 13 9
2 3 13
4 0 3 13 9
4 13 3 10 9
6 13 10 9 7 13 15
7 13 9 0 7 13 9 0
3 13 7 13
1 13
11 10 9 15 1 9 13 7 10 9 1 9
4 3 13 15 9
13 10 13 9 7 13 10 9 15 13 9 7 13 9
10 16 3 9 13 3 13 9 9 7 9
8 15 3 15 13 10 13 10 0
4 13 3 10 13
16 3 7 3 13 1 0 10 9 7 13 3 9 7 13 7 13
6 15 3 13 10 10 3
10 9 3 13 10 1 0 13 3 7 13
22 1 10 13 15 16 10 9 13 7 13 7 13 0 7 0 3 3 13 1 10 9 15
5 15 9 0 0 13
10 13 3 0 13 7 3 13 9 15 13
8 13 13 1 10 9 15 10 13
10 10 9 15 13 7 10 9 15 0 13
22 10 9 15 7 10 9 13 7 10 9 15 1 9 15 13 7 13 10 9 15 3 9
26 6 10 9 10 9 10 13 10 9 15 10 13 1 15 13 7 10 9 10 13 1 10 9 9 8 13
6 13 1 10 9 7 13
7 13 10 9 15 1 9 9
1 13
3 13 10 0
8 13 3 9 1 10 9 10 9
17 6 10 9 13 10 0 9 10 9 13 1 15 16 13 0 7 0
10 13 10 9 15 16 10 9 10 9 13
8 3 13 1 15 9 16 3 13
7 6 10 9 1 10 9 13
16 9 13 9 10 9 7 10 9 10 9 15 13 1 10 9 9
4 6 13 10 13
16 10 9 11 13 7 10 9 9 13 16 0 13 10 9 7 0
15 13 3 15 10 6 6 7 10 3 3 16 3 1 9 13
1 13
2 13 15
1 13
4 13 15 1 15
16 13 10 0 10 9 7 13 1 15 13 9 1 10 9 10 9
13 7 10 9 10 9 13 10 13 7 13 15 10 9
7 3 16 9 13 13 13 15
22 11 9 13 0 15 7 9 13 10 3 13 7 3 13 1 10 9 9 12 7 9 12
15 7 3 13 7 10 9 13 9 7 10 9 13 10 9 15
32 9 15 16 15 1 15 13 1 10 9 7 13 15 15 13 16 10 13 0 1 9 9 15 13 9 15 1 9 7 13 9 9
27 11 9 11 11 0 0 9 11 11 11 11 7 11 1 9 9 9 1 9 9 1 9 7 9 9 11 11
5 9 15 7 9 13
53 0 10 9 7 9 10 9 15 11 11 10 1 10 0 15 9 13 15 1 9 13 1 9 11 11 1 0 1 9 0 7 0 7 0 13 1 9 1 15 10 1 9 9 13 1 9 1 9 0 13 1 9 0
36 1 15 13 0 3 16 9 13 1 0 9 16 10 9 15 10 9 0 9 10 13 1 9 3 13 13 1 9 7 9 7 9 1 9 11 11
4 15 3 13 13
36 1 15 9 13 7 13 9 10 1 10 1 15 9 13 13 1 15 7 15 9 13 10 1 15 9 11 13 10 1 11 9 7 10 1 0 9
28 15 13 16 3 15 15 3 13 15 15 3 13 15 1 10 13 15 1 9 0 13 1 9 1 15 13 9 13
19 3 13 10 9 10 9 15 13 3 13 1 10 13 15 9 1 9 11 11
27 3 9 9 3 13 10 0 1 10 9 15 9 7 1 10 13 15 0 3 0 0 1 15 9 13 16 13
5 0 13 16 15 0
30 10 9 15 13 1 10 9 10 9 1 9 0 1 9 15 13 3 13 3 1 9 0 7 0 1 9 13 9 7 13
12 3 15 9 3 9 7 15 9 15 3 9 9
7 13 10 9 7 10 9 13
34 13 3 15 9 7 15 9 7 9 7 9 7 15 9 3 0 9 10 0 0 9 13 16 1 15 13 1 9 16 13 16 0 10 9
33 1 15 13 9 13 1 9 3 13 1 3 9 0 0 3 0 3 9 13 13 9 0 1 9 0 13 0 9 0 9 1 11 11
4 3 13 1 9
16 6 13 1 11 9 0 0 0 7 10 13 1 15 3 3 13
6 15 3 10 9 10 13
27 13 3 9 15 13 10 13 0 13 1 9 9 7 9 9 7 9 9 15 13 10 9 13 1 15 3 13
25 15 3 9 0 0 9 9 0 9 1 9 16 10 9 13 10 1 9 15 13 1 10 0 15 9
4 3 3 9 9
3 3 3 13
41 0 13 3 0 7 0 13 10 0 9 15 13 1 10 9 10 9 15 1 10 9 13 0 16 16 15 13 15 3 0 1 10 0 9 13 13 10 9 1 9 9
23 13 15 0 9 1 10 9 7 9 3 13 7 9 3 1 15 13 1 9 0 9 3 0
14 3 3 13 10 9 10 9 13 13 10 10 0 9 9
2 15 13
3 10 9 13
3 10 9 13
18 10 9 13 1 15 9 10 9 3 0 10 0 7 0 7 3 10 0
8 15 3 9 16 13 7 13 13
10 7 16 13 7 13 13 0 9 1 9
18 1 0 3 13 16 3 11 13 1 15 15 13 9 16 13 10 9 15
11 15 9 3 13 7 13 9 1 10 9 15
4 15 13 3 13
5 13 3 10 13 3
6 10 13 3 13 10 9
5 7 15 3 13 13
13 15 3 13 1 9 13 3 10 1 10 9 13 9
41 9 11 11 15 13 15 10 9 13 10 9 15 15 13 13 1 9 7 13 13 1 10 9 15 10 9 15 11 15 13 10 9 10 9 7 10 9 11 11 15 13
16 0 10 13 7 10 13 10 9 10 9 7 13 10 1 15 13
4 10 3 9 3
42 9 15 7 9 1 10 13 7 10 13 7 10 13 7 1 10 12 9 15 1 10 9 15 7 1 11 11 10 9 10 0 10 0 10 0 7 10 9 10 9 10 9
35 10 13 15 7 13 15 1 10 9 15 1 10 9 15 7 13 15 9 9 10 9 7 9 15 15 10 9 7 10 9 1 10 9 10 9
1 6
23 6 13 1 10 9 7 13 15 15 9 7 15 15 13 7 13 1 15 15 10 9 10 9
21 15 13 10 9 7 10 9 13 9 10 9 10 13 7 10 13 7 10 13 10 9
33 15 11 10 9 15 7 0 1 10 9 7 9 7 9 1 11 13 1 10 9 10 13 11 1 10 9 10 9 7 1 10 9 11
9 7 13 13 10 9 15 13 1 15
68 10 3 9 15 7 10 9 0 3 9 0 3 9 7 10 9 15 3 9 9 7 10 9 15 0 9 3 1 9 13 7 10 9 15 3 9 9 0 7 13 1 10 0 9 15 9 12 7 1 10 9 15 9 0 0 13 7 10 9 15 3 10 9 13 1 10 9 15
11 7 16 13 15 13 1 10 9 15 3 0
2 3 13
31 15 13 10 0 7 10 0 7 10 13 7 13 0 7 6 13 13 1 10 9 10 9 7 13 10 9 10 9 7 10 11
13 13 3 15 13 7 15 13 7 15 13 13 1 0
20 0 13 10 13 10 12 9 1 10 0 15 10 13 1 0 10 12 9 10 0
30 13 10 9 15 7 10 9 7 10 9 15 7 16 3 13 13 0 7 13 10 13 15 9 7 3 13 7 13 15 0
11 7 13 1 15 16 10 9 15 10 0 13
11 13 3 3 13 7 13 7 10 0 9 13
17 16 3 3 13 15 7 13 10 9 15 1 10 9 15 16 3 13
13 7 0 13 16 13 10 9 10 9 15 3 15 13
10 10 13 9 13 15 10 9 13 10 9
17 10 13 13 15 13 1 10 9 10 9 15 13 1 10 9 10 9
12 0 13 10 0 7 10 0 15 13 0 7 13
5 15 13 15 13 13
16 6 13 13 10 9 1 15 1 9 16 13 7 13 9 9 12
11 13 0 1 9 7 13 15 10 9 10 9
10 10 13 9 13 15 10 9 13 10 9
10 10 13 3 3 13 1 10 9 10 0
8 7 10 9 10 1 11 9 13
10 0 13 10 13 10 9 10 0 10 0
10 3 13 3 15 13 10 9 10 9 3
1 13
16 16 3 3 13 15 0 7 13 1 15 1 10 9 10 9 15
10 10 13 9 13 15 10 9 13 10 9
27 10 13 13 15 10 9 10 13 7 13 15 9 0 7 1 10 9 9 0 13 15 15 13 3 3 10 13
8 7 10 9 10 1 11 9 13
20 0 13 10 9 10 9 10 13 10 9 15 3 9 9 7 10 9 15 0 9
25 13 15 10 9 7 10 9 7 10 9 7 10 9 7 10 9 7 10 9 15 10 0 0 10 0
14 7 13 15 9 16 13 7 3 13 13 1 10 9 15
20 6 13 15 1 9 7 10 13 1 15 1 9 0 16 3 13 1 10 9 15
7 7 10 9 15 13 1 9
21 7 13 15 10 9 16 15 13 10 13 9 7 9 7 13 15 15 1 10 9 15
8 3 15 13 13 16 15 3 13
44 7 10 13 7 10 13 1 9 10 9 15 13 15 9 1 10 9 7 13 15 1 9 0 3 10 9 10 0 13 3 3 15 13 1 10 9 15 7 13 15 10 9 10 0
10 10 13 9 13 15 10 9 13 10 9
8 7 10 9 10 1 11 9 13
9 13 13 7 13 10 0 15 13 13
11 3 3 13 15 10 9 13 1 10 9 15
10 13 3 3 13 7 13 7 13 7 13
16 16 3 3 13 13 3 9 7 3 3 13 15 9 13 1 15
21 7 0 13 9 1 11 15 3 13 10 9 15 7 13 1 15 1 0 16 0 13
33 10 13 3 13 1 9 0 7 3 3 13 10 9 15 1 10 9 10 9 7 13 10 9 15 1 10 9 15 7 1 10 9 15
10 10 13 9 13 15 10 9 13 10 9
21 0 13 10 0 10 0 10 13 10 9 11 10 13 7 15 13 7 13 7 15 13
11 6 13 1 15 9 13 15 15 13 13 15
15 3 0 13 9 7 13 15 10 9 7 3 13 10 9 15
17 6 13 1 10 9 10 11 10 13 15 0 13 7 3 13 7 13
17 6 13 15 16 13 7 13 1 10 9 15 7 13 16 15 13 15
29 16 13 10 9 10 9 15 3 15 15 13 1 10 9 10 9 10 13 13 1 10 9 0 13 10 13 1 10 9
2 13 0
52 10 13 13 15 9 1 10 9 10 9 15 7 3 3 3 13 3 7 13 1 15 10 9 10 9 15 7 10 9 10 9 10 9 15 10 0 11 10 13 1 10 9 1 10 9 15 7 10 9 15 10 0
10 10 13 9 13 15 10 9 13 10 9
16 0 13 10 6 10 9 10 0 7 0 10 9 10 9 10 9
10 13 15 10 9 16 7 0 13 7 0
5 6 0 13 7 0
16 3 16 0 13 7 7 0 7 0 13 15 13 1 10 9 15
59 16 13 16 0 13 7 13 7 15 9 13 7 3 13 16 15 13 10 0 7 0 7 0 7 0 7 0 13 15 13 1 15 9 13 1 9 16 13 7 9 0 16 13 7 3 13 10 9 10 9 15 7 9 13 10 9 15 16 13
4 13 3 7 13
7 6 13 1 10 9 7 13
22 16 15 13 10 9 15 7 13 10 9 7 13 1 15 7 13 1 15 7 15 1 15
10 10 13 9 13 15 10 9 13 10 9
23 1 0 13 7 6 9 13 1 10 9 7 10 9 10 0 15 13 3 9 13 1 15 13
10 13 3 7 13 15 15 13 13 1 0
4 3 13 1 9
24 7 3 10 9 9 12 7 1 10 9 12 0 13 13 1 9 0 7 1 10 9 15 9 0
10 7 1 10 9 13 9 7 9 7 9
24 7 12 9 9 13 1 10 9 15 13 10 12 9 10 9 7 1 10 9 3 9 0 0 9
16 7 1 0 10 9 7 3 10 9 12 9 13 9 3 7 3
17 7 10 12 9 12 1 12 15 13 1 9 12 3 7 3 13 9
8 7 9 3 13 9 7 9 13
16 0 0 0 9 10 9 10 9 10 13 7 10 13 7 10 13
20 7 15 13 1 10 9 7 1 10 9 7 1 10 9 13 10 9 7 13 15
13 7 13 0 16 15 0 13 13 10 9 7 13 15
7 7 12 1 10 0 13 15
2 3 13
20 6 13 10 9 10 1 10 9 11 10 9 11 13 10 9 7 10 12 9 15
12 7 13 7 13 1 10 0 10 13 1 10 9
30 7 16 13 10 9 10 12 9 7 10 12 0 13 1 10 9 13 15 9 7 9 0 13 9 15 13 10 9 10 0
6 7 10 12 9 13 6
6 7 10 0 13 7 13
1 13
23 7 13 7 6 9 0 7 10 13 1 15 13 9 7 13 15 9 7 13 13 7 16 13
1 13
27 7 13 15 9 0 7 10 13 1 15 13 15 13 10 9 1 10 9 7 16 15 13 7 13 15 9 0
1 13
8 7 10 9 7 10 9 3 13
1 13
20 7 13 7 6 9 0 7 10 13 1 15 9 15 9 7 10 11 13 1 15
24 7 13 15 9 1 10 0 10 9 13 1 9 7 1 9 7 1 9 7 1 10 9 10 9
25 7 16 13 10 0 9 13 1 10 9 10 9 10 13 1 10 9 10 9 7 1 10 9 15 13
5 7 13 9 0 13
30 7 13 15 15 9 0 7 13 15 16 13 3 9 0 16 13 7 10 9 15 7 10 9 15 10 13 13 3 3 0
7 7 13 10 9 7 10 9
34 7 1 0 13 12 9 13 1 10 12 9 10 9 13 10 12 9 10 9 16 3 13 9 1 10 9 7 1 10 9 7 1 15 9
6 7 13 10 9 10 13
8 12 9 13 1 15 9 9 11
62 1 9 11 12 9 13 1 9 11 12 9 1 9 11 12 9 1 9 11 12 9 1 9 11 12 9 1 9 11 12 9 1 9 11 12 9 1 9 11 12 9 1 9 11 12 9 1 9 11 12 9 1 9 11 12 9 1 9 11 12 9 13
38 1 0 13 7 6 9 0 15 13 15 15 13 1 15 9 7 9 7 9 7 9 13 1 10 9 7 1 10 9 13 9 0 7 9 1 10 9 15
5 7 13 9 0 13
1 6
1 6
3 7 13 15
4 9 15 15 13
3 7 13 15
27 1 0 13 1 10 9 10 9 7 13 15 9 7 9 1 10 9 15 7 10 13 1 10 9 13 1 15
33 3 13 3 7 13 3 7 3 13 1 15 10 9 7 15 9 16 10 9 10 1 0 10 9 13 15 7 13 15 1 9 9 9
10 7 13 10 9 15 9 1 10 9 15
14 7 3 13 10 9 10 0 13 9 1 10 9 3 9
17 7 13 10 9 10 9 10 9 10 0 1 9 10 9 1 10 9
19 7 13 10 9 10 9 7 13 15 1 10 9 10 9 7 13 1 10 9
9 7 13 9 7 9 7 9 7 9
13 7 10 12 9 10 13 10 12 9 13 15 16 13
4 7 10 0 13
13 7 13 9 7 9 13 1 9 7 13 1 10 9
17 7 10 0 10 9 13 7 10 0 10 9 13 7 15 9 0 13
10 7 3 9 0 9 13 13 1 10 9
5 7 10 0 9 13
23 7 13 1 10 9 9 0 13 3 9 7 13 1 10 0 10 9 7 1 10 9 10 9
8 7 10 9 10 9 13 10 9
18 7 13 10 0 10 9 1 9 7 0 10 9 13 1 10 9 16 13
5 7 10 0 9 13
33 7 13 10 0 10 9 7 10 0 10 9 7 10 0 10 9 16 13 10 0 15 7 10 9 3 13 10 0 15 7 10 9 3
19 7 13 9 1 10 9 13 1 10 9 7 13 15 10 9 10 9 10 9
28 7 13 10 9 10 9 7 13 9 1 10 9 3 9 9 0 7 13 10 9 7 10 9 1 10 9 10 9
30 7 13 15 16 3 13 10 9 10 9 7 15 0 7 15 9 3 3 10 9 15 3 13 10 9 10 9 1 10 9
12 7 13 15 16 3 13 15 7 16 13 9 12
10 7 10 9 15 3 9 9 3 13 9
24 7 1 10 9 0 13 10 9 10 9 7 3 3 13 15 7 13 13 7 13 10 9 1 15
59 7 10 9 10 9 0 9 13 1 9 7 1 10 9 15 3 9 0 9 7 10 9 15 3 9 9 7 13 9 3 9 9 7 10 9 15 3 9 13 7 13 9 3 9 0 7 10 9 10 9 15 3 9 9 9 0 13 1 9
8 13 1 15 9 10 9 10 9
12 15 9 15 3 11 7 1 10 0 9 13 11
5 10 9 10 12 13
5 7 10 0 9 13
22 7 13 10 12 9 10 13 1 10 9 7 9 7 9 7 9 16 13 10 0 10 9
9 7 10 9 10 9 10 0 9 9
4 13 10 9 15
19 7 10 9 10 9 3 9 9 7 1 10 9 15 13 9 7 9 7 9
25 1 10 12 9 0 13 10 0 10 9 1 10 9 7 10 9 7 10 9 10 13 1 10 9 15
15 10 3 9 10 9 1 10 9 15 13 7 1 10 9 15
12 10 3 9 15 0 9 13 9 7 1 15 13
40 7 13 15 9 0 13 1 10 9 13 9 7 10 9 1 10 9 15 7 10 9 15 3 10 9 7 10 9 15 3 9 9 7 13 1 10 9 15 9 13
23 7 13 10 9 15 10 0 1 10 9 10 3 0 1 10 9 7 13 9 0 3 9 13
10 7 16 13 13 10 12 9 10 15 9
7 7 13 9 1 10 9 13
83 7 10 9 15 13 13 1 10 9 7 1 10 9 13 10 9 15 10 0 1 10 9 7 13 1 10 13 1 10 9 10 9 15 13 10 9 7 10 1 15 7 10 9 7 10 1 15 7 10 9 7 10 1 15 16 9 3 13 7 1 10 9 10 9 10 0 9 3 13 13 7 13 10 9 10 9 16 13 10 15 9 10 9
1 13
7 7 13 1 10 9 13 15
4 13 15 10 9
3 7 13 15
7 7 13 15 9 0 9 13
25 7 10 9 10 1 10 9 13 3 7 3 15 13 16 13 10 9 7 10 9 10 0 13 9 12
12 7 13 10 12 9 15 7 13 9 12 13 9
16 0 13 10 12 9 7 10 12 9 10 1 10 9 10 9 13
17 7 16 15 15 13 13 9 13 1 10 9 15 7 13 10 0 15
10 7 16 15 13 15 13 3 13 15 13
35 0 13 9 13 10 9 16 3 9 13 10 9 10 9 15 7 9 13 1 10 9 13 15 1 9 7 13 10 9 1 15 9 3 3 13
23 7 10 9 15 1 10 9 10 9 10 0 15 13 3 11 7 11 3 3 10 9 15 13
26 7 10 13 1 10 9 13 1 15 7 13 7 9 13 15 16 0 10 12 9 13 10 13 1 10 9
29 7 1 10 12 9 7 0 9 9 1 10 9 13 1 15 7 13 1 10 9 15 7 9 0 13 1 10 13 15
9 7 13 9 0 1 10 9 13 15
2 13 3
14 7 13 1 10 9 1 10 9 7 13 15 10 0 15
35 7 1 0 10 9 13 9 0 7 10 0 10 9 13 7 13 1 10 9 9 9 9 12 7 10 0 0 13 7 13 9 10 9 10 9
5 10 9 10 0 13
8 7 13 9 0 1 10 9 13
19 13 10 9 10 9 10 9 15 7 10 11 15 7 13 1 10 9 10 9
24 7 10 12 0 10 1 10 9 15 13 1 10 9 15 13 1 10 9 15 7 13 10 9 13
66 13 15 9 10 9 10 9 10 13 7 10 13 7 16 13 10 9 15 10 0 7 13 7 10 9 13 7 13 10 9 15 7 10 9 10 0 13 7 13 10 9 10 9 15 10 9 7 10 0 7 10 13 10 9 15 10 0 7 10 0 7 13 10 13 10 9
21 7 13 10 9 10 9 10 1 10 9 7 13 10 9 10 9 15 1 10 9 15
12 7 13 9 7 9 7 9 7 9 7 9 0
7 7 9 0 13 1 10 9
29 9 13 10 9 7 10 9 1 10 9 15 7 1 10 9 15 9 9 12 7 1 9 13 7 13 13 7 13 13
17 7 10 9 13 1 10 9 10 13 13 16 3 13 10 9 15 13
13 7 13 9 0 15 13 13 15 10 9 1 9 0
13 7 13 10 9 15 1 10 9 7 1 10 9 15
21 7 10 9 13 1 10 9 3 13 3 9 13 1 10 9 16 3 13 15 9 12
16 7 13 9 1 10 9 10 11 7 10 9 15 13 1 10 9
19 7 10 9 13 7 10 9 15 7 3 13 7 9 13 15 3 1 10 9
11 13 1 10 9 7 10 9 15 1 15 13
8 7 13 9 0 1 10 9 13
9 1 0 13 9 7 10 1 15 13
20 6 10 9 7 10 9 16 13 10 9 1 15 13 9 0 13 16 0 9 13
17 7 16 13 10 9 16 13 1 10 9 13 10 9 15 13 10 0
33 7 13 10 9 10 12 9 10 9 10 0 16 13 1 10 0 1 10 9 15 3 13 3 9 7 9 7 0 9 1 9 10 9
18 7 13 10 9 1 10 9 15 1 10 9 9 3 9 16 15 0 13
25 7 13 10 9 10 9 7 13 10 9 10 9 15 7 13 10 9 15 13 10 9 1 10 9 15
28 7 13 10 9 1 10 9 7 13 13 9 1 10 0 10 9 15 10 13 10 9 10 9 7 13 10 9 11
27 7 13 1 10 9 9 13 13 9 12 7 9 12 7 1 10 9 15 12 9 7 1 10 9 15 9 9
15 7 13 15 10 9 10 9 15 7 10 9 15 7 9 0
23 7 13 0 10 9 1 10 9 7 13 10 9 16 13 10 9 10 9 7 13 10 9 13
10 15 0 10 9 7 15 13 13 1 15
15 7 13 15 9 13 0 7 9 7 13 15 9 13 9 12
23 7 13 10 9 15 1 9 1 10 9 13 10 9 15 7 10 9 15 10 1 10 9 13
24 7 13 15 13 9 1 10 0 7 13 15 7 13 15 9 1 15 9 7 9 7 9 7 9
5 16 15 13 9 13
7 16 15 1 9 1 9 13
9 3 13 10 9 7 10 9 10 0
18 7 13 0 9 13 1 10 9 7 13 9 12 0 9 7 13 3 9
10 7 10 9 10 0 9 15 13 1 15
22 7 13 10 9 7 10 1 15 13 16 13 10 9 10 0 15 13 10 9 10 9 15
18 7 13 9 0 16 3 9 13 13 1 10 9 1 10 9 1 10 9
27 7 13 15 13 9 10 9 10 9 16 3 13 10 9 10 9 7 13 15 3 3 13 10 9 10 9 13
58 7 13 15 10 0 7 10 0 7 10 0 7 10 0 7 10 0 7 10 9 16 13 15 9 1 10 9 15 10 0 7 1 10 9 15 16 3 15 13 13 7 13 3 3 10 13 10 9 10 9 10 9 7 10 9 10 9 15
4 3 10 9 13
4 9 3 9 13
5 7 10 9 15 12
31 7 13 7 6 10 9 13 1 10 9 11 7 1 15 12 9 13 10 9 15 7 10 9 10 9 15 13 1 10 9 15
27 7 13 9 1 10 9 3 9 9 0 7 3 9 9 0 7 10 9 15 13 3 9 13 1 10 9 15
16 7 15 13 13 10 9 3 3 10 12 9 10 13 1 10 9
7 0 13 15 1 9 3 13
3 9 3 13
8 0 10 13 10 9 3 3 13
3 0 3 13
31 7 13 0 9 13 1 9 13 9 0 13 1 10 13 1 10 9 7 1 15 9 7 9 7 9 7 9 13 1 9 0
29 13 10 9 7 13 15 9 16 13 10 9 10 9 15 7 13 10 13 10 9 7 10 9 7 10 9 7 9 9
1 13
17 13 11 10 0 15 1 10 9 10 9 10 9 15 13 15 10 9
10 7 0 9 0 13 15 13 1 9 0
53 16 15 13 10 9 7 10 9 15 7 13 9 1 10 9 15 7 1 10 9 15 3 15 13 1 10 9 10 9 10 9 10 13 0 1 10 9 10 9 15 7 13 1 9 7 9 1 9 0 7 1 10 9
34 7 10 9 10 9 15 1 9 9 13 7 3 13 9 9 7 9 10 13 10 9 7 10 9 15 7 16 15 13 10 9 10 9 15
7 7 13 9 1 10 9 13
1 13
1 6
3 13 10 9
7 10 3 9 15 13 1 15
28 7 13 7 6 9 0 7 1 10 9 13 0 9 9 13 1 10 9 15 9 0 7 1 10 9 15 9 0
16 7 0 9 13 1 10 9 13 1 9 0 10 13 1 10 9
17 13 10 9 15 7 13 16 13 10 9 13 16 13 10 9 10 9
16 7 0 9 13 1 10 9 10 1 10 9 13 3 0 9 0
19 13 15 10 9 10 0 7 13 10 9 10 9 10 9 16 13 10 9 15
27 7 13 10 9 10 9 15 1 10 9 7 13 10 9 10 9 7 13 1 10 9 10 9 10 9 10 0
21 7 13 10 9 1 10 9 7 13 9 1 10 9 1 10 9 10 9 1 9 12
25 7 13 0 9 1 10 9 0 7 0 9 12 13 9 12 10 0 16 1 15 13 10 9 10 9
35 7 13 3 9 0 13 9 7 10 13 1 10 9 7 1 10 9 15 7 1 10 9 10 9 15 13 1 10 9 10 0 13 9 10 9
15 7 13 10 9 11 10 9 10 9 7 10 9 10 9 13
11 0 7 0 10 9 15 9 10 9 10 9
3 3 0 0
9 3 15 10 9 13 7 13 1 15
5 3 10 9 15 13
39 7 1 0 13 7 13 10 9 10 9 10 9 1 10 9 7 13 10 12 9 10 13 10 12 9 1 10 9 13 9 0 0 7 13 1 10 9 9 0
25 7 12 1 10 12 9 13 10 12 9 12 9 0 13 10 9 10 9 10 13 1 10 9 10 9
30 7 13 10 9 9 1 10 9 10 9 7 1 10 9 15 7 15 13 13 1 10 9 16 13 10 12 9 10 12 9
11 7 13 0 9 1 10 9 13 10 12 9
13 13 7 13 10 12 9 10 9 10 9 1 10 9
21 7 13 9 0 7 0 1 10 9 10 13 10 9 10 9 7 10 13 10 9 15
10 7 10 0 13 10 9 15 1 10 9
14 7 13 9 3 0 7 15 9 9 13 10 1 10 9
15 7 10 0 13 10 9 15 1 10 9 7 10 9 10 9
3 7 13 9
7 7 13 10 9 10 9 13
23 0 13 10 13 7 10 13 10 0 16 0 13 16 9 0 7 9 13 7 9 15 13 13
2 0 13
10 7 10 0 13 10 9 15 1 10 9
8 7 13 15 13 10 9 1 9
26 7 13 10 9 9 0 7 13 10 9 10 9 10 13 10 9 1 10 9 0 7 3 13 13 15 9
12 7 10 0 13 10 9 15 1 10 9 10 9
36 7 13 10 9 15 13 7 13 10 9 15 1 10 9 7 13 10 9 10 9 1 10 9 15 7 1 10 9 15 7 3 13 1 10 9 15
13 7 10 0 13 10 9 15 1 10 9 10 0 11
15 7 13 10 9 15 16 13 10 9 10 9 10 1 9 9
27 13 3 9 9 13 9 15 13 1 10 9 10 9 0 13 15 1 10 9 10 9 10 0 10 9 10 9
3 13 3 9
17 0 10 13 7 13 10 9 15 16 3 0 13 7 13 10 9 15
10 7 13 15 1 10 9 10 13 3 11
10 7 10 0 13 10 9 15 1 10 9
11 7 13 9 0 1 10 9 1 10 9 13
1 13
15 7 13 10 9 10 0 1 12 9 7 10 9 10 9 13
19 7 11 10 0 13 1 10 9 13 15 10 9 10 9 10 9 10 9 15
12 7 9 0 3 0 13 1 10 9 1 10 9
18 7 13 10 9 10 9 1 10 9 10 9 16 0 13 10 9 15 3
17 7 13 12 1 10 12 9 10 13 10 12 9 7 13 1 15 13
35 6 13 15 10 9 10 9 10 0 10 13 1 10 9 10 0 1 15 13 10 9 10 9 7 13 10 13 10 9 1 10 9 10 9 15
7 7 13 15 1 0 1 9
39 7 10 9 13 13 0 7 0 7 13 9 7 9 0 7 9 13 9 0 1 10 9 15 13 9 7 10 0 10 9 15 7 1 10 9 15 9 13 9
17 7 13 10 9 13 1 10 9 10 0 7 1 10 9 10 9 11
6 7 13 13 15 9 0
3 1 15 13
22 15 15 13 10 9 10 9 7 10 9 10 13 15 10 13 10 12 9 7 10 12 9
18 10 9 15 13 13 7 3 13 7 13 13 1 10 9 7 1 9 13
30 7 13 10 13 1 10 9 15 3 13 10 9 1 10 9 10 9 1 9 9 13 10 9 16 13 7 3 13 7 13
12 10 12 9 12 9 13 3 10 9 13 1 15
4 7 9 12 13
3 10 12 13
3 10 12 13
21 7 10 9 15 13 7 3 13 3 0 0 13 7 1 10 12 13 7 1 9 13
23 7 10 12 9 15 13 12 9 13 15 9 3 13 7 9 3 9 12 9 13 1 10 9
14 0 12 9 13 7 10 9 7 10 9 15 10 9 13
16 10 9 15 13 3 10 9 13 9 7 9 13 7 9 7 9
28 7 10 12 9 15 13 7 10 9 0 13 10 9 7 13 13 15 7 0 7 10 9 15 13 7 15 13 9
29 10 3 9 13 1 10 9 15 13 10 9 15 7 13 12 9 7 13 10 9 15 10 9 16 13 10 9 10 9
18 7 10 9 15 13 13 10 9 10 0 10 13 9 1 10 9 10 9
20 1 0 13 0 9 13 1 10 9 13 9 0 7 10 9 13 1 10 9 15
1 13
53 13 11 10 0 7 13 9 9 7 9 15 9 0 7 9 15 9 0 7 13 16 1 10 9 10 9 10 9 15 13 15 10 9 7 10 9 10 9 1 15 13 7 10 9 10 9 1 10 9 10 9 15 13
20 13 10 9 15 1 15 16 3 13 10 9 15 7 1 10 9 15 16 3 13
15 3 13 15 10 9 1 10 9 7 13 10 9 10 9 15
14 13 15 3 3 15 13 7 13 10 0 1 10 9 15
8 1 10 9 15 13 13 15 0
11 15 13 15 7 13 0 13 15 9 7 9
7 3 1 10 9 15 13 16
18 1 0 1 12 9 13 10 9 15 9 7 9 7 9 7 1 9 13
33 7 13 7 13 1 15 10 9 10 9 10 1 15 13 7 13 3 13 10 9 10 9 15 1 3 13 1 10 9 10 9 15 13
11 6 6 10 9 10 0 11 10 9 10 0
7 3 12 9 13 10 9 15
85 7 10 9 10 9 13 7 13 1 15 16 10 9 15 15 13 3 9 9 7 9 7 9 0 7 9 7 0 7 9 7 0 7 0 7 15 9 0 7 15 9 0 7 15 9 1 9 0 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 9
27 7 10 9 15 10 9 10 9 13 1 15 7 15 10 0 7 10 0 13 1 15 7 3 3 3 15 13
20 10 9 0 10 13 1 15 1 3 13 1 10 9 10 9 15 13 7 13 13
29 6 6 10 9 10 0 10 13 0 7 0 7 0 7 13 1 9 7 9 0 7 9 16 12 9 13 10 0 9
25 6 6 10 9 10 0 1 15 13 15 10 13 10 9 1 10 9 1 10 9 15 16 12 9 13
22 13 1 15 9 7 10 0 7 10 9 7 10 9 16 13 10 9 10 9 15 1 15
15 7 13 12 9 0 9 3 9 0 7 13 1 10 9 13
12 3 9 13 11 10 0 9 7 3 3 13 3
55 7 9 9 7 0 7 9 7 9 3 3 13 1 15 3 7 15 9 15 9 3 3 13 1 15 3 7 9 9 3 3 13 1 15 3 7 9 9 3 3 13 1 15 3 7 9 9 7 9 3 3 13 1 15 3
33 3 10 9 15 13 10 9 10 9 16 1 10 9 15 13 15 10 9 7 1 15 9 9 7 0 13 7 15 10 13 1 10 9
39 11 9 9 9 0 16 7 10 13 1 9 10 9 0 13 7 9 0 7 7 0 15 3 9 15 3 9 13 0 13 10 7 15 7 1 15 9 13 15
11 9 3 3 10 9 9 0 13 13 10 9
15 10 3 11 0 10 9 13 0 10 1 10 3 11 13 9
12 13 3 10 9 1 3 10 11 0 13 10 9
26 0 3 7 0 9 1 15 13 13 15 3 15 13 1 10 9 9 0 7 0 7 3 3 10 9 9
15 10 3 15 9 13 1 10 15 0 3 9 13 11 10 11
14 0 13 1 9 10 9 13 10 9 15 15 13 9 3
7 7 10 9 13 13 1 15
13 10 3 3 0 10 9 13 10 3 11 1 15 13
9 13 3 1 10 9 13 13 1 11
5 13 3 3 0 9
17 0 3 3 0 1 0 15 13 1 3 0 9 0 10 0 9 13
27 13 3 0 9 1 11 7 10 11 7 1 11 9 3 13 3 10 15 15 1 13 13 10 9 10 9 11
18 13 3 10 9 9 1 10 11 9 13 7 9 10 9 7 13 10 9
14 15 3 13 16 3 0 11 10 0 13 15 9 10 9
5 3 3 15 13 0
26 0 3 13 9 1 0 11 10 11 13 0 13 15 1 10 11 1 9 13 9 13 3 16 3 13 9
19 3 3 13 15 11 10 9 13 0 13 9 13 7 11 7 9 10 9 13
18 1 3 3 0 9 0 13 1 15 10 3 1 0 9 3 3 0 13
12 0 3 13 13 1 10 11 3 15 1 10 11
24 10 3 3 13 9 9 0 13 9 13 10 3 13 9 13 13 0 10 3 15 9 13 13 13
11 0 3 3 16 16 3 0 13 3 3 13
33 15 3 3 0 1 10 11 13 9 13 10 9 9 15 13 9 3 0 1 9 9 0 13 7 3 13 1 10 11 10 11 9 13
9 1 0 3 13 10 0 15 13 0
8 10 3 11 7 10 0 13 13
21 3 3 9 13 13 7 1 10 11 9 13 15 13 10 9 10 9 10 1 10 9
20 3 3 9 15 13 13 13 15 1 11 7 16 1 10 11 13 10 9 10 9
20 16 3 13 0 13 13 10 9 3 3 3 15 10 9 13 16 3 3 0 13
8 0 3 3 9 7 7 9 13
15 15 3 1 3 0 3 13 13 16 3 7 3 3 0 13
26 15 3 13 0 0 13 0 9 1 10 9 0 13 13 1 10 3 10 9 3 0 7 0 9 9 13
9 15 3 1 15 13 0 0 13 0
13 10 0 3 13 9 0 1 10 0 13 13 15 3
33 11 13 9 3 9 9 3 11 9 3 9 10 1 11 9 15 13 1 9 1 0 7 7 9 13 1 9 9 1 10 0 13 11
4 15 3 9 13
12 13 3 9 7 7 9 7 9 10 1 10 11
4 9 3 13 0
9 1 3 10 11 9 15 9 13 0
15 10 3 9 3 13 13 9 1 10 9 10 11 13 3 9
14 13 11 15 10 9 11 13 9 11 9 3 11 10 11
19 11 3 3 10 11 10 11 10 11 0 9 9 13 11 11 3 10 11 0
25 10 3 0 9 13 0 10 9 13 9 9 10 11 1 15 10 9 0 13 10 15 0 0 9 13
9 0 3 3 10 11 13 10 15 9
9 13 3 13 15 13 9 0 15 0
33 3 3 0 13 13 3 15 10 9 11 10 11 13 3 0 10 11 3 10 0 10 9 13 10 11 3 3 3 10 9 10 9 13
13 11 3 3 15 13 13 15 13 1 10 9 10 9
7 9 3 13 9 13 0 9
5 13 16 0 13 0
4 15 3 13 13
13 9 15 13 9 3 0 13 15 9 10 15 13 0
10 3 3 10 0 9 13 1 15 13 13
9 1 15 12 0 13 13 15 10 15
14 15 3 3 13 0 13 13 16 15 15 1 15 13 0
4 15 3 13 0
24 13 11 7 16 13 7 15 16 15 13 13 9 0 7 9 10 15 16 15 15 1 15 13 9
12 9 3 15 13 3 16 7 13 15 13 1 15
14 15 3 15 1 10 9 1 15 13 1 10 13 9 13
12 1 3 15 13 13 3 10 9 10 15 1 9
16 1 0 10 9 1 12 0 13 13 7 1 9 0 13 15 13
9 15 3 3 16 3 13 13 13 0
15 10 3 11 16 13 9 10 9 13 13 10 11 1 10 9
8 7 1 0 3 13 3 10 9
9 13 3 7 13 10 9 13 10 11
20 16 3 1 9 13 13 10 9 1 10 9 13 13 3 7 10 9 13 15 13
19 13 3 10 13 1 10 9 7 13 13 7 13 13 1 9 13 13 10 11
19 1 3 10 9 3 3 3 1 10 0 9 3 9 13 0 1 9 0 13
10 15 3 15 13 15 10 13 13 13 13
9 13 3 3 3 3 10 9 13 13
9 16 3 10 11 13 13 10 9 0
8 3 15 12 9 13 11 13 9
3 15 13 13
32 7 3 11 13 15 7 7 10 9 13 10 9 7 0 15 3 3 13 13 16 3 3 15 13 11 10 0 13 15 3 15 13
19 7 7 0 3 10 0 13 13 13 7 15 10 15 0 13 7 13 3 13
8 10 3 11 3 3 13 10 13
17 3 3 13 7 13 9 3 13 7 10 9 13 7 0 1 0 13
3 13 0 13
4 13 3 13 0
16 16 15 13 9 10 15 13 3 13 13 13 15 3 9 13 15
4 15 3 13 13
15 1 10 0 3 9 10 9 13 3 3 3 0 15 13 0
5 13 3 10 9 13
40 16 3 13 10 9 9 13 3 3 13 10 11 7 15 13 9 15 7 13 7 15 13 7 11 13 1 10 9 10 9 7 15 0 9 13 13 1 10 0 9
9 13 7 3 10 9 7 13 3 11
14 0 3 13 10 11 16 9 9 13 1 10 0 0 11
15 0 10 9 9 7 7 10 9 15 9 15 13 16 3 13
11 10 3 3 9 3 13 10 9 10 9 13
19 11 3 13 13 9 1 11 3 0 7 15 3 9 9 13 15 0 1 11
16 1 3 10 9 9 0 13 0 7 3 15 3 9 0 13 13
6 9 15 9 12 0 13
15 0 3 9 13 3 0 10 0 13 10 9 7 11 10 11
14 13 3 3 7 11 10 0 9 1 15 13 13 13 0
11 13 3 10 9 0 3 3 10 10 11 9
19 10 3 9 0 7 10 9 15 10 11 13 1 9 13 9 1 10 13 9
19 13 3 3 9 3 0 16 13 1 7 11 7 1 11 7 11 10 9 13
14 7 15 3 0 1 15 15 9 13 13 12 13 12 9
5 0 3 13 0 13
32 0 3 11 7 13 1 11 7 13 1 0 7 13 11 0 1 9 1 9 10 9 13 13 1 10 11 7 11 3 10 9 13
18 11 3 13 12 13 12 9 13 11 10 11 7 13 9 12 11 3 11
11 1 3 3 0 3 3 13 13 7 13 3
10 0 3 9 13 13 1 10 9 3 0
8 13 0 13 10 9 1 10 9
7 13 3 13 10 11 9 0
12 16 3 13 1 10 9 9 0 3 13 10 9
19 16 3 1 10 0 13 9 3 10 1 10 9 7 13 7 13 7 9 13
5 13 3 1 9 13
16 15 3 10 7 9 7 10 9 10 1 10 9 16 13 13 3
30 10 3 9 3 13 10 9 0 1 16 13 3 13 10 9 13 7 7 13 10 0 15 3 0 13 13 15 3 13 13
23 0 13 13 9 12 1 15 9 0 0 0 13 1 7 11 9 10 15 13 7 1 11 9
22 10 3 3 12 9 10 12 11 10 11 3 9 13 10 3 13 3 1 10 0 10 9
9 11 0 3 3 10 10 9 13 13
13 10 3 0 0 9 10 9 0 13 3 3 9 0
6 0 3 10 0 13 13
13 3 3 3 0 10 0 10 9 10 1 0 9 13
14 10 3 0 9 9 13 1 10 9 13 15 0 13 9
5 13 3 10 9 13
7 7 10 3 3 9 15 13
10 1 3 10 9 13 1 11 13 10 11
15 7 3 13 15 7 3 15 13 13 10 9 13 1 10 9
24 15 3 10 11 13 1 11 3 13 13 16 3 10 9 10 11 13 15 13 9 10 0 1 11
6 9 13 15 3 13 13
36 0 3 0 13 0 11 10 11 13 11 10 3 11 13 9 1 10 3 13 10 9 10 10 11 13 13 9 13 16 3 15 13 1 10 13 13
6 0 3 3 3 13 13
8 10 3 3 9 1 10 11 13
14 11 3 3 13 15 9 7 13 15 11 13 13 13 0
30 0 3 13 7 7 13 11 0 1 16 3 3 10 9 10 0 13 7 9 0 9 13 7 10 9 1 9 13 13 11
4 15 3 7 13
29 16 3 3 13 7 0 10 9 7 13 1 11 10 9 10 9 13 1 10 11 3 15 13 1 15 15 13 10 9
33 13 3 10 11 9 7 13 0 1 10 11 7 10 9 13 1 10 0 0 13 10 9 13 1 10 11 10 0 9 3 3 15 13
29 3 3 10 7 9 15 13 1 15 7 9 15 13 7 9 7 12 7 1 12 9 10 11 13 10 11 1 10 11
6 15 7 1 10 9 13
12 11 3 13 11 9 0 10 10 11 10 9 13
44 15 3 13 0 13 3 15 0 1 10 9 9 0 13 11 10 0 1 9 13 1 11 13 9 10 3 13 15 0 7 9 0 9 15 15 13 13 7 7 13 7 13 1 11
27 0 10 11 13 10 0 10 9 13 1 11 13 13 1 11 7 7 11 13 3 9 0 13 3 1 11 13
15 13 3 3 1 11 13 3 0 3 3 0 13 9 9 0
12 15 3 1 10 9 13 10 11 13 13 10 9
12 15 3 13 0 13 9 3 15 13 9 3 13
26 3 3 13 15 0 7 13 10 9 7 15 13 15 16 3 9 1 9 13 7 13 1 10 9 10 0
22 13 3 10 11 1 9 13 16 15 3 13 13 15 1 10 9 15 13 1 10 9 13
7 13 1 10 9 1 0 9
35 15 3 13 7 15 10 9 7 13 10 9 13 1 10 9 13 9 10 0 13 3 10 9 13 15 1 10 9 15 3 13 1 10 9 15
6 7 15 3 13 1 11
8 15 3 9 13 13 13 1 11
15 13 3 15 13 1 11 1 10 9 7 13 13 15 10 13
16 11 3 1 9 11 3 1 9 13 3 13 3 3 13 10 9
12 16 3 3 13 15 13 13 16 15 13 1 11
8 7 15 13 3 13 3 13 13
13 7 11 13 9 0 3 0 1 11 1 9 13 9
16 11 3 10 9 10 1 0 9 13 3 13 13 9 12 7 12
40 13 3 13 10 9 0 0 10 9 0 1 11 9 7 0 0 7 9 0 0 9 0 1 15 10 1 11 9 11 10 9 9 15 0 3 15 9 9 9 13
15 13 3 11 13 10 9 11 10 11 9 13 9 12 7 12
6 15 3 9 0 13 9
20 3 3 10 0 13 1 15 13 10 9 10 11 13 1 10 9 9 1 10 9
15 13 3 1 10 7 0 9 15 3 13 7 10 9 12 9
33 0 3 3 0 13 10 11 3 3 1 9 0 9 7 7 9 15 15 9 13 15 3 13 0 13 0 13 15 3 15 3 0 13
16 6 9 9 9 13 0 1 11 7 7 1 15 1 9 13 13
7 11 3 13 13 0 0 13
14 10 3 0 9 13 1 9 9 13 1 9 9 1 9
4 15 3 13 13
13 6 9 3 15 13 13 9 13 13 1 9 9 13
16 3 7 13 11 10 9 7 15 3 3 13 13 13 13 10 9
9 7 3 10 10 9 13 9 9 13
20 13 3 0 9 9 9 9 9 9 9 10 9 7 7 9 9 9 9 9 9
9 0 3 3 0 7 13 15 13 0
13 9 3 0 13 12 9 13 9 15 3 15 11 13
23 0 3 3 0 7 10 9 13 10 11 1 1 11 13 1 11 7 3 3 1 11 1 11
9 13 3 13 1 10 9 1 10 11
23 3 3 9 0 7 0 13 11 10 11 9 13 1 10 9 7 13 15 13 0 7 7 0
16 13 3 15 10 15 7 13 3 15 1 9 13 13 10 11 0
13 3 3 13 15 9 13 15 16 15 3 15 13 0
8 15 3 13 13 9 0 0 13
4 6 9 11 0
7 13 3 11 10 13 13 3
6 15 3 13 11 13 0
3 15 3 13
22 11 0 3 10 9 3 13 9 13 0 7 7 0 7 15 13 0 9 13 7 15 13
17 13 3 0 9 1 10 0 1 11 13 7 9 13 10 0 13 0
13 7 15 0 0 7 13 3 3 3 13 7 13 3
27 16 3 10 1 10 11 13 10 11 10 11 13 0 7 7 0 13 15 0 1 0 13 13 3 0 3 13
4 11 7 7 11
15 0 3 13 9 0 9 7 13 13 7 1 0 9 9 0
12 0 7 0 3 13 7 3 3 13 0 10 9
16 13 9 10 11 10 0 13 3 10 9 15 9 13 1 10 9
14 13 3 10 9 10 9 13 0 1 10 9 13 10 9
8 1 10 9 3 15 13 10 9
10 9 3 12 7 12 13 13 1 10 9
14 0 3 15 13 7 13 1 10 9 9 10 9 0 13
3 0 9 13
35 10 3 9 0 13 10 7 9 7 10 9 13 0 10 9 13 11 7 7 11 10 15 9 15 15 13 3 10 9 13 15 9 13 0 13
24 1 0 3 10 9 16 13 7 7 13 13 1 0 10 9 10 9 3 13 7 1 9 0 13
7 11 3 3 9 0 13 0
4 11 3 13 13
20 6 9 0 10 3 15 9 3 15 13 1 10 15 16 7 9 9 0 15 13
3 15 3 13
16 6 11 13 15 10 9 15 13 0 7 7 0 13 0 9 1
9 1 3 12 9 9 10 9 9 13
15 0 13 9 12 13 9 12 7 12 7 12 0 9 3 13
29 0 10 0 9 10 1 10 12 9 13 12 7 12 7 12 7 12 10 0 15 10 0 9 10 3 15 0 13 9
7 3 3 11 15 13 9 9
12 15 3 15 7 13 0 13 7 9 0 13 9
15 0 3 15 13 15 3 15 15 13 16 13 3 10 9 13
25 3 3 15 0 0 0 3 10 1 9 13 0 13 16 3 15 9 13 15 0 13 3 13 10 9
13 0 3 3 0 9 0 13 0 3 3 13 9 0
10 15 3 9 13 7 9 0 13 13 0
19 16 3 1 0 3 13 10 9 3 0 0 15 15 13 10 0 13 0 13
11 16 3 3 13 13 7 13 3 0 7 0
24 10 15 3 3 0 13 9 13 0 13 3 9 15 13 15 15 13 7 15 3 13 0 3 13
8 15 3 3 10 0 13 0 0
9 3 3 3 9 9 12 15 0 13
4 15 3 3 13
4 0 3 0 13
9 0 3 3 13 9 10 9 0 13
29 0 13 10 11 3 3 7 13 7 9 15 13 15 13 3 13 0 13 15 10 13 0 13 10 9 15 9 13 13
19 1 3 11 13 13 1 9 9 0 11 3 13 16 13 15 13 9 0 0
18 3 3 15 13 13 9 15 15 10 9 13 10 13 13 0 1 10 9
24 13 3 10 11 12 9 15 10 0 3 13 13 3 3 0 10 3 0 10 9 0 10 15 0
5 9 3 15 13 11
16 0 3 3 10 11 13 10 11 10 9 16 13 15 9 0 13
16 15 3 16 13 7 15 9 13 13 10 9 13 3 10 9 9
28 9 3 7 9 7 10 0 15 15 13 1 9 9 1 10 9 13 1 10 9 13 16 15 15 13 10 9 13
14 13 3 0 1 10 11 9 1 9 10 0 0 13 13
4 11 3 15 13
10 13 3 0 10 9 10 9 7 10 9
15 16 3 10 13 13 10 11 13 3 7 7 15 13 13 0
13 6 9 15 7 13 7 3 10 11 13 0 15 13
6 15 7 9 7 9 13
3 15 3 13
14 13 3 9 15 0 13 13 7 1 10 9 7 13 15
5 11 3 15 13 0
25 9 7 0 13 0 13 7 13 1 9 3 13 9 15 13 1 15 9 7 0 3 0 13 13 0
7 15 3 3 9 13 1 11
14 1 3 10 0 9 0 1 10 0 11 9 9 13 0
12 13 3 0 1 10 9 0 10 10 9 9 13
11 3 3 10 9 1 15 13 13 3 0 15
11 9 3 13 1 10 11 10 9 9 13 0
5 0 13 13 3 13
20 3 3 13 15 10 9 7 9 9 7 9 13 15 16 3 15 13 1 10 9
5 15 3 3 0 13
10 11 3 13 10 9 10 9 13 15 0
8 9 3 1 10 15 3 13 3
5 3 3 3 15 13
22 9 3 9 7 10 9 15 13 7 13 10 13 13 3 0 13 15 10 9 1 10 9
2 0 13
16 3 13 3 10 11 10 3 9 15 13 13 1 15 10 9 0
18 6 9 10 0 0 3 7 0 15 13 1 7 9 7 1 9 13 13
14 3 3 15 15 0 13 13 7 15 9 15 13 7 9
14 3 7 15 15 13 9 1 7 9 7 1 9 13 13
13 15 3 15 10 9 13 13 15 3 15 10 0 9
19 15 3 15 7 13 13 1 10 9 7 9 13 16 15 0 13 0 3 13
3 13 11 0
24 6 9 7 9 7 15 15 0 13 15 13 0 7 15 9 9 1 10 9 13 13 15 0 13
28 1 3 10 9 0 10 7 9 15 0 13 7 1 10 13 3 13 9 13 16 3 13 1 10 15 15 9 13
7 12 3 15 0 13 13 9
11 10 3 3 0 13 10 9 3 13 15 13
4 13 10 9 0
14 15 3 3 13 7 13 15 10 9 15 15 0 13 13
10 13 15 10 9 1 9 0 13 15 13
13 9 3 15 3 13 9 15 3 9 0 15 15 13
22 16 3 3 1 9 15 13 13 15 7 0 15 15 15 0 13 13 3 15 13 15 13
11 16 3 3 1 9 15 13 10 9 13 15
2 13 11
11 6 9 13 3 15 13 9 13 1 10 9
9 13 3 0 10 11 13 10 9 11
5 13 3 15 13 0
18 11 15 15 9 13 0 15 15 3 13 13 7 9 13 13 13 15 9
32 3 3 13 3 15 13 0 1 15 0 15 13 9 9 15 10 15 13 13 1 9 13 16 15 1 9 9 0 1 9 13 15
13 1 3 0 7 15 3 0 13 13 3 13 10 9
3 13 10 11
11 6 9 3 3 15 3 3 13 1 9 0
18 3 3 16 15 13 7 13 15 13 13 3 15 13 0 13 13 0 0
13 9 7 15 15 13 13 0 10 13 1 13 15 13
14 0 16 0 13 11 13 1 0 13 9 7 9 7 9
10 13 3 1 10 11 10 9 13 10 9
7 13 3 7 13 15 9 13
19 3 3 10 9 0 3 10 13 10 9 13 3 11 13 10 9 15 3 13
11 15 3 3 13 10 9 13 10 9 10 9
15 13 3 1 10 11 10 7 9 7 10 10 9 9 13 15
18 10 3 11 10 9 10 9 13 3 15 13 16 15 13 15 0 9 13
51 13 3 10 9 3 13 3 1 0 13 15 1 10 9 13 13 13 3 0 7 7 0 10 0 0 13 9 10 3 0 13 16 3 9 13 10 9 9 10 9 13 13 10 3 0 16 9 13 15 13 0
35 13 3 0 1 10 9 13 15 11 13 10 9 13 15 13 10 9 13 10 7 0 15 9 7 16 1 0 10 13 13 13 7 15 13 0
18 11 3 0 13 10 7 11 13 3 13 1 0 0 0 7 13 1 15
12 13 6 9 1 15 15 10 9 16 15 13 9
26 12 3 3 15 15 0 10 0 0 16 3 15 0 13 7 9 3 15 15 15 3 3 13 10 13 13
12 11 3 1 12 9 1 9 0 13 10 9 13
22 3 3 10 11 10 11 9 13 1 11 10 11 7 10 10 9 9 13 9 3 11 13
17 13 3 1 9 16 3 13 16 0 13 10 9 13 15 13 10 9
35 1 3 10 9 0 3 13 10 9 10 7 1 9 7 10 1 11 13 0 3 15 3 1 11 13 15 3 1 11 10 9 15 3 1 11
16 15 3 15 13 1 7 9 7 1 11 15 3 10 0 1 11
11 0 3 3 10 0 9 1 15 13 13 11
7 11 3 1 11 13 15 13
23 13 3 13 10 9 15 15 13 16 16 13 10 9 13 13 15 0 13 16 13 1 9 13
11 15 3 3 0 10 9 13 13 13 1 15
13 15 15 3 3 10 0 10 9 13 3 13 1 0
25 1 3 11 16 13 0 1 10 9 10 9 13 10 9 7 13 10 13 10 11 1 0 9 13 0
16 13 3 15 9 7 9 7 9 9 7 0 13 7 3 13 13
13 9 15 1 9 13 0 9 13 1 9 1 0 9
4 15 9 3 13
3 9 3 13
12 0 10 9 13 10 11 13 13 13 1 10 11
21 13 15 13 0 13 7 7 13 9 7 9 13 3 13 0 1 9 0 0 9 13
9 10 3 3 1 11 3 10 11 13
37 1 3 10 11 10 9 9 3 13 13 15 15 10 9 13 13 1 10 9 10 13 3 3 3 7 0 13 15 3 3 16 3 0 13 9 0 13
10 1 3 0 9 0 10 1 11 9 13
13 9 7 15 13 13 15 15 15 0 15 15 13 0
22 9 3 12 7 12 7 0 0 9 12 0 9 0 13 10 3 15 9 0 9 9 0
11 13 3 3 9 9 9 0 13 9 9 12
5 13 3 15 0 9
36 13 3 3 0 1 10 9 13 7 10 3 0 13 1 10 0 9 13 9 0 9 7 3 12 9 10 3 0 1 10 0 10 9 13 9 12
5 13 3 1 9 11
12 13 3 15 9 11 10 0 9 13 7 15 13
8 3 3 10 13 13 15 9 13
31 3 9 7 0 12 13 15 1 10 0 9 13 7 9 12 13 0 7 7 0 15 10 0 13 0 13 13 9 3 3 13
5 13 3 3 0 11
19 7 10 3 9 1 15 10 9 13 10 9 0 13 3 3 15 3 9 15
31 0 7 9 3 0 0 13 1 0 10 11 7 9 0 0 7 3 3 9 9 0 0 15 9 10 9 10 11 9 13 13
5 0 3 1 11 13
29 10 3 11 13 15 10 7 9 7 10 9 13 9 7 0 15 3 7 9 0 15 0 10 9 10 9 13 3 0
18 10 3 3 0 1 15 13 13 1 11 7 11 1 10 9 10 0 11
30 10 3 13 13 10 9 0 10 9 1 10 9 13 10 11 13 10 9 16 13 1 9 11 7 16 15 9 9 13 9
15 16 3 13 1 15 13 10 9 13 10 9 13 10 9 13
4 15 3 0 13
20 10 3 9 15 1 10 0 10 9 13 13 11 16 13 1 9 0 9 15 13
9 10 3 9 0 13 15 13 9 13
24 9 3 1 0 13 11 7 9 9 7 9 7 9 7 13 10 13 15 13 9 1 10 3 9
9 13 3 10 11 10 11 13 10 0
9 16 3 3 13 10 9 9 13 15
10 13 3 0 13 16 15 0 13 10 9
20 7 3 9 9 9 13 3 3 9 0 0 1 11 13 7 13 7 13 0 13
29 0 13 10 9 10 11 0 15 3 15 13 13 9 0 1 9 13 9 7 3 0 7 10 1 15 13 3 10 9
12 1 3 0 13 13 15 3 9 0 13 13 9
16 13 3 13 0 7 0 13 15 3 10 0 9 15 3 10 0
6 7 15 3 3 3 13
4 15 3 0 3
26 1 3 3 9 9 13 9 10 11 1 3 11 10 9 10 1 10 11 7 7 10 11 9 13 3 11
17 3 3 3 1 10 11 13 7 1 10 11 3 1 11 13 0 13
10 15 3 9 13 10 9 3 13 3 13
67 16 3 0 13 13 13 10 3 3 13 9 10 1 9 11 9 13 15 0 3 13 10 3 9 13 13 3 3 9 10 3 9 13 7 10 11 7 7 11 9 13 1 11 15 0 13 0 7 15 15 0 13 9 10 9 13 16 0 13 13 13 13 10 9 0 9 13
23 16 3 13 3 15 0 10 0 10 0 9 13 0 1 10 9 10 1 9 3 10 9 13
19 7 3 3 7 10 9 0 10 3 15 13 13 0 7 10 9 15 3 0
16 10 3 0 9 3 16 13 3 3 10 0 13 3 15 13 13
27 13 3 1 10 0 13 0 1 0 15 10 9 13 13 1 9 10 9 9 3 13 15 7 15 9 9 0
24 0 3 3 10 9 10 3 0 13 7 7 13 13 10 11 1 11 10 11 0 10 9 13 0
11 11 3 13 9 7 13 10 0 9 13 0
20 13 3 15 10 0 10 9 13 7 9 7 13 0 7 9 1 9 13 7 13
37 11 3 10 0 13 7 13 10 9 13 11 0 3 9 3 13 0 1 10 9 16 3 13 13 0 10 9 13 7 16 15 15 13 13 9 0 13
8 3 0 13 11 13 13 10 11
37 13 15 1 0 10 11 0 15 13 10 0 7 10 1 10 9 0 7 15 3 13 11 10 11 10 3 1 10 9 11 9 13 10 9 13 0 9
23 13 15 7 7 9 13 1 10 9 10 9 3 13 10 0 15 15 13 1 9 13 13 3
22 10 3 9 15 10 0 13 13 15 10 9 13 9 0 15 0 3 3 13 11 0 3
7 9 3 9 13 13 15 3
8 13 3 0 1 11 13 10 9
26 3 3 10 11 13 0 7 9 10 13 13 7 0 13 1 7 10 13 13 10 9 13 3 7 7 3
19 1 3 3 0 9 10 0 13 10 7 10 11 9 7 15 10 11 13 15
15 3 3 9 13 10 0 11 7 10 9 3 3 13 13 13
10 15 3 13 11 3 1 0 1 15 13
24 0 10 9 13 9 1 9 13 7 13 9 15 15 13 0 13 13 13 1 10 9 0 9 13
10 15 10 13 13 13 1 10 9 13 0
6 15 3 3 0 13 13
21 13 3 10 9 9 10 13 10 11 1 10 9 10 1 11 13 13 10 11 10 9
27 15 3 9 7 15 13 9 7 13 0 13 10 9 3 13 15 13 1 10 0 9 9 13 15 3 1 9
8 10 3 3 0 13 0 10 9
15 3 3 7 13 7 3 3 13 10 15 9 15 3 10 9
9 9 3 16 13 13 10 9 10 9
8 13 3 1 11 13 1 10 9
19 11 3 9 13 13 3 10 9 3 13 9 1 10 9 15 15 13 3 15
11 0 3 0 13 9 0 13 10 9 10 9
15 3 3 3 0 9 13 9 13 7 15 15 13 1 10 9
25 7 3 0 0 13 1 11 7 0 15 9 13 9 15 9 13 11 9 0 13 13 7 9 7 9
15 1 9 3 13 1 0 9 13 3 7 0 10 11 13 11
27 1 3 0 10 9 15 13 10 7 1 10 9 9 13 15 7 1 10 9 13 15 10 9 1 9 13 0
4 0 3 3 13
20 3 0 9 13 13 11 11 10 9 0 9 15 15 13 13 1 0 9 0 13
4 13 3 10 9
4 10 3 9 13
6 9 3 13 0 1 9
7 15 3 3 15 13 13 0
13 11 3 13 10 9 7 13 13 10 13 13 10 9
26 0 3 10 1 10 9 1 9 13 13 3 3 7 1 10 9 15 15 15 3 1 9 15 3 1 9
17 13 3 0 9 3 0 11 13 16 7 13 3 10 0 13 7 13
19 15 3 13 10 13 13 10 13 1 11 13 7 13 7 13 0 1 10 15
20 1 15 9 10 9 13 1 0 10 9 15 13 10 0 13 1 0 9 10 11
5 7 11 3 13 11
8 0 3 15 3 1 10 9 13
9 15 3 15 1 9 13 1 10 0
27 10 3 3 0 0 10 9 0 13 10 11 13 10 3 0 1 0 7 0 13 7 13 3 10 9 0 9
18 10 3 3 0 0 7 0 13 3 15 9 1 7 15 10 7 9 0
5 13 3 3 1 9
14 13 6 11 15 1 0 9 11 9 7 15 0 9 13
7 13 7 15 9 13 7 9
8 7 3 3 3 9 13 6 11
17 15 3 3 15 1 0 13 3 13 15 10 11 10 3 13 9 9
18 3 3 0 0 13 11 13 11 9 3 15 13 3 9 1 11 13 0
20 3 3 10 1 9 13 9 7 9 7 9 1 7 0 10 9 7 9 13 11
4 3 3 13 13
8 10 3 11 13 9 13 13 3
6 10 3 11 15 13 0
3 11 15 13
3 0 15 13
3 3 15 13
5 15 3 15 3 13
10 13 15 11 0 13 7 0 9 9 13
11 0 16 13 13 10 0 9 3 10 0 13
15 15 3 9 13 1 9 13 9 0 0 3 3 13 10 9
22 10 3 9 0 1 15 13 3 3 1 15 13 0 1 11 1 10 9 10 9 11 13
13 1 3 3 10 0 9 3 3 3 13 1 10 9
25 1 3 10 1 11 9 7 10 11 7 7 11 9 1 11 3 10 9 0 10 9 13 9 0 13
11 10 3 11 15 13 10 11 10 11 9 13
23 16 3 13 3 0 7 13 10 9 10 11 13 3 10 1 9 13 10 9 1 15 13 11
9 13 3 0 10 0 13 10 11 0
11 3 9 13 0 9 15 15 13 11 9 13
16 10 3 0 13 10 9 13 1 10 9 3 10 0 12 9 0
10 13 3 15 10 9 13 13 13 10 9
25 3 3 3 6 9 9 16 3 13 15 3 15 3 3 13 3 3 3 13 9 13 10 9 10 9
22 1 3 9 3 3 13 0 0 9 10 3 13 15 7 13 10 0 9 0 13 10 9
4 13 3 13 3
8 15 3 3 15 13 15 3 13
15 15 3 13 10 13 13 10 11 1 10 9 0 13 0 13
40 10 9 12 13 9 10 9 13 13 10 3 9 7 10 9 10 7 9 7 10 0 10 3 13 9 10 9 1 9 13 1 0 15 13 16 1 0 9 9 13
9 15 3 1 9 0 13 15 9 13
15 7 1 0 10 9 16 13 15 0 0 10 9 13 10 0
22 0 3 3 15 13 10 11 13 1 11 9 9 7 13 7 13 9 13 7 15 13 13
4 15 3 13 13
12 13 15 11 10 9 7 7 15 9 9 13 0
7 11 3 3 0 1 9 13
23 0 3 13 3 0 10 9 10 11 13 13 7 10 9 10 9 7 13 9 9 1 7 9
11 3 3 15 15 9 13 1 11 0 3 13
21 13 3 10 0 1 11 9 13 1 9 13 13 0 15 3 10 0 1 11 13 11
12 0 10 9 3 13 1 11 1 9 0 13 0
14 3 3 3 3 10 13 13 13 1 11 16 13 1 0
7 1 3 3 10 9 3 13
17 11 3 13 10 9 13 9 1 11 13 13 11 7 7 10 9 9
29 13 3 11 13 1 9 10 15 9 13 3 3 13 0 1 3 0 10 9 7 10 3 9 1 9 13 13 11 0
4 9 15 13 11
28 6 9 1 9 0 13 13 15 0 3 9 0 3 10 0 9 13 13 3 3 15 13 7 15 13 9 13 0
7 3 3 3 9 13 7 13
13 0 3 3 16 13 15 15 13 15 3 3 13 15
8 0 3 16 13 13 15 0 13
9 13 3 10 15 0 13 7 0 13
15 15 3 3 9 13 9 15 3 1 9 13 9 13 1 9
6 0 13 3 13 10 11
11 9 3 16 9 13 13 7 0 7 0 15
7 10 3 9 1 9 0 13
16 13 3 10 0 0 10 3 0 3 9 13 9 0 3 3 11
18 13 3 0 7 13 3 1 9 9 3 3 0 9 13 1 0 3 0
20 3 10 11 9 13 3 15 10 11 10 3 1 9 10 0 11 1 10 0 9
8 13 3 9 0 10 9 0 0
7 9 9 0 9 12 9 13
30 13 3 10 11 1 10 11 0 1 7 9 9 13 1 10 15 9 13 7 3 10 9 0 13 7 13 13 1 11 11
20 11 3 10 11 13 11 3 9 9 3 9 11 10 11 13 13 13 9 11 3
11 9 10 9 9 9 13 13 1 9 10 0
18 3 3 1 0 13 15 9 15 13 10 9 7 13 7 10 9 10 9
17 13 3 15 0 9 10 11 13 3 3 13 9 0 3 3 13 9
45 15 3 0 1 11 13 3 0 15 0 13 13 10 1 15 13 9 12 13 13 3 15 3 13 3 10 9 13 11 13 13 3 9 3 13 3 10 0 13 1 11 10 11 1 11
3 0 7 13
19 7 3 11 7 10 13 9 10 9 0 13 7 10 9 0 13 11 9 13
44 1 3 0 3 3 3 10 11 13 10 9 13 11 9 10 9 7 10 9 13 1 9 12 1 15 3 3 10 9 10 9 13 3 3 10 9 10 9 3 3 3 9 15 13
7 13 3 15 1 0 10 9
24 10 3 9 0 10 9 11 10 0 10 9 13 13 9 13 9 0 1 15 3 3 13 10 9
26 10 3 9 7 7 10 9 16 13 9 1 9 13 10 9 7 13 7 3 15 13 3 0 9 15 13
13 0 15 7 10 9 10 13 13 13 7 9 9 13
11 11 3 13 13 10 9 11 11 10 11 9
9 1 3 9 0 9 0 3 13 13
24 9 3 13 0 10 9 15 3 7 9 7 1 0 16 10 9 13 1 10 9 10 9 13 15
20 0 3 3 10 11 11 13 15 9 13 13 1 9 15 15 1 10 3 9 13
33 16 3 13 1 10 11 9 10 11 10 3 3 3 15 13 1 10 13 9 13 10 9 3 3 10 0 9 9 11 15 10 0 13
45 13 3 11 3 15 13 10 9 10 9 3 3 3 13 3 0 10 9 10 9 0 13 13 10 11 1 10 9 13 15 10 9 1 0 9 13 10 9 3 1 0 13 13 3 3
35 1 10 9 13 9 0 13 13 0 16 3 10 9 13 1 9 13 3 1 10 9 13 1 10 0 9 7 3 13 10 9 1 10 0 13
11 15 3 3 10 3 13 3 10 0 9 13
5 7 0 3 3 13
6 3 3 3 13 13 15
40 11 3 16 13 1 10 9 13 10 11 1 10 11 13 10 3 11 13 10 9 0 10 0 1 11 9 10 1 0 9 3 3 13 3 13 13 10 0 10 9
14 11 3 13 10 15 9 7 13 10 3 13 15 13 11
16 16 3 13 13 10 9 13 9 1 10 9 13 15 1 11 13
5 9 3 3 3 13
17 11 3 16 13 7 13 11 3 1 10 0 9 13 1 10 0 15
7 7 10 3 9 0 3 13
83 11 3 13 1 10 9 10 15 9 13 3 15 10 13 9 0 0 3 10 11 0 13 16 10 0 3 13 13 10 11 13 1 10 11 1 9 13 13 3 0 1 10 9 13 3 3 1 11 13 11 9 0 3 3 1 0 13 3 3 0 3 3 1 0 15 13 9 13 3 10 9 0 10 0 11 13 3 3 0 13 1 9 0
20 13 7 3 0 7 10 15 13 9 13 10 9 13 1 10 9 13 1 10 9
26 10 3 13 7 13 9 9 15 13 15 0 15 13 13 0 13 16 3 3 13 3 3 11 13 1 11
8 0 13 11 10 9 15 9 13
11 13 3 15 10 9 13 10 9 13 13 13
10 13 3 0 11 3 3 13 13 9 13
8 3 3 13 0 1 10 9 9
29 9 3 0 13 9 0 0 13 11 1 10 9 13 3 0 13 10 0 13 9 13 9 9 9 3 0 7 7 9
19 9 3 3 0 13 11 3 13 15 3 13 15 13 1 11 7 7 0 11
9 16 3 15 0 13 3 13 1 9
11 13 3 10 9 1 10 11 15 9 11 13
16 13 3 0 10 9 9 15 1 10 11 7 0 7 0 10 0
16 10 3 9 15 13 1 9 9 7 13 0 7 15 13 13 0
66 1 10 9 3 13 0 15 1 10 9 13 10 0 13 0 7 7 0 1 3 15 9 13 7 15 7 11 13 1 10 0 13 3 11 15 1 9 0 9 11 13 13 1 9 1 11 9 3 10 11 16 13 10 9 1 9 13 13 10 9 13 11 13 9 9 0
25 15 10 9 10 15 13 0 7 7 0 9 0 15 13 7 13 10 9 9 1 15 13 0 9 13
8 10 3 9 13 10 0 9 13
26 16 3 10 15 13 13 10 3 0 9 3 13 13 15 10 3 13 11 3 0 3 13 7 16 13 13
3 0 3 13
9 10 3 9 13 1 10 9 0 1
15 9 9 13 7 3 13 7 10 9 15 13 7 10 9 13
21 15 3 3 0 1 13 16 10 11 0 13 10 0 15 3 15 3 13 13 10 9
26 16 3 3 13 1 10 9 3 3 13 3 10 9 10 9 7 13 15 3 13 13 7 10 11 10 9
22 3 3 10 3 9 10 3 0 13 7 16 13 10 13 13 1 10 9 0 10 9 13
5 15 3 3 13 9
19 11 3 13 15 9 1 0 13 10 9 13 1 10 9 0 9 1 10 9
22 10 3 3 0 13 1 0 9 13 13 1 11 0 3 13 10 0 13 13 3 13 11
13 1 7 3 3 10 0 13 9 7 3 3 1 11
20 10 3 3 0 10 9 1 0 0 10 9 13 9 13 1 0 1 9 13 11
12 10 3 11 0 13 10 0 9 13 13 10 0
25 13 3 3 10 1 9 10 1 9 0 10 7 1 10 9 9 7 10 0 9 7 10 0 10 9
23 13 3 0 10 15 13 3 13 1 9 13 16 12 0 13 15 3 3 13 0 13 10 9
3 13 0 13
5 9 3 0 13 13
20 13 3 15 7 13 0 13 1 9 12 12 0 3 11 7 7 11 0 3 11
5 13 3 0 9 13
12 10 3 3 12 10 0 3 13 13 1 10 11
22 10 3 10 0 11 13 10 0 0 7 13 10 9 1 10 15 9 1 10 9 13 15
6 9 3 0 13 13 0
29 3 3 3 15 0 13 13 13 15 3 16 15 0 13 15 3 15 3 13 13 10 3 15 13 7 13 10 0 0
32 0 3 3 1 0 10 9 13 10 9 0 0 13 13 9 7 7 9 3 0 13 9 0 15 7 10 9 15 13 16 11 13
15 0 3 10 0 0 13 9 3 3 13 1 0 1 0 13
24 10 3 12 13 10 13 10 12 11 13 13 1 11 10 15 9 13 3 15 1 10 11 13 15
14 0 3 10 9 13 9 13 10 0 9 13 11 13 13
9 15 3 3 16 13 10 9 13 13
21 7 15 3 13 7 9 13 0 13 0 9 16 13 10 9 10 9 7 13 11 13
8 3 3 0 3 9 13 0 13
21 16 0 13 9 13 11 11 10 9 10 15 13 9 13 10 0 13 10 9 9 13
9 3 3 13 0 1 0 16 13 3
9 0 7 3 13 3 10 9 7 0
28 3 3 11 10 0 9 11 0 3 13 10 9 15 15 10 9 13 9 13 16 13 10 9 10 9 13 11 0
23 10 3 11 1 10 0 9 13 3 13 0 15 9 10 9 13 0 3 13 0 7 7 0
8 13 3 1 10 11 13 10 9
29 10 3 3 11 0 10 0 13 10 0 10 15 9 1 0 10 9 13 1 9 3 13 7 13 13 7 1 9 13
13 13 3 0 3 3 11 7 13 7 15 10 9 13
6 1 0 3 11 0 13
12 1 10 3 13 9 10 11 10 15 1 15 13
12 15 3 13 7 3 3 1 11 1 15 13 13
6 10 3 11 15 13 0
16 9 9 0 9 0 0 11 3 13 0 9 1 9 13 9 13
7 10 3 15 0 0 3 13
13 13 3 10 9 13 3 10 15 9 13 11 3 13
10 11 3 3 13 13 1 10 13 9 13
6 7 15 15 13 13 13
2 13 3
5 6 9 3 13 11
6 0 3 3 0 0 13
10 1 3 0 3 13 10 15 9 10 9
8 13 3 15 10 9 13 1 11
61 15 3 13 9 0 13 1 15 10 11 7 1 9 13 7 3 12 9 1 15 9 1 9 13 7 3 9 0 13 9 15 3 7 3 9 13 13 7 3 13 10 11 13 0 0 1 13 1 10 9 13 13 16 15 15 9 13 10 3 13 13
5 15 3 3 13 0
28 10 3 11 13 1 10 9 13 3 1 0 13 0 10 10 11 16 15 13 1 9 13 10 15 13 10 13 0
17 7 10 11 13 13 10 9 13 10 11 15 0 13 7 15 13 13
7 11 3 3 3 9 13 13
5 3 3 16 13 13
9 16 3 15 0 13 3 13 10 13
55 13 3 15 7 9 13 13 3 16 13 9 10 11 13 0 7 13 15 10 15 9 13 15 3 13 16 7 15 15 13 3 3 0 13 15 15 3 1 15 13 3 3 1 0 10 0 7 3 10 1 15 0 0 13 13
5 10 3 11 0 13
8 10 3 9 3 13 13 10 9
59 7 10 11 13 10 9 15 11 13 13 7 7 13 16 3 0 9 13 0 9 13 15 9 3 0 13 9 13 1 7 0 13 10 9 7 13 16 15 13 10 1 9 3 13 13 13 10 0 10 13 9 7 13 11 7 7 10 1 11
40 3 13 1 9 11 13 10 11 9 16 13 15 3 9 13 10 9 13 3 3 13 13 10 11 13 16 15 15 13 1 15 13 13 7 13 15 1 10 13 0
6 15 3 13 13 10 9
21 3 3 13 10 11 16 13 10 11 7 0 7 9 0 13 15 1 10 9 13 0
15 11 15 15 9 13 1 9 10 15 13 0 1 9 15 13
3 15 3 13
13 6 9 15 0 13 10 15 3 9 10 15 3 9
10 0 3 0 13 10 9 9 13 15 13
10 15 3 3 0 13 15 9 1 9 13
8 7 0 9 3 0 13 3 13
25 11 3 15 13 13 7 1 15 7 3 1 0 9 13 13 7 13 7 15 7 10 1 0 13 15
6 15 3 9 13 0 13
14 3 3 13 7 7 13 10 9 10 10 9 9 13 13
15 6 9 15 13 1 15 15 13 13 7 13 1 10 13 13
9 11 3 15 13 13 13 15 15 13
5 15 3 15 13 13
9 0 10 0 9 15 0 0 9 13
3 11 3 13
9 7 9 10 15 7 9 10 15 13
6 15 3 15 3 0 13
7 7 13 7 7 13 10 15
7 11 3 0 13 15 11 13
13 13 3 10 15 13 11 15 15 15 13 1 10 13
3 15 3 13
13 16 15 9 13 9 15 13 16 15 13 0 13 15
25 16 3 15 0 13 13 7 13 9 0 0 15 1 15 0 13 15 3 15 0 13 0 13 15 13
10 3 3 13 3 16 15 13 15 15 13
23 13 10 9 1 15 10 9 9 15 13 1 10 13 10 9 13 16 15 3 13 13 10 11
18 7 15 7 15 3 13 9 13 10 9 7 0 13 13 15 0 0 13
10 0 13 10 11 13 16 15 13 3 13
15 13 3 0 7 13 10 9 15 11 13 13 13 1 11 0
17 11 13 15 9 9 0 9 7 9 13 13 9 15 13 15 13 3
3 15 3 13
25 11 3 15 13 15 10 15 9 7 10 9 10 9 7 3 10 9 7 16 13 10 9 13 1 9
12 13 3 0 13 3 13 13 15 10 9 0 13
4 11 3 13 13
13 7 0 13 1 15 11 7 15 15 15 3 3 13
46 16 3 0 13 10 11 13 10 9 1 11 13 13 10 9 1 10 9 10 9 13 16 3 15 13 10 9 13 11 13 1 9 3 13 10 11 9 1 15 15 9 0 13 13 10 9
11 0 7 13 7 16 0 9 13 10 0 9
13 13 3 10 9 7 13 10 13 10 11 13 13 0
24 11 3 0 9 9 13 15 13 9 9 9 0 13 13 10 9 7 13 10 0 9 15 15 13
9 15 3 13 0 13 7 7 13 15
19 12 3 9 13 10 11 9 7 0 13 11 3 0 10 9 0 13 10 13
6 0 3 0 13 15 13
10 1 3 10 9 10 13 3 3 11 13
12 13 3 15 11 16 13 1 9 0 9 15 13
18 15 3 1 0 13 3 13 13 13 13 15 10 15 7 10 11 13 9
9 15 7 10 0 13 13 11 1 9
3 3 0 13
11 1 3 12 3 0 13 9 0 9 3 0
29 15 3 3 13 9 7 11 9 10 9 9 15 3 9 7 13 7 13 1 0 7 3 13 10 0 9 10 15 13
7 0 3 10 11 13 10 9
8 15 3 13 1 11 7 13 11
12 15 3 13 13 15 13 10 9 7 3 10 9
14 11 3 13 0 9 1 10 11 0 7 3 10 13 0
36 1 3 3 11 10 9 9 0 15 13 10 11 10 0 1 3 11 10 7 9 10 0 7 10 9 10 0 1 3 0 10 1 11 9 0 0
8 0 3 3 3 1 15 13 13
19 10 3 1 11 10 0 9 11 3 15 13 0 7 9 7 0 10 1 11
19 10 3 3 1 7 11 7 1 10 11 13 0 7 13 7 10 0 9 9
22 10 3 0 9 1 9 13 9 0 15 15 16 3 13 9 13 13 11 13 10 9 9
12 10 3 11 13 11 3 9 11 3 9 3 0
18 16 3 13 10 9 13 10 9 10 11 10 9 10 13 1 9 13 13
15 10 3 9 15 3 0 13 3 9 10 13 13 1 15 13
6 7 1 3 9 0 13
22 9 3 9 10 11 1 9 3 3 13 15 3 3 0 9 1 10 1 10 11 13 9
20 13 3 11 10 11 9 9 15 10 9 3 13 9 0 10 3 15 9 9 9
13 13 3 15 10 0 9 7 10 9 7 10 13 9
29 9 3 12 13 3 3 1 15 13 1 10 9 3 7 15 9 13 15 0 13 7 13 13 10 10 9 9 13 0
4 13 3 0 15
20 10 3 3 9 10 9 13 9 12 7 12 9 10 3 9 13 9 12 7 12
11 9 3 13 10 9 0 15 13 9 0 13
4 13 3 0 11
5 0 3 3 0 13
5 0 3 3 9 13
17 13 3 0 9 3 10 9 10 3 15 7 7 9 13 15 9 13
19 1 11 10 11 9 9 0 1 10 11 15 13 7 10 9 3 3 13 13
7 3 3 16 3 13 9 13
5 15 3 15 13 15
22 13 3 3 3 7 10 9 7 10 9 7 10 9 7 10 0 15 9 10 9 1 9
8 0 3 3 10 9 3 13 9
7 13 3 3 1 10 9 13
8 0 9 13 1 9 12 13 12
15 13 3 15 10 0 13 1 10 9 13 1 11 7 13 9
34 1 15 13 10 15 15 15 13 0 9 13 1 9 7 7 9 9 16 15 9 0 13 13 1 9 3 15 13 9 7 13 10 1 0
13 1 3 9 13 15 1 10 9 10 9 15 15 13
7 1 0 10 9 13 13 9
6 9 3 3 1 9 13
25 13 3 3 10 3 15 10 9 10 7 11 15 13 10 11 9 13 7 10 9 15 9 13 10 11
29 3 3 9 0 13 10 3 13 13 10 1 11 7 10 13 13 9 1 0 13 13 1 11 3 0 0 9 9 13
12 13 3 0 15 1 10 9 3 3 1 9 13
10 9 1 10 9 13 0 15 9 13 11
4 9 3 13 11
7 0 10 11 13 9 13 0
20 13 10 9 1 9 1 10 15 13 3 0 0 3 3 15 7 0 9 13 13
19 7 0 3 13 9 0 1 15 10 0 13 13 16 10 0 10 0 0 13
15 10 3 1 10 0 9 9 13 15 10 9 9 15 15 13
11 15 3 3 15 13 9 0 7 7 0 13
5 9 3 15 15 13
34 0 3 3 13 10 13 15 13 10 9 13 1 10 13 13 10 11 1 15 15 13 7 13 3 13 3 3 0 13 13 7 13 13 3
12 3 3 15 13 10 15 13 10 3 1 9 13
28 13 3 9 7 9 3 0 3 1 10 9 3 0 13 13 10 9 1 10 15 7 13 15 9 13 1 10 13
10 3 3 15 13 3 13 10 10 11 9
12 3 3 3 9 10 13 13 0 13 13 10 9
5 13 13 15 0 9
16 7 3 10 7 9 13 7 0 1 9 13 3 1 9 0 13
15 15 3 13 15 9 7 15 0 10 9 13 7 13 15 9
5 13 3 0 10 9
22 13 7 3 15 9 0 7 7 0 3 15 13 10 9 7 9 15 13 1 15 9 13
19 15 3 16 13 10 9 10 9 13 12 9 13 7 0 13 10 15 0 13
21 13 3 3 0 10 9 13 9 0 7 7 0 0 15 3 11 13 0 0 3 13
17 13 3 3 0 10 9 16 10 0 10 0 9 10 9 0 13 0
13 0 3 3 15 7 10 9 13 9 13 16 0 13
16 9 3 13 10 0 12 1 3 10 0 10 9 13 7 10 9
23 10 3 3 0 9 10 9 13 0 10 3 0 0 0 3 9 0 0 3 0 0 3 0
9 3 10 12 9 10 9 13 13 9
14 12 3 10 0 13 15 3 13 15 3 13 13 10 9
13 0 3 3 10 11 15 7 13 7 1 10 15 9
9 10 3 0 9 1 13 10 9 13
40 13 3 15 9 0 11 0 13 10 13 3 13 1 9 15 1 9 3 15 13 13 7 9 1 15 1 7 0 3 13 7 7 0 13 3 0 13 0 3 0
14 16 3 0 13 7 13 15 10 9 13 10 0 13 0
15 7 10 7 9 13 3 1 0 13 7 0 13 10 13 13
5 0 3 0 13 15
25 16 15 13 13 0 16 13 1 9 0 9 13 7 15 9 7 7 0 13 1 15 10 9 15 13
11 11 3 3 10 0 9 13 0 7 0 13
11 13 3 9 0 9 9 9 9 9 0 9
6 9 3 3 9 13 0
21 13 3 3 13 0 9 13 7 13 1 10 9 0 7 0 13 7 0 9 0 13
67 3 3 13 12 0 9 7 0 0 13 10 11 1 0 1 0 13 9 16 15 13 1 10 0 7 0 0 15 11 13 7 13 0 15 3 3 13 13 3 9 3 13 3 3 15 3 13 1 0 3 13 10 11 0 7 13 13 12 7 12 9 7 10 9 15 10 0
10 11 3 13 13 11 10 11 10 11 9
8 1 15 3 3 13 15 3 13
23 0 10 10 9 13 13 16 9 10 9 13 15 13 7 10 10 11 9 1 11 15 13 15
21 13 3 10 1 15 13 15 13 1 10 11 13 7 10 9 7 10 9 0 13 13
14 7 15 16 13 13 10 0 13 10 11 13 9 9 0
11 15 13 3 1 10 11 0 13 1 10 11
10 0 3 13 13 3 1 10 0 9 13
17 13 3 1 10 9 10 0 1 11 9 7 1 9 12 9 0 9
19 1 3 10 11 3 0 13 1 10 0 7 12 10 1 0 9 15 13 9
20 3 3 10 3 9 3 13 7 10 3 9 0 0 13 1 0 13 10 0 9
14 3 10 3 9 13 10 9 7 13 10 9 10 9 13
7 10 3 9 10 11 15 13
21 7 16 13 1 10 11 0 11 15 11 9 13 9 7 7 9 13 10 3 3 13
26 15 3 16 13 3 13 10 11 1 11 9 10 0 9 13 0 0 15 15 13 13 10 0 11 10 9
16 13 3 0 10 9 3 15 13 13 15 0 9 15 0 10 9
25 3 3 10 1 11 9 3 13 3 0 0 13 7 10 1 11 9 13 10 13 1 0 10 11 13
20 10 3 10 9 13 10 9 10 1 11 7 10 0 3 9 13 10 9 0 9
23 1 3 3 12 7 12 9 13 10 11 10 9 7 10 15 15 1 7 9 7 9 0 13
10 3 3 3 9 13 1 0 15 0 13
46 7 0 3 10 0 11 7 7 9 13 7 13 13 7 3 13 10 9 9 7 13 15 3 3 0 7 10 7 11 13 3 3 13 1 0 9 13 7 10 0 0 13 1 10 0 9
13 1 3 0 11 3 13 12 9 1 15 9 13 13
7 13 3 11 11 9 10 9
8 7 15 13 9 15 9 13 11
20 15 13 11 1 10 9 13 0 16 13 3 10 15 9 13 3 3 10 11 15
14 13 3 10 9 10 9 10 9 13 1 15 0 0 13
24 15 3 9 13 15 9 13 11 15 13 9 3 13 0 9 3 0 0 1 13 15 0 9 0
18 13 3 15 1 10 9 10 9 0 13 9 10 3 9 13 10 11 15
15 13 3 0 7 13 10 9 13 1 10 9 10 9 9 13
9 13 3 13 13 10 13 1 15 13
20 1 3 15 10 9 10 10 9 9 13 16 13 10 10 9 15 9 13 1 0
26 0 3 3 13 10 11 16 13 10 11 13 11 9 0 7 0 7 9 7 15 9 10 15 13 15 0
20 11 9 15 3 15 13 3 13 7 15 7 13 7 15 13 1 0 15 0 13
5 13 15 11 13 9
3 15 3 13
10 6 9 3 3 3 13 9 0 0 15
11 13 3 1 15 3 1 10 3 9 15 13
14 7 16 15 0 0 3 13 13 3 10 3 15 13 3
18 0 13 10 11 16 15 13 10 9 13 10 1 9 13 13 1 10 9
11 13 3 13 10 15 9 10 15 11 13 9
5 15 3 1 15 13
8 3 3 15 15 1 9 13 13
4 3 3 13 11
21 3 16 13 7 7 13 3 3 3 13 3 15 15 13 10 9 7 1 9 0 13
24 0 3 1 3 13 15 7 16 0 15 0 13 10 9 7 16 11 3 13 9 7 9 0 9
29 16 3 13 0 13 1 10 9 0 13 10 9 15 3 10 9 13 1 15 0 15 3 13 10 3 15 9 10 0
11 7 10 3 0 1 15 13 0 13 10 9
12 13 3 10 15 11 15 9 13 7 3 10 15
20 0 13 7 3 9 13 1 10 9 15 11 15 13 9 7 0 13 7 9 0
4 15 9 13 11
6 10 3 9 13 8 9
28 10 3 9 13 10 9 3 10 9 10 9 13 0 3 10 9 1 11 7 9 10 11 7 1 10 9 10 0
25 3 3 3 10 0 9 1 9 0 13 3 7 0 7 7 9 0 10 3 0 0 9 13 15 0
12 16 3 10 9 9 0 13 13 13 10 11 0
17 13 15 11 10 9 0 13 13 1 10 0 10 9 16 3 3 13
18 7 0 15 13 13 16 3 13 15 7 15 9 13 9 10 0 15 13
5 13 3 13 13 15
21 15 3 3 3 0 10 9 9 13 15 9 3 3 1 9 13 13 10 9 1 9
19 16 3 13 13 15 1 0 13 10 9 13 0 15 15 15 3 3 11 13
3 15 3 13
20 6 9 13 7 1 9 13 7 13 0 7 13 13 7 3 13 1 9 10 15
6 9 3 15 11 9 13
5 15 3 13 13 3
17 3 3 0 13 13 9 13 13 7 7 13 13 9 7 7 9 0
9 7 15 13 13 13 10 15 9 13
8 3 3 3 3 13 3 3 13
36 7 3 3 1 9 13 10 15 9 9 15 15 13 1 9 13 10 9 16 3 11 7 13 9 10 11 9 7 11 10 11 7 15 11 13 13
4 3 7 0 13
9 16 3 0 13 10 9 3 13 13
23 15 3 16 13 10 9 0 7 7 0 13 13 7 13 10 9 10 9 13 15 9 13 15
10 15 3 3 13 0 3 13 3 15 13
12 16 3 3 13 3 10 9 0 13 10 9 0
18 16 3 3 13 15 13 3 13 15 3 3 13 16 3 15 9 13 13
4 13 3 3 15
4 0 3 13 13
11 10 3 10 11 9 9 3 1 15 13 13
13 7 3 7 15 13 13 10 9 7 15 3 13 13
14 10 7 3 13 0 9 13 7 10 13 3 13 10 9
11 15 3 13 13 9 0 3 13 10 15 9
15 10 3 15 13 0 13 13 1 10 9 1 15 13 10 0
15 13 3 10 9 15 10 0 9 13 1 10 0 10 9 13
19 16 3 0 9 10 9 13 13 13 1 9 10 9 10 15 9 9 3 13
19 13 3 10 11 10 15 9 10 0 13 7 1 0 7 13 10 9 10 9
4 7 15 3 13
20 10 3 0 0 11 13 13 13 10 9 10 9 9 15 3 15 7 3 11 13
12 13 1 10 9 0 1 15 13 3 10 9 0
7 13 3 1 0 9 1 9
15 7 10 9 13 13 15 9 13 0 3 10 10 9 9 9
20 15 3 15 13 15 3 9 13 15 3 9 13 10 3 3 15 15 9 9 13
12 10 3 15 10 9 13 13 9 3 0 9 13
6 13 15 10 15 9 13
12 13 3 10 9 10 11 10 9 3 3 13 13
30 13 3 1 9 1 10 9 13 15 1 11 13 13 3 3 11 3 3 3 13 0 10 9 7 1 10 9 10 11 9
36 10 3 11 9 3 13 13 1 10 11 7 3 13 10 9 0 9 13 13 13 6 9 1 10 15 9 9 3 9 3 13 13 10 9 10 9
20 13 3 7 13 11 13 13 10 9 9 10 11 1 13 10 7 9 7 10 9
11 16 3 13 0 13 1 10 11 10 11 13
18 15 3 13 0 0 13 9 13 10 0 9 13 0 1 15 9 0 13
4 15 3 13 3
16 10 3 15 1 10 9 9 15 3 0 13 13 15 0 13 9
8 10 3 3 0 9 10 13 13
13 0 3 13 7 7 9 13 15 16 15 13 10 9
12 16 3 3 0 1 0 15 0 13 0 15 13
36 0 13 10 9 10 11 13 9 15 7 15 10 7 9 10 9 13 13 1 15 7 10 9 0 13 10 7 9 10 9 10 9 10 9 13 13
7 13 3 0 1 9 0 13
16 3 3 3 3 13 13 13 13 10 11 16 10 9 0 13 13
13 11 15 0 13 16 15 7 10 9 10 15 15 13
21 16 3 13 10 9 0 3 0 15 13 10 11 3 13 10 9 7 15 13 10 13
15 15 3 1 15 7 13 13 7 10 13 15 13 3 1 15
21 11 3 15 3 3 13 13 13 1 9 0 13 3 7 13 0 13 10 9 13 15
12 15 3 13 1 10 9 3 3 13 10 13 9
19 13 3 1 9 13 10 9 13 7 13 1 9 3 3 9 15 13 13 15
13 11 3 10 3 9 10 9 13 9 3 3 0 13
10 11 3 3 3 13 13 15 10 9 13
10 16 3 15 13 10 11 13 15 10 11
21 10 3 11 16 13 10 9 3 13 3 13 1 0 9 16 3 13 13 7 13 0
29 6 9 16 13 10 9 13 13 3 15 7 13 1 9 7 15 1 15 13 0 7 9 10 15 7 0 15 13 9
3 13 3 3
15 13 10 9 0 13 10 9 13 15 3 13 10 13 13 15
6 7 13 0 3 3 13
4 15 3 13 3
25 13 3 0 1 0 13 13 15 1 0 9 7 13 13 16 15 13 13 0 0 16 3 0 0 13
21 16 3 13 0 10 13 13 10 9 13 10 9 10 0 7 13 1 0 7 13 15
25 11 3 13 15 15 13 9 1 10 13 0 3 3 3 13 0 1 10 9 10 9 3 13 10 11
17 3 3 16 15 13 13 13 16 13 7 10 9 7 10 13 13 3
21 10 7 3 13 13 13 1 10 9 0 13 3 7 9 10 15 13 3 1 0 13
17 3 3 10 9 3 13 0 3 10 15 9 13 1 10 9 10 0
17 0 3 9 3 10 9 13 13 15 9 9 0 13 13 15 1 9
29 11 3 16 13 0 13 7 0 13 16 7 10 9 15 1 9 13 7 16 1 9 0 1 9 13 13 1 10 9
31 13 3 10 0 13 3 15 9 12 0 9 12 7 12 3 3 13 0 13 13 7 13 1 11 7 13 15 15 3 0 13
22 11 3 16 15 13 10 11 9 13 15 7 1 9 13 15 3 13 15 3 13 10 9
44 16 3 10 9 13 10 9 13 10 7 0 9 7 10 11 10 3 0 7 0 11 13 9 0 9 9 11 3 10 9 10 15 3 9 7 7 0 9 7 7 9 10 0 15
7 0 3 3 13 1 9 13
17 16 3 10 11 13 3 13 10 9 11 13 15 16 13 15 10 9
20 13 3 11 7 3 13 13 15 13 10 9 10 9 13 7 10 9 7 10 9
11 11 3 13 13 13 7 7 13 15 13 15
11 13 3 10 11 7 13 13 10 9 10 9
11 13 3 15 10 11 16 13 15 9 9 13
13 15 3 7 13 13 7 0 13 15 15 3 9 13
10 3 3 13 3 15 13 13 13 10 15
6 11 3 11 9 0 13
15 11 3 1 13 13 10 0 10 9 15 10 9 15 3 13
10 13 3 13 10 11 3 13 15 10 9
18 15 3 1 10 0 13 13 16 13 13 10 9 16 13 7 3 13 0
18 13 7 10 9 7 13 7 15 1 9 13 10 1 10 9 9 13 9
11 15 3 15 15 3 10 0 9 9 13 13
13 7 3 9 7 9 7 9 7 10 0 15 13 13
3 13 10 9
20 16 3 13 7 7 13 10 9 3 1 9 15 13 7 0 1 7 9 13 0
6 3 3 3 10 0 13
19 1 0 3 7 10 9 15 15 13 7 10 3 10 9 13 3 1 0 13
25 3 0 6 9 3 0 9 13 9 13 10 9 13 7 10 9 7 15 10 9 0 13 0 3 15
18 3 3 3 3 13 15 3 13 15 13 0 13 9 7 10 15 7 15
5 13 1 0 10 9
12 6 9 3 0 15 1 0 13 13 9 10 15
16 15 3 13 9 13 9 7 13 10 9 7 9 1 15 0 13
11 3 3 3 15 15 7 10 15 9 13 13
10 7 3 16 0 15 13 15 3 15 13
13 10 3 9 0 1 9 13 1 9 7 7 10 13
13 13 0 10 11 13 7 7 13 10 11 13 15 0
11 6 9 15 3 15 1 9 9 3 0 13
5 10 15 3 9 13
6 3 3 13 13 1 9
18 13 3 3 9 7 7 9 13 3 1 11 7 10 9 7 10 9 15
7 0 13 10 11 13 10 11
21 15 3 15 13 13 1 15 3 3 13 7 13 0 1 9 3 13 15 10 15 9
9 13 3 3 16 9 10 11 13 9
11 1 3 10 3 9 10 15 9 10 9 13
8 13 3 13 1 10 10 9 9
6 13 7 0 13 1 15
10 13 7 15 1 10 9 10 15 10 11
6 3 3 10 9 0 13
11 1 15 3 13 9 3 13 9 13 1 11
13 11 3 13 13 13 9 10 9 10 11 15 15 13
7 1 3 3 0 0 15 13
24 13 10 11 0 1 10 9 13 12 0 10 11 10 0 9 13 16 13 11 13 11 13 10 9
28 13 3 15 0 7 13 0 3 3 10 11 13 1 9 13 11 13 10 15 9 3 3 3 13 3 10 9 13
4 15 3 13 0
20 9 13 7 13 0 10 9 7 15 13 3 3 13 3 13 9 13 15 15 13
9 13 3 1 15 10 9 13 13 13
5 10 3 9 13 0
7 6 9 11 15 3 9 13
8 3 3 3 3 1 0 9 13
7 15 3 11 10 15 9 13
7 1 3 3 10 0 9 13
8 10 3 1 9 7 7 15 13
27 15 15 3 3 13 15 13 15 7 0 1 3 13 7 15 15 1 11 13 16 15 3 13 7 13 10 9
7 9 3 13 13 13 1 9
22 7 16 7 15 1 11 13 9 1 15 13 15 15 15 13 16 7 10 15 0 0 9
13 0 3 0 13 1 0 7 13 1 15 11 13 13
13 3 3 0 10 3 3 13 13 0 7 13 1 9
11 13 0 10 11 13 15 9 0 9 13 13
6 13 3 13 0 0 13
3 13 3 0
9 13 1 9 15 13 9 10 9 13
4 11 3 0 13
5 13 3 9 0 9
12 7 15 3 15 10 11 13 7 13 13 1 9
13 13 3 0 1 15 10 0 15 13 9 9 0 0
16 0 9 13 0 1 15 3 9 13 9 3 10 9 10 9 13
8 0 3 9 13 0 0 0 0
13 0 3 15 9 13 10 3 15 9 9 9 9 0
15 13 3 10 9 10 13 9 0 15 13 1 10 0 13 13
10 13 3 10 0 10 9 13 1 9 13
20 16 3 1 9 13 13 15 10 11 3 15 10 0 13 7 10 13 15 13 0
8 15 3 13 0 13 15 10 0
15 10 3 3 0 9 15 15 0 13 10 3 3 13 15 0
12 13 3 0 10 9 10 11 13 10 15 9 13
5 9 9 3 15 13
6 9 3 13 9 0 13
32 9 3 7 9 7 9 3 1 9 13 13 7 7 10 13 9 13 3 3 15 13 16 3 0 13 10 9 3 3 10 9 13
14 13 3 9 7 7 9 7 9 7 9 7 9 7 9
6 0 3 3 13 0 3
12 13 3 3 10 11 13 1 7 0 13 7 0
12 13 3 0 10 11 11 0 3 11 9 3 11
10 9 3 10 9 1 10 13 9 0 13
9 3 9 13 3 9 3 9 3 9
20 15 3 16 15 13 13 1 9 0 13 10 9 13 10 9 13 10 9 9 3
12 15 3 3 10 13 0 0 3 15 13 13 0
9 1 3 3 10 0 9 3 15 13
25 16 3 13 1 9 10 9 13 10 9 13 9 3 0 3 3 10 9 1 0 13 3 15 10 9
15 13 3 15 9 9 13 13 9 15 3 0 13 13 10 9
10 1 3 3 9 3 15 9 13 9 13
10 9 3 0 3 0 13 13 3 0 13
9 1 0 3 0 9 10 0 13 13
26 1 15 10 0 15 9 7 9 7 9 7 9 13 0 0 1 9 10 3 0 15 10 9 10 9 13
10 9 3 0 13 9 3 0 7 3 0
8 16 3 15 13 13 3 3 13
13 9 3 3 13 7 15 3 13 13 3 13 0 0
5 0 3 3 3 13
18 15 3 3 13 15 13 0 10 0 13 13 10 9 1 15 3 13 13
8 7 16 3 13 3 13 13 15
5 16 3 3 13 13
7 15 3 3 13 13 13 13
15 13 3 15 1 10 9 0 3 15 13 16 0 13 10 13
10 16 3 13 10 0 0 0 10 9 13
11 16 3 0 13 10 0 0 13 13 10 0
6 3 3 1 9 13 13
33 3 3 10 15 3 13 1 9 13 13 15 13 9 0 10 15 0 10 3 0 1 9 10 9 13 10 3 3 13 1 15 0 13
28 1 3 9 13 10 3 13 10 9 15 0 3 9 7 10 3 13 15 0 3 3 10 0 15 3 3 10 13
9 1 10 0 3 9 3 10 9 13
9 13 3 3 10 9 13 7 7 13
7 0 3 0 9 13 9 3
14 7 9 7 0 13 13 7 3 7 1 9 13 9 13
6 0 3 3 0 9 13
14 9 3 0 13 1 10 13 13 0 15 3 0 13 9
11 10 3 10 0 13 9 13 9 1 15 9
6 10 0 3 13 0 13
16 13 3 10 9 1 0 13 1 0 12 0 13 7 13 7 13
17 16 3 3 0 13 3 13 1 9 10 9 7 1 10 9 9 13
15 0 3 1 0 3 13 16 16 13 13 15 9 10 9 13
26 13 3 15 3 13 10 15 9 7 9 7 15 3 0 13 15 9 13 13 0 13 7 0 13 7 0
15 3 3 3 13 9 13 10 3 3 9 1 10 15 9 13
10 15 3 15 13 3 13 0 3 13 13
11 0 3 0 10 13 13 0 3 10 13 9
5 0 3 3 15 1
11 3 3 9 13 13 10 13 3 15 9 13
19 15 3 3 10 9 9 7 9 13 1 9 0 3 13 7 13 10 15 9
10 13 3 15 1 10 9 13 15 0 13
8 3 10 0 9 10 0 9 13
18 1 9 3 7 13 7 13 3 9 13 7 0 15 13 7 13 9 3
15 7 0 15 15 3 13 13 15 9 3 0 13 15 3 3
24 10 9 15 13 0 10 9 7 10 9 13 15 1 10 0 9 15 9 3 8 13 9 3 9
18 1 0 13 13 13 10 9 10 9 3 15 3 15 3 3 7 15 3
8 0 3 3 13 1 15 13 13
26 0 3 3 13 13 7 3 3 1 10 13 16 3 0 13 9 9 10 9 16 3 1 9 7 9 13
7 9 3 3 3 13 0 13
13 9 3 13 0 10 7 0 9 7 10 1 11 9
11 15 3 3 13 0 15 13 3 3 15 13
28 10 3 3 9 9 15 1 9 7 9 13 7 9 0 0 13 13 3 9 7 7 9 7 10 15 9 7 9
11 7 1 3 10 9 0 13 3 3 9 13
6 13 3 1 10 0 9
27 9 3 7 9 16 10 9 3 13 1 9 13 9 1 11 1 11 13 1 10 0 13 15 3 11 13 0
23 15 3 13 15 15 13 13 15 9 9 13 9 13 9 1 10 9 13 13 15 13 1 9
8 15 3 3 9 13 13 15 0
12 1 0 3 0 9 11 13 1 15 3 10 9
14 10 3 0 9 13 0 9 13 9 1 11 13 9 13
26 10 3 9 0 15 3 10 11 13 10 3 9 7 10 9 1 10 0 13 13 9 15 9 15 15 13
41 7 3 10 1 15 9 10 0 13 10 11 7 10 3 7 10 1 10 9 7 10 1 10 9 0 3 1 10 0 7 7 0 13 0 3 1 10 0 7 7 0
11 9 3 3 10 0 0 13 7 9 12 9
14 11 3 15 0 13 9 1 9 3 3 11 7 7 11
11 0 3 10 9 10 0 13 13 1 9 15
3 15 3 13
5 0 9 9 12 13
22 0 3 3 10 9 10 0 3 13 1 9 10 9 9 13 10 3 15 9 13 0 15
12 7 3 9 13 3 9 0 7 0 10 9 9
11 13 3 1 10 0 9 0 1 15 3 15
26 10 3 3 15 9 7 10 0 13 10 9 3 13 9 13 7 3 3 13 15 10 0 15 13 10 9
39 3 3 10 1 10 9 3 9 9 0 3 9 10 15 0 13 13 3 0 13 10 0 9 1 10 0 9 7 3 15 0 10 1 10 9 13 13 10 9
29 1 3 10 9 10 0 11 13 10 3 9 0 10 13 7 0 13 10 13 1 10 9 3 13 7 3 13 10 9
11 9 3 9 15 9 13 11 13 10 9 13
25 1 0 10 9 10 12 9 11 7 11 7 7 11 7 11 7 7 11 13 10 9 10 0 9 11
8 0 3 3 0 0 10 9 13
11 0 12 9 3 0 13 7 3 3 9 13
9 0 3 1 3 10 9 12 9 13
25 9 3 0 15 13 7 0 7 9 7 9 0 7 0 7 9 9 7 9 0 0 7 9 0 13
29 15 3 15 1 10 9 10 0 13 7 13 0 13 9 0 3 3 9 13 1 10 9 7 9 13 15 13 10 9
6 0 3 13 13 1 11
24 9 3 13 15 3 15 0 1 11 10 11 13 15 3 9 0 1 11 10 11 15 3 3 0
12 13 3 15 9 15 1 11 13 7 11 13 9
7 13 3 15 1 0 7 0
13 0 3 0 9 3 13 11 7 0 1 9 15 9
26 10 3 11 13 10 9 9 1 9 9 13 11 3 1 15 13 1 10 9 9 13 9 15 13 9 11
25 13 3 3 0 10 9 9 0 7 3 9 15 3 15 1 10 0 9 13 3 3 10 9 10 9
25 0 3 10 0 9 13 0 3 10 0 11 10 0 13 11 0 9 11 11 11 11 11 11 11 11
6 0 12 9 9 10 0
7 12 3 15 13 11 1 9
15 0 3 10 9 9 3 13 13 0 9 9 3 13 3 3
5 11 3 3 13 9
20 3 3 10 9 10 0 13 10 0 9 3 9 13 11 10 9 13 13 10 9
14 13 3 15 9 9 13 10 9 13 10 9 13 11 9
14 13 3 0 0 13 15 10 12 9 7 13 15 0 9
13 0 3 3 10 0 0 9 1 10 1 10 11 13
3 13 3 0
14 1 11 3 12 13 9 7 1 10 12 9 13 0 12
12 10 3 0 9 13 0 9 13 3 3 0 13
11 0 3 3 3 13 7 13 15 3 13 9
4 15 3 3 13
22 0 3 13 10 9 10 9 3 13 9 9 3 3 15 13 9 10 7 11 9 7 11
30 13 3 0 1 11 13 1 11 15 0 10 0 15 9 13 11 13 11 0 9 9 10 11 15 9 13 3 15 3 13
21 0 13 10 9 13 11 13 10 13 15 9 15 13 9 0 7 15 9 0 15 13
9 13 3 15 13 1 10 9 10 9
13 15 16 15 13 3 10 9 9 13 0 7 10 0
42 1 0 13 10 3 11 11 9 9 10 3 9 10 7 11 7 10 10 0 9 11 9 9 13 13 0 1 11 11 7 3 13 7 10 9 1 15 9 13 10 0 13
28 10 7 3 11 15 13 0 7 10 0 9 7 9 7 7 0 1 15 13 7 13 0 1 3 9 0 13 9
18 16 3 13 10 11 1 10 11 10 9 13 10 11 1 7 11 7 11
24 13 3 1 9 3 10 9 13 15 10 1 10 11 9 7 13 7 10 0 9 13 1 15 13
11 13 3 1 10 11 13 11 13 1 10 9
11 13 3 1 9 0 10 11 13 1 11 0
8 11 15 13 9 10 13 0 15
10 3 13 9 3 13 9 13 7 0 13
16 3 3 15 3 3 13 13 3 16 15 9 13 10 9 15 13
15 3 3 3 15 9 10 3 0 15 3 9 13 15 13 13
12 0 3 9 10 9 13 7 3 13 16 15 13
7 15 3 3 15 3 13 13
10 15 3 13 0 13 16 0 13 10 11
6 6 9 10 3 9 13
19 15 3 3 15 9 13 7 9 0 13 0 13 7 10 0 7 10 3 13
12 10 3 3 0 15 7 13 7 15 9 13 13
14 9 3 9 13 0 15 13 16 7 13 7 0 15 13
8 13 3 15 13 9 0 3 13
11 13 3 15 9 7 13 10 9 7 9 13
12 13 3 15 13 7 7 13 7 13 13 10 9
17 7 3 15 6 9 9 1 9 13 13 16 15 0 15 13 16 13
42 11 3 3 0 15 13 0 0 13 9 3 13 13 15 13 16 16 3 0 9 13 3 13 15 13 13 3 16 3 0 3 10 9 16 10 13 13 13 1 10 9 13
12 11 3 13 10 9 7 13 10 9 13 15 13
13 15 3 3 0 1 10 9 13 13 1 9 10 9
35 11 3 10 9 13 1 10 11 10 11 9 9 15 3 3 13 16 3 13 3 13 10 1 11 1 11 0 3 10 9 13 10 11 9 13
11 1 0 3 9 9 10 15 9 10 9 13
12 11 3 1 0 13 1 10 11 9 13 13 11
15 13 3 3 9 1 0 13 15 9 7 15 7 9 13 13
10 10 3 9 0 13 10 0 1 11 9
17 13 3 10 0 1 10 9 9 13 1 11 15 15 13 9 13 13
9 0 3 16 13 13 10 0 13 13
43 13 3 3 10 9 11 10 9 9 10 9 13 0 13 3 13 0 0 13 7 10 9 7 13 10 9 3 13 3 16 15 10 0 1 11 13 13 15 9 15 3 11 13
23 15 3 13 10 9 9 10 9 1 0 3 13 13 16 3 15 1 15 15 13 3 15 13
4 15 3 0 13
12 15 3 3 10 0 15 9 13 13 13 11 9
8 1 0 10 11 1 9 13 0
17 13 10 9 3 13 10 9 7 0 15 13 13 9 9 1 10 9
6 0 9 15 0 13 13
7 10 9 15 1 10 9 13
7 11 3 3 13 1 0 13
6 0 3 13 10 9 13
5 15 3 3 13 0
18 6 13 16 3 13 0 13 16 3 10 0 1 9 9 13 1 10 9
20 0 16 13 13 10 0 3 13 7 13 13 7 1 15 13 13 13 15 1 11
7 3 3 13 0 3 13 3
3 3 3 13
17 0 3 16 13 0 13 1 10 0 13 9 1 11 13 11 1 11
10 3 3 1 9 11 0 13 1 9 13
10 10 3 11 0 13 9 10 11 11 0
12 11 3 3 13 10 9 13 1 9 13 11 13
27 13 3 9 0 3 0 13 16 9 15 1 10 11 0 7 9 13 9 13 9 15 7 9 13 9 10 3
5 9 3 3 11 13
9 11 3 1 0 13 1 10 13 11
5 7 0 3 11 13
13 0 3 11 9 15 13 9 13 10 9 11 7 3
6 1 3 0 3 9 13
17 0 10 9 3 1 11 9 13 16 13 1 10 11 13 10 9 9
12 16 3 0 13 10 3 9 13 1 10 9 13
9 10 3 9 0 9 0 0 9 13
17 7 10 7 11 7 10 11 7 10 11 7 10 11 0 13 15 13
7 13 3 3 0 9 7 0
16 13 3 1 10 11 0 13 10 9 10 0 15 9 3 13 11
5 13 3 11 12 9
6 13 3 15 12 7 12
25 3 3 16 0 3 3 13 10 9 15 3 13 10 9 1 15 16 13 13 15 9 9 13 10 9
19 3 3 3 10 9 10 9 3 0 9 13 0 3 15 9 0 7 3 13
9 10 3 3 9 10 9 9 0 13
14 10 3 9 13 10 9 13 13 13 9 12 7 3 13
13 16 15 3 13 15 13 0 13 10 9 1 10 9
16 10 3 11 13 13 3 3 15 0 13 13 3 3 15 13 13
58 16 15 3 10 11 1 10 9 13 10 9 10 9 1 0 13 10 9 13 9 7 9 7 9 15 3 3 3 10 9 10 1 10 9 7 10 15 9 1 15 15 9 7 9 7 9 13 10 3 15 15 13 7 0 13 13 1 11
8 10 3 11 13 9 13 10 9
5 11 3 3 3 13
22 13 3 1 10 11 0 13 1 10 11 13 10 9 10 9 15 13 13 1 11 10 9
14 3 3 16 0 15 13 13 0 9 10 13 15 10 9
21 13 3 15 1 10 11 0 10 9 13 9 7 7 9 10 9 7 10 9 10 9
8 0 3 13 13 3 1 10 11
6 15 3 15 10 9 13
5 13 1 10 11 13
18 16 3 1 10 11 13 13 0 1 10 0 13 1 9 12 7 9 13
13 13 3 1 15 0 9 13 9 7 0 9 0 12
17 10 3 9 13 3 15 10 9 13 9 12 13 1 10 0 13 9
10 13 3 10 9 0 15 9 10 9 13
7 10 3 3 12 15 9 13
7 10 3 12 10 13 13 0
4 13 3 10 9
31 13 3 1 10 11 13 10 9 7 10 9 7 10 0 9 15 0 7 13 10 9 15 13 7 3 13 10 11 13 1 11
13 10 3 13 9 10 9 10 7 0 7 10 9 13
10 10 3 0 1 11 13 13 13 10 9
13 10 3 11 15 13 13 15 3 3 10 0 3 13
11 7 3 13 15 3 7 9 0 7 0 13
8 7 0 3 10 9 0 9 13
21 13 3 0 1 9 9 13 16 10 11 15 10 11 13 13 9 13 7 3 10 9
9 11 3 3 1 10 1 11 3 13
6 0 3 0 3 0 13
12 0 3 3 9 0 10 9 3 13 13 10 9
12 13 3 7 13 13 1 9 0 7 10 13 13
13 0 3 3 7 0 15 13 0 11 9 13 9 13
6 3 3 10 0 11 13
20 16 3 10 1 10 9 9 13 11 10 10 9 13 9 13 0 15 0 13 11
27 13 3 9 7 13 15 0 1 10 11 13 9 11 9 9 13 9 0 15 16 13 13 3 15 13 9 3
30 15 13 0 9 9 13 13 1 11 7 3 9 12 13 15 9 3 3 13 15 9 13 9 7 0 0 13 7 13 0
10 0 3 11 10 9 9 1 13 9 13
7 0 3 3 15 9 0 13
12 13 3 0 9 3 13 1 10 9 1 10 9
9 15 3 16 11 13 13 15 10 9
26 3 3 11 7 13 9 0 7 13 10 9 10 0 13 9 0 10 9 0 1 0 3 10 9 0 3
9 7 15 0 9 13 15 10 9 13
26 7 3 1 10 9 9 13 9 13 10 13 7 1 10 9 10 9 13 7 9 9 0 13 10 13 0
21 3 3 10 9 9 0 0 9 7 7 9 13 1 10 9 7 3 1 10 9 13
8 1 3 3 9 3 9 13 13
25 3 3 0 3 13 0 10 9 7 13 0 15 13 0 9 7 10 9 10 0 3 13 15 3 3
10 10 3 11 7 10 11 13 13 11 9
17 0 3 3 13 15 3 13 0 9 0 10 9 13 0 3 3 13
7 10 3 0 0 13 15 13
6 0 3 1 11 13 13
19 15 3 0 13 1 9 7 7 9 3 13 1 9 7 9 7 9 7 9
6 7 0 3 9 0 13
10 15 3 3 0 13 0 10 0 13 0
6 10 3 9 3 9 13
31 16 3 1 11 11 10 11 13 3 0 1 10 9 11 13 1 10 9 1 11 3 3 1 10 11 10 9 0 1 9 13
9 9 3 15 3 0 15 3 0 13
10 12 3 0 0 13 7 0 0 13 9
16 13 3 0 10 0 15 13 13 15 3 7 10 9 13 10 9
17 16 3 9 9 3 10 0 15 9 0 7 9 13 0 10 9 13
24 10 3 3 9 15 0 9 13 13 1 11 7 0 10 9 13 15 7 15 9 0 10 9 13
8 13 3 7 15 7 0 0 0
5 1 3 15 15 13
32 7 3 0 9 13 10 0 3 3 15 7 0 13 13 10 13 10 9 10 7 0 10 9 7 3 10 1 10 9 13 10 9
7 13 1 11 0 13 10 0
6 9 3 3 13 7 13
8 11 3 3 13 9 16 3 13
20 0 3 0 10 11 13 10 7 9 13 7 11 13 1 10 9 3 15 0 13
7 13 3 9 13 1 11 0
18 10 16 15 13 0 13 0 7 7 10 0 10 9 10 11 9 0 13
4 3 15 0 13
5 9 3 3 9 13
31 13 3 7 13 1 10 9 13 1 10 9 10 7 9 7 10 9 7 10 9 7 10 9 7 3 13 10 9 15 0 13
12 0 3 13 7 13 9 0 13 13 15 0 13
14 10 3 3 0 13 0 13 10 0 3 12 9 13 9
11 10 3 12 9 0 13 3 13 7 3 13
14 10 3 3 11 3 13 10 11 3 3 3 10 11 13
9 3 3 10 0 10 0 13 10 0
21 10 3 3 3 10 11 11 0 13 10 3 3 15 0 11 15 9 13 7 15 13
10 11 16 10 15 10 9 0 13 0 13
14 13 1 9 0 9 13 9 0 12 7 12 9 13 0
11 0 9 10 9 10 9 13 0 12 7 0
10 10 3 3 9 0 13 10 9 10 0
9 13 3 3 15 15 9 15 15 13
26 9 3 0 15 0 7 7 0 7 0 9 13 3 3 9 12 3 9 0 13 10 9 9 3 12 9
11 10 3 0 9 10 0 13 9 0 12 9
21 13 3 15 1 0 3 13 3 7 1 10 9 10 9 13 7 10 9 15 9 13
8 13 3 9 0 13 15 1 9
29 3 3 9 13 9 0 7 1 12 9 9 9 9 13 13 0 3 10 9 10 9 0 3 0 10 9 10 0 9
13 1 3 10 9 1 10 0 9 0 13 13 1 15
8 10 0 3 10 9 13 0 9
15 9 3 13 1 10 9 12 0 15 7 9 7 7 9 3
10 13 3 0 9 13 12 9 9 1 11
3 11 9 15
5 3 13 9 3 0
7 13 3 3 10 11 9 0
6 13 3 12 9 10 9
10 10 3 0 15 9 13 15 9 13 11
10 13 3 1 0 13 0 7 0 7 0
7 13 3 0 1 10 0 9
11 10 3 3 9 0 10 9 1 10 9 13
15 10 3 1 0 10 9 1 9 0 10 9 9 9 0 13
20 1 3 3 0 9 1 10 9 10 1 10 9 9 13 15 3 10 9 0 9
7 0 3 3 10 9 9 13
14 0 3 3 9 13 3 0 15 0 10 0 9 0 3
38 1 3 9 0 10 9 13 1 0 1 10 3 10 9 0 0 7 7 0 1 3 10 0 11 11 9 0 3 1 15 3 0 13 12 9 3 13 0
32 1 0 3 10 9 9 0 13 9 7 10 9 7 10 9 7 1 0 10 9 0 9 13 7 0 3 1 0 1 15 12 9
12 9 3 1 15 3 3 1 15 10 9 13 13
17 13 3 3 10 9 13 9 7 7 9 0 1 15 13 13 10 13
14 1 3 10 9 9 0 13 3 13 7 15 9 13 0
34 9 3 3 13 15 3 13 7 9 15 13 9 3 3 9 0 10 0 15 3 10 9 13 1 15 3 13 10 0 13 9 0 10 9
12 3 3 3 3 13 1 10 10 11 10 9 9
9 15 3 0 13 9 0 1 9 13
13 7 3 3 1 11 10 11 10 9 10 9 16 13
7 3 3 3 3 13 9 3
12 16 3 13 3 3 13 10 9 3 1 10 9
22 1 3 10 0 9 3 13 9 12 9 9 0 10 0 3 16 10 9 13 10 9 0
16 13 3 1 10 9 0 3 10 9 0 3 9 12 9 0 0
5 15 3 15 3 13
11 0 10 9 11 3 10 11 13 3 13 13
14 11 3 10 11 13 7 10 9 13 13 3 13 10 9
7 10 3 3 9 0 3 13
6 13 3 3 0 9 0
23 10 3 0 13 10 0 9 12 0 13 15 9 13 11 15 3 13 9 1 10 9 13 0
10 0 3 13 10 9 1 10 9 15 13
25 10 3 3 0 13 0 9 15 9 13 11 15 3 0 13 10 0 13 0 3 9 13 15 15 13
27 0 3 10 9 13 9 0 7 7 3 13 7 0 7 13 9 15 3 3 3 3 10 11 13 15 13 3
11 10 3 9 9 13 1 15 13 10 11 11
27 7 3 15 3 13 1 0 10 9 1 9 13 10 11 9 3 7 1 10 0 0 9 13 7 1 12 9
5 0 3 3 0 13
31 3 3 0 11 13 9 9 0 15 13 1 10 9 9 3 1 10 9 3 13 9 3 10 9 15 13 12 7 7 12 9
15 10 3 13 9 1 0 10 9 13 1 10 9 10 9 13
11 16 3 15 13 9 13 9 3 1 15 13
40 13 3 0 0 10 7 9 0 7 10 9 15 9 16 10 7 9 0 13 1 9 0 13 7 10 9 13 0 1 10 11 1 7 10 9 13 9 10 9 0
27 1 0 3 13 10 9 3 10 7 9 13 7 10 0 10 1 9 9 16 3 13 10 9 13 15 10 9
6 0 3 1 15 9 13
5 0 3 3 0 13
3 13 9 0
21 0 3 1 0 3 3 10 9 10 9 15 13 13 9 13 10 9 9 7 7 9
17 13 3 1 15 16 3 9 13 9 0 1 15 10 9 13 10 0
17 10 3 9 10 9 0 13 0 1 16 3 13 10 9 13 1 15
44 16 3 10 7 13 9 0 13 1 10 9 7 10 1 10 9 13 10 11 9 1 10 0 9 1 10 9 13 7 3 10 13 9 13 1 9 13 13 7 10 9 9 13 13
10 10 3 0 0 9 3 9 0 15 13
8 13 3 1 10 9 9 13 0
8 3 3 3 3 13 3 3 13
3 3 3 0
12 0 10 9 13 0 16 15 1 11 13 10 9
23 11 3 7 0 13 13 10 9 0 15 13 7 9 13 7 0 10 9 13 3 3 13 15
16 10 3 9 0 15 13 0 1 16 1 9 15 13 10 0 13
15 13 3 10 9 13 9 3 3 10 3 0 7 9 13 0
13 16 3 0 7 13 9 7 0 3 3 0 9 13
36 13 3 3 9 10 0 7 9 3 13 1 9 7 9 7 3 3 9 1 10 11 9 3 13 10 1 11 13 15 0 13 9 7 0 15 9
21 0 3 10 11 10 9 13 0 3 9 0 0 13 1 9 0 13 3 3 13 3
7 0 3 15 13 0 13 13
13 1 3 10 9 13 10 1 11 9 13 10 9 3
18 13 3 13 0 13 9 12 7 12 1 0 10 9 10 11 13 15 9
6 13 3 10 9 13 13
9 15 3 9 0 13 13 3 10 9
9 3 3 10 0 15 3 0 13 13
6 10 3 0 13 13 15
19 16 3 13 13 1 10 9 13 7 10 0 7 13 10 9 13 1 10 9
21 15 3 13 3 0 10 11 3 13 7 13 15 15 9 3 13 13 9 9 3 0
8 3 0 3 9 13 10 9 15
15 11 3 9 13 3 9 7 13 0 3 7 15 10 9 13
18 7 3 3 0 15 13 13 7 3 15 13 15 13 15 13 13 3 0
41 13 10 9 0 1 9 10 9 3 1 10 9 13 7 1 3 10 9 13 0 3 13 1 10 9 10 9 13 10 9 3 0 10 9 13 13 13 3 1 10 9
15 3 7 3 13 7 1 0 13 13 0 1 10 0 10 9
32 13 3 0 0 10 9 15 3 13 1 0 0 1 10 9 10 11 9 13 9 3 1 0 9 3 3 1 0 13 1 10 11
26 16 3 3 13 7 13 10 0 10 1 10 11 13 15 3 3 13 10 9 13 1 10 9 13 3 0
29 13 3 3 15 10 1 10 9 9 13 7 0 1 10 9 13 10 1 10 9 10 9 13 13 3 15 3 1 9
8 3 3 1 0 15 13 10 9
7 7 11 3 3 3 0 13
18 10 3 9 10 0 0 3 7 15 13 15 15 13 3 3 3 7 0
18 9 10 0 1 9 15 7 7 10 9 13 1 10 9 9 15 15 13
10 3 0 10 0 9 10 9 10 0 11
8 13 3 0 10 9 0 12 9
25 9 3 0 0 3 15 9 13 16 12 10 1 10 9 9 0 10 0 13 0 10 9 13 9 13
8 0 3 10 9 10 11 13 13
17 10 3 9 10 0 13 3 0 7 0 13 10 9 10 9 13 0
31 13 3 1 10 9 13 7 10 9 7 13 10 9 3 3 3 1 11 0 10 9 13 1 10 9 7 9 7 7 9 13
12 10 3 0 9 15 3 3 10 0 13 1 9
15 10 3 3 0 9 3 13 9 13 7 9 7 9 7 9
16 10 3 10 11 9 3 0 13 13 16 1 12 3 10 3 13
16 10 3 9 3 10 7 9 7 10 9 10 9 13 12 3 9
22 13 3 15 9 13 1 15 10 9 10 0 15 0 1 15 7 9 7 9 7 9 13
37 15 9 9 13 10 7 0 7 9 15 9 9 13 0 10 9 13 10 0 10 9 16 13 7 15 10 9 10 9 13 7 3 13 10 9 10 9
14 9 3 3 13 1 10 11 10 9 3 3 3 10 9
16 10 9 15 13 10 1 10 9 13 1 10 11 13 0 15 0
18 13 3 1 7 12 9 7 12 9 0 13 7 15 3 3 13 10 9
4 15 3 3 13
10 13 3 7 3 0 0 10 9 7 0
12 1 0 3 9 9 0 13 1 3 10 0 0
22 16 3 13 13 1 10 11 7 13 10 9 9 3 10 9 7 10 9 15 1 3 13
11 10 3 9 13 1 10 9 13 1 10 0
16 1 10 9 3 3 3 0 7 13 13 15 9 1 0 10 9
16 16 3 10 9 13 13 3 1 10 0 0 9 10 0 13 9
7 10 3 3 9 15 13 0
10 13 3 10 9 9 13 13 15 10 9
7 9 3 0 13 7 9 0
9 1 3 9 3 15 9 13 13 9
9 0 3 3 15 9 1 10 9 13
5 9 3 15 3 13
9 1 9 0 3 10 9 0 13 0
6 1 3 15 13 9 9
13 13 3 1 12 0 9 13 0 3 10 0 1 15
16 3 3 16 0 13 0 9 13 0 3 13 15 1 0 13 0
4 13 3 1 9
39 16 3 3 13 10 9 13 10 0 10 9 13 3 10 0 7 16 15 15 0 13 7 0 3 13 15 13 0 9 13 13 15 16 15 10 10 0 13 13
18 10 3 3 9 13 1 10 0 9 7 3 10 0 10 0 7 0 13
10 13 3 3 1 0 13 9 10 13 13
15 15 3 15 13 3 13 16 3 13 15 7 1 0 9 13
16 16 3 13 13 7 13 15 15 10 9 9 13 13 10 0 9
6 10 13 1 10 9 13
5 3 3 3 13 9
14 9 3 13 10 13 3 15 13 16 3 13 15 9 13
6 9 3 0 10 1 11
8 3 3 10 9 10 0 0 13
6 9 3 13 13 3 0
7 9 3 15 13 16 3 13
7 10 0 3 0 3 0 13
10 10 3 3 0 10 9 13 10 0 0
15 13 15 9 0 13 1 9 11 3 1 10 9 13 9 9
20 0 3 3 3 13 13 10 15 15 9 13 1 9 1 9 13 1 10 9 13
12 1 9 11 13 9 1 10 9 13 9 0 9
4 15 3 3 13
3 15 3 13
16 0 3 9 15 9 9 13 1 10 9 1 15 10 9 13 13
23 3 16 13 9 3 0 13 1 10 9 3 15 15 9 9 13 1 10 9 13 3 10 9
5 13 3 13 13 0
5 13 15 10 9 11
6 11 3 13 10 11 0
5 3 3 15 9 13
6 13 3 0 0 10 9
8 10 3 0 13 13 7 13 15
10 16 3 13 13 10 9 13 1 10 9
13 7 10 1 0 3 3 0 15 15 13 3 15 13
11 15 3 3 9 7 13 13 7 9 0 13
13 15 3 0 15 13 9 0 13 3 13 10 9 13
8 3 3 0 7 0 0 9 13
10 10 3 9 0 7 0 13 13 7 0
10 13 3 15 3 0 13 0 10 9 13
11 10 3 11 13 7 0 7 0 13 10 11
22 9 3 1 15 9 9 0 0 13 13 1 3 15 9 15 13 3 9 10 9 13 0
15 9 3 1 9 13 15 1 9 13 0 7 0 13 10 0
6 0 3 0 13 9 13
15 9 3 13 12 15 10 15 1 12 1 9 7 7 9 13
14 10 3 12 10 9 10 11 13 1 0 1 10 11 9
20 15 3 3 9 13 15 7 10 3 9 9 10 11 13 7 10 0 12 13 13
24 10 3 11 13 0 1 15 13 9 3 9 9 13 12 9 9 3 3 0 13 15 15 12 9
21 7 10 3 1 10 9 13 10 9 0 10 11 13 13 9 7 9 0 7 9 0
18 9 3 9 0 7 0 1 15 13 10 11 10 0 15 1 9 0 13
22 1 15 3 9 9 0 9 13 13 13 15 13 7 7 13 9 9 15 1 10 9 13
14 10 3 9 3 13 7 13 10 0 9 3 3 13 9
14 10 3 3 1 9 10 9 0 10 11 13 10 11 13
14 10 3 1 9 7 7 9 13 9 13 9 0 1 9
11 0 7 3 15 7 0 10 13 7 13 13
19 0 3 10 9 10 13 0 15 13 9 0 3 10 9 10 1 10 9 13
11 3 3 13 13 11 0 13 0 10 9 13
9 13 3 10 9 13 9 10 9 9
4 11 15 13 9
15 10 3 11 13 3 15 15 13 7 10 9 9 13 10 9
39 11 3 1 0 16 15 9 3 13 13 1 10 11 13 1 10 0 1 10 9 9 9 7 13 1 10 9 9 10 9 7 9 1 9 10 13 10 9 13
12 13 3 15 0 10 9 13 10 11 9 13 0
11 3 3 3 13 16 15 1 9 13 0 13
13 13 3 13 10 15 7 15 13 13 13 15 3 13
12 3 13 9 0 13 7 3 3 3 1 9 13
16 15 3 16 3 13 11 13 13 9 3 15 13 13 10 9 13
14 16 3 15 13 13 3 1 10 15 15 10 0 0 13
9 0 3 13 10 11 13 9 10 0
12 13 3 0 1 0 15 13 10 9 13 15 13
19 15 3 1 10 0 10 9 13 13 13 11 7 7 10 9 15 1 10 9
8 10 3 15 9 13 0 9 13
17 16 3 0 13 13 7 9 0 13 15 3 13 9 9 15 15 13
21 16 3 13 16 9 7 15 13 7 0 0 13 0 0 13 16 9 10 0 13 9
12 3 3 13 9 1 10 13 9 10 0 3 0
15 16 3 13 13 10 0 1 10 9 0 15 1 15 9 13
6 13 3 13 15 10 9
16 0 3 3 16 13 9 3 10 3 13 7 1 9 10 15 13
15 13 3 3 13 0 15 16 13 1 15 0 13 9 13 13
17 1 3 10 13 0 7 3 0 11 3 10 11 9 13 13 10 9
17 3 3 15 13 13 13 15 3 0 13 3 3 0 13 13 0 13
28 0 3 10 9 10 9 3 0 13 7 13 13 1 10 9 10 15 9 3 3 3 9 3 9 0 7 9 0
15 13 3 0 13 10 9 10 0 10 0 3 13 1 10 9
22 16 3 15 9 3 13 0 13 0 0 13 7 1 15 7 15 10 3 13 9 9 0
4 9 3 0 13
18 11 3 13 10 0 9 15 11 3 13 13 11 13 3 15 13 1 0
7 15 3 3 13 3 13 0
28 13 10 11 1 10 9 13 10 11 9 10 0 13 1 10 9 9 7 0 15 3 10 11 15 3 10 11 13
6 3 3 13 3 9 13
12 16 3 3 13 10 11 13 9 15 1 10 9
14 16 3 15 13 0 13 10 9 13 11 7 13 0 13
11 11 9 15 13 15 7 7 10 15 9 13
7 3 3 0 3 13 15 13
9 15 9 13 7 15 15 13 10 13
29 3 3 1 10 13 9 13 13 10 15 9 10 0 13 1 10 9 9 7 0 15 3 10 11 15 3 10 11 13
12 15 3 10 9 13 16 0 3 13 3 3 13
7 10 3 9 15 13 1 11
6 13 3 3 10 11 0
10 6 9 3 13 9 9 13 15 15 13
6 16 3 13 13 3 3
15 15 1 3 9 13 0 9 13 1 3 13 1 0 13 0
23 16 3 15 15 9 13 9 10 15 0 13 1 15 15 15 13 13 15 0 15 15 15 13
16 11 3 0 13 7 13 10 11 13 1 9 13 11 10 9 11
44 1 3 0 11 7 7 9 10 0 9 13 3 1 10 11 13 3 10 0 13 10 9 9 10 9 10 7 13 10 11 9 13 13 7 10 13 13 9 16 13 10 0 13 13
6 13 3 9 7 9 13
8 10 3 9 13 0 3 15 13
19 0 3 3 0 13 7 15 7 10 10 9 11 9 13 9 15 9 13 11
20 15 3 13 10 7 1 10 9 13 7 10 1 10 9 13 9 1 11 13 0
8 3 3 15 3 13 13 10 9
15 13 15 10 9 13 1 0 10 9 0 9 9 10 9 13
11 16 3 0 3 13 9 13 15 10 9 9
25 10 3 10 9 11 9 11 16 15 10 7 9 13 7 13 16 13 0 13 11 1 10 9 13 13
11 16 3 13 7 3 7 10 9 13 13 15
7 7 3 0 3 9 0 13
14 11 3 16 15 11 3 13 13 15 10 15 9 13 11
19 0 10 9 15 3 0 9 9 13 13 0 13 7 3 3 13 3 0 13
9 0 3 3 13 15 13 1 15 13
15 3 3 16 15 10 9 13 13 10 9 7 7 10 0 13
5 9 3 10 9 13
15 9 3 13 9 0 11 13 1 10 13 10 9 10 11 9
10 16 3 13 13 15 10 9 1 10 9
6 13 3 10 9 13 0
15 15 3 15 13 7 7 13 15 9 13 9 10 15 13 9
8 15 3 15 3 3 13 9 13
17 10 3 3 1 10 11 9 10 9 0 9 13 0 15 10 0 13
16 9 3 13 7 0 15 3 13 7 9 7 7 9 9 13 13
7 9 3 7 9 10 15 13
10 15 3 1 9 7 9 7 9 9 13
23 3 3 3 10 9 10 3 1 10 9 0 9 13 10 3 1 10 9 7 9 7 9 9
6 9 3 7 9 13 15
15 7 3 3 15 13 1 10 9 10 3 9 7 10 9 0
4 9 3 13 0
4 0 3 0 13
13 15 3 9 13 9 13 3 9 13 10 13 7 9
14 15 3 13 9 9 9 10 9 13 1 10 9 13 3
17 16 3 9 13 3 10 13 10 15 13 13 15 7 15 9 1 15
5 13 3 10 9 13
6 0 3 10 0 15 13
17 10 3 9 13 3 13 7 9 13 9 13 16 3 13 1 10 13
8 9 3 0 9 13 15 13 9
5 9 3 0 10 9
10 10 9 10 0 15 10 9 10 0 13
24 10 3 0 13 9 13 3 9 13 0 7 3 10 9 15 13 0 3 15 0 3 15 10 9
8 9 3 3 1 15 13 10 11
6 9 3 13 1 15 13
5 13 3 1 10 11
7 13 3 10 9 13 9 0
23 0 3 0 3 0 13 3 13 7 15 0 0 3 3 3 3 13 11 7 7 0 3 11
12 7 10 15 9 13 15 0 13 13 10 9 11
24 13 3 9 10 11 9 3 13 0 7 0 1 10 0 3 13 13 1 9 15 13 13 7 0
20 0 3 16 13 1 10 9 7 10 9 13 10 9 13 10 0 13 3 0 9
12 16 3 13 9 7 0 0 13 13 10 0 9
17 13 3 10 0 10 9 16 1 10 0 13 13 15 10 9 10 9
18 0 13 12 9 15 3 15 0 13 12 15 13 10 0 15 13 1 11
16 13 3 1 10 9 13 13 13 7 10 11 7 15 0 13 13
8 10 3 11 15 1 0 13 0
14 16 15 15 11 0 13 0 3 13 13 3 13 9 15
9 13 3 0 10 1 10 11 13 3
15 3 3 3 15 13 10 9 10 9 16 3 13 1 0 11
6 0 13 10 9 12 9
27 13 3 15 3 10 9 13 1 9 7 10 0 10 9 16 13 10 9 3 13 13 10 9 10 9 9 13
7 13 3 10 9 0 9 11
9 13 3 15 1 9 13 13 11 13
6 9 9 3 15 0 13
5 3 3 10 9 13
32 1 3 3 11 7 10 9 10 9 13 1 12 9 7 10 9 15 11 13 12 9 13 10 0 13 0 15 9 1 10 9 13
18 1 3 10 0 11 10 0 13 9 15 13 13 10 11 13 13 0 11
15 15 3 3 1 11 0 0 13 9 13 3 15 3 13 13
41 13 3 9 0 1 10 11 13 9 0 10 0 9 7 10 9 15 15 9 13 9 15 10 7 9 13 7 13 1 10 0 13 1 11 13 15 0 11 10 11 9
10 15 3 13 9 0 0 13 1 10 11
19 10 3 0 13 1 11 9 7 1 9 11 13 7 10 0 7 13 10 9
19 3 3 3 13 0 10 0 9 7 13 13 3 16 0 15 15 13 1 11
10 1 0 0 3 0 13 11 13 1 15
7 0 3 10 11 9 13 11
31 15 13 0 10 15 9 13 16 15 15 0 13 13 1 0 9 10 11 7 1 15 13 13 9 0 15 3 7 3 11 13
15 3 3 11 1 10 13 7 10 9 7 13 10 0 0 13
12 10 3 9 13 15 13 13 1 10 0 10 9
20 10 3 11 13 13 16 3 1 11 7 10 11 13 13 7 13 10 9 13 15
12 13 3 13 10 0 0 16 12 9 0 3 13
16 1 3 10 9 0 11 3 13 7 7 9 13 10 9 11 13
12 11 3 10 9 10 11 9 13 15 9 13 11
15 13 3 10 9 10 11 10 9 11 0 7 13 7 3 0
17 10 3 0 1 10 13 9 13 1 11 13 15 9 13 0 3 13
18 0 3 10 9 13 1 10 11 7 13 0 0 3 0 13 15 0 13
22 0 3 10 9 11 9 13 7 9 10 0 15 15 0 13 10 9 1 0 10 9 13
9 1 3 3 0 10 11 3 13 13
12 1 3 10 0 9 11 0 9 1 10 9 13
24 11 3 10 11 7 10 0 7 11 3 13 13 1 15 10 9 11 13 7 13 10 10 9 9
7 3 13 13 7 13 1 11
9 10 3 9 15 1 11 10 11 13
14 13 3 1 0 10 11 13 9 15 13 15 1 10 11
19 15 3 13 10 13 0 3 13 3 0 13 0 3 0 10 13 15 13 9
7 0 1 15 3 10 13 13
10 0 15 13 9 10 11 9 0 7 9
4 13 3 3 9
17 13 3 3 10 11 10 0 9 10 11 13 0 9 13 7 3 9
15 10 3 11 0 10 9 13 1 11 13 15 9 1 9 9
6 10 3 11 15 13 0
15 1 3 12 11 7 11 12 12 9 9 13 15 11 13 11
8 15 3 0 13 13 1 10 15
15 16 3 10 9 13 0 9 3 13 10 9 7 13 1 9
10 16 3 13 10 9 3 13 1 10 0
10 16 3 3 13 7 0 7 9 10 13
5 0 10 11 11 13
10 15 3 15 3 10 3 1 10 9 13
11 15 3 15 13 10 11 1 11 13 1 9
13 0 3 3 0 13 1 10 15 13 7 1 11 13
38 13 3 1 13 10 9 13 0 16 15 10 11 3 13 13 1 10 9 10 9 13 13 0 10 10 0 9 13 7 10 13 9 7 13 0 10 11 13
15 13 3 9 0 15 9 3 10 0 10 9 15 9 13 11
24 1 0 13 7 15 0 7 9 7 10 1 11 9 15 13 13 13 3 3 7 10 9 15 11
14 11 3 3 7 0 7 0 13 10 9 13 9 10 15
14 16 3 13 1 10 11 13 15 10 9 13 13 1 11
12 13 3 15 1 10 11 9 1 11 10 11 13
12 0 3 13 10 11 15 11 11 13 7 9 13
23 13 3 1 10 11 10 11 11 9 13 13 15 13 13 9 16 1 10 9 10 9 15 13
23 13 3 7 13 11 13 9 15 13 0 15 3 0 13 9 13 13 0 16 3 13 10 9
11 11 3 3 9 0 13 1 10 0 9 13
16 11 3 9 11 9 10 15 0 13 7 3 13 9 0 10 0
19 16 3 3 13 10 9 10 11 13 1 10 11 9 13 15 13 15 11 13
6 10 3 0 0 13 15
13 13 3 0 10 11 3 3 10 9 13 1 10 11
8 0 3 3 9 9 10 9 13
10 13 3 10 9 3 15 13 1 11 9
6 10 3 0 13 11 15
5 13 3 1 0 9
8 9 3 13 15 3 10 15 9
11 10 3 9 15 9 1 0 10 9 13 0
15 10 9 3 13 10 9 16 13 10 15 0 13 7 3 13
15 0 3 0 9 0 13 7 10 9 0 10 9 13 13 13
10 15 3 3 10 9 0 13 1 0 13
13 13 3 0 10 9 1 11 1 9 15 9 11 13
34 1 3 10 1 0 9 10 7 11 9 13 15 13 10 0 7 1 10 9 11 9 13 7 11 15 10 0 13 7 10 9 13 1 0
7 9 3 13 0 0 10 0
7 9 3 13 10 1 9 9
4 0 1 11 13
6 1 9 3 3 13 9
6 10 3 1 9 0 13
8 9 3 3 3 7 3 9 13
8 9 3 10 0 13 13 10 0
18 9 3 1 0 10 9 13 9 0 9 13 1 9 1 11 9 10 0
10 9 3 10 0 13 10 3 10 1 11
27 9 3 0 10 1 9 13 9 9 13 0 15 10 9 13 1 10 9 10 9 13 1 11 9 13 10 9
9 15 3 0 7 0 13 15 13 0
16 10 3 9 16 13 13 1 10 9 13 7 3 1 9 13 13
16 9 3 13 0 13 0 0 15 10 9 13 9 0 10 3 9
4 16 9 13 13
18 0 3 13 9 9 9 13 10 9 9 10 0 1 15 13 10 9 13
6 9 3 7 0 13 0
15 13 3 10 1 15 9 0 7 0 13 13 0 10 9 13
11 13 3 1 10 9 13 10 9 7 13 13
10 15 3 3 13 1 10 9 9 0 13
4 9 3 0 13
12 1 10 9 13 13 7 0 1 15 10 0 13
5 9 3 0 13 9
4 0 13 9 0
26 15 3 13 0 9 13 1 10 9 13 3 0 15 13 9 7 16 13 1 10 9 13 10 9 13 15
8 13 3 0 13 10 9 10 9
27 0 3 1 1 9 9 1 10 0 13 9 15 15 9 13 7 15 9 7 7 9 13 0 15 7 13 13
6 0 3 3 1 13 9
28 10 3 1 10 9 13 10 1 9 9 15 9 13 10 3 0 10 9 13 13 10 3 3 7 3 13 1 9
9 1 3 10 9 9 0 9 13 9
13 1 3 15 11 9 13 1 9 13 11 1 9 13
8 1 9 3 1 15 9 12 13
6 1 9 0 13 9 13
14 15 3 3 0 13 15 0 13 13 16 1 0 9 13
19 9 3 13 1 10 9 0 10 9 13 9 15 10 9 0 10 9 13 13
10 13 3 1 10 9 0 10 9 3 9
19 9 3 10 1 9 13 9 10 9 3 3 0 13 3 0 3 10 0 13
9 13 3 1 9 0 15 9 11 13
8 1 3 15 9 13 15 9 11
9 0 3 10 9 0 13 9 13 13
26 11 16 15 13 1 10 11 10 11 13 1 15 0 7 9 7 3 3 9 0 13 11 13 1 11 13
15 7 15 16 13 13 1 11 13 9 9 7 13 1 10 11
11 16 3 13 9 1 10 9 13 9 10 11
26 7 15 13 10 9 9 13 13 11 7 13 10 11 15 13 10 9 13 15 7 10 9 13 7 0 13
60 13 3 10 11 3 3 10 7 9 10 9 13 10 11 15 7 10 9 13 1 10 15 0 13 7 10 9 7 10 1 11 13 10 15 9 16 16 10 9 13 10 0 15 10 1 10 11 13 3 12 9 13 1 10 11 9 0 15 13 9
6 0 3 13 10 9 9
10 0 3 7 10 9 1 10 11 9 13
7 10 0 3 15 13 10 11
26 9 3 0 11 10 9 15 3 13 13 1 15 9 7 7 9 10 0 9 13 10 0 13 15 11 13
10 10 3 13 10 9 1 10 9 9 13
8 16 3 13 15 13 0 13 0
19 9 10 13 3 13 9 7 0 7 9 0 7 1 9 13 13 10 9 3
7 13 3 3 0 9 13 15
14 1 3 11 7 10 9 7 10 9 13 13 1 10 9
21 10 3 11 13 11 13 9 7 10 11 9 7 15 13 15 10 9 13 15 10 11
7 10 3 11 15 15 13 9
11 9 3 0 10 9 13 7 13 3 7 13
26 16 3 9 10 9 0 13 13 1 10 0 10 9 0 9 7 15 3 13 10 9 10 9 0 9 13
8 0 3 10 0 10 9 9 13
15 1 3 10 0 9 9 13 13 1 11 10 0 1 0 9
33 1 3 10 9 0 3 1 12 9 9 9 13 9 1 9 0 1 9 7 1 9 0 10 9 13 1 0 10 9 9 0 7 0
13 1 3 15 9 13 0 1 10 0 7 1 10 0
16 0 3 1 11 1 12 9 9 0 13 10 9 1 10 0 11
16 7 3 10 1 11 3 3 0 13 15 0 10 11 10 9 13
5 3 3 13 10 9
18 13 3 10 9 13 10 0 16 3 13 7 10 9 7 10 9 13 0
4 3 3 13 3
9 13 7 0 9 7 13 1 1 9
7 9 3 0 10 9 13 9
27 1 3 0 1 10 9 10 9 1 0 12 9 9 9 7 9 13 0 10 0 7 9 7 9 1 15 13
7 10 3 9 0 9 11 13
10 1 0 10 9 10 9 13 10 9 13
20 7 9 13 1 15 15 9 9 13 9 0 3 15 1 10 9 9 13 3 13
7 1 15 3 10 0 9 13
5 0 3 1 0 13
7 10 9 13 13 1 10 3
5 1 0 3 13 13
14 1 3 10 3 3 0 3 13 13 1 10 9 10 9
18 15 3 15 13 10 0 9 3 3 0 3 10 9 1 9 7 7 9
10 10 9 3 0 10 9 9 13 10 0
12 9 3 15 0 0 13 7 13 3 3 10 9
23 1 3 9 1 0 12 9 9 0 9 7 9 7 9 7 9 1 15 13 15 9 13 9
8 15 0 13 0 9 15 15 13
7 0 3 3 15 13 9 9
7 12 3 0 15 9 15 13
24 0 10 9 13 13 7 1 0 15 10 0 13 16 15 13 13 0 7 10 9 7 10 9 15
16 3 3 1 0 12 9 0 9 9 7 9 7 9 1 15 13
10 13 3 10 9 0 9 15 9 13 11
9 3 3 15 13 9 7 9 7 9
9 0 10 9 10 9 13 10 0 13
9 1 0 10 9 10 9 0 0 13
4 13 3 3 9
9 13 3 7 0 15 13 7 9 13
15 1 3 3 10 9 0 13 10 9 10 1 10 9 13 13
5 10 3 1 0 3
12 13 3 3 10 9 1 0 9 7 10 3 0
7 0 3 3 10 11 0 13
11 3 3 3 13 13 10 9 13 0 16 13
11 10 3 9 3 7 0 7 0 10 9 13
30 1 3 10 9 10 1 9 7 1 0 10 11 0 7 0 7 0 7 0 7 0 13 10 9 7 9 13 1 15 15
22 9 3 3 0 3 10 0 9 13 13 1 10 1 11 11 7 7 9 15 7 9 13
11 10 3 10 0 9 3 9 1 10 9 13
5 0 3 3 3 13
19 10 3 3 10 9 9 16 3 15 3 13 3 0 13 13 3 15 0 0
12 13 3 3 3 10 9 9 15 0 15 15 13
8 16 3 1 0 3 13 3 13
4 0 3 3 13
10 16 3 13 10 9 9 13 13 15 9
6 9 3 9 13 13 15
6 13 3 15 13 0 9
10 16 10 9 13 10 9 13 1 10 9
7 0 3 13 13 10 9 15
17 10 3 3 9 7 10 9 10 9 10 11 1 10 9 13 10 9
14 7 3 3 10 9 13 16 1 11 13 10 9 10 9
12 0 3 13 0 1 10 9 0 10 9 13 9
9 1 3 10 0 0 9 10 9 13
10 13 3 15 3 9 1 9 3 0 13
9 7 12 9 13 1 9 10 9 13
12 13 3 10 13 10 9 3 3 10 9 1 9
15 0 3 13 13 13 16 13 10 9 16 15 13 7 0 13
5 9 3 0 0 13
20 10 3 1 9 10 11 9 11 13 9 3 9 7 9 13 13 15 9 13 9
7 15 10 1 0 10 9 13
5 10 3 1 0 13
8 13 3 0 13 10 1 11 9
23 10 3 9 0 7 7 10 0 10 11 10 1 9 0 0 7 7 0 13 10 10 9 9
22 10 3 3 3 1 10 9 10 11 15 10 9 13 13 0 7 7 0 1 10 11 9
17 10 3 1 0 10 1 9 15 10 9 0 7 3 7 0 7 0
17 0 7 3 3 13 9 7 15 3 10 0 1 9 7 7 9 0
10 9 3 7 9 0 1 11 3 3 13
6 9 3 9 0 3 13
19 0 3 3 9 10 10 9 9 9 13 15 15 13 1 0 0 3 13 13
14 9 3 9 9 13 15 10 9 13 10 9 1 10 9
11 0 3 9 13 1 15 9 0 3 9 13
8 0 3 3 0 13 9 9 13
7 13 3 3 15 0 7 13
27 1 0 3 13 0 13 9 15 9 13 11 9 3 12 9 9 3 0 0 1 10 9 9 7 0 7 9
21 9 3 1 15 13 1 15 10 9 10 0 9 9 13 9 1 10 9 9 13 9
4 15 3 13 13
17 13 3 3 15 3 3 1 11 1 9 3 9 9 13 0 15 13
25 1 0 9 13 1 9 9 13 7 3 13 10 9 9 9 3 13 9 10 3 15 10 0 9 0
8 13 3 1 9 13 1 10 9
12 16 3 13 0 3 1 10 9 1 10 9 13
15 15 15 3 3 13 1 10 9 1 9 13 13 1 10 9
14 3 3 3 10 1 10 9 10 1 11 13 13 13 9
11 13 10 11 9 7 7 9 1 0 9 13
20 1 15 16 13 7 13 10 9 13 15 3 1 10 9 13 1 10 9 13 9
23 10 3 0 13 10 9 13 1 10 9 7 3 1 10 9 9 13 7 13 3 1 10 9
5 10 3 0 13 13
12 7 16 3 13 15 0 10 9 10 9 13 13
10 16 3 3 0 13 3 1 10 9 13
12 15 3 13 0 3 3 13 9 16 15 3 13
22 0 3 13 15 15 13 9 13 7 0 10 0 9 10 9 7 15 3 7 3 13 15
5 9 3 7 9 9
19 13 3 15 3 9 13 15 10 11 0 16 7 11 7 11 13 1 11 0
10 10 3 3 0 9 10 9 10 9 13
15 0 3 0 10 0 9 11 9 13 7 13 15 10 0 11
17 0 7 3 13 7 0 9 7 7 9 13 15 7 9 0 13 13
6 13 3 3 0 10 11
12 10 3 9 10 9 10 0 9 10 0 9 13
21 13 3 3 10 0 9 13 0 0 10 11 15 10 9 13 12 9 1 15 0 9
12 0 3 3 10 9 10 9 13 13 7 7 13
16 0 7 3 13 10 1 10 0 9 10 0 13 13 15 9 13
29 13 7 0 10 0 9 7 10 1 10 0 10 9 13 7 7 13 16 13 7 7 13 10 0 9 7 10 0 13
7 3 1 12 9 0 9 13
6 0 3 3 1 0 13
27 10 3 11 0 9 16 1 10 11 13 1 11 13 1 10 11 13 10 9 13 13 10 0 10 9 10 11
12 15 3 15 3 13 10 9 0 3 13 10 9
11 13 15 1 10 9 13 1 10 9 10 9
9 10 3 3 0 13 0 1 15 13
9 1 3 10 13 13 10 9 10 9
11 13 3 3 3 10 0 13 10 9 10 13
5 0 3 3 3 13
6 10 3 9 13 10 0
21 9 3 3 0 13 7 13 15 0 7 3 0 10 9 11 10 9 10 0 13 0
13 1 3 9 10 9 9 9 13 13 10 0 9 0
10 15 3 3 13 16 15 15 13 9 13
38 10 3 9 13 0 15 1 10 0 9 13 9 16 3 10 9 0 3 13 13 10 9 1 9 7 0 7 13 13 9 9 7 9 15 0 13 1 0
28 1 3 10 9 0 3 13 0 0 7 13 1 10 9 7 10 0 13 13 1 10 9 10 13 10 15 9 13
12 10 3 9 13 10 0 9 13 3 1 10 9
25 13 3 0 1 15 13 9 16 13 13 10 0 9 13 3 10 9 15 3 10 9 13 3 3 13
8 13 3 3 13 10 9 1 9
12 10 3 15 9 10 9 13 13 3 0 10 9
21 10 3 0 10 0 9 13 13 10 9 1 15 15 13 9 7 7 10 9 3 0
11 10 3 3 0 10 0 10 9 13 13 3
17 7 16 1 10 0 9 13 10 0 9 15 13 13 15 1 10 9
15 13 3 10 9 11 3 10 10 0 9 9 13 13 10 9
7 11 3 15 10 0 3 13
7 1 11 3 13 0 0 9
5 10 3 0 3 13
14 10 3 9 15 13 9 13 13 7 15 7 12 9 13
11 13 3 10 9 3 13 1 11 9 13 15
7 13 3 0 13 1 10 11
25 13 3 10 3 15 9 10 7 9 1 7 10 9 10 13 15 7 13 13 16 15 1 10 11 13
10 0 10 9 9 10 11 3 1 11 13
14 15 3 13 10 0 0 3 1 10 11 0 13 1 9
20 15 3 10 9 0 9 13 11 15 3 3 3 1 15 13 13 1 9 10 11
9 3 3 3 10 11 3 10 9 13
16 16 3 3 3 1 10 11 13 10 0 13 1 10 11 13 3
15 13 3 9 13 3 3 9 10 3 0 9 1 9 0 13
30 10 3 1 10 11 10 9 13 1 11 15 10 11 13 0 3 0 0 3 13 0 13 11 13 13 0 3 1 9 3
35 10 3 3 1 11 9 13 10 9 13 1 0 7 16 3 13 13 15 10 0 3 13 15 3 13 16 3 3 13 3 13 13 10 9 0
14 13 3 10 0 1 10 9 3 9 0 1 9 15 13
7 3 3 13 10 9 13 15
3 3 15 9
15 3 10 0 13 13 10 9 7 0 7 13 7 13 15 0
9 10 3 3 1 9 0 13 3 13
18 3 3 9 0 1 10 9 13 10 0 10 9 7 7 10 11 13 9
8 0 3 15 13 1 11 11 13
10 9 3 9 0 13 1 3 9 15 9
10 7 3 0 0 15 7 0 3 3 13
5 13 3 1 0 0
7 9 3 13 0 1 9 0
17 9 3 0 0 15 13 1 15 1 9 7 9 7 10 1 0 13
10 0 3 15 3 9 10 13 13 13 15
13 9 3 10 3 0 15 1 10 0 10 0 9 13
19 10 3 13 13 10 13 13 15 15 13 16 13 13 0 13 10 0 15 9
6 10 3 1 0 13 0
4 13 9 0 0
23 16 3 15 15 13 9 13 0 10 9 7 9 9 0 1 0 15 15 13 3 1 10 9
20 15 3 3 13 7 13 13 1 7 9 7 9 13 1 10 9 1 10 0 15
5 13 3 13 10 9
6 10 3 15 9 0 13
6 9 3 15 0 0 13
12 10 3 9 3 13 7 13 15 0 13 9 13
14 10 3 9 3 13 7 13 10 9 1 10 9 9 0
10 7 10 3 13 0 13 10 3 0 0
7 0 13 0 9 3 9 0
7 10 13 1 9 7 9 0
7 0 3 15 10 0 9 13
10 9 3 13 0 0 11 7 11 7 11
22 10 3 9 15 1 10 0 9 13 11 3 9 7 13 0 0 7 13 13 1 11 15
13 12 3 9 13 10 0 7 0 13 9 13 13 0
8 3 3 13 13 7 3 9 13
15 9 3 13 9 13 0 1 15 10 0 9 13 1 9 9
6 9 3 3 9 13 0
30 10 3 1 11 10 9 3 0 15 13 13 10 0 15 13 9 13 15 7 10 1 3 10 11 0 9 13 13 7 0
17 0 3 13 13 13 1 10 11 9 15 9 13 9 9 3 13 0
30 10 3 9 15 13 0 0 10 9 1 12 9 10 9 10 9 0 3 7 0 7 0 9 13 13 3 1 9 13 0
6 13 3 1 0 10 0
11 3 3 0 9 0 13 15 3 3 13 13
8 13 3 3 15 1 10 0 9
18 3 3 9 13 9 13 10 1 10 11 7 1 0 3 13 13 10 3
9 15 3 3 0 13 13 13 3 13
7 10 3 9 0 13 13 0
12 7 15 10 1 10 9 0 13 13 1 10 9
8 0 3 3 10 9 0 1 13
24 11 3 16 13 3 10 11 13 1 11 13 10 1 11 7 10 0 9 7 10 9 10 0 11
12 10 3 3 11 3 13 10 11 9 3 15 13
10 13 3 11 10 9 13 1 15 9 13
5 0 3 3 0 13
13 10 3 11 15 7 3 9 9 7 13 13 11 13
9 13 3 15 0 3 1 15 13 13
19 11 3 13 9 0 13 13 13 11 9 13 0 13 1 10 11 1 10 11
12 13 3 11 13 1 10 9 10 10 9 13 0
23 13 10 9 3 13 0 1 9 13 9 1 10 9 13 7 1 10 9 9 13 7 13 9
18 7 3 0 13 7 0 10 13 1 10 9 7 1 10 1 10 11 0
18 0 3 16 15 13 10 9 15 13 13 13 15 15 13 10 9 10 9
5 15 3 3 3 13
10 15 3 16 13 1 10 9 13 10 9
29 13 3 7 10 9 10 9 13 10 0 9 13 13 10 9 1 10 9 7 13 1 10 9 10 9 7 13 10 9
14 16 3 13 13 3 10 9 15 3 3 3 9 13 0
16 13 3 10 11 0 13 13 10 9 13 9 7 0 13 15 9
34 15 3 15 13 16 13 3 0 13 15 0 13 3 10 11 1 10 11 9 13 10 3 11 3 1 10 11 13 3 9 10 1 11 0
12 15 3 13 16 3 15 3 10 9 13 3 0
8 15 3 3 0 13 3 3 13
7 0 3 3 0 1 3 13
30 3 11 13 9 11 15 13 1 10 11 9 13 13 1 9 9 7 1 15 13 7 15 7 10 9 7 7 10 9 15
7 13 3 13 10 9 10 11
13 15 3 13 7 13 9 1 10 11 13 1 10 11
19 13 3 10 9 10 9 1 15 13 13 13 1 9 13 3 13 10 9 13
11 10 3 3 9 13 0 10 11 9 13 13
12 13 3 10 9 13 1 10 9 15 13 9 0
6 15 3 0 13 3 13
20 10 3 9 16 13 13 10 9 3 13 1 15 0 13 7 13 15 0 10 9
23 10 3 1 7 11 9 7 9 7 9 7 9 7 0 10 9 10 11 3 13 9 1 11
10 13 3 3 10 1 10 9 13 13 3
18 9 1 9 0 13 1 0 13 10 9 9 1 10 9 0 13 12 9
15 13 1 9 15 9 13 11 1 9 0 10 13 12 9 13
5 13 3 0 0 9
9 10 3 9 7 10 9 13 9 9
28 15 3 9 13 0 16 3 10 9 10 0 13 13 9 9 0 1 10 9 7 3 0 15 9 13 13 0 9
9 9 3 3 10 13 13 1 10 11
22 11 3 16 13 10 9 13 9 1 11 9 12 9 15 1 0 0 13 0 1 10 9
12 13 3 0 1 11 13 9 7 7 9 11 9
11 13 3 1 10 11 9 0 3 1 10 11
18 0 3 3 13 10 9 10 9 1 15 0 0 9 9 11 9 0 13
11 1 3 10 9 11 13 9 13 13 1 11
10 15 3 0 3 13 7 15 1 0 13
10 16 3 1 9 13 13 13 10 9 0
21 0 9 15 9 13 10 9 16 9 13 0 3 3 10 9 7 10 0 9 13 0
22 15 3 16 3 3 3 13 3 3 13 13 3 9 11 9 7 7 9 13 9 10 15
4 13 1 0 11
13 6 9 9 3 15 3 13 3 0 7 13 9 9
11 16 3 15 13 9 13 0 13 15 3 0
7 13 0 10 11 13 10 9
18 0 3 13 3 3 13 10 9 3 13 7 3 13 0 13 9 15 9
6 13 3 10 11 13 13
19 13 3 10 9 3 10 9 9 7 13 15 3 13 7 3 15 3 13 13
13 11 3 3 0 13 3 13 3 13 15 13 10 9
30 11 3 10 11 13 7 7 13 0 3 0 7 13 7 0 0 3 3 13 0 3 13 16 3 3 13 13 1 11 0
14 6 9 15 3 13 10 9 13 7 13 7 13 10 9
11 15 3 13 3 0 15 10 0 13 10 0
12 1 0 13 11 16 0 9 13 13 10 11 13
7 1 3 9 10 15 13 15
13 16 3 10 11 13 0 13 13 10 11 1 10 9
17 9 0 6 0 13 15 0 9 7 16 15 13 13 7 15 3 15
5 0 3 1 0 13
16 3 3 3 3 3 10 9 9 13 15 7 3 13 15 13 9
8 9 0 16 15 0 13 13 13
4 13 3 3 13
14 13 0 0 3 13 10 9 9 3 13 13 1 10 0
6 6 9 13 9 0 13
13 0 13 10 11 13 9 9 9 9 3 9 10 9
10 15 3 16 15 10 9 13 13 13 15
13 7 0 3 0 10 9 13 7 0 7 10 9 15
13 13 3 3 15 3 9 7 9 7 10 15 0 9
7 15 3 0 1 15 0 13
32 3 3 9 3 0 0 9 10 9 0 0 1 10 9 13 7 15 11 13 9 9 7 13 0 7 10 15 9 15 9 13 11
10 10 3 3 10 9 0 9 3 13 13
13 3 3 3 10 10 1 11 13 9 9 3 13 13
23 11 3 13 13 7 13 1 0 0 10 13 9 13 15 13 3 9 9 13 10 9 7 9
17 11 3 16 13 16 13 0 13 7 13 9 7 13 9 13 10 0
6 0 3 3 3 3 13
9 11 3 13 10 9 13 1 10 11
6 3 13 13 1 10 11
51 6 9 15 15 9 13 9 9 0 7 7 0 13 13 9 1 11 16 9 7 0 13 0 7 0 9 7 9 0 9 7 0 3 9 13 0 3 0 15 9 13 13 0 15 3 0 13 7 9 7 9
13 15 3 0 10 9 13 0 13 16 3 0 9 13
11 16 3 15 13 13 16 3 0 1 9 13
13 0 13 10 11 3 13 11 3 3 13 10 13 13
11 3 3 13 9 1 10 11 10 11 13 0
5 11 9 11 0 13
14 15 13 13 15 7 7 10 15 9 13 15 15 9 0
14 3 3 13 3 9 0 13 13 15 3 16 15 15 13
17 0 10 9 13 10 11 7 3 0 13 9 9 13 13 1 10 11
6 13 3 15 13 11 0
52 16 3 13 1 9 7 15 15 13 1 9 15 3 0 9 3 1 0 13 3 15 13 7 7 1 9 15 13 13 16 9 15 13 0 9 9 0 7 7 0 15 15 15 3 0 13 13 13 1 9 10 15
10 3 3 3 3 13 13 0 15 15 13
9 11 3 13 7 10 0 1 11 9
18 15 3 15 13 1 11 13 15 3 3 15 13 15 7 9 13 7 9
17 13 3 15 10 9 9 1 15 13 7 13 10 9 1 15 13 13
25 13 3 10 11 13 9 13 1 10 11 15 13 13 10 9 10 11 13 15 13 1 15 13 9 13
21 0 3 10 11 10 13 1 0 10 9 3 9 13 11 10 9 0 7 13 7 0
8 13 3 11 10 1 10 11 9
16 13 3 1 0 9 13 11 7 7 11 15 3 3 1 9 13
12 10 3 3 0 7 13 3 7 13 1 9 13
15 10 3 13 15 10 9 9 13 11 10 11 10 13 11 9
4 9 3 0 0
20 15 13 7 13 15 3 9 1 9 13 15 3 13 10 11 9 1 9 3 13
5 0 3 0 13 13
20 1 3 3 0 9 9 0 13 7 13 10 0 1 11 7 7 11 9 13 0
9 0 3 3 10 11 9 10 9 13
9 0 3 9 1 15 9 13 10 0
5 13 3 15 3 0
25 13 3 0 7 13 15 10 0 16 15 13 1 13 10 9 9 3 13 13 10 9 10 9 10 9
28 13 3 15 10 9 7 0 13 0 16 3 13 1 10 9 9 13 13 0 3 9 13 15 13 10 9 3 13
13 13 3 13 3 10 0 3 3 15 13 3 10 15
10 10 3 15 0 10 3 13 0 13 13
6 0 3 3 0 3 13
12 3 3 1 0 10 9 3 13 0 13 10 11
5 13 3 13 1 11
23 10 3 11 9 13 11 7 13 0 10 9 13 1 11 16 10 0 13 9 3 13 10 11
21 13 3 10 0 1 10 11 13 10 11 16 3 15 13 9 15 7 13 1 10 15
25 15 3 13 16 16 1 15 13 1 10 9 13 10 11 9 3 13 10 9 10 11 0 15 9 13
10 13 3 12 9 0 13 7 9 0 0
5 13 3 15 9 13
3 13 3 0
5 11 15 13 13 9
9 0 3 13 10 9 13 15 3 13
44 0 13 10 11 13 10 11 13 3 13 0 7 13 9 13 7 9 10 9 3 0 13 9 0 13 3 13 1 10 11 15 13 10 0 15 3 0 13 3 3 3 10 15 9
11 10 3 9 0 10 11 15 3 13 1 11
28 13 3 10 11 1 10 11 13 1 10 11 16 11 13 9 9 3 3 0 3 3 0 7 7 0 7 1 11
6 9 3 13 0 7 9
14 15 3 1 0 10 9 13 13 1 15 10 9 1 15
17 7 15 0 13 0 3 13 0 1 15 9 0 1 10 9 10 9
9 0 3 3 0 15 10 13 13 13
18 3 3 13 3 13 11 9 0 7 7 0 3 0 11 7 3 0 13
7 13 3 12 9 0 15 13
5 15 3 13 15 0
19 15 1 9 10 9 9 13 9 0 7 0 3 13 15 1 10 9 10 9
11 1 3 12 9 12 15 0 13 1 10 9
8 13 3 0 3 0 9 0 13
12 10 3 3 11 16 0 13 0 13 13 1 11
34 10 3 11 16 15 13 1 11 7 13 10 1 10 11 13 0 3 0 11 13 13 3 12 9 0 3 3 9 9 7 7 10 0 9
21 13 3 10 11 10 7 11 1 10 11 7 10 0 9 7 10 0 13 9 1 11
18 16 3 13 1 11 13 10 9 1 11 16 3 9 9 1 10 11 13
9 7 3 3 13 0 10 9 0 13
4 9 0 13 13
13 13 11 10 1 10 9 9 1 9 0 13 15 13
35 15 3 0 15 13 13 10 9 13 10 9 0 10 9 15 9 13 11 0 13 1 0 13 10 9 1 0 3 3 9 13 3 3 10 9
17 13 3 10 11 13 15 10 11 16 10 9 15 10 0 11 13 13
8 13 3 15 15 13 0 13 13
3 15 3 13
8 15 3 3 0 10 9 15 13
12 3 15 13 11 15 13 7 13 3 3 15 13
3 15 0 13
4 0 13 10 11
20 15 3 13 0 16 9 13 13 1 11 9 9 13 10 0 15 10 13 15 9
25 16 3 13 3 3 13 10 1 10 9 1 10 9 13 3 3 13 7 9 7 0 7 10 9 13
19 15 3 16 13 1 10 11 10 9 1 10 11 1 13 13 7 13 9 12
9 11 3 3 13 10 9 10 11 13
25 3 3 13 15 10 9 10 9 13 13 7 10 9 13 3 7 11 13 13 7 10 9 10 11 13
6 13 3 0 0 13 9
17 13 3 3 10 13 10 9 13 1 11 1 11 13 13 11 1 9
18 10 3 11 13 10 11 13 13 3 3 3 13 3 13 3 13 10 9
27 16 3 13 3 13 1 11 13 15 15 3 15 16 3 13 1 11 13 11 13 15 10 9 13 1 10 9
10 10 3 9 13 3 3 0 15 13 9
14 0 3 10 11 13 9 13 0 10 15 9 10 1 11
13 3 3 0 15 13 10 11 0 1 15 13 3 13
8 11 3 3 0 13 13 10 9
9 11 3 13 10 0 9 15 0 13
16 13 3 1 10 9 13 10 7 15 9 7 10 1 10 11 13
25 11 3 10 9 0 3 3 13 9 9 10 9 13 13 10 7 9 15 15 13 11 7 10 9 15
12 16 3 3 13 0 13 13 16 9 10 9 13
9 3 3 3 3 13 13 13 13 0
8 13 3 10 9 10 0 13 0
14 10 3 9 13 0 0 3 13 15 1 10 0 10 9
7 0 3 3 3 13 10 9
28 13 3 3 13 12 7 15 13 1 11 1 10 9 10 1 10 11 13 13 3 13 13 10 1 10 9 13 9
18 7 0 3 9 13 10 9 9 13 10 11 16 3 0 15 10 0 13
11 3 3 3 1 10 0 11 10 0 0 13
32 15 3 13 10 9 15 3 13 9 1 10 9 10 13 1 11 0 3 0 13 13 10 9 13 0 1 0 9 13 3 13 0
9 11 3 3 0 16 3 13 13 13
6 0 3 10 15 15 13
8 9 3 3 9 13 1 10 9
23 11 3 10 0 16 10 9 13 9 1 0 10 9 13 0 13 0 0 1 11 9 9 13
12 10 3 11 11 3 10 11 3 13 13 7 13
14 11 3 10 11 13 10 9 3 1 9 13 7 1 9
15 11 3 13 9 9 15 9 7 13 0 15 0 9 3 13
9 0 3 0 13 10 9 13 13 15
17 16 3 15 15 3 13 7 15 0 13 3 13 9 10 11 13 0
11 15 3 15 3 13 9 16 15 3 13 13
5 7 13 0 9 13
3 7 15 13
11 1 0 10 9 7 10 9 13 13 11 0
25 16 3 3 13 15 13 15 13 9 15 3 0 13 7 3 13 0 16 3 15 0 1 15 9 13
9 9 3 15 13 3 13 15 10 9
16 15 3 0 7 15 15 3 13 13 7 0 1 0 13 9 0
6 0 3 13 13 10 11
11 3 3 9 13 12 0 9 13 13 3 0
18 13 3 15 0 9 10 10 13 9 0 13 13 13 15 13 3 13 13
16 0 3 13 15 10 9 13 1 9 10 9 13 10 9 13 13
14 15 3 16 13 11 3 13 11 7 1 0 3 13 11
9 15 3 3 0 13 11 7 11 13
18 10 3 11 13 7 10 0 13 9 13 9 9 10 11 3 13 10 0
12 10 3 3 11 3 13 13 7 3 0 0 7
17 10 3 11 13 10 9 15 0 3 7 13 1 9 0 13 10 9
53 3 3 3 13 16 10 7 11 13 7 10 0 13 10 9 13 9 10 0 11 10 11 0 7 13 7 3 13 1 11 13 13 9 9 13 1 9 7 10 1 11 9 13 1 15 9 13 13 7 13 15 10 13
5 13 3 10 9 0
12 13 3 1 11 13 9 0 10 9 1 11 9
14 13 3 3 0 9 1 9 7 9 7 0 13 1 11
26 3 3 15 11 9 0 13 1 10 11 9 11 10 1 11 13 13 10 11 9 15 13 9 0 11 13
16 15 3 13 0 1 11 13 13 10 9 16 13 1 15 13 9
6 10 3 11 15 13 13
14 13 3 11 10 9 15 3 1 11 13 13 1 10 11
10 13 7 3 1 11 11 7 13 10 11
19 1 11 10 9 9 13 13 1 15 16 15 10 0 3 13 0 13 1 11
4 0 3 0 13
6 9 3 0 0 13 0
21 9 3 9 7 7 9 13 1 10 0 11 15 13 13 10 9 11 13 11 0 0
15 0 3 0 11 10 9 9 0 13 16 1 10 13 13 13
27 16 3 3 3 13 15 1 15 3 13 13 13 3 10 0 9 7 13 13 7 3 0 7 7 10 9 13
32 10 3 3 9 13 11 3 10 0 0 1 9 10 0 0 13 15 3 1 15 3 13 10 11 9 11 3 7 10 11 9 15
14 13 3 11 3 15 9 9 11 7 11 7 11 7 11
9 0 3 11 10 9 13 0 10 9
18 13 3 0 10 9 10 13 13 11 10 0 9 7 13 0 10 9 11
14 3 3 16 0 13 0 9 13 11 7 13 9 1 0
11 10 3 15 0 13 13 13 1 11 0 9
19 13 3 11 7 13 11 10 11 9 9 15 13 11 10 9 9 13 1 11
8 13 3 10 9 13 13 1 11
11 1 3 10 15 9 13 1 0 15 15 0
10 1 3 10 9 15 9 13 9 15 13
13 16 3 13 13 1 11 7 13 1 11 13 3 11
18 3 3 15 0 9 13 10 11 7 13 0 9 0 13 15 9 13 11
15 13 3 3 10 11 10 11 9 1 10 11 11 13 10 9
24 15 3 1 9 13 3 0 13 13 0 9 1 15 9 0 9 13 7 9 7 15 7 9 15
10 13 3 1 9 10 11 13 1 15 0
5 10 3 13 13 0
13 9 9 9 13 1 0 9 7 9 0 3 0 15
9 3 3 10 0 15 15 13 10 11
8 3 3 15 0 0 7 13 13
28 7 3 10 0 0 13 15 7 10 1 10 9 1 10 0 13 9 1 10 7 9 15 13 0 9 7 9 0
12 9 3 13 13 1 10 9 7 9 1 10 9
4 3 0 13 13
19 13 3 15 13 3 15 13 9 3 0 0 9 13 7 9 0 7 0 13
15 13 3 13 0 1 10 9 10 9 15 13 1 10 9 13
22 9 3 13 13 10 11 0 13 9 10 1 10 9 0 7 13 15 15 15 13 7 0
8 9 3 13 9 15 15 0 13
8 15 12 9 9 10 0 9 13
10 9 3 0 13 0 0 3 0 13 0
6 0 3 9 9 0 13
12 13 3 0 10 9 13 3 10 11 9 1 13
44 7 1 3 9 3 3 0 7 3 0 7 9 0 0 13 15 9 13 1 7 0 13 0 7 9 7 7 0 15 7 9 13 13 15 7 9 15 1 3 15 13 9 13 13
10 13 3 10 11 15 13 3 15 15 13
4 11 3 0 13
4 11 3 13 0
5 3 3 1 0 13
28 16 3 10 0 9 13 10 9 7 13 1 10 13 13 10 11 10 11 15 9 1 9 10 9 9 13 1 9
14 0 3 15 3 13 10 13 13 3 9 13 1 10 11
9 13 3 3 12 9 13 13 10 9
15 15 3 13 10 0 9 15 10 11 13 13 1 10 9 13
9 6 9 0 13 1 11 1 13 9
14 15 3 9 0 13 0 13 15 1 9 12 9 9 13
9 10 3 11 0 13 13 1 10 9
12 13 3 3 3 13 13 13 10 11 13 10 9
13 0 3 15 3 0 9 13 13 9 12 7 12 9
12 11 3 13 15 13 15 13 7 13 10 9 1
14 3 3 10 11 13 1 12 9 13 16 15 13 15 13
20 13 3 10 11 13 10 9 13 10 11 16 15 12 7 9 13 7 10 9 13
9 9 13 15 10 9 16 3 13 13
35 10 7 3 11 13 10 9 10 9 13 1 0 9 7 10 11 13 10 3 1 10 11 7 15 13 1 0 3 13 1 10 9 10 1 9
7 13 3 1 10 9 0 3
27 13 3 1 10 11 10 11 9 1 15 9 7 13 15 13 15 9 7 3 13 10 9 7 9 0 1 15
20 13 3 1 10 11 7 3 13 1 9 10 0 9 12 13 13 12 9 3 12
13 1 3 10 0 9 0 7 9 13 7 0 9 13
17 0 3 13 7 1 10 11 9 13 12 13 9 9 3 12 7 0
12 9 3 11 7 10 11 13 9 0 15 9 11
18 1 3 10 11 9 3 13 9 12 9 3 12 7 0 7 9 1 15
12 9 3 0 12 1 0 13 15 15 9 13 13
22 0 3 11 3 3 0 7 7 0 10 0 13 3 10 0 13 9 7 1 10 0 13
6 0 10 15 9 13 12
11 9 3 3 9 0 13 1 11 1 11 13
35 16 3 3 13 10 9 10 0 10 9 7 10 9 13 12 9 3 0 3 13 0 1 11 9 13 1 10 9 10 0 13 12 9 13 12
13 12 3 7 12 9 1 9 0 13 13 9 3 12
19 3 10 0 11 13 1 11 10 0 13 12 9 10 9 10 1 9 3 13
12 16 3 15 10 0 0 3 13 15 3 0 13
10 10 3 1 11 1 11 9 13 13 0
19 7 3 13 9 13 10 15 1 9 10 0 1 11 0 3 0 9 13 12
40 16 11 10 11 11 3 10 9 9 13 9 9 10 15 9 0 13 11 7 11 9 13 10 3 0 1 0 13 0 1 9 12 15 0 7 3 3 3 1 15
9 10 3 3 9 10 11 9 13 0
19 1 10 0 9 10 9 13 10 11 9 15 13 0 7 0 13 0 10 9
6 13 9 0 13 13 9
6 15 9 13 9 3 13
10 0 3 16 9 13 3 0 13 13 9
12 3 3 13 10 9 13 10 9 1 15 3 13
18 3 3 15 13 13 13 9 10 1 11 13 9 1 9 10 3 11 13
17 3 3 0 0 13 1 0 10 0 0 0 1 9 13 13 1 11
17 0 3 15 1 0 13 15 0 13 9 0 15 7 3 0 13 13
13 3 3 9 13 1 10 9 13 3 10 9 10 9
24 13 3 15 10 0 10 9 0 10 9 9 9 15 13 9 1 10 9 10 9 13 15 0 13
15 13 3 13 3 3 10 0 13 13 9 1 10 11 0 13
21 7 10 9 9 13 1 10 0 10 9 16 3 1 9 9 13 9 0 7 7 0
27 13 3 3 0 0 9 1 10 9 10 11 10 0 1 11 10 9 1 9 15 13 10 0 0 13 10 0
8 10 3 3 12 10 9 9 13
12 0 9 13 3 1 11 10 11 10 11 10 11
7 0 3 9 1 0 9 13
10 11 13 15 0 11 13 13 15 0 9
27 11 3 3 13 10 11 16 3 0 3 13 10 13 7 3 0 10 0 9 13 15 11 9 1 11 10 11
8 0 3 9 13 3 0 1 0
17 1 0 3 10 11 10 11 13 13 0 1 0 7 13 1 10 9
10 10 3 0 13 0 1 9 13 1 11
28 7 15 0 13 1 11 13 15 15 13 10 0 0 15 7 13 10 0 0 7 3 3 11 11 9 7 7 9
16 13 3 1 0 3 13 15 1 9 13 13 9 3 9 13 0
69 11 13 7 13 0 1 10 11 9 9 9 13 0 7 13 9 16 15 1 10 0 0 9 13 1 10 0 3 13 9 7 13 3 13 13 7 7 13 10 11 11 10 1 11 13 3 10 9 15 1 10 9 13 1 9 10 9 13 10 1 11 10 3 13 3 3 3 0 13
34 15 3 9 3 13 7 13 9 0 3 3 10 7 9 13 10 9 0 10 7 0 7 13 15 0 9 13 10 9 0 10 3 15 13
31 3 3 3 10 0 13 0 10 9 1 11 13 13 10 11 9 16 13 9 9 7 0 9 7 0 13 13 15 10 11 13
10 10 3 10 9 0 13 3 10 10 9
6 13 3 0 1 9 9
9 15 3 3 13 1 11 10 9 13
9 10 3 9 13 0 13 1 11 9
19 9 3 15 13 13 0 9 13 12 7 9 7 10 9 10 15 11 9 0
8 15 16 13 9 10 9 13 0
16 13 10 11 10 9 7 0 13 0 10 9 13 10 9 10 9
8 10 3 13 15 1 10 9 13
22 10 3 3 0 9 1 11 3 13 7 11 13 9 10 11 11 1 10 11 10 1 11
25 3 3 0 0 9 13 13 1 10 11 9 10 9 13 9 11 10 11 3 1 9 13 7 1 9
23 10 13 1 10 11 9 10 10 9 9 0 13 7 3 1 0 13 7 15 13 1 12 9
9 10 3 13 13 3 13 3 1 11
9 7 15 15 3 3 13 9 10 0
22 7 3 9 13 13 10 7 9 9 7 0 3 13 13 7 3 9 0 13 1 10 11
10 13 3 1 10 9 10 9 10 9 13
9 0 3 16 13 15 15 10 9 13
19 13 3 1 9 10 9 1 15 13 10 0 16 1 12 9 13 1 10 11
42 3 3 13 1 11 10 1 10 11 13 3 0 1 9 12 13 3 3 0 3 0 7 7 9 1 10 0 13 3 10 1 11 7 7 11 15 0 9 13 13 0 9
21 1 0 3 3 10 0 9 13 11 10 9 13 10 11 1 10 11 11 13 10 9
5 3 3 0 9 13
31 1 3 15 12 9 13 11 7 9 9 15 3 3 9 13 10 11 13 7 11 11 9 3 13 0 3 10 3 3 13 13
6 0 10 9 13 1 9
7 13 3 10 11 10 9 13
28 3 3 0 13 0 0 13 10 11 9 11 7 11 7 11 7 11 13 10 9 13 3 0 9 9 0 1 11
9 0 3 3 0 7 0 9 13 13
15 0 3 13 15 13 10 11 0 10 15 9 11 10 11 9
24 11 3 0 13 0 3 9 13 1 11 13 10 0 9 1 16 0 7 7 11 10 0 15 13
26 0 3 9 3 13 7 13 1 0 10 9 10 0 11 10 11 0 13 10 11 13 0 13 1 10 9
17 16 3 10 9 0 3 3 13 13 3 13 9 15 0 10 11 13
16 16 3 15 13 13 13 1 11 10 0 13 13 13 11 10 11
4 10 3 0 13
20 13 3 10 11 10 11 9 15 13 1 0 10 9 7 15 13 3 1 10 0
26 13 3 10 11 10 11 3 3 0 13 13 3 0 13 11 15 10 7 9 15 11 13 7 10 9 11
15 16 3 15 10 9 13 9 7 7 9 11 13 13 10 11
9 10 3 0 13 3 3 13 10 11
6 10 3 9 13 0 11
8 9 3 11 13 13 11 10 9
26 10 7 3 15 10 0 13 10 11 7 3 3 10 9 15 0 9 13 10 3 11 3 13 10 3 11
12 11 3 9 3 10 11 13 10 3 0 9 11
6 0 3 1 11 15 13
19 9 3 10 9 16 3 3 10 0 13 10 0 7 10 0 13 1 15 9
6 3 3 0 13 10 0
17 1 3 9 7 7 9 10 9 13 0 10 0 13 1 10 15 9
9 0 3 10 9 1 10 15 9 13
13 3 3 9 15 13 13 1 10 9 7 9 7 9
14 0 3 15 13 1 10 11 9 11 10 9 13 13 9
7 0 3 3 10 0 11 13
35 10 3 3 0 11 13 10 0 10 9 7 10 9 1 0 13 13 15 3 0 13 9 16 3 15 10 0 13 9 3 9 10 0 11 13
23 16 3 3 10 0 9 0 13 3 15 1 10 15 9 13 10 9 13 7 13 0 1 0
7 12 7 3 9 1 12 13
9 3 3 3 10 9 13 1 10 9
9 1 10 9 3 13 10 11 13 0
11 10 3 11 13 9 13 1 10 11 10 9
22 10 3 3 0 13 10 11 1 10 11 9 13 11 7 1 15 15 0 0 15 0 13
8 0 3 13 13 1 9 10 11
13 10 3 3 9 7 10 9 15 13 9 10 9 0
8 0 3 3 13 7 10 9 15
6 10 3 0 0 3 13
4 0 1 9 13
9 13 3 9 10 9 13 10 9 13
16 0 13 3 10 9 10 9 15 3 13 3 10 11 0 1 9
6 13 3 15 9 13 9
6 0 1 10 11 9 13
13 11 3 16 13 13 11 7 10 0 11 3 0 13
14 3 3 15 0 13 1 10 11 10 11 3 1 0 9
8 0 3 13 0 10 9 13 13
8 12 3 10 11 9 10 9 13
21 13 3 10 9 7 3 13 13 10 7 11 7 10 11 7 10 9 15 13 10 9
12 10 3 0 0 13 1 10 9 15 13 15 0
6 13 3 10 11 10 9
18 16 3 13 1 10 9 13 3 15 13 13 1 10 0 10 9 3 13
14 10 3 9 13 1 10 9 16 3 10 9 15 13 13
6 3 3 0 9 13 3
3 15 3 13
8 6 9 7 3 9 13 7 0
16 15 3 3 10 9 15 13 13 7 7 3 3 13 1 0 0
23 0 3 1 0 11 7 10 12 0 10 13 1 11 13 13 9 1 11 9 13 13 1 9
8 13 3 15 0 7 7 11 13
8 13 3 1 10 9 13 15 0
7 16 3 3 13 13 15 13
13 10 3 9 1 15 0 13 13 13 13 10 9 13
10 0 3 3 13 1 10 15 9 0 13
31 11 3 13 13 9 7 9 1 0 13 1 15 11 9 3 13 1 15 13 13 7 13 10 9 10 0 7 11 13 9 13
7 13 3 15 0 1 10 9
14 0 3 3 9 13 9 3 7 9 1 0 13 9 13
9 0 3 13 1 11 1 13 10 9
4 3 3 0 13
11 13 3 0 10 0 13 3 10 9 10 0
11 1 15 3 3 3 0 0 0 15 13 13
26 3 3 1 10 11 13 10 0 10 9 10 7 9 10 0 3 13 7 0 13 10 9 13 3 0 13
21 0 3 0 1 10 11 13 9 3 7 1 9 13 7 3 1 0 10 9 10 0
6 0 3 16 3 11 13
12 0 3 7 0 16 1 9 9 13 1 11 13
15 13 3 10 9 0 3 3 0 13 13 0 9 13 1 9
8 9 3 10 9 13 1 10 11
13 0 3 13 10 9 13 0 10 9 3 10 9 13
10 13 7 3 10 9 10 0 7 0 13
7 3 3 0 13 12 15 13
15 10 3 0 0 9 10 0 13 1 10 11 13 3 10 9
12 13 3 3 0 12 9 1 10 9 10 9 13
6 9 3 13 15 0 13
11 10 3 9 15 1 15 13 13 1 10 9
24 15 3 3 3 1 15 13 13 13 1 9 13 9 1 10 9 1 3 10 9 10 1 9 13
9 7 10 9 10 0 13 13 0 0
14 15 3 0 9 13 0 13 1 10 0 10 1 10 9
4 13 3 15 0
16 9 9 7 9 13 9 0 9 1 9 9 1 0 0 13 9
6 15 9 0 11 0 13
27 13 3 3 1 12 0 7 3 10 9 16 13 9 0 16 3 0 13 3 0 10 15 13 13 10 0 0
6 13 3 9 0 0 13
10 13 3 0 16 13 3 13 3 9 13
7 13 3 0 0 15 13 13
5 0 3 3 0 13
10 0 3 1 0 1 9 13 13 13 0
12 10 3 11 1 15 3 0 3 13 15 13 9
9 13 3 10 0 13 10 9 9 13
11 7 0 3 1 15 3 13 3 13 10 9
5 15 13 0 3 13
8 7 3 3 3 0 13 10 9
7 0 13 13 3 3 13 15
10 15 15 13 13 15 13 13 15 10 9
8 11 13 13 9 11 7 7 11
12 0 9 13 13 15 9 13 10 9 13 9 13
13 3 13 13 9 13 1 10 9 15 13 3 13 0
24 13 3 10 0 1 10 9 10 9 7 3 13 1 10 0 3 10 0 13 10 3 9 15 13
4 10 3 9 13
20 9 3 9 7 0 13 7 9 0 13 13 1 0 3 0 13 9 0 0 13
21 13 3 15 9 13 0 9 1 10 11 3 3 13 11 3 3 10 0 0 0 9
6 13 3 0 3 0 13
14 10 3 9 10 13 1 0 1 10 9 13 1 9 0
10 1 0 3 10 9 10 0 13 1 11
16 10 3 11 15 13 11 7 7 11 9 13 7 15 13 0 13
10 10 3 11 15 0 13 7 9 0 9
14 13 3 10 0 0 9 15 13 13 0 3 0 13 13
15 13 3 3 16 9 13 3 9 3 1 9 0 3 1 11
20 15 3 1 0 13 13 1 15 13 9 0 10 11 7 10 11 0 7 10 11
18 13 3 1 0 10 0 15 7 13 13 7 9 1 10 9 0 13 13
27 0 3 3 10 9 7 1 15 9 0 13 10 7 0 7 9 13 1 11 13 7 7 13 1 15 10 9
14 10 3 1 0 9 7 13 7 9 13 13 1 10 0
40 3 3 13 0 13 15 3 9 13 7 3 3 10 9 0 10 7 11 7 10 11 13 15 7 15 13 7 7 13 10 15 9 1 10 0 15 11 3 13 9
21 13 3 1 0 10 9 9 7 15 7 9 0 0 13 9 13 0 10 9 12 9
12 3 3 13 10 9 9 3 15 10 3 0 9
8 13 3 3 10 0 10 0 9
6 13 3 15 3 0 9
7 13 3 10 0 13 10 0
7 15 3 13 9 16 3 13
29 15 3 3 9 13 10 9 1 10 9 13 15 13 16 3 13 15 3 0 13 13 3 7 10 13 15 9 13 13
10 1 0 10 0 1 11 13 13 10 9
37 0 3 3 13 1 10 9 13 9 12 10 9 0 15 13 1 10 0 7 13 1 11 10 9 0 3 15 9 13 13 1 10 9 13 16 15 13
24 3 13 3 0 10 9 15 13 13 9 13 10 9 7 15 13 9 7 7 1 10 9 9 13
8 10 3 9 10 13 1 0 13
7 9 3 3 12 9 13 0
17 12 3 3 7 0 0 12 3 16 15 3 13 13 9 13 3 3
8 7 0 9 13 15 1 10 9
7 0 3 15 13 7 3 13
17 0 3 3 16 15 15 1 9 13 13 1 10 9 13 1 10 9
5 0 3 3 0 13
15 15 3 9 13 13 10 0 16 13 1 15 13 0 0 13
9 13 3 3 1 0 7 7 9 0
14 13 3 3 1 0 12 0 10 13 15 1 10 11 13
17 3 0 3 13 15 10 0 9 13 10 12 0 13 0 3 10 9
10 13 3 3 0 10 12 7 13 9 0
8 13 3 1 10 11 13 10 9
36 13 3 10 9 10 1 11 13 9 0 15 13 0 0 1 0 13 3 10 9 0 13 7 13 10 9 10 9 13 0 15 3 13 10 15 9
13 0 3 3 10 9 0 15 13 13 10 10 9 9
8 10 3 9 13 15 1 10 0
14 13 3 3 1 15 10 10 0 9 9 0 10 0 0
11 13 3 1 10 0 9 16 3 9 3 13
31 13 3 0 9 13 3 0 0 10 9 10 0 7 0 16 10 3 0 9 15 10 0 10 9 10 0 13 15 3 0 13
23 0 3 3 7 9 10 9 1 0 1 9 10 0 9 3 3 1 15 13 0 3 1 15
14 10 3 9 10 1 9 1 0 13 9 1 15 13 13
16 3 3 0 13 3 10 1 10 9 13 13 10 9 13 10 9
18 0 16 13 13 10 0 10 3 11 9 13 0 15 3 1 10 9 13
14 12 3 9 3 13 13 16 0 13 13 13 1 9 0
11 1 9 3 13 15 1 0 9 13 0 13
44 13 3 0 10 1 10 9 1 10 11 13 7 0 1 10 11 1 15 7 7 10 9 9 13 0 16 7 9 9 15 13 13 1 10 0 7 16 0 13 9 15 13 1 0
29 3 7 1 0 13 15 10 9 13 0 7 7 0 13 15 1 0 15 0 3 13 0 3 3 11 13 1 11 13
16 13 3 10 11 1 10 0 9 10 9 15 13 3 0 10 9
6 13 3 13 1 10 9
5 13 3 10 11 13
8 9 9 13 0 15 3 13 3
30 13 3 0 9 9 9 13 15 10 3 7 13 0 13 10 11 0 1 10 9 13 7 3 13 0 9 0 13 10 9
14 15 16 1 15 13 13 15 3 7 10 9 15 13 13
14 9 3 13 13 16 13 3 3 10 0 15 9 7 9
7 3 3 15 3 0 13 13
12 16 3 0 13 13 3 13 15 1 15 13 13
29 0 3 0 1 0 7 11 13 7 15 1 10 9 16 0 7 9 7 0 9 13 15 1 10 11 13 15 3 13
4 15 3 0 13
5 0 3 11 13 0
49 3 3 10 7 9 1 13 10 9 7 10 9 0 1 10 9 7 9 9 1 9 13 7 9 15 0 9 16 3 15 6 0 9 13 9 1 10 9 13 13 15 7 0 13 15 1 9 7 0
26 16 3 3 0 3 13 15 13 0 16 13 10 9 0 0 9 13 1 15 0 3 3 10 0 13 13
19 3 3 0 9 0 13 7 13 0 0 1 10 11 16 13 13 1 10 9
18 16 3 15 0 13 3 3 15 13 3 1 15 9 0 13 3 3 3
6 0 3 13 9 9 0
9 13 9 7 0 9 13 13 10 9
9 11 3 13 0 10 9 13 9 0
6 0 9 3 15 13 13
16 13 11 10 11 9 3 13 1 11 3 10 3 9 7 7 9
11 1 3 15 0 10 9 7 1 0 9 13
6 13 3 1 11 1 9
10 13 3 15 3 10 11 13 0 10 9
6 11 15 15 13 0 13
3 13 3 9
5 1 3 13 9 0
30 0 13 10 11 13 3 10 9 15 10 3 0 13 9 1 11 13 0 13 7 1 10 0 3 10 10 11 7 13 3
4 9 1 9 13
5 13 3 9 0 0
5 0 3 3 9 13
13 0 3 3 13 0 15 1 0 11 13 7 0 11
16 3 3 10 11 13 16 13 3 3 10 0 13 13 0 10 11
14 13 3 3 0 13 1 9 13 10 13 11 13 9 13
21 16 3 13 10 9 3 13 15 0 12 1 10 9 1 15 13 10 11 13 10 9
22 10 3 11 13 7 15 15 1 0 13 7 13 15 9 10 9 1 13 13 13 15 12
13 15 3 3 13 1 9 10 0 15 13 10 9 13
23 16 3 13 13 10 11 10 13 10 9 0 9 13 10 9 7 10 13 0 9 15 13 13
9 13 3 13 10 0 0 3 10 0
41 13 3 3 10 13 10 9 7 13 3 13 1 10 9 15 13 13 7 3 10 0 13 16 3 13 1 10 13 16 15 3 15 9 13 13 3 13 15 10 9 13
9 13 3 1 10 11 9 11 0 13
11 10 11 3 15 0 13 13 1 0 10 9
32 13 3 16 15 13 7 10 0 13 10 9 13 13 13 1 10 0 15 13 13 1 9 13 16 16 13 1 9 13 15 13 13
21 13 3 7 13 15 16 3 13 13 13 7 13 1 10 13 16 15 13 15 0 13
6 15 3 3 13 13 0
20 11 3 1 0 10 9 13 7 15 13 0 10 9 1 10 9 9 11 9 13
5 10 3 9 0 13
20 0 0 9 15 15 9 13 11 9 9 0 11 0 7 9 9 3 3 3 9
6 10 3 3 9 0 13
9 13 3 10 11 0 3 15 9 13
4 0 3 0 13
10 10 3 11 1 9 3 13 0 10 9
14 16 3 13 1 9 11 10 11 9 0 3 13 11 0
11 11 3 10 13 1 10 11 13 1 10 9
30 13 3 1 9 13 3 7 13 10 9 13 7 7 13 10 9 1 10 1 11 9 7 13 3 3 15 13 10 9 13
15 13 3 13 16 15 10 9 10 0 7 7 0 13 9 0
11 13 3 10 9 7 13 9 15 13 10 9
14 13 3 10 9 1 10 11 13 0 13 10 9 10 11
28 15 3 15 15 13 11 13 13 7 15 1 15 15 9 13 3 0 7 7 10 15 0 13 15 3 1 11 13
11 15 3 11 13 13 7 7 13 11 15 13
29 13 3 15 1 9 1 11 9 9 1 10 9 9 1 0 7 13 13 10 11 13 7 13 1 15 13 9 10 9
6 13 7 3 7 13 0
10 15 3 15 13 9 9 13 15 3 13
17 9 3 15 13 16 0 0 13 16 1 0 10 9 11 10 9 13
33 0 3 16 3 13 10 11 0 3 15 13 10 9 15 9 13 11 13 3 3 1 10 9 9 13 1 10 0 13 15 10 0 9
11 15 3 3 3 1 9 13 9 10 0 13
15 15 3 13 10 9 13 15 15 3 10 7 0 7 10 0
11 0 3 15 13 10 9 6 0 7 0 9
35 15 3 10 0 3 3 9 0 13 16 15 13 13 11 3 7 3 3 3 13 13 0 13 7 13 15 9 10 0 3 13 9 1 10 9
9 3 13 7 13 1 10 0 13 11
6 13 15 0 3 3 13
7 11 3 1 11 13 13 0
25 11 3 15 13 10 0 13 9 0 3 3 0 3 15 13 9 3 15 13 9 10 0 13 1 0
10 11 3 0 13 15 10 9 0 9 13
12 10 3 0 10 9 3 3 13 1 9 15 0
12 7 11 3 13 1 3 15 3 9 0 9 11
10 15 13 10 9 0 13 10 1 9 9
17 3 3 10 9 10 1 11 9 9 13 13 0 13 7 13 10 9
10 7 3 1 3 11 3 13 10 9 13
8 13 3 1 9 13 15 1 11
5 7 13 3 10 9
4 13 3 0 13
27 7 0 15 10 9 13 15 7 0 3 3 3 3 9 13 9 0 7 9 13 7 1 11 10 0 0 13
19 3 3 0 3 10 3 13 10 9 13 15 0 1 9 11 3 13 13 15
21 9 3 10 0 9 13 3 3 15 13 13 1 11 15 3 0 10 1 9 9 13
8 0 3 9 15 15 13 1 0
7 13 3 3 0 3 1 9
16 3 11 11 3 10 0 9 9 0 11 3 10 11 10 11 9
11 3 3 16 3 10 9 13 13 3 13 13
23 16 3 3 13 10 11 3 15 13 13 10 9 10 0 10 11 1 10 15 9 13 10 9
9 11 3 13 11 7 13 15 0 13
8 0 3 3 13 15 13 13 13
5 11 3 3 13 11
49 9 3 11 16 13 11 13 13 1 7 0 7 9 10 3 9 13 10 9 16 0 13 10 0 11 0 3 13 15 16 13 0 9 15 9 13 3 13 16 0 3 3 13 13 13 15 13 10 0
6 3 3 13 13 10 9
6 6 11 13 15 0 13
14 13 3 0 13 12 10 9 9 13 15 1 3 3 13
17 13 3 0 13 13 1 9 11 10 0 15 10 11 13 9 3 0
14 13 11 9 10 15 15 15 11 13 0 1 15 13 9
8 3 3 3 15 0 13 13 3
9 3 3 1 10 15 9 0 15 13
8 13 16 1 0 15 1 9 13
4 13 1 0 11
18 9 15 13 9 15 13 9 1 15 15 15 7 0 7 0 13 0 13
18 7 16 3 15 0 15 15 13 13 10 15 9 13 15 1 15 13 13
20 9 3 15 3 13 10 9 16 15 0 7 10 15 9 0 13 1 9 10 15
22 16 3 3 15 0 13 3 15 10 13 13 6 9 13 15 9 13 15 1 9 0 13
9 15 3 3 13 1 11 15 9 13
28 3 3 3 9 13 15 13 1 11 16 15 0 7 15 13 1 10 0 7 10 11 9 0 10 0 13 0 13
30 0 3 1 9 10 15 13 9 13 10 0 3 3 0 13 15 13 9 13 1 11 16 3 15 11 9 10 0 0 13
5 11 3 13 0 13
38 1 15 3 10 9 7 1 10 11 1 9 13 7 11 10 1 10 9 13 11 1 9 13 7 11 13 1 11 13 1 9 1 0 15 10 9 13 0
19 13 10 0 11 0 13 9 9 0 13 0 11 9 9 0 1 10 11 13
12 13 3 0 10 11 9 13 1 10 11 13 15
9 9 3 3 1 3 13 13 0 9
13 10 3 9 10 9 13 10 9 15 13 11 10 11
14 0 3 0 13 13 10 9 10 11 13 10 9 10 9
15 9 9 9 15 13 15 10 0 15 13 13 7 9 7 9
4 13 9 1 0
21 15 3 13 10 0 10 9 13 10 9 7 3 16 0 10 9 13 0 3 9 13
10 15 3 3 1 15 13 3 13 13 0
14 15 3 0 13 13 15 13 13 1 10 9 13 9 0
4 9 3 0 13
9 0 3 7 0 13 10 0 13 9
9 11 3 10 9 10 9 9 13 11
24 13 3 0 10 11 13 3 15 9 9 3 9 10 3 0 3 0 7 3 9 0 13 1 0
15 13 10 11 9 13 0 7 9 7 9 13 1 15 3 13
15 15 3 13 13 3 15 13 13 13 7 10 9 7 0 11
6 13 1 0 10 9 15
19 6 9 0 3 15 13 13 7 0 7 10 0 15 7 3 15 3 15 13
10 3 3 15 13 13 10 15 9 0 13
23 16 7 3 13 9 9 0 15 13 7 0 16 15 0 15 3 13 1 0 3 13 0 9
6 15 15 10 9 15 13
12 15 3 15 13 16 15 9 3 3 15 13 1
10 0 13 7 3 13 10 9 3 7 9
16 9 3 3 9 0 13 0 10 9 13 10 9 7 0 0 13
8 3 3 16 13 10 9 13 13
7 1 3 10 9 0 0 13
23 16 13 1 10 11 10 11 1 10 9 13 10 11 1 15 13 10 9 13 13 0 10 11
17 13 3 3 10 0 11 9 13 11 13 13 9 9 1 15 3 0
8 10 3 9 0 13 13 0 0
15 13 3 10 9 3 3 10 0 0 9 10 0 10 9 13
9 13 3 0 0 13 10 9 10 0
43 13 3 10 9 15 7 13 0 7 3 3 11 7 10 11 15 3 10 0 9 13 7 10 0 9 11 10 11 11 3 0 15 11 10 0 13 1 11 1 9 13 9 3
19 11 3 3 0 16 15 13 13 10 9 13 1 11 7 15 13 1 10 9
16 13 3 10 9 7 3 13 0 9 9 13 1 15 9 15 13
31 0 3 13 0 13 3 1 15 10 0 13 15 10 3 9 13 13 11 3 13 3 9 1 15 9 7 15 13 0 0 13
41 9 3 10 1 11 13 16 13 10 9 10 11 13 7 10 9 10 0 13 10 0 1 11 0 3 11 10 0 9 10 0 13 3 13 10 9 0 13 1 10 11
21 10 3 1 11 9 13 9 1 0 13 11 15 3 13 10 9 0 9 13 10 9
10 0 3 3 9 0 13 3 1 0 13
40 11 3 13 11 9 7 11 7 7 11 15 9 9 13 3 0 11 9 13 10 1 11 13 9 7 13 15 1 10 9 10 9 16 13 10 3 13 10 9 13
21 11 3 13 1 10 1 11 9 13 3 11 13 3 11 7 7 11 7 11 7 11
6 0 3 1 9 0 13
19 1 3 11 13 15 1 11 9 13 9 10 9 10 0 9 13 13 1 9
11 13 3 1 10 11 13 10 9 1 10 11
28 13 3 10 9 3 13 9 15 7 0 7 0 3 13 13 15 11 10 11 9 9 15 10 9 9 11 13 9
35 0 10 9 10 9 13 13 10 11 10 9 7 1 9 13 10 9 3 13 16 3 13 3 13 10 9 3 7 13 13 13 3 0 10 9
35 0 3 3 3 13 10 9 7 10 9 1 9 13 10 11 3 3 15 3 16 9 10 9 13 7 13 10 9 16 3 13 1 10 9 13
28 3 3 13 7 13 10 11 10 9 3 1 10 11 9 13 7 10 9 10 9 7 9 13 0 7 1 9 0
5 9 3 13 1 9
11 9 3 3 13 9 1 12 9 3 1 12
18 3 3 10 13 15 13 1 11 1 11 0 9 0 7 7 0 9 9
22 13 3 3 0 3 13 1 9 15 7 13 15 0 9 7 13 10 3 10 11 0 13
9 3 3 15 3 0 10 9 13 13
7 15 3 3 13 1 9 13
13 7 13 7 10 9 13 7 13 1 0 3 0 13
8 13 3 10 15 0 3 0 13
11 1 3 0 10 9 13 7 7 13 10 9
34 13 3 16 13 13 10 9 1 10 9 15 13 10 1 11 9 1 15 13 10 9 9 13 7 0 7 10 9 15 11 7 11 7 11
10 10 3 9 0 9 13 9 11 9 9
7 0 3 3 10 9 3 13
39 0 3 13 16 13 10 11 13 11 7 13 1 11 13 10 11 1 10 11 13 10 9 7 13 3 9 15 15 10 11 13 13 3 9 10 13 10 0 9
12 0 7 11 13 0 10 9 9 13 1 10 11
5 0 3 3 3 13
19 11 3 10 11 9 7 11 10 0 9 13 1 10 11 7 10 0 11 13
8 11 3 3 11 13 9 3 11
9 3 3 15 3 0 13 9 11 13
4 0 13 10 11
29 11 3 3 10 11 9 9 0 3 1 15 13 13 10 9 1 11 3 10 9 9 13 9 13 16 13 1 10 11
5 0 3 3 11 13
11 0 3 11 10 0 9 13 1 10 11 13
10 10 3 3 11 13 11 9 10 9 0
17 0 3 13 15 10 13 13 1 10 11 7 13 10 9 1 15 13
7 11 3 3 11 13 3 13
11 11 3 10 11 9 13 1 11 13 1 11
17 13 3 15 1 10 11 13 11 10 11 9 1 15 15 13 9 13
16 15 3 3 13 13 13 7 10 13 3 15 3 10 13 9 13
8 3 15 11 13 1 0 10 9
6 0 10 9 13 3 15
3 13 3 11
17 11 3 13 3 13 11 1 10 0 13 9 13 1 9 9 11 13
16 15 11 9 10 0 13 13 13 10 9 10 9 10 1 11 9
17 13 3 1 11 13 1 9 13 1 15 0 13 9 1 15 1 11
13 13 3 10 9 10 15 9 16 0 13 9 13 15
33 3 3 13 1 10 9 10 11 1 15 15 3 3 13 10 11 13 1 9 7 0 0 13 9 13 10 3 13 15 9 3 3 13
9 15 15 3 0 9 13 13 10 9
22 3 3 10 11 1 9 13 11 9 9 10 1 11 13 9 13 9 3 13 15 9 1
6 13 3 13 10 9 11
30 15 3 13 15 10 13 13 10 11 10 3 1 10 11 13 13 15 3 13 10 3 0 10 1 10 9 13 11 15 13
10 0 3 13 0 13 3 0 9 10 11
6 1 11 3 3 13 9
13 11 3 0 13 10 9 9 13 1 11 0 11 13
19 10 3 0 0 13 3 11 3 0 13 0 9 13 1 10 9 15 9 13
7 13 10 9 1 15 10 0
10 15 3 13 12 9 13 1 11 1 11
20 3 3 13 10 1 10 11 13 10 9 13 1 3 15 15 11 13 0 13 13
7 11 3 3 7 0 13 0
11 1 3 11 0 0 0 7 0 13 9 0
20 13 3 10 9 10 9 7 12 13 9 13 1 10 11 10 0 9 1 0 13
7 10 3 0 9 3 13 0
11 13 3 7 0 3 13 7 9 7 7 0
41 13 3 0 1 0 10 9 7 13 13 0 3 9 15 13 0 9 7 10 9 13 0 0 10 3 0 13 13 15 10 9 13 3 13 10 0 1 11 13 10 11
12 10 3 11 13 9 0 1 10 9 10 0 13
18 1 3 0 13 10 9 13 10 9 1 3 15 3 9 15 10 11 13
3 13 3 3
12 10 3 1 10 9 13 9 0 0 9 13 12
22 13 3 0 9 12 9 7 0 12 9 0 3 0 13 12 9 0 3 13 9 12 9
16 1 3 0 0 7 13 7 9 0 3 12 9 13 9 3 12
6 9 3 13 0 9 12
13 15 3 0 10 15 9 13 12 7 12 7 12 9
13 0 3 9 13 10 3 9 10 9 10 9 13 12
50 16 3 3 0 13 1 10 0 7 10 0 15 0 13 3 10 9 9 13 10 9 10 0 9 13 16 3 0 13 13 7 3 3 10 11 0 3 13 13 3 3 13 9 1 7 11 13 0 15 13
35 0 13 13 10 9 10 9 15 1 11 3 10 0 13 10 9 13 1 9 13 3 3 13 1 10 11 0 10 9 10 13 13 13 15 0
11 9 9 3 15 15 3 13 13 10 9 9
12 10 3 15 0 15 9 13 13 1 10 0 0
28 13 3 13 0 16 13 7 0 15 1 10 9 7 15 7 10 9 7 10 0 13 7 0 13 15 3 0 13
45 16 3 0 3 3 13 15 3 3 1 9 13 0 3 15 13 13 15 3 15 13 16 13 10 9 13 7 16 15 10 9 9 13 10 3 9 0 1 11 7 16 10 9 0 13
18 10 3 9 1 15 3 13 0 10 9 9 7 13 7 3 13 10 9
9 15 3 0 13 0 0 10 9 13
11 0 3 3 3 13 1 10 11 10 9 13
17 3 3 10 9 13 1 10 11 13 9 7 3 3 15 3 0 13
10 3 3 3 3 10 9 9 11 13 0
19 1 9 3 9 13 15 10 9 9 9 7 13 0 7 9 7 0 3 9
14 3 3 15 16 3 13 9 13 10 3 3 9 15 13
19 16 3 9 7 7 9 13 15 15 13 9 16 3 13 15 9 9 10 9
17 7 15 15 9 10 0 13 13 7 3 13 10 0 7 13 0 13
9 0 13 10 9 13 15 0 10 11
38 15 3 13 3 1 9 10 9 16 10 9 13 9 13 10 9 1 15 7 10 9 13 10 0 10 9 10 9 13 1 9 13 7 10 9 9 1 9
11 1 3 3 9 12 13 7 7 13 10 13
21 10 3 1 0 10 9 15 0 13 9 0 13 7 9 7 7 9 13 1 15 0
5 15 9 13 0 13
6 13 10 0 3 13 15
28 0 13 7 1 0 3 13 15 13 7 3 9 9 7 13 1 10 9 13 7 13 3 13 1 10 9 7 13
10 3 3 13 15 13 0 10 9 9 13
24 9 3 13 16 3 13 10 9 3 13 13 0 1 9 13 13 10 7 9 10 15 7 10 0
16 10 3 11 1 15 10 9 13 10 0 9 3 13 11 10 11
18 9 3 13 11 1 10 0 11 13 10 9 3 3 10 0 10 11 9
15 3 3 16 13 10 9 10 9 13 3 0 10 9 1 9
3 15 3 13
23 13 3 0 3 1 10 13 1 10 11 13 10 9 13 1 10 9 1 10 11 1 12 9
10 0 3 10 9 13 7 13 13 10 9
12 13 3 3 0 10 0 13 10 0 13 10 0
11 3 3 3 10 0 10 9 13 10 0 0
17 10 3 13 1 10 9 13 0 9 3 13 7 9 0 7 3 13
19 13 3 3 3 3 0 13 9 12 7 1 0 15 9 12 10 9 9 13
11 9 3 3 10 0 10 9 13 1 10 15
18 15 3 10 9 0 13 10 9 1 9 0 3 16 13 13 1 10 11
7 9 3 3 3 3 13 13
7 15 3 3 13 1 10 9
29 11 3 10 9 16 13 10 9 10 9 13 9 13 12 10 0 13 1 3 11 3 3 13 16 13 1 10 0 11
8 15 3 3 16 13 13 1 11
11 9 3 3 13 7 9 13 0 13 1 11
27 13 3 0 1 11 1 9 10 9 10 15 13 0 9 10 3 1 0 10 0 13 10 3 9 13 1 0
15 10 3 3 1 10 0 13 16 1 0 13 10 9 3 13
9 15 3 10 0 3 13 13 13 3
14 7 3 3 11 0 0 9 0 9 7 7 0 9 13
7 15 3 9 0 9 13 9
17 3 3 0 10 0 13 16 9 3 10 0 13 1 10 9 13 9
8 9 3 7 9 1 9 9 13
13 10 3 1 10 9 0 9 3 9 3 10 9 13
8 3 10 13 10 0 13 1 11
25 9 3 15 11 0 15 0 13 13 1 10 0 13 9 1 11 9 1 15 11 9 13 1 9 13
16 10 3 0 9 0 3 10 9 13 10 1 10 9 7 10 9
7 10 3 0 13 9 9 13
20 13 3 0 0 1 9 3 13 10 0 9 15 11 7 7 11 13 10 9 13
10 9 3 0 3 3 15 15 13 15 13
5 11 3 3 0 13
18 0 3 10 15 13 10 3 1 10 9 1 10 9 10 15 13 3 13
25 0 3 10 1 11 10 0 9 0 13 1 10 11 9 13 10 9 1 0 9 13 3 9 13 9
15 10 3 0 0 9 13 13 3 9 1 3 11 13 10 11
14 0 3 13 10 0 0 9 13 1 3 15 0 10 13
7 1 15 0 3 15 13 13
28 0 3 13 1 11 13 1 9 10 0 7 0 0 7 7 10 9 15 15 9 13 11 13 9 10 9 13 13
6 13 3 3 15 0 9
33 16 3 15 7 10 11 1 10 9 13 13 11 3 10 9 10 0 3 13 10 9 10 11 13 7 10 9 15 11 1 11 9 13
13 10 3 0 0 13 10 0 7 9 13 7 13 13
29 9 3 15 13 13 0 1 10 0 15 10 9 7 9 10 0 13 10 1 10 9 10 3 1 10 9 15 11 13
12 10 3 3 0 10 0 0 1 9 9 13 13
9 10 3 9 15 12 13 10 0 13
7 3 3 10 3 0 13 0
12 11 3 10 10 0 9 1 10 11 13 1 11
15 7 15 13 11 15 9 0 13 15 1 10 11 1 15 13
24 7 3 13 9 1 11 13 7 3 1 10 11 3 1 9 16 15 9 0 0 13 13 1 9
9 0 3 13 9 3 9 0 11 13
26 1 3 10 9 10 1 11 13 9 13 9 13 1 11 11 10 11 3 0 7 0 13 15 7 0 13
22 7 0 0 10 13 1 11 1 10 9 10 9 1 10 9 7 10 9 7 10 9 13
8 11 3 13 3 11 13 10 9
10 15 3 3 10 9 13 15 3 9 13
5 0 3 3 3 13
20 0 3 13 0 1 11 13 7 9 9 3 13 15 13 1 11 13 10 0 9
26 0 7 3 13 0 7 10 0 9 3 3 13 1 10 9 10 11 13 10 0 13 1 11 10 9 13
14 13 3 3 13 16 3 13 0 0 7 9 7 9 13
8 7 3 9 1 0 9 0 13
13 0 3 15 13 1 11 9 9 12 12 0 0 13
7 10 3 12 15 9 13 13
26 0 3 1 10 9 10 0 0 9 0 1 10 9 9 9 13 13 10 9 16 1 12 9 12 0 13
11 1 3 0 10 9 13 1 9 10 9 13
8 13 3 10 9 9 3 15 13
12 3 3 10 11 13 1 11 13 9 7 9 0
17 13 3 15 11 13 9 16 10 9 13 1 10 11 1 10 0 11
7 13 3 0 11 3 0 13
10 0 3 1 10 11 13 13 15 10 9
27 1 11 3 13 15 10 9 3 13 1 10 11 3 13 10 9 10 7 3 7 10 1 11 9 10 10 9
16 15 15 13 13 0 7 11 9 13 7 10 9 15 10 0 13
5 13 3 10 11 3
8 10 3 9 0 13 13 10 9
27 10 7 3 9 10 9 0 13 7 13 10 9 10 11 13 3 13 1 9 1 10 13 9 9 0 15 13
24 16 13 7 13 1 9 9 7 16 13 1 15 13 13 0 9 13 13 15 16 13 11 10 0
25 16 3 3 16 13 13 13 1 9 11 15 3 7 3 13 0 15 13 15 13 7 3 15 10 9
37 3 3 15 0 7 0 1 7 16 3 13 3 0 1 9 13 11 7 10 11 9 7 10 13 11 16 13 13 1 11 10 3 15 9 3 3 13
37 11 3 13 0 7 13 10 0 13 16 15 3 13 13 1 9 10 15 10 9 10 11 13 7 7 13 3 13 13 3 9 3 15 7 7 9 9
6 10 3 1 11 3 13
28 10 3 0 9 10 9 13 1 11 10 0 9 16 13 13 3 10 9 10 1 10 9 13 11 7 11 7 11
5 13 3 0 10 9
23 9 9 13 10 9 1 9 10 0 1 10 0 13 7 3 1 15 10 9 13 13 10 9
13 13 3 3 10 1 10 9 9 10 0 1 10 0
5 3 3 13 10 9
15 3 9 10 9 3 13 10 9 15 13 10 9 13 0 15
11 0 7 3 13 7 10 9 13 0 10 9
16 3 7 10 0 9 13 0 3 1 9 3 3 3 3 1 9
15 1 3 11 13 10 0 9 10 1 0 13 10 11 13 15
29 13 3 10 1 10 11 0 10 11 11 7 1 15 9 0 13 7 11 7 10 9 10 1 11 7 11 7 7 11
27 0 3 3 7 10 3 0 3 13 13 10 9 7 13 13 10 15 3 1 10 0 9 7 3 9 11 13
15 10 3 9 13 0 10 9 10 13 13 1 7 11 7 11
6 1 3 11 3 13 3
19 0 3 9 3 0 10 9 9 13 1 9 11 10 11 13 10 1 11 9
12 10 3 11 1 11 9 10 0 15 13 10 9
20 13 3 15 1 3 11 10 11 10 11 13 10 9 0 0 11 10 11 9 0
6 13 9 9 10 11 0
22 10 3 11 15 13 9 13 1 10 9 0 15 3 15 13 1 10 9 0 1 0 13
13 13 3 10 9 10 0 9 1 9 7 7 9 13
11 1 3 10 11 3 13 3 10 15 9 11
33 3 13 3 3 11 10 11 13 9 0 10 3 3 1 11 7 7 11 13 10 3 0 0 11 10 11 9 13 0 10 9 0 0
27 0 10 11 13 1 10 9 10 15 13 10 9 13 9 13 3 0 7 9 13 7 15 13 13 9 7 0
11 15 3 13 7 13 1 15 13 15 10 9
8 13 3 13 15 10 9 15 13
17 11 3 13 3 13 10 9 3 13 7 10 11 9 7 13 3 13
32 13 3 3 10 11 3 3 11 10 11 0 13 0 0 0 3 13 0 15 10 13 13 10 9 13 1 10 9 7 13 10 9
25 15 3 0 3 13 10 9 10 11 1 11 9 1 11 16 3 13 15 10 0 13 13 1 10 9
10 13 3 0 9 12 7 7 12 10 9
14 1 3 10 9 0 10 11 3 15 13 9 12 10 9
19 13 3 10 9 10 11 10 11 7 10 0 9 0 13 10 0 0 13 9
7 7 15 10 9 13 13 9
10 13 3 10 11 11 10 9 1 9 13
11 13 3 10 11 0 13 13 10 9 13 11
8 13 3 10 9 11 13 13 11
6 0 3 3 1 11 13
17 3 3 13 9 10 9 7 7 10 9 13 11 10 11 9 9 0
21 7 15 13 9 13 3 9 9 7 9 0 7 7 0 13 1 15 9 15 13 13
29 9 3 13 1 9 3 11 13 13 9 13 10 9 9 1 10 9 1 9 0 3 10 9 0 3 7 0 10 9
49 13 3 3 11 9 0 3 11 10 11 11 3 10 13 9 13 10 9 1 11 13 9 10 9 15 15 3 1 11 13 3 3 3 13 3 10 9 11 15 10 9 15 15 1 0 9 13 3 13
14 11 3 13 1 10 11 13 1 9 10 9 11 3 13
13 10 3 9 13 0 13 1 15 10 9 10 13 3
18 11 7 3 13 10 11 12 13 9 7 13 11 10 9 9 10 9 11
11 0 3 10 11 11 3 3 13 1 10 11
9 13 3 15 13 0 10 13 9 0
8 0 3 3 9 1 0 9 13
15 9 3 10 9 13 1 9 11 13 7 13 1 10 11 0
19 0 13 3 13 10 11 13 11 16 15 10 7 9 13 7 0 9 13 3
11 0 3 3 0 9 0 13 10 3 15 13
18 3 3 13 13 10 9 1 11 13 9 12 9 10 13 13 1 10 11
12 0 3 3 11 1 10 12 10 9 13 1 11
10 10 3 15 0 10 9 13 13 10 9
23 10 3 9 0 13 10 11 9 10 0 9 11 3 1 10 11 10 9 13 9 7 1 0
45 7 0 1 10 9 13 10 9 7 15 13 16 13 11 9 13 1 9 13 9 0 13 16 3 11 9 13 1 10 9 13 13 10 9 16 10 9 13 13 10 9 13 1 10 15
17 11 3 16 10 9 11 10 11 13 13 0 3 15 11 0 3 0
18 7 3 9 7 9 13 7 0 9 1 15 15 9 13 15 1 9 13
8 11 3 1 11 13 1 10 11
26 11 10 11 9 13 9 1 10 9 9 15 0 10 9 13 13 16 0 13 7 3 15 13 7 7 13
9 13 3 3 1 10 0 3 0 13
6 7 15 0 3 0 13
37 1 3 10 9 10 0 13 9 1 9 11 10 11 13 1 9 9 0 3 3 0 3 13 0 3 0 9 7 0 13 7 3 13 9 11 9 11
22 13 3 10 9 0 10 11 16 13 1 10 11 0 3 13 1 9 13 1 10 0 9
10 9 3 10 0 0 9 13 1 10 11
44 16 3 13 10 11 13 10 11 1 10 11 3 0 9 13 10 3 13 9 9 10 12 11 9 13 16 0 13 13 9 10 3 9 10 9 13 15 10 11 9 13 1 10 9
29 16 3 13 3 9 0 9 13 3 3 0 9 0 13 10 9 10 11 13 1 10 11 13 3 1 7 11 7 11
8 0 3 3 15 9 13 10 9
10 0 3 10 0 9 1 15 13 9 13
11 10 3 1 9 9 15 15 13 3 0 13
12 1 3 3 11 13 3 1 10 9 13 1 11
7 1 3 11 13 10 11 13
21 13 3 15 13 9 9 0 7 7 0 3 3 13 9 0 10 9 13 1 10 11
24 3 3 0 13 10 9 0 10 1 10 11 15 3 1 10 9 13 13 15 3 1 10 9 13
13 15 3 15 13 3 13 7 1 0 13 15 3 9
7 10 3 3 0 9 3 13
6 7 15 0 13 10 9
4 11 3 0 13
8 3 3 3 0 9 13 1 9
15 3 3 3 0 13 1 10 9 0 11 16 3 15 0 13
11 0 3 3 10 9 3 13 13 1 10 11
29 0 3 9 0 10 11 0 3 0 13 1 10 0 16 9 13 13 9 13 15 10 9 13 7 10 9 1 11 13
26 10 3 3 0 3 1 11 7 10 0 13 7 9 13 0 13 10 9 9 7 13 0 7 9 0 13
13 10 3 9 15 13 1 7 10 9 7 1 10 9
34 13 3 3 0 10 9 0 7 0 13 15 0 15 10 9 13 15 1 11 13 10 9 0 15 3 1 10 11 0 10 9 10 9 13
25 10 3 9 10 0 0 13 10 11 1 11 7 9 13 7 11 0 3 11 9 0 13 1 10 9
5 0 3 3 13 0
20 1 3 0 13 10 11 10 9 15 15 1 9 13 3 13 15 7 13 15 0
16 13 3 9 15 3 13 1 10 11 13 13 9 9 7 7 9
7 0 3 3 1 10 11 13
19 0 3 9 13 1 10 15 0 9 10 0 13 9 7 0 7 0 9 13
28 0 7 3 13 0 7 10 13 1 10 11 9 0 3 9 13 15 13 13 10 9 15 3 9 1 15 13 13
39 13 3 15 0 3 0 13 13 7 1 15 13 10 9 13 16 1 10 9 1 15 13 7 0 9 13 13 7 1 10 11 13 10 9 15 13 13 10 11
19 1 0 3 10 9 11 10 11 9 13 9 13 1 11 13 13 9 10 0
12 1 3 15 9 10 0 13 0 1 0 13 9
9 1 3 3 15 10 0 9 13 13
7 13 3 0 1 9 10 11
15 11 3 13 1 10 11 13 10 11 15 15 15 13 10 9
6 15 3 15 10 13 13
6 10 3 11 1 15 13
28 1 3 10 11 0 10 9 13 11 10 11 13 10 11 13 9 3 0 9 9 3 10 0 1 0 3 15 0
8 1 9 3 3 13 3 10 11
29 0 3 13 15 9 13 0 11 10 11 10 11 10 11 13 13 15 1 0 10 9 15 3 13 7 3 10 11 9
13 1 3 9 3 0 11 13 10 9 15 9 13 11
12 9 3 15 13 13 11 10 11 10 11 10 11
4 0 3 13 0
8 13 3 10 11 10 9 9 13
14 0 3 10 3 13 13 1 9 9 10 9 10 0 13
6 15 3 3 0 13 13
14 13 3 3 10 3 13 0 13 3 16 3 0 13 9
5 10 3 3 0 13
11 13 3 13 1 11 13 15 15 13 10 9
15 10 3 11 15 13 0 10 9 13 9 13 3 3 10 0
7 10 3 3 11 0 15 13
18 10 3 0 13 15 0 3 13 15 10 0 13 9 0 15 9 13 11
18 13 3 0 10 11 0 10 0 13 10 13 15 10 9 0 13 7 13
22 16 3 13 3 0 3 13 0 15 13 16 7 0 0 15 13 1 0 7 13 15 9
31 3 3 10 9 1 10 10 0 9 13 10 9 10 11 9 13 1 10 0 13 10 0 7 9 7 9 3 13 15 1 13
16 13 3 10 9 10 13 1 10 13 3 13 0 13 1 10 0
8 7 15 9 13 11 15 3 11
22 0 13 0 7 9 13 13 0 13 10 15 9 10 9 15 7 10 1 0 13 3 13
6 0 3 0 13 0 9
31 0 3 1 10 13 1 9 15 13 0 10 9 9 1 3 3 11 10 11 10 9 13 13 3 1 9 7 13 16 13 9
7 3 3 3 1 9 0 13
20 1 3 11 10 11 13 10 3 3 9 15 13 3 13 10 10 9 9 0 0
8 0 3 3 1 15 9 13 13
19 3 3 10 1 9 9 13 0 10 11 13 0 13 9 7 3 10 11 9
18 10 3 11 3 9 13 1 9 11 15 0 3 13 3 3 9 13 0
7 7 0 3 3 1 0 13
8 15 3 15 3 13 0 9 13
24 9 7 3 0 10 9 9 13 9 12 11 7 11 7 11 0 7 9 13 1 15 3 13 9
8 16 3 3 15 1 10 9 13
3 0 3 13
8 12 3 9 9 1 9 13 15
10 9 3 13 1 10 9 15 3 3 13
12 10 3 13 15 10 9 7 7 10 9 13 15
4 0 3 10 0
9 10 3 15 10 0 1 0 15 13
31 9 3 15 7 0 13 10 9 13 1 10 0 9 0 0 1 11 7 9 9 7 9 0 0 7 1 10 9 15 9 0
15 7 0 13 0 13 15 3 13 10 9 7 0 13 12 0
21 3 13 3 10 9 1 10 9 13 15 1 10 9 9 7 12 9 0 7 9 9
5 13 3 0 15 13
11 10 0 3 0 3 1 9 13 1 9 13
7 10 3 9 10 13 0 13
5 13 3 3 10 0
10 7 16 15 0 9 13 13 9 1 13
9 7 13 13 10 9 13 12 13 12
22 16 3 3 13 10 3 15 10 9 13 13 10 10 9 9 12 9 13 0 3 10 15
8 9 13 10 13 1 15 10 0
8 1 3 10 9 9 13 9 13
16 16 3 0 13 0 9 1 9 0 0 12 13 9 7 7 9
7 3 13 3 0 9 0 13
15 10 3 3 9 10 0 10 0 9 13 1 10 9 10 9
19 16 3 13 9 0 1 15 13 11 1 9 9 10 0 0 1 10 9 13
38 0 3 7 10 9 7 0 9 16 13 1 10 0 0 9 3 10 9 13 7 10 9 3 7 9 13 0 13 10 0 3 13 10 9 0 3 13 0
17 15 3 3 1 9 10 9 13 0 3 9 13 1 9 3 13 13
7 13 3 15 0 0 10 9
20 16 13 10 9 0 13 9 0 10 13 13 15 15 9 10 9 7 10 0 13
14 1 3 3 9 10 13 9 10 13 9 13 10 9 15
22 10 9 15 7 9 7 9 13 10 0 9 7 9 7 9 13 7 9 9 7 9 9
12 3 1 9 13 15 15 13 7 1 10 0 13
5 0 3 3 3 13
26 3 3 10 11 13 1 10 11 7 0 10 11 0 13 10 11 13 3 9 3 13 3 9 7 9 13
18 11 3 13 1 11 13 10 11 13 10 9 1 9 0 9 1 15 13
8 7 3 3 13 0 0 13 0
3 13 0 9
13 13 15 9 10 9 9 15 13 10 9 3 10 11
19 0 10 9 13 13 9 0 0 10 1 11 9 7 0 3 0 1 0 13
33 13 3 15 10 9 0 10 9 15 3 9 7 0 9 7 0 13 3 3 3 13 10 9 9 10 9 15 13 0 0 13 13 0
10 13 15 1 15 9 1 10 10 11 9
11 15 3 13 1 10 11 13 1 10 0 9
19 16 3 13 10 9 1 7 10 9 13 7 13 10 9 13 10 9 10 9
10 13 3 13 15 15 15 13 1 10 9
5 15 3 13 15 13
4 15 3 3 13
8 13 3 15 1 10 13 15 13
6 15 3 3 15 13 13
15 13 3 10 9 1 0 13 13 3 3 10 9 13 10 9
15 15 3 13 10 9 10 9 13 16 13 15 10 1 11 9
9 1 3 3 0 10 9 13 10 9
10 10 3 11 13 3 10 9 0 10 9
3 13 3 0
30 0 7 10 9 15 13 10 9 0 13 9 13 10 15 15 12 15 3 0 0 13 7 10 9 15 13 3 10 0 13
14 15 3 15 13 1 10 9 13 13 3 11 9 13 0
5 1 0 3 9 13
36 3 3 0 7 10 11 13 0 15 15 3 13 15 13 10 9 10 11 10 11 7 0 10 0 13 13 1 0 3 3 10 9 10 9 13 13
9 15 3 1 0 0 10 15 13 13
12 13 3 10 7 9 7 10 9 10 9 13 13
19 1 3 15 9 0 7 3 13 10 12 9 10 9 0 13 0 3 10 11
16 7 15 15 10 9 1 9 13 1 10 9 13 16 15 9 13
18 15 3 13 7 10 9 15 13 10 9 7 1 9 13 10 9 13 13
4 3 3 15 13
5 0 13 3 10 9
6 9 3 15 13 10 3
10 10 3 9 13 7 10 11 10 13 13
10 9 3 10 11 1 10 3 15 13 13
8 1 0 3 15 10 9 11 13
6 9 3 13 11 3 13
5 11 3 13 10 9
29 13 3 13 10 11 13 11 10 11 10 11 13 9 10 0 11 16 15 7 16 15 13 9 1 11 13 15 1 9
12 10 3 11 13 0 10 11 3 13 1 9 0
23 13 11 11 10 11 10 11 9 10 11 13 13 11 10 9 13 0 10 11 13 7 13 9
12 1 0 3 10 11 10 9 10 1 10 11 13
20 1 3 10 9 13 13 0 10 9 15 13 11 3 16 15 13 10 9 9 13
33 0 3 13 10 9 10 11 13 10 11 7 1 11 13 7 3 13 11 10 9 9 13 0 15 3 13 0 7 13 7 13 0 11
20 9 3 13 1 15 9 13 9 13 10 9 10 1 11 16 11 13 9 10 11
21 0 3 13 1 9 10 11 1 10 11 3 13 11 11 10 11 9 1 11 13 0
12 10 3 11 11 10 9 13 15 11 13 13 13
13 3 3 10 11 13 10 9 13 3 11 13 11 9
19 0 3 9 0 13 0 7 11 7 13 1 9 7 11 10 9 13 10 9
10 13 3 11 1 11 1 9 1 0 9
10 1 10 9 10 9 10 11 13 13 9
31 13 3 10 11 10 11 13 3 9 0 1 0 13 10 9 1 9 7 7 9 13 10 11 15 15 13 10 13 1 10 13
27 15 3 13 10 9 13 13 0 3 15 3 13 0 3 3 10 3 9 0 13 0 7 0 9 7 0 9
13 0 3 13 7 13 13 1 10 9 1 10 15 9
7 3 3 13 13 10 11 9
5 13 3 10 9 13
24 6 9 9 15 10 7 0 13 13 7 10 0 11 0 13 15 10 9 15 15 13 9 0 9
18 11 3 3 13 1 10 9 13 13 15 1 10 0 9 3 13 1 11
20 15 3 3 10 0 9 13 13 15 13 1 10 9 10 9 7 15 0 13 9
14 7 3 16 3 13 15 10 13 0 3 13 1 0 3
12 10 7 9 0 1 11 16 11 9 0 3 13
8 13 3 3 15 3 10 0 9
5 15 3 3 0 13
15 6 9 16 15 9 13 13 10 9 15 1 15 13 10 0
16 16 15 13 11 1 15 9 0 1 10 0 13 15 9 13 11
8 13 3 10 9 15 13 15 13
4 7 15 3 13
12 16 3 15 13 13 9 13 15 13 15 10 13
4 15 3 13 0
4 15 3 3 13
11 0 3 15 0 13 7 13 13 15 10 9
12 13 3 15 13 10 11 13 16 0 13 10 9
20 7 0 3 10 9 13 13 1 10 9 10 1 10 9 10 0 13 15 13 11
10 0 3 10 9 10 0 0 9 13 13
10 3 6 9 13 15 15 15 3 13 13
7 1 3 15 10 9 0 13
40 3 3 15 3 13 10 0 13 16 0 10 11 16 15 15 13 13 0 13 3 13 15 15 13 10 9 3 10 12 9 3 13 9 10 0 0 0 13 10 9
7 15 3 15 6 9 0 13
16 13 3 3 0 10 11 3 1 0 9 16 9 10 9 13 0
9 9 3 0 1 9 10 15 3 13
5 10 3 0 15 13
14 1 3 9 0 7 11 7 10 0 13 13 10 9 9
5 15 3 3 0 13
7 0 3 13 11 9 13 13
12 13 3 10 0 15 7 13 7 10 9 15 13
16 3 3 3 3 13 15 10 0 3 13 1 10 11 1 9 11
12 15 3 13 7 15 3 7 9 7 7 9 13
19 3 13 1 10 11 11 7 0 13 9 15 7 0 0 9 7 7 9 13
19 3 3 3 3 0 15 13 0 13 0 0 15 3 10 13 9 1 11 13
20 11 3 10 11 11 13 13 10 9 7 15 13 9 11 15 3 11 15 9 13
6 0 10 11 3 13 11
13 3 3 3 11 13 1 11 7 9 0 15 11 13
4 13 0 1 11
9 13 3 15 15 0 13 13 9 0
23 1 0 3 13 3 1 10 9 13 9 0 9 13 1 11 1 9 13 7 10 9 15 13
8 13 3 1 11 7 13 1 0
6 0 3 3 13 9 0
26 3 3 16 10 11 13 10 1 10 11 9 3 13 11 13 1 10 9 0 15 15 0 1 10 9 13
27 3 3 3 10 9 15 10 9 13 1 15 13 3 13 0 3 13 9 12 9 10 0 0 7 9 7 9
14 13 3 15 1 9 10 0 9 13 1 10 0 9 0
16 1 3 0 11 0 13 13 1 11 9 13 9 7 13 1 11
45 3 3 13 1 10 11 0 13 9 13 10 9 1 10 11 15 7 9 13 15 3 3 13 15 15 3 3 13 7 3 3 1 11 9 0 13 10 9 10 13 13 13 10 11 9
19 1 3 0 10 9 13 13 1 10 9 10 11 9 7 3 3 13 0 15
8 9 0 13 1 9 13 1 9
7 10 3 9 9 15 13 9
16 10 3 11 1 15 10 9 0 13 13 9 13 10 11 1 11
18 13 3 11 0 0 13 13 15 13 1 10 0 1 11 15 3 0 13
11 13 3 15 0 7 13 13 10 13 1 9
11 15 3 13 10 9 13 13 10 0 13 9
28 3 13 3 10 0 10 9 13 13 15 15 3 13 16 15 13 10 9 10 9 13 3 10 15 9 13 15 9
11 11 3 13 10 9 13 1 10 9 15 13
13 13 3 1 9 10 9 13 1 10 9 1 10 9
77 1 3 10 9 1 7 10 9 7 10 9 16 15 1 10 9 13 7 0 13 13 9 0 3 3 10 0 13 9 16 10 11 13 10 1 11 13 13 3 3 0 0 13 16 1 11 13 13 10 9 10 9 3 3 0 16 1 9 15 10 11 0 10 13 1 10 9 13 13 7 0 10 9 1 9 13 13
8 11 3 13 1 11 13 11 13
7 7 3 3 13 3 13 15
15 13 3 10 9 9 9 15 13 1 7 10 0 9 7 11
7 0 3 13 13 0 1 9
23 16 3 1 3 13 10 11 9 3 1 0 15 13 11 9 0 3 0 13 13 0 10 0
16 3 3 10 0 10 3 1 10 0 9 3 13 7 16 9 13
22 7 3 3 15 1 0 10 9 13 10 9 15 0 13 10 11 0 7 7 0 13 3
18 7 3 10 0 10 0 13 13 7 9 1 0 13 0 0 0 3 13
6 0 9 0 13 9 13
8 0 3 15 13 10 0 9 13
5 9 3 15 13 0
14 16 10 9 9 13 15 0 13 3 10 0 10 0 0
29 13 3 10 11 13 10 0 15 15 10 15 9 13 13 15 3 13 10 9 13 9 3 13 10 9 13 1 10 0
7 0 3 13 0 1 10 0
14 9 3 13 10 0 1 10 9 13 7 0 3 13 15
6 3 3 10 11 13 0
25 13 0 9 7 13 0 13 13 9 3 13 10 0 10 1 10 9 13 13 3 13 15 13 10 9
11 9 3 13 0 12 9 13 1 9 0 13
11 0 3 3 13 13 10 0 10 1 10 9
26 3 3 0 13 10 9 3 13 10 3 10 3 15 15 13 16 3 3 15 15 13 1 9 13 10 13
5 3 3 3 13 13
13 3 3 10 11 13 15 15 10 9 13 9 10 9
12 13 3 3 13 10 15 0 15 13 9 10 9
5 15 3 13 11 13
7 15 3 16 13 13 0 13
10 6 11 0 3 3 15 13 13 11 13
13 1 3 0 10 11 10 3 0 9 13 13 1 11
11 12 3 0 13 10 9 13 1 10 0 13
17 13 3 15 13 1 10 9 10 9 13 13 3 0 13 9 3 13
7 13 3 0 13 1 10 11
20 13 3 15 13 10 0 1 10 9 13 15 13 3 13 10 11 13 3 15 13
15 16 3 3 1 10 9 10 9 13 13 3 1 9 10 9
14 0 13 0 7 7 9 13 9 13 7 13 0 10 13
24 11 3 9 13 3 16 10 9 15 13 15 10 9 9 7 7 13 16 15 13 10 10 13 9
7 13 3 10 9 9 13 11
8 3 3 3 15 13 0 1 15
7 0 10 9 13 13 10 9
16 1 0 3 9 15 13 1 9 0 16 15 3 3 10 0 13
10 0 3 3 1 0 11 13 13 13 3
20 0 3 9 13 1 9 3 15 13 11 9 3 13 15 9 13 7 1 0 13
21 11 3 13 13 10 9 1 0 13 15 3 13 3 3 10 13 13 10 9 1 15
7 1 0 3 13 15 13 9
7 3 3 9 10 1 11 13
18 13 3 11 16 13 9 13 1 11 9 13 11 1 10 1 11 9 13
22 0 3 9 13 13 13 9 1 11 7 15 13 0 13 1 11 1 10 1 11 13 9
17 13 3 13 10 9 10 11 13 15 11 10 11 13 1 11 0 9
5 15 13 13 9 9
7 0 13 10 9 13 10 9
12 9 3 13 0 13 11 1 11 13 9 10 9
10 3 13 3 13 10 0 13 15 11 0
17 13 15 10 9 13 1 10 11 1 0 9 10 1 15 11 11 9
26 0 10 9 13 10 7 0 15 13 10 0 7 3 3 13 0 9 1 15 15 10 11 0 10 9 13
8 13 3 15 1 9 13 0 13
12 9 0 13 1 11 13 15 13 1 9 13 0
3 13 3 0
8 13 3 10 15 11 13 9 13
26 0 7 3 13 7 13 13 15 10 0 15 10 9 13 13 1 15 3 13 16 15 13 13 1 15 0
13 15 3 15 7 10 9 13 7 0 10 9 13 13
9 10 3 3 1 11 13 9 0 13
9 11 3 13 10 9 1 10 13 9
14 9 3 0 13 13 1 11 0 10 13 10 9 10 9
13 13 3 1 9 10 11 7 13 10 9 13 10 9
5 15 3 13 13 0
18 7 3 16 13 3 13 7 16 3 9 3 13 9 10 9 13 1 15
10 0 3 15 13 13 1 0 9 1 0
11 10 3 3 0 9 13 13 3 13 10 9
12 11 11 10 3 3 0 3 9 13 7 9 13
8 13 16 9 3 3 0 13 9
10 7 9 9 13 0 7 13 9 7 9
13 0 3 13 16 15 3 15 13 13 9 7 9 0
6 9 3 0 9 3 0
12 0 13 10 11 9 10 9 13 15 13 10 13
13 10 3 11 13 10 13 10 9 7 10 13 0 13
13 15 3 1 10 9 0 6 0 13 13 1 15 13
12 11 3 13 0 16 15 3 3 13 10 0 13
17 10 3 9 16 10 0 9 13 9 15 1 0 13 0 13 13 0
11 13 10 0 7 13 13 3 13 10 0 13
9 7 13 3 3 10 0 9 1 11
11 13 3 10 9 9 13 0 9 10 0 0
5 13 3 10 9 13
11 7 13 3 11 11 13 1 10 11 9 0
14 1 0 13 3 1 15 13 0 10 11 10 0 13 9
13 1 15 3 0 13 13 15 9 1 0 13 10 9
22 10 3 0 13 3 15 0 10 9 9 1 10 3 0 13 13 12 9 13 3 0 13
8 9 3 1 10 9 3 13 13
24 0 7 3 13 10 0 7 10 15 13 12 9 10 0 13 1 10 11 7 13 9 12 10 13
17 11 3 16 10 0 1 10 9 3 13 1 9 13 13 1 10 11
13 3 3 0 13 13 7 7 13 10 1 10 9 9
5 0 3 3 0 13
17 9 3 10 0 13 10 9 15 1 11 13 7 3 15 13 13 13
9 12 3 3 10 9 13 13 3 13
12 12 3 15 0 13 10 9 13 1 9 11 0
5 13 3 10 9 13
16 15 3 16 15 13 3 0 3 13 13 13 15 10 9 13 3
8 0 3 3 15 0 10 9 13
6 0 3 13 13 9 12
10 13 3 10 9 13 10 0 3 0 0
11 7 15 1 0 13 9 12 9 13 12 0
7 9 3 7 13 13 7 0
11 13 3 15 9 9 15 9 11 9 9 13
12 0 10 0 3 13 3 7 13 1 0 1 11
8 1 3 10 0 11 10 11 13
18 9 3 13 0 10 0 13 10 9 13 7 15 9 12 0 10 9 13
7 0 3 3 9 13 1 9
10 11 3 3 3 13 10 9 13 10 9
22 15 3 9 13 13 1 7 11 7 11 11 7 13 9 9 7 11 10 11 9 9 15
37 16 3 10 9 0 10 13 13 1 9 13 10 11 1 10 11 9 3 13 0 9 0 7 7 3 13 3 13 13 3 10 0 15 9 10 13 0
16 13 3 3 10 0 9 15 10 0 9 13 10 15 0 11 13
49 3 3 3 1 10 9 13 10 9 3 10 7 11 7 10 11 7 1 11 13 1 7 0 7 1 9 10 9 13 3 3 15 13 13 3 10 9 10 11 16 10 0 9 13 3 10 9 3 13
10 3 3 3 10 11 15 13 0 3 13
31 16 3 1 10 0 9 13 13 10 11 1 0 3 3 0 13 13 10 9 13 10 0 10 0 1 10 9 13 13 7 13
8 0 3 13 1 10 0 9 13
17 16 15 3 0 0 13 10 0 13 3 0 10 11 13 13 1 11
20 10 3 9 13 10 11 13 3 13 10 9 1 10 11 13 7 3 1 10 11
10 9 0 15 13 13 3 0 13 1 15
12 3 3 7 13 1 10 15 15 7 10 9 13
5 0 3 13 10 0
10 3 3 9 12 9 13 1 10 9 13
19 11 3 3 0 13 13 1 10 9 1 10 11 0 3 13 7 9 7 9
13 7 0 3 3 9 9 10 13 13 0 13 10 9
10 3 15 13 0 13 11 10 3 13 0
8 7 1 9 13 13 1 15 3
14 0 3 3 10 9 3 3 3 1 9 10 15 9 13
12 10 3 0 16 13 1 10 11 13 1 10 9
11 3 3 9 7 13 7 9 10 9 9 13
15 9 3 13 10 9 10 0 1 15 13 0 13 15 0 13
20 0 3 3 13 10 9 7 10 12 10 13 10 9 9 10 9 0 15 13 0
8 10 3 9 13 3 15 0 9
4 15 13 3 0
4 13 3 0 9
12 15 3 15 0 9 13 1 10 9 13 9 13
33 13 3 0 0 3 13 11 10 11 13 10 9 10 0 13 10 13 0 15 10 13 15 9 13 7 13 15 1 10 15 16 3 13
7 10 3 0 0 11 13 13
9 7 0 3 13 1 11 13 15 0
16 10 3 9 13 13 10 9 10 0 9 1 11 7 11 7 11
15 13 3 0 10 9 3 9 7 13 7 13 3 13 10 0
10 10 3 9 13 3 7 13 3 13 9
16 16 3 3 13 10 9 0 15 1 13 16 13 3 13 10 9
18 15 3 13 1 10 9 0 3 10 9 13 13 13 10 1 11 13 9
9 0 3 10 9 13 1 10 11 9
28 13 3 10 11 7 13 0 9 13 1 9 10 0 13 7 0 7 13 10 0 10 0 13 15 3 10 9 13
14 7 13 3 10 11 0 9 10 11 13 7 3 10 11
7 1 0 15 13 11 10 11
11 0 3 16 13 0 13 7 0 1 10 11
10 13 3 15 9 12 15 10 0 13 11
21 7 15 13 9 13 0 13 7 0 3 10 9 13 15 10 0 13 10 0 9 11
18 7 15 13 10 0 9 0 9 13 13 1 10 11 9 3 13 0 11
10 13 3 0 15 1 10 9 9 13 9
12 13 3 11 1 10 9 1 10 1 11 13 9
11 3 3 15 10 9 13 0 10 12 9 13
15 13 3 3 15 9 3 10 0 0 11 11 0 3 0 0
36 10 3 3 0 10 9 10 11 11 13 3 1 10 9 11 13 1 10 11 10 3 0 1 0 11 1 11 9 13 1 10 9 10 11 11 11
19 3 3 3 10 9 15 15 13 1 11 1 0 13 13 7 7 13 1 9
31 3 3 13 7 0 7 13 1 10 15 13 7 13 1 9 3 10 3 15 10 0 13 1 9 15 13 13 9 10 1 11
25 7 0 3 13 3 1 10 9 10 9 13 1 11 9 11 0 3 9 3 3 9 7 7 0 13
20 15 3 3 0 7 13 11 7 0 13 1 10 0 9 10 1 11 10 11 13
32 13 3 10 9 10 11 10 11 0 13 13 1 15 15 15 15 9 13 13 0 0 7 3 13 15 3 0 15 3 3 3 13
30 7 0 3 0 13 15 3 3 10 9 13 13 0 13 1 10 9 11 9 7 15 1 0 10 9 9 0 7 9 13
25 3 3 13 1 10 9 10 11 0 16 3 15 13 3 10 11 13 0 1 10 0 9 13 1 11
20 6 0 0 15 13 15 13 7 3 13 9 0 1 10 9 9 13 1 9 9
13 7 3 3 11 7 13 7 9 0 10 11 13 0
7 15 3 3 15 10 13 13
13 0 3 15 13 10 3 13 0 3 13 13 10 9
6 13 3 13 10 9 0
11 0 3 3 13 13 3 3 0 13 10 9
6 0 3 3 10 0 13
8 13 10 11 10 9 10 15 13
18 13 3 1 10 9 13 1 10 11 7 13 10 9 13 1 10 15 0
7 1 3 3 10 9 13 0
19 3 3 13 0 3 10 9 10 1 11 13 1 10 9 10 9 13 3 11
13 7 15 0 13 13 13 7 7 13 3 3 3 13
10 3 3 15 0 13 10 9 10 0 13
9 0 3 12 10 9 13 1 9 13
12 16 3 3 13 15 10 9 13 13 1 10 9
11 10 9 0 3 15 13 7 15 13 0 13
9 15 3 15 15 9 13 10 9 13
8 11 3 3 3 10 9 13 13
10 0 3 13 1 9 11 13 13 9 3
3 13 3 3
16 13 1 0 10 9 13 0 13 11 7 10 11 7 0 15 0
13 15 3 3 7 13 7 15 0 15 13 3 9 0
9 13 3 3 3 13 3 15 13 15
15 13 3 15 13 15 0 0 0 7 9 7 13 13 3 0
19 0 13 10 0 3 1 10 9 3 10 9 3 13 10 0 13 9 13 9
6 0 3 3 9 0 13
19 15 3 3 13 7 0 0 13 10 12 9 9 13 1 10 9 13 15 0
4 0 3 15 13
20 13 3 7 13 13 15 13 10 9 1 0 13 0 9 10 3 13 1 9 13
6 0 3 3 0 13 13
5 0 3 13 13 9
5 13 3 13 10 9
24 13 3 10 0 15 10 0 13 9 13 9 0 13 10 11 0 13 9 0 1 9 13 7 11
11 13 3 3 10 11 15 0 0 9 10 13
6 13 3 3 1 11 13
11 3 3 3 1 15 13 0 1 9 13 0
12 7 16 3 3 13 10 9 13 15 13 13 11
14 16 3 13 0 10 9 0 7 13 0 10 0 9 13
23 3 3 3 0 0 7 13 13 7 3 1 15 3 0 13 10 9 10 9 13 3 13 13
16 15 10 9 13 12 3 13 10 9 15 3 13 15 3 3 13
11 0 3 15 1 15 3 13 7 1 15 13
19 16 3 15 9 10 15 13 13 15 9 7 0 7 9 0 10 1 10 11
16 16 3 10 10 13 10 9 13 13 15 15 15 13 0 10 0
8 13 3 10 9 10 9 13 13
18 3 3 10 9 15 10 9 13 13 16 0 15 13 9 10 9 11 13
13 15 3 13 3 3 9 13 16 3 3 15 9 13
13 16 3 1 0 13 3 3 13 3 10 0 3 13
8 10 3 0 9 13 10 9 11
14 10 3 9 3 13 3 10 0 10 9 13 9 10 0
10 13 3 0 13 3 13 10 9 13 15
8 0 3 13 13 10 0 9 9
6 10 3 9 0 13 9
10 13 3 9 3 0 10 0 15 3 12
6 0 3 3 10 0 13
10 0 3 16 0 13 10 9 13 3 9
12 0 3 3 9 15 15 15 13 9 1 0 13
12 0 3 13 9 7 0 13 7 10 9 0 13
12 3 3 13 10 9 3 10 9 10 9 9 13
13 1 0 3 3 13 10 0 7 13 13 1 10 0
9 13 3 10 3 13 10 9 13 13
14 10 3 10 0 13 15 13 10 9 0 13 7 13 0
19 13 3 10 9 13 13 16 15 1 10 9 13 9 7 13 7 13 10 9
13 7 0 3 1 0 10 9 10 9 13 9 13 0
8 3 3 13 10 9 11 10 11
23 0 3 11 10 11 3 13 10 9 9 10 9 13 9 13 0 3 15 0 0 7 7 0
28 10 3 0 10 0 13 7 13 1 10 9 1 15 13 10 1 11 9 13 11 13 13 10 0 13 1 10 9
11 9 3 13 1 0 1 9 9 15 0 13
5 0 3 3 13 11
24 10 3 0 10 9 13 11 0 3 13 9 3 10 0 1 0 13 10 9 13 3 1 10 11
21 1 0 10 1 9 9 13 10 9 1 12 7 12 9 0 3 12 7 12 7 12
4 13 3 15 0
23 13 3 15 1 10 9 13 0 15 9 9 15 13 9 13 0 15 10 9 10 9 15 13
5 10 3 15 9 13
6 0 3 3 11 13 13
18 11 3 13 1 10 9 1 10 11 16 13 1 11 13 9 1 10 9
10 15 3 16 9 3 13 9 13 10 9
12 13 3 1 9 0 9 11 13 13 3 13 13
12 13 3 1 15 13 9 13 10 15 9 1 11
35 7 13 3 3 10 0 3 1 10 9 13 7 1 10 9 10 9 7 13 10 0 13 10 9 1 11 10 0 15 3 13 1 9 11 3
19 10 3 9 0 0 3 13 7 15 1 9 12 0 0 1 9 13 1 11
18 10 3 10 9 13 11 7 7 11 16 13 1 10 11 13 13 1 11
45 16 3 13 15 13 1 15 7 15 0 13 13 0 15 15 7 15 10 0 9 13 1 9 15 15 9 13 11 1 3 11 12 7 0 9 13 12 3 1 10 9 15 13 0 9
12 7 3 9 7 9 7 9 13 1 15 9 0
7 1 3 9 0 9 15 13
9 13 3 0 13 7 3 13 1 9
9 1 3 0 1 15 13 13 0 9
8 10 3 9 10 9 13 0 9
7 13 3 0 7 9 13 0
18 3 10 9 13 9 11 15 3 1 15 13 10 9 0 13 10 0 9
7 10 3 3 1 9 13 3
23 0 3 13 1 10 11 12 1 10 0 13 9 0 13 3 16 0 1 11 13 1 10 11
6 13 3 1 10 11 13
10 3 3 13 0 7 10 9 15 13 3
13 15 3 7 3 11 10 11 11 3 9 13 0 13
30 11 7 3 0 0 0 13 16 11 13 1 10 11 10 9 15 13 1 10 0 13 7 10 0 10 0 1 15 15 13
10 11 3 0 0 3 9 13 15 15 13
11 0 3 3 10 13 3 9 0 13 10 9
6 0 3 15 1 11 13
17 9 13 0 3 0 13 11 3 0 13 13 1 10 9 15 9 0
12 16 3 13 9 0 13 15 9 0 0 7 13
10 7 10 9 3 7 15 0 0 13 0
23 9 3 3 13 16 3 0 3 3 13 10 10 11 13 13 0 13 10 11 3 15 0 13
11 7 3 3 15 13 0 10 9 13 10 9
15 3 3 3 13 15 15 0 1 3 0 9 7 15 3 13
13 3 3 9 13 13 1 3 3 0 9 1 0 9
10 13 3 3 9 7 0 3 13 3 13
2 13 3
10 1 3 11 7 3 11 13 3 3 0
42 0 3 3 11 10 11 10 1 11 9 1 11 13 1 10 9 10 1 11 9 7 13 7 13 3 7 15 11 13 10 9 10 1 10 9 13 15 3 13 13 1 11
12 13 3 13 9 0 3 13 10 15 9 13 3
11 10 3 11 1 10 9 13 0 0 13 13
24 13 9 0 7 9 0 13 10 9 9 7 15 13 0 13 13 13 1 10 9 1 15 15 13
17 13 3 1 9 9 0 3 13 1 10 9 10 9 15 13 10 9
8 15 10 7 9 13 7 15 13
19 13 3 10 11 9 13 7 15 15 7 0 13 7 3 0 13 3 0 0
14 11 3 10 11 10 11 10 11 13 9 15 9 13 11
10 0 13 9 0 13 10 0 0 9 13
40 0 3 13 7 13 1 15 0 10 11 9 13 15 9 15 13 11 9 13 13 1 0 9 7 3 0 1 11 3 13 11 10 9 1 9 1 10 0 13 9
12 3 9 15 15 7 0 13 7 9 13 13 9
11 15 11 7 9 7 9 13 1 0 0 13
33 1 3 3 11 13 11 10 11 9 15 1 0 3 9 12 9 13 10 3 11 13 0 10 9 3 7 9 11 11 10 0 13 9
14 0 3 1 11 13 1 3 10 9 10 0 11 11 0
6 0 3 1 10 0 9
38 0 7 3 9 7 11 11 9 1 11 7 9 1 11 9 11 11 10 13 7 3 9 1 11 13 10 9 9 7 1 0 13 15 9 7 0 11 11
7 0 3 3 1 0 11 13
22 1 3 11 13 11 7 10 11 0 10 1 11 13 7 0 11 11 9 7 9 13 0
8 1 3 11 13 0 10 9 11
5 0 3 1 11 0
5 0 3 13 10 9
19 13 3 0 1 10 13 9 10 11 0 3 10 9 7 15 13 7 9 0
33 16 3 10 0 13 10 9 10 7 9 10 9 7 9 0 11 15 13 1 15 13 9 12 10 11 13 0 7 10 9 7 0 15
16 13 3 10 9 13 0 10 15 10 11 13 15 10 9 13 9
5 13 3 10 9 13
6 7 3 15 3 3 13
8 10 11 3 13 0 10 9 13
10 3 3 13 10 11 9 13 15 9 13
15 13 3 10 9 0 3 1 15 13 0 9 1 3 0 0
30 11 3 10 3 0 7 10 0 13 13 9 3 15 3 13 11 1 10 7 9 7 10 9 13 15 3 13 13 1 15
10 16 3 13 10 9 13 3 13 13 13
5 10 3 11 13 13
3 3 9 11
5 1 0 3 0 13
8 11 3 9 13 13 1 0 0
28 9 9 10 15 9 15 7 15 15 13 7 15 15 16 0 7 13 13 3 7 12 15 0 13 7 10 0 13
8 13 3 13 11 13 10 9 11
14 1 3 9 10 9 0 13 7 3 9 13 1 10 11
22 0 3 13 13 11 7 10 10 9 7 10 9 0 13 13 10 9 1 10 9 10 0
14 15 13 7 11 10 11 7 0 13 13 9 1 10 9
16 1 3 10 1 11 9 13 11 3 0 13 1 0 3 3 13
5 0 3 0 13 13
23 13 3 10 11 10 9 13 1 11 9 13 16 10 0 13 0 13 9 1 11 1 10 9
33 13 3 1 15 13 10 11 10 9 13 0 13 1 9 7 13 9 13 12 9 13 16 15 3 13 3 13 10 9 16 3 13 15
11 10 3 0 16 3 15 13 11 9 7 13
11 11 13 13 1 9 0 9 13 3 0 9
11 9 3 15 13 11 13 3 9 10 0 9
5 3 3 15 3 13
22 13 3 13 1 10 9 15 15 3 13 3 7 13 15 10 0 7 15 15 3 3 13
15 1 10 9 7 13 7 3 9 15 13 3 10 0 9 13
7 15 3 15 10 9 13 13
25 11 3 3 3 13 13 3 7 9 0 13 7 11 13 7 13 7 12 7 12 9 7 13 10 9
26 0 3 13 16 10 9 10 9 11 11 13 13 15 1 0 13 0 13 1 11 16 15 9 10 9 13
25 13 3 13 16 13 10 9 10 9 10 13 10 0 10 9 9 7 10 1 9 9 0 0 13 11
24 10 3 11 3 13 13 3 11 13 10 9 0 7 13 3 11 13 3 3 13 15 10 0 9
29 0 3 1 11 11 13 13 1 9 10 7 15 7 3 11 10 11 15 9 13 1 10 9 11 13 10 0 9 1
7 11 3 0 3 13 3 13
31 13 3 15 1 9 13 10 9 10 9 7 10 1 11 13 0 13 7 10 11 9 16 13 11 7 7 13 10 9 13 0
28 13 3 10 9 15 1 10 9 10 9 13 3 1 10 9 12 9 11 3 1 0 13 7 10 9 7 13 13
9 10 3 12 9 13 10 9 15 11
7 11 3 11 10 11 3 13
7 3 3 0 0 13 3 13
11 13 3 10 9 1 10 11 3 13 13 0
13 3 3 13 0 10 9 15 3 7 10 0 9 9
15 7 0 3 15 3 13 13 7 9 3 13 9 13 1 0
13 15 3 3 3 13 15 7 13 9 7 3 3 11
5 0 3 3 11 13
4 0 3 0 13
30 10 3 9 0 11 3 13 7 13 10 0 13 3 7 13 10 0 9 9 13 13 11 1 11 13 9 10 10 0 9
14 3 3 13 0 0 13 13 7 15 1 11 13 9 13
18 16 3 9 0 10 9 13 9 7 10 0 7 9 10 0 13 10 9
30 7 15 13 0 15 13 16 3 13 15 7 13 10 9 1 10 0 9 10 9 7 0 3 13 13 15 3 13 3 13
11 3 13 15 13 10 9 10 1 10 0 9
3 13 3 0
6 13 3 15 3 10 9
29 1 0 3 10 9 7 10 0 0 15 13 10 9 10 1 11 9 15 13 13 1 10 11 10 0 9 15 0 13
24 13 3 10 9 10 15 9 7 7 9 7 9 9 13 7 9 7 7 9 3 13 3 1 15
14 13 3 9 7 9 1 11 13 9 15 13 10 13 0
14 10 3 11 15 13 0 9 13 0 15 3 0 0 13
25 0 3 1 10 9 9 13 3 13 0 7 9 0 0 15 13 13 10 9 10 9 15 13 3 13
24 10 3 9 13 13 16 9 9 0 13 9 1 10 15 1 10 15 3 13 13 0 13 0 13
9 10 3 11 1 9 13 0 10 11
3 3 3 0
48 9 3 3 0 0 0 16 10 11 10 1 11 13 1 0 11 10 11 9 9 13 9 13 1 11 10 1 11 1 11 13 13 1 10 9 10 9 13 15 10 9 15 0 13 15 10 9 13
4 9 3 3 13
14 0 3 3 13 13 10 11 0 13 16 15 3 0 13
9 3 3 10 11 13 0 7 7 11
24 13 3 11 3 0 3 13 13 12 9 1 10 0 9 11 9 7 13 1 11 10 11 0 12
10 10 3 3 0 13 11 10 3 13 11
30 11 3 3 13 3 9 13 1 10 0 0 7 11 10 11 13 1 11 13 7 10 1 11 9 7 9 13 15 1 11
13 3 7 9 13 7 0 0 15 10 9 13 1 15
15 13 3 11 10 11 9 13 10 11 16 13 0 9 15 13
11 13 3 15 3 1 0 10 9 13 3 11
7 10 3 11 13 10 15 9
24 7 3 1 0 7 7 11 9 10 0 9 13 13 0 11 13 10 15 12 7 7 12 9 13
12 13 3 11 10 9 13 1 10 9 10 0 11
13 10 3 11 1 3 10 11 3 0 13 1 9 13
6 1 3 11 13 9 9
24 13 3 7 13 1 15 0 9 11 10 11 15 13 11 3 9 11 3 9 9 0 9 13 13
16 9 3 9 13 0 13 0 3 0 9 3 3 13 9 15 13
12 7 16 10 3 3 0 13 15 3 1 9 13
7 0 3 15 10 9 13 0
28 0 3 10 9 9 13 0 16 10 11 0 13 9 7 9 0 13 10 0 9 7 0 9 7 0 9 0 13
11 13 3 3 0 15 0 13 1 10 13 11
18 0 3 1 10 11 1 10 9 13 9 13 9 15 9 13 1 10 11
7 10 3 9 0 13 11 9
25 0 3 9 15 13 1 11 10 7 0 9 13 15 3 10 9 7 3 15 1 0 3 0 13 15
15 13 11 9 0 0 7 7 9 9 10 11 13 10 9 13
9 3 13 15 10 11 0 13 10 3
19 3 3 13 16 13 1 9 10 9 13 10 9 1 15 0 9 13 10 9
32 16 3 15 13 9 13 10 0 15 3 13 15 15 3 10 0 13 13 10 7 11 16 13 0 13 1 9 9 10 7 9 13
23 16 3 13 11 13 1 10 11 3 0 3 9 1 10 9 10 11 0 9 13 1 10 13
22 0 3 3 13 7 11 15 0 0 13 3 1 11 13 13 11 9 3 15 11 3 9
13 11 3 3 13 11 9 3 13 11 10 11 9 9
6 16 3 13 13 11 0
19 3 3 15 13 10 0 0 3 13 16 13 10 9 0 1 9 11 13 11
14 7 9 7 3 13 7 15 15 0 13 13 1 10 0
21 15 3 3 11 7 7 11 9 7 15 11 13 7 13 9 13 3 3 3 15 13
22 15 3 16 13 10 9 0 13 3 3 13 10 0 13 1 9 0 7 0 13 9 9
11 3 15 3 15 13 16 15 13 13 13 15
24 13 13 10 11 13 9 1 10 11 1 10 11 16 0 13 15 3 13 9 7 7 9 10 15
14 13 3 3 3 9 10 15 11 13 13 1 10 9 0
20 0 3 1 11 13 1 11 10 0 9 3 15 13 13 10 7 9 7 10 9
19 0 3 15 15 13 1 10 15 13 16 11 7 7 11 13 15 13 3 15
8 0 3 3 1 13 1 15 13
7 0 3 1 15 0 13 13
22 16 0 7 7 10 0 0 13 15 9 10 11 13 9 9 10 0 13 10 11 9 13
11 3 10 7 15 0 13 0 9 10 7 0
7 15 3 3 15 0 13 13
17 15 3 3 13 13 13 9 0 13 15 9 15 0 13 13 1 15
6 13 3 3 0 13 3
17 16 3 3 13 15 13 13 10 9 1 0 9 13 15 10 13 13
3 0 13 13
5 1 15 3 11 13
35 6 9 3 0 13 10 13 9 0 7 7 10 13 15 10 7 0 13 13 0 7 0 7 9 10 1 10 11 13 3 13 13 15 13 0
2 15 13
4 15 3 9 9
18 13 3 15 9 13 0 15 1 10 15 13 9 7 7 9 7 9 13
31 13 3 3 0 3 13 1 10 9 0 1 9 10 15 13 7 15 1 11 13 7 0 13 1 0 11 13 15 13 1 9
14 3 3 13 9 3 13 0 9 13 1 7 9 7 9
22 16 3 15 9 13 13 10 0 9 7 0 1 0 13 13 16 1 0 0 10 13 13
7 1 3 10 13 3 13 9
4 0 3 3 13
18 9 3 3 0 9 13 15 13 1 11 9 3 13 1 0 9 16 13
21 15 3 3 13 15 6 9 13 9 13 13 7 9 10 1 10 11 7 9 10 0
12 3 3 15 13 3 1 0 9 13 10 9 9
22 16 3 3 15 13 9 7 0 13 9 13 15 1 9 13 3 16 13 9 0 10 0
5 13 3 3 15 0
10 0 3 15 7 1 9 15 9 13 13
8 11 3 0 13 10 11 9 13
26 13 3 10 0 9 7 3 13 9 13 0 10 13 11 10 11 9 13 11 15 3 7 0 13 13 0
22 15 3 6 9 13 1 9 13 0 0 3 9 15 1 9 7 0 7 1 9 13 13
10 15 3 15 13 0 15 15 0 13 13
12 13 13 10 11 13 9 1 10 11 1 10 11
17 7 3 3 13 15 7 1 9 7 3 1 9 13 7 3 1 0
6 10 3 9 13 13 0
4 3 3 15 13
22 7 16 10 9 13 7 13 9 13 1 10 11 7 3 13 10 9 0 3 9 13 0
30 15 3 15 9 0 0 0 13 7 15 3 15 0 13 13 9 16 9 15 13 11 10 0 13 3 9 11 13 1 9
14 3 3 9 13 0 1 9 3 12 15 10 9 9 13
15 15 3 3 13 1 9 15 0 13 15 9 13 7 15 13
6 3 3 10 9 0 13
14 3 3 3 15 13 13 1 15 13 15 15 13 13 0
8 10 3 3 13 9 0 13 13
11 16 3 3 13 15 13 13 3 15 0 3
7 13 3 1 10 9 10 9
6 0 3 15 15 3 13
6 10 3 0 15 15 13
15 13 3 16 1 9 10 0 3 7 9 10 0 13 10 9
8 13 3 10 9 10 13 15 13
24 3 3 3 9 0 1 0 13 1 0 16 15 10 9 13 9 13 7 9 1 15 13 3 15
10 3 3 13 13 0 10 9 0 3 15
13 13 3 3 15 9 13 9 1 15 9 0 13 13
7 15 3 3 0 6 9 13
17 15 3 6 9 11 11 13 13 9 0 1 9 3 13 0 3 13
9 0 3 0 1 13 15 15 9 13
4 3 3 3 13
4 9 3 13 0
11 1 15 12 3 13 10 13 1 3 10 13
16 10 3 3 13 13 3 13 13 15 3 13 13 16 3 3 13
12 7 16 3 13 3 3 1 10 9 0 13 13
8 9 3 0 1 9 10 9 13
20 15 3 15 13 10 9 13 0 15 13 7 9 15 13 7 13 9 15 15 13
16 16 3 3 15 13 10 15 0 13 1 3 15 3 15 16 13
4 11 3 0 13
5 11 3 13 13 0
6 11 9 13 10 15 9
22 7 15 0 10 9 13 13 0 7 0 7 13 15 1 10 11 3 7 13 1 10 9
10 15 3 3 1 15 15 3 13 0 13
58 3 3 13 1 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 13 3 13 0 3 13 16 16 15 9 13 7 3 0 7 3 3 13 1 10 15 16 13 13 10 13 1 0 15 11 7 13 7 13 1 10 11
23 3 13 0 3 13 7 13 7 13 13 9 16 7 0 15 1 9 7 0 15 1 9 13
5 0 3 1 0 13
11 3 3 9 7 13 7 11 13 10 11 9
14 9 3 9 13 3 13 15 3 9 13 13 1 10 11
11 13 10 11 9 15 13 0 7 7 0 13
15 3 3 13 6 9 9 3 13 1 10 11 13 13 9 9
10 7 3 13 13 3 7 10 13 15 13
8 15 3 0 13 13 10 11 13
9 9 3 13 9 3 0 9 15 13
8 9 9 9 15 13 16 0 13
18 9 7 3 1 10 15 0 3 13 7 10 13 0 13 15 9 15 13
7 9 3 16 13 0 13 13
12 9 3 13 3 10 0 9 10 11 13 13 13
24 6 9 11 7 3 13 1 9 7 13 10 9 7 10 15 9 1 15 13 9 3 1 15 13
4 3 3 0 13
10 16 3 3 3 13 0 15 1 15 13
16 16 7 0 7 0 13 1 0 9 3 3 0 3 1 9 13
6 13 3 15 13 11 0
6 1 3 3 0 9 13
9 13 3 0 15 13 13 15 15 13
7 3 0 3 13 0 13 13
14 13 3 3 7 13 13 9 13 15 3 13 13 15 0
5 3 3 3 13 13
27 16 3 9 13 10 13 7 15 3 1 9 13 13 9 1 11 13 3 15 10 0 0 9 3 3 15 13
28 13 3 3 3 13 0 16 13 10 15 9 15 7 13 1 0 13 1 10 15 9 7 3 1 9 10 15 13
16 0 0 6 9 1 15 13 13 7 3 7 10 13 0 13 13
26 15 15 3 0 13 9 0 9 13 3 3 10 15 0 9 9 9 13 9 13 3 13 9 10 15 13
48 15 3 13 1 15 3 3 0 13 9 15 9 12 13 9 15 3 9 13 15 3 13 7 13 16 0 13 13 10 9 0 15 13 3 13 10 13 0 13 9 16 10 0 15 7 7 9 13
25 3 3 16 13 1 10 0 13 15 13 10 1 9 9 13 9 9 15 9 3 13 15 13 10 9
7 7 7 0 13 6 9 0
17 9 3 10 1 9 13 0 13 15 15 15 13 9 15 0 0 13
15 15 3 10 1 15 9 0 10 9 3 10 3 13 1 9
20 16 3 3 3 13 0 0 15 15 13 7 15 10 0 13 15 15 0 13 13
30 3 3 3 1 0 3 9 13 0 15 15 3 3 13 0 13 15 1 10 9 16 13 15 13 15 13 10 15 9 13
27 16 3 15 3 1 15 9 13 7 13 13 7 16 10 15 9 13 7 16 10 15 7 13 0 3 13 13
12 16 3 3 13 3 3 13 3 3 0 0 13
28 16 3 15 3 13 13 7 3 15 7 15 13 7 3 13 15 1 9 15 13 13 0 1 15 13 13 3 15
7 1 3 0 10 13 9 13
11 0 13 11 13 11 13 13 15 13 10 13
27 13 3 10 11 9 7 13 1 10 0 9 16 1 0 9 13 13 15 13 10 0 9 15 3 1 11 13
5 13 3 10 11 13
9 11 3 15 13 13 13 0 0 13
15 0 7 13 11 10 9 13 7 0 9 13 15 13 10 9
54 15 3 6 9 3 9 13 3 0 7 7 0 13 9 1 0 3 13 15 10 15 10 9 13 13 3 0 13 10 0 13 13 3 10 1 9 11 9 3 13 13 3 3 10 1 9 10 11 13 3 3 11 1 9
11 13 0 9 13 13 15 0 13 1 15 9
23 16 3 0 15 13 9 7 9 3 13 13 15 9 0 15 3 3 0 13 7 10 9 13
10 15 3 13 3 9 10 1 10 9 13
11 13 3 13 10 1 15 0 13 1 10 9
27 0 3 13 3 13 10 9 16 9 13 3 11 7 13 0 9 7 11 15 0 13 0 13 3 13 0 13
5 10 3 9 13 0
24 13 10 11 13 9 9 1 3 10 9 10 9 9 15 13 3 3 13 1 10 9 13 10 9
42 13 3 0 10 9 9 7 10 13 3 15 9 1 10 9 15 13 13 9 15 1 10 13 13 0 0 10 13 9 13 7 11 10 9 3 9 13 9 15 13 10 9
17 1 3 11 9 1 3 12 9 0 13 9 7 7 10 0 10 9
8 0 3 9 13 13 9 0 9
14 0 10 15 3 3 0 1 0 13 9 12 0 3 0
11 15 3 13 15 9 3 13 1 10 0 9
5 15 3 3 9 13
24 15 3 9 13 15 3 0 9 3 13 15 3 1 10 9 0 9 13 15 3 9 7 7 9
21 7 0 3 3 13 10 0 13 1 10 11 13 1 12 9 3 3 10 1 10 11
7 1 3 11 10 11 13 9
9 3 3 13 13 1 9 0 10 9
3 9 3 13
13 11 3 10 11 7 11 10 11 9 9 13 10 9
15 10 3 11 13 9 0 7 7 0 1 9 13 13 1 9
16 3 3 13 1 10 9 10 9 0 7 13 7 9 3 12 9
14 1 3 10 9 0 1 15 13 10 11 11 9 0 13
18 15 3 1 11 3 3 10 11 13 15 3 10 9 0 1 0 13 13
8 13 3 0 11 11 11 11 11
7 9 3 0 15 10 11 13
22 0 3 13 10 3 13 9 0 3 13 1 9 15 3 3 13 0 16 13 1 10 3
6 0 3 13 7 7 13
14 10 3 3 0 1 9 13 10 9 10 9 9 0 13
17 3 3 10 7 3 9 7 10 3 10 0 9 13 13 15 0 13
22 13 3 9 15 15 13 13 10 3 3 9 10 9 13 0 3 15 13 0 10 9 13
6 13 3 10 9 13 3
10 3 7 3 13 7 13 10 15 10 9
9 9 3 15 0 13 1 10 11 13
18 3 3 15 13 13 9 1 15 11 13 13 13 7 9 13 7 9 13
16 10 3 0 0 15 3 3 10 9 13 3 10 11 9 13 13
5 0 3 3 3 13
33 13 3 3 9 1 10 9 0 7 7 9 13 9 7 7 0 7 9 10 9 13 16 3 13 10 9 7 10 9 13 1 10 11
11 10 3 3 0 1 0 9 13 10 11 13
22 15 3 1 11 10 0 15 3 1 11 0 3 1 11 10 1 11 15 3 1 11 13
18 15 3 3 10 9 9 0 13 13 10 13 1 9 13 9 3 13 13
9 7 3 9 1 9 0 1 13 13
44 0 3 16 13 10 11 9 13 10 11 1 15 13 13 1 11 3 9 13 11 9 7 0 3 0 3 11 15 9 13 13 11 15 1 15 10 9 10 11 13 1 10 11 13
18 1 3 3 10 10 9 11 9 13 15 1 9 9 13 1 11 13 13
28 1 0 10 9 13 11 10 11 9 9 13 10 9 9 15 0 0 7 0 11 9 7 13 13 1 10 9 13
20 13 3 9 11 13 11 9 10 13 15 7 13 9 11 7 15 9 13 13 0
17 6 9 0 13 15 15 10 9 11 13 10 9 10 0 7 10 9
15 13 3 10 9 10 0 11 0 0 13 11 15 15 13 9
3 15 3 13
18 6 9 7 15 13 7 13 10 3 13 10 15 9 7 13 15 3 13
37 16 3 3 15 13 1 9 13 10 0 13 15 13 1 10 9 9 13 7 13 13 9 3 12 9 13 15 9 9 3 0 9 9 0 13 12 9
5 7 0 15 15 13
11 0 3 15 1 9 7 7 9 13 13 9
4 15 3 0 13
12 15 3 7 13 3 9 10 15 7 9 0 13
8 15 3 15 1 15 9 0 13
36 9 7 15 13 15 7 10 12 9 15 10 9 13 1 15 13 10 12 9 16 3 15 0 13 10 12 9 12 9 7 13 15 9 1 15 13
12 13 7 0 15 3 0 13 13 7 13 3 0
13 3 3 15 0 13 7 1 10 13 7 1 9 13
10 0 3 13 7 0 13 13 10 3 3
18 11 3 13 9 9 13 7 9 1 15 9 13 13 1 11 9 0 11
9 1 15 11 9 1 9 9 13 13
29 1 3 11 10 9 13 1 10 9 10 9 7 9 13 1 11 9 3 9 13 13 3 1 11 13 1 9 10 9
21 13 3 1 11 0 3 13 9 1 10 11 13 9 7 7 9 7 13 9 9 13
15 3 7 1 11 7 1 11 13 1 9 9 10 3 0 3
11 0 3 1 10 0 13 1 9 7 7 9
12 15 0 3 13 11 13 0 3 13 3 13 13
7 13 3 0 0 13 3 13
8 1 3 0 13 3 13 1 11
13 15 3 1 0 10 11 13 1 10 11 1 10 11
21 1 0 3 10 9 1 11 13 13 15 13 10 3 9 9 10 3 0 10 0 0
9 13 3 12 9 1 11 1 10 3
14 7 3 13 10 9 13 9 0 13 7 0 15 7 13
20 16 3 13 11 0 13 10 11 13 12 13 9 9 7 13 1 10 9 9 9
12 3 3 13 16 3 9 1 0 13 13 10 11
9 13 3 3 13 13 0 7 7 0
16 6 0 9 9 15 9 13 0 16 15 13 15 1 0 0 13
15 15 3 1 9 3 15 9 13 3 13 7 0 7 0 9
11 7 15 3 0 13 15 13 0 10 0 9
5 15 3 15 9 13
40 13 3 3 9 7 9 13 1 3 10 1 10 0 11 12 7 7 12 1 3 10 0 12 7 12 10 3 11 0 10 3 11 1 9 16 13 10 9 10 9
32 13 3 9 13 0 15 3 1 10 11 10 0 10 9 1 10 3 13 10 3 0 1 9 7 7 10 0 9 7 7 9 1
24 9 3 9 13 10 9 7 9 16 7 1 10 9 13 10 13 13 9 0 7 1 10 11 3
26 0 3 13 13 1 9 13 9 0 10 9 3 3 0 13 7 12 3 9 13 1 0 12 3 10 0
22 16 3 13 10 9 9 9 13 7 13 0 10 9 10 9 9 13 1 10 9 10 9
6 13 3 3 3 3 13
25 13 3 15 10 9 13 10 1 10 9 9 0 13 7 0 13 9 7 10 3 1 9 7 9 13
18 13 3 7 13 0 10 11 0 13 7 13 10 9 15 13 13 10 9
19 15 3 13 16 9 13 10 9 9 10 9 13 9 13 9 9 9 3 15
9 0 13 10 11 0 13 13 10 9
23 16 3 13 10 9 11 10 9 13 10 1 10 9 9 13 7 10 9 13 1 11 13 0
19 11 3 15 3 13 15 13 3 15 13 13 7 13 7 3 13 13 15 13
8 15 3 16 0 13 13 13 0
17 6 9 13 15 9 13 12 7 15 13 15 1 15 13 1 10 11
8 3 7 13 10 11 7 13 0
35 6 0 9 15 13 15 13 0 1 10 11 7 13 9 15 7 9 7 0 7 9 13 1 15 9 13 15 9 15 13 9 0 10 9 13
26 3 3 0 13 16 1 10 9 10 9 13 10 9 15 0 3 13 9 13 10 9 0 3 0 13 13
13 16 3 3 0 13 0 0 13 9 9 3 13 13
11 15 3 3 7 10 12 10 9 13 10 0
9 10 3 12 15 13 3 10 9 13
38 16 3 0 13 3 13 15 13 0 13 10 11 9 13 10 0 0 13 13 3 10 9 13 15 3 1 0 10 9 15 3 1 0 7 3 13 10 9
9 13 3 0 0 1 0 13 10 9
35 13 3 3 9 12 1 9 15 13 3 3 9 12 7 0 1 15 13 10 9 3 1 10 9 13 3 3 0 0 13 9 12 13 3 0
6 0 3 13 9 1 0
9 13 9 0 10 0 15 9 13 11
16 1 3 0 10 12 9 9 11 0 13 15 9 3 13 0 12
11 1 3 3 10 9 13 3 9 13 10 9
9 15 3 3 1 0 10 9 9 13
9 0 3 1 0 11 1 9 9 0
12 13 3 15 9 15 9 13 11 11 9 9 9
11 13 3 16 15 9 13 1 10 9 1 9
16 15 3 1 9 9 10 0 7 7 0 12 1 9 10 9 13
10 1 3 10 9 1 10 0 9 13 0
3 0 0 13
18 7 0 12 3 1 10 9 1 10 9 9 13 0 7 3 13 10 15
9 10 3 12 1 0 13 0 9 13
18 13 3 0 9 3 10 1 10 9 13 10 9 7 9 10 3 13 11
7 10 3 0 13 9 9 0
32 13 3 10 9 1 10 11 10 9 1 7 9 11 7 9 10 0 1 3 11 13 11 9 13 1 0 1 10 11 1 11 9
12 10 11 3 13 1 0 9 13 1 10 11 9
21 7 0 3 15 1 10 11 9 13 9 7 7 9 13 7 15 3 3 0 9 13
13 13 3 7 13 0 0 10 11 10 0 13 9 12
7 9 3 10 9 10 9 13
9 0 3 13 9 9 1 10 9 13
26 1 9 3 13 3 1 0 3 13 11 9 7 11 7 11 15 3 3 11 0 13 1 0 3 11 0
12 16 3 13 1 11 0 13 11 13 15 10 9
14 3 16 13 13 1 10 9 13 7 10 0 7 10 9
8 13 3 13 10 9 9 13 13
15 16 3 13 7 7 13 9 0 13 7 10 9 7 10 9
26 16 3 13 15 3 10 11 1 10 9 13 15 3 10 9 7 10 9 9 0 9 3 10 11 15 13
4 1 3 0 13
12 6 9 3 0 15 13 13 3 7 7 0 0
4 13 3 15 13
3 15 3 13
4 15 3 13 13
7 0 0 1 10 9 13 0
28 1 3 3 0 9 15 3 9 13 0 13 7 0 7 10 0 15 3 13 3 7 3 3 13 13 3 3 13
18 10 7 3 9 13 7 10 9 13 3 0 13 0 13 13 13 10 9
13 3 10 3 9 0 13 10 9 9 0 10 9 13
12 10 3 9 0 13 10 9 0 1 15 13 13
4 11 3 13 13
22 11 9 3 3 0 1 13 0 15 3 15 13 13 13 7 0 13 0 13 9 1 9
1 13
4 0 15 3 13
4 15 3 13 13
12 6 9 9 3 10 13 10 9 3 13 0 13
27 15 3 3 3 1 0 9 13 0 7 1 15 15 7 0 13 7 3 3 13 15 12 10 0 15 13 0
6 11 3 1 0 13 0
9 0 9 15 0 13 13 12 15 0
18 16 3 15 3 13 0 13 10 15 9 9 3 0 15 10 0 9 13
16 6 9 7 9 0 15 3 9 13 13 3 7 10 9 10 9
13 16 3 0 13 10 12 15 15 13 0 3 0 13
9 10 3 12 0 13 9 7 7 9
24 3 3 10 9 13 9 0 3 3 15 13 15 13 9 13 15 0 10 0 0 13 13 10 9
17 3 3 12 0 13 13 10 9 7 1 15 10 9 1 15 3 13
12 7 3 10 12 15 10 0 13 10 0 13 13
18 16 13 15 15 0 13 0 15 13 0 15 3 13 3 10 3 3 13
7 9 3 3 13 9 15 9
20 9 3 3 3 13 0 16 13 3 13 15 13 13 9 1 3 10 9 0 13
3 13 11 0
8 11 3 3 15 3 0 0 13
8 3 7 15 13 7 15 3 13
17 16 3 3 13 1 10 3 13 9 10 15 3 13 13 3 0 15
21 16 3 13 1 15 10 13 3 10 0 13 13 13 1 15 3 3 10 0 0 13
6 0 3 3 1 0 13
8 13 3 9 13 3 13 10 0
11 10 3 13 13 3 10 3 13 13 10 9
10 10 3 13 7 15 7 13 3 3 13
8 13 10 9 9 1 15 9 13
30 16 3 0 10 1 15 13 9 9 13 0 3 15 7 3 13 9 0 15 9 13 0 3 3 3 13 15 1 0 13
7 0 3 9 0 9 13 13
26 15 3 13 0 9 7 10 9 0 13 7 13 15 10 11 13 3 7 9 13 3 7 15 0 15 13
8 0 3 3 0 0 9 13 13
13 0 3 15 3 3 13 9 7 9 0 10 9 13
4 13 11 1 0
12 6 9 16 13 15 13 9 15 3 15 9 13
9 3 3 13 1 0 9 0 9 13
12 0 3 10 9 13 15 15 9 13 1 10 9
11 3 3 1 0 0 3 13 10 0 0 13
14 7 3 15 16 13 13 0 13 13 10 9 7 0 13
9 0 3 3 13 15 9 0 15 13
11 0 3 13 0 3 13 3 10 15 9 13
4 13 1 0 11
18 1 3 0 1 10 15 13 9 7 9 7 9 3 13 13 0 15 13
10 15 3 15 0 1 15 9 10 15 13
13 0 13 7 11 13 1 11 0 13 11 9 10 0
7 16 3 15 13 13 15 0
33 6 9 0 15 15 13 13 9 7 13 0 7 3 13 10 3 13 9 13 0 7 7 0 0 7 12 7 0 7 10 0 9 13
6 0 3 15 0 0 13
8 0 3 1 13 13 10 9 3
8 0 3 10 9 13 1 10 9
35 16 3 13 10 9 13 1 0 9 11 1 10 9 13 1 10 9 15 15 9 0 13 15 15 13 13 10 11 0 3 1 9 10 0 13
17 13 3 13 10 9 1 10 11 7 0 9 7 0 9 15 9 13
27 0 3 13 3 13 7 16 10 9 13 13 1 10 9 7 16 13 15 10 11 13 7 1 0 10 9 13
34 16 3 0 15 13 13 1 3 10 0 10 9 10 1 10 11 10 0 7 7 10 9 0 1 3 10 1 10 0 10 9 7 10 9
5 0 3 10 9 0
14 10 3 0 0 3 10 7 9 7 10 10 9 3 13
4 13 3 3 0
6 1 3 0 10 0 9
8 7 10 9 3 13 1 10 0
8 3 3 13 3 0 13 9 15
13 11 3 16 13 1 10 11 13 10 9 1 9 13
15 13 3 10 9 15 1 12 9 7 1 12 9 13 15 9
10 3 13 11 3 13 10 11 9 13 0
21 6 11 15 3 9 13 9 7 9 1 11 11 13 0 10 11 13 13 13 15 9
8 3 3 1 0 13 15 13 0
4 9 3 13 9
27 0 3 0 0 13 16 13 3 13 9 1 10 11 11 3 7 3 3 3 1 15 13 13 1 10 0 9
9 13 3 3 0 15 9 13 1 11
13 9 3 13 9 0 13 9 10 3 0 10 3 0
6 3 3 13 10 10 0
14 10 15 9 15 13 10 3 13 1 3 15 10 0 9
15 10 3 0 1 10 11 13 1 9 13 10 0 13 10 0
18 15 3 3 1 9 13 1 0 9 13 10 9 1 15 15 13 13 13
11 10 3 11 13 10 11 9 7 7 9 0
7 1 3 15 13 9 0 11
27 1 15 9 7 13 0 0 15 3 11 13 7 9 9 1 15 13 1 11 1 0 10 9 16 1 9 13
17 13 3 10 11 10 9 13 0 13 7 7 13 10 9 7 13 0
29 10 3 3 9 10 15 13 1 11 10 9 13 11 1 10 9 10 0 11 13 1 15 11 7 0 13 9 7 9
6 13 3 3 11 9 0
8 10 3 9 0 10 0 13 9
12 15 3 1 10 11 0 10 9 10 9 9 13
6 3 3 13 1 0 9
13 0 3 10 9 10 0 10 9 13 12 7 12 9
5 13 3 0 10 9
16 13 7 1 12 9 9 9 7 13 0 3 3 13 13 3 9
17 13 3 7 13 10 12 9 13 1 10 9 9 13 9 1 10 9
15 0 3 13 15 13 1 10 13 16 15 15 0 10 9 13
5 10 3 13 0 13
4 9 3 3 13
4 3 3 9 13
21 9 3 0 13 9 3 0 9 3 0 3 3 9 1 10 0 9 13 1 10 9
10 7 9 13 11 10 11 9 10 11 9
15 13 3 3 1 3 9 9 1 3 15 0 7 10 0 9
26 16 3 11 10 11 7 7 11 13 1 11 10 11 7 13 15 10 9 11 13 15 9 15 9 13 11
8 13 3 0 13 10 11 0 9
6 1 0 3 10 9 13
7 9 3 10 0 0 13 13
9 10 3 9 9 3 13 11 9 9
6 13 3 3 1 15 9
16 13 3 11 10 0 1 11 1 10 9 0 13 3 0 10 9
6 0 1 15 3 13 9
14 9 3 3 3 9 13 9 13 11 10 11 0 0 13
13 0 3 1 3 9 13 0 1 3 10 9 0 13
4 0 3 1 0
6 13 3 15 11 10 11
15 9 3 10 9 1 3 10 9 9 1 0 13 0 13 13
3 9 3 13
11 9 3 0 7 9 3 3 3 9 9 13
8 10 3 9 15 10 9 13 9
13 0 3 7 9 13 11 10 11 7 7 11 10 11
15 9 3 9 3 13 1 9 13 9 3 0 13 7 9 0
4 3 3 9 13
6 13 3 3 13 3 9
13 9 3 9 3 13 13 0 10 3 15 3 3 0
6 9 3 13 11 10 11
4 0 3 13 0
7 11 3 7 0 11 10 11
5 9 3 11 10 11
7 0 3 7 11 11 10 11
13 0 3 9 7 13 7 9 0 0 13 7 9 13
10 0 3 3 13 9 13 11 10 11 9
11 9 3 1 9 13 13 9 3 7 9 0
11 9 3 0 7 13 7 9 0 13 7 9
7 11 3 9 13 11 10 11
12 9 3 7 9 7 7 9 13 13 3 3 9
4 0 3 13 0
7 9 3 7 9 11 10 11
5 9 3 11 10 11
5 0 3 9 13 13
12 1 3 9 13 9 0 13 15 3 10 9 13
4 3 3 9 13
9 3 3 9 9 13 0 13 9 9
5 13 3 3 9 0
16 10 3 9 10 3 0 13 9 13 1 9 10 3 15 0 9
27 0 3 7 9 10 1 11 13 13 11 10 11 7 11 10 11 9 15 3 13 10 9 11 9 0 0 13
10 10 3 3 1 11 9 7 0 13 11
24 10 3 1 9 9 9 0 3 3 13 13 10 9 13 9 3 15 10 0 9 3 7 9 0
10 10 3 1 10 11 0 9 13 15 9
14 0 3 10 1 10 11 9 10 3 0 3 3 9 13
15 0 3 9 13 1 10 9 1 7 10 9 13 7 10 9
7 7 1 3 9 10 9 13
8 10 3 9 10 9 0 13 13
7 9 3 1 9 13 9 9
11 9 3 9 3 0 13 13 9 3 0 13
6 9 3 13 11 10 11
21 9 3 3 7 9 11 10 11 13 9 3 7 9 7 0 11 10 11 7 7 11
9 9 3 3 10 0 9 13 0 13
15 10 3 9 3 9 13 13 9 9 15 0 13 0 13 9
14 13 3 1 10 11 1 10 9 3 10 9 13 1 9
9 0 3 3 3 9 13 13 9 0
7 0 0 13 11 11 13 9
7 9 3 3 10 0 13 9
11 1 3 11 10 11 13 10 9 13 10 9
4 9 3 13 0
5 0 3 13 9 0
6 1 11 3 9 13 9
14 9 3 7 9 13 11 10 11 15 1 11 13 1 11
38 9 3 1 3 10 9 9 13 13 1 3 10 9 9 3 3 9 13 0 1 3 10 9 7 7 10 9 9 9 3 3 9 7 7 9 7 9 0
20 0 3 13 3 1 10 11 13 9 10 3 0 13 3 0 13 0 13 1 11
10 9 3 10 1 10 11 13 11 10 11
11 1 3 10 9 9 7 7 9 13 9 0
6 10 3 9 9 0 13
7 1 0 10 9 11 13 9
23 9 3 10 9 0 3 13 10 0 9 13 9 15 15 16 1 10 9 9 13 13 3 13
9 9 3 9 7 0 13 7 9 13
14 13 3 15 9 15 0 1 3 10 9 1 9 13 9
14 9 3 1 3 10 9 9 0 13 9 3 7 9 0
4 9 3 13 0
11 9 3 7 9 7 9 3 3 9 13 13
19 9 3 1 3 10 9 9 0 9 3 0 0 9 7 0 3 3 9 13
8 9 3 7 9 13 11 10 11
9 0 3 7 9 3 3 9 13 13
6 0 3 11 10 11 13
19 0 3 10 9 13 11 10 11 15 1 11 13 0 9 0 13 1 10 9
13 0 13 10 1 9 13 7 9 7 13 1 10 0
23 0 3 10 9 13 3 0 15 3 13 7 10 13 7 13 0 13 7 9 7 7 9 13
6 9 3 7 9 10 9
8 13 3 3 0 15 3 13 9
54 13 3 0 7 7 10 0 9 10 0 11 7 10 11 7 11 10 11 10 9 13 3 13 1 11 7 11 10 11 11 0 0 9 9 11 3 13 9 7 11 10 11 7 7 11 9 7 11 10 11 7 11 10 11
9 0 13 9 10 0 0 1 10 12
8 13 3 0 10 9 0 1 0
22 16 15 15 13 10 9 7 9 13 7 9 0 9 13 7 13 0 7 0 12 7 0
11 9 3 0 13 1 15 9 7 0 0 13
7 9 3 0 13 15 3 13
23 3 3 9 7 0 7 0 13 13 9 7 3 13 3 3 9 7 9 0 7 7 3 13
5 13 3 0 10 9
8 3 3 15 13 9 7 0 0
13 3 1 10 9 13 15 15 7 0 7 0 13 9
12 13 3 15 9 9 0 13 9 3 0 3 9
11 9 3 1 13 13 10 7 0 7 10 0
5 15 13 3 9 12
11 9 3 3 13 13 7 0 7 0 1 9
6 13 3 9 13 1 9
7 10 3 9 0 10 9 0
13 15 3 3 13 16 7 9 16 7 9 1 15 13
6 15 3 1 9 13 13
10 0 3 0 10 9 7 13 1 10 9
12 9 3 10 3 1 10 0 13 9 7 0 3
11 9 3 9 3 13 10 0 3 1 10 0
5 13 3 9 7 9
9 1 3 10 9 13 9 7 9 0
6 13 3 3 0 15 9
12 3 3 3 0 7 0 13 3 3 1 10 0
11 0 3 9 3 13 10 0 3 1 10 0
8 13 3 15 9 9 3 13 9
5 0 10 9 0 13
13 9 3 10 9 13 12 9 1 10 9 7 10 9
8 10 3 3 15 9 13 1 9
4 0 3 0 13
9 9 3 13 11 7 7 11 11 9
10 10 3 0 15 9 11 13 1 11 13
9 16 3 13 1 11 1 9 13 0
23 13 3 15 1 10 9 10 9 13 9 7 10 9 3 13 13 7 7 13 0 13 10 11
11 13 3 9 7 13 7 1 9 13 10 9
9 10 3 9 3 1 9 13 3 13
18 13 10 9 1 10 9 1 15 3 13 10 9 1 10 9 13 10 9
6 11 3 3 13 10 9
11 9 3 1 9 10 1 10 11 12 3 13
23 1 3 10 9 9 13 3 13 9 10 0 13 3 9 0 9 3 9 3 13 13 7 9
14 0 3 10 9 10 0 13 3 0 13 1 10 0 9
9 3 3 13 10 11 13 10 1 9
13 10 3 11 0 10 9 7 10 1 11 15 11 13
5 0 3 9 13 12
23 0 3 13 1 3 10 9 9 0 9 3 0 10 9 0 13 7 9 7 0 7 9 0
4 9 3 0 13
9 0 3 13 9 12 7 12 13 3
8 10 3 9 13 9 10 9 15
5 10 3 15 13 9
6 10 3 15 3 3 9
5 0 3 0 9 13
26 15 3 1 11 7 11 15 3 1 11 15 3 1 11 15 3 1 11 15 3 1 11 3 10 0 13
20 0 3 3 1 3 10 9 9 0 9 3 13 1 9 0 13 7 9 0 13
12 12 3 9 0 7 9 13 3 10 0 9 13
10 1 3 11 10 11 9 9 13 10 9
8 9 3 12 13 9 0 9 13
13 10 3 9 0 13 10 1 11 13 1 11 7 9
10 0 3 13 9 12 0 7 13 7 0
25 13 3 9 0 7 9 0 0 7 9 3 3 9 9 1 10 9 13 1 3 10 9 9 9 13
7 0 3 9 13 1 11 13
10 1 3 11 10 11 9 0 13 10 9
17 9 3 10 1 10 11 12 13 9 13 7 0 9 7 13 1 11
7 10 3 15 3 3 9 13
6 13 3 7 9 7 9
11 0 3 15 0 13 1 10 0 10 9 13
8 9 3 12 9 13 13 3 9
4 7 0 0 9
15 0 3 0 13 1 10 0 9 3 10 9 9 10 1 11
17 9 3 12 9 13 13 7 3 9 7 10 3 13 9 3 9 9
5 13 3 13 3 9
11 13 3 1 15 10 9 9 7 9 7 9
10 0 3 0 13 13 9 9 7 9 0
24 0 15 7 10 1 10 0 13 15 13 0 0 9 15 15 3 3 9 13 1 9 9 3 13
11 13 3 3 3 9 7 3 10 15 13 9
19 3 9 3 15 10 15 13 9 7 9 10 9 0 15 15 13 9 13 15
36 10 3 0 13 11 7 10 11 7 11 10 11 7 11 10 11 7 11 10 11 10 3 0 7 7 0 9 11 10 11 7 9 7 10 11 9
9 0 3 13 11 11 13 1 15 9
7 10 3 0 9 13 10 12
53 10 3 13 1 3 10 9 0 13 0 0 11 11 7 0 11 11 7 0 11 11 7 9 11 11 7 0 11 11 7 0 11 7 10 11 7 11 10 11 7 9 11 7 10 11 7 11 10 11 7 11 10 11
21 10 3 3 0 3 13 9 3 3 13 11 3 15 3 9 13 1 10 11 13 9
21 9 3 3 13 15 11 9 3 13 11 9 3 1 11 10 1 9 10 3 3 9
14 13 3 9 7 7 0 7 0 7 7 0 12 9 13
19 7 0 10 9 1 3 10 0 9 0 13 15 7 10 9 9 0 9 13
19 15 3 13 9 13 15 10 9 13 15 13 0 9 3 0 10 3 15 0
7 1 3 0 10 0 9 13
14 11 3 16 13 7 7 13 10 9 13 0 15 13 13
16 7 13 10 9 16 1 0 1 0 13 7 10 9 7 10 0
28 10 3 9 10 9 13 15 7 12 9 1 10 9 13 10 9 1 9 13 15 3 7 13 10 9 3 1 9
10 15 3 1 10 9 13 13 7 10 9
19 16 3 7 0 13 7 13 1 10 9 13 11 10 11 13 15 1 10 11
5 13 3 15 13 0
10 11 3 15 15 0 15 13 13 15 13
24 15 13 9 7 7 3 15 13 15 7 7 10 0 9 10 15 1 9 13 9 7 0 7 0
11 3 3 15 0 13 16 9 13 9 15 13
4 15 3 0 13
4 15 3 13 13
8 9 3 9 13 1 15 7 9
14 15 3 15 9 13 13 13 15 15 0 13 3 0 13
7 16 3 0 13 11 13 0
35 9 16 9 13 3 13 0 13 15 3 13 15 0 1 15 13 10 11 9 3 3 3 0 13 9 3 0 13 1 7 9 13 7 9 0
11 15 13 10 11 10 7 9 13 7 10 9
12 13 3 3 15 9 10 1 0 10 0 9 13
13 9 3 1 3 13 15 15 13 0 13 0 3 13
17 16 7 3 13 13 12 0 13 15 16 7 0 0 16 7 3 0
5 0 13 11 13 13
9 11 15 13 9 9 12 9 0 13
1 13
2 13 15
8 15 13 0 10 9 9 0 13
9 15 3 13 3 3 1 9 12 13
30 16 3 0 7 13 7 9 0 15 15 7 7 15 1 15 13 9 1 9 13 0 13 16 3 9 10 9 0 13 13
2 3 13
4 13 15 10 13
23 3 3 13 12 7 3 0 7 3 12 13 3 0 15 3 7 3 1 12 13 9 0 13
13 3 3 0 1 12 0 13 3 12 13 0 12 9
27 1 3 3 12 13 1 9 10 15 13 3 13 0 3 1 10 15 9 0 7 13 13 9 1 0 0 13
10 13 3 1 10 0 3 3 13 0 15
17 7 1 15 3 0 0 13 15 15 13 13 3 3 3 0 7 0
6 15 15 13 0 0 13
4 1 0 11 13
11 6 9 3 13 16 9 13 3 0 15 13
13 15 3 16 13 13 10 9 10 0 13 10 13 9
25 3 16 15 13 10 3 0 13 0 0 3 13 15 15 9 7 7 9 13 0 9 7 7 9 13
10 9 3 15 13 9 7 15 7 9 13
18 15 3 7 12 9 13 0 7 13 13 7 12 0 7 13 3 3 13
25 16 3 9 13 7 0 15 10 13 9 13 3 15 3 12 0 10 9 15 9 0 13 12 0 13
7 0 3 13 3 15 0 13
14 13 3 15 9 9 15 13 0 3 3 3 10 15 15
6 13 3 15 3 0 13
5 13 3 10 0 3
16 3 13 13 15 9 9 1 9 7 13 1 10 9 13 7 13
4 3 7 13 13
6 13 3 1 9 15 9
5 15 3 3 0 13
31 0 3 1 9 13 11 7 9 1 10 11 0 13 11 10 11 10 3 1 11 13 13 13 10 9 1 10 11 1 10 11
15 13 3 3 0 0 10 9 9 1 10 11 7 10 11 3
21 0 3 15 10 7 1 11 7 10 11 1 10 1 11 1 9 0 0 10 9 13
11 10 3 1 11 11 0 3 13 13 0 13
19 10 3 13 1 9 15 9 11 13 13 9 0 3 3 11 0 10 1 11
21 0 3 13 3 13 7 10 13 15 1 9 9 13 3 16 3 0 9 0 13 11
30 15 16 13 1 0 7 11 10 11 13 15 0 13 7 13 1 10 11 3 13 16 9 13 13 9 7 13 1 10 0
30 16 3 15 3 9 13 1 10 9 13 9 0 13 10 9 7 10 9 7 10 9 7 10 9 7 3 13 1 10 9
8 13 3 0 15 13 1 10 9
11 3 3 0 3 13 3 3 1 0 1 9
9 11 3 1 10 11 13 1 10 11
22 13 3 3 3 0 15 13 10 1 11 15 7 13 1 9 0 11 7 13 7 0 11
20 13 3 13 1 11 0 3 10 0 9 15 0 13 1 9 9 15 9 13 11
6 13 3 0 0 9 11
20 1 3 15 10 0 11 9 13 15 3 3 13 10 9 13 10 11 9 7 13
11 10 3 9 0 3 3 13 11 3 3 11
15 13 3 10 11 9 10 9 13 9 0 0 13 11 11 11
32 0 7 3 13 7 1 0 9 0 0 11 3 1 7 11 13 11 1 3 11 11 1 15 9 12 13 10 9 11 7 7 11
28 1 3 0 10 9 13 10 0 9 13 15 1 12 9 13 13 3 12 9 3 3 10 9 0 7 7 3 0
6 0 10 9 0 13 13
7 10 3 9 0 9 13 11
15 0 3 3 10 9 10 0 7 7 0 1 0 9 13 13
17 9 3 9 1 15 10 9 9 13 0 9 9 9 0 0 9 9
28 0 15 3 1 9 13 1 10 9 13 10 3 15 10 0 13 13 3 1 15 1 9 10 15 15 3 13 13
16 13 7 3 9 0 9 7 0 7 9 0 7 13 10 0 0
31 10 3 9 0 13 3 1 10 9 10 0 9 3 10 9 13 10 13 10 9 9 3 10 13 3 3 1 11 7 15 0
20 13 3 10 11 10 13 0 0 13 9 10 9 15 12 11 13 9 7 0 11
39 3 3 3 1 0 10 9 10 9 13 1 0 9 10 11 9 13 13 0 7 7 0 1 15 0 7 7 0 13 9 15 13 9 7 7 9 7 3 9
39 13 3 10 11 1 11 9 9 9 7 7 9 13 13 1 9 16 15 13 1 9 7 11 7 9 11 15 3 0 13 13 11 15 3 0 0 0 9 13
32 10 3 9 0 10 1 10 11 9 13 11 13 10 3 1 9 1 9 11 13 1 10 11 10 3 1 9 13 1 0 10 11
8 1 15 10 9 13 13 9 0
24 13 3 0 1 10 9 7 15 0 1 0 1 12 9 10 9 13 1 10 9 10 11 13 13
8 0 3 7 10 1 0 13 11
56 3 3 9 10 1 11 1 0 9 13 13 1 11 9 13 11 9 0 13 7 13 1 11 3 13 0 0 10 9 7 10 1 10 11 9 13 3 3 15 0 13 10 3 1 9 13 13 1 9 13 10 3 1 9 3 13
21 10 3 9 0 15 9 11 10 9 13 7 13 9 7 13 13 7 3 10 1 15
33 16 3 3 1 10 11 13 9 7 10 11 10 0 13 7 13 15 9 0 13 7 13 7 15 0 13 1 10 9 7 10 9 13
5 13 3 15 10 9
13 0 3 10 11 13 0 1 9 3 9 13 10 9
8 9 3 3 11 13 11 13 9
20 10 3 13 9 10 9 7 13 11 1 15 0 13 3 16 0 1 10 9 13
20 11 3 7 10 0 9 13 1 10 11 10 0 13 10 9 13 1 10 11 13
27 13 3 1 10 0 7 0 1 9 11 15 1 0 13 13 1 11 9 7 13 1 10 9 10 1 11 9
12 16 3 1 10 11 13 10 11 13 3 10 9
39 13 3 10 9 3 13 10 1 9 9 0 13 1 11 9 7 10 11 1 11 7 9 7 11 15 13 9 10 0 7 7 0 1 10 0 9 10 9 13
9 13 3 3 1 0 10 9 10 0
17 10 3 13 0 9 1 0 13 11 0 3 13 10 9 13 7 13
13 10 3 3 9 3 13 7 7 13 13 1 10 11
17 10 3 9 9 1 10 9 1 10 9 10 9 0 13 1 11 9
26 13 3 7 13 16 15 10 9 13 13 1 10 9 13 0 1 11 10 9 13 3 15 13 0 13 13
11 3 3 15 13 12 1 0 7 11 10 11
4 15 3 1 13
7 10 3 11 13 15 13 0
14 0 9 0 0 9 3 10 0 13 13 13 7 9 13
5 9 3 10 9 13
6 0 3 10 11 13 0
9 3 1 3 10 0 13 10 9 15
20 9 3 13 9 13 0 3 10 9 13 16 3 15 10 9 13 1 0 10 9
24 3 3 9 13 13 16 3 15 13 1 10 13 0 15 9 1 10 9 16 10 0 13 0 0
15 10 3 9 10 1 10 11 1 10 13 1 10 9 13 0
7 1 3 9 13 1 10 0
17 1 3 9 15 13 13 7 3 13 15 3 13 12 9 0 3 12
10 3 0 13 10 1 11 15 13 10 9
40 3 3 10 0 13 3 13 10 9 10 9 7 13 3 1 10 9 13 3 15 13 0 13 7 10 9 1 13 9 13 1 10 0 9 16 3 3 13 3 0
7 0 3 0 0 0 1 13
5 13 3 0 13 13
7 9 0 9 11 0 15 13
18 15 13 9 13 1 15 15 13 9 11 10 11 13 1 10 11 9 11
6 3 3 3 13 15 9
23 7 3 15 9 1 10 15 9 13 7 15 0 13 15 0 13 7 1 15 0 9 13 13
15 13 3 0 3 0 10 9 13 15 9 0 9 0 13 0
20 13 1 11 10 0 13 0 9 1 9 0 11 7 10 11 7 10 1 0 13
32 0 3 10 0 0 9 13 3 0 1 11 9 13 11 10 11 16 15 3 13 13 15 1 11 9 13 7 13 1 15 13 0
39 16 3 3 11 7 13 0 13 9 1 11 7 0 9 13 1 11 13 11 1 9 3 13 3 13 7 15 9 1 15 13 0 3 3 15 3 0 0 13
31 13 3 0 16 16 15 9 10 0 0 1 0 13 13 13 10 0 13 3 1 10 10 3 0 3 0 15 13 3 15 13
6 3 3 3 0 0 13
33 3 3 0 13 16 3 0 13 10 13 10 9 1 10 11 16 15 1 10 0 3 10 9 13 15 3 13 15 13 1 10 13 9
19 1 3 10 11 15 7 13 9 1 10 9 13 11 7 3 3 1 0 11
17 10 3 11 0 9 9 10 1 11 13 1 9 11 10 1 11 13
13 15 13 11 1 0 7 10 1 11 7 11 3 13
21 1 9 3 15 10 9 13 9 10 0 9 13 13 11 12 15 10 9 13 9 0
16 0 3 10 11 13 1 11 13 15 9 9 7 0 0 10 9
12 3 3 15 13 7 0 13 0 3 3 13 13
16 0 3 3 0 13 13 16 15 3 10 9 15 9 10 9 13
19 10 0 3 9 3 1 10 15 9 13 13 7 1 9 7 0 7 9 0
7 0 3 3 13 0 10 9
23 13 3 11 10 9 10 11 13 11 10 9 9 0 1 0 7 11 10 11 15 13 9 11
13 1 3 3 0 9 1 9 13 15 10 9 13 9
30 13 3 11 9 7 7 0 7 0 7 7 9 7 3 0 7 7 10 9 0 9 13 1 0 10 9 13 10 11 0
6 0 3 13 11 10 0
53 16 3 3 11 13 0 9 10 9 11 13 13 1 9 11 13 1 10 9 3 3 10 11 10 9 13 10 11 9 11 7 7 11 3 13 10 9 0 3 13 10 9 16 13 9 10 9 13 0 13 10 11 9
13 10 3 9 10 10 0 13 11 13 10 9 7 15
17 15 3 16 13 10 11 11 3 13 9 0 13 13 15 11 9 15
11 15 3 10 11 13 7 13 15 15 10 11
8 15 3 3 3 7 13 7 13
11 10 3 3 0 0 1 10 11 13 9 13
5 11 3 10 9 13
29 9 3 10 1 11 16 13 1 9 13 10 3 15 0 13 7 9 15 7 13 13 1 0 13 1 10 11 9 13
11 10 0 3 0 3 9 10 1 11 13 13
10 13 3 0 0 0 13 9 13 9 0
8 0 3 9 9 13 0 10 11
17 3 3 16 10 9 10 9 13 1 10 11 13 15 1 9 13 0
12 13 15 0 7 10 0 9 13 15 1 10 0
46 15 3 13 1 10 11 3 3 13 16 9 9 13 13 10 11 7 13 15 10 0 9 1 10 11 13 1 10 11 9 3 13 16 1 11 13 1 9 3 13 15 10 11 1 15 13
15 0 3 3 13 15 10 0 9 0 13 7 0 13 10 13
5 13 3 15 15 13
12 10 3 3 13 9 9 3 10 3 0 13 13
4 15 3 0 13
6 11 3 0 13 13 0
13 9 9 9 13 0 13 15 9 1 10 0 13 13
57 0 3 15 0 13 0 9 13 16 15 1 0 9 13 13 7 10 11 10 11 1 0 9 13 13 7 10 9 13 1 15 15 0 9 7 7 9 13 7 15 1 13 13 7 10 11 9 13 10 7 1 15 0 0 1 9 13
9 7 3 3 15 7 1 10 0 13
15 3 3 16 13 10 9 7 13 1 15 3 3 11 9 13
11 9 3 0 10 9 9 16 3 13 13 13
12 1 0 3 9 7 3 0 13 7 3 15 13
9 0 13 7 13 10 11 13 7 0
17 3 3 0 13 10 9 11 13 9 10 9 13 1 11 7 7 0
17 1 0 10 11 16 13 13 10 9 10 11 10 0 15 0 13 9
10 6 9 9 9 13 9 13 13 10 9
15 15 3 13 9 1 10 9 3 15 13 0 1 10 9 13
14 7 16 15 10 9 3 0 13 15 15 13 10 0 9
12 7 7 0 15 0 13 13 7 13 9 0 0
5 11 3 3 0 13
10 13 3 10 0 9 10 0 13 15 0
14 6 9 0 3 9 13 10 11 13 15 1 15 7 9
12 15 3 16 3 9 13 3 13 10 11 3 13
5 16 3 13 15 13
27 15 3 3 15 10 9 9 13 13 13 15 10 0 9 13 13 16 10 9 0 15 13 13 3 1 15 13
10 3 16 10 9 13 15 13 15 15 13
7 0 3 3 13 13 3 13
5 0 3 13 15 13
27 3 3 3 3 0 9 9 0 13 13 16 0 13 0 13 10 9 0 3 9 13 0 3 13 3 9 9
16 15 3 11 10 9 9 0 13 1 9 13 13 7 7 13 9
8 3 3 9 15 15 13 13 0
3 13 11 0
27 16 3 15 13 13 10 15 13 3 3 13 10 0 3 13 7 13 10 11 16 1 10 9 10 9 15 13
9 0 3 10 9 10 9 15 13 13
11 10 3 3 10 9 9 0 10 11 13 13
35 11 3 1 0 13 3 1 10 9 16 3 13 10 0 13 0 3 7 3 0 13 13 1 11 13 1 0 13 11 9 0 3 10 9 13
4 15 3 0 13
56 16 3 0 13 10 9 13 10 11 13 9 12 11 10 11 9 0 1 11 13 9 0 7 0 9 13 10 9 3 13 7 16 3 10 0 13 10 7 9 15 13 7 9 7 7 9 15 13 10 11 16 3 10 9 3 13
47 10 3 11 0 0 0 13 1 9 9 0 3 13 0 7 13 7 0 13 15 7 1 9 1 0 0 13 10 9 13 1 11 3 1 0 13 7 7 13 9 11 10 1 11 13 10 9
15 15 1 10 0 0 10 1 15 13 3 0 3 0 0 13
36 13 3 0 9 15 15 11 13 13 13 3 13 7 16 10 9 13 10 9 7 11 13 13 7 3 3 0 13 1 10 11 3 15 10 9 13
9 11 3 13 9 11 15 9 13 11
28 3 3 3 0 13 16 13 10 0 9 1 7 10 11 11 7 11 13 11 10 0 7 1 11 10 9 10 9
27 10 3 11 0 13 1 9 3 3 0 13 7 1 9 0 16 10 9 7 13 7 16 13 10 9 13 13
8 7 3 13 7 13 13 3 9
6 10 15 3 13 13 11
7 1 0 3 13 13 10 9
20 10 3 11 1 0 10 9 13 1 10 9 13 7 13 1 9 0 9 0 13
16 13 3 9 10 15 13 16 13 13 10 0 13 15 1 10 9
4 3 3 13 13
15 0 3 9 13 1 15 10 9 10 0 1 0 7 0 11
5 10 3 1 11 0
8 0 3 0 13 10 9 0 13
18 15 3 3 3 13 13 7 7 13 13 16 3 15 13 13 10 11 13
13 16 3 13 15 3 15 15 3 13 10 0 10 9
6 7 13 13 1 10 0
4 13 3 3 0
9 16 3 13 13 15 13 13 9 12
10 13 3 3 16 13 1 10 9 13 0
33 6 9 15 13 10 9 15 1 10 9 0 13 9 3 0 7 9 0 13 3 7 0 1 3 0 3 13 15 13 7 15 0 13
8 15 3 3 3 13 3 15 13
12 1 3 10 9 15 9 13 15 3 3 3 13
22 13 3 10 9 16 3 13 13 13 3 12 9 1 3 9 9 13 11 3 0 3 13
11 3 3 13 1 11 7 15 9 13 10 9
6 0 3 3 13 10 9
12 9 3 16 15 13 10 1 0 13 9 13 0
4 10 3 11 13
9 0 10 9 16 13 13 13 10 9
16 13 3 11 1 9 11 13 1 11 10 3 11 13 13 0 9
29 1 3 9 9 9 15 13 15 1 9 7 7 0 13 9 0 1 11 13 1 9 12 9 11 15 1 15 0 13
12 9 3 3 13 7 13 7 13 9 13 13 13
14 16 3 1 11 13 13 13 15 9 0 13 1 10 9
12 13 3 10 9 15 3 15 3 9 1 11 13
14 3 11 9 13 13 7 7 13 1 3 9 13 9 0
6 0 3 9 3 13 9
26 10 3 11 9 13 11 9 11 13 0 15 3 13 1 11 7 11 10 9 13 13 1 11 10 0 9
13 7 10 3 1 9 7 7 9 10 9 15 9 13
15 1 3 10 11 13 3 13 0 13 15 7 9 7 3 9
18 0 3 9 1 11 13 13 10 0 1 15 3 0 13 13 9 0 11
11 10 3 3 11 13 0 13 13 13 10 9
17 9 3 1 9 10 0 13 3 13 16 3 15 13 15 10 9 13
16 16 3 13 0 13 13 10 9 1 10 11 13 1 10 9 9
9 13 3 1 0 10 9 10 9 13
20 9 9 13 13 10 9 10 0 16 11 7 7 10 0 13 11 1 9 10 9
6 15 3 3 0 13 13
16 13 3 13 3 15 9 0 16 16 3 13 13 15 13 10 9
14 3 3 15 13 0 1 10 0 11 0 1 15 13 13
11 13 3 3 13 9 15 15 0 3 13 13
6 0 3 9 9 0 13
7 15 3 13 0 15 9 13
8 16 3 13 10 9 13 1 11
43 13 3 10 11 1 11 13 13 1 11 10 9 3 13 7 13 1 10 11 1 10 9 15 3 1 11 10 3 1 11 13 1 9 11 1 3 11 7 9 13 7 10 11
14 3 13 10 9 1 12 9 13 7 15 13 10 9 9
22 13 3 0 3 11 10 11 1 10 9 13 9 3 13 3 10 9 0 3 11 10 11
5 13 3 0 9 3
32 13 3 9 1 11 10 11 9 9 13 15 13 7 13 1 10 9 13 1 10 9 10 13 13 10 9 7 10 9 7 10 9
18 16 3 0 15 0 13 0 3 13 13 7 15 0 13 13 10 9 13
12 13 3 10 9 1 10 9 3 13 1 10 9
20 9 3 13 9 3 3 13 3 7 3 3 16 1 10 9 13 9 9 13 0
23 10 3 9 16 13 1 10 9 13 1 10 13 1 11 3 7 13 10 9 7 1 15 9
10 10 13 3 9 13 10 1 11 9 13
12 0 3 13 13 15 1 11 7 3 0 10 15
23 0 3 13 13 10 9 3 13 1 10 11 10 0 10 3 0 9 13 9 10 11 1 11
4 0 3 10 11
11 1 3 10 0 10 11 3 10 11 13 9
4 3 3 11 9
17 10 3 11 10 3 1 9 9 0 7 7 0 0 13 1 10 11
11 10 3 1 10 9 10 9 9 13 7 9
19 13 3 1 10 9 0 0 9 15 11 13 10 0 7 9 13 11 1 15
13 13 3 9 1 0 10 9 7 10 3 0 9 13
18 13 3 9 10 9 13 16 9 13 1 9 13 9 10 0 15 3 13
18 10 3 3 9 10 0 1 0 7 13 7 10 0 15 3 1 9 13
12 10 3 3 13 13 3 13 1 10 11 10 0
8 9 3 13 3 10 9 11 9
10 10 3 3 9 0 10 9 13 13 0
23 15 3 13 7 13 16 7 9 13 13 10 0 7 9 3 15 13 13 10 13 1 10 11
25 16 3 13 10 9 13 1 11 13 1 10 9 13 15 15 3 1 11 3 15 3 1 9 1 11
8 10 3 3 9 1 9 13 13
7 0 3 0 13 10 11 9
26 9 3 13 10 9 0 3 9 10 13 13 0 13 10 13 15 7 15 3 13 10 0 13 9 0 13
34 1 3 0 10 9 10 9 9 7 13 1 11 3 3 10 11 9 11 10 9 13 1 15 3 10 9 0 10 9 13 7 9 15 13
12 9 3 3 1 10 9 3 3 3 10 9 13
10 13 3 0 10 9 10 9 1 9 13
35 10 3 3 0 15 13 11 3 13 13 10 9 7 3 10 9 15 10 13 13 1 10 9 10 9 13 0 13 15 13 10 9 0 7 0
7 10 3 13 0 9 13 11
21 10 3 0 15 13 11 3 15 15 9 13 11 10 11 13 9 0 13 0 10 9
13 15 16 10 9 13 1 0 13 13 16 15 13 0
35 16 3 13 3 13 7 13 0 10 9 15 3 13 1 10 9 1 9 10 0 13 15 1 0 13 9 7 13 10 9 7 9 0 9 13
16 7 15 16 3 13 1 10 15 9 13 13 15 10 9 13 3
12 10 3 15 15 13 1 10 9 0 13 3 9
26 10 3 0 15 13 11 9 0 13 13 1 10 9 10 11 7 10 3 9 13 10 9 10 3 9 3
16 16 3 3 0 13 10 9 10 0 13 1 11 13 13 1 11
22 13 3 7 13 1 10 11 13 1 11 13 3 10 11 13 3 0 1 10 0 10 11
21 10 3 12 9 10 9 12 13 1 10 9 10 1 13 11 7 7 11 13 3 11
34 3 10 0 16 9 9 13 13 1 10 9 13 0 1 11 16 15 10 3 13 0 13 15 10 9 12 9 13 1 10 9 9 1 11
11 10 3 9 15 13 13 1 9 3 11 0
24 0 3 13 10 0 13 10 11 9 1 11 7 7 10 9 10 1 11 7 9 13 7 0 9
64 1 3 3 0 10 9 7 11 0 7 0 13 10 9 7 9 13 3 3 3 15 13 13 10 3 1 10 9 10 1 10 11 13 12 7 12 7 12 10 3 0 0 10 9 13 9 12 7 12 9 7 1 9 7 7 12 3 1 0 9 13 1 0 9
13 0 0 9 13 12 7 12 7 3 12 7 7 12
10 13 3 0 10 9 3 3 0 13 12
11 3 3 9 3 13 1 15 12 9 7 12
15 0 3 3 10 1 10 11 0 13 0 13 12 9 7 12
12 9 3 13 1 0 12 7 3 9 12 7 9
13 10 3 0 12 7 12 9 13 10 3 9 12 9
18 13 3 3 0 10 9 10 13 0 7 0 10 9 9 9 13 12 9
29 7 3 10 7 1 10 9 7 10 0 9 13 13 12 7 9 7 12 7 12 7 3 9 12 7 9 12 7 9
4 9 3 13 13
20 9 3 3 10 1 11 9 7 10 1 10 9 10 13 10 11 13 12 7 12
11 1 3 3 0 10 9 9 12 7 12 13
45 0 3 15 9 13 7 9 7 9 7 0 7 10 0 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 7 0 7 15 10 11 10 0 13 0 10 9 12 9 13 13
22 0 3 10 9 0 13 10 1 10 11 13 10 15 9 10 0 9 12 7 12 7 12
7 13 3 0 9 12 7 9
40 10 0 3 0 13 9 0 10 9 10 13 0 7 10 1 10 0 9 13 7 3 1 10 0 9 10 1 13 10 9 0 10 0 9 3 13 13 0 7 0
13 3 3 15 13 0 0 13 7 7 0 7 0 15
26 3 12 7 9 7 12 7 12 7 9 12 7 9 12 7 9 12 9 13 11 10 11 1 11 7 11
9 0 3 3 10 0 10 11 9 9
12 9 3 0 7 9 7 9 15 3 13 0 9
24 3 3 9 7 7 10 0 9 10 0 7 9 0 10 13 3 3 0 1 9 15 3 13 9
22 3 15 15 9 13 13 10 9 10 9 13 15 7 3 3 10 9 13 9 15 9 0
28 13 3 13 16 9 9 0 10 9 13 7 15 0 12 9 9 13 1 9 0 7 3 12 7 0 9 7 12
10 9 3 7 9 7 9 7 9 3 13
20 9 3 13 0 9 9 7 1 7 9 15 15 0 13 0 11 13 0 10 9
30 1 3 9 1 9 7 7 9 10 9 13 13 15 9 7 0 7 0 9 9 15 3 9 13 10 1 0 10 9 13
29 15 3 3 15 13 13 10 9 7 15 3 13 9 15 3 13 10 9 13 10 9 7 0 7 13 7 10 9 15
7 15 3 1 0 10 11 13
10 15 3 1 11 9 15 3 1 11 13
6 13 3 10 9 9 0
18 13 3 9 16 0 10 9 1 9 13 13 15 0 9 10 9 9 13
12 9 3 1 10 9 9 13 9 0 11 10 11
13 16 3 3 1 0 10 9 13 9 13 3 13 13
19 1 0 10 9 9 15 0 13 13 12 3 0 9 7 0 9 7 9 0
15 3 11 10 11 9 9 13 1 11 3 10 9 0 13 0
11 7 15 3 10 15 3 13 9 0 0 13
9 13 3 15 3 0 0 9 13 0
11 0 3 9 7 10 0 9 13 3 13 9
19 3 13 10 9 10 0 9 16 15 13 13 10 9 9 0 1 10 9 13
31 9 3 0 7 13 7 13 9 10 9 10 9 1 7 0 7 10 11 7 10 9 13 13 0 9 7 3 3 0 13 13
6 15 3 3 0 9 13
24 15 3 16 13 11 9 13 7 9 13 10 0 3 13 1 10 11 13 0 15 15 0 13 9
20 15 3 3 10 0 13 1 10 11 13 11 9 9 1 0 3 7 1 0 13
35 13 3 9 1 10 9 0 10 11 3 13 10 9 13 1 11 7 7 10 9 1 10 11 1 9 13 16 1 10 9 13 1 11 10 0
8 3 3 13 13 1 10 9 13
8 1 0 3 10 9 9 13 11
19 12 3 10 9 0 13 7 0 0 13 7 3 13 10 1 11 10 9 9
14 13 7 3 10 15 13 10 0 7 13 13 1 10 0
26 15 13 10 1 11 10 0 9 11 10 11 15 3 0 0 9 11 1 9 0 13 13 13 10 0 9
17 13 3 15 13 10 11 13 15 0 0 10 9 13 1 9 10 0
15 13 3 0 10 11 7 13 16 0 0 3 0 13 13 13
12 3 3 1 10 9 13 13 3 10 0 13 13
16 16 3 15 13 13 10 9 13 15 10 13 9 13 3 15 13
19 10 3 3 0 10 10 9 9 1 10 12 9 15 13 11 13 13 1 11
38 11 3 7 10 0 13 1 11 7 11 13 13 3 3 0 1 9 1 11 3 9 13 9 10 7 15 13 7 10 11 9 13 16 0 13 10 1 9
7 3 3 10 0 9 13 0
15 10 3 3 1 11 9 11 0 3 13 10 9 10 9 13
48 1 11 3 10 11 13 11 10 9 10 9 13 10 15 13 13 15 0 9 10 1 10 0 10 0 11 3 11 10 11 13 11 9 1 11 13 3 3 3 1 9 0 13 10 0 9 9 0
15 15 3 13 10 9 0 0 0 13 13 10 11 0 9 13
7 11 3 13 10 9 10 0
12 3 13 7 13 9 15 13 7 3 1 9 13
33 0 3 13 10 11 10 11 9 9 16 9 10 9 13 0 1 9 11 10 11 7 13 15 13 13 0 10 11 1 11 10 0 13
11 13 3 0 10 13 1 15 9 10 9 13
9 0 3 10 1 11 7 10 1 11
22 1 3 0 10 9 13 1 10 11 1 9 9 1 15 9 7 7 9 1 15 9 13
16 1 3 10 9 9 0 7 0 13 15 10 11 9 0 9 13
22 0 3 3 9 13 1 10 9 13 1 11 11 1 15 11 9 13 1 9 1 9 13
18 3 3 3 0 13 15 10 9 0 1 10 9 1 9 1 15 11 13
9 12 7 3 7 12 9 10 9 13
14 10 3 9 15 13 10 9 10 0 13 9 1 9 11
12 1 3 10 9 11 9 13 1 10 9 10 9
21 13 3 0 11 9 3 0 1 9 10 11 15 1 10 9 0 13 1 10 11 13
7 1 3 10 11 9 0 13
10 1 3 10 11 9 12 9 13 1 11
17 9 3 3 11 13 10 11 1 10 0 10 3 3 9 1 10 9
18 13 3 10 9 0 1 3 10 0 9 11 1 3 10 0 7 0 11
8 13 3 3 0 1 0 10 9
25 13 3 15 3 10 1 9 9 13 15 1 11 15 3 10 1 9 7 9 13 10 1 0 10 9
37 13 3 0 9 10 13 10 9 1 0 10 9 9 7 12 9 7 9 7 9 12 0 0 1 11 7 10 11 12 7 12 7 1 10 0 11 12
3 0 3 9
11 1 3 11 12 7 1 11 12 7 0 12
50 0 3 15 10 9 13 13 1 9 16 0 3 13 0 10 0 10 3 0 10 9 0 15 13 9 10 9 7 15 13 1 9 1 0 7 13 7 9 7 10 1 10 0 9 13 7 15 13 0 15
11 3 3 9 13 10 13 1 10 11 7 9
18 13 3 0 15 7 13 15 0 1 9 13 3 13 10 3 0 15 0
13 13 3 3 10 13 3 13 0 1 10 9 13 3
8 15 3 0 13 13 1 10 11
10 0 13 3 3 3 15 9 1 9 0
59 10 3 13 3 7 15 10 9 13 0 13 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 10 11 13 10 9 1 11 1 0
16 0 3 15 13 0 9 11 7 7 11 13 10 9 1 10 9
12 0 3 13 0 11 9 7 3 3 13 11 9
16 15 3 13 1 11 13 9 7 10 13 12 7 15 13 9 13
16 13 3 13 3 0 15 1 10 9 13 13 15 13 11 10 11
15 0 3 1 0 9 13 11 0 9 13 16 15 3 13 13
18 13 3 1 10 9 13 13 7 13 7 3 13 1 10 0 10 9 9
4 15 3 13 13
23 0 3 10 1 11 0 13 9 16 0 13 10 15 9 13 7 3 0 13 16 15 13 13
19 3 3 11 3 15 13 3 13 13 7 9 13 1 10 11 1 9 13 3
13 3 13 1 9 3 13 10 1 11 9 13 10 0
6 0 3 3 3 13 13
16 10 3 1 11 9 16 3 13 10 9 10 9 13 13 1 9
14 10 3 3 0 0 13 13 1 11 10 9 13 1 9
30 11 3 9 7 9 13 10 9 0 3 7 13 13 13 7 9 1 10 9 13 15 13 3 13 15 0 9 10 9 13
14 0 13 15 13 11 9 9 13 15 13 7 15 15 13
24 13 3 3 13 1 11 16 13 13 3 9 0 7 10 9 16 13 0 7 7 11 13 9 9
16 10 3 3 13 10 9 15 13 13 1 9 3 0 3 13 13
8 13 3 0 10 9 0 3 13
12 15 3 3 13 13 10 9 15 3 10 9 13
8 0 3 13 13 7 10 9 13
8 13 3 15 3 13 3 1 9
8 7 3 15 13 9 7 13 0
9 13 7 13 1 11 15 3 13 15
6 7 15 0 3 13 13
8 13 11 10 11 13 1 10 9
3 15 3 13
14 13 3 3 0 15 16 13 1 10 11 1 10 9 0
12 13 3 9 15 13 13 3 3 13 13 9 0
11 15 3 10 9 13 1 15 9 9 0 13
4 13 3 3 3
6 9 3 15 13 3 13
9 16 13 13 10 9 3 10 9 13
22 13 3 16 0 3 7 10 13 1 11 13 13 15 15 9 9 15 15 9 13 9 13
20 3 7 3 11 0 13 10 13 13 7 0 13 15 9 0 13 10 15 9 13
3 15 3 13
16 6 9 15 13 3 9 9 16 3 0 3 3 13 3 15 13
6 0 13 3 13 10 11
30 0 3 16 3 13 7 15 13 9 7 7 9 13 13 13 1 15 9 7 7 0 13 13 15 13 13 1 9 10 15
11 16 3 13 13 1 10 9 10 9 13 0
9 15 3 13 7 3 13 3 3 13
18 0 3 13 15 15 7 3 3 0 9 16 0 3 9 13 0 3 9
10 16 3 10 9 3 13 3 0 3 13
18 10 3 9 13 13 15 0 13 9 15 13 11 3 3 0 3 3 13
36 16 3 3 0 13 10 9 15 0 13 10 9 10 0 7 10 0 3 1 0 7 9 13 7 9 0 13 3 3 10 9 7 3 13 9 13
10 10 3 0 13 13 9 7 7 9 13
9 15 3 3 13 13 0 13 10 9
7 13 3 13 9 0 10 9
8 13 3 3 0 10 9 3 0
18 16 3 15 13 13 10 9 10 9 13 7 1 9 7 3 13 13 3
4 3 3 3 13
8 10 3 0 10 0 15 0 13
18 10 3 9 1 9 7 7 1 9 13 13 7 1 9 0 13 1 9
9 0 3 1 10 9 13 13 10 9
12 16 3 15 13 0 10 9 3 10 0 13 13
42 13 3 9 15 15 13 10 13 9 11 10 9 9 9 13 15 1 9 15 0 15 1 9 13 13 13 7 10 9 15 1 10 9 13 1 11 7 13 10 3 13 9
21 0 3 13 0 13 1 11 7 15 13 1 10 9 10 9 1 10 11 13 9 13
12 9 3 0 13 3 1 11 13 1 11 9 0
6 13 3 1 0 15 0
32 13 3 0 13 9 16 11 7 10 11 9 0 7 11 9 13 10 13 1 9 0 10 9 7 13 10 9 10 9 3 15 0
29 0 3 3 0 13 13 16 10 10 9 9 13 3 1 11 7 7 11 9 7 1 11 10 0 3 3 10 0 13
8 0 3 13 11 0 10 9 13
29 13 3 3 3 3 13 3 9 0 10 9 11 16 10 9 0 13 13 7 11 3 13 10 13 10 9 1 10 9
3 0 0 13
18 11 3 16 13 15 13 10 11 13 3 0 13 13 11 7 15 13 11
8 13 3 1 9 9 1 10 9
9 1 7 0 3 13 13 15 0 9
6 13 3 3 10 9 0
11 13 3 1 10 11 9 10 1 10 9 13
12 9 3 10 9 0 7 10 9 10 0 13 11
9 13 3 10 11 0 1 9 10 9
28 13 3 1 7 11 9 0 13 10 0 1 10 0 7 1 11 7 13 9 7 1 9 9 3 3 10 0 13
29 1 0 3 10 9 7 3 13 10 9 10 11 13 13 15 10 9 1 0 3 13 9 10 0 1 0 3 10 0
11 9 7 3 13 7 15 13 1 9 10 9
9 10 3 3 3 9 13 1 15 13
11 10 3 1 10 9 9 9 9 13 11 13
7 13 3 15 10 9 3 13
11 13 3 13 10 9 10 9 15 13 9 0
4 13 3 3 9
26 9 3 13 0 3 9 13 9 13 1 10 9 3 7 13 10 9 7 13 10 9 7 3 10 0 13
9 16 3 13 9 13 9 1 9 13
8 13 3 15 15 13 0 13 9
28 10 3 9 16 13 10 9 0 7 7 0 13 13 1 10 9 10 9 13 16 1 15 13 9 7 13 3 13
5 0 3 3 0 13
12 10 3 1 11 7 11 9 9 3 15 9 13
7 15 3 13 10 9 1 9
22 10 3 1 11 9 0 3 10 9 11 13 1 10 0 13 10 13 13 1 9 15 9
11 3 3 3 0 13 10 13 10 9 10 9
5 0 3 3 9 13
9 3 13 10 9 7 15 13 10 9
3 15 3 13
13 1 3 0 13 15 3 13 7 13 1 9 0 13
8 15 3 15 1 11 13 3 13
11 13 3 3 16 0 15 13 11 16 13 13
17 15 3 7 9 10 13 3 13 3 13 10 9 1 15 13 13 9
12 13 3 15 9 0 13 7 10 11 9 3 13
9 0 3 15 1 9 0 13 13 3
27 15 3 6 11 9 0 7 0 9 0 1 9 9 13 7 15 3 3 1 11 3 9 13 9 13 11 9
4 11 3 13 9
10 3 15 13 13 16 0 0 3 15 13
23 0 7 3 13 11 7 13 9 13 0 9 13 10 9 3 3 9 13 3 3 13 10 13
45 9 3 15 7 0 3 0 0 1 13 16 3 10 9 15 13 10 9 0 11 10 9 13 13 10 3 1 11 0 13 1 10 0 10 13 15 13 0 13 11 13 16 3 13 15
7 15 3 13 0 3 3 13
12 10 3 3 9 10 13 13 7 13 7 13 11
8 9 3 7 0 13 0 1 0
9 0 3 0 3 0 13 7 3 13
5 13 3 15 11 11
16 11 3 16 9 13 9 13 13 9 1 9 3 3 9 9 13
6 7 3 13 1 11 3
21 1 3 10 9 10 9 0 7 13 7 0 10 9 0 3 3 10 9 7 7 9
7 10 3 3 9 10 9 13
11 15 3 1 10 0 9 13 1 10 0 13
11 3 3 13 1 10 0 13 9 0 10 9
16 3 3 10 9 10 9 13 9 13 15 9 3 1 10 3 13
8 0 3 3 0 13 0 1 15
6 13 3 9 15 10 13
25 3 3 13 10 13 15 13 9 1 10 13 10 9 13 9 15 13 0 1 10 0 13 7 7 13
7 15 3 10 9 13 10 9
26 7 11 3 1 0 10 9 13 9 13 0 7 0 1 15 0 9 15 15 3 9 0 13 13 10 9
6 13 3 3 0 10 12
10 3 3 9 13 3 15 7 0 7 0
18 3 3 3 3 11 12 9 11 7 7 11 1 10 11 9 11 13 11
18 15 3 13 10 9 11 10 9 15 10 15 13 3 0 15 13 0 9
34 11 7 3 12 9 3 13 13 7 1 10 9 10 11 9 7 7 0 9 13 0 16 15 0 7 9 10 9 13 7 13 10 0 3
12 16 3 0 13 13 10 9 3 3 13 10 9
24 1 7 3 10 0 10 9 13 3 7 13 10 9 13 13 1 10 9 15 0 10 15 1 0
15 10 3 9 13 1 10 9 3 3 10 0 9 13 1 11
13 0 3 7 9 0 13 3 13 9 0 13 9 11
4 0 9 15 13
37 15 3 3 13 0 13 1 9 13 10 9 9 16 15 15 0 10 0 9 13 16 13 10 9 10 9 1 9 13 1 15 10 9 7 3 1 9
14 1 3 0 13 13 0 12 9 11 7 7 11 11 9
21 13 3 15 3 3 3 3 13 7 10 0 13 3 1 11 13 13 13 9 13 0
9 9 3 0 12 13 1 9 9 12
10 0 3 3 10 15 13 10 3 9 0
11 6 9 13 0 16 0 13 10 0 9 13
8 0 3 3 0 10 3 9 0
23 9 0 0 11 15 3 9 11 9 13 13 9 15 3 11 13 3 13 3 13 11 9 13
16 9 3 3 7 9 3 3 10 10 9 9 9 13 15 10 13
7 15 3 13 1 10 9 13
4 11 3 13 13
23 3 3 15 3 15 13 15 3 10 3 0 13 9 3 13 3 13 3 15 13 13 3 11
43 15 3 3 3 13 13 11 1 11 7 1 9 0 15 3 9 13 1 10 9 13 15 13 10 9 13 3 13 7 13 1 10 9 13 10 3 9 15 13 1 10 9 13
11 13 3 1 11 10 11 13 9 7 7 9
4 13 3 0 13
8 7 15 9 15 13 9 7 13
7 9 3 13 10 13 11 13
16 13 3 3 0 13 9 1 11 10 12 0 13 15 9 13 11
8 13 3 0 1 11 16 13 13
21 10 3 0 15 10 11 13 3 3 1 10 9 13 13 1 9 13 1 10 9 9
4 3 0 13 13
8 13 3 3 9 0 10 9 9
6 3 3 10 3 15 13
13 16 3 15 13 10 0 13 15 3 15 3 13 13
14 10 3 0 15 13 11 13 9 0 13 1 10 9 11
7 11 3 13 11 13 13 3
4 11 9 13 0
4 13 3 10 9
6 15 3 13 0 13 3
3 15 3 13
11 6 9 9 3 0 15 10 0 7 9 0
5 15 3 13 13 13
9 10 3 3 15 0 0 3 3 0
4 13 1 0 11
8 11 15 9 0 10 9 0 13
1 13
1 13
11 15 3 13 15 10 9 10 9 3 9 13
3 15 3 13
11 16 10 0 9 9 12 13 1 10 11 9
52 13 3 1 15 9 13 15 9 13 11 15 11 9 1 15 0 13 9 0 3 13 13 9 1 10 9 13 3 3 13 3 15 13 1 15 0 13 15 15 15 13 3 10 15 9 13 7 15 3 13 9 9
20 0 3 9 15 13 0 15 0 13 15 16 10 0 11 13 1 10 0 13 0
11 13 3 10 0 11 0 3 10 0 0 13
9 16 3 0 3 13 0 15 13 13
5 13 10 11 9 0
17 1 0 10 9 15 0 13 1 15 9 0 0 10 13 13 13 15
24 13 1 0 11 9 7 13 11 7 10 0 9 9 13 7 10 9 7 13 16 13 11 13 0
18 6 9 13 15 9 13 9 15 13 15 3 13 7 3 13 9 10 15
9 7 3 3 3 9 0 13 9 13
23 16 3 1 10 13 9 15 9 13 12 0 1 10 9 12 13 13 11 0 15 13 10 0
30 0 3 13 10 0 9 0 7 15 13 7 9 3 0 15 13 7 15 10 0 10 0 13 7 10 0 10 0 3 13
11 16 3 13 7 15 13 0 0 7 0 15
25 10 15 3 13 3 9 13 10 10 0 3 13 9 3 7 13 10 9 15 7 13 15 7 9 13
13 0 3 16 13 1 9 1 9 15 10 13 9 13
3 13 11 0
9 11 3 7 15 13 13 7 13 0
9 11 3 13 3 15 0 13 13 15
52 3 3 3 0 3 13 16 3 13 10 15 9 10 7 13 0 1 0 13 7 10 13 16 9 3 9 3 13 13 7 13 0 10 9 3 3 13 10 9 9 9 10 0 15 13 13 13 16 3 3 9 13
5 0 3 13 10 0
14 9 3 9 3 13 13 0 15 13 7 3 13 10 0
22 0 13 11 13 1 10 0 7 11 13 16 9 7 13 7 9 0 13 13 10 9 13
24 0 15 0 3 7 0 9 1 3 3 0 3 3 13 16 9 11 15 3 3 9 13 13 11
22 3 3 3 3 1 10 0 0 13 16 13 3 13 15 15 13 9 9 9 0 10 0
8 15 3 3 0 13 15 13 13
10 13 3 3 10 9 3 15 10 0 13
4 13 3 9 0
20 11 3 10 11 13 1 9 3 3 15 13 7 10 13 15 13 3 13 0 0
19 16 3 11 13 13 1 10 11 13 1 11 10 11 7 13 0 13 0 13
6 3 3 3 3 13 13
5 0 3 13 16 13
4 15 3 13 0
18 9 0 13 10 9 0 13 7 3 1 10 9 10 9 13 10 9 9
21 13 3 0 3 13 10 9 1 10 9 16 13 0 10 9 15 9 13 1 10 9
5 13 3 13 7 13
6 0 3 3 3 13 13
