485 11
6 13 16 13 13 10 0
4 13 16 13 13
7 3 13 16 13 13 10 0
7 9 1 9 7 9 1 9
10 16 3 13 10 13 15 12 15 9 13
30 7 15 13 9 3 13 0 15 15 13 0 15 16 13 10 9 15 1 9 7 9 15 15 13 1 9 13 15 1 9
8 9 15 15 1 9 13 9 15
9 7 16 13 3 13 3 10 0 0
5 7 1 9 15 13
4 13 1 0 9
20 3 15 15 13 15 9 9 13 1 9 9 7 10 13 9 9 15 10 1 9
12 7 13 16 13 11 0 9 13 9 1 9 15
20 13 16 9 3 13 7 13 15 15 13 9 7 13 9 15 13 11 1 9 15
8 7 1 9 15 13 0 7 13
13 7 13 11 1 9 11 7 13 9 15 13 1 9
8 0 7 3 9 15 13 1 15
6 7 10 9 13 15 13
9 7 13 11 9 15 13 1 10 0
5 3 13 1 10 0
6 7 11 13 13 1 15
12 7 13 9 3 13 1 15 10 9 7 3 13
12 7 6 9 13 12 9 13 3 13 9 9 15
15 3 16 13 13 10 9 13 3 13 9 15 7 13 10 9
9 7 13 15 9 7 13 15 11 13
13 3 9 3 13 13 15 3 13 7 0 15 3 13
8 3 13 16 13 13 9 1 9
10 7 13 16 13 11 13 10 12 9 15
4 9 1 9 13
3 6 13 15
4 13 7 3 13
10 11 7 11 0 13 1 9 9 3 15
10 3 3 13 12 0 0 9 15 15 13
4 7 15 13 13
7 3 0 13 1 11 10 9
7 1 9 9 12 9 13 15
7 7 10 9 13 10 9 13
2 15 13
11 13 3 15 1 9 13 1 15 9 15 13
10 7 3 1 9 0 13 11 9 0 13
26 7 3 9 9 13 1 12 3 1 3 7 9 13 7 9 13 7 9 13 7 0 9 10 13 0 13
8 7 15 13 13 10 9 13 0
19 13 7 3 11 13 9 9 7 9 0 1 9 15 7 13 9 7 9 0
24 7 1 16 13 13 11 13 11 1 11 13 9 9 9 13 16 13 10 9 7 13 15 9 9
13 7 13 1 11 7 3 9 9 13 1 9 13 15
8 13 7 13 3 1 0 9 0
16 9 3 13 3 13 9 13 1 15 15 10 0 13 7 9 13
16 7 13 1 15 9 13 13 15 7 9 13 7 13 1 15 16
5 7 13 1 15 3
3 7 13 15
6 3 13 13 0 7 0
8 3 9 13 9 0 1 9 0
10 9 1 9 13 13 3 9 1 9 9
14 7 13 15 1 9 0 1 9 9 15 13 1 10 9
13 7 13 1 9 7 13 15 13 15 7 13 1 15
5 3 13 11 11 13
16 7 13 3 9 15 7 9 15 7 3 13 13 1 15 13 15
5 15 13 9 13 13
10 7 0 13 10 1 9 13 10 9 13
11 1 15 9 13 13 15 7 13 15 10 13
15 3 9 9 15 16 13 1 9 0 15 9 13 10 1 9
6 9 3 9 15 16 13
7 7 13 1 9 1 9 11
6 13 9 0 1 10 9
17 7 13 9 10 0 13 1 10 9 7 13 10 9 1 9 1 9
5 13 15 1 9 13
12 3 15 13 13 1 10 9 13 16 9 15 13
3 7 13 15
5 7 13 15 13 13
16 7 13 10 12 7 13 15 13 12 15 7 13 15 9 9 0
25 7 13 9 11 0 3 13 9 15 7 13 16 11 10 9 1 0 13 7 3 13 0 9 1 15
38 7 13 9 0 3 11 9 9 15 9 13 10 0 15 7 9 7 10 0 11 7 13 3 9 11 7 13 7 13 11 7 10 13 13 9 1 0 9
16 7 0 13 10 9 1 10 9 7 1 10 13 3 13 15 13
1 7
15 7 16 13 1 9 1 10 9 13 15 9 15 1 10 9
19 13 7 3 0 9 9 9 0 9 7 13 15 16 10 9 13 1 9 15
16 7 3 13 1 9 11 7 11 13 1 9 11 1 0 9 11
11 7 16 13 15 0 1 9 15 13 1 9
5 7 13 1 10 9
3 6 13 15
10 3 3 13 7 13 16 0 13 9 15
9 7 1 9 13 9 15 13 1 15
30 7 13 13 15 16 13 9 9 3 13 7 13 13 13 1 10 0 7 10 0 9 7 9 7 13 7 1 12 9 13
7 7 15 13 9 9 9 15
18 9 0 13 15 3 13 7 13 9 12 15 12 7 11 12 7 12 11
5 7 13 15 13 16
4 15 13 1 0
5 7 13 15 1 15
3 7 13 13
6 7 1 9 13 13 15
1 9
8 7 16 9 15 13 15 13 15
13 7 13 9 13 15 13 3 13 9 9 13 13 15
11 7 1 9 3 9 15 1 10 0 13 15
9 7 13 15 13 9 1 0 13 15
3 3 13 9
8 7 15 13 1 0 9 13 0
13 7 13 3 10 12 13 15 13 15 13 15 13 16
14 13 3 13 9 15 15 13 7 9 15 15 13 16 13
11 7 15 15 13 13 0 1 15 13 15 9
6 7 13 11 13 13 15
5 7 11 13 1 15
8 7 15 10 3 13 13 1 15
14 7 13 15 1 9 3 13 9 13 1 11 1 10 12
10 7 3 13 16 15 13 9 1 10 9
15 7 1 9 13 15 13 1 15 10 0 9 7 9 7 0
5 7 3 3 13 15
22 9 13 9 7 13 15 9 7 13 9 1 9 7 13 9 7 13 15 9 7 13 3
4 0 13 10 9
8 13 3 16 1 15 10 9 13
7 7 15 13 7 13 1 15
10 7 10 0 13 9 7 13 3 13 9
17 7 1 0 16 13 3 13 1 9 11 1 9 3 15 13 9 13
7 7 13 11 13 13 1 9
9 7 6 10 9 7 13 1 0 9
11 7 9 9 13 13 7 9 10 1 9 13
2 13 0
9 7 15 13 13 7 13 15 9 13
4 7 13 10 9
2 9 9
5 7 13 15 10 9
14 7 13 10 9 9 1 0 13 9 7 13 1 9 9
21 7 13 11 1 9 3 13 12 9 10 0 9 7 13 11 13 15 13 1 15 13
7 7 15 13 13 7 13 16
2 15 13
7 13 3 13 15 10 9 9
2 13 15
4 7 15 3 13
14 3 7 10 0 9 13 15 1 15 3 1 10 9 13
7 7 11 13 16 15 3 13
4 13 3 0 3
6 3 15 13 3 13 15
20 1 0 3 13 10 12 13 7 13 9 15 7 9 16 10 13 15 13 3 13
17 7 0 13 13 1 15 1 9 9 7 10 9 13 1 10 13 9
33 13 3 16 13 15 1 9 9 15 1 9 9 1 9 9 9 15 13 1 13 13 1 9 9 7 15 9 13 9 13 3 9 9
11 15 3 13 0 7 9 15 0 1 9 15
33 3 3 1 9 0 13 13 9 11 1 9 1 9 11 15 13 11 1 9 1 9 9 15 9 11 1 9 11 7 9 10 9 11
6 7 13 1 15 10 9
9 6 3 1 0 3 13 15 15 9
16 7 13 9 7 9 15 16 13 9 9 15 1 15 7 13 15
12 13 3 9 15 3 7 9 15 7 13 13 9
13 13 3 1 9 0 13 9 1 9 11 13 15 9
4 7 0 15 9
20 7 13 15 10 9 13 7 13 9 1 15 15 13 7 13 3 13 13 1 15
10 7 13 15 11 7 13 1 11 9 15
4 15 16 13 15
4 0 13 9 15
5 7 13 15 9 13
4 7 13 1 15
10 15 13 9 15 10 0 1 15 3 13
6 7 13 1 15 10 9
5 3 13 9 9 15
6 13 3 13 1 15 16
6 15 15 3 15 11 9
9 13 3 1 10 9 13 1 9 11
6 3 15 13 1 15 16
6 7 1 9 15 13 9
11 7 13 10 9 1 9 13 15 13 1 15
8 7 15 13 13 1 9 7 13
7 15 13 13 9 7 12 9
4 13 0 0 9
10 7 9 0 1 9 0 13 7 12 13
14 7 13 1 15 16 9 13 10 9 9 3 10 9 9
7 7 13 15 15 13 1 15
9 7 15 13 9 15 1 9 15 13
7 6 16 3 15 13 15 9
12 7 3 13 16 13 15 9 3 15 13 15 3
5 3 13 7 3 13
15 7 15 13 9 1 9 9 15 7 9 1 15 9 3 13
5 0 13 15 13 0
8 7 1 9 15 13 0 7 13
4 7 13 13 9
11 7 13 12 9 15 11 13 15 1 11 13
5 15 13 1 9 13
14 6 15 13 9 15 1 9 15 15 13 9 15 1 15
13 13 3 11 10 9 7 9 13 7 9 13 7 13
6 7 13 11 13 1 11
4 1 15 13 15
58 7 13 3 16 7 15 13 1 9 7 9 13 7 13 9 9 7 10 12 1 15 7 9 15 13 13 9 0 7 9 7 11 15 13 13 11 1 15 13 9 12 7 11 9 11 9 11 7 11 7 0 0 15 13 15 1 9 15
4 15 13 0 9
24 7 10 1 10 0 9 0 13 0 15 1 9 0 7 0 13 10 9 13 7 9 13 1 9
6 13 3 1 12 10 9
4 13 3 1 15
9 3 13 9 10 0 13 1 10 9
14 13 3 10 13 10 13 13 7 13 1 9 7 1 9
3 3 15 13
4 3 13 10 9
2 9 13
10 7 1 15 9 13 3 13 7 3 13
5 3 9 3 13 13
7 7 13 3 7 13 13 15
4 13 3 11 13
13 13 15 10 3 13 15 3 13 9 16 13 9 9
4 13 3 11 13
11 13 3 9 1 15 10 15 3 15 0 13
17 13 3 1 16 13 9 9 15 7 15 9 15 13 1 13 1 11
6 13 15 3 3 13 9
7 7 15 13 7 13 9 9
1 13
6 3 13 1 9 1 9
11 3 11 7 11 0 13 1 9 9 3 15
7 9 15 13 9 0 9 13
5 3 15 13 15 9
9 7 16 13 9 13 0 0 0 0
3 10 0 13
8 7 13 10 9 13 9 15 0
15 7 15 3 13 9 15 7 13 1 15 3 13 13 15 9
5 15 13 9 13 13
8 13 1 15 16 13 9 15 13
8 9 13 1 9 7 1 9 15
6 3 15 13 1 15 16
17 9 15 13 0 15 13 9 7 0 13 13 1 15 16 13 9 15
9 7 13 15 9 9 15 13 10 0
4 7 13 1 15
7 3 15 9 13 12 9 13
15 15 10 13 9 15 7 13 0 13 7 15 15 13 13 13
7 7 3 16 13 15 13 15
4 11 9 13 15
4 7 13 1 15
2 3 13
1 13
4 12 13 13 3
5 7 3 13 0 9
5 12 9 7 0 9
5 13 3 9 13 15
16 15 15 13 13 7 13 0 7 13 9 1 9 7 13 13 15
3 13 3 11
7 13 3 15 16 11 9 13
3 9 16 13
15 7 16 13 1 0 9 13 3 11 13 15 7 13 1 15
23 1 13 3 15 0 13 13 9 1 16 1 11 13 7 13 15 16 3 13 13 9 9 13
4 7 13 1 15
4 7 13 1 15
3 7 15 13
8 13 15 16 16 0 13 9 13
13 7 10 0 9 7 9 13 15 13 7 10 0 9
5 7 3 3 13 15
5 7 13 13 0 9
7 13 15 16 15 13 10 9
6 7 1 15 13 13 15
5 15 13 9 7 9
10 13 9 9 11 7 9 11 7 9 11
12 13 1 0 15 16 15 13 9 15 9 9 15
12 7 13 15 9 3 16 13 9 15 13 1 0
12 13 9 12 3 15 13 12 9 0 7 12 9
10 3 10 9 13 15 13 9 11 13 16
17 3 13 15 13 1 9 7 3 10 9 13 1 9 1 15 15 13
5 0 3 9 13 9
4 3 13 15 11
21 3 9 13 13 1 15 16 9 15 13 15 13 15 7 15 13 15 1 10 0 9
13 0 13 9 15 1 9 13 16 15 0 13 3 13
16 10 3 9 15 1 9 13 9 7 10 9 15 1 9 13 9
3 0 15 13
6 3 13 11 1 10 12
9 0 3 13 15 13 12 13 10 12
5 9 15 3 3 13
8 7 9 0 1 15 13 1 9
6 12 9 13 7 15 13
9 7 11 16 13 3 9 13 3 13
13 3 0 9 1 15 13 7 3 13 1 10 13 15
12 0 3 13 1 9 15 13 13 10 13 1 15
7 15 3 3 15 13 13 15
9 7 0 9 15 3 13 9 13 13
5 15 1 15 15 13
2 13 11
7 0 13 1 15 13 7 13
20 16 15 13 1 9 15 1 9 9 15 13 7 13 9 7 10 9 0 15 13
5 13 16 9 11 13
3 3 13 15
5 3 13 9 1 15
12 15 9 3 13 7 13 9 15 7 15 13 15
3 3 9 13
12 11 9 15 13 3 13 9 15 7 13 7 13
6 3 0 13 15 13 13
6 7 15 13 7 13 13
5 13 3 15 10 9
4 7 13 15 13
14 3 3 13 15 9 16 16 15 15 13 11 1 9 13
5 3 13 1 15 3
7 13 10 9 7 13 1 15
4 13 0 7 13
18 7 16 10 0 9 13 1 15 13 7 10 9 15 13 16 13 9 15
10 9 3 13 3 16 13 7 13 7 13
13 3 15 13 0 1 15 7 15 13 0 1 15 15
8 13 3 9 1 11 7 9 13
10 7 15 9 0 13 15 7 3 13 3
3 13 15 11
6 7 13 0 1 15 3
4 13 1 11 3
10 13 3 3 11 3 9 3 1 9 12
9 13 16 13 1 9 1 10 0 9
10 7 0 16 13 13 3 7 13 1 15
3 7 13 11
4 9 3 0 13
3 11 13 3
18 7 11 13 9 9 9 0 0 7 13 9 11 7 13 9 15 9 15
20 13 3 3 3 10 0 9 16 3 11 13 16 0 1 0 13 9 7 13 11
10 16 9 9 13 1 9 13 15 12 13
5 13 3 9 1 9
9 0 7 3 13 13 0 9 13 13
10 0 13 11 7 13 7 13 15 1 15
13 15 13 1 15 3 13 1 15 7 1 10 13 15
14 16 3 13 9 15 7 13 9 15 13 3 13 1 15
8 16 0 13 0 13 16 13 0
9 6 6 13 15 16 12 15 13 15
19 13 15 7 3 13 1 9 16 3 15 13 15 3 13 13 3 15 13 3
7 9 3 3 13 15 13 3
7 7 3 16 13 13 15 9
6 7 11 13 7 1 15
10 13 15 16 15 1 9 7 9 1 15
4 3 13 15 9
21 16 15 15 13 9 15 13 7 9 15 13 15 7 1 15 13 7 9 1 15 13
5 13 7 13 1 15
8 3 13 15 9 3 15 13 15
33 3 15 15 13 7 15 13 15 7 13 15 16 15 13 7 9 13 7 9 15 1 9 13 16 15 3 13 9 1 9 15 13 15
9 16 13 7 13 1 15 9 3 13
4 1 9 13 15
10 3 16 15 3 13 9 3 13 1 15
6 15 15 13 9 15 13
12 6 6 13 15 16 13 7 13 15 7 9 13
16 7 13 9 15 15 3 3 1 9 13 7 3 1 9 13 15
17 0 3 13 10 0 9 16 13 15 12 0 9 7 15 13 11 11
13 7 15 15 15 13 7 15 15 7 13 13 1 0
12 1 10 9 3 13 3 15 1 10 9 3 13
4 7 15 15 13
4 3 13 15 11
7 16 3 15 13 13 0 13
15 13 7 3 11 15 13 9 16 0 13 12 9 13 1 9
10 7 3 13 1 15 11 13 7 13 15
7 0 9 13 15 13 11 9
4 3 13 15 11
4 3 15 9 13
6 15 13 16 9 13 15
4 6 0 7 11
5 6 0 13 10 9
9 7 13 1 9 3 7 13 1 11
4 7 9 13 13
6 3 1 9 9 13 0
4 15 13 3 13
22 7 13 0 9 1 9 15 13 9 9 15 7 13 15 1 9 9 10 13 1 9 15
10 7 9 9 9 7 9 9 9 7 9
5 1 15 13 15 9
5 9 3 9 0 13
4 1 11 3 13
6 3 13 9 1 10 13
3 3 13 13
5 0 13 11 3 13
7 15 10 13 1 15 3 13
5 7 3 15 13 9
3 3 11 13
2 3 13
28 7 16 15 10 9 13 7 15 0 9 13 13 13 1 15 7 0 10 9 7 9 9 13 3 13 1 10 9
4 3 3 15 13
30 13 3 1 9 9 15 13 13 15 15 13 1 15 3 3 13 16 13 13 7 13 1 3 13 15 3 9 13 9 9
2 9 13
3 13 1 13
2 15 13
10 10 3 9 3 13 9 0 9 7 0
4 13 3 15 13
13 7 0 13 10 9 16 9 13 15 3 1 9 13
7 15 15 13 15 13 0 9
13 15 3 1 0 13 11 3 13 9 7 13 13 9
3 7 3 13
8 13 15 11 9 15 7 15 9
7 15 13 3 3 10 11 9
22 16 3 1 9 9 3 13 10 9 1 9 9 13 9 1 10 9 10 9 13 10 13
7 7 3 9 13 15 1 9
9 15 0 1 11 7 15 0 1 11
19 3 13 3 1 9 0 7 3 1 9 9 7 9 7 1 9 9 7 9
7 7 10 0 15 13 3 9
6 7 3 1 15 9 13
10 15 3 1 9 13 13 9 9 9 13
3 13 13 9
3 3 13 0
8 15 13 9 7 9 0 3 13
8 13 10 0 3 0 16 0 13
2 0 13
20 7 16 15 13 15 10 13 7 13 13 15 15 13 15 13 3 9 13 1 9
11 13 3 3 15 13 16 15 9 9 11 13
8 7 9 9 13 7 13 10 13
9 0 9 10 0 9 13 1 15 9
26 3 9 3 12 13 7 9 13 0 10 7 3 9 15 1 9 10 12 0 13 12 13 9 3 3 11
18 3 3 13 9 13 1 9 15 3 13 7 3 9 1 9 15 3 13
2 3 13
4 9 3 3 13
14 3 13 1 9 13 9 13 16 1 9 9 1 15 13
10 1 15 9 13 15 13 13 16 3 13
8 7 16 9 0 13 3 11 13
11 3 3 1 11 15 13 3 1 11 15 13
12 3 15 13 10 13 1 0 16 3 0 3 13
4 1 9 15 13
4 6 9 15 13
12 7 9 9 15 13 15 9 1 9 15 11 11
5 15 15 1 9 13
9 16 15 3 13 9 11 11 13 9
12 9 15 7 9 1 9 9 15 7 9 11 11
32 7 0 9 13 3 13 1 15 16 0 9 13 7 1 15 13 1 11 7 3 1 11 13 1 15 7 1 15 13 15 1 11
3 16 9 13
17 7 3 15 16 15 13 13 1 15 1 9 11 16 3 13 1 11
5 13 3 15 15 13
25 13 3 0 9 0 9 13 7 3 3 11 13 9 1 9 16 16 3 13 9 11 1 9 10 13
15 0 3 15 1 15 16 9 13 1 0 9 13 1 9 9
14 7 13 7 13 3 13 1 10 9 7 0 13 1 9
10 3 15 1 10 3 3 15 13 1 9
12 9 3 13 0 13 15 7 1 9 9 13 15
10 7 10 0 9 3 9 13 13 3 15
3 13 9 9
3 13 13 9
24 13 3 0 10 1 9 13 15 0 13 15 9 7 9 7 9 7 9 7 9 7 9 7 9
23 1 0 3 9 15 9 1 0 9 16 3 0 9 13 1 15 9 16 13 9 3 13 13
15 7 9 9 15 7 15 9 1 15 1 15 13 1 9 9
1 13
49 1 9 3 13 3 1 9 13 16 9 15 9 3 0 7 0 9 1 9 9 9 13 7 15 9 13 1 9 9 7 13 15 9 7 1 9 11 13 7 3 13 1 13 15 9 16 13 15 9
18 3 3 3 3 13 1 15 9 13 15 16 3 1 15 13 1 9 11
12 13 3 3 9 15 0 13 10 1 0 13 9
20 7 15 13 3 13 13 16 13 9 10 13 9 16 1 15 13 13 3 3 15
8 1 9 13 3 16 15 0 13
6 15 13 7 15 3 13
10 1 15 12 9 9 13 16 13 1 15
16 15 3 13 0 0 13 1 0 9 3 16 15 0 3 13 15
5 3 15 13 15 11
20 3 0 0 9 3 3 3 13 10 1 13 7 0 15 16 16 13 3 3 13
16 3 16 15 13 13 7 16 15 10 0 13 7 15 3 13 13
8 7 9 9 7 9 13 1 15
1 6
9 3 16 13 15 1 11 1 9 13
11 3 16 15 13 0 3 13 13 15 0 13
3 3 0 13
8 3 15 15 12 13 1 11 11
8 7 16 9 3 9 9 1 11
12 13 3 15 16 16 0 13 9 15 13 13 15
7 7 3 10 1 9 1 9
10 16 0 9 10 0 3 3 10 13 9
11 7 10 13 15 0 13 10 9 15 15 13
4 7 9 1 9
9 15 3 9 13 7 3 13 9 11
7 7 10 0 13 3 13 0
8 3 15 9 11 1 9 15 13
115 3 3 15 13 15 9 1 9 11 11 7 9 1 15 10 0 13 13 1 15 9 13 1 9 15 16 9 9 15 11 11 9 9 13 15 9 9 7 9 1 9 15 13 9 9 15 16 13 15 15 13 9 9 15 0 7 9 9 9 15 1 0 7 15 9 9 9 15 1 15 10 13 1 9 9 9 15 15 13 1 11 13 15 1 0 7 13 1 0 15 1 9 1 15 9 7 9 7 9 7 9 7 15 9 13 3 3 1 0 9 7 3 1 10 0
12 7 13 13 9 15 15 3 7 9 0 15 3
78 1 0 13 9 15 1 9 9 15 11 11 1 15 15 9 1 9 7 1 9 13 16 13 15 1 9 9 15 9 13 1 9 15 1 0 9 13 11 1 9 1 9 15 16 1 9 13 7 13 13 13 1 15 10 0 15 13 9 7 9 7 9 7 9 13 10 9 0 10 9 9 11 16 13 1 15 9 9
14 7 3 13 10 0 9 9 1 15 13 13 1 9 9
5 7 3 13 9 9
10 13 9 0 13 1 9 7 9 7 0
13 9 9 7 9 1 9 1 9 9 7 9 11 11
9 3 15 9 7 9 7 9 11 13
47 3 3 9 11 13 16 7 13 7 13 15 7 3 13 1 15 16 13 1 12 9 12 9 3 13 9 9 7 3 1 9 13 1 10 9 15 13 15 9 9 7 15 9 7 0 1 9
10 3 3 0 13 1 9 7 9 15 13
9 16 15 0 13 13 1 9 15 3
6 3 3 13 1 9 3
14 3 16 1 9 13 16 15 13 15 1 15 13 13 13
24 3 13 1 11 10 0 9 15 15 13 0 1 15 9 11 11 15 7 13 15 15 9 1 9
22 9 9 1 9 11 13 15 1 9 1 15 3 13 1 9 9 9 15 13 15 1 0
10 15 3 13 13 3 0 15 1 9 13
28 13 15 3 3 13 9 0 7 0 9 9 9 9 9 9 9 13 15 3 7 13 0 16 15 1 15 13 9
5 9 13 9 1 15
4 0 3 13 13
61 15 3 13 13 9 9 9 10 13 1 11 1 11 11 16 10 0 13 3 15 1 15 9 3 3 15 1 9 15 7 9 13 11 7 0 9 7 15 13 7 9 3 13 7 15 9 0 13 13 15 1 9 13 16 13 7 1 13 15 9 3
22 3 7 15 3 3 13 13 1 13 9 15 16 3 13 15 10 13 7 3 13 9 15
17 1 7 0 3 15 13 3 9 13 7 9 15 13 9 15 0 15
12 7 1 10 9 7 9 9 3 13 16 15 13
14 1 7 0 13 15 3 7 13 15 15 15 3 3 13
3 1 15 13
6 13 9 15 1 9 0
94 9 0 9 9 1 0 13 15 9 9 1 15 3 13 3 16 0 13 1 9 13 10 13 15 9 7 15 13 9 1 15 1 9 9 15 11 1 9 1 9 9 15 1 9 9 13 9 3 13 9 7 3 13 9 9 15 11 11 15 9 13 9 0 1 9 9 7 1 9 9 15 16 13 13 1 10 0 15 7 13 1 15 10 13 3 13 13 9 15 1 15 1 9 0
10 7 3 3 9 15 13 7 13 3 9
11 9 9 9 1 9 9 7 11 11 9 15
1 6
13 7 13 9 3 13 7 13 1 9 7 13 1 9
17 13 3 15 9 0 13 1 10 3 16 3 13 1 9 7 9 9
13 3 15 9 9 0 7 3 9 1 9 1 9 13
17 3 13 0 10 1 15 9 15 13 13 15 1 9 1 9 9 9
9 7 10 13 1 9 3 13 0 13
16 3 3 3 9 0 0 13 7 15 3 15 13 13 3 13 13
24 7 15 13 0 13 13 1 9 7 9 9 7 9 0 0 7 0 15 13 9 1 9 7 9
58 13 9 15 15 13 1 9 1 0 9 3 13 13 1 15 9 1 9 15 9 7 9 13 15 13 13 9 15 16 9 13 9 13 10 15 13 1 15 0 9 15 13 3 1 9 15 11 7 9 15 11 13 7 3 16 3 1 15
10 7 3 3 1 11 13 15 3 15 13
20 1 0 15 13 1 10 13 16 3 0 9 13 15 13 1 11 11 1 9 0
6 7 10 0 0 9 13
46 7 0 13 16 1 0 9 13 9 0 7 13 9 15 13 0 9 0 13 9 0 0 0 0 0 13 13 15 0 0 13 0 13 13 9 15 3 3 9 13 9 9 7 9 15 13
26 15 9 0 9 7 0 1 9 1 9 1 9 1 9 1 9 16 13 13 9 9 1 15 9 0 13
3 11 1 11
4 7 15 15 13
4 0 13 9 0
10 16 3 15 13 1 9 13 0 3 15
9 13 15 11 10 13 15 1 11 11
