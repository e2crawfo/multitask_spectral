720 11
30 13 11 16 13 9 0 15 1 9 10 9 7 10 9 10 1 9 10 9 9 9 2 9 0 1 9 0 10 9 2
14 13 9 0 1 9 1 10 9 10 1 9 0 9 2
18 13 9 9 1 1 7 13 15 3 1 9 15 7 13 15 9 1 2
55 16 13 2 1 15 2 14 13 10 9 11 10 9 11 14 11 1 9 1 1 10 9 2 13 0 9 3 16 10 9 14 13 1 9 1 11 10 9 9 0 3 10 9 10 10 9 9 1 9 10 9 1 10 9 2
24 9 2 11 14 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2
25 13 15 1 1 10 9 14 13 1 9 10 9 9 14 9 1 10 9 10 9 9 14 9 3 2
5 11 13 15 15 2
22 1 9 2 14 13 9 1 9 9 1 9 1 9 9 1 9 14 9 7 14 9 2
17 13 0 14 13 9 10 1 11 2 1 9 7 8 2 1 9 2
23 14 13 9 14 9 14 13 9 1 9 9 0 1 9 9 15 14 9 0 1 12 9 2
3 11 11 2
13 1 9 1 14 12 1 9 14 13 3 10 9 2
5 13 9 1 3 2
23 2 15 1 14 13 15 9 1 9 1 2 7 13 15 10 9 9 14 0 1 10 9 2
15 9 0 1 9 10 11 14 13 1 9 9 14 13 1 2
31 16 16 14 13 15 1 15 16 13 1 9 9 14 13 15 1 9 1 15 2 13 15 1 9 0 14 13 10 9 1 2
9 10 9 1 9 1 11 11 11 2
34 10 9 14 13 1 11 7 1 15 7 9 0 9 14 9 1 9 2 7 6 2 1 9 9 2 14 13 1 10 9 1 10 9 2
6 14 13 15 10 9 2
7 13 9 10 1 10 9 2
34 13 0 13 0 11 1 9 10 9 7 11 1 9 7 1 9 1 9 9 13 9 0 1 10 9 14 13 10 9 1 9 0 10 2
30 9 10 1 9 10 13 15 0 1 9 1 2 13 0 2 13 9 9 0 1 10 9 0 14 13 15 1 10 9 2
16 1 9 7 12 3 0 14 13 15 1 9 10 9 1 9 2
8 11 2 15 13 1 9 1 2
28 13 9 1 10 9 10 16 13 9 1 9 16 14 13 10 9 10 1 1 9 14 9 3 1 10 9 0 2
20 13 0 3 1 9 10 9 1 13 10 9 13 3 13 9 7 9 10 9 2
8 13 0 1 11 1 9 10 2
9 13 11 10 9 14 13 1 9 2
4 9 13 15 2
4 14 13 11 2
23 16 16 14 13 1 1 9 2 14 13 9 11 11 11 2 13 1 9 1 9 14 9 2
82 9 12 16 13 9 7 9 10 9 9 14 9 1 10 9 9 14 9 1 9 1 9 10 9 9 2 13 10 9 10 15 14 9 0 1 9 10 9 9 2 1 10 9 2 16 13 9 7 9 10 9 9 14 9 1 10 9 9 14 9 1 9 1 9 10 9 9 2 13 10 9 10 15 14 9 0 1 9 10 9 9 2
7 13 1 9 9 13 15 2
29 1 9 10 2 1 10 9 1 9 2 7 14 13 15 0 1 10 9 1 9 1 10 9 9 13 0 3 1 2
7 9 1 10 9 1 9 2
22 9 10 11 13 1 10 9 16 13 11 9 10 12 9 14 13 1 2 1 10 9 2
1 2
36 13 9 1 9 1 9 1 9 10 14 13 1 11 11 15 11 1 10 9 10 16 13 9 9 14 9 1 1 15 15 2 9 14 13 9 2
20 14 13 15 1 10 11 9 11 11 7 13 15 1 9 1 9 1 10 11 2
13 13 0 1 11 14 13 9 9 0 1 9 0 2
19 14 13 15 9 1 9 1 2 1 15 2 13 15 1 9 10 9 1 2
14 13 3 1 9 1 9 0 10 9 8 14 13 15 2
30 13 9 1 10 9 14 9 1 9 14 0 1 11 14 11 2 9 0 10 9 9 2 14 13 9 1 9 1 9 2
15 13 15 1 16 9 1 10 9 2 13 15 10 9 1 2
29 9 16 13 15 1 9 2 13 1 9 10 9 14 13 1 10 9 14 9 1 9 0 7 1 9 0 1 9 2
24 9 7 9 1 9 10 9 1 11 11 15 11 14 11 14 13 1 11 10 9 2 9 11 2
44 13 15 1 9 9 2 9 2 9 2 14 13 9 1 1 11 14 9 1 9 2 14 9 1 9 1 9 14 9 1 10 9 1 9 10 11 1 10 12 7 10 12 9 2
10 2 9 1 9 11 0 13 15 15 2
81 8 1 9 13 1 9 1 9 8 2 8 16 9 15 13 1 9 8 8 14 13 15 2 13 9 15 13 9 0 10 9 14 13 10 9 2 7 8 16 9 15 13 1 9 8 8 14 13 15 2 13 9 15 14 13 10 9 1 9 9 12 7 14 13 10 9 1 9 1 9 9 12 7 13 9 15 1 14 13 1 2
9 13 9 1 10 9 14 10 9 2
37 13 0 1 15 2 3 2 10 9 9 0 15 14 9 1 9 1 9 14 9 1 10 9 0 14 0 14 13 9 0 10 2 9 10 12 9 2
23 2 13 9 13 0 1 9 9 10 1 9 3 1 14 9 1 9 10 9 9 3 1 2
41 14 13 15 2 1 15 15 2 9 1 10 9 14 13 1 9 1 9 2 2 16 13 9 1 9 9 15 9 1 9 14 13 10 9 2 13 15 1 9 2 2
4 2 14 13 2
20 14 13 15 3 14 0 1 10 9 1 10 9 10 9 16 14 13 9 1 2
36 13 9 1 9 1 10 11 11 1 9 9 10 11 7 15 1 9 10 9 14 9 3 1 9 10 9 1 9 11 2 9 14 13 1 9 2
21 13 10 12 9 2 11 7 11 0 0 7 14 13 9 1 10 9 13 9 15 2
16 13 15 11 8 11 13 9 1 10 9 14 9 1 9 12 2
5 13 1 10 9 2
13 11 0 14 13 1 1 10 9 14 0 14 9 2
21 13 15 3 0 1 10 9 7 13 9 15 9 14 13 10 9 1 1 10 9 2
6 13 10 9 1 9 2
28 16 14 13 11 10 9 1 16 15 1 9 10 9 14 9 13 15 10 9 1 9 7 14 13 10 9 1 2
49 13 11 1 9 13 0 10 9 14 13 10 9 0 10 2 11 9 2 1 9 10 9 2 13 15 15 2 1 10 9 14 13 1 2 16 14 13 9 10 10 9 14 0 0 1 11 9 2 2
8 1 9 10 9 14 13 15 2
8 13 11 11 1 9 1 11 2
71 16 14 13 15 1 12 9 10 9 16 14 13 1 9 3 0 16 14 13 2 14 13 2 16 14 13 11 13 1 15 14 13 16 16 13 15 14 13 15 3 2 16 13 1 9 1 14 13 15 15 7 16 13 15 15 10 9 10 9 14 9 2 9 16 14 13 9 0 2 0 2
15 13 10 9 1 10 15 10 9 1 15 15 14 9 3 2
15 12 9 13 1 8 7 12 9 2 9 2 9 2 9 2
25 13 9 14 13 9 1 15 2 3 9 2 1 14 13 0 1 1 9 9 1 9 0 10 9 2
4 9 1 9 2
25 13 15 9 10 9 14 9 1 9 9 10 9 1 9 0 2 7 9 10 9 1 10 9 10 2
11 11 13 10 9 1 10 9 2 14 9 2
34 13 9 10 1 9 10 9 2 11 11 11 2 14 13 3 1 12 12 1 9 9 1 9 0 16 14 13 10 9 9 1 9 12 2
28 16 14 13 1 9 10 9 0 14 9 13 1 9 7 1 9 0 0 15 1 10 9 0 2 13 9 0 2
35 13 8 1 9 1 10 9 1 1 9 9 9 0 7 9 10 9 11 16 13 0 3 1 9 8 12 1 9 1 10 9 11 14 9 2
7 13 15 1 9 1 9 2
5 6 2 14 9 2
17 1 9 10 13 15 9 9 1 1 9 10 9 0 10 1 11 2
7 15 15 10 9 3 15 2
13 14 13 15 15 9 9 1 10 9 2 1 11 2
10 13 9 0 1 1 9 9 0 9 2
36 16 15 1 9 10 9 10 1 9 11 2 13 9 1 3 15 14 13 1 10 12 9 7 1 10 9 14 0 14 9 0 1 9 10 9 2
14 7 1 9 14 9 13 10 9 10 9 3 10 9 2
19 13 10 9 11 2 8 11 2 2 9 0 9 2 1 1 10 9 10 2
35 14 13 15 10 9 1 9 1 2 14 13 9 0 0 1 11 2 10 9 0 2 3 12 9 9 1 15 7 14 13 15 1 9 9 2
15 16 13 15 1 9 3 1 9 9 7 13 12 9 1 2
2 11 2
11 15 13 1 9 10 9 9 10 9 10 2
26 13 15 14 13 11 11 1 10 9 9 2 16 14 13 10 12 9 1 11 7 10 11 1 9 12 2
7 9 1 2 14 11 0 2
7 9 9 9 14 13 1 2
5 13 9 9 1 2
4 13 15 0 2
29 1 9 10 2 13 9 1 11 14 11 2 10 9 14 13 9 10 9 1 9 9 14 13 15 1 11 1 9 2
35 13 0 14 13 15 10 9 10 3 2 16 13 15 0 14 0 1 9 11 14 13 10 11 14 13 1 9 1 9 9 14 9 1 9 2
33 9 11 9 11 13 9 9 15 11 11 2 1 9 2 9 14 13 1 9 0 1 9 9 2 7 13 9 15 1 10 9 9 2
16 2 13 1 9 3 2 2 14 13 15 3 7 9 1 9 2
19 1 10 9 9 14 13 1 9 13 9 10 9 1 1 9 11 9 0 2
18 13 0 9 1 1 9 14 9 1 10 9 15 14 13 9 13 9 2
18 13 10 9 10 9 1 7 13 14 13 10 9 9 9 0 1 11 2
26 13 10 9 0 2 1 13 9 0 14 13 15 2 13 15 1 9 0 16 9 9 0 14 13 15 2
24 2 13 12 9 15 15 2 2 13 10 9 10 7 14 13 15 1 10 9 14 9 1 9 2
24 2 14 13 15 9 2 13 10 9 2 7 14 13 15 9 2 13 10 9 2 2 13 11 2
22 13 9 10 11 9 9 1 9 14 13 10 11 1 9 1 10 9 10 1 9 9 2
44 13 1 9 14 13 1 10 9 15 2 16 13 10 9 1 1 9 0 0 15 14 13 15 1 1 9 0 2 7 13 9 10 3 15 1 9 0 10 9 14 13 14 9 2
10 13 15 3 16 14 13 10 9 3 2
8 2 13 15 2 2 13 15 2
1 2
54 13 10 9 1 11 1 10 11 11 11 7 13 15 9 14 13 9 1 9 10 9 0 2 13 1 9 10 9 1 10 9 2 14 13 9 1 10 9 14 9 1 10 9 9 1 16 13 1 10 9 0 1 11 2
22 13 11 0 0 1 1 11 3 2 11 0 1 10 9 1 11 14 11 1 9 11 2
112 8 13 9 14 13 1 9 13 9 15 1 13 7 1 13 1 10 9 7 1 9 1 9 8 1 9 1 9 9 14 13 1 9 10 9 1 10 9 1 9 9 14 0 14 13 7 14 13 3 2 13 10 9 10 1 9 1 10 9 2 1 14 13 10 9 2 1 10 9 14 13 10 9 0 1 9 8 1 9 9 14 9 9 1 9 1 9 8 7 1 9 7 1 9 8 13 10 9 0 1 9 8 1 9 9 14 9 1 9 0 3 2
28 13 10 9 1 9 1 14 13 10 9 2 12 9 1 15 2 1 9 14 13 1 9 9 0 0 14 9 2
14 13 9 9 7 9 1 3 0 1 9 1 10 9 2
34 7 1 9 14 13 15 10 9 1 9 10 11 1 14 12 10 9 9 2 13 14 0 1 7 13 15 1 9 1 9 10 9 9 2
22 13 10 9 1 9 1 10 9 9 1 11 2 15 0 1 9 9 9 11 1 11 2
17 13 15 14 13 9 1 9 10 11 16 14 13 1 9 10 9 2
16 13 10 9 0 1 1 9 1 9 9 14 13 1 14 0 2
19 2 13 9 14 13 9 9 1 15 10 9 10 1 2 2 14 13 15 2
5 13 7 14 13 2
37 9 10 9 9 14 13 1 9 9 14 13 15 9 1 9 1 9 14 13 9 1 1 16 14 13 1 11 0 1 9 10 9 1 11 11 9 2
24 13 9 10 9 0 1 3 2 1 7 1 2 7 13 10 9 15 1 10 9 1 9 15 2
6 14 13 15 3 3 2
21 10 9 14 13 1 9 1 14 9 16 9 14 9 7 9 1 10 9 1 9 2
8 1 9 3 1 10 9 9 2
14 11 15 9 1 16 10 9 1 1 9 1 9 1 2
35 1 10 12 9 3 2 13 10 9 10 1 9 10 9 1 9 10 9 10 0 7 9 10 9 0 2 13 9 1 15 1 9 10 9 2
28 14 13 10 11 1 10 9 10 7 13 1 9 3 1 12 9 1 14 13 1 10 9 2 11 11 2 9 2
19 14 13 9 1 10 12 9 14 9 2 15 15 15 7 15 14 13 1 2
9 10 9 1 10 9 1 9 11 2
55 14 9 11 11 2 16 13 10 9 14 9 1 10 9 16 14 13 1 9 11 2 13 15 1 9 1 14 13 15 1 9 1 10 9 1 9 10 9 13 15 10 9 15 14 13 10 9 0 1 9 0 14 13 1 2
27 2 9 2 16 14 13 10 9 10 9 0 2 7 10 9 0 2 9 9 1 10 9 13 9 1 15 2
18 13 15 9 16 13 0 3 1 2 9 14 13 3 1 9 10 9 2
14 13 10 9 14 13 10 9 9 1 9 1 9 9 2
7 14 13 1 10 9 3 2
21 9 0 1 12 9 3 2 13 9 11 11 1 9 14 0 1 9 9 14 9 2
26 14 13 16 12 1 9 1 1 12 16 13 9 14 11 1 9 9 1 9 9 14 9 1 10 9 2
57 2 11 0 10 13 15 11 14 11 2 9 10 9 10 2 10 9 1 9 2 2 9 14 13 9 10 9 1 2 7 9 14 13 9 1 9 2 1 9 7 1 9 13 0 1 9 10 11 2 16 14 0 1 9 10 9 2
15 13 10 9 9 9 1 1 9 0 1 15 9 9 15 2
28 2 13 9 16 9 1 10 9 14 13 1 9 1 9 11 14 13 14 13 15 15 1 9 10 9 0 3 2
31 16 14 13 1 11 14 11 15 13 10 9 10 9 14 9 1 9 7 9 1 9 15 10 9 14 13 10 9 1 9 2
4 2 11 3 2
3 10 9 2
19 9 14 13 1 2 8 1 9 16 14 13 15 7 16 14 13 9 1 2
6 7 13 9 0 1 2
19 13 15 9 14 9 3 7 13 15 10 9 9 1 9 1 9 10 9 2
6 13 15 13 9 15 2
46 14 13 14 13 10 9 9 14 13 1 9 1 9 1 9 0 14 13 1 9 10 9 7 13 9 1 9 14 13 9 0 1 9 1 9 10 9 10 7 14 0 10 9 10 1 2
26 13 11 11 7 9 9 10 10 9 14 9 7 13 11 1 9 14 13 9 14 9 1 10 9 9 2
17 13 10 9 1 9 1 10 9 1 1 10 9 14 9 1 9 2
8 14 13 9 1 9 1 9 2
6 9 1 11 14 9 2
9 13 15 15 10 9 2 9 2 2
24 13 15 10 9 10 9 1 10 9 1 9 9 14 9 1 9 2 11 2 7 1 10 9 2
28 13 12 9 11 1 3 2 2 9 0 0 7 9 0 0 2 2 2 12 2 8 14 13 15 1 9 12 2
10 13 10 9 0 14 13 15 3 0 2
58 13 9 0 1 9 0 1 9 1 15 1 9 1 2 9 10 9 2 2 2 9 9 10 9 2 7 2 1 11 1 9 2 2 1 9 7 9 2 7 1 2 9 10 9 2 7 2 1 9 1 9 2 2 10 9 0 2 2
52 1 10 9 2 13 9 1 10 9 15 1 9 1 9 16 10 9 0 2 7 13 13 0 1 9 13 15 9 10 9 10 11 14 11 13 1 9 1 9 10 9 10 3 2 10 12 9 2 16 13 15 2
66 13 10 9 1 1 9 14 9 1 9 10 9 9 1 15 14 13 15 1 9 2 2 13 1 9 1 11 11 10 9 7 13 10 9 1 3 14 13 9 1 10 9 9 7 14 13 9 1 1 9 2 2 14 13 11 11 2 9 1 10 9 1 12 9 3 2
5 13 15 1 9 2
8 13 9 14 13 15 1 11 2
7 14 13 15 10 9 1 2
8 3 1 14 13 15 1 9 2
20 13 15 14 13 7 14 13 10 9 1 11 7 9 1 10 9 14 9 3 2
21 2 9 2 9 9 10 9 0 13 1 9 3 1 9 12 9 14 11 1 9 2
37 13 0 10 9 10 1 9 9 7 9 1 12 12 9 16 13 15 0 1 9 3 1 9 1 9 9 1 9 10 9 7 1 9 1 9 0 2
10 13 15 3 1 10 9 7 9 9 2
6 2 9 9 0 2 2
8 13 0 1 9 3 14 11 2
37 1 9 9 3 2 13 10 11 9 1 9 11 1 9 1 14 0 1 9 10 9 1 9 0 10 8 2 16 0 7 8 16 15 9 10 2 2
22 14 13 12 9 1 9 10 9 0 7 14 13 2 9 9 7 14 13 9 9 15 2
14 13 10 9 9 7 15 1 9 9 14 13 10 9 2
8 13 9 0 1 9 1 9 2
7 15 0 7 0 7 0 2
28 13 10 9 9 1 9 0 10 16 13 9 1 9 9 2 1 9 7 13 13 9 0 1 9 0 1 11 2
3 14 13 2
30 13 0 14 13 9 11 2 15 1 9 7 1 11 11 1 9 10 2 1 9 0 1 11 2 7 9 9 14 0 2
5 14 13 15 0 2
14 11 0 15 11 14 13 1 9 14 0 9 11 11 2
4 9 7 9 2
8 13 15 1 9 7 1 9 2
3 2 9 2
9 13 10 9 3 1 9 14 0 2
24 13 9 10 9 2 11 14 11 2 1 9 10 9 2 8 10 11 2 9 10 9 1 15 2
13 13 9 1 10 9 1 11 11 1 12 9 9 2
67 16 14 13 15 9 1 11 14 9 14 13 10 9 9 9 1 2 11 1 9 1 11 14 13 9 1 1 10 9 15 7 15 7 11 1 9 1 2 13 9 13 15 1 9 9 11 1 11 1 9 7 13 9 9 1 10 9 13 0 1 9 16 13 0 1 15 2
24 9 14 9 1 9 9 14 13 9 1 10 9 0 7 14 13 9 1 9 9 9 1 9 2
28 13 9 1 10 9 2 11 11 2 9 1 9 14 9 1 9 10 10 9 7 13 15 9 9 1 1 0 2
33 13 9 0 14 13 1 9 1 2 9 8 14 13 1 9 9 0 14 9 1 8 13 1 10 9 14 13 1 9 10 9 9 2
17 9 14 13 15 1 10 11 11 7 13 15 0 1 9 10 9 2
15 13 11 14 11 1 9 1 10 9 14 0 7 14 0 2
10 9 9 1 9 1 2 9 0 2 2
17 1 9 10 14 13 10 9 14 9 3 1 9 1 9 0 9 2
22 9 14 13 1 9 0 14 13 10 9 9 1 15 2 9 9 2 9 7 9 0 2
12 13 15 10 9 1 9 1 9 1 9 10 2
15 13 10 9 14 13 1 11 14 11 1 9 7 9 1 2
6 13 15 10 9 1 2
18 13 9 9 3 1 9 7 13 15 1 9 10 9 1 9 1 9 2
4 2 13 1 2
22 13 9 14 13 1 9 3 1 10 9 8 7 9 1 9 10 9 14 13 1 9 2
13 10 9 13 1 7 2 8 8 2 8 8 8 2
5 9 9 9 8 2
15 7 13 2 1 9 9 9 14 13 10 11 9 11 1 2
24 13 10 9 14 13 15 1 9 1 2 11 10 9 1 9 9 14 13 0 9 10 9 10 2
24 13 9 1 14 13 15 1 10 9 13 0 16 13 9 1 3 1 2 1 9 7 1 11 2
36 13 15 10 9 14 0 2 1 9 2 14 13 10 9 9 0 1 9 1 9 10 11 7 14 13 1 1 9 10 9 14 13 9 10 9 2
48 1 9 10 9 2 9 10 9 1 10 9 7 9 10 9 7 13 10 9 1 1 9 2 1 9 9 13 10 9 1 9 1 16 9 1 10 9 3 1 9 10 9 7 1 9 1 9 2
34 13 15 10 9 14 13 1 7 13 9 14 13 12 9 0 1 9 9 1 13 1 9 2 1 9 9 10 9 7 1 9 9 9 2
14 13 9 15 10 9 1 2 9 2 9 7 9 9 2
49 9 13 10 9 1 9 0 13 1 9 10 9 1 9 14 13 1 10 9 2 16 13 10 9 11 11 2 14 13 10 9 14 9 1 9 7 9 2 14 13 15 1 9 1 9 0 1 8 2
11 13 9 0 10 9 1 9 1 10 9 2
2 11 2
7 13 15 13 1 9 1 2
6 3 13 15 1 9 2
15 10 12 9 0 2 10 9 3 2 13 2 10 9 3 2
9 14 13 10 9 14 13 10 9 2
8 13 10 9 14 14 13 15 2
22 2 9 0 3 13 2 2 9 9 11 11 2 1 9 3 1 10 9 9 10 9 2
20 15 15 10 9 14 13 1 10 9 1 9 11 13 0 14 13 10 9 9 2
33 13 15 9 2 3 2 1 9 2 0 2 10 9 2 12 2 2 14 13 2 16 13 15 1 9 0 1 9 2 2 12 2 2
44 13 15 9 0 1 15 2 1 9 10 9 1 9 2 7 1 9 14 0 16 13 13 1 10 9 14 13 15 2 7 2 1 10 9 2 14 13 13 1 9 14 13 15 2
26 1 9 0 2 13 9 10 9 7 9 10 9 7 9 10 9 1 7 10 9 1 10 9 15 1 2
39 13 15 11 14 9 14 13 10 9 7 16 9 13 9 0 1 11 1 9 1 9 7 13 9 1 1 9 10 9 0 14 14 13 15 9 9 1 15 2
25 2 13 9 1 9 1 9 0 13 1 9 1 9 16 13 1 14 9 1 9 1 11 11 9 2
24 13 15 9 1 9 7 1 9 10 9 9 2 16 13 15 0 3 1 9 2 1 15 15 2
31 15 1 14 13 15 1 9 1 15 15 14 9 1 9 10 1 14 13 10 9 14 13 10 9 11 1 9 1 9 10 2
6 14 13 15 10 9 2
7 13 10 9 2 0 2 2
37 13 9 0 2 1 9 10 9 7 13 15 9 2 1 9 10 9 10 9 9 7 9 2 0 1 9 7 14 13 15 1 9 2 1 9 0 2
28 13 1 12 3 14 13 9 1 9 0 1 9 0 14 13 9 1 9 10 8 7 14 13 1 9 10 11 2
6 9 11 11 1 9 2
33 8 13 9 0 1 9 9 1 9 9 14 13 1 9 10 11 16 13 15 7 15 1 9 9 10 9 10 14 9 1 7 1 2
86 9 9 2 9 14 13 1 9 0 0 8 9 0 14 0 0 8 9 0 14 0 0 8 9 0 14 0 0 8 9 0 14 0 0 9 2 8 9 0 14 0 0 8 9 0 14 0 0 8 9 0 14 0 0 0 9 0 14 0 0 8 9 0 14 0 0 8 9 0 14 0 16 9 0 15 13 0 15 7 13 8 1 1 9 9 2
20 2 1 9 2 9 0 9 9 0 9 9 9 1 9 11 9 11 8 11 2
34 8 1 9 14 13 9 1 10 9 1 9 10 2 13 10 11 9 10 2 0 2 1 1 9 10 9 14 13 14 9 1 9 9 2
20 13 10 12 9 1 9 9 1 9 12 7 1 9 12 13 12 9 1 9 2
26 13 15 0 14 13 15 3 0 2 1 9 9 1 9 9 2 1 9 14 13 7 9 9 14 9 2
38 8 1 9 9 8 1 9 10 2 13 15 14 13 1 10 9 9 10 9 9 13 0 1 10 9 7 13 9 13 9 1 9 14 9 1 10 9 2
22 13 15 14 13 1 9 1 10 9 10 7 9 0 10 9 1 9 14 13 1 9 2
37 2 8 2 10 9 14 13 2 1 9 0 2 10 9 1 9 1 9 10 2 13 10 9 12 9 9 9 14 13 0 1 14 9 7 14 9 2
11 13 15 3 14 0 16 14 14 13 1 2
26 13 10 9 9 10 0 1 10 9 0 14 9 1 9 2 14 13 10 9 9 10 9 10 1 9 2
6 13 2 13 7 13 2
213 3 1 9 12 9 1 1 9 11 9 1 9 2 13 10 9 10 9 10 14 13 2 1 9 1 1 9 1 10 9 9 16 13 1 9 12 2 8 9 1 9 14 9 2 1 9 9 12 2 14 13 10 9 1 9 2 13 15 1 9 1 9 7 1 9 1 12 9 2 1 9 9 0 1 2 8 9 1 9 0 10 9 14 9 14 13 2 8 9 7 9 9 14 13 10 9 7 9 1 9 1 1 9 1 9 1 9 10 2 8 9 1 9 1 9 9 0 13 0 16 12 9 2 14 13 2 8 9 10 12 9 14 13 1 10 9 9 14 9 1 9 1 1 9 9 0 1 7 9 10 12 9 14 13 10 9 0 1 9 10 2 8 10 9 9 7 10 9 1 9 1 9 9 2 8 9 0 1 9 2 8 9 1 9 9 2 8 9 1 9 3 10 9 14 13 9 9 1 9 12 9 1 9 10 9 1 9 13 0 16 12 9 2
14 16 13 1 11 1 9 2 13 11 11 3 1 9 2
67 9 9 10 11 2 11 11 2 10 9 0 2 11 11 2 9 0 10 11 2 11 11 2 9 10 9 0 2 11 11 2 9 0 10 11 2 11 11 2 11 10 11 2 9 14 11 2 11 11 2 11 10 11 2 9 11 2 11 11 2 11 9 11 2 11 2 2
37 13 0 9 1 9 9 10 9 7 10 9 1 14 9 14 13 10 9 1 9 10 3 0 1 16 13 9 10 9 1 9 9 10 9 1 9 2
10 13 10 9 10 3 0 2 3 0 2
22 9 10 9 2 9 1 14 13 10 9 0 1 1 9 0 7 10 14 9 1 9 2
42 13 0 1 0 7 0 0 1 9 7 14 9 0 1 10 9 13 1 9 1 16 13 15 1 9 2 1 9 2 7 1 9 1 10 9 1 2 13 1 9 15 2
5 13 1 10 9 2
7 9 9 0 0 1 9 2
27 1 9 16 13 9 0 10 1 9 1 10 9 13 1 9 1 9 13 10 9 1 9 14 9 14 0 2
19 2 13 10 9 1 11 1 9 3 1 10 9 7 14 13 15 1 3 2
10 2 1 9 2 13 15 14 9 3 2
25 2 13 10 9 2 2 13 11 2 2 13 9 15 2 14 9 11 2 7 13 0 1 9 15 2
7 7 9 1 9 9 10 2
7 7 13 1 16 14 13 2
24 13 15 10 9 0 1 9 7 9 7 1 9 14 9 1 9 2 7 9 14 9 1 9 2
6 13 0 1 1 9 2
23 1 10 9 2 14 13 9 1 12 9 14 13 9 9 0 14 9 1 10 9 1 9 2
9 7 13 3 3 3 1 9 9 2
6 13 15 13 9 15 2
184 12 1 9 9 12 2 16 9 15 2 8 14 13 10 9 7 9 1 9 12 1 9 12 1 9 1 9 9 1 9 9 2 1 9 9 15 7 15 13 0 1 9 9 2 1 9 9 0 1 9 10 12 9 1 11 2 12 2 7 1 9 2 1 9 0 2 7 8 14 13 10 9 7 10 9 10 1 9 1 9 0 10 9 9 14 9 1 9 1 9 2 3 2 16 9 15 2 1 9 1 9 9 1 1 9 13 10 9 7 10 9 10 1 9 2 13 9 0 1 9 1 10 9 9 10 9 9 2 13 0 9 10 9 7 9 1 9 10 14 13 1 9 1 9 1 9 9 12 12 7 9 14 13 1 10 9 8 12 12 1 9 13 15 8 9 9 7 9 9 0 10 9 9 1 9 9 16 13 9 12 12 1 9 2
60 16 13 9 10 9 11 1 9 10 11 14 9 13 0 13 1 10 12 9 7 13 0 14 13 11 11 1 9 14 0 1 9 1 10 9 9 16 3 0 14 14 13 11 1 11 1 12 9 1 9 7 10 9 1 9 12 9 1 15 2
20 14 13 10 9 1 3 14 13 9 1 9 1 16 10 9 9 7 10 9 2
38 14 11 14 9 13 10 9 1 1 14 13 15 15 1 9 0 1 9 2 1 9 2 1 9 7 1 9 0 7 14 13 15 15 10 9 14 0 2
5 13 9 1 3 2
8 16 13 15 13 9 14 9 2
29 2 13 15 12 9 10 9 9 1 11 1 9 10 9 1 9 7 12 9 10 9 3 1 9 1 9 1 11 2
25 2 13 1 9 3 14 13 11 1 10 11 9 10 9 0 14 13 11 11 1 9 1 11 11 2
35 13 15 1 9 1 10 9 7 13 15 15 1 9 14 0 1 9 15 2 13 13 9 1 16 1 9 9 3 1 9 1 9 15 9 2
3 13 3 2
51 14 13 15 1 13 10 9 7 9 14 13 1 9 0 10 1 9 1 10 9 9 1 10 9 1 9 9 1 11 2 1 9 1 10 9 14 13 1 9 1 9 10 9 3 3 1 9 10 12 11 2
15 14 13 15 1 9 1 16 15 14 9 1 9 1 9 2
32 15 14 13 15 1 9 11 11 14 9 2 16 9 9 14 9 1 2 14 13 15 0 15 14 9 7 13 10 9 0 9 2
22 1 1 9 1 11 8 15 9 9 7 9 1 9 10 9 3 7 13 15 3 8 2
5 11 2 9 9 2
30 12 13 0 9 14 9 1 9 1 9 1 9 3 2 9 14 0 7 13 15 9 10 9 14 9 1 9 3 3 2
27 3 13 15 13 9 1 9 0 14 13 1 9 1 2 7 9 7 9 1 1 14 13 7 14 9 3 2
15 2 11 11 2 9 14 13 9 1 1 9 9 1 11 2
10 14 13 10 9 14 13 9 10 9 2
31 13 1 10 9 14 11 2 13 10 9 11 1 9 14 13 15 14 0 1 10 9 1 8 7 10 2 9 2 1 8 2
50 13 9 1 9 9 1 9 11 7 13 9 1 14 13 10 9 9 0 1 9 9 2 16 14 13 9 0 15 7 14 13 15 3 3 1 9 14 13 15 3 2 11 2 12 2 12 2 12 2 2
42 13 9 0 1 11 2 9 9 10 9 0 2 1 10 9 1 9 0 3 7 13 10 11 1 9 14 13 9 9 14 9 1 16 13 10 9 2 0 2 1 9 2
42 9 9 0 3 13 11 10 9 16 14 13 15 1 12 8 2 13 15 1 12 9 1 9 2 7 1 12 9 1 9 9 14 13 15 10 12 8 9 1 12 9 2
19 1 9 11 2 13 11 11 1 9 9 0 1 9 10 9 7 10 9 2
18 15 0 10 12 9 3 14 13 10 9 10 1 10 9 1 9 9 2
16 13 15 9 1 9 10 11 14 13 9 7 9 1 9 0 2
6 16 13 13 14 13 2
20 13 10 9 2 9 12 2 16 14 13 10 9 10 1 9 1 12 7 12 2
19 13 9 1 14 13 9 1 1 9 2 1 16 13 1 15 1 10 9 2
15 3 13 10 9 12 9 1 9 13 9 1 1 9 10 2
6 13 11 1 9 12 2
9 2 3 1 14 13 15 1 9 2
19 7 1 10 9 13 15 15 1 10 9 1 9 7 15 1 10 9 0 2
15 13 9 1 10 9 7 13 9 1 10 9 1 10 9 2
35 1 9 10 9 14 13 1 13 11 11 2 11 11 2 11 14 11 2 11 11 2 11 11 2 11 14 11 2 11 11 2 7 11 11 2
22 7 1 14 12 10 9 13 10 9 9 11 14 11 1 9 1 9 1 9 0 8 2
8 13 10 9 14 13 10 9 2
5 14 13 8 15 2
6 10 9 3 14 0 2
55 10 9 0 14 13 10 9 1 9 1 9 7 1 9 7 1 10 9 9 7 9 2 13 10 9 9 14 9 2 9 14 9 2 9 14 9 2 9 0 14 9 7 9 14 9 1 10 9 10 14 13 1 9 1 2
35 16 13 15 1 10 9 1 9 9 13 9 1 11 11 1 9 9 1 13 11 11 2 0 1 9 11 2 9 0 1 9 1 9 10 2
11 3 2 13 0 1 10 9 14 9 3 2
26 13 0 1 14 13 9 0 1 14 13 1 9 15 7 13 9 1 14 13 15 9 1 9 9 0 2
6 13 10 9 1 11 2
14 13 10 9 7 9 1 9 1 9 1 9 0 10 2
35 14 13 9 1 10 9 15 13 9 1 10 9 16 13 10 9 1 15 9 14 13 15 1 2 2 15 2 15 3 14 9 0 10 9 2
7 2 14 13 9 1 1 2
38 16 14 13 15 9 1 9 1 13 15 10 9 14 13 1 13 10 9 15 1 9 9 14 14 13 9 1 9 14 13 10 9 9 1 9 10 9 2
12 8 11 0 1 9 1 9 7 11 1 9 2
41 13 1 9 1 10 9 10 9 9 14 13 10 9 1 9 9 10 9 1 10 9 11 14 13 1 10 9 0 7 9 7 1 10 9 1 9 9 7 9 9 2
34 11 10 9 1 1 9 2 14 11 1 9 11 2 13 9 1 10 9 3 1 11 7 13 11 1 9 10 9 9 2 8 2 1 2
12 13 10 9 1 11 11 1 9 11 11 3 2
6 8 9 9 1 9 2
4 13 9 15 2
7 13 0 1 9 14 9 2
47 13 9 15 9 14 13 1 2 16 13 1 16 13 9 0 0 2 13 1 9 14 13 15 2 1 14 13 1 9 8 13 9 1 9 15 14 9 1 3 13 0 1 9 1 10 0 2
11 9 2 8 2 1 10 9 12 14 9 2
17 13 10 9 10 13 9 0 10 9 10 1 9 10 12 9 9 2
41 13 11 1 9 14 0 1 9 1 12 7 12 7 14 13 3 0 15 1 14 13 10 9 1 9 1 10 9 13 0 1 9 2 16 1 11 1 11 9 9 2
34 7 14 13 9 1 9 1 15 14 13 10 9 7 14 13 3 1 9 1 9 9 9 2 9 9 9 2 1 9 1 10 9 10 2
14 1 9 9 2 9 10 9 0 14 13 9 9 1 2
23 13 15 1 9 1 9 1 9 9 1 9 1 9 0 14 13 9 9 1 10 9 0 2
35 13 8 1 1 9 7 8 12 9 1 9 9 2 8 13 2 13 2 13 15 8 13 2 13 2 13 15 8 13 2 13 2 13 15 2
29 11 14 13 1 9 1 9 7 9 0 1 9 10 9 10 1 12 9 1 12 2 7 12 9 9 1 9 8 2
4 13 14 0 2
41 9 3 0 1 10 9 0 10 1 9 14 11 2 13 9 11 11 2 9 1 9 1 9 10 9 2 11 2 1 2 11 11 2 11 11 9 9 11 11 2 2
13 16 3 13 10 9 10 14 0 1 0 7 0 2
34 7 2 1 9 1 9 2 13 0 10 9 14 13 15 1 9 14 11 1 9 10 9 9 2 14 9 14 13 15 15 1 12 9 2
24 6 2 13 9 0 1 9 0 10 9 3 15 7 9 10 9 0 1 9 10 9 1 12 2
29 13 1 12 7 15 1 9 1 10 9 1 9 11 2 8 11 7 1 9 1 9 1 14 13 1 9 1 8 2
9 13 9 0 1 9 1 10 9 2
16 14 13 15 1 9 9 0 1 9 14 9 14 0 10 9 2
24 2 1 10 9 0 2 13 9 10 9 0 14 13 1 9 1 10 9 9 1 9 1 9 2
28 1 9 1 15 13 9 0 1 10 11 11 7 13 15 10 9 2 14 9 9 7 10 9 15 1 10 9 2
40 13 9 1 9 15 9 9 14 13 1 10 9 10 1 9 14 13 0 1 12 9 2 9 2 12 9 7 9 14 13 10 9 9 1 7 14 13 1 9 2
15 15 9 13 1 1 9 1 9 10 1 9 13 3 1 2
20 13 10 9 11 9 0 1 9 9 14 13 0 1 9 9 1 9 9 9 2
25 2 13 0 14 13 9 1 10 9 15 14 9 1 10 9 7 9 14 13 1 9 15 14 9 2
15 13 1 10 9 1 9 12 13 1 9 12 2 13 1 2
23 13 9 1 11 7 1 10 9 2 11 2 1 9 10 9 2 3 12 9 3 1 9 2
17 14 13 15 1 1 14 13 10 9 9 10 9 9 14 13 15 2
57 13 1 9 14 13 10 10 9 1 10 9 1 9 2 7 1 9 1 9 13 0 9 9 14 9 1 9 2 7 9 0 7 10 9 2 16 13 9 0 10 9 0 1 10 10 9 1 14 12 9 7 12 9 9 1 9 2
127 13 15 15 10 2 9 9 2 1 9 1 9 1 10 9 9 14 13 9 0 9 12 3 7 1 10 9 9 15 15 10 9 1 9 1 9 10 2 9 2 1 9 2 9 12 3 2 13 0 10 9 2 13 15 1 9 10 2 9 2 14 9 14 13 2 10 2 9 1 9 2 7 1 9 0 2 2 13 15 9 14 13 0 1 9 14 9 9 0 2 14 13 10 9 14 0 3 0 2 13 15 10 9 3 1 7 13 15 1 9 1 9 1 9 2 13 15 9 1 9 0 1 9 1 10 9 2
6 13 11 1 11 3 2
33 15 10 9 2 13 0 14 13 1 9 14 0 1 9 10 8 2 13 13 1 11 14 13 9 12 1 10 9 10 1 10 11 2
13 15 10 14 13 1 9 1 2 1 9 13 3 2
6 10 9 14 13 11 2
3 10 8 2
9 16 13 0 2 9 0 13 1 2
4 16 13 15 2
8 8 10 9 3 2 14 11 2
7 15 14 14 13 10 9 2
10 15 13 1 14 12 0 14 13 1 2
16 16 3 13 9 9 13 1 9 16 13 9 0 1 8 3 2
16 8 2 12 8 2 14 13 11 2 9 12 2 1 9 8 2
9 2 8 10 9 14 0 1 9 2
9 2 2 15 14 13 10 9 1 2
12 2 2 6 2 13 15 3 0 8 1 9 2
5 14 0 1 9 2
10 9 9 1 9 2 9 2 12 2 2
36 8 13 1 15 9 12 2 9 8 2 1 14 13 2 1 9 8 2 9 12 2 13 10 9 2 8 2 8 2 8 1 10 9 1 9 2
38 13 9 7 12 1 3 1 9 13 10 2 8 2 3 1 1 9 14 13 10 9 1 16 1 14 13 9 14 13 1 9 3 3 1 10 9 0 2
7 1 12 9 1 14 9 2
50 10 9 14 13 15 2 7 13 15 0 14 13 9 9 1 16 14 13 15 13 11 14 13 1 9 1 2 7 9 11 7 9 2 16 9 0 2 16 1 9 7 9 9 2 10 9 0 2 2 2
9 2 8 2 16 14 13 15 15 2
32 13 9 7 9 10 9 1 11 1 12 9 3 1 10 9 1 9 2 1 13 8 1 12 1 10 9 14 0 1 10 9 2
21 14 0 7 14 13 10 9 13 9 0 0 3 1 15 1 9 9 14 9 1 2
23 7 13 0 9 0 0 0 14 13 15 10 9 9 16 14 13 15 1 10 9 10 1 2
24 13 15 3 10 9 10 7 9 1 14 13 10 9 3 1 9 9 1 14 12 10 9 9 2
6 9 14 0 14 9 2
12 1 12 2 3 2 13 9 1 9 9 9 2
40 11 11 2 9 2 9 2 14 9 2 7 13 11 14 13 1 9 1 9 9 14 11 9 7 13 15 15 15 1 9 9 2 9 14 9 10 9 1 9 2
19 13 15 9 1 3 0 7 14 13 15 7 3 0 3 7 14 13 15 2
17 13 9 9 0 14 9 1 12 9 2 1 9 0 7 9 0 2
17 2 9 2 14 13 10 9 10 9 2 13 1 7 14 13 3 2
15 2 6 13 9 1 2 13 11 2 15 7 10 9 9 2
30 9 2 8 13 9 0 1 10 9 10 2 7 13 9 1 9 0 9 7 9 0 9 0 1 9 3 0 14 9 2
41 9 1 9 9 1 9 9 1 11 14 11 0 1 9 9 10 11 0 11 12 13 15 9 9 10 11 14 13 10 9 9 10 1 11 14 11 1 9 10 9 2
13 13 9 2 3 2 10 9 9 14 9 1 9 2
13 2 1 13 15 3 1 9 2 2 14 13 11 2
33 2 13 9 10 9 9 1 9 1 9 2 11 11 2 1 11 11 7 8 9 10 3 9 9 1 9 9 9 14 9 1 9 2
31 1 10 9 14 13 1 13 9 9 2 11 11 2 11 11 2 11 11 2 11 11 11 7 9 10 1 9 0 10 9 2
9 2 7 9 10 3 1 11 11 2
16 16 13 9 14 0 2 14 13 10 9 0 9 9 1 15 2
16 9 1 10 9 2 9 10 9 0 2 0 2 1 9 0 2
32 2 1 9 10 2 9 10 9 16 0 10 9 2 13 9 0 1 7 13 15 1 9 14 13 10 9 1 9 9 1 9 2
16 13 12 1 11 15 2 9 13 3 0 1 9 10 11 3 2
28 13 10 9 14 11 10 9 14 13 9 1 9 7 9 7 9 1 9 9 7 11 1 9 10 12 9 9 2
52 13 1 9 14 13 15 9 2 13 10 9 0 2 7 14 0 10 9 14 13 1 10 9 1 9 1 9 0 2 1 9 1 10 9 7 10 9 2 7 13 9 16 14 13 14 0 1 9 15 2 2 2
12 1 10 12 9 3 2 13 10 9 0 1 2
2 11 2
3 2 2 2
10 16 13 9 0 9 1 10 9 10 2
6 16 14 13 9 1 2
6 11 2 13 0 15 2
9 1 9 2 1 9 2 1 9 2
20 15 1 3 15 2 2 7 15 1 9 15 1 9 14 13 9 10 9 1 2
27 14 9 1 15 9 13 1 9 1 14 9 1 9 7 13 3 1 9 9 1 11 1 9 7 1 10 2
11 3 14 13 11 2 11 1 10 9 10 2
10 14 13 3 1 11 13 15 1 15 2
10 16 13 15 2 9 1 9 9 3 2
4 2 12 2 2
14 2 16 14 13 15 0 13 9 1 9 1 9 1 2
2 8 2
22 13 9 1 14 13 1 9 10 9 16 9 0 1 9 9 2 9 2 9 7 9 2
38 2 2 3 2 14 11 2 2 14 13 15 2 2 13 15 1 9 10 9 10 1 9 14 9 9 0 16 13 9 13 9 10 14 13 1 1 9 2
17 13 15 13 1 9 1 10 9 0 14 9 13 9 9 15 2 2
13 9 0 7 15 13 15 9 0 14 13 1 15 2
11 2 16 13 10 12 9 1 1 9 8 2
42 11 1 9 9 9 0 1 9 2 15 1 9 0 9 0 9 7 13 0 1 2 10 10 9 0 1 10 9 1 9 7 9 1 9 10 9 1 9 9 0 1 2
9 1 9 1 9 13 11 3 3 2
16 13 0 1 9 16 10 9 2 11 11 2 7 11 14 11 2
37 16 13 11 0 7 15 1 9 10 9 7 10 9 1 9 1 10 9 2 10 8 1 10 9 1 9 10 9 9 1 9 1 9 1 10 9 2
28 2 13 15 9 1 10 9 0 16 13 15 1 9 12 7 3 9 9 10 14 9 3 16 13 10 9 9 2
7 14 13 9 0 1 9 2
26 13 1 9 13 15 13 0 1 9 0 1 14 13 2 9 2 2 9 14 13 0 1 9 14 0 2
37 13 9 1 14 13 14 0 1 1 11 1 9 9 7 16 9 1 9 9 8 10 9 0 1 9 10 14 9 1 9 13 1 2 1 9 9 2
20 16 13 9 7 9 1 9 14 13 1 9 1 9 13 10 9 9 1 9 2
20 2 11 2 2 13 11 7 2 1 9 10 9 1 9 11 2 13 15 1 2
25 13 10 9 1 11 14 13 10 9 1 9 1 3 1 9 9 14 13 9 0 1 1 10 9 2
5 13 15 15 0 2
15 1 10 9 0 15 14 13 10 9 14 13 1 9 15 2
48 16 14 13 15 3 2 13 9 7 9 15 14 0 1 9 1 10 9 2 14 13 9 0 0 1 16 14 13 1 15 2 1 9 3 1 9 2 1 9 1 9 9 9 1 2 13 1 2
66 7 14 13 1 2 2 13 15 2 2 7 13 15 1 9 2 7 3 2 3 14 13 15 2 2 13 15 2 2 7 13 15 14 9 3 3 1 10 9 2 2 13 15 2 2 1 9 2 1 9 1 9 2 2 13 15 2 2 14 13 15 1 9 10 9 2
36 2 10 9 13 0 14 13 10 9 1 10 9 2 2 14 13 11 2 2 16 0 7 0 15 2 14 13 10 9 10 10 9 1 9 0 2
124 9 12 9 0 13 8 7 9 9 0 2 2 9 14 9 1 9 9 7 1 9 9 1 9 10 7 2 16 0 2 1 9 0 2 2 10 9 9 9 0 7 9 0 14 9 7 14 9 1 9 7 9 2 13 10 9 2 9 9 0 2 9 7 10 9 10 1 9 10 9 7 1 9 9 2 13 0 15 9 14 13 15 2 2 10 9 7 13 1 9 10 14 9 7 14 9 2 2 10 9 9 9 14 9 1 9 1 9 9 7 1 9 0 14 13 9 1 9 14 9 7 14 9 2
44 13 9 10 11 11 2 10 9 1 11 7 11 1 9 3 1 11 10 11 3 0 1 9 9 13 1 11 7 11 11 10 9 14 13 10 9 11 11 8 9 14 9 0 2
26 2 9 2 16 13 9 1 3 2 13 1 9 2 16 1 10 9 10 13 10 9 9 1 10 9 2
8 16 13 15 15 14 13 15 2
28 2 16 15 1 14 13 14 9 14 13 9 7 9 1 10 11 10 1 11 11 7 11 2 11 11 14 11 2
7 2 9 1 9 13 1 2
18 9 9 11 2 11 11 2 11 11 2 11 2 11 11 7 8 11 2
9 2 3 13 9 1 15 14 9 2
11 16 3 14 13 15 2 10 9 14 9 2
13 16 13 15 10 10 9 1 9 14 13 1 9 2
19 2 14 9 1 13 15 10 9 1 15 13 9 10 9 16 13 0 1 2
4 13 15 11 2
24 2 13 10 9 10 9 1 1 9 10 9 1 9 2 9 7 9 0 2 2 14 13 11 2
26 3 10 14 0 10 9 14 13 10 9 1 9 10 11 9 10 10 9 0 14 9 3 0 10 1 2
8 13 15 13 0 10 9 10 2
21 16 13 1 10 9 2 15 13 0 9 0 14 9 1 9 1 15 14 13 15 2
28 13 10 9 1 9 1 11 12 1 10 11 11 1 9 10 1 7 15 1 9 3 1 11 12 2 12 2 2
13 9 0 1 9 12 1 11 2 13 15 0 1 2
11 13 0 14 13 9 1 15 15 14 13 2
16 13 9 9 1 1 9 14 9 1 9 10 9 14 9 1 2
7 11 1 9 9 0 11 2
7 15 14 13 15 1 11 2
12 13 15 7 13 15 10 9 1 9 1 15 2
12 16 9 1 11 11 13 9 10 9 10 0 2
24 13 15 9 0 1 9 11 1 9 1 9 9 7 9 14 13 10 9 1 15 1 9 11 2
27 13 3 15 1 9 14 13 9 10 9 14 10 9 2 12 2 2 7 1 9 10 9 10 2 12 2 2
35 1 9 10 9 13 15 13 10 9 16 13 15 14 9 1 9 3 1 9 3 2 9 14 13 1 9 16 9 10 9 7 1 9 0 2
10 3 13 0 16 14 13 10 9 1 2
15 11 15 10 9 7 13 1 9 1 10 9 1 10 9 2
20 10 9 14 13 15 3 0 2 16 3 14 13 15 15 7 13 15 1 9 2
10 9 10 9 13 9 9 1 11 11 2
48 13 15 15 9 9 0 1 9 1 10 9 7 1 9 2 13 0 14 13 12 0 9 0 1 7 14 13 15 15 10 9 9 9 13 0 16 13 8 1 1 15 16 9 7 9 1 9 2
31 9 0 1 9 10 9 14 13 1 9 9 1 2 1 9 9 2 1 9 9 7 9 2 1 9 2 13 15 0 3 2
26 2 9 2 7 2 9 2 1 2 10 9 2 7 2 10 9 2 14 13 1 10 9 7 10 9 2
29 13 15 1 9 10 9 7 1 9 1 9 1 9 9 14 9 7 14 0 13 9 10 9 1 9 1 10 9 2
24 13 9 1 14 11 11 1 9 12 7 3 1 9 2 13 15 1 9 1 9 1 11 3 2
38 16 13 9 1 10 9 1 9 2 7 16 13 10 9 15 1 10 9 13 3 13 2 13 15 1 9 1 9 2 16 0 0 10 9 1 9 15 2
19 14 13 9 1 9 1 10 9 15 15 1 9 0 14 9 1 9 1 2
52 1 9 0 10 13 11 0 12 9 1 9 1 7 13 1 15 14 13 2 1 9 12 13 9 10 9 9 1 9 10 9 1 9 7 9 3 1 9 10 9 14 13 10 9 10 1 9 14 9 1 9 2
25 13 1 9 14 13 9 9 3 0 3 3 7 13 15 1 9 2 7 10 9 10 9 0 1 2
25 13 11 14 0 7 9 1 9 1 9 11 11 2 11 12 2 1 9 2 1 9 7 1 9 2
259 8 1 9 9 8 1 9 10 2 14 13 10 9 14 14 13 1 9 10 1 9 2 8 1 9 9 1 9 14 13 1 9 8 2 8 7 8 1 9 8 1 9 10 9 0 2 8 1 9 14 13 10 9 9 1 15 15 1 9 7 13 15 10 9 14 0 7 1 9 10 9 9 7 13 0 7 12 9 9 0 7 9 9 0 10 9 2 16 1 2 7 10 9 14 13 15 2 7 12 9 1 9 14 13 10 9 13 15 9 10 9 15 2 7 8 1 10 9 10 2 7 9 1 9 14 13 10 9 13 15 9 10 9 15 2 8 1 9 9 1 9 14 13 1 9 8 1 9 8 1 9 10 2 7 9 1 9 14 13 10 9 13 15 9 10 9 15 2 8 1 9 9 1 9 14 13 1 9 8 1 9 8 1 9 10 2 7 8 1 9 9 1 9 14 13 1 9 8 1 9 8 1 9 10 2 7 8 1 9 9 14 13 9 0 7 12 9 1 2 7 12 9 2 8 1 9 9 14 13 12 9 1 2 7 12 7 12 9 2 7 8 1 9 9 14 13 12 9 7 9 0 1 2 7 12 7 12 9 2
10 2 15 9 9 13 1 9 3 3 2
28 13 9 1 9 1 10 8 1 9 9 7 9 10 9 7 9 7 13 3 14 0 14 13 7 14 13 15 2
27 1 11 13 12 9 1 9 3 2 16 13 9 1 9 1 9 0 8 1 8 2 7 1 8 1 8 2
16 10 9 16 9 2 13 15 14 9 7 14 13 15 3 1 2
8 3 3 13 9 0 1 11 2
132 8 1 9 9 14 9 2 10 9 14 13 9 1 1 9 1 9 10 14 13 1 9 1 9 16 1 10 7 1 9 16 13 1 9 8 7 2 16 16 14 13 2 16 1 7 1 9 9 10 9 13 1 9 14 13 1 9 15 1 9 8 2 2 10 9 2 2 2 13 9 1 7 13 9 1 16 1 10 7 1 9 10 7 2 16 16 14 13 2 16 1 10 7 1 9 2 16 14 13 9 1 7 9 1 9 1 9 10 9 10 14 13 16 15 1 9 10 9 14 13 1 10 9 10 1 9 1 10 9 0 10 2
21 3 0 1 15 2 13 9 14 11 1 10 9 0 9 9 9 0 1 10 9 2
54 13 3 1 9 0 10 9 15 7 13 11 2 1 9 11 0 2 7 11 1 11 2 9 1 1 9 10 9 1 9 9 2 10 9 9 0 13 1 9 1 2 9 9 2 9 0 2 9 2 9 2 8 2 2
12 13 15 3 8 0 2 9 2 2 1 9 2
12 13 15 1 10 9 9 7 10 9 14 0 2
39 10 9 0 0 13 0 1 9 0 10 14 13 9 7 9 16 0 1 9 7 9 0 10 9 2 7 1 14 13 15 9 1 9 14 9 14 0 0 2
27 16 13 1 9 10 9 14 13 15 1 9 15 1 10 9 14 13 15 1 7 15 1 9 1 9 15 2
42 13 15 0 14 0 2 1 15 2 14 13 11 1 9 9 9 11 1 12 12 9 3 14 9 2 13 15 1 9 1 8 12 1 8 2 9 10 9 2 11 0 2
25 2 9 0 1 9 11 2 0 2 14 13 1 9 1 10 9 2 14 14 13 9 0 10 11 2
5 13 15 3 9 2
10 14 0 2 13 10 9 1 12 9 2
80 16 13 9 9 7 9 9 1 11 1 9 1 9 1 2 9 2 1 9 1 11 2 16 13 8 1 9 1 9 1 8 1 9 10 9 9 11 1 9 0 8 1 10 9 2 9 13 1 9 14 9 1 9 10 9 14 11 2 13 1 2 13 0 9 3 1 10 9 1 9 14 13 9 10 9 1 11 1 9 2
44 10 12 9 10 14 13 1 9 7 9 14 9 1 9 2 10 9 10 1 2 1 9 9 7 9 1 9 1 9 10 9 10 2 14 13 2 13 3 15 2 1 9 1 2
68 1 9 9 7 9 8 9 10 11 10 9 0 0 9 10 1 2 7 1 14 13 1 9 1 9 1 2 16 14 13 9 0 1 1 9 0 2 14 13 9 10 9 7 10 9 1 10 9 1 2 9 14 13 1 9 1 9 1 3 16 13 1 2 3 0 1 9 2
21 13 9 3 1 9 1 9 1 9 10 9 14 0 7 13 9 1 15 1 9 2
29 9 12 9 14 12 12 16 14 13 10 9 10 0 2 15 14 13 0 1 10 9 11 1 9 1 0 2 9 2
16 10 9 11 2 9 2 9 0 7 1 9 10 1 10 9 2
16 13 15 9 10 0 1 2 16 15 14 13 3 1 10 9 2
32 13 10 9 14 11 1 1 9 14 13 10 9 10 1 1 10 9 1 12 1 9 9 3 1 9 1 10 9 9 1 9 2
32 13 15 14 0 1 10 9 7 13 15 3 9 8 1 10 9 13 9 0 1 7 13 10 9 9 1 14 13 9 10 9 2
38 2 13 9 11 1 9 12 9 1 9 1 10 9 3 16 13 9 16 13 9 1 9 11 0 1 8 9 1 9 1 9 7 16 13 9 1 9 2
11 16 14 13 10 9 0 0 10 16 9 2
47 13 9 1 2 7 1 16 14 13 10 9 1 9 13 10 9 1 9 9 1 9 1 9 7 16 14 13 9 9 9 14 13 0 1 9 16 12 9 1 9 7 12 9 10 1 9 2
39 9 1 9 14 9 1 9 0 0 9 1 9 2 9 1 9 0 14 13 1 2 14 13 16 13 15 2 13 15 10 10 9 7 13 15 1 9 9 2
308 10 9 1 9 9 1 14 13 3 1 9 0 2 1 9 2 13 9 0 1 9 9 10 9 9 2 10 9 7 10 9 1 7 13 15 0 1 9 9 1 3 9 9 1 9 1 9 9 2 1 9 2 13 10 9 1 9 13 1 9 1 9 16 14 13 15 1 9 0 9 9 9 14 13 9 1 10 9 2 13 15 9 9 9 0 7 3 1 12 9 1 10 9 2 16 13 15 1 9 9 0 1 9 2 1 9 1 9 14 13 10 9 2 13 10 9 10 9 1 9 7 13 15 1 10 9 1 9 9 0 2 3 1 9 0 1 9 2 14 13 10 9 1 0 14 13 1 9 10 2 13 9 9 14 9 1 9 9 2 9 7 9 10 9 1 14 13 9 1 9 2 13 15 15 2 10 9 9 14 13 1 10 9 2 13 15 10 9 8 10 9 9 9 1 9 14 13 9 7 14 13 9 1 2 13 9 9 14 9 1 10 10 9 7 9 2 13 10 9 9 2 9 7 9 1 9 3 1 12 9 9 2 13 9 9 0 14 9 1 9 10 1 9 7 9 9 0 13 15 9 0 10 9 7 0 2 0 7 0 2 13 9 0 16 14 13 10 12 9 1 9 1 9 2 16 14 13 12 9 0 1 9 13 9 1 10 9 0 2 9 9 2 9 7 9 2 13 15 9 0 9 7 0 2 0 7 0 2
51 14 10 9 1 9 13 10 9 2 9 7 9 2 14 13 9 1 9 1 9 0 1 9 10 9 2 9 13 0 14 13 9 9 1 3 2 9 9 2 9 14 13 1 9 0 1 9 0 14 9 2
17 13 15 0 9 9 9 10 9 12 7 1 1 10 9 9 0 2
38 16 9 15 13 9 1 9 10 9 10 9 0 14 9 1 9 10 9 13 1 9 2 13 0 1 10 9 2 10 9 2 14 13 15 0 14 0 2
29 13 9 0 1 9 9 10 11 0 2 1 9 9 0 1 3 12 9 7 3 9 10 9 0 2 8 2 8 2
17 3 16 14 13 10 9 14 13 15 2 7 14 13 15 10 9 2
27 13 9 1 1 9 0 7 9 10 1 9 0 1 9 10 9 14 13 3 1 9 7 14 14 13 9 2
27 13 10 9 10 9 1 10 9 1 9 7 1 9 11 2 11 11 2 11 11 2 11 11 7 10 8 2
27 2 2 14 0 2 13 11 11 2 9 9 10 9 9 9 2 9 16 13 10 9 10 1 9 1 9 2
5 1 11 14 11 2
10 13 10 9 15 1 3 2 1 9 2
23 2 16 13 10 9 10 9 1 2 10 9 14 13 15 3 0 1 10 9 14 13 1 2
18 13 8 0 2 0 7 9 10 9 1 2 16 14 0 1 9 9 2
18 13 15 8 14 0 1 9 16 7 13 1 9 1 16 9 10 9 2
89 8 13 9 1 9 7 1 9 1 9 8 9 1 9 14 9 1 9 9 9 9 7 9 14 13 0 1 7 1 1 9 10 7 13 15 7 15 2 16 13 7 10 9 14 13 10 9 11 3 1 7 1 15 2 9 0 1 9 14 9 1 9 1 12 9 7 9 1 9 10 7 13 15 7 15 1 9 10 9 1 9 10 14 9 1 9 1 11 2
16 7 16 14 13 15 1 9 9 2 13 9 9 14 13 1 2
51 10 9 10 0 13 15 9 0 10 9 1 9 9 7 13 15 1 9 2 9 1 9 2 0 2 1 9 0 2 7 9 1 9 10 9 0 14 13 9 3 0 1 1 2 9 2 7 2 9 2 2
51 13 10 9 1 9 1 1 9 3 2 9 9 0 2 9 10 9 0 2 1 10 9 9 14 9 2 16 14 13 1 9 1 10 9 1 9 0 0 1 9 0 2 9 13 9 1 10 9 14 9 2
27 3 13 15 1 9 1 10 9 2 9 1 10 11 2 10 9 0 0 0 10 14 13 1 11 1 11 2
33 2 16 13 15 10 0 2 9 1 9 1 9 9 9 1 10 9 13 0 14 13 1 9 0 2 7 13 0 1 10 9 10 2
25 14 13 9 7 12 1 15 14 9 1 9 9 16 13 1 10 9 9 9 9 14 13 9 1 2
42 2 13 15 1 9 1 9 13 0 9 14 13 10 9 14 9 9 16 13 9 14 13 15 10 9 9 0 2 16 13 0 15 14 9 1 10 9 1 9 14 9 2
76 16 13 0 2 13 9 0 9 1 13 10 9 0 1 9 9 9 2 1 9 11 11 2 11 11 7 12 9 1 9 10 9 12 1 8 1 15 2 16 14 13 11 9 0 1 10 9 7 10 9 2 13 15 10 9 2 13 2 1 9 1 9 14 13 1 9 1 10 9 2 1 9 14 13 9 2
65 12 10 9 0 14 13 9 1 0 1 9 14 13 7 14 13 9 0 1 9 14 13 1 9 2 13 1 0 9 0 1 9 9 2 13 1 9 14 13 10 9 0 8 2 7 3 10 9 9 14 13 8 9 10 9 1 11 1 10 9 9 10 14 13 2
54 13 1 14 13 15 1 9 1 10 9 13 0 1 8 2 9 9 14 9 1 9 10 11 7 9 1 2 15 1 1 2 9 2 7 9 0 10 9 2 14 13 2 10 9 10 1 9 1 9 7 1 9 2 2
20 9 9 14 13 1 9 9 0 2 1 9 7 1 9 9 7 9 0 0 2
49 2 13 2 1 9 1 8 2 14 13 10 9 9 10 9 9 1 9 0 10 9 7 14 13 9 1 9 2 10 9 7 10 9 9 9 0 2 2 14 13 10 8 11 14 11 2 9 9 2
3 13 15 2
24 1 9 10 9 1 2 13 15 1 11 1 9 0 10 9 7 1 9 1 10 11 11 11 2
18 9 9 9 14 13 1 14 13 1 9 1 9 9 0 9 1 9 2
27 13 10 11 0 1 9 1 9 10 11 14 13 12 12 1 2 1 10 9 2 1 9 1 9 10 11 2
33 16 15 10 9 14 0 14 13 9 1 9 7 13 1 13 0 10 9 9 14 9 1 10 9 14 13 3 0 1 10 9 0 2
61 1 9 13 9 1 9 0 1 10 9 10 2 13 11 9 0 1 10 11 1 9 14 9 1 9 9 2 9 14 13 2 9 15 2 9 1 9 0 10 9 2 7 13 15 10 9 10 3 1 9 0 7 0 14 9 1 10 9 1 9 2
57 13 0 2 13 0 7 13 0 10 9 14 13 11 1 9 9 10 9 2 10 8 1 9 2 1 9 14 13 15 0 1 9 2 7 1 9 13 1 9 1 10 9 9 14 0 1 9 7 9 9 2 14 0 2 11 11 2
19 1 9 10 9 10 0 2 13 9 0 1 1 9 7 9 10 9 3 2
19 8 13 9 1 9 10 9 2 7 13 0 15 1 10 9 9 3 0 2
35 13 15 0 1 9 9 9 14 9 1 9 9 1 9 0 0 14 13 1 9 1 10 9 1 9 10 11 1 11 11 2 12 9 9 2
16 14 13 1 13 15 10 9 0 15 1 11 10 12 9 10 2
16 12 13 10 12 9 1 11 7 13 1 12 1 9 14 9 2
16 2 13 15 10 9 3 3 0 7 14 13 1 10 9 15 2
29 7 14 13 15 1 10 9 10 16 14 13 15 1 10 9 9 14 13 1 9 10 9 14 13 11 1 9 1 2
36 13 9 1 16 9 1 9 10 12 9 14 8 1 12 7 12 7 14 13 1 10 12 9 9 2 1 9 14 9 1 9 1 10 9 0 2
20 2 13 9 1 8 10 9 14 13 10 9 2 16 1 10 9 13 10 9 2
37 8 1 10 9 9 0 14 9 0 2 13 9 14 14 13 1 9 10 9 7 9 14 13 1 10 9 10 16 14 13 14 9 1 9 9 0 2
17 13 10 9 1 14 0 7 2 14 0 2 9 9 9 10 9 2
24 13 15 0 15 16 13 1 9 1 10 12 9 0 10 1 14 13 1 9 10 11 1 9 2
28 1 9 2 1 9 2 14 13 9 1 3 2 7 9 14 0 1 9 10 1 9 2 7 13 10 10 9 2
7 13 0 1 9 14 9 2
14 13 10 9 9 1 9 1 2 13 10 9 0 0 2
7 13 9 1 9 1 8 2
28 13 0 9 10 9 14 9 1 9 2 1 9 9 1 9 14 0 2 1 9 1 10 9 7 10 9 9 2
32 13 15 14 13 9 9 1 9 1 11 7 14 13 15 15 14 13 9 0 10 9 14 9 14 0 7 15 9 3 1 9 2
25 14 13 10 9 9 1 9 1 7 13 0 13 0 1 15 2 16 13 9 1 9 14 9 1 2
11 14 13 14 11 9 11 1 9 1 9 2
15 13 9 1 9 7 9 1 9 14 13 1 9 10 8 2
15 1 9 7 13 1 9 0 14 13 10 9 1 9 3 2
39 16 1 9 16 14 13 15 14 9 13 9 1 9 10 9 3 7 13 15 1 9 1 9 1 7 16 14 13 10 9 0 14 13 15 1 1 10 9 2
43 13 15 9 10 9 1 9 1 9 7 13 15 9 9 1 9 9 10 9 1 9 1 10 9 1 9 9 10 9 7 1 9 10 9 1 9 10 9 1 9 10 9 2
40 13 9 1 9 1 9 9 10 11 1 9 9 2 0 1 9 12 2 1 9 11 0 2 13 10 9 10 1 9 14 9 1 10 9 10 1 9 10 2 2
20 13 10 11 11 13 0 10 11 14 9 1 15 14 13 10 11 1 9 1 2
40 13 1 9 10 13 0 1 11 14 9 0 1 10 9 1 9 14 13 15 9 10 9 1 11 14 9 1 9 9 10 9 10 1 9 14 9 1 10 9 2
8 9 7 9 13 0 14 13 2
29 16 13 10 9 10 16 13 9 9 2 13 9 14 13 15 9 0 10 9 16 13 15 0 9 10 9 14 9 2
29 2 1 10 9 0 13 9 9 1 9 2 7 14 13 10 9 1 15 10 9 13 1 9 1 10 11 14 9 2
21 9 7 9 0 0 2 9 0 0 2 10 9 0 1 9 0 1 9 10 9 2
17 11 9 3 13 9 9 1 9 1 9 0 10 9 1 9 9 2
34 13 0 14 13 1 10 9 10 2 16 13 15 1 9 14 13 1 9 1 9 1 10 9 10 2 7 13 9 10 9 10 1 1 2
27 13 10 9 1 10 9 2 3 2 14 13 15 9 0 7 13 10 9 13 9 9 14 9 1 10 9 2
33 13 9 10 9 2 11 11 1 11 1 11 2 14 13 12 9 9 1 9 1 9 1 10 9 1 9 2 16 13 1 10 9 2
38 10 9 10 1 9 10 11 13 15 15 7 11 11 9 9 1 9 1 10 9 9 14 0 9 14 13 1 9 1 13 9 11 2 11 7 11 1 2
5 13 9 0 15 2
10 13 15 10 9 14 13 15 1 11 2
5 15 9 9 10 2
5 13 14 13 1 2
5 13 0 9 15 2
5 13 11 10 9 2
35 13 10 9 15 1 9 1 2 10 9 0 14 0 1 9 10 9 2 9 7 9 2 9 0 1 10 9 7 10 9 10 1 9 1 2
30 13 15 9 9 1 9 1 10 9 1 15 16 13 15 3 1 9 0 1 9 12 16 14 13 15 12 9 1 9 2
6 13 10 9 1 9 2
6 7 1 1 9 1 2
12 13 15 10 9 11 10 9 1 9 1 11 2
12 13 15 14 13 15 10 9 10 3 0 15 2
6 2 13 0 1 15 2
12 9 1 9 0 10 2 10 9 0 1 15 2
6 13 0 9 7 9 2
20 13 15 10 9 3 1 9 9 14 13 10 9 0 3 1 9 9 1 11 2
7 13 10 9 1 10 9 2
7 14 13 9 10 9 1 2
7 13 9 1 10 9 1 2
7 9 10 9 14 13 1 2
16 13 10 9 1 13 1 9 10 9 14 13 10 9 9 0 2
8 3 1 10 9 1 9 0 2
8 13 10 9 12 1 9 11 2
8 13 15 1 9 1 9 10 2
25 13 15 10 9 14 13 10 9 0 1 9 7 14 13 15 10 9 14 13 14 11 1 2 9 2
17 13 9 0 0 0 1 9 0 7 1 9 1 9 10 9 0 2
10 13 0 9 14 13 1 9 1 8 2
20 2 13 0 1 10 9 9 14 9 7 10 9 14 9 1 10 9 1 9 2
11 2 2 9 9 10 11 2 2 8 2 2
24 13 3 14 13 10 9 1 9 10 9 1 9 1 9 2 9 14 13 10 9 10 1 9 2
12 13 9 9 15 14 0 14 13 15 1 11 2
9 13 10 9 1 9 1 10 9 2
7 13 9 14 13 9 1 2
4 14 13 11 2
5 13 14 0 15 2
12 2 16 13 15 14 9 1 9 1 10 9 2
7 2 14 13 15 10 9 2
12 14 13 10 9 1 9 1 9 1 10 9 2
5 12 9 9 9 2
8 13 15 1 9 11 1 11 2
5 13 11 7 9 2
81 3 1 9 1 9 1 9 10 9 14 13 9 11 1 11 1 9 1 1 10 9 0 13 9 3 2 2 13 10 9 2 8 11 11 11 1 9 2 8 9 2 9 9 2 8 2 8 2 2 13 10 9 7 10 9 1 9 1 9 1 9 1 9 14 9 1 9 2 13 13 15 10 10 12 9 1 9 9 9 1 11
61 13 1 15 2 1 9 14 9 1 1 9 0 1 10 9 14 9 1 9 14 8 9 1 9 1 15 1 11 11 1 9 10 9 3 16 14 13 10 9 2 14 13 9 7 12 1 1 10 9 2 1 9 14 0 1 9 9 1 11 11 2
40 2 16 13 9 9 2 16 13 1 10 9 2 13 7 13 2 10 9 0 2 2 10 9 14 13 9 10 9 10 1 1 10 9 1 15 2 1 12 9 2
16 9 1 11 14 11 14 13 10 9 2 11 11 9 1 11 2
24 2 7 2 14 11 2 13 15 10 9 0 2 2 2 10 9 0 2 0 0 2 14 11 2
16 13 1 7 1 2 3 2 9 1 10 9 1 1 13 9 2
40 2 8 2 14 13 9 1 9 8 1 9 14 13 1 9 9 0 1 9 1 9 1 9 14 13 1 9 12 8 1 9 1 9 9 11 11 11 2 12 2
27 13 1 9 9 9 14 0 14 13 9 1 9 7 9 9 2 16 13 9 10 1 9 9 1 2 3 2
38 12 9 9 10 12 9 2 13 9 14 9 2 16 13 9 10 1 15 10 9 2 7 13 13 1 9 16 14 13 7 14 13 1 9 0 10 9 2
19 1 15 13 11 11 11 2 9 14 13 1 9 1 11 1 9 10 9 2
11 13 10 9 14 13 3 15 1 14 0 2
25 2 2 13 11 15 12 9 1 9 9 2 1 11 11 1 12 7 1 12 2 12 10 12 9 2
14 13 10 9 9 10 1 0 3 3 1 9 11 11 2
29 1 14 9 0 1 10 11 13 11 1 10 9 16 14 13 7 13 1 9 9 1 9 14 13 1 9 1 3 2
32 13 11 7 9 11 16 3 1 9 1 9 1 9 7 13 9 0 11 2 11 2 16 3 1 9 1 9 10 9 1 9 2
44 13 10 9 0 16 10 9 1 10 9 11 14 11 7 10 9 11 14 11 2 9 14 13 3 1 9 2 7 14 13 1 9 9 7 14 13 9 9 1 10 9 1 9 2
44 9 1 10 9 7 10 9 10 13 0 1 9 2 9 1 9 2 1 9 2 1 9 9 2 9 16 0 2 2 1 10 9 13 1 9 7 1 9 9 13 1 1 9 2
62 13 10 0 1 9 1 9 10 9 7 13 0 15 1 9 1 9 2 7 1 15 14 13 1 9 1 9 7 1 9 9 7 9 2 7 14 0 1 9 1 9 9 7 9 9 0 9 2 14 13 9 1 9 0 0 2 14 9 7 14 9 2
21 13 9 10 9 9 10 11 1 10 9 1 9 2 9 7 9 9 0 10 8 2
18 13 9 2 9 7 9 1 9 14 0 0 1 10 9 7 9 1 2
15 16 14 13 15 1 9 14 9 1 11 1 9 1 9 2
3 9 12 2
9 13 9 1 9 1 9 14 0 2
9 13 1 9 10 9 14 13 15 2
9 1 9 9 1 2 9 10 11 2
15 16 9 1 10 9 14 9 13 0 1 9 14 9 1 2
37 14 13 10 12 9 1 2 7 10 9 14 9 1 10 9 2 15 7 14 9 3 1 9 2 7 13 0 10 9 15 10 9 14 13 9 9 2
34 13 0 9 1 9 3 14 13 9 10 9 9 0 1 1 3 16 13 0 14 9 13 1 11 14 13 15 10 9 9 9 1 15 2
25 13 1 10 9 2 13 10 9 1 14 11 7 10 9 9 16 14 13 9 9 1 9 10 9 2
22 3 9 9 1 9 14 13 3 7 13 9 1 10 9 14 0 1 9 10 9 10 2
32 2 13 12 9 10 1 9 10 9 3 1 11 11 7 11 11 14 13 15 9 15 15 14 9 3 1 9 0 9 3 11 2
13 8 10 9 14 13 15 10 2 2 9 2 1 2
34 13 10 9 0 15 15 1 15 14 9 1 10 9 2 13 1 9 2 1 9 14 13 9 1 15 14 9 3 15 7 15 1 9 2
24 13 9 1 16 13 9 14 13 11 10 11 14 11 3 1 11 1 9 10 9 14 9 3 2
7 13 13 8 14 13 15 2
7 13 9 14 13 15 3 2
14 14 13 15 10 9 10 1 9 1 14 13 0 3 2
7 13 11 12 9 1 9 2
7 9 2 9 9 1 9 2
18 13 15 11 14 14 13 1 10 12 9 2 9 0 2 14 13 15 2
18 13 10 9 0 16 14 13 15 7 14 13 15 1 9 3 1 9 2
22 13 0 9 14 9 1 9 9 1 9 1 9 0 9 9 14 9 1 9 9 11 2
22 13 9 10 9 0 2 9 0 2 1 12 9 14 13 1 9 1 2 9 7 9 2
37 9 14 13 14 0 13 1 11 14 13 9 10 11 9 7 12 1 9 1 9 9 2 7 13 1 10 9 10 13 9 10 11 0 7 1 9 2
15 13 10 9 0 1 9 14 13 10 11 7 9 9 10 2
30 1 9 0 13 8 14 11 9 1 10 9 0 1 10 9 1 9 10 11 7 10 9 13 1 9 0 1 9 9 2
19 16 13 1 9 10 14 9 10 9 9 2 1 10 9 14 9 1 9 2
19 13 15 3 14 13 9 1 9 1 10 9 7 9 10 9 9 1 9 2
42 14 13 10 11 10 9 1 10 9 10 2 7 13 0 14 13 10 11 15 1 9 10 9 9 2 13 9 2 14 13 9 1 9 1 1 10 9 9 15 1 9 2
63 13 15 0 1 10 9 1 9 9 1 9 1 9 9 13 0 3 1 9 14 13 0 1 10 9 7 1 10 9 9 8 10 9 9 2 9 14 13 1 9 1 9 1 10 13 9 2 1 11 7 1 9 10 11 2 2 14 13 10 9 14 11 2
12 13 10 9 0 3 1 9 13 0 1 9 2
8 11 11 3 2 14 9 0 2
4 9 1 9 2
4 9 10 9 2
16 16 13 9 15 10 9 14 13 10 9 0 1 0 1 9 2
8 13 11 14 13 11 14 0 2
12 16 9 10 9 2 13 1 9 14 13 1 2
21 8 14 13 10 9 15 0 15 9 14 13 1 9 7 14 13 15 1 9 9 2
9 2 14 13 10 9 9 14 9 2
9 9 9 15 15 2 9 0 9 2
18 13 1 2 1 9 10 2 13 1 9 10 9 1 9 0 1 9 2
14 13 15 3 14 0 7 10 9 1 9 1 9 1 2
19 2 13 10 9 1 10 9 10 3 1 9 7 1 9 10 11 14 0 2
24 13 15 10 9 15 9 16 14 13 15 1 9 15 2 0 1 10 9 0 10 2 11 11 2
29 14 13 9 11 1 9 10 9 15 0 14 13 10 9 1 1 9 10 11 1 9 9 7 14 13 12 9 1 2
39 14 13 3 1 9 3 16 13 14 13 9 10 9 11 0 1 9 1 10 9 2 7 14 13 1 9 1 3 16 10 9 14 9 1 10 9 14 9 2
39 16 13 10 9 1 14 13 15 15 7 10 11 1 2 13 0 9 10 13 1 9 1 9 0 14 13 9 1 9 1 9 7 1 9 10 11 0 1 2
25 14 0 1 9 10 9 13 9 1 9 14 13 9 14 9 1 9 10 2 7 9 1 9 10 2
30 13 1 10 9 10 9 13 0 3 1 10 11 14 9 7 14 13 10 9 1 9 13 9 0 10 1 9 10 11 2
10 2 13 0 14 13 9 1 9 1 2
10 14 11 14 9 1 9 1 10 9 2
37 13 0 1 10 9 13 1 10 11 1 9 9 1 9 1 9 0 1 9 9 1 15 7 10 9 12 16 14 13 9 1 10 9 1 9 3 2
27 13 11 14 11 7 11 14 11 1 10 12 9 1 9 10 11 10 0 1 3 1 11 11 1 11 11 2
11 14 13 15 9 10 9 1 9 9 3 2
28 13 9 9 11 1 9 9 9 7 9 1 11 3 1 9 14 9 1 10 9 10 1 12 1 12 9 9 2
23 13 1 2 3 2 14 13 9 9 1 9 11 13 0 15 14 9 1 9 0 1 9 2
6 9 9 1 9 9 2
6 2 13 9 1 2 2
18 2 9 0 2 16 9 15 14 13 10 9 1 9 1 9 1 9 2
12 1 9 14 13 10 9 10 9 1 10 9 2
12 9 0 15 15 0 1 9 1 9 14 0 2
6 13 15 1 10 9 2
24 13 15 10 9 14 0 14 13 9 1 10 9 10 14 13 13 9 1 9 10 11 15 10 2
31 13 9 15 9 14 13 10 9 1 10 9 9 0 1 9 16 14 13 15 0 14 13 10 9 1 9 1 9 10 11 2
19 13 10 9 0 10 2 2 13 11 1 9 1 9 1 9 10 9 2 2
19 1 10 9 1 10 9 2 13 15 1 9 3 3 1 10 9 1 9 2
27 13 1 10 9 0 1 9 2 9 0 1 9 9 2 1 9 3 1 10 9 1 10 9 3 2 3 2
7 13 1 9 1 9 3 2
21 13 15 10 9 11 11 1 12 7 13 15 1 9 1 1 9 9 1 9 15 2
14 13 10 9 10 10 9 14 13 9 12 1 9 9 2
36 8 14 13 9 1 9 10 9 10 1 9 10 9 9 14 13 1 9 7 1 9 9 0 16 0 10 9 14 13 10 9 10 1 9 0 2
22 1 12 1 9 1 10 12 9 10 2 13 10 9 1 9 14 0 1 9 10 9 2
15 13 9 0 1 9 16 14 13 9 9 16 13 0 1 2
15 13 15 1 9 1 11 9 1 9 0 1 9 1 12 2
8 13 10 9 14 14 13 15 2
33 14 13 9 9 1 10 9 2 16 13 0 14 13 15 1 2 7 9 1 10 9 13 15 1 9 1 9 10 9 3 1 9 2
9 13 0 10 9 14 9 1 15 2
18 13 10 9 10 9 1 9 14 13 9 3 3 10 9 9 14 9 2
9 13 1 14 9 1 9 9 9 2
18 13 10 9 10 9 11 2 16 14 13 15 16 1 9 1 10 9 2
28 9 9 1 9 15 13 10 9 1 10 9 9 3 1 9 0 14 9 1 9 14 13 0 1 1 10 9 2
10 13 1 10 9 16 14 13 1 9 2
10 13 10 9 14 13 10 9 1 9 2
11 13 15 14 13 10 9 10 9 1 11 2
35 14 13 10 11 1 9 16 3 0 2 7 11 2 7 11 2 7 11 2 7 11 2 9 14 13 0 14 0 1 9 12 9 1 15 2
4 1 9 3 2
8 13 9 1 9 0 10 9 2
5 14 13 10 9 2
14 13 9 9 3 7 13 9 1 9 1 9 10 9 2
5 9 2 5 2 2
