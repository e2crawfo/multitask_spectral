6174 11
9 9 1 12 12 9 13 9 0 0
65 8 8 2 9 0 2 12 2 12 2 8 8 2 2 9 9 13 1 9 0 8 8 7 13 1 15 9 15 1 9 0 7 13 15 1 7 15 13 12 12 9 7 1 7 15 13 0 1 9 9 1 12 9 1 9 9 1 9 9 8 8 1 9 8 2
32 7 13 8 2 12 9 2 9 9 9 0 1 9 8 2 9 9 2 1 7 13 9 9 9 8 0 15 13 9 9 0 2
26 7 13 8 8 0 9 2 14 7 15 13 7 13 9 15 1 9 0 1 9 14 9 7 13 0 2
24 7 1 15 7 9 13 9 13 9 0 7 9 0 7 9 0 7 13 1 15 9 15 0 2
18 7 14 13 1 0 1 15 9 9 9 7 9 9 7 15 13 9 2
25 7 13 1 9 0 13 14 13 2 9 13 15 9 9 2 2 2 2 2 14 15 9 1 9 2
7 14 13 0 1 9 2 2
45 7 1 7 13 9 15 7 9 1 9 7 9 9 15 13 13 1 9 15 1 9 13 1 9 7 13 8 8 0 1 9 12 8 9 8 8 1 7 13 1 15 1 12 9 2
28 7 13 9 1 8 8 8 8 7 15 9 0 1 9 15 13 1 15 8 8 9 9 1 9 1 9 0 2
33 7 13 2 1 9 0 13 9 15 0 1 9 13 9 9 1 9 15 1 9 2 1 9 1 9 15 9 7 9 15 1 9 2
36 7 1 12 9 13 8 8 1 9 9 0 7 9 0 15 13 13 15 0 7 13 1 15 13 9 15 7 13 1 15 9 9 7 9 9 2
30 7 13 13 9 1 9 0 13 1 9 9 8 8 7 13 15 9 9 1 9 9 0 9 9 1 9 9 7 9 2
30 7 13 9 0 1 9 8 8 1 12 12 9 1 15 12 12 9 7 14 13 9 0 1 9 15 1 1 12 9 2
39 7 13 8 8 15 13 1 9 0 1 9 0 1 9 8 8 7 9 8 8 13 9 1 0 14 7 8 13 1 9 0 13 1 9 9 0 1 15 2
29 7 13 2 7 8 8 13 1 9 14 13 0 1 9 15 7 15 13 9 13 9 0 9 1 9 9 15 2 2
26 1 9 13 8 7 15 14 13 1 12 12 9 7 13 1 9 15 9 1 8 1 9 1 9 15 2
31 14 9 7 1 7 13 7 9 0 1 0 7 13 12 12 9 13 9 1 9 8 1 9 8 1 9 1 9 15 3 2
27 7 13 1 15 9 9 9 7 15 13 1 9 2 1 15 7 14 13 7 15 0 1 15 1 9 2 2
14 9 9 0 1 9 1 9 9 0 7 13 9 9 0
60 8 12 2 12 2 8 8 2 2 13 7 9 0 15 13 1 9 9 0 12 1 9 0 9 9 1 9 8 8 1 9 1 8 13 9 9 9 0 7 14 13 0 1 9 0 9 7 13 13 0 9 9 0 0 2 8 8 8 2 2
43 7 9 1 9 1 9 9 9 9 2 13 9 9 9 1 9 0 1 9 9 8 8 15 13 0 1 9 8 8 2 7 15 13 9 1 9 1 9 1 2 9 2 2
41 7 13 2 8 9 1 9 12 1 9 3 9 1 9 9 7 13 13 2 1 1 8 8 2 9 2 2 7 15 9 15 13 15 9 1 9 1 9 9 2 2
10 7 13 7 2 9 9 13 1 8 2
12 7 14 8 1 9 9 9 7 13 9 15 2
7 7 13 1 15 9 2 2
60 7 7 9 8 13 13 2 7 1 1 9 2 13 9 1 9 9 9 9 9 9 0 7 13 9 2 7 13 9 1 9 7 13 9 15 13 1 9 15 1 9 1 9 2 7 13 12 1 15 1 9 7 14 13 0 14 1 9 2 2
28 7 9 1 9 1 15 7 13 3 9 7 14 2 13 9 0 7 2 9 9 13 0 1 9 1 9 9 2
16 7 13 1 0 9 7 13 9 7 14 13 1 9 15 2 2
28 7 13 9 0 13 1 9 1 9 9 9 0 8 8 9 15 7 9 13 9 0 1 9 8 8 9 8 2
25 7 1 9 15 2 13 9 1 9 9 9 0 8 8 9 9 0 0 1 9 8 1 9 9 2
26 7 13 9 8 2 8 1 9 0 0 1 8 7 9 0 9 9 1 9 2 1 10 1 10 9 2
37 7 13 2 8 2 8 2 13 9 3 1 9 1 9 0 9 15 7 15 1 0 9 7 13 9 0 1 9 9 1 8 7 8 8 2 8 2
33 7 13 9 9 13 1 9 8 8 1 9 0 7 15 14 13 9 0 9 1 9 9 1 12 9 2 9 7 1 9 9 0 2
7 9 8 0 2 9 9 8
51 8 2 8 2 12 2 12 2 8 8 8 2 2 13 9 9 8 8 2 8 2 9 15 1 9 9 8 0 2 9 0 1 9 9 1 9 8 8 2 9 0 2 2 15 13 9 9 1 9 8 2
47 7 13 8 2 15 13 1 9 0 1 9 8 9 0 1 9 8 2 13 1 9 1 9 15 13 15 1 9 1 9 2 7 15 14 13 1 8 1 9 9 0 1 15 13 9 8 2
29 7 14 13 9 9 1 8 9 8 8 9 8 1 9 9 9 2 15 14 13 0 9 15 1 9 9 8 8 2
8 9 13 9 0 1 9 1 9
48 9 12 2 12 2 8 8 2 2 13 9 9 8 8 1 9 0 9 15 1 8 9 1 9 1 9 2 7 9 9 1 15 15 13 1 9 1 8 7 9 0 1 9 9 0 1 12 2
39 7 13 9 2 8 2 0 1 9 0 9 9 2 1 12 9 1 9 2 13 9 7 9 9 0 1 9 9 1 9 9 9 0 15 13 1 9 2 2
43 7 1 9 2 7 14 9 9 1 9 13 1 9 9 9 9 0 7 0 13 9 2 7 9 15 15 13 9 0 1 9 2 1 9 1 9 1 9 1 9 9 15 2
15 7 13 9 7 2 12 9 0 0 8 1 9 0 2 2
39 7 14 13 1 9 1 9 0 9 1 9 0 7 9 13 9 7 0 7 9 1 9 9 9 0 9 15 9 1 9 9 0 0 1 8 7 9 0 2
24 7 13 0 1 12 9 9 15 1 9 0 7 9 9 0 7 0 2 13 9 1 9 0 2
6 9 8 2 8 1 9
52 8 2 8 2 12 2 12 2 8 8 8 2 2 13 8 2 9 9 2 9 9 1 9 9 8 1 9 9 1 9 15 1 8 12 2 9 1 9 0 1 9 9 9 0 15 13 1 8 2 8 2 2
43 7 13 9 8 1 9 0 8 8 8 8 1 9 8 8 7 8 8 12 2 12 2 12 2 12 2 7 12 2 12 7 12 2 12 7 12 2 12 7 12 2 12 2
50 7 13 8 13 12 2 8 1 9 0 15 13 1 9 0 7 13 8 8 1 8 12 2 12 7 12 2 12 7 12 2 12 2 8 8 1 8 8 12 2 12 7 12 2 12 7 12 2 12 2
26 7 13 9 9 0 1 0 14 13 9 15 1 9 8 2 7 13 8 1 8 2 7 8 1 8 2
36 7 13 8 1 9 0 1 12 1 12 9 0 2 9 0 1 9 0 7 8 15 13 1 9 9 1 12 1 12 0 1 8 2 8 2 2
22 7 14 13 9 8 8 0 7 15 13 1 12 9 7 12 9 1 9 8 7 8 2
12 9 7 12 9 1 9 9 9 1 9 9 0
44 9 12 2 12 2 8 8 2 2 13 9 0 0 9 7 9 9 9 15 13 9 9 1 9 9 0 15 13 1 9 9 9 14 13 1 9 9 7 9 12 1 9 9 2
37 7 13 9 9 9 7 15 1 9 9 7 9 1 9 8 2 13 8 8 2 12 9 2 1 9 9 1 8 8 2 12 9 2 7 13 15 2
21 7 13 1 9 9 9 8 8 9 9 8 13 1 9 9 1 9 7 13 15 2
35 7 13 7 15 1 1 8 13 9 9 1 9 1 8 8 13 1 9 9 1 15 15 13 1 9 12 1 15 1 15 9 1 9 9 2
15 9 7 9 13 7 13 9 1 8 15 13 1 9 0 2
15 7 13 9 9 15 9 0 12 1 7 15 2 0 2 2
23 7 13 9 0 13 9 9 1 9 12 7 9 12 0 1 15 9 7 9 0 1 9 2
62 1 9 15 13 1 9 8 8 8 9 9 9 9 0 2 9 2 7 9 9 9 0 0 15 13 9 2 7 9 0 1 9 15 0 0 1 9 9 1 9 2 1 10 9 2 0 1 9 15 15 13 15 9 9 0 15 13 15 9 1 12 2
7 9 8 2 8 1 9 9
50 8 2 8 2 12 2 12 2 8 8 8 2 2 13 9 8 8 0 0 9 9 9 1 9 8 0 0 1 9 9 1 9 15 1 9 8 8 8 12 2 12 7 12 2 12 7 12 2 12 2
64 7 13 9 9 15 2 0 8 8 1 9 15 1 9 8 8 12 2 12 7 12 2 12 7 12 2 12 2 7 9 8 8 1 9 15 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 9 8 8 12 2 12 7 12 2 12 2
9 9 8 1 9 1 9 9 9 0
43 9 12 2 12 2 8 8 2 2 13 9 0 0 7 9 9 9 0 1 9 2 8 2 8 8 2 9 9 0 2 13 9 9 9 1 9 1 2 9 9 0 2 2
35 7 13 9 7 8 8 13 1 9 9 9 9 0 1 9 14 13 1 9 9 0 8 8 2 8 1 7 13 15 9 8 8 1 9 2
40 7 13 9 0 1 8 8 8 8 9 1 9 9 7 9 8 2 13 1 9 0 9 1 9 9 9 9 1 8 0 9 15 1 9 2 9 1 8 2 2
19 7 13 8 1 9 1 9 9 1 8 1 9 1 9 9 7 9 9 2
24 7 14 13 1 9 9 7 9 7 9 0 0 7 9 7 14 13 1 9 1 8 7 8 2
39 7 13 8 13 9 9 0 1 9 15 0 8 8 7 13 1 15 2 9 15 1 9 8 2 0 1 9 9 1 8 1 9 9 9 0 1 9 0 2
28 7 1 0 1 9 2 9 13 9 15 13 0 9 1 9 1 9 15 1 9 9 15 12 12 9 1 9 2
35 8 13 7 9 9 9 14 13 1 9 1 8 7 14 13 8 3 9 7 9 14 13 9 0 13 7 13 1 15 9 0 9 1 8 2
46 14 9 15 13 0 0 1 8 7 13 1 9 0 1 9 15 0 7 13 1 9 15 0 9 1 9 2 9 1 7 15 13 12 12 9 1 9 1 15 12 12 9 0 1 9 2
28 7 13 9 7 9 9 9 0 1 9 0 0 2 1 9 9 0 2 8 8 1 9 9 0 1 9 0 2
11 9 9 9 1 9 9 1 9 15 1 9
41 8 12 2 12 2 8 8 2 2 13 9 9 9 1 9 9 0 1 9 9 0 7 13 13 1 9 9 9 1 8 2 9 2 2 1 15 13 9 9 9 2
15 7 14 13 9 7 15 9 0 1 9 2 8 2 8 2
34 12 2 1 9 12 8 8 1 9 9 0 1 9 12 9 1 9 8 0 1 9 9 8 15 13 9 1 15 1 9 1 12 9 2
18 7 13 9 9 8 8 7 9 0 15 13 1 9 15 13 1 8 2
29 7 13 9 14 13 1 9 15 1 9 1 9 1 9 0 1 9 9 2 7 13 1 9 9 9 15 7 13 2
26 13 1 7 9 9 1 9 2 2 12 9 1 9 1 12 9 2 2 13 1 9 9 9 1 9 2
22 7 13 9 9 7 15 13 9 9 9 7 9 9 15 2 7 14 13 13 9 0 2
24 7 14 13 9 9 9 0 1 8 1 9 1 9 8 7 13 1 9 9 1 1 10 9 2
28 7 13 1 9 9 9 12 9 9 7 12 1 9 0 1 9 9 9 1 9 9 1 12 9 1 9 9 2
23 7 14 13 9 1 9 9 1 9 0 1 15 8 7 9 7 9 7 8 7 9 0 2
12 9 8 8 14 13 9 1 1 9 9 1 8
42 9 12 2 12 2 8 8 2 2 13 9 1 9 9 9 0 8 8 1 9 1 9 0 0 9 9 7 9 0 0 0 1 8 8 7 15 8 9 14 13 9 2
49 7 13 9 8 8 2 14 8 8 9 9 15 14 13 15 10 9 1 9 2 7 15 14 13 9 0 9 0 1 15 2 8 8 8 8 7 9 9 13 9 0 1 9 9 9 1 9 2 2
43 7 13 10 9 0 1 9 9 0 1 8 8 7 2 9 13 2 1 9 9 2 9 9 15 1 9 9 8 8 9 9 0 1 9 2 14 7 15 13 1 9 2 2
35 7 1 1 8 2 2 7 13 3 0 9 1 9 9 9 12 7 12 9 0 1 9 14 13 9 1 0 9 1 9 9 8 1 9 2
9 7 0 15 9 1 9 0 2 2
25 7 1 0 7 13 9 0 9 0 1 9 7 14 13 1 9 12 2 9 0 12 7 8 2 2
13 7 13 7 13 1 9 0 1 12 9 2 9 2
48 1 9 0 2 13 9 0 0 7 9 0 14 13 0 2 1 1 15 13 15 9 1 9 0 1 8 8 2 1 9 15 1 9 0 2 1 9 9 7 9 9 0 2 1 9 9 0 2
31 7 13 9 7 15 7 1 9 10 9 2 14 13 9 8 1 9 2 9 2 1 9 9 1 9 9 9 1 9 15 2
37 7 14 13 9 0 7 0 7 0 1 9 9 1 9 0 7 1 9 0 1 9 9 1 9 1 9 15 13 13 1 9 2 1 1 9 0 2
47 7 13 9 8 8 1 9 0 1 9 9 9 0 13 15 9 0 9 1 9 0 2 8 8 7 13 9 0 8 8 1 9 1 9 1 9 13 10 9 0 2 1 9 0 1 9 2
39 7 13 9 0 0 1 9 0 9 15 7 9 9 0 7 0 13 2 1 9 0 2 9 1 9 1 9 0 1 9 9 0 7 9 9 9 0 0 2
9 9 13 9 1 9 1 9 8 8
43 9 12 2 12 2 8 8 2 2 13 9 2 9 2 0 9 9 9 1 9 9 15 1 9 0 0 1 8 8 7 15 13 2 1 1 9 1 2 9 2 9 0 2
47 7 13 9 7 2 9 0 0 1 9 9 15 7 9 9 1 9 2 9 7 2 1 9 0 9 1 9 9 7 9 12 7 12 9 1 10 9 13 7 13 1 9 9 7 9 2 2
35 7 13 2 13 1 9 15 13 15 7 15 9 9 7 9 7 7 1 9 7 13 9 9 0 7 9 0 7 13 1 9 9 9 2 2
46 7 13 9 9 0 8 8 13 1 9 9 1 8 8 1 9 0 8 8 2 12 9 0 2 13 9 9 0 9 1 9 0 1 9 9 0 0 7 1 15 9 7 9 9 0 2
17 7 13 9 2 10 9 13 0 9 0 7 13 9 9 0 2 2
35 7 13 1 7 2 9 0 15 13 8 1 9 15 14 13 1 9 7 9 7 9 7 14 13 1 15 1 9 1 9 9 1 9 2 2
14 12 9 1 9 1 15 12 9 1 9 9 2 9 2
39 9 12 2 12 2 8 8 2 2 13 9 0 9 9 7 12 9 1 15 12 1 9 9 9 13 7 13 12 0 1 9 7 9 1 9 9 1 9 2
42 7 13 9 2 8 2 7 12 9 13 7 13 12 0 9 9 9 1 9 13 15 9 0 0 1 9 15 1 8 1 9 8 8 2 12 8 1 9 9 0 2 2
34 7 13 9 9 7 9 1 9 13 7 13 0 1 9 9 1 9 13 15 9 0 0 1 8 1 8 2 12 8 1 9 9 2 2
28 7 13 9 8 7 15 13 9 1 9 9 13 1 9 1 12 9 2 9 1 9 1 8 1 8 9 0 2
25 7 13 9 7 9 13 1 9 1 9 7 8 8 8 7 13 0 1 9 9 1 9 9 0 2
23 7 13 9 9 1 7 9 0 1 8 13 9 1 9 9 0 1 7 13 9 1 9 2
32 7 13 9 3 7 12 9 13 1 9 3 9 1 9 9 13 1 9 9 1 9 8 1 9 2 12 8 1 9 9 2 2
35 1 15 13 12 0 0 9 1 9 1 9 9 1 9 2 12 8 1 9 9 2 7 1 9 2 12 8 1 9 9 2 1 1 9 2
37 7 13 9 1 9 9 2 9 9 0 1 9 9 13 12 9 1 0 1 15 1 12 0 0 2 7 1 12 9 1 1 9 13 9 1 9 2
12 7 14 13 9 7 7 15 14 13 10 9 2
9 9 9 0 2 9 0 13 9 15
39 9 12 2 12 2 8 8 8 2 2 13 9 9 0 9 15 1 9 1 9 9 0 0 1 9 9 15 13 15 9 1 12 1 12 9 2 9 0 2
68 7 13 1 10 9 0 7 0 9 9 9 9 7 9 9 0 1 9 9 2 7 13 9 9 9 9 0 15 13 1 9 7 13 9 0 0 2 7 13 9 0 1 9 9 9 0 15 13 1 9 7 13 9 8 3 2 7 14 13 8 0 0 9 9 9 1 15 2
52 7 13 9 1 9 1 1 9 1 9 8 2 9 9 2 15 13 15 9 1 15 1 9 9 15 1 9 9 0 9 2 7 13 9 0 1 9 0 2 9 9 9 0 2 7 13 1 15 12 2 12 2
34 7 13 9 1 9 9 0 1 7 13 1 15 9 15 0 0 8 8 0 2 9 1 7 15 14 13 1 15 1 9 9 1 9 2
19 7 13 8 15 13 13 1 9 0 1 9 0 7 13 9 1 9 0 2
72 7 13 9 9 13 1 9 0 9 9 1 9 0 1 9 9 9 1 9 9 2 7 13 0 8 8 1 12 12 9 7 9 8 8 1 9 9 0 7 9 8 7 15 13 9 1 9 9 0 9 8 8 7 9 8 8 8 8 8 8 1 7 13 9 1 15 1 9 9 9 15 2
56 7 13 9 9 3 1 9 9 9 15 13 9 0 1 9 0 1 9 9 0 9 9 1 9 15 13 15 1 9 0 7 1 15 11 8 8 13 8 9 1 9 15 7 11 8 8 8 8 8 8 13 9 9 9 8 2
17 7 13 10 9 9 9 0 9 1 9 9 8 8 8 8 8 2
43 7 13 9 9 9 1 9 9 1 12 9 2 1 12 12 9 2 7 9 1 9 12 9 2 1 12 12 9 2 7 13 9 9 9 12 12 9 2 12 12 9 2 2
58 7 13 9 8 9 13 1 9 9 9 0 8 8 1 8 9 2 9 9 2 1 1 9 1 12 12 9 2 12 2 12 8 2 2 7 15 0 9 1 9 9 0 1 9 7 15 13 1 15 9 0 1 9 9 0 9 0 2
20 7 13 1 9 7 13 1 9 0 1 0 8 8 8 8 8 8 8 8 2
72 7 1 9 0 1 9 0 2 7 14 9 14 13 13 9 1 9 0 7 0 8 1 9 15 13 1 15 9 15 7 1 9 15 0 0 9 1 9 8 8 9 2 0 2 7 13 15 9 0 7 9 15 0 1 8 9 8 1 9 0 1 9 8 12 1 9 0 13 0 1 9 2
39 7 1 9 9 9 2 13 9 9 1 9 9 1 9 9 9 1 9 9 0 0 12 1 9 7 13 9 9 1 9 12 12 9 2 1 12 9 2 2
112 13 7 9 15 0 9 13 9 15 1 9 9 9 9 0 7 13 9 9 0 15 13 1 9 9 12 2 7 9 15 0 1 9 7 13 1 9 12 9 2 7 13 1 9 0 12 9 9 12 7 12 7 12 2 7 9 9 2 9 9 9 0 2 9 9 12 7 12 2 7 9 9 9 0 12 9 9 12 7 12 7 12 2 7 9 9 9 0 9 9 12 7 12 2 7 9 9 0 9 9 12 7 12 2 7 9 9 0 0 9 12 2
12 9 8 2 9 8 13 9 0 0 1 9 0
44 9 12 2 12 2 8 8 8 2 2 13 9 8 8 8 9 0 0 1 9 9 0 1 9 15 12 2 12 8 1 9 0 0 1 9 8 1 9 9 15 13 15 9 2
27 7 13 9 0 7 15 12 2 12 8 1 9 8 1 9 7 13 15 1 12 9 2 9 0 1 8 2
27 7 13 8 9 8 8 0 2 12 2 12 8 2 7 8 8 1 8 0 2 12 2 12 8 3 2 2
75 7 13 9 9 0 1 9 12 9 2 12 0 7 12 0 7 12 0 2 2 13 15 9 1 9 12 9 2 12 0 7 12 0 7 12 0 2 2 7 9 1 0 12 9 2 12 0 7 12 0 7 12 0 2 2 1 1 13 9 0 1 9 12 9 2 12 0 7 12 0 7 12 0 2 2
15 9 9 9 1 9 13 1 2 9 0 2 1 9 9 9
36 9 12 2 12 2 8 8 2 2 13 9 9 9 0 8 8 9 9 2 9 0 2 15 13 15 9 0 1 9 9 9 9 9 1 9 2
40 7 13 8 1 9 0 2 3 9 13 2 14 13 1 9 15 9 9 1 9 1 10 9 1 9 1 9 9 13 1 9 12 9 1 1 9 9 9 2 2
22 7 13 1 7 9 9 13 1 9 1 9 7 13 1 2 9 13 1 9 0 2 2
17 13 1 7 9 9 0 15 13 9 9 0 13 1 9 9 9 2
30 7 13 9 9 9 7 2 9 0 0 1 12 9 1 9 9 13 9 9 1 9 0 2 1 1 9 9 1 9 2
24 7 13 9 1 9 13 1 9 9 0 1 9 1 9 9 1 9 9 9 13 1 9 0 2
25 7 13 10 9 9 0 1 9 0 1 9 2 9 12 13 0 1 12 9 1 9 0 7 0 2
39 7 13 9 9 9 0 15 13 15 9 7 13 15 9 12 9 1 9 9 0 1 9 0 1 9 9 9 0 0 0 1 9 1 8 8 1 9 0 2
6 8 13 1 9 9 15
40 8 12 2 12 2 8 8 2 2 13 9 9 0 1 9 8 8 8 15 13 1 15 1 12 9 2 9 1 9 0 2 9 9 1 9 9 15 1 9 2
42 7 13 8 15 13 1 15 9 1 9 0 13 15 1 9 9 1 12 9 9 9 9 9 9 8 8 2 1 9 7 9 9 15 9 0 1 2 9 9 0 2 2
43 7 13 7 2 0 9 0 1 9 14 13 15 9 8 8 8 9 1 9 0 1 0 9 2 2 8 1 9 1 8 8 1 7 9 13 9 2 8 8 9 0 2 2
22 7 13 9 15 13 9 0 1 9 0 13 9 9 1 9 0 1 9 9 1 8 2
17 7 13 9 9 7 0 15 1 9 1 7 13 9 15 1 9 2
23 7 14 13 9 0 10 9 1 9 9 1 9 8 9 1 9 15 13 1 9 8 8 2
38 13 1 7 9 9 13 1 9 0 7 7 9 9 13 1 9 0 1 9 15 0 9 15 13 12 5 1 9 0 7 13 1 9 0 1 9 9 2
14 8 8 13 0 9 1 9 0 13 9 1 9 8 2
26 7 1 0 7 13 9 0 0 8 8 8 0 1 8 8 9 9 9 0 1 9 9 1 9 9 2
11 9 9 9 0 2 9 0 1 8 7 8
64 8 2 9 0 2 12 2 12 2 8 8 8 2 2 13 9 0 8 8 8 8 9 0 1 9 9 9 9 0 1 8 8 2 8 8 8 1 9 0 1 9 9 9 12 8 1 9 7 9 1 7 13 12 2 12 8 7 12 2 12 8 1 9 2
16 7 13 8 9 0 7 13 0 0 9 1 15 1 9 0 2
52 7 13 8 2 9 14 8 8 2 8 9 9 1 0 1 12 9 1 9 9 8 1 15 0 2 2 0 2 8 8 0 1 9 9 9 2 8 8 8 13 7 15 8 8 8 9 12 2 12 9 2 2
30 7 13 8 2 8 1 9 9 0 2 9 1 15 13 1 9 15 1 9 9 15 0 1 9 15 12 9 10 9 2
22 7 13 8 8 2 9 9 12 15 13 8 10 9 2 0 1 9 12 2 12 8 2
16 1 9 15 2 13 8 9 0 9 0 0 9 1 9 0 2
11 9 8 12 2 8 2 9 9 9 13 9
48 8 12 2 12 2 8 8 8 2 2 13 9 9 9 0 1 9 9 9 1 9 9 8 2 8 0 8 8 8 8 2 0 1 9 9 12 1 9 9 0 9 15 1 9 7 8 0 2
48 7 13 1 9 9 9 12 9 13 1 12 9 2 13 8 8 7 8 7 8 7 8 7 8 2 7 0 8 8 8 8 8 7 8 8 8 2 7 0 8 7 8 7 8 7 9 0 2
17 7 13 9 1 9 9 7 9 7 13 9 9 9 0 1 9 2
6 9 9 0 1 9 8
48 8 2 8 2 12 2 12 2 8 8 2 2 13 9 9 9 1 8 1 9 9 0 1 9 9 0 0 8 2 8 8 13 9 0 1 12 9 1 9 15 7 13 9 15 12 9 0 2
21 7 13 8 9 9 9 8 8 13 1 12 9 2 9 1 9 12 1 9 15 2
20 7 13 9 9 9 0 1 9 12 7 12 7 13 9 12 9 7 9 9 2
33 7 13 9 0 9 8 1 15 9 8 1 9 0 1 9 1 9 9 9 1 9 9 7 13 9 9 15 1 9 15 9 12 2
12 9 0 1 8 13 9 1 9 15 2 9 2
39 8 2 8 2 12 2 12 2 8 8 2 2 13 9 9 9 8 1 9 15 9 0 1 9 15 15 13 9 9 0 1 9 0 1 9 10 9 0 2
29 7 13 2 9 0 2 0 9 15 13 1 9 1 9 9 1 9 10 9 0 0 1 9 0 1 9 8 8 2
24 7 13 9 9 0 8 8 1 9 8 8 2 7 9 8 15 9 0 1 9 9 0 2 2
34 14 7 10 9 13 7 13 1 7 9 13 7 13 2 0 9 2 7 2 9 9 0 2 1 9 14 13 9 1 15 1 9 0 2
18 7 13 8 2 14 9 1 9 1 9 0 1 9 1 9 8 8 2
32 7 9 0 7 13 7 13 1 9 14 13 9 8 8 2 9 13 0 1 9 2 0 1 9 9 1 9 9 1 8 2 2
26 7 13 9 8 13 1 9 0 1 9 0 1 8 7 8 8 2 9 9 2 1 7 13 1 15 2
31 7 13 10 9 1 9 2 9 0 1 9 9 0 0 7 13 8 1 9 9 7 13 9 9 8 8 1 9 8 8 2
30 7 13 9 9 8 8 2 12 12 9 2 0 1 9 1 9 9 8 1 9 9 9 1 9 1 8 9 1 9 2
56 7 13 8 8 2 7 8 1 9 9 14 13 0 1 9 7 3 9 0 1 9 15 13 10 9 1 9 9 15 13 15 1 8 2 9 2 0 2 7 9 2 9 0 15 9 2 7 9 0 1 9 7 9 0 2 2
23 7 13 2 8 0 8 9 0 2 0 1 15 2 7 15 14 13 3 9 1 9 2 2
54 7 1 9 1 9 9 9 7 1 9 0 1 9 13 1 9 13 9 7 9 8 8 2 12 9 2 2 8 9 0 7 0 8 8 3 1 9 0 7 1 9 13 9 8 8 8 1 8 8 9 9 8 2 2
27 7 13 9 0 0 0 9 9 9 8 8 1 8 15 3 1 9 9 1 9 0 0 0 1 9 8 2
31 7 13 9 9 9 0 0 8 8 7 9 14 13 7 2 13 1 9 2 7 9 9 13 15 1 15 13 1 9 0 2
34 7 13 8 8 9 1 9 8 10 9 7 13 7 12 1 12 1 9 1 8 13 9 1 9 0 1 8 1 12 1 12 13 9 2
39 7 13 9 9 7 1 9 8 0 7 13 9 1 9 15 1 9 9 1 9 15 15 14 13 1 9 8 7 13 1 2 9 2 9 1 8 8 8 2
17 7 13 9 1 9 7 9 9 15 13 1 9 9 9 1 9 2
29 7 13 9 1 8 1 9 0 1 9 12 12 9 14 7 15 13 1 9 9 9 0 1 9 7 13 1 9 2
24 14 7 9 9 8 8 13 7 9 0 2 8 8 1 9 15 1 9 2 14 13 9 0 2
13 7 15 9 13 15 3 9 9 9 1 9 0 2
14 9 8 0 1 9 15 0 13 1 9 9 2 9 2
47 8 2 8 2 8 2 12 2 12 2 8 8 2 2 13 9 1 9 8 0 1 9 9 0 1 10 9 0 0 1 9 9 7 8 1 9 9 7 1 0 9 9 0 0 1 15 2
21 7 1 9 15 0 14 13 1 9 8 0 15 13 1 9 0 1 12 12 9 2
33 7 15 13 1 9 0 0 1 9 9 0 1 9 9 7 13 9 15 1 9 12 0 1 9 14 12 15 13 1 15 8 0 2
56 7 13 8 8 9 1 9 0 1 9 9 1 8 1 9 8 8 2 9 12 13 15 1 12 12 9 9 15 1 9 15 13 1 9 0 2 8 8 2 7 1 12 9 3 14 7 15 13 1 7 13 10 9 0 2 2
67 7 13 1 8 7 13 2 9 9 2 1 0 9 0 0 2 12 9 1 15 9 8 0 2 7 9 9 13 9 0 1 9 8 2 7 9 0 0 13 1 12 9 1 9 8 2 7 9 0 13 9 0 1 9 2 9 1 9 8 1 9 15 0 1 9 0 2
22 7 1 9 9 0 1 9 9 1 10 9 0 15 14 13 9 9 15 14 9 9 2
41 7 1 9 9 9 9 7 9 9 1 0 9 15 7 9 2 14 7 13 0 1 9 9 7 9 7 14 13 9 15 1 9 8 9 0 1 9 1 9 8 2
36 7 13 9 10 9 9 7 1 9 9 9 1 15 13 1 15 1 9 0 7 0 1 9 2 14 9 0 7 14 13 1 9 1 9 0 2
36 7 13 9 8 2 15 13 1 0 0 2 9 9 1 9 8 15 8 1 15 1 9 15 1 9 7 9 7 9 7 9 2 2 2 8 2
11 14 9 15 7 15 9 13 1 9 0 2
13 7 13 10 9 0 9 1 9 1 9 9 0 2
24 7 13 9 9 0 9 1 9 8 7 13 9 1 12 9 0 1 9 0 1 9 9 8 2
14 7 13 9 9 9 0 1 9 9 1 9 9 9 2
28 7 13 9 1 9 9 0 1 9 9 9 8 8 7 13 1 9 15 7 13 15 9 9 1 9 15 0 2
15 7 13 9 1 9 7 9 0 12 8 7 12 9 0 2
26 7 13 8 9 9 2 7 9 9 13 0 1 9 9 7 9 7 9 15 13 9 15 1 9 2 2
26 7 13 9 1 9 1 9 1 9 9 7 13 1 15 9 0 13 9 9 9 1 15 1 12 9 2
24 1 9 13 9 1 15 13 8 8 9 1 15 9 1 9 9 1 9 0 9 0 1 9 2
26 14 7 9 9 9 14 13 7 13 9 0 14 1 9 9 9 15 13 1 9 9 1 10 9 0 2
34 7 9 1 9 1 8 13 12 9 7 9 9 13 1 15 9 7 9 9 1 9 1 9 8 2 8 7 9 10 9 13 1 9 2
17 7 14 13 1 10 9 1 9 0 7 14 13 15 9 9 9 2
10 8 13 8 8 1 9 15 9 1 8
49 8 12 2 12 2 8 8 2 2 13 9 0 8 8 9 9 9 1 9 0 8 8 1 9 9 15 9 1 9 13 1 15 1 15 7 2 13 9 9 1 9 9 8 1 9 7 9 2 2
70 7 13 1 9 9 15 13 15 9 9 0 8 7 9 8 9 15 2 9 7 9 1 9 1 9 2 9 0 8 8 0 2 8 1 9 0 1 7 15 14 13 9 1 10 9 7 14 13 0 9 1 0 9 2 1 9 10 13 1 15 9 15 1 9 7 9 7 9 2 2
61 7 13 8 2 8 0 9 0 0 15 13 15 1 8 0 1 9 9 8 8 8 8 1 9 15 1 9 7 9 9 15 0 9 0 1 9 2 7 1 9 15 9 15 1 9 7 9 9 2 7 9 9 15 0 7 9 15 9 0 2 2
65 7 13 8 1 2 9 1 9 9 9 2 7 9 9 8 9 7 9 9 1 9 0 2 7 13 0 9 7 9 1 9 9 0 2 0 1 9 1 9 8 8 8 1 8 8 1 9 9 9 8 8 1 9 15 0 2 7 13 0 0 1 9 15 2 2
41 7 13 8 8 1 12 1 12 1 9 1 9 0 15 13 9 0 7 13 1 15 9 1 9 15 15 13 1 0 1 9 2 9 1 7 13 8 1 12 9 2
10 9 9 1 9 0 1 8 8 1 9
41 9 12 2 12 2 8 8 2 2 13 9 8 8 9 9 7 8 13 9 1 9 0 9 1 9 8 8 15 13 1 9 0 1 9 13 1 9 1 9 0 2
51 7 14 13 9 1 9 9 13 15 9 8 7 13 1 15 12 9 0 9 13 1 15 9 9 7 9 1 9 0 1 9 9 8 8 2 7 13 0 1 9 9 0 7 9 9 0 1 9 0 0 2
59 7 13 1 10 9 9 13 2 7 9 8 14 13 1 10 9 1 9 15 9 1 9 9 7 9 0 15 13 8 8 7 13 1 9 0 8 8 8 8 8 8 8 1 9 8 8 8 0 8 8 8 8 13 9 9 8 0 2 2
65 7 13 9 2 7 9 9 7 9 15 9 13 0 15 7 13 1 9 1 9 9 0 9 15 0 7 0 1 9 1 0 9 1 9 9 7 9 0 1 9 9 1 9 15 7 15 13 9 7 9 1 9 15 9 15 1 9 9 9 7 15 13 9 2 2
47 7 13 9 8 2 9 0 0 7 9 2 0 8 2 8 1 9 9 15 1 9 0 1 10 9 0 7 9 1 9 9 0 9 9 1 9 9 9 7 15 13 1 15 1 9 2 2
22 7 13 9 0 1 9 8 1 9 9 9 1 9 12 9 1 9 1 9 9 9 2
41 7 13 9 9 0 13 1 15 2 9 9 0 2 7 13 9 9 1 8 8 1 9 1 9 9 12 0 1 9 0 1 9 0 7 15 13 9 9 7 9 2
8 1 9 1 9 1 9 8 8
10 8 12 2 12 2 12 2 6 8 2
52 1 0 9 8 8 1 9 9 0 7 8 9 0 0 1 0 9 1 2 9 0 2 7 2 9 0 2 7 2 1 14 9 2 7 2 9 0 2 7 9 15 1 10 9 1 1 7 8 8 1 9 2
41 13 8 8 1 9 7 8 9 1 9 9 2 1 9 15 0 2 1 9 15 2 8 14 8 7 8 9 0 1 10 9 1 9 9 0 8 8 1 9 9 2
13 1 9 0 7 8 8 0 15 9 7 13 9 2
17 7 15 13 1 9 0 1 9 0 14 13 1 9 9 1 9 2
58 7 13 10 9 13 9 9 1 9 15 0 2 7 15 15 13 1 15 1 13 2 1 9 9 9 1 9 9 7 9 1 12 7 12 9 13 15 1 9 15 1 9 2 7 9 9 1 9 0 7 12 7 13 9 15 1 9 2
37 7 1 15 14 13 9 1 8 8 9 15 7 13 9 0 2 7 9 8 8 13 9 15 1 10 9 1 9 9 7 13 1 9 9 9 0 2
11 9 9 0 2 8 8 14 13 9 9 15
41 9 12 2 12 2 8 8 8 2 2 13 9 0 1 9 9 0 8 8 9 9 8 7 9 0 8 8 14 13 1 9 0 9 9 15 13 15 9 9 12 2
34 7 13 8 1 9 2 9 2 0 7 15 14 9 1 2 9 2 1 9 8 1 9 1 9 15 9 9 9 15 1 9 9 9 2
21 7 13 2 9 8 14 13 7 13 1 9 13 1 15 9 15 1 9 15 2 2
35 7 13 9 15 9 1 9 1 9 7 13 9 9 0 0 8 8 1 9 9 8 8 1 9 9 9 8 1 9 0 7 1 9 0 2
41 7 13 9 1 9 1 9 0 0 1 9 8 1 9 9 15 1 9 9 15 1 1 13 8 1 9 0 1 9 0 1 9 1 9 0 1 9 2 9 12 2
25 7 13 9 0 1 7 8 0 1 9 9 9 1 9 0 2 7 13 9 0 8 8 0 2 2
22 7 13 7 9 0 0 1 8 8 14 13 9 1 9 0 1 9 9 0 8 8 2
65 7 13 2 8 8 15 13 1 9 8 8 0 1 9 8 8 8 15 14 13 1 15 8 1 9 12 15 13 1 15 2 1 9 1 2 9 0 2 15 13 15 8 8 1 9 1 9 0 8 8 15 13 9 9 0 9 1 9 9 7 9 1 9 0 2
67 7 9 1 9 1 9 2 9 9 0 9 0 1 9 1 9 12 1 9 9 2 1 9 10 13 1 15 9 8 0 15 13 9 0 1 9 1 9 9 1 12 9 1 9 2 13 8 2 10 1 9 7 9 9 1 9 9 1 1 8 8 15 8 1 15 2 2
22 9 7 15 13 2 10 9 1 9 13 0 7 14 9 1 9 1 9 7 9 2 2
38 7 1 0 7 13 8 8 15 13 9 0 12 1 9 0 1 9 12 1 12 1 9 2 9 0 1 9 9 1 9 7 13 9 0 1 9 15 2
12 9 13 9 9 1 9 9 1 9 0 9 0
39 9 12 2 12 2 8 8 2 2 13 9 0 0 9 9 9 1 9 0 9 1 12 9 2 9 1 9 1 7 15 14 13 9 0 1 9 9 0 2
41 7 1 9 13 15 9 9 0 9 9 13 7 9 2 13 1 9 9 1 9 9 9 15 1 9 15 13 1 12 9 2 9 7 9 1 9 0 1 15 2 2
82 7 13 9 7 15 2 13 9 1 9 9 0 1 9 9 9 9 2 9 7 9 7 9 7 9 1 9 9 0 1 15 7 9 15 1 9 7 9 0 1 9 15 7 9 1 9 9 1 9 7 9 0 1 15 1 9 9 1 9 7 9 0 9 9 7 9 9 9 9 7 9 0 9 2 9 1 0 1 9 2 9 2
26 7 13 10 9 1 9 9 13 1 9 2 9 1 9 9 15 14 13 1 9 0 0 1 9 9 2
27 7 13 13 9 13 9 15 1 12 9 2 9 7 13 1 9 1 10 9 1 9 9 1 1 0 9 2
24 7 9 9 1 10 9 2 13 9 0 1 12 12 9 0 1 9 9 0 1 9 2 9 2
33 7 13 9 2 9 2 13 9 7 9 0 13 12 12 9 13 1 12 9 2 1 15 12 9 2 13 9 0 1 9 9 0 2
34 7 13 9 1 12 9 1 9 15 14 13 1 9 0 0 13 1 9 0 1 12 12 9 9 15 1 9 7 9 1 1 9 0 2
16 8 2 9 9 0 1 9 2 14 13 1 9 1 9 9 2
43 9 12 2 12 2 8 8 2 2 13 9 9 0 11 8 8 1 9 0 13 9 9 7 9 9 0 1 9 1 10 13 12 9 2 14 13 1 9 1 9 9 2 2
45 7 13 8 1 9 1 9 2 9 2 15 13 8 8 1 9 1 15 7 2 9 1 15 9 0 1 7 9 9 14 13 1 9 1 9 9 15 13 8 0 1 10 9 2 2
12 7 13 8 7 2 9 14 13 1 9 9 2
17 8 8 8 8 9 1 9 7 1 9 0 1 9 9 0 2 2
38 7 13 9 9 0 1 9 9 14 12 1 9 9 8 0 1 9 2 7 9 0 1 9 13 1 9 7 1 9 9 9 7 9 9 9 0 2 2
57 7 13 13 2 1 9 13 10 9 0 1 7 9 9 1 9 14 13 0 9 1 9 9 9 7 14 3 12 1 12 2 2 0 1 2 9 9 0 1 0 1 9 7 9 9 9 0 7 9 9 9 1 9 9 0 2 2
10 9 13 1 9 0 0 1 9 8 12
40 9 12 2 12 2 8 8 2 2 13 9 0 7 15 13 2 1 9 2 9 9 9 0 1 9 9 2 9 2 8 12 2 15 13 8 8 1 12 9 2
32 7 13 9 1 9 9 0 1 9 9 7 2 9 0 5 8 12 5 13 1 9 0 1 9 1 9 15 1 9 0 2 2
27 7 13 13 1 9 2 9 12 1 9 0 9 1 10 9 15 13 7 13 9 9 9 7 1 15 9 2
35 7 13 10 9 0 9 9 9 15 7 9 0 2 13 1 9 9 9 0 0 7 14 13 1 0 9 1 9 0 9 1 9 0 2 2
24 7 13 2 7 9 15 9 9 0 1 9 1 9 8 9 2 7 15 14 13 9 9 9 2
13 7 14 13 9 9 0 9 9 0 7 9 9 2
34 7 13 9 0 13 1 9 2 9 12 7 9 14 13 1 9 9 2 8 2 12 2 7 15 9 0 1 9 2 8 2 12 2 2
17 7 13 9 9 8 8 7 9 1 9 0 14 13 9 9 0 2
48 7 13 9 0 0 13 7 15 14 13 1 9 0 9 9 2 9 13 1 15 9 2 9 2 7 15 9 0 1 9 0 0 1 9 2 8 2 8 2 7 2 8 2 8 2 0 9 2
14 7 13 9 0 7 15 13 9 9 0 1 9 9 2
3 1 9 9
72 8 12 2 12 2 8 8 2 2 1 15 13 9 9 0 0 1 9 9 2 9 2 9 9 13 9 0 7 9 15 13 1 9 9 1 9 13 7 13 9 9 0 2 7 9 9 1 15 15 13 1 9 1 8 7 9 0 7 13 9 0 14 13 1 15 1 9 13 1 9 9 2
39 1 9 12 8 8 8 2 9 8 13 9 9 0 8 8 1 8 9 0 9 0 1 9 0 0 0 15 13 8 9 0 2 1 9 9 9 0 2 2
8 9 9 0 13 1 9 1 9
42 8 12 2 12 2 8 8 2 2 13 9 0 7 9 0 8 8 11 8 13 9 9 9 9 8 11 8 1 9 1 9 0 8 8 8 1 9 9 1 9 0 2
38 7 13 9 9 15 7 9 0 0 13 2 9 0 2 1 9 9 0 13 2 1 9 9 9 1 9 9 1 9 9 0 7 0 9 9 0 2 2
57 7 13 9 11 8 1 12 9 1 9 15 13 1 15 9 9 0 9 15 8 8 15 13 9 9 0 9 0 1 9 8 8 1 2 9 0 2 7 14 3 9 9 0 2 15 13 9 7 8 7 9 7 8 7 8 2 2
44 7 13 10 9 0 15 8 9 12 9 1 12 1 9 9 0 0 1 9 7 9 1 12 1 9 0 15 13 15 9 9 12 7 13 1 9 15 9 8 0 1 9 9 2
42 7 13 8 1 9 9 9 8 1 9 2 9 7 9 2 9 7 13 8 0 9 0 8 8 7 9 0 8 15 13 1 9 15 1 9 9 0 1 9 9 15 2
35 7 13 9 0 1 9 0 8 8 9 9 7 9 8 1 9 9 0 1 9 0 8 8 1 9 0 1 9 9 0 1 9 9 9 2
10 9 8 9 1 9 8 1 9 9 9
48 8 12 2 12 2 8 8 2 2 13 9 0 9 9 7 9 9 1 8 2 0 2 8 9 15 13 15 9 10 9 1 9 9 9 0 0 8 8 1 9 13 1 15 1 9 1 9 2
28 7 14 13 9 8 8 2 12 9 2 1 9 0 2 9 2 1 9 9 9 2 1 9 9 13 12 9 2
24 7 13 8 7 9 9 2 13 9 9 0 8 8 8 7 1 3 9 1 8 9 9 2 2
47 7 13 9 15 13 9 15 8 8 8 8 8 7 8 13 9 9 1 9 15 1 9 2 7 9 0 7 0 1 9 15 13 15 2 9 2 13 14 13 1 9 1 8 9 0 2 2
50 7 13 9 13 1 9 2 9 12 1 9 12 9 1 8 7 9 15 1 9 0 9 0 1 9 15 1 9 9 1 2 9 8 2 2 8 2 1 0 7 13 9 15 0 0 0 1 9 0 2
34 7 13 1 12 1 9 9 2 0 2 9 9 0 0 7 9 9 9 1 7 15 13 2 9 2 1 9 1 9 15 9 9 0 2
26 7 13 9 9 8 8 8 1 9 9 1 8 0 14 15 1 7 15 2 9 0 2 1 9 9 2
15 9 13 7 15 1 0 1 9 15 9 9 0 1 9 8
48 9 12 2 12 2 8 8 2 2 13 9 7 9 9 0 8 8 2 8 13 9 9 7 9 0 1 9 9 0 1 9 2 8 2 14 13 0 1 9 15 9 1 9 0 1 9 0 2
28 7 13 9 9 9 0 1 9 1 9 0 1 9 8 9 8 8 8 13 9 9 9 1 9 0 1 9 2
29 7 13 9 0 1 9 2 8 8 7 9 8 14 13 0 1 9 15 8 8 13 7 8 8 8 9 9 2 2
46 7 13 8 2 8 2 7 9 0 1 9 0 13 9 1 9 9 2 0 1 2 7 15 13 1 0 9 8 9 1 9 9 2 1 1 7 13 9 9 9 1 9 0 1 9 2
41 7 14 13 9 0 8 8 1 9 0 1 9 9 9 9 9 9 9 1 9 2 8 2 1 2 9 3 1 9 9 1 9 0 1 9 9 7 9 15 2 2
54 7 13 8 1 9 1 9 0 1 9 9 9 1 9 2 8 2 7 9 9 0 8 8 2 13 7 3 9 13 1 9 9 1 9 7 9 7 9 1 9 9 9 7 13 9 14 13 9 15 1 9 0 2 2
20 7 13 8 8 9 1 9 1 9 9 9 8 0 1 9 2 9 1 8 2
45 7 13 8 1 9 1 9 9 1 8 1 9 1 9 9 7 9 9 13 1 9 15 9 7 9 7 9 0 0 7 9 1 7 13 1 8 7 8 1 9 9 15 1 9 2
34 7 1 0 1 9 2 9 13 9 2 0 9 1 9 1 9 2 7 15 0 1 9 9 15 1 9 1 9 12 12 9 1 9 2
14 9 7 15 14 13 9 1 9 8 1 9 9 9 2
23 7 13 8 13 3 9 7 9 0 14 13 9 0 9 1 8 7 13 7 13 9 0 2
40 7 13 9 2 0 0 9 1 9 1 8 7 13 9 15 12 12 9 1 9 1 15 12 12 9 0 1 9 2 0 9 1 9 1 9 15 1 9 9 2
31 7 13 9 7 9 9 9 0 1 9 0 9 15 2 9 9 0 2 7 9 9 1 9 9 0 15 13 9 1 9 2
15 9 8 7 9 9 9 1 12 9 1 8 1 9 9 9
41 8 12 2 12 2 8 8 2 2 13 9 9 0 9 9 7 0 13 9 15 7 7 9 9 13 1 12 9 9 1 9 9 0 1 9 0 9 9 7 9 2
34 7 13 8 8 9 1 9 7 9 13 15 9 0 1 8 2 9 2 13 8 1 14 12 2 15 9 0 1 9 9 0 1 9 2
45 7 13 8 7 9 15 13 9 15 1 12 9 1 9 13 0 1 12 9 9 1 9 0 7 13 1 9 9 1 9 0 1 8 8 8 8 15 13 0 8 1 9 9 0 2
33 7 13 7 9 9 8 15 13 9 15 8 9 1 9 1 10 9 13 9 1 12 12 9 9 1 9 0 1 9 7 9 8 2
26 7 1 9 9 2 9 0 13 9 1 9 9 1 8 2 9 2 7 9 1 9 8 2 9 2 2
18 7 13 9 9 9 1 9 8 2 9 2 9 1 9 9 9 0 2
35 7 13 9 0 9 1 9 9 1 9 8 1 9 0 2 9 2 7 13 9 9 1 9 1 9 15 13 1 9 12 0 9 0 0 2
19 7 13 9 9 7 9 13 1 9 9 9 9 9 0 0 1 9 9 2
7 9 0 0 1 9 8 8
51 8 2 9 0 2 12 2 12 2 8 8 2 2 13 9 0 8 8 7 9 9 0 8 8 7 9 0 8 8 9 9 9 9 0 15 0 1 9 9 8 8 2 7 13 9 1 9 0 9 9 2
30 7 13 9 7 9 15 13 15 9 13 1 15 8 1 9 9 9 1 0 13 1 12 2 12 8 2 1 9 9 2
25 7 14 13 9 15 13 1 9 9 9 0 1 9 7 0 9 2 7 14 13 0 9 1 15 2
16 7 13 9 9 0 7 8 13 9 9 9 9 1 9 15 2
18 7 13 9 0 0 1 8 8 1 9 9 1 9 1 9 9 9 2
40 7 13 8 9 1 10 9 0 9 9 9 9 1 8 8 8 7 9 9 9 12 1 9 7 1 9 14 13 1 9 0 9 1 9 12 9 9 1 9 2
16 7 13 8 1 9 9 0 0 1 8 8 8 9 1 9 2
19 7 13 9 0 9 0 1 9 8 8 9 9 13 7 13 9 9 9 2
10 9 9 0 2 9 0 1 9 0 9
71 9 12 2 12 2 8 8 8 2 2 13 9 0 9 9 15 0 1 9 9 2 15 13 1 9 9 2 12 2 12 2 9 0 12 2 12 2 9 9 1 9 9 9 1 9 1 9 9 0 1 9 1 9 9 1 9 9 8 11 8 15 13 15 9 1 12 9 2 9 0 2
52 7 13 9 1 0 1 0 9 1 15 1 9 7 13 9 15 0 1 9 12 2 12 2 1 1 13 7 13 9 9 9 15 0 1 9 15 13 1 9 12 2 12 9 0 1 9 1 9 0 1 9 2
38 1 9 15 2 13 9 9 15 0 1 9 7 13 1 1 9 7 13 1 9 12 2 12 2 7 9 12 2 12 2 7 9 12 2 12 1 9 2
48 7 13 9 0 1 9 1 9 9 12 2 12 7 9 13 9 1 9 12 1 12 2 12 1 7 13 8 8 8 9 12 2 12 1 9 12 7 9 0 13 0 1 9 9 12 2 12 2
23 7 1 9 0 13 9 9 0 1 9 1 9 0 15 13 9 1 12 9 12 2 12 2
103 7 13 1 9 8 8 2 12 9 2 8 8 8 2 12 2 8 8 8 8 2 12 2 8 8 8 2 12 2 8 8 8 2 12 2 7 11 8 2 12 2 8 8 8 2 12 2 2 7 1 9 8 8 8 2 12 2 8 8 8 2 12 2 8 8 8 8 2 12 2 8 8 8 8 2 12 2 8 8 8 2 12 2 8 8 8 2 12 2 8 8 8 2 12 2 8 8 8 8 2 12 2 2
17 7 13 9 13 9 3 1 9 12 2 12 2 12 2 12 2 2
8 9 9 8 2 8 1 9 0
47 8 12 2 12 2 8 8 8 2 2 13 8 1 9 0 1 9 9 9 0 1 9 9 15 13 8 9 15 9 12 1 9 15 1 8 12 2 9 1 9 9 0 9 9 1 8 2
14 7 13 8 8 2 12 2 8 8 2 12 2 9 2
9 7 13 8 13 9 8 2 12 2
8 9 9 8 2 8 1 9 0
48 8 12 2 12 2 8 8 8 2 2 13 8 1 9 0 1 9 9 9 0 1 9 9 15 13 8 9 15 9 12 1 9 15 0 1 8 12 2 12 1 9 9 0 9 9 1 8 2
50 7 13 8 8 2 12 2 8 8 2 12 7 12 7 12 2 8 8 2 12 7 12 2 8 8 2 12 1 9 9 2 7 8 8 2 12 2 9 8 2 8 8 2 12 7 12 2 9 8 2
9 7 13 8 13 9 12 2 8 2
8 9 9 8 2 8 1 9 0
48 8 12 2 12 2 8 8 8 2 2 13 8 1 9 0 1 9 9 9 0 1 9 9 15 13 8 9 15 9 12 1 9 15 1 8 8 12 2 12 1 9 9 0 9 9 1 8 2
31 7 13 8 8 2 12 7 12 7 12 2 7 8 8 8 2 12 2 9 8 2 8 8 8 2 12 2 9 8 8 2
9 7 13 9 13 9 12 2 12 2
8 9 9 8 2 8 1 9 0
50 8 2 8 2 12 2 12 2 8 8 8 2 2 13 8 1 9 0 1 9 9 9 0 1 9 9 15 13 8 9 15 9 12 1 9 15 1 8 12 2 12 1 9 9 0 9 9 1 8 2
25 7 13 8 8 2 12 2 8 8 8 2 12 2 9 8 2 8 8 8 2 12 2 9 8 2
9 7 13 8 13 9 12 2 12 2
15 9 8 0 1 9 1 9 1 9 9 0 1 9 9 0
52 8 12 2 12 2 8 8 2 2 13 9 0 8 8 8 1 9 15 1 9 1 9 1 9 15 14 13 9 8 1 9 0 0 2 1 0 2 7 9 14 13 1 15 1 9 1 9 9 1 10 9 2
54 7 13 9 8 1 9 13 15 1 9 15 13 13 15 1 8 1 8 1 9 2 8 8 2 0 9 9 7 15 13 2 9 0 1 9 9 0 2 0 7 2 8 15 8 8 8 1 15 15 9 1 8 2 2
38 8 8 1 9 9 9 0 14 12 15 13 1 9 8 15 13 1 12 1 12 1 9 2 9 8 9 8 1 9 0 15 13 15 9 0 8 8 2
32 7 13 9 0 2 14 8 8 8 1 9 3 7 15 14 13 8 8 9 13 7 13 1 0 15 1 9 9 0 8 2 2
45 7 13 2 14 9 0 15 7 9 9 2 1 8 13 9 0 9 7 13 9 0 9 1 13 9 0 2 8 1 7 15 2 8 8 7 8 1 7 9 9 9 13 0 2 2
64 7 13 8 2 7 1 0 7 15 14 13 1 9 9 7 12 15 14 13 9 0 1 9 0 2 0 2 15 0 0 1 9 1 9 1 9 10 9 7 14 3 7 7 15 14 13 9 1 9 9 7 1 10 9 15 14 13 15 1 9 9 15 2 2
38 7 13 7 13 9 9 9 9 1 9 9 0 1 0 7 15 13 12 9 2 1 9 0 1 8 1 1 9 0 7 9 2 1 7 13 9 9 2
16 8 8 1 9 15 1 9 2 14 13 8 2 1 9 0 2
62 8 12 2 12 2 8 8 8 2 2 13 9 0 0 8 8 1 9 15 1 9 1 9 2 15 13 1 15 9 9 2 7 9 1 8 8 7 14 13 1 9 0 1 9 9 9 1 9 0 7 13 1 7 15 14 13 2 1 9 0 2 2
17 7 14 13 8 9 8 8 15 13 9 0 9 1 0 8 8 2
23 7 13 1 9 0 9 15 8 8 8 15 14 13 9 1 15 1 9 0 1 9 0 2
61 7 13 8 7 15 13 9 1 9 8 2 2 8 8 9 1 8 7 8 8 1 9 9 0 1 9 15 13 1 8 9 9 0 7 13 13 9 0 2 7 8 1 9 3 1 9 9 0 1 9 7 1 9 9 9 8 8 11 8 2 2
53 7 13 8 9 0 1 7 15 2 14 13 9 8 1 9 0 0 1 9 0 1 9 0 2 2 7 13 0 9 1 9 15 1 15 14 13 1 15 8 1 9 15 2 14 13 15 9 7 4 9 3 2 2
39 7 13 2 1 8 8 1 9 9 8 8 9 9 8 8 8 1 9 1 9 1 9 1 9 9 9 15 8 1 15 8 8 1 9 8 8 0 2 2
51 7 13 9 8 0 2 14 8 8 1 9 9 13 1 12 9 8 8 8 1 9 0 13 1 9 9 7 9 1 8 8 1 9 8 8 8 9 9 1 9 0 7 0 7 0 8 8 8 9 2 2
8 9 9 0 1 8 2 0 2
39 8 12 2 12 2 8 8 2 2 13 9 8 8 8 9 9 9 1 9 7 15 13 9 0 1 9 0 1 9 2 9 0 14 13 0 1 9 9 2
36 7 13 9 15 13 1 9 0 15 13 9 0 7 13 1 15 9 0 1 9 0 2 12 9 13 9 1 9 0 0 1 8 2 9 0 2
15 7 13 9 0 1 12 9 7 12 1 9 9 1 9 2
57 7 13 9 15 13 15 9 8 1 9 0 7 9 0 13 12 9 0 1 9 15 13 9 0 1 9 0 1 1 15 9 9 13 8 8 13 1 9 9 9 7 9 0 1 9 13 1 15 9 9 0 14 13 1 15 9 2
36 7 13 8 8 2 7 15 1 9 0 2 9 1 9 7 9 1 1 14 13 9 0 13 9 1 9 9 1 9 9 0 9 0 9 9 2
15 7 1 9 13 8 8 1 9 9 7 8 8 1 9 2
29 7 13 8 8 15 13 9 1 9 0 1 9 0 9 0 7 13 9 9 0 8 8 9 1 9 7 9 0 2
54 7 14 13 9 0 1 9 0 0 2 15 13 9 15 0 1 9 9 2 1 12 9 1 9 9 14 12 9 1 12 15 13 9 15 9 9 2 7 13 9 1 12 9 1 15 12 1 9 9 0 0 9 9 2
33 7 14 13 9 9 0 1 9 7 7 9 0 13 1 9 1 9 9 7 9 9 1 9 0 9 9 0 7 13 9 9 9 2
23 7 1 9 15 13 9 9 0 15 13 9 1 9 2 1 9 9 15 9 1 9 0 2
40 7 13 8 1 9 7 9 0 0 2 13 9 8 8 0 7 13 1 9 9 9 9 9 2 0 2 7 9 1 9 0 0 7 7 9 9 14 13 2 2
33 7 13 9 0 13 12 9 1 15 1 15 9 9 15 14 13 1 9 15 9 9 2 7 1 0 7 8 9 8 9 9 0 2
12 9 13 9 15 1 9 9 9 9 1 9 9
51 9 12 2 12 2 8 8 2 2 13 9 0 9 9 7 15 14 13 1 15 7 13 14 13 9 1 9 9 9 0 1 9 9 15 13 9 2 7 15 7 13 14 13 1 9 0 1 9 1 9 2
42 7 13 9 9 0 8 8 8 7 15 2 1 9 7 8 9 9 9 9 0 1 9 9 2 9 2 1 9 15 13 1 15 9 9 9 9 9 1 10 9 2 2
36 7 13 9 13 1 12 9 2 9 0 9 9 1 9 9 9 0 1 12 9 2 9 0 1 9 9 9 1 9 9 9 9 0 1 9 2
30 7 1 9 2 9 0 13 9 9 0 1 9 9 9 1 9 8 0 1 9 9 9 2 0 1 15 9 9 9 2
33 7 13 8 7 2 9 9 0 13 9 1 10 1 15 8 7 13 9 13 1 9 9 1 9 9 9 1 9 9 9 9 2 2
26 7 13 7 9 13 8 8 1 10 9 1 9 9 9 1 9 0 1 9 0 1 9 0 8 8 2
27 7 13 13 2 8 8 1 9 0 0 9 1 9 0 9 9 15 7 9 9 15 13 9 9 9 2 2
42 7 13 1 7 15 14 13 1 9 9 0 1 9 2 8 2 15 14 13 9 1 9 2 9 9 9 9 1 9 0 1 9 9 7 13 9 0 0 1 9 9 2
32 7 13 8 0 1 12 9 1 8 0 9 9 1 9 9 9 1 12 9 1 9 0 1 9 9 0 7 9 1 9 9 2
8 9 9 9 9 8 2 9 2
34 9 12 2 12 2 8 8 2 2 13 9 0 7 9 13 9 9 9 1 9 13 9 0 9 1 1 7 13 1 9 9 7 9 2
10 7 13 9 7 9 9 14 13 1 2
14 7 13 1 9 9 9 0 9 1 9 1 9 9 2
8 9 8 2 8 8 1 9 9
78 8 2 8 2 12 2 12 2 8 8 8 2 2 13 9 8 8 0 0 7 9 8 8 0 9 9 9 1 9 8 0 0 1 9 9 0 9 9 15 12 12 9 8 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 12 2 12 2 12 2 12 2 7 12 2 12 1 9 9 9 2
15 7 13 9 0 1 9 9 9 1 9 9 1 9 9 2
60 7 1 9 0 2 13 9 8 8 0 0 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 0 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 8 8 8 12 2 12 7 12 2 12 7 12 2 12 2
8 0 12 9 1 9 9 1 9
33 8 12 2 12 2 8 8 2 2 13 12 9 9 9 9 1 9 9 7 8 0 1 9 9 7 13 9 9 1 9 8 8 2
10 8 13 9 0 1 9 15 0 1 8
52 8 2 8 2 12 2 12 2 8 8 2 2 13 9 2 8 2 0 1 8 9 9 7 9 8 13 9 9 0 1 9 15 0 1 8 1 9 9 0 15 13 15 0 9 0 8 8 1 9 8 0 2
28 7 13 9 0 7 9 8 13 9 1 9 15 1 9 8 0 15 13 15 1 8 1 9 12 1 9 0 2
27 7 13 9 0 9 9 8 1 0 1 9 2 9 9 0 1 9 1 9 0 13 1 15 9 0 0 2
31 7 13 10 9 1 9 9 8 1 9 2 7 13 9 9 10 9 12 12 1 1 12 12 1 8 2 1 1 8 2 2
36 7 13 9 0 15 13 1 9 9 0 1 9 0 1 7 9 9 0 14 3 9 7 9 2 14 13 1 9 9 0 7 3 9 0 2 2
38 7 13 9 8 0 7 9 7 10 9 2 13 15 2 9 1 8 2 8 8 8 0 7 9 9 15 1 9 0 7 9 1 9 15 9 0 2 2
6 9 9 0 13 1 9
38 8 12 2 12 2 8 8 2 2 13 9 9 0 8 11 8 9 9 1 9 9 0 9 1 9 0 8 8 11 8 1 9 15 0 8 8 8 2
23 7 13 11 8 1 9 1 9 7 9 15 13 1 9 9 0 1 9 7 9 9 0 2
21 7 14 13 9 8 1 9 9 0 1 9 1 9 13 0 1 9 0 1 12 2
24 7 13 9 9 9 9 0 7 9 1 9 9 0 1 9 0 15 13 15 9 0 7 0 2
13 9 9 0 2 9 0 1 9 1 9 12 2 12
62 9 12 2 12 2 8 8 8 2 2 13 9 9 0 7 0 1 9 12 2 12 2 9 0 12 2 12 2 9 9 1 9 9 9 1 9 1 9 0 0 1 9 1 9 9 1 9 9 8 11 8 15 13 15 9 1 12 9 2 9 8 2
58 7 9 15 0 1 9 1 9 2 0 13 1 9 9 12 2 12 2 7 15 13 13 1 9 12 2 12 2 1 1 14 13 1 9 9 1 9 0 1 15 1 9 1 9 0 1 9 9 0 1 9 15 12 2 12 9 0 2
10 12 9 1 9 9 1 9 1 1 9
34 9 12 2 12 2 8 8 2 2 13 9 9 1 9 8 8 7 12 9 0 13 9 9 9 1 9 9 7 13 0 1 9 9 2
18 7 13 9 7 9 13 1 9 9 9 1 9 7 9 1 9 15 2
24 7 13 9 13 1 9 0 7 9 13 1 9 9 9 0 7 13 9 9 0 7 9 9 2
15 7 13 9 7 10 9 14 13 1 9 0 7 14 0 2
23 2 7 13 9 9 8 0 1 9 0 1 9 0 1 9 8 8 1 8 10 9 2 2
42 7 13 9 1 9 9 8 2 7 0 1 8 8 0 2 13 9 1 9 9 1 9 12 1 9 0 2 12 8 2 7 13 1 15 12 9 9 1 9 12 9 2
25 7 13 9 8 7 8 13 1 2 9 0 2 7 7 9 1 9 9 13 7 13 1 9 2 2
11 9 12 9 1 9 1 9 1 9 1 9
48 9 2 9 0 2 12 2 12 2 8 8 2 2 13 8 12 9 1 1 15 12 9 9 9 7 13 1 12 9 0 1 9 1 9 1 9 0 7 9 2 1 15 13 9 9 8 8 2
27 7 13 9 9 7 13 13 9 15 13 1 9 1 9 0 15 14 13 0 2 1 15 13 9 9 15 2
38 7 13 9 9 0 0 9 9 1 9 2 9 0 1 9 9 9 1 9 1 9 8 1 9 15 1 9 15 7 9 9 7 9 1 9 0 2 2
37 7 13 9 1 9 9 0 1 9 0 8 15 8 1 9 15 9 1 9 8 9 0 7 1 8 8 13 9 15 1 9 1 1 12 12 9 2
13 8 13 9 9 0 1 9 9 9 2 8 2 0
58 8 12 2 12 2 8 8 2 2 13 9 9 0 2 8 8 8 2 1 9 15 0 9 2 7 9 8 8 13 9 9 0 2 8 8 2 1 9 1 9 9 0 2 8 12 2 1 9 9 0 0 1 9 2 8 8 2 2
45 7 1 9 2 9 0 2 13 9 0 1 9 2 8 8 2 15 13 9 8 0 2 1 2 8 8 2 8 13 9 0 2 8 12 8 2 0 9 0 1 9 8 1 9 2
17 7 13 9 9 0 0 13 1 9 12 0 7 13 12 12 9 2
37 7 13 9 9 1 7 9 8 13 7 9 9 0 1 9 9 8 12 13 1 9 9 0 0 1 8 7 13 1 9 9 8 8 9 1 8 2
16 7 13 1 9 1 9 9 9 0 7 13 9 9 10 9 2
71 7 1 12 9 2 9 2 13 9 9 0 8 8 1 7 9 0 1 9 9 12 1 8 8 7 9 9 0 2 1 8 8 8 1 9 9 1 8 7 9 12 9 8 12 1 12 9 2 13 9 1 9 9 0 7 13 1 2 9 9 2 7 13 15 9 2 8 8 2 0 2
13 9 10 14 13 1 12 9 1 9 1 9 9 8
35 8 12 2 12 2 8 8 2 2 13 9 0 9 9 7 15 14 13 1 12 9 13 1 9 13 9 1 9 1 8 1 9 7 0 2
38 7 13 9 1 9 9 1 9 8 8 7 9 15 13 9 1 9 1 9 8 1 8 2 7 9 1 0 2 13 3 1 9 9 1 9 1 9 2
19 7 13 9 9 7 13 0 13 9 9 0 1 9 7 15 13 1 9 2
14 7 13 9 1 9 9 7 13 9 1 9 9 0 2
12 7 14 13 9 9 1 1 9 1 9 9 2
8 10 9 1 9 12 9 2 9
13 12 2 9 0 13 1 9 0 9 0 1 8 2
42 12 2 9 0 0 2 9 9 0 13 9 9 0 13 1 9 2 9 1 9 0 7 13 1 9 9 1 12 9 1 9 9 9 0 7 0 1 15 13 15 2 2
23 12 2 8 2 9 8 0 13 1 9 1 9 15 8 1 9 0 0 13 1 9 15 2
21 12 2 9 0 0 8 8 13 1 8 1 7 13 1 9 15 1 9 12 9 2
17 12 2 9 0 13 12 9 0 2 8 2 1 9 9 0 0 2
23 12 2 9 9 9 9 9 1 9 8 8 13 9 1 9 1 9 8 8 1 9 0 2
8 12 2 9 9 0 8 8 2
9 12 2 9 9 8 8 8 8 2
22 12 2 9 9 0 9 8 8 13 9 9 0 1 9 7 9 1 9 13 12 9 2
21 12 2 9 9 9 0 8 8 8 1 9 15 7 9 15 9 1 9 8 0 2
24 12 2 9 13 1 12 1 9 1 8 8 12 9 1 9 9 9 0 0 1 9 9 0 2
8 10 9 1 9 12 9 2 9
10 12 2 9 9 7 9 0 8 8 2
14 12 2 9 0 13 9 8 8 8 7 9 9 15 2
24 12 2 9 9 8 1 9 9 0 7 8 7 9 0 15 13 9 9 0 1 9 0 0 2
28 12 2 9 8 8 1 9 1 9 12 1 9 9 0 0 0 9 1 9 0 7 9 9 8 8 1 12 2
21 12 2 1 9 9 0 0 1 9 2 13 9 0 1 9 1 9 1 9 8 2
23 12 2 9 0 1 9 13 9 8 8 8 7 9 9 9 13 8 8 8 9 1 9 2
21 12 2 9 0 9 8 13 9 15 13 1 9 0 1 9 9 1 15 1 9 2
20 12 2 9 2 9 1 9 0 2 1 9 8 0 1 9 7 9 0 0 2
25 12 2 8 2 9 8 13 1 9 1 9 13 12 9 1 0 7 13 1 9 1 12 12 0 2
32 12 2 9 9 0 1 8 7 9 1 9 9 9 0 1 8 8 8 9 1 9 1 9 9 1 9 13 1 12 1 8 2
37 12 2 8 1 8 1 9 0 1 12 9 7 9 13 12 9 2 7 1 9 9 15 2 13 9 0 1 0 9 1 12 9 2 8 9 0 2
53 12 2 9 13 9 1 9 9 0 2 9 13 1 12 1 9 9 15 9 2 9 2 13 1 9 12 0 7 9 12 0 1 9 2 7 1 12 1 9 9 15 2 13 9 1 9 1 9 9 1 10 9 2
9 9 0 13 9 9 9 1 8 8
58 8 2 9 0 2 12 2 12 2 8 8 2 2 13 9 0 9 3 9 9 15 1 9 9 9 9 0 0 1 9 8 8 1 9 1 9 1 9 1 9 0 1 9 0 1 9 1 9 9 8 8 1 9 9 12 9 0 2
31 7 13 9 9 1 9 9 0 8 8 8 2 13 1 7 15 14 13 1 9 10 9 7 13 1 9 0 1 9 2 2
29 7 13 2 14 8 8 1 9 1 9 1 9 15 13 9 9 0 2 1 9 0 2 1 9 9 1 8 2 2
58 7 13 9 0 7 13 9 9 9 0 1 9 1 0 9 1 15 1 9 12 2 9 0 0 12 7 8 2 15 14 13 1 9 8 7 14 13 1 8 9 1 12 0 2 7 14 13 1 9 9 9 0 1 9 0 8 8 2
27 7 13 9 0 13 3 1 7 9 9 8 8 13 1 9 0 0 1 9 0 1 9 9 0 1 0 2
16 9 2 9 0 1 9 0 13 12 5 1 9 7 12 1 9
33 8 12 2 12 2 8 8 2 2 13 9 13 15 3 9 9 0 1 9 7 9 0 1 9 0 13 9 9 9 1 9 15 2
49 7 13 10 9 15 13 1 12 12 9 7 12 12 9 2 7 1 12 5 1 9 7 12 5 1 9 13 9 0 1 9 15 1 9 7 9 0 1 9 9 2 0 7 0 2 7 9 0 2
48 7 13 9 0 1 9 7 1 12 5 1 9 7 12 5 1 9 15 13 15 9 2 7 15 13 12 12 9 7 12 9 1 9 9 2 13 1 10 9 1 9 1 9 12 15 13 9 2
35 7 1 9 0 2 3 9 13 1 9 9 9 9 1 9 2 7 9 13 1 1 10 9 12 12 9 9 7 9 12 12 9 1 9 2
35 7 0 13 9 1 7 12 5 1 9 15 13 1 9 0 1 1 9 9 2 13 1 9 1 9 15 1 9 0 1 12 5 1 9 2
11 9 1 9 0 1 9 0 1 9 8 8
47 8 8 2 8 2 12 2 12 2 8 8 2 2 13 9 0 1 8 9 1 9 0 1 9 13 15 9 1 8 8 1 8 2 8 2 8 8 3 1 9 0 1 12 9 1 9 2
40 7 13 9 1 9 9 9 7 7 9 9 15 13 1 9 9 7 9 15 13 1 12 2 14 13 1 9 9 3 14 1 9 9 9 9 1 9 1 9 2
47 7 13 9 9 7 1 15 8 2 14 13 13 1 9 1 9 7 7 9 1 9 13 13 1 15 1 9 8 1 9 2 7 13 9 1 9 0 0 2 8 8 2 14 9 0 2 2
12 7 1 9 2 13 12 7 15 1 9 0 2
8 9 0 13 1 12 8 1 8
39 8 12 2 12 2 8 8 2 2 13 9 9 0 3 9 1 9 2 8 8 2 1 9 0 0 2 1 12 8 1 8 2 7 13 9 1 9 9 2
25 7 13 1 10 9 15 13 9 15 1 12 12 8 2 1 9 13 0 1 8 7 0 1 8 2
25 7 13 9 1 9 9 9 0 8 8 2 7 8 13 1 12 9 0 1 8 13 1 9 9 2
23 7 13 9 9 15 1 7 9 9 12 7 15 9 0 7 9 2 13 7 13 9 9 2
18 7 1 9 10 9 2 13 1 12 8 1 8 1 9 8 8 0 2
11 9 1 8 7 8 1 9 1 9 9 9
46 8 12 2 12 2 8 8 2 2 13 9 2 8 8 2 9 9 7 9 7 8 13 9 9 1 9 9 8 8 0 9 1 9 12 9 0 9 0 9 0 1 9 1 9 9 2
46 7 13 9 1 7 9 0 13 9 9 1 9 1 9 9 0 13 13 9 9 1 9 9 15 13 1 15 0 1 12 9 2 9 1 7 13 9 15 1 9 9 1 8 1 8 2
37 7 13 8 8 1 9 0 9 15 7 9 0 13 9 9 1 9 9 8 1 9 1 9 0 1 9 1 8 1 9 12 1 8 1 10 9 2
58 7 13 9 2 7 15 2 0 2 13 7 8 8 8 9 8 8 14 8 1 15 1 9 1 0 1 9 9 2 7 13 1 0 7 8 9 9 7 7 0 13 9 2 7 13 2 14 15 9 0 13 1 9 9 1 9 2 2
32 7 13 9 1 7 8 14 13 1 9 0 1 9 1 8 1 9 9 9 1 9 0 1 9 1 9 8 14 13 1 9 2
42 7 13 8 8 7 9 0 13 1 9 9 9 9 7 7 15 13 1 9 1 9 9 1 15 1 9 1 9 9 15 1 9 8 1 9 1 8 1 9 0 0 2
6 8 1 8 1 9 9
32 8 12 2 12 2 8 8 2 2 13 9 9 0 7 9 0 8 8 13 9 9 1 8 1 9 9 1 8 1 9 9 2
16 7 13 9 9 15 7 8 14 13 9 15 0 8 8 8 2
36 7 14 13 9 8 0 1 9 15 13 15 1 9 12 9 7 13 1 15 1 8 9 1 9 9 9 0 1 12 9 2 9 1 9 0 2
31 7 13 8 13 1 9 9 8 8 1 12 9 2 9 8 1 1 7 13 1 15 13 1 9 0 1 9 9 9 0 2
17 7 14 13 8 0 0 1 9 9 0 8 1 9 1 9 9 2
34 7 13 8 8 1 9 2 9 12 7 13 8 15 13 1 9 13 1 9 9 1 9 0 1 9 15 1 9 9 15 0 1 9 2
16 7 13 8 9 0 1 9 0 1 9 1 9 2 9 0 2
21 7 1 0 7 13 8 3 9 1 8 8 7 13 7 8 1 10 13 9 8 2
7 13 8 9 9 1 9 8
65 8 12 2 12 2 8 8 2 2 13 9 9 8 9 9 0 1 9 9 9 15 13 15 9 1 9 9 2 7 13 9 0 1 9 0 0 2 8 0 2 1 9 8 9 9 7 13 0 9 0 0 13 1 8 0 1 9 0 15 13 1 12 1 12 2
54 7 13 9 7 15 1 9 8 12 13 12 9 2 7 14 13 12 1 0 0 1 9 9 1 9 1 9 7 0 1 9 9 1 15 8 1 8 0 7 14 13 9 1 15 1 9 0 2 7 9 1 9 9 2
23 7 14 13 9 9 15 1 8 7 1 9 15 12 0 0 1 9 9 1 9 8 0 2
23 7 10 9 0 1 9 0 1 12 14 13 1 0 9 1 9 0 1 9 2 9 0 2
33 7 14 13 9 0 0 8 8 2 8 7 9 8 0 8 8 2 8 3 1 9 9 9 9 1 9 7 9 1 9 9 9 2
10 8 13 9 1 9 9 1 9 1 8
35 9 12 2 12 2 8 8 2 2 13 9 9 0 8 8 9 9 7 13 9 7 9 1 9 9 13 1 15 9 0 1 9 1 15 2
19 7 13 9 0 0 7 8 13 7 13 10 9 2 1 9 9 0 2 2
23 7 13 7 9 14 13 1 9 9 0 7 13 1 9 0 0 1 9 9 0 1 9 2
33 7 13 8 15 13 0 9 1 9 9 7 9 0 14 13 13 1 9 1 1 10 9 1 9 15 13 15 2 9 0 0 2 2
47 7 14 13 9 0 1 9 7 9 1 9 9 0 1 9 9 1 12 9 2 9 0 13 1 9 9 7 13 2 7 9 0 13 1 10 9 1 9 9 1 9 1 9 0 1 9 2
39 1 9 0 13 9 8 8 9 9 0 15 13 9 1 9 9 9 7 8 2 13 15 13 1 9 9 1 9 2 1 9 7 13 15 13 9 1 9 2
29 7 13 9 8 1 9 13 9 1 9 8 0 1 7 9 1 8 13 1 9 7 15 0 1 9 1 9 9 2
7 9 8 2 8 1 9 0
53 8 12 2 12 2 8 8 8 2 2 13 9 8 8 9 0 1 9 8 0 0 1 9 9 0 9 15 12 2 12 12 9 1 9 15 1 8 8 1 8 12 2 12 7 12 2 12 2 12 2 12 2 2
163 7 13 9 8 8 1 9 8 8 12 2 12 2 12 2 12 2 7 12 2 12 7 12 2 12 2 7 9 8 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 8 8 8 12 2 12 7 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 0 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 8 1 0 8 8 12 2 12 7 12 2 8 7 12 2 12 2 8 8 8 1 9 8 8 12 2 12 7 12 2 12 2
122 7 13 9 8 8 1 0 8 8 12 2 12 7 12 2 12 7 12 2 12 2 7 9 8 8 1 0 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 2 12 2 12 2 7 12 2 12 7 12 2 12 2 12 2 12 2 2 7 9 8 8 1 9 15 8 8 8 12 2 12 7 12 2 12 7 12 2 12 2 7 9 9 8 8 1 0 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2
11 9 8 2 9 8 7 9 8 1 9 0
54 8 2 9 0 2 12 2 12 2 8 8 8 2 2 13 9 8 9 9 0 1 9 8 0 0 1 9 9 0 9 15 12 12 9 1 9 15 1 0 8 8 12 2 12 2 12 2 12 2 7 12 2 12 2
24 7 13 9 0 8 8 0 1 9 1 9 15 1 9 8 8 12 2 12 7 12 2 12 2
94 7 13 9 8 8 1 0 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 0 8 8 12 2 12 2 12 2 9 2 7 12 2 12 7 12 2 12 2 7 0 8 8 1 9 8 8 12 2 12 7 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2
119 7 13 3 8 8 1 8 1 9 15 8 8 12 2 12 7 12 2 8 2 7 9 8 8 1 8 8 8 12 2 12 7 12 2 12 2 12 2 12 2 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 8 8 8 8 1 9 8 8 12 2 12 7 12 2 12 7 12 2 12 2 12 2 12 2 2 7 9 8 8 1 9 15 8 8 12 2 12 7 12 2 12 2 7 9 8 8 8 1 0 8 8 12 2 12 7 12 2 12 2
11 9 9 0 0 0 14 13 0 7 9 0
64 8 12 2 12 2 8 8 2 2 13 9 9 8 1 9 9 9 0 9 8 8 9 9 7 9 12 7 12 12 1 9 9 0 0 8 15 13 1 9 12 9 1 9 2 14 13 0 1 9 2 7 9 0 7 9 13 0 1 9 1 9 9 2 2
35 7 13 8 7 2 9 9 9 9 1 0 9 1 9 0 1 9 1 9 2 2 0 7 9 9 1 9 9 0 1 9 1 9 2 2
39 7 13 7 2 14 9 9 15 13 15 9 7 9 9 0 7 9 9 7 9 9 9 2 9 15 9 13 1 9 0 1 15 1 9 1 9 9 2 2
31 7 13 13 2 14 9 9 0 1 9 10 13 7 14 13 15 1 9 15 1 9 9 9 1 9 1 9 9 0 2 2
18 7 13 1 7 15 14 13 0 9 1 9 9 7 9 1 9 9 2
21 7 13 9 0 13 1 9 0 9 7 9 0 1 9 8 13 1 9 9 9 2
20 7 13 9 8 7 2 9 0 9 7 9 9 14 13 7 13 9 15 2 2
33 7 13 1 7 9 9 13 0 1 9 2 7 14 13 1 9 9 9 2 15 13 9 9 7 13 0 1 9 15 1 9 0 2
25 1 9 0 13 9 9 9 8 8 7 9 13 9 9 9 14 7 9 13 0 1 9 1 15 2
34 7 13 2 14 9 0 2 7 15 13 9 9 15 13 1 15 8 0 2 8 8 9 9 0 0 7 15 13 0 7 1 9 2 2
37 7 13 9 1 9 9 9 1 7 0 9 0 14 13 0 1 9 1 9 2 8 7 15 13 1 0 2 9 0 2 7 9 1 9 9 8 2
29 7 13 8 1 9 1 9 9 9 8 8 9 15 2 14 15 13 1 0 0 9 1 9 0 2 1 9 9 2
42 7 13 9 9 1 7 9 9 14 13 1 0 9 0 1 9 9 9 2 7 13 8 1 9 7 2 9 1 9 13 1 9 8 8 8 1 9 9 9 0 2 2
24 7 13 1 0 7 13 9 1 9 1 9 15 1 9 7 9 7 9 1 9 9 1 15 2
20 7 13 9 0 7 9 0 1 12 9 8 7 0 1 15 14 13 9 0 2
38 7 14 13 8 7 15 1 0 9 9 0 1 9 12 8 9 1 9 8 1 9 12 9 9 7 12 9 9 2 1 9 0 13 1 8 8 8 2
26 7 13 9 0 1 9 1 9 0 2 8 2 1 7 15 14 13 9 0 9 0 1 9 3 9 2
35 7 10 9 15 13 1 15 9 15 13 9 1 15 1 12 2 15 0 1 9 9 0 8 8 9 8 1 12 7 13 1 9 12 9 2
9 8 0 13 1 9 0 1 8 0
36 8 12 2 12 2 8 8 2 2 13 9 8 0 8 8 8 9 9 1 9 9 1 9 9 1 0 1 9 1 9 1 9 0 1 15 2
32 7 13 8 1 9 13 15 1 9 9 0 7 12 1 9 1 9 0 1 9 9 1 12 9 1 9 0 1 9 9 0 2
37 7 13 7 15 1 0 9 9 1 9 9 1 9 0 9 1 9 1 9 9 0 0 1 9 12 7 15 13 9 2 12 2 12 2 1 0 2
30 7 13 1 9 9 15 1 7 10 9 1 9 0 13 7 13 1 1 9 9 1 9 12 12 9 0 1 8 0 2
31 7 13 8 2 7 9 0 13 9 1 9 9 13 3 1 9 8 9 9 7 3 1 9 9 9 1 9 9 8 2 2
42 7 13 8 0 1 9 0 1 8 8 8 7 8 8 8 1 9 2 9 0 9 9 0 0 0 1 9 0 9 1 9 2 14 7 8 8 14 13 1 1 9 2
14 9 0 2 9 7 9 2 0 2 1 9 1 9 9
29 9 12 2 12 2 8 8 2 2 13 9 9 0 8 8 9 7 9 7 9 2 0 2 1 9 1 9 9 2
25 7 13 8 1 9 1 9 0 0 2 8 8 0 1 9 7 0 7 8 1 0 9 13 2 2
40 7 13 9 15 13 13 1 9 9 1 8 15 13 15 0 2 14 9 13 1 9 9 9 7 9 3 2 1 15 13 7 15 15 9 0 1 9 9 2 2
45 7 13 8 8 13 9 9 9 8 1 9 12 13 1 9 2 9 8 2 8 9 9 2 13 9 7 14 13 9 1 9 0 1 9 2 1 1 7 13 0 9 1 10 9 2
47 7 13 8 7 15 13 9 1 9 1 9 1 9 9 0 8 8 15 13 9 15 1 9 1 12 9 2 9 1 7 13 9 15 0 1 9 0 2 14 13 0 1 9 7 9 2 2
28 7 1 0 7 13 1 15 9 9 9 0 1 9 8 11 8 1 9 9 0 0 8 8 2 8 8 2 2
27 7 13 8 9 1 9 9 1 9 0 0 9 1 9 9 1 9 9 9 8 8 1 9 9 0 0 2
34 7 13 9 3 9 1 9 9 0 8 8 8 7 9 9 9 0 1 9 9 0 8 8 2 8 8 2 7 0 9 0 8 8 2
27 13 1 7 9 9 13 9 0 1 9 1 9 1 9 8 8 15 13 1 9 1 12 9 2 9 0 2
32 7 13 9 9 2 9 15 0 15 14 13 9 15 2 7 13 9 9 9 0 1 9 15 13 15 9 9 12 9 1 15 2
7 8 13 8 1 9 9 0
32 8 12 2 12 2 8 8 2 2 13 9 9 0 7 9 0 8 8 13 8 9 9 1 9 9 9 1 8 1 9 9 2
13 7 14 13 8 1 9 9 15 0 8 8 8 2
22 7 9 1 9 0 0 1 8 7 14 8 14 13 9 1 8 8 7 13 7 8 2
32 7 13 8 13 1 9 9 8 8 1 12 9 2 9 12 9 1 1 7 13 1 15 13 1 9 0 1 9 9 9 0 2
34 7 14 13 8 0 0 1 9 9 0 8 1 9 1 9 9 2 7 13 8 9 9 7 13 1 9 9 0 2 1 9 0 2 2
34 7 13 8 8 1 9 2 9 12 7 13 8 15 13 1 9 13 1 9 9 1 9 0 1 9 15 1 9 9 15 0 1 9 2
16 7 13 8 9 0 1 9 0 1 9 1 9 2 9 0 2
17 8 13 1 9 9 15 1 8 7 8 13 9 9 15 1 9 9
53 8 12 2 12 2 8 8 8 2 2 13 9 8 1 9 9 1 9 9 15 7 13 8 1 9 0 0 1 8 9 9 2 1 1 13 8 9 9 7 8 1 9 9 15 7 13 9 1 9 9 1 8 2
63 7 13 8 1 9 0 1 9 15 0 1 9 0 1 9 9 9 0 1 8 8 8 1 9 2 9 0 7 15 9 9 1 12 9 9 1 9 15 1 8 8 2 12 9 1 7 0 13 0 9 15 7 1 9 15 8 8 0 9 1 9 0 2
58 7 14 13 9 0 1 9 9 0 8 8 7 8 8 9 8 8 15 14 13 9 1 12 9 2 9 9 12 2 9 9 0 2 7 7 10 9 13 0 1 9 7 9 9 0 13 1 7 15 14 13 0 9 0 1 9 0 2
42 7 13 1 9 0 9 15 8 8 15 14 13 9 1 9 13 1 15 1 9 8 2 7 3 9 9 8 8 8 8 15 14 13 9 1 9 1 9 1 9 9 2
25 7 14 13 8 9 0 1 9 15 13 15 1 9 8 7 15 13 9 9 9 8 0 8 8 2
29 13 7 8 8 0 9 0 0 1 9 9 0 2 12 9 2 13 1 9 8 7 3 9 1 9 1 8 8 2
47 14 9 8 8 8 8 7 13 1 12 9 1 9 15 13 9 8 7 15 8 8 8 8 8 8 8 7 8 2 7 13 9 1 9 9 0 9 9 9 8 8 7 9 9 8 8 2
43 7 13 8 9 8 8 8 8 1 7 13 1 15 1 9 2 7 0 13 1 9 0 1 8 0 9 0 7 13 15 1 9 8 8 8 7 13 9 0 0 1 9 2
47 7 1 9 8 1 8 13 9 8 1 9 1 9 9 0 15 9 8 8 2 8 0 2 7 9 8 8 2 8 8 0 2 2 1 1 13 1 9 0 0 8 8 7 0 8 8 2
22 7 14 13 9 0 1 9 8 8 8 15 13 9 15 9 0 1 9 0 1 9 2
29 7 13 9 8 8 8 9 9 15 15 13 9 9 8 7 13 9 1 9 15 1 8 1 9 0 12 2 12 2
26 7 13 3 9 9 7 9 1 8 7 13 0 1 9 9 8 0 1 9 1 9 0 2 9 0 2
61 7 1 9 0 2 13 8 1 9 1 8 2 7 8 1 9 1 8 2 7 9 1 8 1 9 2 8 8 1 8 1 8 2 8 1 9 1 8 2 7 8 1 8 1 8 2 7 9 8 1 9 1 8 2 7 8 1 8 1 8 2
11 9 8 14 13 1 9 9 9 1 9 8
49 8 12 2 12 2 8 8 2 2 1 0 1 12 9 1 9 1 9 9 1 9 8 0 2 14 13 9 8 15 13 9 15 9 3 14 1 9 0 9 9 9 14 13 1 9 9 9 0 2
25 7 13 9 8 8 8 15 13 9 9 2 9 0 1 9 1 9 1 9 12 8 1 9 9 2
46 7 13 1 9 7 2 9 13 9 1 9 15 1 9 9 9 9 1 7 15 9 0 15 13 7 13 1 9 9 1 8 7 15 13 1 9 9 15 1 9 9 9 9 9 2 2
46 7 13 2 9 9 0 1 9 8 1 9 1 12 8 1 9 9 7 13 9 9 9 15 1 9 9 15 1 12 8 1 0 1 9 9 9 1 9 9 15 13 9 1 15 2 2
55 7 1 15 13 1 9 9 9 0 2 12 9 7 12 12 9 2 15 13 9 1 9 9 9 9 2 13 9 9 9 8 1 2 9 9 1 9 9 0 1 8 7 9 1 9 0 1 9 9 0 1 9 0 2 2
40 7 13 9 1 2 9 15 2 1 2 9 0 1 9 2 9 0 0 0 9 9 9 9 2 7 13 9 0 1 9 9 0 14 3 1 9 9 9 0 2
28 7 13 7 2 9 1 9 9 8 13 9 15 1 9 8 8 15 13 15 9 9 0 7 13 15 8 2 2
24 7 13 2 9 8 1 9 9 1 9 15 1 9 9 0 1 9 0 1 9 9 0 2 2
38 7 13 9 9 0 1 3 1 8 1 9 9 1 9 8 8 8 8 8 1 1 7 13 1 0 9 2 1 1 9 15 13 9 2 0 9 2 2
35 7 13 9 0 1 9 0 1 7 8 14 13 13 9 9 9 0 1 9 15 13 1 15 9 15 7 13 15 7 13 3 1 9 9 2
17 14 7 8 13 9 7 2 9 9 0 13 15 7 13 9 2 2
41 7 13 1 9 8 7 0 15 9 8 8 8 7 8 8 8 7 8 0 1 8 9 2 1 9 1 9 0 12 7 0 15 9 8 8 8 7 8 8 8 2
27 7 13 9 9 9 9 1 9 8 9 9 14 3 9 9 8 8 8 7 8 8 8 7 8 8 8 2
39 7 13 9 0 1 9 9 0 8 8 8 7 9 9 0 0 1 8 8 8 9 9 1 9 15 13 1 9 9 1 9 0 15 13 15 8 1 9 2
11 0 9 0 1 8 10 9 1 9 12 8
44 8 12 2 12 2 8 8 8 2 2 13 8 8 8 8 0 9 0 1 15 10 9 1 9 12 8 15 12 2 12 9 3 9 1 9 0 8 7 13 1 9 2 9 2
45 7 14 13 8 2 12 9 2 9 1 0 9 0 1 9 0 2 0 1 3 9 7 9 15 1 8 8 9 0 7 9 9 15 8 8 13 9 1 9 15 1 9 12 8 2
74 13 7 8 9 12 9 1 9 0 7 9 9 7 9 0 2 13 1 9 0 1 9 9 9 8 1 8 8 9 0 1 8 0 12 8 12 9 2 7 9 9 8 8 8 13 1 9 9 15 1 8 9 1 8 8 9 9 0 2 8 13 9 1 9 12 8 2 7 13 9 14 13 1 2
46 7 13 8 9 0 7 15 14 13 1 9 15 1 8 7 7 15 14 13 9 12 7 12 8 1 8 2 7 13 2 8 8 8 0 2 2 7 13 15 1 15 9 15 8 8 2
50 7 7 8 8 9 8 13 1 9 9 15 7 9 0 1 10 9 13 1 9 9 2 15 14 13 9 9 15 0 1 9 9 0 7 15 13 1 9 9 9 1 0 12 0 1 9 9 7 9 2
46 7 13 9 0 13 8 1 12 9 2 9 9 12 1 9 9 15 9 1 9 8 1 9 15 13 1 15 1 9 8 0 2 7 15 13 9 9 15 0 1 9 9 1 9 9 2
71 7 13 9 9 1 9 0 8 1 9 9 9 1 12 9 2 9 0 1 9 9 9 13 9 15 8 0 7 1 1 12 9 1 0 9 1 15 1 12 9 2 9 12 1 9 8 0 7 13 9 0 1 9 12 8 2 12 2 12 9 2 7 12 8 2 12 2 12 8 2 2
47 14 0 9 0 1 8 1 9 15 7 13 1 12 9 2 9 0 1 9 8 0 7 13 12 2 12 9 7 13 1 9 0 0 1 9 8 8 15 13 9 1 9 12 2 12 9 2
41 7 13 8 9 15 9 0 1 9 8 2 9 9 8 0 2 0 12 2 12 7 13 0 1 9 8 8 8 8 2 9 9 1 9 12 7 12 8 1 9 2
6 8 1 8 1 8 8
40 9 2 8 2 12 2 12 2 8 8 8 2 2 13 9 0 8 8 15 13 15 8 8 8 0 1 9 15 1 9 8 8 0 2 8 14 13 0 9 2
54 7 13 8 13 1 9 8 1 12 9 7 13 9 15 8 8 8 9 1 9 2 7 13 9 15 1 9 2 9 0 1 9 9 7 9 15 1 9 13 0 1 9 8 8 15 13 9 9 8 9 8 8 8 2
36 7 14 13 8 9 8 8 9 8 8 0 7 13 0 1 9 0 2 7 13 3 9 0 0 8 8 2 15 13 9 1 8 9 9 8 2
7 9 8 13 8 1 9 9
38 8 12 2 12 2 8 8 2 2 13 9 8 8 8 8 9 9 7 15 13 9 9 0 0 8 8 3 2 1 7 13 9 0 8 8 9 9 2
31 7 13 8 2 0 9 0 1 9 1 7 9 9 2 1 9 1 9 15 1 9 1 9 0 1 9 9 1 9 0 2
33 7 13 8 1 9 2 8 8 9 3 1 8 2 8 8 14 8 9 1 9 9 7 8 14 13 1 9 9 1 9 9 2 2
19 7 13 7 9 8 1 9 9 13 2 1 9 0 7 9 9 0 2 2
31 7 14 13 8 9 0 1 9 2 7 13 7 9 15 13 1 9 8 1 8 13 13 1 8 9 9 9 0 1 9 2
31 7 13 9 8 1 8 1 9 12 2 12 8 2 0 1 8 7 9 7 13 1 9 8 1 9 9 0 1 9 0 2
40 7 1 9 9 8 8 1 12 9 2 9 0 2 13 8 1 1 12 9 1 1 7 13 1 9 0 1 9 9 0 1 9 0 1 12 9 2 9 0 2
48 7 13 9 9 0 8 8 7 9 15 13 1 7 13 9 7 9 1 9 1 9 9 0 2 7 13 2 8 7 13 2 9 2 9 2 9 0 2 8 8 8 8 8 1 9 0 2 2
23 7 13 8 7 2 8 0 9 0 1 8 7 1 0 1 0 7 13 8 8 9 2 2
27 13 7 12 5 1 9 8 2 12 12 9 2 1 9 2 7 8 15 0 9 1 9 1 7 9 9 2
10 9 0 0 13 1 9 1 9 9 8
47 9 12 2 12 2 8 8 2 2 13 9 1 9 9 9 9 0 0 1 9 9 9 0 8 8 1 9 9 0 8 8 8 9 1 9 8 1 9 7 15 13 9 15 1 9 0 2
28 7 13 1 9 9 9 7 9 0 1 9 8 12 8 9 0 13 9 0 7 9 1 9 9 1 9 9 2
39 7 13 9 8 1 9 1 9 15 7 9 0 0 9 9 1 9 15 14 13 9 15 9 9 13 1 9 8 2 7 8 14 8 1 9 0 1 9 2
12 9 9 0 0 0 1 9 1 9 15 9 9
38 9 12 2 12 2 8 8 2 2 13 9 9 0 9 8 8 8 9 1 9 8 1 9 7 15 0 1 7 15 14 13 9 1 9 15 9 9 2
39 7 13 9 1 9 9 7 15 1 9 9 1 9 15 1 9 0 0 1 9 9 1 9 9 9 0 8 8 1 9 9 15 13 9 15 1 9 0 2
41 7 13 8 8 1 8 8 2 8 8 0 2 8 14 13 9 15 13 9 8 9 2 8 8 8 1 9 9 1 9 15 1 9 2 3 8 9 8 9 2 2
30 7 13 7 9 15 9 8 8 0 1 9 1 9 9 15 1 12 9 14 13 1 8 1 9 15 7 9 1 9 2
34 7 13 9 2 8 8 2 0 9 9 7 9 0 15 13 15 8 8 9 9 0 9 8 8 13 12 12 9 1 9 1 12 9 2
10 9 0 2 9 9 0 2 9 0 2
42 8 12 2 12 2 8 8 2 2 13 8 8 9 9 0 1 9 0 1 9 0 7 9 9 0 13 2 9 0 1 9 9 9 9 7 9 1 9 15 0 2 2
22 7 13 9 9 1 9 8 8 2 10 9 13 9 1 9 0 7 1 9 8 2 2
23 7 13 7 2 9 13 9 0 1 9 9 0 7 9 9 13 0 1 9 7 9 2 2
41 7 8 15 13 9 15 13 1 9 9 1 8 2 8 2 15 13 1 0 1 9 2 9 2 13 1 7 9 0 14 13 9 1 9 1 9 0 15 14 13 2
30 7 13 7 9 9 1 9 15 14 13 1 15 9 0 0 9 15 2 1 9 9 7 9 9 7 9 9 9 2 2
40 7 13 1 9 0 15 13 9 1 9 9 8 8 8 8 2 9 9 0 14 13 1 9 15 9 13 9 15 1 8 2 9 9 2 7 9 9 1 8 2
14 7 13 9 9 0 9 13 9 1 9 2 9 0 2
11 9 1 9 9 14 13 1 9 9 0 0
52 8 12 2 12 2 8 8 2 2 13 9 9 9 0 9 8 8 1 9 13 15 9 9 8 9 9 7 13 2 9 1 9 0 1 9 2 1 9 9 0 8 0 1 9 12 9 1 9 8 1 9 2
22 7 13 8 13 1 9 0 7 3 0 1 9 0 13 1 9 7 0 1 9 9 2
26 7 13 9 8 8 1 9 0 1 9 9 7 9 9 0 1 9 9 14 13 9 9 9 1 15 2
25 7 13 9 0 7 9 7 9 0 1 9 14 13 9 15 7 13 3 9 7 9 1 9 15 2
34 7 13 9 8 9 9 7 9 9 7 9 0 9 1 9 1 8 1 9 8 13 9 9 0 13 1 9 9 9 1 9 9 0 2
20 7 13 9 0 13 9 9 9 9 1 9 0 14 13 0 1 9 9 9 2
24 7 13 12 9 1 9 9 0 1 9 1 9 8 9 9 8 7 14 13 9 13 9 15 2
25 8 12 2 8 8 13 2 2 1 9 0 15 13 1 9 7 9 1 9 9 9 1 9 9 2
84 9 12 2 12 2 8 8 8 2 2 14 13 9 9 0 1 9 9 8 12 8 8 0 9 1 7 9 1 9 0 0 15 14 13 9 10 9 0 1 12 1 12 9 0 2 14 13 0 1 9 0 15 7 9 0 9 13 9 7 9 1 9 10 13 1 9 1 9 9 7 9 1 9 12 15 13 10 9 0 0 1 9 0 2
80 7 13 9 7 15 3 9 9 9 9 0 1 9 2 8 2 8 2 8 2 15 13 9 9 0 1 9 9 1 9 9 9 7 13 1 9 1 9 8 8 2 2 14 9 7 9 2 7 1 9 0 1 9 9 9 2 13 1 12 9 2 7 10 9 15 13 1 1 9 13 0 7 13 1 9 2 9 0 2 2
38 7 13 2 8 7 8 9 1 7 9 1 9 1 15 15 13 1 9 7 9 7 13 9 9 3 7 13 9 9 9 0 13 12 9 1 12 2 2
22 7 13 2 8 7 9 9 1 9 9 8 13 1 9 9 7 9 9 1 9 2 2
34 7 13 9 15 13 1 9 9 9 0 9 1 9 1 7 15 2 13 0 7 15 13 9 7 13 9 13 9 9 7 13 9 2 2
52 7 13 9 9 7 9 13 9 1 9 9 0 1 9 9 9 1 12 9 2 9 0 2 15 13 1 9 0 1 9 9 1 9 3 9 1 9 9 15 0 8 8 1 9 9 1 9 1 9 15 0 2
37 7 13 8 1 7 9 13 9 9 9 9 7 9 7 9 9 1 9 0 1 9 15 1 9 9 9 1 9 9 0 7 9 0 1 10 9 2
28 13 7 9 9 8 8 13 1 9 9 1 9 15 9 9 9 9 7 13 9 10 9 9 1 9 9 0 2
77 7 13 9 0 13 1 9 9 2 9 0 9 0 1 9 9 1 9 9 0 1 9 9 0 7 9 9 9 9 1 15 9 7 7 9 9 14 13 9 9 9 0 7 1 15 9 0 0 15 13 1 12 12 9 0 7 13 1 9 0 7 15 9 9 15 15 8 1 15 9 1 9 0 9 9 12 2
31 7 13 9 1 9 9 1 9 9 15 13 12 9 7 1 0 9 7 9 15 0 9 7 9 1 9 14 13 9 9 2
54 7 1 9 15 14 13 15 9 0 13 8 2 2 3 12 9 0 1 9 9 0 8 8 7 9 1 9 1 12 1 9 8 2 7 14 13 9 1 9 0 7 3 9 7 9 7 15 1 1 9 9 0 2 2
39 7 13 2 14 13 10 9 0 1 0 9 0 1 9 9 8 8 7 9 2 2 7 1 9 1 9 7 7 10 9 14 13 1 9 0 1 9 8 2
26 7 13 9 0 13 9 15 0 9 9 0 2 7 15 14 13 9 15 1 9 0 9 1 9 9 2
23 7 13 9 9 0 13 8 0 1 9 9 1 9 7 13 9 1 9 0 1 9 0 2
3 1 8 8
71 8 12 2 12 2 8 8 2 2 1 9 0 1 9 9 2 9 2 0 2 9 2 9 8 2 13 8 8 9 9 0 9 9 9 15 1 9 0 2 1 8 1 8 8 2 7 14 13 3 9 1 9 12 9 0 2 7 9 9 14 13 13 1 9 9 9 0 1 9 9 2
6 1 9 12 8 8 2
45 8 2 9 8 2 13 9 0 0 7 9 13 2 0 2 1 9 0 0 9 9 0 1 12 9 2 9 0 7 7 9 9 7 9 13 9 9 0 0 1 9 9 9 15 2
6 1 9 12 8 8 2
43 9 2 0 2 9 2 9 8 14 13 9 0 9 9 8 1 9 1 9 8 2 7 13 8 2 9 15 2 1 9 8 7 1 9 0 0 13 15 1 0 9 15 2
6 1 9 12 8 8 2
59 9 2 0 2 9 2 9 8 8 2 1 9 9 0 1 9 0 15 13 9 15 0 1 8 8 2 13 8 8 9 9 1 9 9 15 0 7 13 1 9 9 15 13 1 15 9 15 7 2 9 15 2 0 1 9 0 8 8 2
6 1 9 12 8 8 2
6 9 0 13 9 9 8
55 8 12 2 12 2 8 8 2 2 13 9 9 9 9 7 9 0 8 1 9 15 1 9 7 9 1 9 12 9 1 9 8 0 13 9 9 1 1 9 12 8 8 1 9 8 9 9 8 8 13 9 15 1 15 2
26 7 13 9 9 1 9 12 9 1 9 8 8 0 1 9 12 9 1 8 8 2 8 9 8 0 2
11 7 14 13 9 1 9 7 9 1 9 2
11 7 13 9 9 1 0 12 9 1 9 2
13 9 9 9 1 9 13 1 9 1 9 1 9 9
32 9 12 2 12 2 8 8 2 2 13 9 9 9 1 9 8 8 9 9 9 7 9 0 1 9 9 1 9 1 9 9 2
30 7 13 8 1 9 0 1 9 7 15 2 1 0 9 1 9 9 9 1 9 9 0 7 9 0 13 1 9 2 2
41 7 13 2 8 7 15 8 8 8 1 1 7 8 9 7 9 7 8 10 9 1 9 0 8 8 9 9 1 9 15 9 9 1 1 9 15 1 9 0 2 2
27 7 13 13 2 14 13 3 9 1 9 9 7 9 9 9 2 7 13 9 9 0 1 9 1 9 2 2
34 7 1 0 7 13 8 9 9 0 1 8 1 9 9 13 12 9 1 9 2 13 1 15 1 9 0 9 9 2 9 1 9 2 2
26 7 13 9 15 13 9 1 15 1 0 12 1 9 9 9 0 1 9 0 1 9 9 0 7 9 2
29 7 13 9 1 9 1 9 1 9 9 15 13 9 15 1 9 9 7 9 9 9 9 1 9 15 13 15 9 2
33 7 1 9 13 1 12 9 2 9 0 2 13 9 9 0 11 8 8 7 9 15 13 9 9 1 9 9 15 13 1 9 15 2
28 8 7 8 13 1 9 15 1 9 1 0 1 9 2 9 7 9 0 13 2 9 2 9 1 9 9 9 2
11 8 8 14 13 9 9 15 0 1 9 0
40 8 12 2 12 2 8 8 2 2 13 8 8 9 9 0 9 9 9 15 1 9 0 2 1 8 1 8 8 2 7 14 13 3 9 1 9 12 9 0 2
15 7 9 9 14 13 13 1 9 9 9 0 1 9 9 2
57 7 14 13 9 8 8 2 8 8 2 2 9 2 8 2 8 8 2 0 7 9 1 9 15 8 2 8 2 8 2 8 8 2 7 2 8 8 2 15 13 12 9 0 0 2 1 12 12 9 2 7 13 9 13 1 8 2
58 7 13 9 2 8 8 2 1 9 12 9 9 1 9 0 1 9 2 8 2 2 7 13 9 0 12 0 9 1 15 2 1 9 1 8 7 8 8 7 8 8 8 2 8 8 8 7 8 7 8 8 8 8 8 7 8 8 2
34 7 14 13 9 2 8 8 2 1 8 2 9 2 7 1 8 8 2 9 2 1 9 1 9 1 10 9 0 7 13 12 12 9 2
43 7 13 9 9 9 2 8 8 2 8 8 1 9 15 1 9 2 7 13 1 9 2 14 15 14 13 1 8 8 7 8 8 9 0 1 9 14 13 9 9 15 2 2
49 7 13 2 13 1 9 8 7 13 1 9 1 12 1 0 9 0 2 8 7 8 8 7 8 2 2 7 13 7 9 13 9 1 2 9 8 1 9 0 7 9 9 7 9 0 7 9 2 2
68 7 13 2 8 8 2 0 0 9 9 0 2 1 9 8 2 8 2 8 2 9 8 8 2 2 7 8 2 8 2 8 2 8 8 2 7 8 2 8 2 8 2 8 2 2 7 13 3 9 0 0 13 9 2 8 8 2 13 9 8 2 8 2 8 1 9 0 2
46 7 14 13 10 9 0 1 9 1 9 0 15 13 9 1 9 2 7 9 1 9 9 7 9 9 2 7 13 9 2 8 2 9 2 8 8 2 15 13 9 15 9 8 2 8 2
34 7 13 9 1 9 12 12 9 9 7 12 12 9 1 9 9 1 9 0 1 8 8 13 12 12 9 0 1 9 2 8 8 2 2
58 7 14 13 9 9 1 9 8 2 8 12 9 9 7 12 9 0 1 8 8 2 7 14 13 9 8 2 8 1 12 9 9 9 7 9 0 1 8 8 1 12 7 12 1 12 9 2 15 13 9 1 9 12 1 12 1 9 2
35 7 13 9 1 9 2 8 8 8 8 2 0 8 8 1 9 1 9 8 8 7 9 0 8 2 8 2 14 13 1 9 9 9 2 2
35 7 13 2 8 8 2 1 9 9 9 1 9 0 1 9 9 7 9 13 1 7 9 0 14 13 9 0 1 12 1 12 1 9 0 2
31 7 14 13 9 1 9 1 9 0 1 9 15 13 9 9 1 9 0 7 13 9 2 9 9 1 0 2 1 9 15 2
23 7 1 0 7 13 9 1 9 9 2 9 12 14 7 14 13 1 9 9 0 1 9 2
8 12 9 1 9 9 9 1 8
41 8 12 2 12 2 8 8 2 2 13 12 9 9 15 1 9 9 9 1 9 9 8 9 7 13 13 9 1 15 1 9 9 0 2 7 13 9 0 9 9 2
42 7 13 9 2 8 8 2 7 2 8 8 2 7 9 9 2 0 1 9 13 1 9 12 9 1 9 9 12 0 2 13 1 8 1 9 1 8 1 9 8 8 2
28 7 13 9 9 9 0 0 7 12 9 9 13 13 9 9 1 9 1 9 15 1 9 15 0 7 13 9 2
20 7 1 9 2 13 12 9 1 0 9 1 9 9 1 9 9 9 1 15 2
33 7 13 8 8 0 9 9 0 15 13 9 9 1 9 1 9 15 1 9 0 7 15 13 12 5 1 9 9 0 0 1 8 2
21 7 14 13 9 9 1 9 9 9 0 7 9 1 8 1 9 1 9 1 9 2
13 0 9 9 9 1 9 0 9 9 0 1 9 15
73 8 12 2 12 2 8 8 8 2 2 13 0 9 9 9 1 9 0 8 8 9 0 1 9 1 9 9 1 9 13 9 15 7 13 15 9 8 8 0 2 7 7 15 14 13 9 1 9 0 9 9 15 1 9 0 9 0 1 8 8 0 1 12 9 2 9 1 12 9 0 2 9 2
42 7 13 8 7 15 9 9 0 1 9 1 12 9 9 9 1 9 9 8 13 15 8 8 1 9 8 2 7 15 1 9 0 13 1 9 9 9 15 1 9 0 2
44 7 13 8 2 8 1 9 0 1 9 1 9 9 9 1 9 9 2 2 7 13 2 14 13 8 0 9 0 1 9 1 9 9 0 2 8 8 1 9 10 1 8 2 2
21 7 14 13 8 2 15 13 3 9 9 8 2 9 0 0 1 12 9 1 8 2
54 7 13 8 1 7 13 9 0 9 0 8 1 9 15 2 9 1 7 9 0 1 15 1 9 8 1 9 7 13 1 9 9 2 7 13 1 10 9 2 14 13 9 9 1 9 13 0 1 9 8 1 9 2 2
32 7 13 8 13 1 9 8 8 9 1 9 1 1 0 9 0 1 9 15 1 9 9 7 13 9 8 2 13 0 9 2 2
54 7 13 1 8 7 13 9 1 9 1 9 15 12 9 1 9 7 13 1 10 9 2 2 7 13 9 9 8 8 9 2 7 14 8 8 8 9 0 2 8 9 8 8 0 1 8 8 1 9 1 9 9 2 2
32 7 13 8 1 9 12 1 9 9 1 9 9 8 8 0 2 7 13 1 8 1 9 1 9 9 9 9 0 0 8 8 2
9 9 0 13 9 1 9 9 1 9
45 8 12 2 12 2 8 8 2 2 14 13 9 0 9 9 8 1 9 1 9 8 2 7 13 9 2 9 15 2 1 9 8 0 7 1 9 0 0 13 15 1 0 9 15 2
37 7 13 9 0 15 13 15 8 1 9 9 15 1 9 9 0 1 9 9 15 14 13 1 15 1 8 0 1 9 8 14 9 9 7 13 9 2
49 7 13 9 9 9 9 8 8 8 0 1 9 9 0 2 7 10 9 0 1 9 9 2 7 9 9 14 13 9 15 1 7 9 14 8 2 8 8 8 9 13 2 7 9 13 7 13 2 2
33 7 13 9 1 9 2 15 13 7 9 2 0 2 15 13 9 0 0 1 9 9 0 2 15 1 9 15 1 9 1 0 9 2
32 7 14 13 9 0 0 1 9 9 1 0 8 8 1 9 2 9 0 1 9 9 3 7 13 1 15 0 1 12 12 9 2
40 7 13 9 9 0 2 1 8 8 8 1 8 8 2 9 0 9 7 9 0 9 1 9 8 7 13 8 9 9 1 9 9 15 13 15 8 1 9 8 2
37 7 13 8 8 9 9 8 8 8 1 9 2 7 13 10 9 9 15 14 13 1 15 9 9 15 15 13 15 9 9 1 9 12 7 12 2 2
45 7 13 9 9 1 9 8 7 9 15 1 9 0 2 8 2 8 2 1 9 9 2 7 7 13 9 0 2 7 13 9 15 3 9 1 9 2 7 3 13 9 9 9 0 2
32 7 13 9 8 8 8 9 0 1 9 2 9 0 1 9 9 8 2 9 2 15 13 9 9 7 9 15 9 1 8 0 2
57 7 1 9 2 14 13 9 2 8 2 8 2 8 8 2 15 13 9 2 8 2 1 9 9 7 9 2 8 2 0 1 9 9 0 2 1 9 1 9 2 1 9 9 1 9 2 9 9 2 2 9 9 2 1 9 8 2
53 7 14 9 1 9 1 9 2 7 9 8 1 8 8 2 14 13 9 15 9 8 1 9 2 9 1 9 7 14 13 9 15 13 15 7 13 1 15 9 1 9 0 1 9 0 1 9 7 9 0 1 8 2
49 7 13 9 0 1 9 2 8 2 8 2 9 0 1 9 2 8 2 8 2 8 2 8 2 2 1 9 2 13 3 9 1 9 0 2 1 9 15 0 2 13 1 9 15 13 15 3 2 2
33 7 1 15 0 2 14 13 9 9 0 1 9 8 2 7 9 9 0 1 9 0 1 9 15 2 7 9 9 1 9 0 0 2
29 7 13 8 8 9 1 9 15 2 8 8 1 9 15 9 13 2 7 14 13 1 15 9 7 9 7 9 2 2
66 7 7 3 9 14 9 1 9 15 2 14 14 13 9 2 2 9 1 10 9 2 13 8 8 7 2 13 9 9 2 2 14 9 8 8 7 13 7 2 9 0 1 9 14 13 9 1 12 9 1 9 9 0 2 2 7 9 14 13 1 9 8 8 0 9 2
46 7 15 1 9 2 2 1 10 9 13 8 8 0 1 9 2 8 2 8 2 0 1 9 8 1 9 2 1 12 9 2 14 13 9 10 7 13 9 15 13 1 9 15 0 2 2
5 2 9 1 9 2
78 9 9 0 2 9 13 9 9 12 2 12 2 8 8 8 2 2 13 9 0 9 9 0 0 1 9 0 15 13 15 1 12 0 1 9 15 9 0 1 9 7 13 1 9 9 15 0 12 2 12 2 9 12 2 12 7 12 2 12 7 12 2 12 7 12 2 12 7 12 2 12 2 1 9 0 9 9 2
18 7 13 9 9 15 1 12 9 7 13 9 0 7 1 15 12 9 2
40 7 1 9 0 2 13 9 9 15 0 7 13 1 9 9 9 12 2 12 2 12 2 12 7 12 2 12 7 12 2 12 7 12 2 12 7 12 2 12 2
15 7 13 9 9 9 1 9 0 2 7 9 9 1 9 2
5 2 9 1 9 2
52 9 9 2 8 8 13 0 8 2 9 0 2 12 2 12 2 8 8 8 2 2 13 9 8 8 0 1 9 0 0 1 9 9 9 0 0 9 9 1 8 1 9 15 1 9 9 9 8 8 3 9 2
35 7 14 13 8 1 9 0 1 9 9 15 9 9 7 15 13 9 15 13 15 1 9 8 8 0 1 12 9 1 7 13 12 9 0 2
27 7 13 9 0 1 8 9 12 0 7 13 9 8 8 9 0 7 13 9 0 7 0 1 9 8 8 2
31 7 14 13 9 8 8 2 15 13 1 9 9 9 8 8 1 8 1 9 2 1 9 9 1 9 8 8 8 8 8 2
9 9 0 2 9 0 13 12 9 9
43 9 12 2 12 2 8 8 2 2 13 9 9 9 7 12 9 13 9 1 9 1 9 9 0 0 1 9 8 2 12 9 9 9 2 7 8 2 12 9 1 9 2 2
37 7 13 9 9 7 9 13 1 9 13 15 9 0 1 9 9 9 1 8 1 8 1 1 7 9 0 0 13 0 0 1 8 1 9 9 15 2
31 7 13 9 13 9 1 9 1 8 1 9 9 0 0 13 9 15 1 9 9 0 1 15 13 9 2 8 8 8 2 2
32 7 13 9 7 9 9 13 0 0 12 1 9 0 1 9 9 13 1 12 9 1 9 8 1 8 2 12 9 9 9 2 2
17 7 13 9 2 9 2 7 9 9 13 1 9 9 1 12 9 2
39 7 1 9 9 13 12 9 1 15 12 9 0 1 9 13 1 9 1 9 13 15 9 2 7 13 9 9 2 9 0 1 9 0 1 9 1 12 9 2
4 2 9 8 2
61 9 9 9 0 2 8 1 9 0 7 8 13 1 8 8 2 9 0 2 12 2 12 2 8 8 8 2 2 13 9 0 9 8 8 9 15 1 9 0 1 9 15 0 1 9 9 12 9 9 1 9 0 1 9 9 9 0 1 8 8 2
56 7 13 8 9 9 1 9 9 12 7 12 9 7 12 9 1 12 1 9 2 7 13 1 9 9 0 8 8 15 13 12 8 12 8 12 9 2 7 13 9 0 9 0 1 9 8 8 2 12 8 12 8 12 9 2 2
29 13 7 8 0 1 9 12 9 15 0 9 0 13 1 9 9 1 9 12 8 9 7 15 7 13 1 0 12 2
24 7 13 8 1 9 15 1 9 8 8 0 2 0 1 9 9 15 1 7 9 15 0 9 2
48 7 1 9 12 8 0 2 13 8 8 2 12 8 12 8 12 9 2 7 8 8 2 12 8 12 8 12 8 2 8 8 1 8 1 1 13 8 8 2 12 8 12 8 12 8 2 0 2
58 7 1 9 2 13 9 9 8 8 1 0 8 8 2 12 9 2 1 9 12 8 0 7 13 9 1 9 12 8 12 9 2 8 12 8 12 9 1 0 15 13 0 2 1 1 13 8 8 1 9 0 2 12 8 12 9 2 2
12 7 13 8 8 8 1 9 12 8 0 3 2
44 7 1 9 9 12 8 9 2 13 9 1 8 8 2 12 8 12 8 12 9 2 1 8 8 2 12 8 12 8 12 8 2 7 8 8 2 12 8 12 8 12 8 2 2
12 13 7 9 9 0 7 0 3 13 1 8 2
11 9 9 9 0 13 7 13 1 9 9 9
46 8 12 2 12 2 8 8 2 2 13 9 0 0 9 7 9 9 9 9 0 15 13 1 9 9 8 7 1 9 15 12 9 2 13 7 13 1 9 9 9 1 9 9 9 0 2
45 7 13 9 9 9 0 8 8 15 13 9 15 13 15 9 1 9 1 9 9 7 9 13 1 9 1 9 1 9 0 7 2 14 13 1 15 9 9 2 2 7 13 9 8 2
30 7 13 9 8 2 8 1 9 1 9 9 9 15 13 1 15 9 7 9 9 14 13 1 9 7 13 9 9 0 2
17 7 14 13 9 15 13 15 9 8 1 9 0 9 9 1 9 2
29 7 13 8 7 9 9 0 1 9 0 9 0 1 9 7 9 13 1 9 9 9 9 1 0 9 0 1 9 2
6 9 9 9 9 1 9
31 8 12 2 12 2 8 8 2 2 13 9 0 0 9 9 7 9 9 9 9 8 11 8 8 8 13 9 9 1 9 2
41 7 13 9 0 0 8 8 7 9 0 8 8 13 1 9 0 15 7 1 1 15 9 9 8 8 8 8 8 8 7 9 9 8 8 8 7 9 9 8 8 2
26 7 13 8 7 8 7 9 9 9 13 9 8 1 9 9 13 15 1 9 0 9 9 0 7 0 2
43 7 13 9 0 9 8 11 8 11 8 8 8 9 9 8 8 11 8 8 9 9 7 9 9 11 8 8 9 9 7 9 8 8 11 8 8 9 9 7 9 7 9 2
36 7 13 9 8 1 9 15 7 9 15 1 8 15 2 1 9 9 8 8 7 9 9 9 9 1 8 1 9 15 1 9 9 0 0 2 2
23 13 1 7 9 15 9 0 1 9 13 1 15 9 9 14 13 15 3 1 9 7 9 2
27 7 13 9 9 0 7 9 8 14 13 1 9 10 9 1 9 9 1 0 9 7 9 9 1 9 0 2
23 7 13 9 8 13 9 9 0 7 9 7 8 15 13 1 9 8 8 1 9 8 8 2
6 9 8 13 1 9 8
42 8 12 2 12 2 8 8 8 2 2 13 9 8 1 9 9 9 0 1 9 8 0 8 8 2 12 9 2 1 8 8 9 0 2 7 13 1 0 1 9 15 2
61 7 13 9 9 8 8 9 9 7 8 2 15 13 0 1 9 12 8 1 9 9 9 1 12 9 2 9 0 2 14 13 9 1 9 9 0 14 1 9 9 12 2 9 9 9 9 12 0 7 9 15 7 9 9 15 1 9 1 9 15 2
54 7 14 13 8 2 9 12 9 0 1 9 0 7 9 9 7 9 0 7 9 1 0 9 0 0 2 8 1 3 9 7 9 15 1 8 8 9 0 7 9 9 15 8 8 13 9 1 9 15 1 9 12 8 2
30 7 13 8 9 15 13 1 9 9 8 1 8 9 1 8 8 9 9 0 2 15 2 13 9 1 9 12 8 2 2
41 7 8 13 9 0 2 8 7 13 9 0 2 8 8 14 8 8 8 8 8 1 8 8 8 8 8 9 12 7 12 8 1 8 2 8 8 8 8 0 2 2
35 7 13 9 9 0 1 9 1 8 1 9 9 9 0 1 9 8 15 13 1 9 0 9 14 13 9 1 9 15 13 1 15 1 9 2
32 7 1 9 8 2 14 13 8 1 9 12 8 1 8 1 9 9 12 8 7 15 1 9 8 8 7 8 8 7 8 8 2
8 9 0 13 8 1 9 1 9
40 9 12 2 12 2 8 8 2 2 13 9 9 0 1 9 8 8 9 9 9 9 8 8 1 9 1 9 2 7 15 1 9 0 1 9 13 1 9 0 2
24 7 13 8 1 9 8 0 1 9 9 9 2 14 14 13 3 1 9 0 1 9 0 2 2
42 7 13 7 9 9 2 14 13 13 9 1 9 1 9 15 13 15 9 0 2 0 2 7 15 14 13 1 9 0 7 14 1 9 1 9 7 14 3 9 9 2 2
31 7 13 8 1 7 2 9 0 1 9 1 0 0 1 15 1 9 7 9 7 15 14 13 9 0 7 9 0 0 2 2
27 7 13 9 0 0 1 8 7 13 1 9 9 1 9 1 9 8 8 15 13 1 12 9 2 9 0 2
12 7 13 9 9 9 9 0 1 9 8 8 2
57 7 13 9 15 13 7 9 0 1 10 1 10 9 0 15 13 15 7 13 15 9 12 15 9 15 2 0 2 2 13 1 9 0 1 9 8 8 7 13 9 1 9 9 0 1 9 0 15 13 9 0 0 1 9 0 12 2
14 7 13 9 1 9 1 9 1 9 0 1 0 15 2
8 9 8 9 1 9 1 9 9
37 9 12 2 12 2 8 8 2 2 13 9 9 0 9 9 7 9 9 8 8 8 2 9 9 9 8 8 13 9 1 9 0 1 9 9 0 2
29 7 13 8 1 9 9 9 2 0 8 2 0 7 9 9 0 15 13 1 15 7 13 9 9 9 1 9 12 2
35 7 9 8 13 0 7 9 9 13 13 7 13 8 8 8 9 9 9 1 10 9 7 15 8 13 1 9 9 9 1 9 0 1 9 2
21 7 14 13 8 8 9 1 9 9 7 9 1 9 1 15 13 1 9 9 9 2
16 7 13 9 8 9 0 9 0 1 0 0 0 1 9 0 2
41 7 13 9 8 1 10 9 1 9 13 15 12 9 1 9 12 1 9 9 0 2 9 0 1 8 2 2 9 1 9 0 1 9 8 1 9 2 9 12 2 2
28 1 9 0 13 9 8 8 8 2 9 2 8 8 8 8 8 2 0 2 9 8 8 1 9 0 1 9 2
28 13 1 7 8 7 15 9 9 9 5 8 5 0 15 13 9 0 9 15 2 13 9 0 9 9 0 0 2
54 7 13 9 5 8 5 13 1 9 0 2 9 0 1 9 9 0 15 13 1 9 5 8 5 15 13 1 9 2 9 12 7 13 9 15 1 9 0 7 0 14 0 1 15 1 9 0 13 12 9 1 9 0 2
21 7 14 13 9 9 9 0 8 1 9 2 9 0 1 9 13 15 1 15 9 2
23 7 13 8 13 1 9 9 9 9 1 9 7 13 1 9 0 1 9 13 15 9 12 2
11 8 9 13 8 9 9 9 9 1 9 0
32 9 12 2 12 2 8 8 2 2 13 8 9 7 9 0 9 8 8 9 9 8 8 1 9 9 9 9 0 1 9 0 2
38 7 13 8 1 9 1 9 8 8 2 8 8 8 1 10 9 1 12 9 8 8 8 8 9 0 1 9 9 1 9 0 1 9 1 9 9 2 2
36 8 8 7 9 9 13 1 9 9 1 9 0 0 13 7 12 9 0 13 1 9 1 9 0 1 9 0 1 12 1 9 9 1 9 0 2
43 7 13 8 7 9 9 1 9 1 9 9 0 2 13 9 1 9 0 1 9 0 7 9 9 9 1 15 1 9 9 9 15 0 2 7 13 2 7 15 9 9 2 2
27 7 13 9 8 8 0 0 0 13 1 9 9 9 0 1 9 9 0 7 14 3 9 7 9 7 9 2
10 9 9 0 1 9 9 0 2 9 2
43 8 12 2 12 2 8 8 2 2 1 9 9 9 9 0 2 8 2 15 13 1 9 9 8 1 0 1 3 9 1 1 9 0 7 9 9 7 9 9 0 1 9 2
26 7 13 9 9 9 0 8 8 7 9 14 13 1 15 9 9 15 14 13 9 1 15 1 9 9 2
89 9 0 2 13 9 2 8 8 2 1 8 8 9 1 9 9 0 7 2 1 9 9 9 1 9 0 7 15 8 1 9 8 0 1 9 7 9 2 7 13 9 1 9 9 9 9 2 8 2 7 1 9 9 7 13 1 9 1 0 9 2 8 7 15 14 13 1 9 9 7 9 9 14 13 8 1 12 9 7 14 13 1 15 9 9 9 8 2 2
19 7 13 7 2 9 12 9 14 13 9 1 9 1 9 1 9 8 2 2
32 8 7 9 2 8 2 13 1 7 2 9 9 8 2 12 0 1 9 9 8 13 1 9 1 9 12 9 1 9 12 2 2
31 9 1 2 9 2 0 1 9 0 1 9 9 1 9 15 1 9 2 7 13 9 9 9 12 1 12 9 1 9 9 2
30 9 1 9 9 8 1 9 0 1 9 2 7 1 9 9 1 0 15 7 13 1 9 1 9 9 9 15 1 9 2
13 9 0 0 1 0 9 9 0 1 9 8 7 9
49 9 12 2 12 2 8 8 2 2 13 9 9 7 9 0 0 1 9 9 0 1 9 9 0 15 13 1 9 9 8 1 0 9 9 13 1 15 9 0 1 9 0 8 1 9 8 7 9 2
51 7 13 8 8 9 9 9 9 9 7 9 0 0 1 9 8 8 2 7 15 9 1 9 13 1 15 9 0 1 9 9 13 9 9 0 1 9 1 0 9 9 0 1 9 0 1 9 0 8 2 2
91 7 13 9 8 8 14 13 1 7 0 9 9 0 1 9 9 1 9 15 1 9 2 14 13 1 9 1 9 7 13 0 9 15 13 9 9 12 9 2 9 1 9 2 8 2 1 9 15 1 9 7 9 7 13 9 7 9 15 1 1 13 9 9 0 7 9 15 1 9 1 8 1 9 15 9 2 7 14 13 12 1 9 1 9 8 8 0 1 9 2 2
44 7 13 9 14 13 9 1 9 0 1 1 15 8 8 7 9 15 7 1 3 9 0 9 7 9 7 7 9 7 9 8 9 8 9 15 1 9 7 8 7 13 9 0 2
55 7 13 8 9 15 13 1 15 9 14 13 9 9 9 7 13 9 0 1 10 9 2 9 7 9 0 7 9 0 2 1 9 9 9 1 9 0 7 13 9 15 9 9 1 9 1 8 8 7 8 8 7 9 15 2
110 7 13 9 1 9 9 7 13 9 0 13 1 9 8 0 7 13 8 1 9 9 9 0 13 9 9 15 7 15 9 15 13 7 13 1 9 9 7 7 13 9 0 1 7 13 1 9 1 9 9 8 7 11 1 9 0 1 9 8 7 1 9 1 9 0 15 13 9 9 8 1 9 9 0 9 12 1 9 9 1 9 7 13 9 9 8 8 9 1 9 9 15 13 9 15 1 9 7 9 7 13 1 8 9 12 9 2 9 12 2
8 9 0 13 1 9 9 1 9
38 9 12 2 12 2 8 8 2 2 13 9 9 8 8 9 7 0 9 0 8 8 9 9 1 2 9 9 15 13 9 7 9 0 1 9 9 2 2
49 7 13 8 1 9 13 15 1 8 2 9 2 7 2 9 7 9 7 9 2 0 2 7 9 9 2 8 8 2 14 13 9 7 14 8 1 9 9 0 7 14 3 9 9 1 9 9 2 2
41 7 13 8 8 13 9 15 9 9 0 0 9 0 14 15 2 1 9 9 9 2 0 2 13 7 14 8 9 9 1 9 0 2 1 1 7 13 0 9 0 2
59 7 13 8 7 15 9 1 9 7 2 9 1 9 1 9 7 9 1 9 7 9 9 1 1 13 15 9 0 1 15 1 9 9 1 15 2 7 13 1 7 15 2 7 13 9 1 9 7 14 15 14 13 1 9 9 15 0 2 2
13 7 13 9 9 0 8 9 9 9 14 3 9 2
23 7 13 9 9 1 12 5 1 9 0 9 15 12 12 7 9 15 1 8 0 7 12 2
14 7 13 13 9 0 1 9 15 13 0 1 12 9 2
26 7 14 13 2 9 9 2 7 15 9 9 0 9 1 9 0 2 1 9 9 0 1 9 0 2 2
30 7 1 9 9 13 9 9 0 7 9 0 9 9 7 13 0 1 9 2 7 13 9 10 9 1 9 9 9 15 2
25 7 13 9 7 9 0 0 9 1 9 14 13 9 15 1 9 9 2 1 9 9 7 9 0 2
13 9 0 13 9 1 9 7 1 9 2 2 9 2
39 8 12 2 12 2 8 8 2 2 13 9 9 9 9 0 8 1 9 8 9 1 9 0 9 9 9 8 7 9 14 13 13 9 9 9 1 9 0 2
42 9 9 2 13 9 9 0 0 8 8 9 15 9 9 9 9 1 9 9 2 7 13 9 0 13 1 9 9 15 9 9 1 9 9 13 9 1 9 0 9 9 2
34 7 13 9 0 1 9 0 7 9 9 15 1 9 9 7 1 9 1 9 9 7 9 1 9 1 9 0 1 9 1 9 9 9 2
39 7 14 13 9 9 13 1 9 9 9 7 3 1 9 9 13 1 9 9 0 1 9 2 7 1 0 7 9 9 13 9 1 9 9 9 1 9 15 2
16 7 13 9 9 9 1 7 9 13 9 1 9 1 9 9 2
50 9 9 2 13 15 9 1 9 1 9 9 9 2 8 7 15 13 9 15 1 9 2 7 14 13 9 0 1 7 9 2 8 2 13 1 9 0 13 1 2 9 2 9 0 1 9 8 1 9 2
18 7 13 8 9 9 7 9 9 2 1 1 9 2 15 14 13 9 2
35 14 7 0 9 0 14 13 9 9 9 15 9 9 9 2 7 14 13 9 0 9 1 9 1 9 0 9 14 13 1 9 9 1 9 2
5 8 13 9 9 9
36 8 12 2 12 2 8 8 2 2 13 9 9 0 8 8 7 9 0 13 9 9 9 9 12 9 8 1 9 0 0 8 1 9 9 8 2
29 7 13 9 9 9 9 13 1 9 1 9 9 9 2 7 13 9 9 9 9 9 1 9 9 9 1 9 9 2
31 7 13 8 7 15 14 13 1 15 7 13 3 9 1 9 9 9 15 13 1 9 9 9 9 0 1 9 1 15 13 2
33 7 13 9 9 9 8 8 15 13 9 9 15 13 15 9 1 9 2 1 9 7 13 9 13 1 9 0 1 0 9 0 0 2
40 1 9 0 13 8 8 0 9 9 9 15 13 9 7 9 8 13 15 7 13 1 9 9 1 9 0 0 7 9 13 9 9 13 1 9 9 1 9 9 2
9 9 9 0 0 9 9 2 9 2
28 8 2 7 13 8 1 8 2 8 1 8 2 7 8 1 8 2 7 9 1 8 2 7 8 1 9 8 2
10 12 9 13 1 9 13 1 9 1 9
45 8 8 12 2 12 2 8 8 2 2 13 9 9 8 8 7 12 9 0 1 15 9 7 9 13 13 1 9 1 9 0 1 9 9 2 13 9 9 1 9 1 9 1 9 2
33 7 13 9 10 9 1 9 15 13 1 9 0 1 9 2 8 8 8 8 1 9 15 13 9 15 9 7 13 1 8 8 2 2
65 7 13 9 15 13 7 15 9 0 1 9 9 9 0 9 1 9 2 15 15 9 15 13 15 9 15 7 9 15 7 13 9 0 1 9 1 9 1 9 2 14 15 13 9 1 9 3 7 7 13 14 13 1 15 1 9 7 15 13 9 1 9 15 2 2
16 7 13 9 15 13 9 9 7 13 9 0 2 9 0 0 2
19 7 13 9 0 1 15 9 0 1 9 8 9 1 9 0 0 1 9 2
38 7 13 12 12 9 9 9 15 1 9 8 7 9 15 13 1 9 1 12 9 2 9 0 1 9 9 0 9 1 9 0 1 9 9 9 0 0 2
17 7 14 13 12 1 15 1 9 7 13 9 9 1 15 1 9 2
13 7 13 9 0 1 12 9 1 9 9 1 9 2
31 7 13 9 1 9 8 8 9 7 12 9 2 14 7 9 0 7 1 15 9 9 9 8 8 13 1 15 1 9 0 2
11 9 9 0 1 8 1 9 9 9 1 9
51 9 12 2 12 2 8 8 2 2 13 9 0 7 9 15 13 9 0 0 13 9 9 1 9 2 7 14 13 9 1 9 9 0 8 8 9 9 1 9 7 15 13 7 13 1 15 1 9 7 0 2
25 7 13 9 15 13 15 9 9 0 8 8 9 1 0 0 7 9 1 9 1 9 9 8 8 2
11 9 13 1 9 0 9 9 0 1 9 15
35 9 12 2 12 2 8 8 2 2 13 9 1 9 9 0 0 1 9 9 1 9 13 1 9 0 1 9 0 1 9 7 9 9 15 2
41 7 14 13 9 0 1 9 9 9 7 13 1 15 9 1 9 9 9 15 13 1 9 1 9 8 13 9 9 9 7 9 0 2 1 9 10 13 15 9 0 2
19 7 13 9 7 1 10 9 7 15 8 2 13 9 7 9 1 9 0 2
27 7 13 9 7 9 0 13 9 9 1 9 0 1 9 1 9 8 1 9 0 1 9 1 9 7 9 2
46 7 13 10 9 1 9 8 8 7 9 1 9 0 0 1 9 0 1 9 2 13 9 9 9 1 9 0 2 7 7 15 13 1 9 0 1 9 9 0 1 9 9 0 1 9 2
44 7 13 8 9 9 10 9 7 13 2 1 1 9 2 9 9 8 15 13 1 12 9 2 7 13 9 1 9 15 10 9 3 7 13 2 7 13 2 9 8 1 9 0 2
23 7 13 7 13 9 0 1 12 9 2 9 1 9 1 9 0 1 9 9 15 1 9 2
41 7 14 13 9 0 9 0 9 0 1 8 8 8 1 9 8 0 7 13 9 1 9 12 9 7 9 12 9 1 9 1 9 9 0 0 7 9 1 9 0 2
11 9 9 0 1 8 1 9 9 9 1 9
39 9 12 2 12 2 8 8 2 2 13 9 0 0 9 9 1 9 1 9 9 0 8 8 9 9 1 9 7 15 13 7 13 1 15 1 9 7 0 2
72 7 13 9 9 0 9 9 0 8 8 2 8 7 9 0 9 8 8 7 9 15 8 9 2 9 9 8 0 2 1 15 13 15 1 9 9 9 9 1 9 15 0 2 0 2 8 0 8 8 8 1 8 2 7 13 9 0 9 1 0 9 1 9 9 8 8 7 9 0 1 9 2
18 7 13 9 0 0 7 9 9 0 9 0 8 8 0 3 1 9 2
25 7 13 9 8 7 15 1 0 7 13 9 9 1 9 9 1 8 9 9 7 1 15 12 0 2
16 7 13 9 0 9 9 1 8 1 9 9 1 8 1 9 2
10 9 12 12 1 9 7 9 0 1 8
47 8 2 8 2 12 2 12 2 8 8 2 2 13 9 0 1 9 8 9 9 7 15 13 12 9 0 1 9 1 9 7 9 0 13 1 15 15 13 9 15 1 12 7 12 12 9 2
36 7 13 9 1 9 15 7 15 13 9 1 9 1 9 9 0 0 7 13 9 9 9 9 15 13 13 9 0 1 8 9 8 2 9 2 2
14 7 13 9 7 9 9 0 13 0 1 8 1 8 2
19 7 13 9 0 1 8 1 9 0 1 8 7 13 9 1 9 9 15 2
8 7 14 13 9 7 9 9 2
24 7 13 9 1 9 9 8 1 9 8 8 2 14 9 14 13 0 7 14 8 9 0 2 2
12 9 13 9 1 9 9 0 1 9 9 1 9
43 8 12 2 12 2 8 8 2 2 13 9 9 0 8 8 8 9 9 9 1 9 1 9 1 9 9 7 1 9 1 9 9 15 1 9 0 1 10 9 0 1 9 2
40 7 13 9 0 1 9 0 1 9 1 9 9 9 7 9 14 13 9 14 13 1 9 0 9 8 1 7 15 14 13 2 8 0 2 1 9 13 9 15 2
32 7 13 8 2 14 9 9 14 13 7 13 1 9 2 0 7 15 1 0 1 9 0 7 12 9 9 2 1 9 9 2 2
29 7 1 7 13 1 9 9 8 1 9 13 8 9 8 1 9 8 8 8 1 9 1 9 1 9 9 1 9 2
22 7 13 2 9 13 15 15 0 1 9 9 9 1 9 7 15 15 15 13 9 2 2
29 7 13 9 9 9 2 1 9 13 9 9 1 9 7 1 9 0 13 1 9 9 7 9 7 9 1 9 2 2
44 7 13 9 9 0 9 0 0 1 9 13 9 1 9 9 1 9 0 1 0 7 12 1 9 2 9 0 7 13 7 13 9 15 1 15 1 9 0 9 9 1 9 9 2
24 7 1 9 9 9 15 13 9 9 1 9 9 13 8 1 9 9 15 1 9 9 1 9 2
27 7 13 9 7 9 8 7 9 15 9 14 13 1 9 15 7 7 0 9 0 7 15 13 1 9 0 2
28 1 9 15 13 9 9 1 2 9 9 2 1 9 2 9 9 2 1 9 7 13 1 9 15 1 9 9 2
11 9 8 12 2 8 7 8 1 0 9 0
44 8 12 2 12 2 8 8 8 2 2 13 8 7 8 2 9 0 2 9 9 1 8 9 9 0 0 1 9 9 9 1 9 9 15 13 15 9 7 8 0 3 9 12 2
57 7 13 8 9 9 0 12 9 0 1 9 15 1 7 13 9 0 1 12 7 12 9 2 9 0 7 13 1 9 9 15 8 0 9 1 9 9 1 9 1 9 8 2 7 8 9 0 1 15 1 8 2 7 9 1 8 2
34 7 0 9 1 9 9 0 14 13 1 8 7 8 2 9 0 2 2 7 9 8 2 9 0 2 7 8 8 8 2 9 0 2 2
71 7 13 9 0 9 0 7 12 9 14 13 1 9 15 9 9 12 9 1 12 0 1 9 9 15 13 1 15 12 9 1 9 9 0 1 9 9 13 1 9 9 2 7 13 0 9 13 9 0 1 0 8 2 7 14 13 1 9 9 1 12 0 1 9 9 9 1 8 0 9 2
11 7 13 9 9 0 1 9 12 9 0 2
11 9 0 1 8 7 8 1 9 8 1 8
48 8 12 2 12 2 8 8 2 2 13 8 7 9 0 8 8 7 9 9 0 8 8 13 0 9 9 1 9 9 1 9 0 7 9 0 1 8 15 13 1 15 9 9 0 0 8 8 2
27 7 13 8 1 9 7 8 13 3 8 1 15 13 1 15 7 1 9 0 8 8 1 9 15 0 9 2
22 7 13 9 7 8 7 8 13 1 8 8 1 9 9 9 0 2 0 9 1 9 2
35 1 9 0 13 9 8 2 8 0 1 9 1 9 0 1 8 8 8 8 9 15 9 7 8 13 9 9 15 1 8 2 0 9 2 2
10 9 13 1 9 0 1 9 0 7 0
46 9 12 2 12 2 8 8 2 2 13 9 1 9 1 9 0 1 9 0 0 15 13 9 0 1 9 9 7 13 1 9 9 7 12 9 1 9 15 13 9 9 0 0 9 9 2
68 7 13 9 9 0 8 8 8 1 9 9 13 15 1 9 0 1 9 0 8 8 7 8 7 8 2 14 13 0 1 9 8 8 1 9 7 13 13 1 9 1 8 8 0 7 13 8 8 1 9 9 0 0 1 9 9 9 9 7 9 9 0 7 9 15 0 2 2
32 7 13 0 7 13 12 0 1 9 13 15 9 0 7 0 9 9 7 9 1 9 0 1 9 1 9 9 1 15 13 9 2
45 7 13 8 1 9 15 15 13 15 3 1 9 0 1 9 9 0 7 2 9 15 13 15 9 0 7 0 1 10 9 13 9 0 1 9 13 9 9 0 7 9 9 15 2 2
45 7 13 8 7 2 10 9 13 9 0 1 9 1 9 1 1 9 15 1 9 0 15 13 15 9 0 7 0 7 9 9 1 10 9 15 13 1 9 0 1 9 7 9 2 2
72 7 13 1 7 9 0 2 13 1 9 15 0 7 0 15 13 15 1 15 9 9 0 7 9 9 0 7 9 0 1 9 9 0 1 9 9 1 9 7 9 9 9 7 9 9 15 7 9 1 9 1 9 0 7 0 7 0 15 13 1 15 1 10 9 0 9 1 9 9 0 2 2
49 7 1 9 10 2 13 9 9 9 0 8 8 9 9 2 9 8 9 0 0 1 9 15 1 9 0 1 9 9 15 13 15 9 8 8 1 0 1 9 0 1 9 9 9 9 1 9 2 2
53 7 13 9 9 0 1 9 9 15 7 2 9 13 9 7 9 7 9 9 7 9 7 9 15 7 9 15 0 13 1 9 1 9 7 13 9 15 7 13 9 15 1 9 7 9 7 9 9 9 7 9 2 2
37 7 13 8 7 2 9 9 9 1 9 9 9 1 15 9 9 0 7 9 9 1 9 7 9 1 9 9 1 9 7 9 9 1 9 15 2 2
28 7 13 9 9 0 1 9 9 12 1 9 7 9 0 7 0 15 13 9 9 0 1 9 9 7 9 15 2
17 7 14 13 9 1 10 9 15 14 13 1 9 15 0 9 0 2
35 7 13 9 0 0 7 0 1 9 0 1 9 12 9 7 0 1 12 9 1 12 1 9 13 15 9 8 8 1 9 1 9 0 0 2
11 9 9 7 9 9 1 9 1 8 1 9
44 8 12 2 12 2 8 8 2 2 13 9 0 0 8 8 9 9 7 15 13 9 0 1 9 7 9 9 1 9 1 9 0 1 8 1 9 9 0 1 9 8 9 0 2
50 1 9 0 13 9 2 8 8 8 2 1 9 9 1 9 8 8 8 9 15 7 9 9 0 15 13 1 9 1 9 8 1 9 8 13 1 9 0 9 15 12 8 1 9 2 8 8 8 2 2
39 7 13 7 9 0 13 1 9 1 9 7 9 7 15 9 9 15 15 13 1 9 9 15 13 1 9 2 9 12 1 12 9 1 8 7 9 0 0 2
24 8 8 0 7 9 9 8 9 0 13 12 9 1 15 12 9 7 12 9 14 13 1 9 2
14 9 8 8 13 9 9 15 1 8 8 1 10 1 12
52 8 2 8 2 12 2 12 2 8 8 8 2 2 13 9 9 0 0 8 8 2 12 9 2 7 15 13 9 9 15 1 9 8 8 15 13 1 9 0 1 9 9 1 9 9 0 1 10 1 9 12 2
33 7 13 8 1 9 0 13 9 9 2 8 1 9 8 8 1 10 1 12 2 9 0 1 9 8 8 8 9 7 8 8 2 2
34 7 13 8 0 1 9 8 1 9 9 1 9 0 2 7 15 13 1 7 13 1 9 1 9 14 13 9 1 9 9 1 9 15 2
32 7 13 0 0 13 1 9 8 1 8 9 12 9 1 12 12 9 2 7 13 1 0 12 8 1 9 13 1 15 12 9 2
9 9 9 0 2 8 13 9 9 9
51 8 12 2 12 2 8 8 2 2 13 9 8 1 9 1 9 9 0 8 8 9 15 7 9 0 13 1 9 9 9 9 9 12 9 8 1 9 0 0 2 8 2 1 9 12 9 1 9 9 8 2
29 14 7 9 9 0 9 8 8 13 1 9 7 9 2 9 1 9 2 0 1 9 9 9 15 13 1 9 8 2
30 7 13 7 9 9 9 1 9 0 14 13 1 9 9 2 12 8 8 2 1 0 9 7 13 9 0 1 9 15 2
36 7 13 9 9 9 9 13 1 9 1 9 9 9 2 7 13 9 9 9 9 9 1 9 9 9 1 9 9 15 14 13 9 1 9 15 2
28 7 14 13 0 9 0 1 9 9 9 9 2 7 7 9 9 9 9 0 13 0 9 1 15 1 9 0 2
18 7 13 9 8 9 7 15 13 1 2 9 0 2 1 9 9 9 2
35 7 13 9 7 2 9 9 1 9 0 1 9 9 13 1 9 0 1 9 1 9 2 15 13 9 0 1 0 15 2 7 13 9 0 2
32 7 13 1 7 9 9 13 2 1 9 1 9 2 2 1 15 2 9 0 0 7 9 9 0 7 9 7 9 9 9 2 2
30 7 1 9 9 2 8 2 9 0 1 9 9 9 7 13 9 1 9 0 0 15 13 13 1 9 2 8 8 2 2
38 7 14 13 9 2 8 2 9 9 9 1 10 13 2 7 13 9 8 7 2 9 1 9 9 0 2 13 9 1 9 7 13 1 9 15 1 9 2
34 7 13 9 9 9 0 8 8 15 13 9 9 15 13 15 9 1 9 2 1 9 7 13 9 13 1 9 0 1 0 9 0 0 2
13 7 14 13 3 1 15 9 9 9 1 9 0 2
37 1 9 0 2 13 9 0 9 9 9 0 2 0 7 0 2 15 13 1 9 9 15 13 12 9 8 9 0 1 9 0 1 9 9 9 0 2
33 7 14 13 9 2 8 2 1 9 13 12 8 1 9 8 0 1 12 8 8 7 12 8 8 2 1 9 0 1 8 8 8 2
54 7 10 9 15 13 9 0 9 9 0 7 15 13 14 13 0 1 9 0 0 1 0 1 12 9 2 13 9 9 1 9 9 9 0 7 13 9 0 1 8 1 9 8 8 15 13 9 9 15 1 9 0 0 2
12 9 9 0 2 9 9 8 0 13 1 9 0
44 8 12 2 12 2 8 8 2 2 13 9 1 9 9 9 9 9 7 9 15 13 15 9 9 0 8 2 8 8 2 1 9 9 9 15 8 13 1 9 0 1 9 0 2
38 7 13 8 8 9 9 9 1 9 0 9 1 9 9 8 0 15 13 1 12 9 2 9 0 1 8 7 10 9 14 13 9 1 15 9 9 0 2
31 7 14 13 9 8 8 9 7 15 14 13 9 9 9 9 15 8 15 13 9 15 1 9 9 8 1 9 9 9 0 2
9 11 8 2 9 0 1 9 9 0
35 8 8 12 2 12 2 8 8 2 2 13 9 9 0 1 9 8 11 8 9 9 1 8 8 7 9 13 0 1 9 9 9 1 9 2
43 7 13 11 8 1 9 0 1 9 9 2 14 9 0 1 9 9 0 1 9 1 7 13 9 9 9 0 2 7 1 9 0 8 8 8 2 9 0 2 7 9 2 2
43 7 13 9 0 1 9 9 8 8 1 0 7 12 1 9 2 9 0 1 12 9 2 14 7 15 14 13 1 15 13 1 9 1 9 0 1 9 9 0 1 9 0 2
22 7 13 9 1 9 15 1 9 0 0 1 9 9 9 15 1 9 9 9 8 8 2
19 7 13 11 8 8 8 1 9 0 1 9 9 9 0 1 9 7 9 2
10 8 13 9 1 12 12 9 1 9 9
37 9 12 2 12 2 8 8 2 2 13 9 0 8 8 9 9 7 15 13 9 1 12 12 9 13 15 2 9 0 2 1 9 9 0 1 9 2
57 7 13 8 1 9 1 9 2 8 2 0 2 7 9 0 13 1 9 12 12 9 9 1 9 9 1 9 2 8 8 8 2 7 10 9 13 9 0 0 1 9 2 7 10 9 15 9 9 0 1 9 15 13 8 8 2 2
20 7 13 8 2 3 9 9 0 1 9 1 9 9 8 13 13 9 15 2 2
25 7 13 7 2 9 0 0 2 0 1 9 9 9 14 13 1 9 7 14 13 15 1 9 2 2
45 7 13 9 7 9 8 13 7 2 9 9 0 14 13 9 15 1 9 9 0 2 0 1 9 9 7 3 9 1 9 1 9 9 1 9 9 1 9 5 9 9 5 2 9 2
48 7 13 8 7 10 9 15 13 1 9 8 8 2 12 1 12 9 2 9 2 0 2 0 2 13 1 9 7 8 1 9 8 8 2 8 8 13 9 0 1 9 0 7 0 7 0 2 2
22 7 13 1 9 1 12 12 9 9 15 1 9 0 15 13 1 15 9 9 1 12 2
10 8 8 8 13 1 9 2 9 1 8
44 9 12 2 12 2 8 8 2 2 13 9 0 8 8 8 9 9 1 9 7 15 14 13 9 15 0 8 8 1 9 2 9 0 1 8 1 9 9 9 0 1 9 0 2
23 7 13 9 0 1 9 13 1 9 12 1 9 9 1 9 1 9 9 0 0 1 9 2
10 9 9 0 13 2 9 0 2 1 9
34 9 12 2 12 2 8 8 2 2 13 9 9 0 0 8 8 8 8 8 2 9 0 1 9 0 2 1 9 8 1 9 9 9 2
45 7 13 9 8 0 9 9 1 9 9 9 15 2 1 9 9 13 1 9 0 9 9 9 1 8 8 1 9 7 9 7 9 5 8 8 8 5 0 9 1 9 7 9 2 2
35 7 13 8 8 8 9 0 1 9 0 8 8 8 1 9 8 0 1 9 9 0 7 0 2 1 9 1 9 10 2 1 9 10 9 2
34 7 13 9 0 2 14 9 0 9 1 9 0 2 1 9 7 9 7 9 8 8 8 2 13 1 9 9 1 9 8 2 9 9 2
30 7 13 2 14 8 7 8 10 9 0 1 15 7 1 9 14 13 9 0 1 15 7 13 7 1 9 9 9 2 2
20 7 13 9 0 0 1 9 9 8 1 9 9 9 1 9 9 1 9 0 2
18 7 13 9 2 8 0 2 1 9 0 9 9 7 9 9 1 9 2
23 7 13 2 13 0 12 9 9 1 9 2 14 9 9 13 1 9 1 9 9 9 2 2
23 7 13 9 9 10 1 9 9 0 1 9 1 9 9 0 1 9 9 1 9 1 9 2
45 7 13 9 9 0 7 0 1 9 9 8 9 8 8 8 1 9 9 2 9 0 7 9 7 9 9 13 1 9 0 1 9 9 15 13 2 0 9 2 1 9 0 7 0 2
38 7 13 2 14 9 9 1 9 13 1 9 0 7 13 9 1 9 9 9 1 9 12 1 12 7 13 9 9 1 9 9 14 12 1 12 0 2 2
16 7 13 9 9 9 12 12 9 1 15 12 12 1 12 9 2
8 9 0 0 1 9 9 1 9
29 9 12 2 12 2 8 8 2 2 13 9 0 7 9 0 1 9 9 1 9 13 1 9 0 9 9 1 9 2
55 7 13 9 15 13 9 9 9 15 7 9 0 15 13 15 8 8 2 8 8 2 9 9 9 0 1 9 9 0 13 3 8 8 2 8 8 2 9 9 0 0 8 8 8 8 9 9 8 8 9 0 9 9 0 2
27 7 13 9 0 9 7 0 1 9 9 9 0 8 11 8 14 13 8 1 7 13 9 7 9 10 9 2
33 7 9 1 9 1 9 8 8 8 9 9 9 0 13 9 1 9 9 0 1 9 2 14 2 14 13 9 0 9 1 9 2 2
28 7 13 9 1 9 1 15 7 13 1 0 9 9 0 1 9 1 9 0 2 14 9 8 8 1 15 2 2
41 7 13 9 0 0 13 3 9 7 9 9 0 8 8 13 1 8 0 9 1 9 15 9 9 1 9 9 0 1 9 1 9 9 8 8 1 12 9 2 9 2
24 7 13 9 0 7 9 0 14 13 9 9 9 1 7 13 9 15 1 9 1 9 0 0 2
22 7 13 9 1 9 1 9 8 8 7 2 9 9 0 1 9 0 13 1 9 2 2
23 7 13 9 0 1 9 1 9 7 9 2 9 2 7 13 9 0 1 9 0 8 8 2
30 7 9 1 9 0 7 7 9 9 0 14 13 9 1 9 14 13 2 1 0 9 2 1 9 0 1 9 8 8 2
21 7 13 9 0 7 0 7 0 9 9 15 1 9 0 1 9 1 9 7 9 2
11 9 9 1 9 9 1 9 9 9 0 8
54 8 12 2 12 2 8 8 2 2 13 9 8 1 9 1 9 8 8 9 9 0 9 15 7 9 13 1 9 1 9 9 9 9 9 2 8 2 9 9 9 1 9 9 9 1 9 9 7 13 1 9 9 0 2
28 7 13 9 9 0 8 8 13 1 9 9 7 9 0 13 2 9 9 2 9 9 9 2 8 2 14 12 2
29 14 7 9 9 0 9 8 8 13 1 9 7 9 2 9 1 9 2 0 1 9 9 9 15 13 1 9 8 2
30 7 13 7 9 9 9 1 9 0 14 13 1 9 9 2 12 8 8 2 1 0 9 7 13 9 0 1 9 15 2
59 7 9 2 9 2 15 14 13 9 15 1 9 9 15 9 1 9 13 1 9 9 9 9 9 15 13 1 9 2 7 10 9 15 14 13 9 15 1 9 0 2 13 1 9 1 9 9 1 9 7 13 1 9 9 1 9 1 15 2
19 7 13 9 3 9 0 1 9 7 9 1 9 9 1 10 2 9 2 2
26 7 13 9 7 2 0 15 7 13 9 0 2 2 0 1 7 9 14 14 13 1 9 14 13 9 2
45 14 7 9 9 8 9 8 8 13 9 1 9 1 9 2 8 8 8 2 0 1 7 2 9 9 1 9 9 1 9 15 1 9 12 9 2 14 13 10 9 0 1 9 2 2
20 7 13 7 15 2 1 0 0 7 13 9 1 9 9 1 1 10 9 2 2
7 9 0 0 13 9 9 8
41 8 12 2 12 2 8 8 2 2 13 9 0 0 2 8 8 2 9 9 9 9 9 8 9 2 7 15 9 1 9 1 9 9 0 1 9 1 8 7 8 2
37 7 13 9 0 1 9 2 8 8 2 8 8 7 10 9 13 7 9 9 0 9 7 9 13 1 9 9 9 1 9 8 9 1 9 9 8 2
44 7 13 8 7 9 0 1 9 1 9 0 2 8 8 10 9 7 15 1 9 9 0 0 14 13 9 2 9 2 1 9 1 9 15 0 1 9 9 9 0 1 9 2 2
18 7 14 13 9 1 2 8 8 2 9 9 15 13 1 9 10 9 2
23 7 13 2 8 8 1 9 1 9 0 0 7 13 8 8 7 15 0 1 10 9 2 2
66 7 13 2 1 8 8 9 15 8 1 8 9 9 8 8 15 13 1 9 13 9 9 2 7 1 10 9 8 9 8 5 8 8 12 5 8 1 8 2 0 2 7 9 10 9 7 9 9 5 8 8 12 5 1 9 8 8 8 1 8 13 1 9 0 2 2
27 7 13 9 1 9 9 1 9 1 9 8 8 7 15 2 1 0 9 2 1 15 14 13 9 9 8 2
42 7 13 8 8 13 9 9 9 8 15 13 15 1 9 0 1 9 8 0 1 9 2 8 8 2 8 13 1 8 1 12 9 2 9 0 7 13 1 9 12 9 2
35 7 1 10 9 13 9 8 0 1 9 0 1 9 0 2 7 0 7 2 8 8 2 7 2 8 8 2 8 9 0 15 13 9 8 2
16 1 9 8 9 9 9 8 0 1 9 9 0 0 1 9 2
9 14 9 1 9 8 9 2 0 2
46 8 2 8 2 12 2 12 2 8 8 2 2 13 9 0 1 9 0 0 8 8 9 9 7 9 9 8 8 13 9 9 1 9 15 13 15 1 9 8 1 9 2 9 0 2 2
20 7 13 8 13 1 9 0 1 9 7 9 14 13 9 1 9 9 1 9 2
33 7 9 15 13 1 9 2 14 13 9 9 9 2 9 2 2 1 1 7 13 15 15 2 9 0 15 13 9 15 1 15 2 2
21 7 13 7 8 14 13 1 15 9 1 9 9 1 9 2 1 9 9 0 2 2
33 7 14 13 12 9 7 9 7 9 7 9 13 9 0 7 9 9 7 0 8 9 1 9 8 8 1 1 12 9 1 9 8 2
28 7 13 1 10 9 12 9 0 1 9 2 8 12 2 0 8 9 1 0 1 9 2 9 9 1 12 9 2
38 7 13 9 1 9 1 9 1 9 14 12 0 1 9 8 2 7 14 13 9 0 9 9 1 8 7 14 13 1 9 1 8 1 9 9 1 9 2
41 7 14 13 9 1 9 9 0 0 1 9 9 9 0 8 8 1 9 9 0 8 8 2 7 13 9 9 1 0 9 7 9 9 8 8 7 9 0 1 9 2
17 7 13 1 8 9 9 0 9 8 8 8 1 9 9 9 0 2
36 7 1 8 13 9 1 9 9 9 0 7 9 9 8 8 14 13 1 9 1 9 9 9 0 1 8 2 8 2 1 8 1 9 8 8 2
20 7 13 9 9 0 8 8 1 9 8 8 7 15 14 13 0 9 1 9 2
30 7 13 8 15 3 9 1 9 9 1 9 8 0 1 9 12 9 1 8 1 9 9 15 12 9 1 9 8 8 2
59 7 14 13 0 9 1 9 9 9 1 9 9 1 9 2 7 13 9 7 9 0 13 15 8 8 9 9 0 9 8 8 14 13 13 12 12 9 1 1 9 1 9 7 9 0 1 8 9 8 0 1 8 2 8 8 13 10 9 2
54 7 13 7 13 9 8 8 9 12 12 9 1 9 1 12 9 0 7 9 0 8 8 1 15 13 9 0 2 7 13 1 9 0 13 1 9 2 8 8 2 1 1 9 13 15 9 9 1 9 0 13 1 9 2
11 8 13 1 8 9 1 9 1 9 8 0
29 8 12 2 12 2 8 8 2 2 13 9 9 0 8 8 9 9 1 8 1 9 9 1 12 9 1 8 8 2
18 7 14 13 9 8 9 1 8 9 1 9 8 8 7 8 8 8 2
16 7 9 1 10 9 9 9 0 7 9 9 0 1 9 9 2
35 7 13 9 0 1 8 8 8 7 9 8 0 9 1 9 8 2 13 1 9 0 1 8 1 9 9 8 0 1 9 0 7 12 2 2
10 8 8 8 13 1 9 2 9 1 8
44 9 12 2 12 2 8 8 2 2 13 9 0 8 8 8 9 9 1 9 7 15 14 13 9 15 0 8 8 1 9 2 9 0 1 8 1 9 9 9 0 1 9 0 2
27 7 13 8 1 10 9 1 9 0 0 1 9 0 8 8 8 13 9 1 9 1 9 9 1 9 8 2
33 7 13 8 13 9 9 1 9 15 8 1 9 8 1 9 9 9 9 0 1 9 0 9 15 1 9 9 2 9 0 1 8 2
17 7 13 7 2 9 13 2 1 9 8 8 13 2 9 0 2 2
26 7 13 9 13 9 15 0 1 9 9 12 1 7 13 9 1 9 9 0 1 9 0 0 1 9 2
8 0 9 9 1 9 0 1 9
49 8 2 8 2 12 2 12 2 8 8 2 2 13 9 9 8 8 0 1 8 7 9 0 0 13 9 9 1 8 2 8 2 8 9 9 1 9 12 9 13 15 9 9 9 0 7 13 9 2
18 7 10 9 15 0 1 9 0 1 9 9 9 8 8 8 1 12 2
53 7 14 13 9 9 9 1 9 9 0 1 9 15 13 15 9 1 9 9 2 7 14 13 9 1 9 9 15 9 0 7 13 1 9 9 10 9 0 2 7 13 7 15 14 13 9 1 10 9 14 9 9 2
38 7 13 9 0 1 9 15 1 9 9 0 1 9 9 0 7 9 9 9 0 7 13 9 15 7 9 15 1 9 0 9 1 9 15 13 7 13 2
18 7 14 13 9 0 8 8 8 2 9 8 1 9 2 1 9 9 2
25 14 9 9 1 9 0 7 9 9 9 7 9 15 13 9 9 9 9 7 14 13 1 9 0 2
11 8 2 8 7 8 8 8 13 7 13 8
46 9 12 2 12 2 8 8 2 2 13 9 8 8 8 9 9 1 9 7 9 9 7 8 8 8 13 7 13 9 8 1 9 0 1 9 9 9 0 1 8 1 9 2 9 0 2
31 7 13 8 1 9 0 13 15 1 9 7 2 9 9 8 1 9 9 0 1 15 2 14 13 1 9 9 9 0 2 2
39 7 13 8 13 1 9 9 1 9 0 9 1 15 1 9 9 15 1 9 8 15 13 15 1 0 1 9 2 9 1 9 0 0 1 9 1 9 8 2
11 8 2 0 9 2 1 9 1 8 7 8
34 8 12 2 12 2 8 8 2 2 13 8 9 9 1 2 9 15 0 2 1 9 0 1 9 1 9 0 7 9 9 8 7 0 2
27 7 13 9 1 9 9 0 7 2 8 13 1 9 0 9 9 15 13 1 9 0 1 8 7 8 2 2
41 7 13 9 1 9 0 15 13 1 9 9 9 8 7 0 2 7 13 7 9 10 9 2 0 2 1 9 0 9 2 9 1 9 0 2 13 7 13 1 9 2
27 13 1 7 9 1 0 0 1 8 7 9 0 1 8 7 8 13 12 9 7 9 1 9 0 1 9 2
39 7 9 0 2 13 9 9 0 1 9 2 9 1 9 0 2 9 1 9 9 9 1 9 8 8 12 0 9 1 9 9 7 15 8 8 8 8 8 2
14 9 13 1 7 9 9 9 1 9 13 1 9 9 9
43 8 12 2 12 2 8 8 2 2 13 9 0 1 9 8 8 9 9 7 9 9 9 1 9 0 13 9 1 15 9 10 9 9 7 9 7 7 9 9 9 1 9 2
41 7 13 9 8 8 15 13 9 9 7 9 9 0 2 13 1 15 9 13 9 0 7 13 1 9 0 7 13 1 9 9 9 1 9 0 15 13 1 9 2 2
35 7 13 1 12 5 1 9 0 1 9 0 1 9 9 2 7 14 13 9 8 0 1 9 1 12 5 3 1 9 9 8 8 8 8 2
56 7 13 9 15 13 12 9 13 9 9 7 13 9 15 1 9 2 8 8 8 8 2 7 9 9 9 0 0 1 9 9 9 1 9 14 13 1 12 5 2 14 8 9 9 7 14 13 1 9 1 9 15 1 9 15 2
26 7 13 9 8 7 2 15 13 1 9 9 15 13 7 15 13 9 1 9 10 9 9 7 3 2 2
32 7 13 7 2 9 1 9 9 7 9 0 1 0 2 7 12 1 9 1 9 9 0 1 9 3 7 7 13 9 0 2 2
33 7 13 7 2 9 7 0 13 7 13 1 9 1 9 15 13 9 7 7 13 8 8 9 0 7 0 7 13 1 9 15 2 2
23 7 13 9 0 13 15 9 8 8 13 1 7 8 9 13 1 9 9 7 9 1 9 2
5 8 13 9 1 9
28 9 12 2 12 2 8 8 2 2 13 9 9 0 8 8 9 9 9 1 9 1 9 1 9 9 1 9 2
42 7 13 8 1 9 0 1 9 9 2 7 9 13 8 8 9 0 9 2 8 1 7 13 9 1 9 9 7 1 7 13 9 9 13 8 8 9 0 1 9 2 2
24 7 13 10 9 1 9 9 1 8 7 8 8 9 9 0 1 9 0 0 1 9 8 8 2
40 7 13 8 1 9 0 7 15 1 9 9 1 9 1 9 1 8 8 7 7 10 9 13 9 9 2 7 14 9 9 1 9 9 9 2 7 13 1 9 2
8 9 0 0 1 9 1 9 8
46 8 12 2 12 2 8 8 2 2 13 9 1 9 0 8 7 9 9 0 13 0 13 1 9 15 1 9 9 0 9 0 1 9 8 15 13 1 9 12 9 7 9 1 12 9 2
30 7 13 9 8 1 9 1 9 9 15 7 15 13 9 9 1 8 0 15 13 1 8 2 7 13 9 15 1 9 2
27 7 13 12 9 1 9 9 15 13 1 9 1 9 1 8 1 9 8 1 9 8 1 0 1 9 0 2
25 8 7 9 1 9 14 13 1 15 13 9 8 2 8 1 9 1 9 9 0 1 9 1 9 2
22 7 13 9 9 1 9 8 7 9 0 1 9 9 15 12 8 1 9 8 8 8 2
13 9 8 12 2 9 7 9 13 1 9 0 1 9
48 9 12 2 12 2 8 8 8 2 2 13 9 7 9 9 9 1 9 0 1 9 9 9 8 1 9 9 0 1 9 9 9 0 1 8 1 12 9 0 2 9 1 12 9 2 9 0 2
75 7 13 9 9 9 1 9 9 9 7 13 1 9 9 9 0 15 13 8 7 9 0 7 8 7 8 7 8 2 7 13 9 9 0 1 9 9 0 1 12 9 2 9 0 1 8 8 1 0 9 9 9 8 15 13 15 9 7 13 8 0 7 9 7 9 9 7 13 9 15 1 9 8 3 2
30 7 13 9 13 1 9 9 3 9 1 9 12 2 12 2 7 13 9 8 12 2 12 2 7 13 0 1 9 0 2
89 7 13 9 9 0 9 7 9 2 7 13 9 9 0 7 0 1 9 8 8 9 9 0 15 13 12 9 9 1 9 2 7 13 9 9 7 8 1 9 9 1 12 9 1 9 15 1 9 9 0 1 9 9 9 0 15 13 9 15 7 13 9 1 9 1 9 1 12 1 0 9 2 7 14 13 14 1 9 9 0 1 9 9 7 9 9 1 9 2
42 7 13 9 13 1 9 15 12 1 9 0 2 1 9 12 2 12 2 7 9 12 2 12 2 7 8 12 2 12 2 7 15 0 15 13 1 9 9 15 1 9 2
32 1 9 2 14 13 9 0 0 9 1 9 15 2 7 13 1 9 12 2 12 2 7 13 1 9 12 2 12 1 9 0 2
50 7 13 1 0 9 1 9 0 1 9 9 7 8 9 0 9 1 8 8 13 1 0 1 9 0 2 7 13 9 8 8 9 9 15 1 9 1 8 9 1 1 9 9 0 1 0 9 9 8 2
16 13 7 9 13 1 9 9 9 0 15 13 1 9 9 0 2
14 8 2 13 1 9 9 9 15 3 1 1 9 1 9
49 8 2 9 2 12 2 12 2 8 8 2 2 13 9 9 0 8 8 9 9 1 9 9 1 9 9 7 9 0 0 8 8 7 15 13 1 9 9 9 15 2 3 1 1 9 2 1 9 2
35 7 13 8 1 9 9 9 1 8 1 9 9 0 1 9 11 11 7 2 9 13 1 9 8 0 7 15 13 1 9 9 9 15 2 2
54 7 13 9 0 15 13 9 0 1 8 7 13 9 15 2 14 9 0 1 9 1 9 7 9 1 9 14 13 1 9 9 9 2 2 2 2 2 8 7 15 13 1 9 9 9 15 3 1 1 9 2 1 9 2
24 7 13 8 1 2 9 9 1 9 7 9 1 9 1 9 1 0 12 1 9 2 9 2 2
16 1 9 15 13 8 7 2 9 9 9 0 0 2 1 9 2
51 7 13 2 13 9 9 1 9 15 1 15 7 13 9 1 9 7 9 0 2 2 0 7 2 9 7 9 13 2 1 9 2 9 12 1 9 2 1 9 0 12 1 9 2 9 2 1 9 9 0 2
20 7 13 8 13 8 9 1 7 13 9 9 0 1 8 1 15 13 9 0 2
13 9 9 9 0 1 9 8 9 1 9 7 14 9
39 9 12 2 12 2 8 8 2 2 13 1 9 0 1 9 7 9 9 13 9 0 13 9 9 1 9 8 8 7 13 9 9 9 15 13 1 9 15 2
44 7 13 8 8 1 9 0 1 9 8 8 7 9 2 8 2 9 9 13 1 9 15 1 8 7 13 1 9 7 13 1 9 15 1 9 12 8 1 8 8 1 9 0 2
44 7 13 8 7 15 13 9 9 10 13 1 9 15 7 13 9 9 1 9 0 1 1 9 9 2 7 9 1 9 9 2 13 1 9 9 3 8 8 9 9 2 7 9 2
39 8 7 9 0 1 9 2 9 2 8 8 8 8 8 2 2 13 1 9 1 9 8 8 7 15 13 9 9 10 13 1 9 9 7 9 15 12 9 2
20 7 13 9 9 15 7 9 9 9 14 12 1 9 9 14 13 1 9 15 2
7 9 9 0 1 9 1 8
43 8 12 2 12 2 8 8 2 2 13 9 8 8 0 1 9 12 2 12 8 2 1 9 9 8 1 8 1 9 9 15 0 1 9 1 9 9 0 14 12 1 9 2
36 7 13 1 12 12 9 0 8 1 9 0 1 9 2 7 13 1 9 0 1 9 15 9 1 9 1 9 15 13 1 15 1 9 1 9 2
31 7 1 0 7 13 8 9 0 1 7 13 1 9 15 9 0 0 1 8 7 13 15 1 12 12 9 1 9 9 9 2
11 8 13 9 15 1 9 0 1 9 9 8
55 9 12 2 12 2 8 8 2 2 13 9 0 8 8 1 9 9 9 9 13 12 9 13 1 15 9 9 9 0 1 9 2 8 2 2 0 1 9 15 1 9 9 15 14 13 15 9 1 8 1 9 2 9 0 2
26 7 13 8 1 9 7 2 9 9 8 0 2 7 9 9 1 9 9 2 13 15 8 8 8 2 2
25 7 13 7 15 13 1 7 15 2 0 9 2 1 9 10 9 2 1 9 9 1 9 8 2 2
31 7 13 8 1 9 0 13 15 1 9 7 2 9 9 8 1 9 9 0 1 15 2 14 13 1 9 9 9 0 2 2
48 7 13 1 7 9 13 1 2 9 1 9 8 8 2 7 7 8 2 0 1 9 8 8 7 1 9 9 9 0 2 2 7 13 7 15 2 14 13 7 8 9 13 8 8 10 9 2 2
31 7 13 1 9 2 8 0 2 0 1 2 9 1 9 9 0 2 7 13 9 1 10 9 9 9 7 9 0 1 9 2
31 7 13 8 7 9 9 7 8 8 8 13 7 13 9 8 1 9 0 1 9 9 9 0 1 8 1 9 2 9 0 2
17 7 13 0 7 9 9 9 8 13 7 13 9 12 7 12 9 2
18 7 13 7 12 9 9 9 1 9 8 13 9 15 9 0 1 8 2
39 7 13 7 9 0 8 8 7 9 0 8 8 7 9 0 8 7 9 9 9 8 8 8 13 1 9 0 7 7 15 14 13 9 2 1 8 9 2 2
44 7 13 8 9 9 8 1 2 9 0 2 9 0 0 1 9 9 9 9 15 13 9 9 12 9 2 7 13 1 9 2 9 0 1 9 9 9 7 9 1 9 0 2 2
6 9 0 13 9 0 0
42 9 12 2 12 2 8 8 2 2 13 9 0 8 8 8 8 9 9 1 9 1 9 0 0 9 8 11 8 8 1 9 9 0 7 13 9 9 0 2 8 2 2
43 7 13 9 7 8 7 9 8 2 15 13 1 9 1 9 9 9 0 15 13 15 9 1 12 9 2 9 0 2 13 9 9 9 0 1 0 9 7 9 9 9 0 2
19 7 13 9 7 9 8 13 1 8 9 0 1 9 0 0 8 8 8 2
23 7 1 9 9 13 9 0 0 1 9 9 0 1 9 9 9 0 1 9 9 1 9 2
20 7 13 9 0 9 9 7 9 9 9 9 15 8 9 9 1 9 9 0 2
23 7 14 13 10 9 9 1 9 13 8 1 9 15 13 9 1 15 1 9 9 12 9 2
13 8 13 9 9 0 1 9 9 9 1 0 9 0
32 9 12 2 12 2 8 8 2 2 13 9 0 9 9 9 9 0 1 0 9 0 1 9 9 9 1 9 9 9 8 8 2
20 7 13 9 1 9 8 8 8 7 9 14 13 1 0 7 12 1 9 0 2
21 7 13 9 0 7 8 14 13 9 1 9 9 1 9 7 15 13 9 1 8 2
24 7 0 7 8 13 9 1 8 1 9 12 1 9 15 7 9 12 9 1 9 0 15 8 2
22 7 13 9 9 0 1 9 8 8 9 9 8 1 9 1 9 1 9 0 1 8 2
23 7 13 8 1 9 8 0 1 9 9 9 2 8 13 3 1 9 0 1 9 0 2 2
11 9 8 14 13 1 12 1 12 9 2 9
48 9 12 2 12 2 8 8 2 2 13 9 9 0 1 9 9 9 9 0 1 9 2 8 2 1 8 1 9 1 12 1 12 9 2 9 0 7 13 9 0 0 0 13 9 9 1 9 2
57 7 13 9 15 13 1 9 9 9 0 8 8 1 9 2 7 15 13 9 9 9 15 13 0 9 1 12 1 12 9 2 9 9 1 9 8 7 13 1 9 15 8 8 9 9 9 0 1 9 15 1 12 1 9 9 15 2
35 7 9 1 9 8 13 12 9 9 9 15 1 9 0 1 9 1 8 9 12 7 15 9 7 9 7 9 7 0 7 0 7 9 9 2
21 7 13 9 8 7 9 7 8 7 9 7 9 14 13 1 9 2 0 9 2 2
12 7 13 9 0 1 9 13 1 9 9 12 2
12 7 13 9 0 9 9 9 0 1 9 15 2
7 8 13 9 9 8 1 8
34 8 12 2 12 2 8 8 2 2 13 9 8 8 0 9 9 9 1 8 9 9 0 14 12 0 1 15 2 9 9 7 9 2 2
42 7 13 8 0 1 9 15 1 1 12 12 9 0 13 15 1 9 1 9 9 8 1 8 2 13 8 13 9 15 9 2 13 15 1 9 2 13 8 7 9 2 2
13 7 1 0 7 13 10 9 1 12 1 9 0 2
42 7 13 9 15 13 1 9 0 1 9 15 9 1 9 1 9 15 13 1 15 1 9 1 9 2 13 1 9 15 9 0 0 9 0 1 10 9 0 1 9 2 2
16 7 13 8 9 0 1 9 15 13 15 1 9 9 1 9 2
32 7 1 7 13 9 15 0 13 1 9 9 15 0 2 8 2 1 9 8 0 7 13 15 1 12 12 9 1 9 9 9 2
54 7 13 8 9 15 13 15 1 9 15 9 1 9 8 1 9 0 2 9 12 0 2 14 8 2 13 9 8 0 2 13 9 15 7 9 15 7 9 15 7 9 15 7 9 15 7 13 15 13 1 9 15 2 2
42 7 13 0 2 14 2 14 8 2 2 15 8 1 0 7 12 1 9 0 2 9 12 2 8 8 9 1 9 9 8 8 8 9 9 7 9 13 1 9 15 2 2
10 9 9 14 13 9 1 9 1 9 8
40 8 12 2 12 2 8 8 2 2 13 9 9 0 9 8 8 9 9 9 7 9 9 14 13 9 1 9 1 9 8 1 7 15 2 13 0 1 15 2 2
28 7 13 9 1 9 9 9 0 8 2 8 2 8 2 14 8 9 1 9 1 9 7 14 1 9 15 2 2
60 7 13 2 14 8 1 9 15 13 1 9 2 7 9 0 0 15 7 3 0 13 9 2 8 0 2 14 1 9 1 9 7 14 8 8 13 9 1 9 7 9 13 1 7 15 1 9 9 12 9 2 9 14 13 8 14 13 9 2 2
52 7 13 9 7 15 1 9 14 13 1 9 2 9 0 2 1 9 1 9 1 9 2 7 13 7 9 0 15 13 1 15 13 9 9 1 9 9 2 8 2 13 1 15 9 9 1 1 9 1 9 9 2
21 7 13 9 0 0 1 9 9 1 8 9 9 0 1 9 9 9 9 9 9 2
8 9 9 0 1 9 9 9 0
42 8 12 2 12 2 8 8 2 2 13 9 0 0 1 9 9 0 9 9 0 1 9 9 9 8 0 9 9 9 1 9 9 15 13 15 9 7 13 9 8 8 2
36 7 13 9 0 7 9 9 8 1 9 12 2 12 8 8 2 9 0 1 9 9 9 13 1 9 15 13 1 9 12 9 1 9 9 8 2
33 7 13 9 7 9 14 13 1 9 9 12 7 12 9 0 7 15 13 9 9 1 9 9 7 9 1 9 9 1 9 9 15 2
18 9 0 2 9 13 1 8 1 9 2 9 0 2 1 9 15 1 9
50 8 12 2 12 2 8 8 2 2 13 9 2 8 8 2 0 1 9 15 15 13 9 7 9 0 8 8 13 1 8 1 2 9 0 2 1 9 15 1 9 9 1 9 9 1 9 8 1 9 2
44 7 1 9 15 14 13 9 15 7 7 2 9 9 13 1 7 8 13 1 9 9 9 9 15 2 2 7 1 15 2 13 8 1 9 8 1 9 1 9 0 2 1 9 2
31 7 13 9 7 9 0 1 9 9 0 13 9 9 9 0 7 13 1 9 9 15 1 2 9 0 0 2 1 9 8 2
44 7 13 9 7 9 13 7 13 1 15 8 9 0 1 9 1 9 0 2 0 0 1 9 0 2 9 0 1 8 2 7 1 0 7 13 8 1 10 9 1 9 9 3 2
40 7 13 8 1 8 7 13 9 15 1 9 0 2 1 9 9 9 9 0 0 2 1 9 15 7 7 2 13 0 8 8 2 8 13 9 9 1 9 8 2
23 7 9 1 9 1 9 8 8 13 9 1 9 9 9 0 9 1 10 13 15 9 0 2
5 9 9 9 1 9
41 9 12 2 12 2 8 8 2 2 13 9 9 9 8 11 8 8 8 9 9 9 1 9 0 1 9 1 9 0 1 9 9 1 15 14 13 15 3 1 9 2
52 7 13 9 0 0 7 9 9 8 8 13 1 9 9 9 1 9 15 1 9 0 2 0 2 7 13 15 9 9 8 8 1 9 0 1 9 15 1 9 8 1 8 9 7 13 1 15 1 8 9 9 2
27 7 1 0 7 13 9 9 9 1 9 15 8 1 15 9 1 9 9 0 8 8 7 9 9 8 8 2
31 7 13 9 9 1 9 0 2 9 0 9 9 9 0 2 7 14 13 9 9 8 1 9 9 9 1 9 1 9 0 2
34 7 13 9 9 13 1 0 9 0 1 15 1 9 1 9 2 9 12 2 7 14 13 3 1 9 0 9 9 1 9 1 0 9 2
39 7 13 9 13 1 9 9 15 12 12 9 1 9 0 1 12 9 2 7 13 9 1 12 12 9 1 9 1 9 1 9 9 9 9 13 15 9 0 2
21 7 13 1 12 12 9 1 9 7 13 1 12 12 9 0 9 15 0 1 9 2
8 8 12 2 8 13 9 1 9
52 9 12 2 12 2 8 8 8 2 2 13 9 9 9 8 8 8 1 9 9 8 8 7 15 13 9 1 9 9 8 0 12 1 9 1 12 1 12 9 0 2 9 0 1 9 9 9 15 9 1 9 2
36 7 13 8 2 8 9 1 9 1 8 12 1 9 8 8 9 1 9 2 7 14 8 8 8 1 9 7 8 9 1 9 9 9 9 2 2
67 7 13 8 13 1 9 1 9 9 1 9 2 9 0 7 13 13 1 9 9 8 0 7 9 1 9 9 15 1 9 1 9 9 9 8 8 15 13 1 9 8 12 2 12 2 9 1 7 15 13 9 2 7 13 1 9 0 1 8 7 13 1 9 15 1 9 2
61 7 14 13 9 0 1 9 0 9 1 9 0 1 9 9 9 9 1 9 2 7 15 0 1 9 9 0 1 9 2 7 13 7 9 0 13 15 0 9 1 9 9 2 0 1 9 0 2 9 9 12 2 7 0 1 9 0 2 9 0 2
34 7 13 9 9 0 8 8 13 8 1 9 15 14 13 1 9 1 8 1 12 1 12 9 2 9 0 1 9 9 15 1 9 9 2
42 7 13 9 9 0 9 1 9 15 1 9 9 9 0 1 9 1 0 9 0 1 9 2 7 14 13 9 0 1 9 9 15 14 13 15 9 0 9 2 9 0 2
101 13 7 8 13 1 9 1 9 0 1 9 9 7 9 0 9 12 7 13 9 1 0 1 9 12 9 1 15 12 1 8 9 2 7 13 0 1 9 9 0 0 12 9 2 7 7 15 13 9 1 9 1 9 9 15 1 9 12 9 1 9 9 0 1 9 7 9 9 9 9 1 9 8 0 1 9 8 8 2 12 9 2 7 9 1 9 8 8 7 0 8 8 7 0 8 8 2 12 9 2 2
8 9 0 8 9 15 0 1 9
49 8 2 9 0 2 12 2 12 2 8 8 2 2 13 9 0 9 9 9 9 15 0 1 9 1 12 9 7 15 1 7 13 10 9 1 9 1 9 9 15 13 9 0 7 9 1 9 0 2
39 7 13 9 1 9 9 0 1 9 0 8 8 7 9 0 2 0 1 7 13 7 9 0 8 9 2 12 9 2 9 2 9 9 15 0 1 9 2 2
44 7 13 9 8 8 8 8 8 7 8 2 13 1 9 15 13 15 1 9 0 2 8 8 2 7 15 13 1 9 9 9 1 9 9 9 7 9 1 9 8 8 8 2 2
45 7 13 9 7 9 0 2 13 1 9 0 7 9 9 0 7 1 9 15 1 9 0 1 9 15 1 9 9 9 1 9 0 7 0 0 15 13 9 0 9 9 15 0 2 2
31 7 13 9 8 8 8 8 1 12 7 15 13 1 1 9 1 9 7 9 0 9 9 0 1 9 15 13 15 9 0 2
10 9 8 1 9 2 13 1 9 7 9
54 9 12 2 12 2 8 8 8 2 2 13 9 7 9 1 8 7 9 12 2 9 7 12 2 12 1 9 9 9 1 9 9 9 0 1 9 8 1 9 9 1 9 2 1 12 9 2 15 13 1 9 8 0 2
48 1 9 0 2 13 8 8 2 12 2 8 8 8 2 12 2 9 9 2 7 1 0 2 13 8 8 2 12 2 8 8 11 8 2 12 2 9 9 2 8 8 8 2 12 2 9 9 2
14 9 9 0 2 9 13 0 1 12 12 9 1 9 9
38 9 12 2 12 2 8 8 2 2 13 9 9 0 8 8 8 9 9 7 9 13 0 1 12 12 9 1 9 9 0 1 15 1 9 2 9 12 2
29 7 13 9 9 0 9 1 9 7 2 9 0 0 1 9 1 12 9 13 1 9 9 13 1 12 12 9 2 2
27 7 13 2 7 1 9 13 2 9 2 9 15 13 1 9 9 1 9 12 12 9 1 9 7 9 2 2
85 7 13 9 9 2 14 15 13 9 15 13 1 9 9 9 1 9 1 9 1 9 12 1 9 9 0 2 15 13 1 7 15 2 7 13 9 1 9 0 7 0 13 15 9 7 0 9 0 9 13 7 14 13 9 1 9 0 2 7 13 9 0 0 0 1 9 9 0 2 7 7 1 9 10 9 9 9 9 0 1 9 10 9 2 2
16 7 13 9 1 9 0 1 9 15 9 1 9 2 9 12 2
41 7 1 9 0 2 13 1 15 9 0 1 9 0 2 9 12 7 1 9 9 2 9 1 9 2 2 1 9 9 0 1 9 15 0 1 9 9 0 7 9 2
32 7 13 9 1 9 9 0 7 8 1 9 9 9 0 7 9 7 3 9 9 9 0 1 9 0 0 1 9 9 1 12 2
7 9 0 7 0 13 9 9
26 9 12 2 12 2 8 8 2 2 13 9 0 0 7 9 0 7 0 13 9 9 9 0 9 9 2
50 7 13 9 9 0 0 1 9 9 15 7 2 12 8 0 13 9 0 1 9 8 8 7 8 1 7 13 1 9 1 9 8 0 0 8 13 1 15 7 13 15 1 9 1 9 15 1 8 2 2
40 7 14 13 9 15 13 15 10 9 1 9 9 12 1 9 0 1 9 12 9 7 9 1 12 9 1 9 2 1 9 13 15 8 8 9 1 9 0 0 2
41 7 9 9 13 9 1 9 1 9 0 1 9 0 9 15 13 9 0 1 9 9 7 13 9 7 9 1 9 9 7 12 9 1 9 10 13 9 9 0 0 2
91 7 13 9 9 0 8 8 8 1 9 9 13 15 1 9 0 1 9 0 8 8 1 7 9 0 2 13 1 9 15 0 7 0 15 13 15 1 15 9 9 0 7 9 9 0 7 9 0 1 9 9 0 1 9 9 1 9 7 9 9 9 7 9 9 15 7 9 1 9 1 9 0 7 0 7 0 15 13 1 15 1 10 9 0 9 1 9 9 0 2 2
11 9 9 2 9 9 8 8 0 1 9 9
49 8 12 2 12 2 8 8 8 2 2 13 9 9 9 9 0 0 1 9 9 15 13 1 12 9 2 9 0 2 7 13 9 9 8 8 0 1 9 9 2 13 15 9 8 0 8 8 0 2
44 7 13 1 9 12 9 13 1 12 9 2 13 8 0 8 8 0 8 8 0 2 7 0 8 7 9 0 8 8 0 2 7 0 8 0 7 9 9 8 8 0 8 0 2
26 7 13 1 0 7 13 1 9 3 9 8 0 8 8 0 8 8 13 1 9 0 1 9 9 9 2
14 9 0 2 9 13 9 1 1 12 12 9 1 9 12
46 9 12 2 12 2 8 8 2 2 13 9 0 7 9 9 9 0 13 12 12 9 2 7 1 9 0 1 12 12 9 0 2 1 9 9 1 9 2 9 1 9 2 1 9 12 2
45 7 13 9 9 0 1 9 7 2 9 9 0 13 0 1 12 12 9 2 1 9 0 13 12 12 9 1 9 9 1 0 1 9 2 9 12 1 9 5 9 1 9 5 2 2
34 7 13 9 0 1 9 7 9 2 13 1 9 15 9 15 12 12 9 1 9 9 0 1 10 9 1 0 1 9 2 9 2 0 2
33 7 9 13 9 9 2 9 1 9 2 8 8 9 7 9 0 1 9 9 1 9 1 9 10 9 0 1 9 0 0 1 9 2
29 7 13 8 1 9 0 13 1 9 2 1 0 9 9 10 9 1 9 9 0 7 9 0 7 1 9 0 2 2
39 7 13 9 1 9 1 9 1 9 9 15 13 1 15 1 9 10 9 7 1 9 9 9 1 9 9 0 1 9 1 9 0 7 0 1 10 9 9 2
29 7 13 8 2 15 13 1 9 1 0 9 0 2 7 9 0 13 9 9 2 9 2 1 9 1 9 9 15 2
7 7 13 8 9 9 9 2
15 9 1 9 0 7 9 0 13 9 9 0 1 9 9 9
34 9 12 2 12 2 8 8 2 2 13 9 0 9 9 7 9 1 9 0 7 9 0 13 0 8 8 1 9 9 7 13 9 0 2
63 7 13 9 0 1 9 7 2 9 1 9 0 1 9 1 9 0 13 1 9 9 0 8 8 2 12 9 2 1 8 9 8 7 13 9 1 9 15 13 1 15 1 9 7 13 1 9 15 7 9 15 1 9 9 9 7 14 13 7 13 9 2 2
64 7 13 1 9 1 9 9 1 9 0 7 15 2 1 9 9 9 13 9 1 9 0 13 15 9 1 9 9 0 8 8 1 9 8 1 9 9 7 0 1 9 0 2 7 13 1 9 9 1 1 9 7 13 1 9 1 9 7 13 1 9 15 2 2
30 7 13 9 7 2 9 1 0 15 13 1 15 1 1 9 0 7 14 13 9 9 13 1 9 9 7 9 9 2 2
38 13 9 7 9 0 1 9 12 9 0 1 9 9 9 7 9 1 9 7 9 7 9 1 9 7 9 9 0 7 9 9 0 7 9 9 9 9 2
14 9 8 12 2 9 9 13 9 9 1 9 12 2 12
78 9 12 2 12 2 8 8 8 2 2 13 9 1 9 12 2 12 1 9 1 9 9 0 1 9 12 2 12 2 9 0 12 2 12 2 9 9 1 9 9 9 0 7 0 1 9 9 9 8 1 9 9 15 13 1 9 7 0 1 9 9 9 0 1 8 1 12 9 0 2 9 1 12 9 2 9 0 2
23 7 13 9 9 1 9 9 2 7 13 9 9 1 15 1 15 1 9 15 1 9 9 2
44 7 13 9 9 9 13 1 9 9 0 8 8 8 1 9 0 1 9 9 9 2 7 15 13 1 15 1 14 7 13 9 9 7 13 1 9 1 9 0 9 1 9 15 2
81 7 1 9 2 7 7 13 9 9 13 9 0 1 9 0 1 9 9 8 8 8 1 9 2 13 9 9 13 9 15 8 8 2 7 13 1 9 1 9 9 1 9 1 15 7 13 9 9 9 9 1 9 0 13 1 15 8 7 9 9 7 9 9 7 13 9 0 1 9 7 13 1 15 12 9 1 7 13 8 9 2
16 13 7 9 13 9 9 3 3 9 1 9 9 9 7 8 2
13 9 12 1 9 1 9 0 7 9 9 0 1 9
57 9 12 2 12 2 8 8 2 2 13 9 0 0 9 9 1 9 8 8 7 9 1 9 13 9 9 1 9 0 7 9 1 9 9 0 0 1 9 0 1 9 8 9 9 2 7 13 1 9 12 1 9 0 7 9 0 2
31 7 13 9 0 7 9 1 9 1 9 14 13 9 15 2 13 1 9 13 1 15 9 9 1 9 1 7 13 9 0 2
35 7 13 9 7 15 13 1 9 9 7 9 9 9 0 1 9 9 9 15 1 9 9 1 9 9 0 2 7 13 3 9 0 1 9 2
21 7 13 9 0 1 8 1 8 9 1 9 8 8 9 7 13 9 9 1 0 2
49 7 13 9 9 15 1 7 9 9 9 13 9 15 1 9 7 13 9 15 1 15 1 1 9 9 0 0 0 1 9 0 2 7 13 7 2 9 9 0 13 1 9 0 1 7 13 9 2 2
11 9 0 7 9 9 13 1 9 9 9 0
61 9 12 2 12 2 8 8 2 2 13 9 0 1 9 9 7 9 9 0 2 0 0 1 9 8 2 1 0 9 7 8 1 15 1 9 8 8 1 2 9 9 1 9 1 10 9 7 14 7 7 9 14 13 1 9 0 13 1 9 2 2
38 7 13 1 2 9 9 9 9 0 1 0 9 1 9 9 0 1 9 8 8 2 7 13 1 7 2 9 9 0 13 7 13 9 1 9 9 2 2
40 7 1 9 0 13 9 7 9 1 2 9 1 9 1 9 9 0 1 9 9 0 0 7 9 8 8 1 9 7 9 1 9 9 15 1 9 9 15 2 2
33 13 1 7 9 0 7 9 0 1 8 13 13 1 9 9 0 0 15 13 9 1 9 9 9 0 0 1 12 9 2 9 0 2
13 9 8 12 2 8 2 9 8 1 8 12 2 12
60 8 8 12 2 12 2 8 8 8 2 2 13 9 8 8 0 0 8 8 9 9 15 8 1 9 1 8 12 2 12 1 8 8 9 9 9 1 9 9 0 1 9 9 0 1 9 9 0 8 8 2 8 0 8 8 7 9 8 2 2
18 7 13 8 9 8 2 12 7 12 2 2 8 2 12 2 9 8 2
10 9 8 2 9 9 13 9 1 9 0
44 8 12 2 12 2 8 8 2 2 13 9 9 0 9 9 7 9 1 9 9 13 9 9 9 1 8 9 7 13 1 9 1 9 9 9 9 0 8 0 1 9 9 8 2
38 7 13 9 7 8 14 13 1 9 0 2 0 1 7 9 9 13 1 9 9 3 1 9 0 1 0 1 9 9 1 9 0 1 8 2 8 2 2
10 9 0 0 13 1 9 1 9 9 0
41 9 12 2 12 2 8 8 2 2 13 9 0 0 9 8 11 8 8 9 9 1 9 15 1 9 9 1 9 13 1 9 1 9 9 9 0 15 13 15 9 2
36 7 13 9 9 0 7 9 8 13 9 0 1 9 9 0 0 0 0 1 9 9 9 7 9 1 9 9 9 0 1 12 9 2 9 0 2
20 7 13 1 9 13 1 9 9 7 9 2 13 1 9 0 1 9 9 2 2
21 7 13 9 7 9 0 7 0 9 13 1 9 9 8 7 9 15 0 8 8 2
25 7 13 9 7 9 0 14 13 1 0 1 9 1 9 1 9 9 9 0 1 9 1 9 9 2
30 14 9 0 0 9 9 7 9 1 9 9 15 14 13 9 15 1 9 9 1 9 9 0 7 14 13 3 9 15 2
35 7 14 13 8 9 8 13 1 9 0 8 9 9 8 9 1 9 1 9 9 0 7 1 9 9 0 7 13 9 9 0 2 8 2 2
12 8 2 9 0 1 9 1 9 0 14 13 0
49 8 12 2 12 2 8 8 2 2 13 9 0 0 1 9 0 8 8 9 9 7 9 0 14 13 0 1 9 1 9 9 0 1 9 1 9 8 9 7 13 9 7 9 0 1 9 9 0 2
45 7 13 8 1 9 1 12 9 13 1 9 7 9 0 7 9 0 0 1 9 1 9 0 1 9 9 8 8 0 2 0 15 13 1 12 1 12 9 2 9 0 1 9 8 2
32 7 13 8 7 2 9 2 8 2 8 13 9 9 15 1 9 9 7 9 1 0 7 15 13 7 15 0 1 9 9 2 2
26 7 14 13 9 9 0 8 8 7 9 9 0 8 8 1 9 1 8 8 7 9 13 1 9 9 2
22 7 8 13 7 9 13 0 13 0 1 9 0 1 9 0 1 9 7 9 9 0 2
24 7 13 7 2 9 15 14 13 0 13 9 15 2 2 2 2 2 7 13 9 9 9 2 2
22 7 1 0 7 13 8 9 8 1 9 9 2 7 14 13 9 9 1 9 9 15 2
8 10 9 1 9 12 9 2 9
13 12 2 9 0 0 8 8 2 13 1 12 2 2
43 12 2 8 9 8 8 8 13 1 9 7 1 15 1 8 1 9 13 15 9 9 8 8 2 7 1 12 9 13 9 0 1 9 1 9 13 8 7 13 8 1 9 2
10 12 2 9 13 9 1 9 9 0 2
16 12 2 9 0 1 9 9 9 9 0 13 1 9 9 8 2
14 12 2 9 9 9 0 8 8 2 13 1 12 2 2
21 12 2 9 0 13 1 8 1 9 1 9 8 8 1 9 8 8 0 1 8 2
8 10 9 1 9 12 9 2 9
11 12 2 9 8 8 9 1 9 1 8 2
5 12 2 9 8 2
13 12 2 9 9 0 8 8 2 13 1 12 2 2
9 12 2 9 9 0 1 8 0 2
11 12 2 9 9 8 0 8 8 1 8 2
8 12 2 9 9 0 8 8 2
14 12 2 8 2 8 8 13 0 9 9 9 1 8 2
9 9 9 0 1 9 9 1 9 8
60 8 12 2 12 2 8 8 2 2 13 9 9 8 2 8 2 8 8 1 9 0 9 15 7 9 0 1 9 9 14 12 1 9 0 0 8 1 9 8 14 8 1 9 9 9 9 7 9 9 14 13 1 9 1 9 1 9 9 9 2
34 7 14 13 9 1 9 8 1 9 9 12 3 2 7 14 13 9 15 13 9 1 1 9 9 0 2 1 9 15 1 9 9 9 2
20 13 7 9 0 1 7 8 1 9 1 9 7 9 1 9 1 9 9 15 2
10 9 9 9 1 9 0 8 1 9 9
86 8 12 2 12 2 8 8 2 2 9 2 0 2 9 2 0 2 13 9 0 0 1 9 0 8 8 7 9 0 14 13 0 1 9 1 9 9 0 1 9 1 9 8 9 7 13 9 7 9 0 1 9 9 0 2 7 13 7 2 9 2 8 2 8 13 9 9 15 1 9 9 7 9 1 0 7 15 13 7 15 0 1 9 9 2 2
56 9 2 9 2 13 9 9 0 8 8 9 1 9 1 9 1 9 9 1 9 2 7 13 2 7 9 13 8 8 9 0 9 2 8 1 7 13 9 1 9 9 7 1 7 13 9 9 13 8 8 9 0 1 9 2 2
37 7 13 9 9 0 1 9 8 11 8 1 9 15 1 9 1 9 9 0 1 9 1 9 9 2 9 7 9 9 2 9 13 1 9 9 0 2
63 9 2 8 2 9 2 0 2 13 9 9 0 8 8 1 9 9 1 9 9 7 9 0 0 8 8 7 15 13 1 9 9 9 15 2 3 1 1 9 2 1 9 2 7 13 7 2 9 13 1 9 8 0 7 15 13 1 9 9 9 15 2 2
62 9 2 9 2 13 9 0 1 9 9 7 9 9 0 2 0 0 1 9 9 2 1 0 9 7 9 13 1 9 9 9 0 2 7 13 9 1 9 1 2 9 9 1 9 1 10 9 7 14 7 14 9 14 13 1 9 0 13 1 9 2 2
102 9 2 9 2 0 2 9 2 13 9 0 7 9 9 9 0 13 12 12 9 2 7 1 9 0 1 12 12 9 0 2 1 9 9 1 9 2 9 1 9 2 1 9 12 2 1 9 15 2 13 9 9 0 8 8 8 7 9 13 0 1 12 12 9 1 9 9 0 1 15 1 9 2 9 12 2 7 13 2 1 9 13 2 9 2 9 15 13 1 9 9 1 9 12 12 9 1 9 7 9 2 2
50 9 2 8 2 8 2 13 9 9 0 1 9 9 9 9 0 1 9 2 8 2 1 8 1 9 1 12 1 12 9 2 9 0 7 13 9 0 0 0 13 1 9 9 9 0 8 8 1 9 2
45 7 13 9 7 15 13 9 9 9 15 13 0 9 1 12 1 12 9 2 9 9 1 9 8 7 13 1 9 15 8 8 9 9 9 0 1 9 15 1 12 1 9 9 15 2
72 8 2 8 2 13 9 0 0 2 8 8 2 9 9 9 8 9 2 8 8 9 1 9 1 9 9 0 1 9 1 8 7 8 2 7 13 9 0 1 9 2 8 8 2 8 8 7 10 9 13 7 9 9 0 0 7 0 13 1 9 9 8 9 1 9 8 9 1 9 9 8 2
97 9 2 9 2 13 9 0 8 8 7 15 13 9 1 12 12 9 13 15 2 9 0 2 1 9 9 0 1 9 2 7 13 2 7 9 0 13 1 9 12 12 9 9 1 9 9 1 9 2 8 8 8 2 7 10 9 13 9 0 0 1 9 2 7 10 9 15 9 9 0 1 9 15 13 8 8 2 2 7 13 2 3 9 9 0 1 9 1 9 9 8 13 13 9 15 2 2
101 9 2 9 2 13 9 9 0 8 8 8 9 1 9 1 9 1 9 9 7 1 9 1 9 9 15 1 9 0 1 10 9 0 1 9 2 7 13 1 9 1 9 9 9 7 9 14 13 9 14 13 1 9 0 8 8 1 7 15 14 13 2 9 0 2 1 9 13 9 15 2 7 13 2 7 9 9 14 13 7 13 1 9 2 0 7 1 0 1 9 0 7 12 9 9 2 1 9 9 2 2
7 9 1 9 8 9 1 9
46 8 2 8 2 12 2 12 2 8 8 2 2 13 9 0 9 0 7 9 1 9 0 1 9 8 2 9 8 2 13 9 9 0 9 9 1 9 15 8 0 0 1 12 9 9 2
39 7 13 8 8 1 9 1 9 9 7 15 14 13 0 1 7 9 8 8 14 13 1 9 15 7 13 12 1 9 14 12 2 9 1 9 9 2 9 2
30 7 13 7 15 14 13 1 9 2 7 13 9 0 2 1 9 14 13 1 9 1 9 9 1 12 9 2 9 0 2
48 7 1 9 10 9 2 13 8 1 9 0 2 7 15 9 0 13 9 0 1 9 8 2 0 1 9 8 8 1 9 2 7 13 7 10 9 2 13 9 5 8 5 2 9 9 8 8 2
48 7 13 8 7 15 14 13 1 9 8 1 9 0 13 15 9 0 8 8 1 9 1 9 1 2 9 2 9 0 9 1 15 1 15 9 0 12 15 13 9 0 7 13 13 1 9 9 2
14 7 13 9 0 1 9 1 9 0 1 9 7 9 2
12 9 9 8 1 8 1 9 9 0 1 9 15
34 8 12 2 12 2 8 8 2 2 13 9 0 9 9 7 9 9 0 8 8 1 8 14 13 9 9 1 9 9 0 1 9 15 2
33 7 13 9 0 8 8 1 9 8 8 7 9 13 2 9 1 9 9 2 9 15 13 14 13 8 1 8 8 1 8 1 8 2
17 7 13 9 8 0 1 9 12 1 9 0 2 12 8 8 2 2
22 7 13 9 9 15 7 9 0 14 13 9 15 1 8 1 7 13 9 9 1 9 2
16 7 1 9 0 2 13 8 14 13 9 9 9 8 8 8 2
33 7 1 9 9 8 8 0 0 1 12 9 2 9 0 13 8 1 9 12 9 9 1 9 1 9 1 9 9 0 1 9 0 2
33 7 13 9 9 0 8 8 9 0 7 8 2 0 9 0 1 9 2 13 1 7 13 9 7 9 1 9 1 9 9 0 0 2
21 7 13 2 8 7 13 9 9 9 0 7 1 0 7 8 1 15 8 8 2 2
6 9 8 13 9 1 8
37 8 12 2 12 2 8 8 2 2 13 9 9 9 9 8 11 8 8 9 9 1 8 9 7 9 0 13 8 8 12 12 9 13 15 9 0 2
15 7 13 12 1 9 9 9 9 15 13 1 12 12 0 2
30 7 13 1 9 9 1 9 0 9 0 1 9 0 1 9 8 8 8 15 13 3 1 8 7 13 1 9 1 9 2
21 7 13 9 12 12 9 1 9 1 9 1 15 12 12 1 9 0 1 9 15 2
13 9 9 1 2 0 9 2 1 9 9 7 9 15
39 9 12 2 12 2 8 8 2 2 13 9 0 9 9 7 9 13 9 9 0 1 9 15 13 1 9 0 1 9 1 9 9 7 9 15 1 10 9 2
47 7 13 9 2 9 2 1 9 9 9 8 2 9 2 1 9 9 8 8 9 15 7 9 13 7 9 2 9 2 15 13 15 13 9 9 0 1 9 9 1 11 9 1 9 9 0 2
34 7 13 9 9 8 8 8 8 13 9 9 9 0 0 1 9 8 8 2 9 0 1 9 9 8 8 8 2 1 9 1 10 9 2
23 7 13 8 7 2 0 1 9 2 14 13 9 15 13 7 2 14 13 9 15 9 2 2
61 1 9 0 2 13 9 0 1 9 2 12 8 9 9 2 9 9 8 0 1 9 9 15 13 1 7 15 13 1 9 1 9 9 0 7 9 9 9 7 13 1 9 9 13 8 8 8 8 2 12 9 2 7 9 0 1 12 9 1 9 2
32 7 13 9 9 0 1 9 0 1 9 9 15 9 1 9 0 1 9 9 1 9 1 9 7 9 9 1 9 1 9 0 2
45 7 13 8 1 9 1 9 2 8 2 13 15 9 7 9 9 13 2 9 1 9 2 0 1 9 0 0 1 9 13 9 2 9 9 0 7 9 9 7 9 9 7 9 2 2
14 7 13 2 8 7 13 9 1 9 0 1 9 2 2
11 9 9 0 1 9 9 0 12 12 9 0
36 8 12 2 12 2 8 8 2 2 13 9 0 1 9 9 0 15 13 9 9 1 7 9 9 0 1 9 0 8 8 13 12 12 9 0 2
25 7 13 8 9 9 15 9 15 13 1 0 15 0 8 8 15 13 9 15 1 9 2 9 0 2
36 7 13 9 9 0 1 7 9 8 15 13 13 9 0 1 9 7 9 9 13 1 12 12 9 1 9 0 7 12 12 1 9 9 7 9 2
47 7 14 13 9 9 9 9 0 15 13 1 8 9 1 15 1 9 1 9 0 2 7 13 9 1 9 9 1 9 9 8 8 7 15 14 13 15 7 13 13 1 8 9 9 1 8 2
49 7 13 9 1 9 15 7 9 9 1 15 2 14 13 1 9 1 9 0 13 15 9 9 1 9 1 9 0 2 2 0 7 10 9 2 14 13 0 7 14 13 0 1 9 9 0 0 2 2
31 7 13 9 1 7 15 13 9 1 10 9 7 13 1 9 15 0 9 0 1 9 9 1 15 1 9 9 9 1 9 2
9 9 0 1 8 8 8 9 1 8
51 8 2 9 0 2 12 2 12 2 8 8 2 2 13 9 0 7 1 9 0 7 9 9 0 8 8 7 9 15 0 8 8 14 13 1 9 0 9 9 9 2 1 9 0 2 1 9 9 1 9 2
29 7 13 9 9 15 7 9 14 13 1 9 0 2 12 5 12 2 1 9 0 1 9 9 1 9 0 7 8 2
19 7 13 9 0 7 9 14 13 0 1 9 9 0 7 0 1 12 9 2
19 7 14 13 9 0 9 1 9 1 12 1 9 9 1 9 0 1 9 2
23 7 13 9 1 8 9 0 1 9 14 3 0 7 9 0 15 0 1 9 9 0 0 2
18 14 7 9 13 8 8 0 7 0 1 9 9 0 8 8 1 12 2
27 7 1 0 7 13 9 0 1 9 0 8 8 9 1 9 15 14 13 1 9 0 1 9 0 1 9 2
46 7 13 9 0 8 8 9 0 9 15 13 15 8 1 9 0 2 1 15 13 15 9 9 1 9 2 7 13 8 0 1 9 15 13 15 8 1 2 9 1 9 2 9 9 9 2
35 14 7 8 13 1 9 9 0 1 8 7 13 9 0 9 1 9 15 1 9 12 15 13 1 9 8 1 9 1 9 1 9 9 0 2
13 8 9 0 1 9 9 9 0 1 9 0 7 0
36 8 12 2 12 2 8 8 2 2 13 9 0 8 8 9 9 1 9 0 9 1 9 9 0 1 9 0 1 9 0 1 9 9 9 0 2
34 7 13 8 9 1 9 13 15 9 1 9 9 9 2 9 1 9 0 7 0 15 14 2 0 1 7 15 13 1 9 9 9 0 2
39 7 13 7 9 15 13 15 9 9 0 1 9 8 12 12 9 0 7 9 15 13 1 10 9 2 13 0 1 9 1 9 1 9 1 9 2 9 0 2
37 7 13 9 0 7 15 2 13 9 9 0 2 7 13 7 15 2 14 13 9 9 15 1 9 1 9 0 1 9 0 1 9 1 9 0 2 2
59 7 13 8 8 1 9 1 9 9 0 0 1 9 0 2 9 2 9 9 0 1 9 1 9 9 9 2 1 9 0 1 9 7 1 9 9 0 13 1 9 1 9 9 7 9 9 0 1 9 15 13 15 1 9 9 1 1 9 2
13 8 2 2 14 8 8 2 1 9 9 1 9 0
49 8 12 2 12 2 8 8 2 2 13 9 0 8 8 9 9 1 0 1 9 1 9 9 1 9 0 0 1 9 2 9 9 0 2 1 9 15 13 0 1 9 0 7 9 7 9 1 8 2
46 7 13 8 1 9 2 8 8 9 2 9 13 1 9 7 14 8 8 14 7 8 13 9 1 9 7 9 7 15 13 1 7 1 15 0 1 9 8 13 8 8 15 8 8 2 2
40 7 13 8 1 9 1 9 0 1 9 9 0 8 8 8 2 2 13 7 13 1 9 15 0 1 9 7 1 7 15 14 13 0 9 1 9 7 9 2 2
16 8 2 9 2 9 2 9 0 14 13 1 2 9 2 9 0
42 8 2 8 2 12 2 12 2 8 8 2 2 13 9 9 0 9 1 9 8 8 9 9 1 7 9 2 9 2 9 0 1 9 14 13 1 2 9 2 9 0 2
39 7 13 8 0 1 9 1 9 1 9 9 1 9 1 8 2 8 2 1 9 9 0 0 1 9 9 8 8 2 8 8 1 9 1 9 8 8 2 2
47 7 13 9 1 9 8 8 1 8 9 9 9 1 9 7 8 13 7 15 14 13 9 1 9 8 0 1 12 9 2 9 0 2 1 9 9 9 1 9 0 7 9 13 15 9 2 2
46 7 1 1 13 8 0 1 9 9 13 9 9 0 1 9 8 8 9 9 9 1 9 1 12 9 1 9 8 8 2 1 9 1 12 8 9 8 2 13 9 15 9 9 1 9 2
11 9 8 0 9 1 9 9 15 8 1 8
36 8 12 2 12 2 8 8 8 2 2 13 9 8 8 0 0 9 8 8 0 9 1 9 9 15 8 8 1 9 9 9 9 1 8 0 2
19 7 13 9 9 0 3 9 8 0 8 8 7 9 9 8 0 8 8 2
42 7 13 8 9 8 1 8 8 0 3 9 1 9 9 0 1 9 9 9 0 2 12 2 9 2 1 9 0 1 9 9 0 7 13 9 0 1 9 15 8 8 2
37 7 13 8 9 1 9 8 9 9 0 13 15 1 15 1 9 1 8 2 7 7 15 13 1 0 7 13 9 0 1 9 1 15 9 9 9 2
67 7 13 8 1 9 0 1 8 8 8 1 9 9 15 1 9 7 13 0 2 8 12 9 8 1 9 9 2 8 7 8 15 15 9 15 0 1 9 1 8 8 7 9 15 0 2 2 7 13 2 7 15 13 1 9 0 2 8 8 1 7 8 1 9 0 2 2
61 7 13 8 2 9 8 0 0 2 13 9 15 1 9 9 1 9 8 7 13 1 15 1 9 9 9 0 1 8 7 13 1 0 2 7 13 1 8 2 13 8 2 1 9 9 2 7 13 1 9 15 9 8 0 0 8 8 1 9 9 2
77 7 13 8 1 15 1 9 8 9 12 1 7 13 1 8 1 9 1 8 1 9 12 9 7 13 1 15 1 9 0 7 13 15 1 9 1 9 9 2 7 13 15 7 13 1 8 8 15 13 13 1 9 0 1 9 1 9 0 0 1 9 0 15 13 1 15 1 7 13 1 9 0 1 9 9 0 2
17 7 13 8 1 1 9 1 7 13 9 0 1 9 2 9 0 2
1 9
13 13 9 7 9 0 1 15 1 9 9 1 15 2
18 13 9 0 1 9 7 1 15 7 1 9 15 2 7 9 1 15 2
13 1 9 9 2 13 15 9 1 0 1 9 0 2
9 9 15 1 9 1 9 7 9 2
9 0 9 15 10 9 15 9 9 2
1 9
19 14 14 13 9 1 9 0 7 13 15 1 9 1 9 0 1 9 9 2
10 9 15 0 0 1 9 7 9 9 2
8 15 1 9 1 9 7 9 2
11 9 1 0 9 1 15 9 0 9 9 2
9 0 9 15 10 9 15 9 9 2
1 9
11 13 9 7 9 7 9 1 9 7 9 2
6 13 9 1 9 15 2
9 13 0 7 14 13 1 9 0 2
8 13 9 1 9 0 7 0 2
9 0 9 15 10 9 15 9 9 2
1 9
10 14 13 1 9 0 1 9 9 15 2
17 9 15 14 13 15 1 9 1 9 14 13 1 9 1 9 15 2
17 14 13 9 10 13 1 15 1 9 9 1 15 13 15 10 9 2
8 9 0 7 13 1 9 15 2
9 0 9 15 10 9 15 9 9 2
1 9
12 13 7 14 13 1 9 15 1 9 10 9 2
11 14 13 9 15 0 13 7 13 1 15 2
13 8 9 1 9 15 7 13 0 9 1 9 9 2
16 13 7 13 8 8 1 15 7 13 9 7 13 15 1 15 2
9 0 9 15 10 9 15 9 9 2
1 9
9 13 1 15 1 15 1 9 9 2
20 13 15 9 9 9 0 1 9 10 9 7 13 1 15 9 0 1 9 15 2
15 9 15 1 9 0 14 13 1 9 15 7 14 13 9 2
11 9 0 1 9 13 7 13 0 1 9 2
9 0 9 15 10 9 15 9 9 2
1 9
12 13 15 9 9 1 1 9 9 1 9 15 2
16 9 15 1 9 9 9 0 14 13 15 1 9 1 9 0 2
17 14 13 9 0 15 14 13 15 0 9 1 9 15 13 1 15 2
15 13 15 9 9 0 1 9 15 7 9 15 7 9 15 2
9 0 9 15 10 9 15 9 9 2
1 9
13 13 9 7 9 0 1 15 1 9 9 1 15 2
18 13 9 0 1 9 7 1 15 7 1 9 15 2 7 9 1 15 2
13 1 9 9 2 13 15 9 1 0 1 9 0 2
9 9 15 1 9 1 9 7 9 2
9 0 9 15 10 9 15 9 9 2
1 9
32 14 14 13 9 15 1 9 9 9 15 0 8 8 1 7 13 15 1 9 1 10 7 14 15 14 13 8 1 9 8 8 2
8 9 15 13 9 10 1 15 2
16 15 1 9 1 9 1 9 9 7 13 9 15 0 1 9 2
5 13 0 1 9 2
9 0 9 15 10 9 15 9 9 2
1 9
8 14 14 13 9 9 1 0 2
11 1 15 1 9 0 1 10 13 1 15 2
25 14 15 9 0 9 1 9 15 7 9 13 8 9 7 13 9 1 9 15 7 9 15 1 0 2
10 14 13 0 1 15 13 15 1 9 2
9 0 9 15 10 9 15 9 9 2
1 9
9 13 9 9 1 9 1 9 0 2
8 14 13 9 1 9 1 0 2
11 14 13 9 15 0 7 13 9 15 0 2
14 13 9 0 7 13 1 9 0 1 9 1 9 9 2
9 0 9 15 10 9 15 9 9 2
1 9
23 9 15 15 13 15 1 15 9 9 15 0 1 15 9 14 13 9 0 1 9 1 15 2
16 9 9 15 9 7 9 9 14 13 1 9 15 1 9 0 2
12 13 1 9 0 0 1 1 9 15 1 9 2
15 13 9 1 0 9 1 9 9 1 1 9 1 9 9 2
9 0 9 15 10 9 15 9 9 2
1 9
7 9 1 9 14 13 9 2
11 14 13 7 7 13 7 13 9 15 0 2
6 13 1 9 9 0 2
13 14 13 1 9 0 1 9 15 1 9 9 0 2
9 0 9 15 10 9 15 9 9 2
13 1 9 13 9 0 2 7 13 1 9 15 1 9
10 12 0 1 9 9 7 9 1 12 9
37 13 9 9 9 0 1 9 0 8 8 1 9 9 0 9 13 1 15 2 0 2 0 1 12 9 13 1 15 9 9 7 14 13 1 9 9 2
33 9 9 13 7 9 0 13 1 9 9 13 1 15 9 0 1 9 9 0 8 8 9 9 0 1 9 0 2 9 1 9 0 2
56 7 13 9 1 9 7 13 1 9 0 1 9 9 15 0 7 13 1 7 15 13 13 1 9 1 8 8 9 8 0 1 9 9 8 1 9 9 7 13 1 9 13 1 9 15 9 0 7 13 1 9 15 1 9 0 2
52 7 1 7 13 1 9 0 1 15 13 9 9 0 0 7 13 1 15 9 7 13 1 15 9 9 7 9 9 0 1 15 13 1 9 0 1 9 9 0 1 9 1 9 9 0 1 7 13 9 1 15 2
43 7 9 1 10 9 13 9 9 9 0 8 8 1 9 9 7 13 1 9 1 7 13 1 9 9 0 1 9 15 1 10 13 9 1 9 13 15 9 0 1 15 0 2
34 7 9 1 15 13 0 9 0 1 9 1 9 9 9 0 9 1 9 15 0 9 9 0 1 9 0 8 8 1 9 9 1 9 2
52 7 13 1 9 9 13 15 1 9 1 9 0 1 15 7 14 13 9 0 12 7 13 9 1 15 13 1 15 7 13 9 12 1 15 9 15 13 1 15 7 1 0 7 13 1 0 9 1 9 9 0 2
2 8 8
6 1 9 9 9 0 2
7 9 0 1 9 0 1 9
27 9 2 9 9 2 13 9 1 9 9 0 0 1 9 9 9 15 1 9 1 9 9 9 0 1 9 2
43 7 13 9 9 9 0 1 9 8 15 13 12 9 1 9 1 9 9 7 12 0 1 9 9 0 0 13 9 15 1 9 9 9 9 0 1 9 15 7 15 13 15 2
48 7 13 9 9 9 9 9 15 7 15 13 15 0 9 15 7 13 13 1 9 2 1 9 1 9 1 9 9 9 7 1 9 1 9 9 0 15 14 13 15 1 0 9 1 9 9 15 2
24 7 13 9 13 13 15 9 15 1 9 7 9 0 14 13 15 1 9 9 15 1 10 9 2
11 7 14 13 9 9 0 9 7 13 15 2
49 7 13 9 0 1 10 13 9 15 9 0 9 9 9 9 1 9 1 9 9 15 1 15 7 9 15 1 9 9 0 1 9 9 7 13 1 9 9 0 1 9 7 9 0 0 1 9 9 2
69 7 13 9 8 7 9 9 9 9 0 7 15 13 1 9 1 9 8 9 9 9 0 0 0 1 9 0 1 9 0 7 1 9 0 13 13 15 12 1 9 0 9 9 0 0 1 10 9 15 13 9 0 7 9 13 1 15 1 9 9 15 0 7 0 15 15 13 9 2
1 0
12 12 9 9 12 9 1 9 0 1 9 9 9
15 9 2 9 1 9 0 0 1 9 9 9 7 9 15 2
75 13 9 9 9 9 9 0 1 9 9 1 9 9 9 9 9 9 1 9 1 9 13 1 15 9 9 12 9 7 14 13 9 1 9 9 0 1 10 9 1 9 0 13 9 15 1 12 9 1 9 15 1 9 7 9 0 1 9 9 1 10 9 7 10 9 0 1 9 9 0 1 9 1 9 2
7 9 9 1 9 0 1 9
50 7 1 9 9 3 13 9 9 9 9 9 1 9 9 0 1 9 1 9 9 9 9 1 9 1 9 0 1 10 9 7 14 13 9 0 1 9 9 1 9 9 1 13 9 9 1 9 1 15 2
5 9 1 9 9 0
42 7 13 9 0 1 9 1 9 9 9 0 7 1 10 9 13 9 9 1 9 1 9 9 9 13 1 15 9 9 9 0 13 1 9 9 12 1 9 9 9 0 2
35 7 13 7 9 0 1 9 9 9 3 1 9 1 9 9 7 9 1 9 1 9 9 7 15 9 1 9 0 1 9 1 9 7 9 2
2 8 8
4 9 9 0 2
8 9 0 13 1 9 9 1 8
40 8 8 2 9 9 2 13 9 9 7 9 0 1 9 9 0 1 9 9 13 9 1 9 9 1 9 9 14 13 1 9 9 15 13 15 9 9 8 8 2
39 7 13 9 13 3 7 15 13 9 0 1 9 13 9 9 0 9 1 9 1 9 9 0 14 1 0 9 1 9 9 9 9 0 8 8 7 9 15 2
48 7 14 13 9 0 0 1 9 8 7 9 9 15 8 8 1 9 0 7 9 1 9 0 2 7 13 9 8 1 9 9 1 9 15 7 9 9 13 1 9 9 1 9 9 7 9 9 2
34 7 13 9 1 9 9 9 9 1 9 9 8 2 1 1 15 9 8 8 9 9 0 1 9 0 2 8 8 8 8 9 9 0 2
51 7 13 9 0 7 8 13 1 9 0 9 9 0 1 9 8 7 9 9 9 0 2 8 8 9 1 9 8 1 9 9 0 1 9 2 7 0 10 8 13 1 9 1 9 9 7 9 1 9 0 2
42 7 9 9 9 0 1 9 9 8 1 9 9 2 14 7 15 13 1 9 9 9 9 9 0 1 9 0 15 14 13 1 9 9 9 0 1 9 8 8 8 8 2
29 7 13 8 13 1 9 9 0 1 9 9 0 2 8 12 9 1 9 1 9 15 2 7 15 14 13 10 9 2
17 7 13 9 0 7 8 13 1 9 0 1 9 9 1 9 15 2
21 7 13 10 9 9 0 1 9 9 0 7 8 2 7 9 0 1 9 15 9 2
36 7 13 8 8 9 9 9 0 1 9 15 1 9 1 9 9 7 9 9 13 9 15 1 9 13 1 9 2 7 0 13 1 9 9 15 2
29 7 13 9 8 1 9 8 1 9 9 1 9 7 14 13 9 1 9 15 1 9 13 15 14 12 1 9 0 2
29 7 13 9 0 9 9 0 8 9 9 7 9 0 14 13 0 1 9 9 9 1 9 0 7 0 7 0 9 2
3 1 9 0
8 9 1 12 9 9 0 1 9
47 13 9 0 0 1 9 0 1 9 0 1 9 7 9 0 1 9 9 9 9 9 1 9 0 7 13 9 15 9 1 12 9 0 9 0 13 1 9 15 1 2 8 2 1 9 0 2
44 8 8 7 9 9 13 9 1 10 9 0 9 0 1 9 9 0 8 1 7 13 0 1 9 9 0 1 9 0 8 8 1 9 9 7 9 9 0 1 10 9 1 15 2
40 7 13 9 0 7 9 0 1 9 9 13 1 9 9 9 9 7 9 9 0 0 0 1 9 9 15 7 13 9 2 8 2 8 0 1 9 1 9 0 2
64 7 13 9 1 15 7 13 9 1 9 1 9 15 1 9 8 7 1 9 9 1 15 1 9 9 9 9 0 1 9 0 8 8 13 0 1 15 15 13 9 15 1 14 12 9 7 14 12 9 7 15 13 1 9 0 1 9 9 8 8 8 8 8 2
41 7 13 7 15 13 1 9 9 9 9 1 9 15 7 13 15 9 12 1 15 12 9 7 13 1 9 0 1 9 9 1 7 13 9 7 13 1 15 9 0 2
3 8 2 8
2 1 9
7 13 9 9 7 13 1 9
41 13 9 9 1 9 9 0 1 9 9 0 1 9 9 13 1 9 1 12 9 13 9 15 1 9 9 1 1 9 0 7 13 0 0 1 7 15 13 9 0 2
38 7 14 0 1 10 9 7 15 7 7 8 9 0 7 1 15 0 13 1 9 1 9 7 13 1 15 7 13 0 1 9 1 13 9 15 12 9 2
76 7 14 1 9 9 7 14 9 0 7 0 1 15 13 1 7 0 13 13 1 9 9 0 7 13 1 15 7 13 9 15 7 1 9 9 9 15 13 15 7 15 13 13 1 9 1 9 14 1 9 9 9 15 1 9 7 13 1 7 9 0 7 13 1 9 1 9 7 13 1 15 13 15 9 15 2
73 0 9 13 1 9 0 1 9 9 13 9 9 15 0 7 13 9 7 15 15 13 1 15 0 7 13 1 9 7 13 1 0 7 1 9 9 7 13 1 9 9 7 9 15 0 13 15 1 9 9 15 13 15 1 9 9 15 1 9 9 15 7 13 15 1 9 7 15 13 13 1 9 2
49 7 1 9 13 8 1 9 7 13 9 9 7 13 1 9 9 15 13 9 15 1 9 9 1 9 9 1 15 7 14 13 1 15 13 1 15 7 13 9 15 1 9 1 9 9 1 9 15 2
7 9 9 13 14 12 9 2
15 9 9 0 1 9 2 7 9 8 1 9 1 9 1 9
57 8 2 8 8 2 13 9 0 3 9 15 1 9 9 7 13 12 1 15 1 12 9 13 8 13 9 9 0 7 15 13 1 9 15 2 0 2 1 9 0 8 8 8 2 1 1 13 9 9 1 9 1 13 1 9 9 2
31 7 1 9 13 9 0 9 9 7 9 12 0 1 9 1 9 15 13 15 9 9 3 1 9 0 1 9 1 9 9 2
18 7 13 9 9 0 1 9 9 0 2 1 15 9 7 12 9 2 2
17 7 13 9 9 1 9 7 2 9 0 2 1 0 13 1 9 2
35 7 13 7 9 7 15 0 1 9 15 1 12 9 13 9 0 1 9 0 7 13 1 9 9 1 9 15 13 1 9 9 1 1 15 2
16 7 13 9 1 2 7 9 0 1 9 0 13 7 13 2 2
40 7 13 9 9 7 12 7 12 9 13 1 9 15 8 8 15 13 9 0 13 0 1 9 1 9 9 1 9 12 1 9 0 3 7 15 14 13 9 9 2
38 7 14 13 9 0 3 9 0 1 8 9 13 9 0 7 15 13 15 1 12 7 12 9 13 7 7 13 7 15 13 13 9 9 9 0 1 15 2
5 1 0 9 7 9
24 7 1 9 15 13 9 0 1 9 8 0 9 7 12 0 0 13 9 3 1 9 9 0 2
37 7 14 13 1 9 0 0 9 1 10 9 15 13 9 0 7 15 13 1 9 9 9 2 15 13 1 0 9 1 9 1 9 0 7 9 0 2
21 7 13 9 0 7 0 7 15 13 1 9 9 9 8 0 1 9 0 8 8 2
50 7 1 9 9 13 9 0 1 9 9 15 13 9 1 9 0 1 9 0 7 9 2 7 13 9 0 7 0 14 13 7 10 9 13 9 9 9 7 9 1 9 9 0 15 13 1 15 0 0 2
28 7 13 9 0 7 0 9 9 2 7 13 9 9 7 9 1 9 0 0 1 9 9 9 9 9 1 9 2
46 7 13 9 9 1 9 0 15 13 1 15 9 9 0 15 13 1 9 9 0 7 15 13 9 0 7 9 15 13 0 1 12 9 2 1 15 12 5 1 0 2 7 1 12 9 2
32 7 13 9 1 9 9 0 1 9 9 1 9 1 7 15 0 2 7 13 2 1 9 9 7 9 13 9 1 9 9 2 2
8 13 8 7 9 7 8 8 8
8 9 0 1 8 1 8 9 0
44 8 2 7 1 2 2 13 9 1 9 9 0 8 8 8 3 7 9 0 13 8 7 9 7 8 7 8 1 8 2 9 9 2 14 13 1 8 2 1 12 9 8 2 2
44 7 13 8 8 7 2 9 0 1 8 14 13 1 9 8 8 13 9 9 0 2 7 14 13 2 9 7 9 0 15 1 15 9 1 10 9 7 9 7 8 7 8 2 2
22 7 13 7 9 0 1 9 9 1 10 9 15 2 14 13 1 12 9 1 8 2 2
39 7 13 9 0 13 1 9 9 1 9 0 8 8 7 9 9 9 0 9 8 8 8 8 8 8 9 9 9 9 8 8 7 15 9 9 0 9 0 2
25 7 13 8 1 12 9 9 0 7 9 0 0 13 1 12 12 9 7 1 12 12 9 1 8 2
37 1 9 0 2 13 9 0 8 8 13 3 9 7 15 14 13 15 7 13 9 9 15 7 7 15 0 1 9 1 9 2 9 7 4 9 2 2
69 7 1 8 13 15 1 9 9 0 0 13 9 8 14 15 2 0 1 9 1 9 9 2 1 9 2 9 7 4 9 2 8 8 1 9 1 9 9 9 0 1 9 9 8 8 9 9 1 9 1 9 1 9 9 1 9 9 9 9 1 9 0 9 1 9 9 15 0 2
25 7 13 9 9 15 13 0 7 13 1 9 7 9 1 9 9 9 1 9 7 9 0 1 9 2
22 7 13 8 7 15 2 13 1 9 9 0 1 9 7 14 8 9 0 9 0 2 2
43 7 13 2 13 1 15 0 9 1 9 7 15 9 9 0 2 14 3 7 2 9 1 9 9 0 1 9 7 15 1 9 9 0 1 9 7 7 13 9 9 0 2 2
49 7 13 7 2 9 9 13 9 9 2 1 1 7 13 1 15 9 7 15 2 14 13 7 8 9 1 9 9 1 9 2 0 0 0 7 9 15 1 9 2 7 9 15 15 13 9 9 2 2
41 8 8 13 8 7 2 0 1 9 0 1 8 14 8 1 15 7 9 9 1 15 9 0 1 9 9 0 2 0 0 7 2 9 10 13 0 1 9 0 2 2
2 8 9
39 9 0 2 13 9 8 8 9 0 7 9 0 1 9 0 12 1 9 9 9 9 0 1 9 9 1 9 1 9 0 7 0 0 1 9 12 9 8 2
4 1 9 0 2
40 13 9 9 0 1 9 0 7 0 9 0 1 9 9 0 1 9 2 7 13 9 9 13 9 0 13 15 9 1 0 9 2 7 13 1 9 15 9 0 2
20 7 1 0 7 13 8 9 1 9 9 9 14 13 9 15 7 9 15 0 2
4 9 1 9 2
24 8 7 9 0 1 9 13 9 1 9 9 1 9 9 14 13 9 15 1 0 1 9 0 2
24 7 14 13 10 9 9 9 0 1 9 9 1 9 9 15 1 9 9 9 0 9 9 0 2
3 9 0 2
34 13 9 0 1 8 9 0 0 1 15 1 9 0 2 7 15 9 13 7 13 15 9 1 9 9 15 1 9 0 1 9 9 15 2
29 7 13 9 0 0 7 9 0 0 7 9 9 0 2 0 0 1 9 1 9 9 15 1 12 9 1 9 9 2
3 8 2 8
4 9 9 9 9
10 0 9 9 1 9 10 14 13 15 9
33 8 2 8 13 1 9 9 9 9 12 9 8 0 1 12 8 9 9 9 1 0 9 9 1 9 9 9 9 1 9 12 8 2
87 7 1 9 0 1 15 1 9 0 7 14 9 9 1 9 7 9 7 9 13 9 9 1 9 0 9 7 12 9 1 9 8 0 9 7 12 9 1 9 9 2 7 14 13 9 9 9 1 9 9 1 9 0 1 9 12 9 13 1 15 9 0 1 9 7 9 9 1 9 9 15 1 12 9 7 12 9 7 12 9 7 9 9 1 9 9 2
59 7 7 14 13 9 9 9 9 9 7 14 9 15 14 13 1 15 13 14 12 9 1 9 9 9 9 1 9 0 2 9 7 9 9 9 9 9 13 1 9 9 0 7 0 1 10 9 9 7 9 9 7 9 9 1 9 7 9 2
47 0 7 1 9 1 9 0 7 1 15 13 1 9 8 7 14 9 9 1 0 9 1 9 0 1 8 9 9 9 13 1 9 1 9 9 1 9 0 9 7 10 9 13 9 1 9 2
19 0 7 14 9 9 0 1 9 0 1 8 9 1 9 0 13 1 9 2
58 7 0 7 1 9 1 9 0 8 1 9 9 1 8 1 9 7 14 9 9 9 9 14 13 9 9 1 9 9 1 7 13 13 1 9 8 9 9 9 0 1 9 9 7 9 0 0 1 9 9 7 13 1 9 15 9 0 2
81 7 1 9 9 13 7 9 0 7 13 9 1 9 1 7 13 9 0 1 9 7 9 9 7 15 15 13 9 9 9 0 7 9 9 1 9 7 9 7 9 9 0 1 15 7 9 9 9 9 0 14 13 0 1 9 15 7 7 13 9 9 13 9 9 7 1 8 8 8 1 8 9 14 13 9 9 9 12 9 0 2
2 8 8
11 9 0 2 9 12 9 0 1 9 7 9
43 9 2 9 2 12 9 0 0 1 9 7 9 1 9 9 0 7 9 13 9 1 9 15 0 1 9 9 0 1 15 1 9 0 0 7 9 1 9 15 7 9 15 2
50 1 9 9 0 7 15 9 0 1 9 0 7 9 0 7 14 8 1 15 9 9 7 9 0 9 1 9 9 0 15 1 9 15 9 9 7 9 9 9 0 7 9 0 9 8 8 1 15 9 2
67 1 9 0 13 9 0 1 9 9 9 7 9 0 9 1 9 1 9 9 9 7 9 7 9 1 9 0 1 9 0 7 9 9 0 1 9 9 0 7 9 9 9 7 13 10 9 1 9 9 9 15 1 9 15 9 0 1 9 9 9 1 9 0 7 0 0 2
38 14 9 0 7 15 0 1 9 9 0 7 9 7 9 0 9 15 1 9 15 9 9 9 7 9 0 0 7 0 8 8 8 0 7 0 7 0 2
38 1 1 13 9 0 0 9 15 9 1 9 0 9 7 9 0 9 0 1 9 9 7 9 9 0 7 9 9 15 7 9 15 7 9 8 9 15 2
48 7 13 0 9 1 9 9 15 1 9 15 1 9 1 9 7 9 0 1 15 13 9 0 1 9 15 7 9 15 9 7 7 15 13 1 10 9 9 9 0 9 9 0 0 7 9 0 2
7 1 9 8 8 1 9 0
6 9 9 9 0 1 9
51 9 2 9 9 2 2 13 8 8 13 15 9 0 8 8 9 7 13 1 15 9 0 7 9 0 9 12 15 13 1 9 9 0 1 9 9 1 9 9 9 7 13 9 0 9 1 9 9 9 0 2
50 7 13 9 8 9 1 9 1 9 9 8 0 0 0 1 8 13 1 9 9 2 1 8 9 8 8 13 9 0 1 9 9 9 0 12 7 9 9 0 2 0 15 13 9 2 1 9 2 2 2
37 7 13 8 9 0 9 1 9 8 1 9 1 9 9 0 8 8 0 2 7 14 9 1 10 14 13 1 9 1 9 9 1 9 9 15 2 2
33 1 9 15 13 9 8 9 9 9 9 9 0 1 9 9 1 8 8 2 7 8 13 9 12 13 0 1 9 0 1 9 2 2
45 9 1 7 9 15 13 1 12 9 13 1 9 9 9 0 7 9 9 1 7 15 9 0 0 15 13 1 9 15 1 9 0 2 12 2 12 2 1 9 9 0 1 9 9 2
43 1 9 13 1 9 0 9 9 1 9 12 7 14 13 1 15 9 2 9 9 9 2 7 15 9 15 13 15 9 9 8 8 0 1 8 7 0 1 9 15 1 8 2
46 7 13 8 1 9 9 8 1 1 7 13 15 0 7 8 13 9 12 1 9 9 0 1 9 9 1 2 9 2 15 13 13 1 15 2 1 9 9 7 9 7 9 9 0 2 2
36 7 1 9 0 1 9 15 1 8 13 9 8 1 9 10 9 0 9 0 2 1 9 9 9 0 1 9 9 7 9 0 1 9 15 2 2
27 7 13 8 7 9 12 13 1 2 9 9 0 2 1 9 9 1 9 7 8 2 8 1 9 0 2 2
39 7 13 9 9 0 0 9 9 1 9 9 1 10 9 15 13 9 1 9 9 0 1 9 7 1 7 13 9 9 1 9 15 1 9 0 1 10 9 2
35 13 7 8 13 1 0 9 1 9 9 9 0 1 9 15 1 9 13 1 15 1 12 12 9 7 13 1 9 1 12 12 1 9 15 2
35 14 9 9 0 7 13 1 8 8 2 9 9 2 7 13 9 9 0 1 7 15 13 9 9 0 15 13 15 9 1 9 12 7 12 2
45 13 1 7 9 9 15 13 15 9 2 7 15 13 1 9 9 0 15 13 1 15 0 9 0 8 8 2 7 3 9 1 9 9 7 9 8 8 8 8 8 13 9 9 0 2
39 7 13 9 0 1 9 9 9 7 8 13 9 8 13 9 9 15 13 9 9 15 7 13 8 8 14 13 1 9 9 1 9 1 7 13 9 9 0 2
35 7 13 9 0 1 7 9 9 13 1 9 2 1 8 2 2 13 9 0 1 9 2 7 8 7 1 15 9 8 1 8 9 9 0 2
2 1 8
14 9 12 9 1 9 9 1 9 0 7 9 12 9 0
36 13 9 9 9 0 8 8 1 9 0 1 9 7 9 0 12 9 1 9 9 1 9 13 7 15 0 1 9 1 9 0 0 1 9 9 2
38 7 13 1 10 9 9 9 8 8 7 9 13 15 9 1 9 9 9 0 1 9 9 1 9 7 12 9 0 14 13 9 1 9 15 0 7 0 2
34 8 8 7 9 1 0 12 14 13 0 1 9 9 9 9 0 8 8 1 9 1 9 9 0 1 9 0 8 2 9 9 15 2 2
34 9 9 13 7 9 0 13 9 9 9 0 8 8 9 15 9 12 9 13 7 15 0 1 9 9 1 9 1 9 0 1 9 9 2
53 7 9 1 9 9 7 14 13 9 1 9 9 1 9 0 1 15 7 13 0 1 15 7 13 1 15 9 1 9 9 7 13 1 15 12 9 0 14 13 9 15 1 7 9 15 7 9 8 8 7 9 0 2
36 7 1 9 15 1 9 0 14 13 0 1 15 1 9 7 8 1 9 9 7 7 9 0 1 9 15 0 7 13 9 1 15 13 1 15 2
73 7 13 7 15 13 1 15 1 15 1 9 1 9 1 10 9 1 9 15 1 9 9 0 0 1 15 7 13 0 1 15 12 2 9 15 0 9 8 7 9 1 8 7 0 15 1 8 2 7 15 13 1 9 7 13 9 15 1 9 9 9 7 8 9 15 9 7 15 13 9 15 13 2
2 8 8
10 9 9 11 8 1 9 9 9 9 2
14 8 8 7 13 9 9 7 9 7 13 9 9 7 9
60 8 2 8 2 1 9 9 9 9 0 13 9 8 8 11 8 9 3 1 9 0 1 9 1 10 13 9 15 2 2 8 9 8 9 13 8 8 1 8 9 0 9 9 0 13 15 9 1 15 7 1 9 9 1 9 7 0 7 9 2
42 14 15 9 9 8 8 15 13 1 8 8 9 9 7 0 9 7 13 1 8 8 9 9 7 9 8 8 8 1 9 9 7 9 0 7 9 8 8 1 9 0 2
43 7 14 8 1 10 9 0 1 9 9 9 7 9 1 1 15 13 15 9 7 9 9 7 9 1 0 9 1 9 1 0 9 7 9 9 9 1 0 15 1 0 9 2
34 7 8 1 10 9 1 9 9 0 7 9 0 1 9 9 8 8 9 7 9 9 0 9 8 8 8 0 8 8 8 0 7 0 2
47 7 14 8 8 8 8 10 9 0 1 9 0 13 1 15 9 7 13 9 14 9 1 8 8 1 7 13 9 9 7 9 7 13 1 15 9 9 7 9 1 9 9 7 9 7 9 2
2 8 9
2 8 9
41 8 1 15 9 1 15 9 0 0 1 9 7 13 15 1 9 7 9 1 9 0 7 0 1 9 7 1 15 7 1 8 9 7 9 1 9 9 7 9 15 2
7 7 9 9 7 9 1 9
11 7 9 9 7 9 0 1 0 2 2 2
1 2
2 9 0
8 12 9 0 1 8 2 2 2
7 7 8 13 1 9 9 0
36 9 2 9 9 2 2 13 9 9 9 9 15 1 9 8 7 13 9 1 9 8 8 9 1 9 9 0 1 9 8 8 8 8 8 9 2
50 7 14 13 9 9 1 9 9 1 9 13 1 9 12 9 1 0 1 15 9 9 9 9 9 0 1 9 9 2 7 9 1 12 1 9 15 7 13 9 15 7 15 1 0 7 12 1 9 0 2
34 7 13 9 0 7 9 8 8 13 1 9 0 1 0 0 1 9 8 1 9 9 13 1 15 9 9 1 9 8 8 8 1 9 2
16 7 13 9 9 12 9 0 1 9 0 7 0 1 9 9 2
17 1 9 13 9 1 9 9 8 7 9 9 15 1 9 9 0 2
17 7 13 9 1 9 1 15 7 9 14 13 9 0 1 9 9 2
34 7 13 9 9 9 9 9 0 1 9 0 7 13 1 9 8 9 9 8 8 2 9 9 9 0 0 15 13 1 8 8 9 0 2
24 7 13 8 3 9 9 0 1 9 8 7 13 9 0 7 15 2 8 9 2 1 9 15 2
37 7 13 8 1 9 0 0 1 9 13 15 1 9 9 0 7 9 15 13 9 15 9 1 9 0 2 14 13 9 7 13 9 0 1 9 2 2
43 7 13 9 2 8 2 0 13 3 7 9 0 1 9 0 13 1 8 9 9 0 1 9 8 7 13 7 15 2 8 9 1 9 15 2 1 9 9 9 2 9 2 2
48 7 13 9 2 9 9 13 13 1 9 9 0 1 9 9 8 7 9 13 1 10 9 9 9 9 7 9 15 13 15 1 8 8 8 8 8 8 8 15 13 7 13 8 8 1 9 2 2
34 1 9 0 13 9 0 1 9 7 2 9 9 9 9 0 7 9 9 1 9 9 8 14 13 1 9 0 9 9 8 1 9 2 2
7 15 13 1 9 0 0 2
36 9 2 9 13 7 15 13 9 9 13 1 9 9 9 9 0 0 2 1 15 13 9 0 7 9 15 13 9 1 9 15 1 9 7 9 2
40 7 14 13 9 1 9 9 9 9 1 9 0 2 1 9 9 15 9 9 2 2 9 0 2 7 15 15 13 1 9 0 3 7 7 13 9 9 15 0 2
27 7 13 9 1 9 1 9 2 13 1 9 15 1 9 9 9 2 9 1 7 9 1 9 1 9 9 2
55 9 7 9 0 0 2 14 13 9 15 13 9 1 9 9 0 2 7 15 15 13 9 9 0 2 13 9 1 15 2 9 8 8 2 9 9 9 1 9 15 13 15 9 1 9 1 9 9 9 0 0 1 10 9 2
3 9 9 2
82 7 13 1 9 15 13 1 2 9 2 7 9 13 1 9 1 9 7 9 9 0 2 7 9 13 7 13 9 9 0 2 7 1 9 1 9 2 13 9 9 9 9 1 9 9 1 10 2 7 9 0 1 9 2 13 14 13 3 1 9 9 0 2 13 1 15 9 0 9 1 9 0 2 7 13 1 9 0 1 9 15 2
42 7 13 7 9 1 9 9 7 9 9 14 13 1 9 0 2 1 7 13 9 1 9 10 9 1 9 0 1 9 1 7 9 13 1 9 0 15 13 1 9 0 2
30 13 7 9 8 8 9 0 1 9 0 0 13 13 9 0 9 9 0 2 13 1 15 9 9 15 1 9 0 0 2
2 8 8
7 9 0 1 9 9 11 8
53 8 2 8 2 13 9 3 1 9 9 1 9 9 0 0 1 9 9 8 0 9 0 1 9 9 0 0 7 1 9 9 0 1 9 7 9 8 8 9 1 9 15 0 1 9 8 9 11 8 1 9 0 2
44 7 13 9 8 0 1 9 9 15 9 0 15 13 15 9 8 9 11 8 1 9 9 7 9 0 0 1 7 9 9 15 13 9 15 1 9 1 10 9 14 13 12 9 2
58 7 13 9 0 1 9 9 0 9 7 9 15 13 1 9 9 7 9 0 1 15 9 9 9 1 12 9 9 12 1 12 0 7 9 0 1 12 1 12 9 1 9 9 15 9 1 9 9 9 0 7 9 0 7 3 9 0 2
30 7 13 1 9 0 8 1 9 9 0 1 9 7 9 0 1 10 9 1 13 9 0 7 0 1 9 8 9 0 2
89 7 1 9 0 13 9 8 0 1 9 0 1 9 8 9 11 8 1 9 0 12 2 12 7 13 7 10 9 0 13 0 7 0 8 8 9 7 0 1 9 7 9 9 9 9 0 7 13 1 7 9 0 1 10 9 0 13 9 0 1 9 9 0 7 9 1 9 9 7 9 9 0 1 9 0 1 9 0 9 1 9 1 9 0 1 9 9 0 2
53 7 13 9 0 1 9 9 1 9 9 15 9 0 1 9 0 1 9 9 9 12 9 8 7 9 1 9 8 9 11 8 9 1 9 9 0 0 7 1 9 9 0 0 9 8 7 9 7 9 0 1 9 2
86 7 13 9 8 8 8 9 9 0 1 9 7 9 0 13 1 9 15 7 9 12 9 14 13 9 13 1 15 0 9 15 1 9 9 8 9 11 8 7 9 1 9 9 7 9 1 9 15 1 10 13 15 8 1 9 9 15 0 1 9 7 9 15 9 9 7 9 9 0 7 9 9 7 9 9 0 7 9 7 9 7 9 0 7 0 2
4 9 0 1 9
13 2 9 1 9 0 7 9 9 9 0 1 9 0
74 1 9 12 0 1 9 0 1 1 9 12 1 9 8 0 15 13 9 0 1 12 9 1 0 9 7 9 7 9 7 9 13 9 0 0 9 1 8 9 1 9 9 1 9 8 8 8 0 1 9 9 9 7 15 13 15 9 15 1 9 0 7 0 1 15 9 15 15 13 1 10 9 0 2
4 9 0 1 9
47 1 10 9 13 0 9 1 1 9 1 9 9 9 1 9 0 15 13 9 0 0 1 9 0 1 9 8 0 1 9 10 1 9 9 7 7 9 0 14 13 9 1 9 9 0 0 2
30 2 2 2 8 8 2 12 1 10 9 15 13 9 0 0 1 9 0 9 1 9 15 1 9 0 9 7 0 9 2
55 10 9 9 8 8 8 8 8 7 14 13 15 9 9 1 8 9 0 1 9 9 2 7 7 2 9 9 2 1 9 0 8 8 13 9 1 9 15 1 9 9 1 8 7 13 1 9 9 1 0 1 9 0 0 2
74 2 2 9 2 9 9 2 8 8 8 8 7 15 13 9 9 1 9 0 1 9 0 1 12 9 7 9 9 14 13 15 0 1 9 1 9 0 9 0 0 1 8 7 8 7 9 0 0 1 7 8 9 2 9 9 0 2 8 8 8 7 15 13 9 15 1 8 1 9 9 0 2 2 2
25 1 1 7 0 9 8 8 2 9 8 2 13 9 15 1 9 0 9 1 9 9 9 0 0 2
5 9 7 15 7 15
69 14 1 15 13 1 9 0 7 7 9 8 8 8 7 15 13 9 0 1 9 9 1 8 1 9 0 1 9 8 0 13 9 15 1 9 0 1 9 9 0 9 15 1 15 9 9 2 15 7 15 2 1 8 8 7 15 14 13 1 9 15 1 9 1 9 0 1 9 2
27 2 7 1 9 9 7 7 8 8 14 13 2 8 2 8 8 8 14 13 2 1 8 8 2 2 2 2
3 8 11 8
6 9 9 0 1 9 13
10 9 12 9 0 7 9 0 1 12 9
84 9 2 9 9 2 2 13 9 9 0 1 9 7 13 9 3 1 9 0 13 1 9 0 1 9 9 0 8 1 9 0 7 9 9 1 9 7 13 9 0 1 9 15 9 7 9 12 0 1 9 12 1 0 15 9 8 9 9 0 3 7 13 9 1 9 0 7 12 1 9 9 13 3 1 9 13 1 15 1 9 8 8 9 2
6 9 1 9 1 9 0
35 7 1 9 2 13 0 9 1 9 0 3 1 9 0 13 0 1 9 0 2 7 13 9 0 1 9 9 7 9 1 0 0 7 0 2
22 7 14 13 9 0 1 8 1 0 9 1 9 9 9 9 9 1 9 1 9 9 2
27 7 13 12 9 14 13 7 13 9 0 1 9 9 0 3 1 9 0 1 0 9 7 9 0 1 9 2
32 7 13 9 9 2 15 13 1 15 9 0 7 0 0 9 0 2 1 9 0 0 8 8 9 9 0 1 9 0 8 8 2
12 7 9 9 13 7 9 0 14 13 1 0 2
25 7 1 8 13 9 9 9 0 1 9 0 9 3 7 13 0 1 9 15 1 0 9 10 9 2
28 7 1 8 8 9 13 9 0 7 9 13 7 13 0 1 9 1 9 9 9 9 3 1 9 1 10 9 2
2 9 0
32 7 1 9 0 0 13 0 1 9 0 9 9 9 9 0 3 2 7 13 1 9 9 0 7 9 12 0 1 9 8 8 2
14 7 13 9 0 0 7 9 13 1 9 9 9 0 2
29 7 1 15 13 9 0 9 12 9 0 7 9 7 9 9 0 1 9 1 9 13 9 1 9 0 1 9 0 2
12 7 13 9 0 1 9 1 9 9 8 9 2
23 7 13 9 1 7 9 0 13 15 14 13 1 12 9 1 9 15 9 1 9 9 0 2
4 9 12 9 0
25 1 9 0 2 13 9 1 9 0 3 7 12 1 9 9 13 1 9 1 9 8 0 0 8 2
31 7 13 10 9 7 9 9 9 13 1 9 7 13 13 9 9 0 1 9 2 15 13 1 12 9 1 9 1 9 0 2
28 7 13 9 9 8 7 8 13 1 9 13 9 15 1 9 2 7 13 1 9 9 15 1 9 9 15 0 2
21 7 13 1 7 8 13 9 9 15 13 1 15 9 0 0 1 9 0 1 9 2
5 9 0 8 8 9
41 7 13 10 9 7 13 9 0 3 0 1 9 9 2 9 9 0 2 0 7 1 2 0 2 7 13 1 2 15 14 9 2 9 9 9 2 9 1 15 2 2
54 7 13 9 9 1 9 9 0 1 9 13 9 8 8 9 1 15 2 8 8 9 7 9 9 9 1 9 9 0 7 9 9 0 9 1 10 9 7 15 13 15 1 9 9 13 9 9 7 9 1 8 8 2 2
69 7 13 9 2 13 1 9 7 13 7 15 14 13 1 9 9 1 9 7 9 15 14 1 9 0 7 1 8 9 9 0 2 0 7 2 9 9 9 9 8 8 7 9 9 9 7 9 9 1 15 15 1 9 15 13 1 9 9 15 7 9 9 15 1 10 14 9 2 2
46 7 13 9 0 7 2 9 14 13 0 1 9 9 7 9 8 8 9 1 9 0 9 1 9 8 2 2 2 2 2 7 9 0 7 0 13 8 8 9 9 7 9 15 0 2 2
7 9 0 13 9 9 8 8
39 8 2 9 9 2 2 13 9 0 9 1 9 9 0 1 9 1 9 8 0 1 8 13 9 10 9 7 7 15 13 9 9 0 7 13 9 9 0 2
33 7 13 9 2 8 8 2 1 9 1 9 7 9 0 7 9 9 0 1 9 13 1 9 0 1 9 0 7 9 1 9 0 2
61 7 13 10 9 13 9 9 1 9 15 1 9 9 0 7 13 8 8 7 9 15 1 9 0 1 9 7 13 1 9 1 9 8 8 8 0 13 1 9 9 0 1 9 15 13 1 15 9 0 9 1 8 9 15 1 9 13 1 12 9 2
28 7 13 9 10 13 1 10 9 7 15 13 1 15 1 9 9 1 9 0 1 15 1 9 9 9 9 8 2
2 9 9
26 1 9 13 9 8 9 1 10 9 7 13 9 0 1 9 9 13 9 9 9 0 7 0 1 8 2
41 7 13 9 0 0 1 8 8 9 15 0 1 9 7 9 7 0 1 9 0 1 9 1 10 13 15 8 9 2 0 7 0 2 1 8 8 9 2 9 2 2
31 7 13 0 9 0 0 9 9 10 9 0 15 13 8 9 15 9 9 9 7 13 9 0 1 9 9 9 0 7 0 2
35 7 13 9 1 9 1 9 9 15 1 8 7 13 9 15 1 9 1 9 0 7 13 15 1 15 13 1 8 7 9 0 7 0 3 2
36 7 13 1 7 9 9 9 0 1 9 0 1 9 2 8 2 13 9 1 9 0 1 9 0 1 8 9 1 9 9 1 9 0 1 15 2
1 9
9 9 9 0 13 1 15 9 0 2
11 13 7 13 0 9 0 1 10 13 15 2
15 13 15 9 0 1 9 0 7 13 0 1 9 1 9 2
19 8 1 9 1 9 1 1 9 1 9 9 9 1 9 0 1 9 9 2
9 0 9 15 10 9 15 9 9 2
1 9
12 13 0 1 9 15 1 9 15 13 8 0 2
17 14 14 13 1 9 15 13 1 15 10 9 1 9 7 9 9 2
17 9 15 0 7 0 7 14 13 3 9 9 0 1 9 9 15 2
14 9 13 1 15 1 0 1 9 7 13 9 15 0 2
9 0 9 15 10 9 15 9 9 2
1 8
14 14 13 1 9 15 13 1 15 7 13 9 9 0 2
27 13 1 9 15 13 1 1 15 8 1 9 7 13 3 1 9 9 8 15 13 8 8 1 9 1 15 2
9 14 13 3 9 1 9 7 9 2
12 1 15 1 9 1 9 9 1 9 9 9 2
9 0 9 15 10 9 15 9 9 2
1 9
8 1 15 9 1 9 10 9 2
10 14 13 7 13 1 15 9 9 15 2
15 0 9 0 1 9 14 13 0 15 14 13 1 9 15 2
8 1 15 1 9 1 9 15 2
9 0 9 15 10 9 15 9 9 2
1 9
11 14 13 1 9 0 9 9 15 0 0 2
15 13 15 9 0 13 15 1 1 15 9 9 0 1 9 2
14 13 9 9 9 1 9 7 9 15 14 13 15 0 2
5 8 0 9 0 2
9 0 9 15 10 9 15 9 9 2
1 9
12 14 13 9 9 1 9 9 9 7 9 0 2
26 13 1 9 1 9 9 9 7 9 0 0 7 1 9 9 15 1 9 1 9 7 15 0 1 15 2
10 9 14 13 1 8 0 7 9 9 2
9 14 13 1 9 1 9 7 9 2
9 0 9 15 10 9 15 9 9 2
1 9
11 9 9 0 7 9 0 1 9 9 0 2
9 13 1 9 9 0 1 10 13 2
11 14 13 1 9 0 1 9 9 1 10 2
12 15 13 1 9 0 1 9 15 1 9 15 2
9 0 9 15 10 9 15 9 9 2
1 9
9 9 9 0 13 1 15 9 0 2
11 13 7 13 0 9 0 1 10 13 15 2
15 13 15 9 9 1 9 0 7 13 0 1 9 1 9 2
19 13 1 9 1 9 1 1 9 1 9 9 9 1 9 0 1 9 9 2
9 0 9 15 10 9 15 9 9 2
1 9
8 9 13 1 9 9 9 0 2
9 14 13 15 1 9 7 9 0 2
12 13 7 14 13 1 9 15 1 9 10 9 2
14 13 7 15 13 1 9 9 0 1 7 13 0 9 2
9 0 9 15 10 9 15 9 9 2
1 9
15 13 9 1 9 0 1 15 7 14 13 1 15 1 9 2
10 13 9 15 0 1 9 9 9 9 2
13 13 1 9 9 9 7 13 13 1 9 0 15 2
16 14 9 1 9 9 1 10 13 7 14 13 3 9 1 9 2
9 0 9 15 10 9 15 9 9 2
1 9
12 14 13 9 15 13 1 15 1 9 9 15 2
13 14 14 13 0 1 9 0 1 9 15 13 15 2
9 14 13 0 1 9 7 9 9 2
29 14 13 15 7 13 9 9 15 1 9 7 13 9 1 15 7 7 13 9 15 7 7 15 14 13 15 1 9 2
9 0 9 15 10 9 15 9 9 2
1 9
12 14 13 0 13 1 15 7 13 1 9 15 2
23 13 0 1 9 15 7 7 13 9 15 13 15 1 9 9 7 1 9 1 9 1 15 2
7 14 14 13 9 9 15 2
9 14 13 1 9 1 9 7 9 2
9 0 9 15 10 9 15 9 9 2
1 8
6 13 9 1 9 0 2
13 13 15 9 1 9 0 1 9 9 1 9 0 2
16 14 13 9 0 0 1 0 9 7 14 13 1 0 9 0 2
12 13 1 9 0 1 9 15 7 9 15 0 2
9 0 9 15 10 9 15 9 9 2
13 9 0 1 8 9 0 9 1 9 1 9 7 9
66 13 9 9 0 1 9 9 0 1 9 0 1 9 9 8 9 11 8 1 0 9 15 13 15 0 9 15 7 0 9 15 7 13 1 9 1 9 9 8 13 1 9 7 9 7 13 0 0 13 1 9 0 9 7 9 7 9 0 1 9 9 8 0 7 9 2
53 7 7 13 9 9 0 9 9 9 0 1 10 13 9 15 1 9 9 15 0 0 2 7 9 0 15 9 0 10 9 15 13 9 7 13 9 1 9 9 0 1 9 9 1 15 13 1 15 1 12 12 9 2
87 7 13 9 9 9 8 9 11 8 1 9 7 9 7 9 7 9 1 9 9 15 7 13 1 9 9 0 1 9 10 9 1 9 10 13 1 15 1 9 0 7 9 0 1 1 9 15 1 9 7 9 7 9 7 9 7 9 9 15 13 15 9 9 15 7 9 15 1 9 15 0 7 0 7 0 1 0 9 1 9 9 0 1 9 7 9 2
62 7 13 9 9 15 10 9 1 9 9 1 9 7 13 9 15 1 9 1 9 0 1 0 9 9 2 0 9 1 10 9 0 0 15 13 1 9 7 9 9 0 1 9 7 9 7 13 1 15 9 9 0 1 9 0 9 9 0 1 9 0 2
58 7 9 10 9 13 1 9 9 9 15 13 1 15 10 9 0 1 15 15 9 1 9 9 0 13 9 0 7 0 1 9 0 0 0 1 9 15 7 9 15 7 0 1 9 15 7 0 15 1 9 9 15 1 0 9 7 9 2
68 7 13 9 1 9 15 13 1 9 0 1 9 8 1 0 8 11 8 1 9 7 0 9 9 8 8 15 13 9 9 8 9 11 8 1 9 9 0 1 9 15 9 9 8 9 2 9 9 9 1 15 1 10 1 10 1 9 1 9 7 9 1 9 1 9 7 9 2
43 14 9 9 1 9 10 0 7 15 9 9 15 1 9 0 9 1 8 7 15 9 15 13 1 9 9 1 9 15 7 13 9 9 9 7 9 15 13 1 10 9 0 2
3 1 9 9
9 8 13 1 9 1 9 0 1 8
33 8 2 8 8 2 2 13 9 1 9 0 7 8 13 1 9 9 3 1 9 9 0 1 9 13 1 8 9 9 15 1 9 2
30 7 13 9 7 15 14 13 13 8 1 9 9 7 13 9 1 9 1 9 1 9 1 9 13 9 9 9 14 12 2
14 7 9 9 0 0 1 9 13 9 9 1 10 9 2
29 7 13 9 9 15 13 15 8 7 9 0 9 1 9 9 9 0 1 9 9 13 1 8 9 9 15 1 9 2
20 7 13 9 7 2 9 9 13 1 9 7 13 9 9 0 2 1 9 0 2
24 7 13 9 9 1 9 0 1 9 0 8 8 9 9 1 9 9 12 9 1 9 9 8 2
17 7 13 9 1 9 1 9 8 8 7 9 9 10 9 14 13 2
23 13 1 7 9 13 9 0 9 1 9 9 9 0 0 1 9 9 1 9 0 14 12 2
23 7 13 8 9 9 1 12 9 1 0 7 9 9 9 9 1 0 1 9 12 0 9 2
47 7 13 9 9 0 14 13 1 9 9 9 0 1 9 15 13 15 9 0 1 9 0 8 8 7 13 1 15 1 9 9 8 1 9 9 0 15 13 15 1 9 9 0 0 1 9 2
25 7 14 13 9 12 15 13 15 8 7 9 0 3 1 8 9 9 1 9 15 1 9 0 0 2
30 7 9 8 10 9 1 0 1 9 13 9 9 0 1 9 9 1 9 9 9 9 8 8 0 8 1 9 12 9 2
32 7 13 9 0 8 8 13 1 12 9 0 1 9 0 9 0 7 0 1 9 15 1 9 1 9 7 9 1 9 15 0 2
21 7 14 13 8 13 1 1 12 12 9 1 9 1 9 9 13 15 1 9 9 2
4 0 1 9 0
7 9 9 0 1 9 0 9
44 9 2 9 2 14 13 9 0 9 0 1 9 0 7 1 9 9 12 7 13 7 13 9 9 0 0 7 13 12 5 1 9 9 7 15 15 9 15 7 13 9 0 0 2
71 9 0 0 7 14 13 15 1 1 9 9 1 9 1 9 0 1 9 0 1 9 9 7 9 7 9 9 1 9 9 9 0 1 9 1 9 1 9 9 7 7 9 9 9 1 9 14 13 9 9 9 1 9 0 1 15 13 9 0 1 9 1 9 13 1 9 0 1 9 0 2
3 9 0 9
69 1 10 9 14 13 9 9 1 9 1 9 9 0 1 10 13 1 9 9 0 7 9 0 0 9 7 9 1 15 14 13 9 1 8 9 0 1 9 0 1 1 9 14 13 1 9 1 15 2 7 1 9 9 8 7 15 1 9 9 12 14 13 9 9 9 1 9 9 2
5 9 0 1 9 0
101 7 1 9 0 7 9 1 9 9 9 0 7 0 1 9 9 7 14 13 7 13 9 1 15 9 0 7 14 13 9 9 0 1 0 1 9 9 9 7 9 9 7 9 9 7 9 9 1 9 0 1 9 9 2 13 1 10 9 7 15 14 13 9 0 1 9 9 1 9 9 7 14 13 9 9 0 1 9 9 9 7 9 7 9 9 2 9 1 9 9 0 1 9 0 7 0 7 9 1 15 2
3 9 9 9
81 7 1 9 14 13 9 1 7 13 9 9 9 7 0 0 1 7 13 9 15 1 9 7 9 1 15 13 1 9 1 9 9 1 15 1 12 9 1 9 12 9 2 7 14 13 9 9 1 9 0 13 1 9 9 7 9 9 1 9 9 0 1 9 9 9 7 9 9 1 9 1 9 9 1 9 9 0 14 0 9 2
45 7 1 9 9 1 9 14 13 9 1 0 9 0 1 1 9 9 0 15 13 1 15 7 15 10 13 1 9 9 9 1 9 9 0 1 9 1 15 13 9 0 1 9 0 2
5 9 0 1 9 9
35 7 10 9 0 15 13 1 9 12 1 9 9 11 8 0 13 1 15 1 9 9 0 1 9 9 13 1 15 1 0 9 9 2 2 2
46 7 14 13 9 9 0 1 9 9 0 1 0 1 9 15 13 9 15 0 0 1 8 7 9 7 9 0 1 9 10 13 1 9 0 9 1 9 9 1 10 13 1 9 9 0 2
2 8 8
7 15 14 13 9 0 1 2
50 9 2 9 2 13 9 1 9 7 1 9 7 9 0 1 9 9 1 9 0 7 9 0 13 9 1 9 7 13 9 1 9 7 9 1 9 1 9 1 9 1 9 0 7 0 15 13 1 9 2
62 7 13 10 9 7 13 9 9 1 9 0 1 9 9 7 7 10 9 15 13 1 15 9 0 13 1 9 0 1 9 0 0 1 9 9 9 7 3 1 9 9 9 7 15 15 13 1 9 9 7 9 9 1 9 0 7 1 9 7 9 0 2
4 9 1 8 0
70 7 13 9 9 1 9 14 13 1 9 9 9 7 1 9 0 1 9 1 9 9 1 9 9 9 1 9 9 9 15 1 9 0 7 13 9 9 0 1 15 7 3 7 14 13 9 9 0 1 9 1 9 0 9 1 9 7 9 1 9 0 7 13 1 9 1 0 1 9 2
71 7 9 7 9 9 13 1 9 7 9 1 9 14 7 15 7 1 1 9 1 9 9 9 14 13 9 9 1 9 0 7 7 9 0 7 3 9 9 0 14 13 1 9 15 1 9 1 9 3 7 13 9 1 9 15 13 1 9 1 9 7 15 13 9 1 15 1 9 9 0 2
3 9 1 9
52 7 1 9 2 9 2 9 9 13 9 0 1 9 1 9 0 1 9 1 9 1 9 9 9 7 7 13 9 13 0 1 9 7 9 9 13 13 1 9 7 9 9 10 9 0 7 13 1 9 7 9 2
35 8 9 9 15 8 8 1 9 13 9 9 1 9 1 9 9 9 9 9 1 9 9 7 3 1 9 0 15 8 1 15 9 3 0 2
2 8 8
1 9
7 9 9 1 9 7 9 9
57 1 9 9 9 0 13 9 0 1 9 9 1 9 1 9 1 9 9 9 8 7 0 1 9 9 1 9 2 2 9 0 7 9 0 2 9 1 15 13 9 1 9 9 0 0 7 9 9 9 9 7 9 9 1 9 9 2
44 7 14 13 9 9 1 9 1 9 9 0 7 9 9 9 1 9 7 9 1 9 9 9 1 9 9 0 1 9 9 1 9 7 9 1 15 1 9 7 9 9 1 9 2
81 7 13 9 1 9 0 0 7 0 1 9 1 9 0 0 1 9 7 15 13 9 15 1 9 0 7 9 9 9 0 7 9 9 0 1 9 0 1 9 9 1 9 1 9 7 9 1 9 9 0 10 13 15 1 9 7 9 9 0 0 9 9 9 0 9 0 7 3 9 9 9 15 13 9 15 9 0 7 9 0 2
72 9 1 7 9 13 1 9 1 9 0 0 0 1 9 9 12 7 9 15 2 9 1 9 9 9 7 9 1 9 9 0 13 1 15 0 9 9 7 9 9 1 9 9 7 9 7 9 7 9 9 7 9 1 9 15 1 9 9 1 9 7 9 0 9 9 9 9 0 7 9 0 2
50 1 9 0 13 9 1 9 0 1 9 1 9 1 1 9 8 9 9 9 0 0 1 9 9 1 9 9 1 9 9 7 9 7 9 9 7 13 9 1 9 9 1 9 0 7 1 9 0 0 2
3 8 8 2
2 1 8
8 13 9 15 7 13 9 9 0
19 13 9 9 8 8 1 9 12 9 13 9 15 1 9 9 1 9 0 2
40 7 14 13 9 13 7 13 8 15 13 1 15 9 13 7 15 13 9 1 12 9 13 9 0 1 9 1 9 7 13 1 15 1 7 15 1 9 7 0 2
46 9 10 9 13 9 9 13 1 9 15 7 9 15 9 15 13 15 1 9 9 1 12 9 13 9 15 1 9 0 1 9 14 7 15 13 1 9 0 9 9 10 1 9 15 0 0
80 7 1 9 9 0 1 15 12 13 9 15 0 1 9 9 7 13 1 9 9 9 1 9 9 1 9 0 7 13 9 15 7 1 9 1 9 13 1 15 13 1 15 7 14 13 9 15 7 14 13 9 1 9 15 1 9 9 9 0 13 15 1 9 1 9 9 0 7 13 13 15 1 9 9 1 9 15 13 15 2
21 7 14 13 0 12 1 9 0 1 12 9 13 1 15 9 9 1 12 12 9 2
24 7 1 9 9 1 0 13 9 15 9 9 9 1 9 9 7 13 15 15 9 1 9 15 2
1 8
21 7 13 9 1 15 1 9 1 9 1 9 15 2 9 2 9 9 9 0 1 9
156 7 13 0 13 9 0 1 9 9 9 9 15 1 12 9 0 2 7 13 1 9 9 0 1 0 1 12 9 2 7 13 0 1 7 9 0 9 1 9 9 0 14 13 9 9 0 7 13 1 9 0 1 9 9 2 9 2 0 1 9 15 2 7 13 9 0 9 9 1 9 9 1 9 0 13 1 9 9 9 9 1 0 2 1 9 7 9 0 1 9 9 13 2 7 13 7 9 1 9 1 9 1 12 9 0 1 9 0 1 9 0 13 1 9 1 9 12 0 7 13 9 15 1 9 1 9 9 0 1 9 9 0 2 7 7 0 13 1 9 1 9 0 1 9 9 2 1 9 0 12 9 2 13 10 9 2
59 7 13 2 9 2 7 9 1 9 13 9 1 9 10 13 1 9 9 9 15 7 9 1 0 9 1 9 9 0 7 9 1 9 9 9 0 0 7 9 9 9 9 1 9 9 7 13 15 1 9 9 0 0 13 9 9 1 15 2
12 9 0 13 1 9 1 9 1 9 1 9 8
2 8 8
61 13 9 9 1 9 9 1 9 9 9 9 1 9 2 9 8 0 2 15 13 9 1 9 9 2 7 14 13 9 2 9 0 9 2 15 13 9 9 9 9 1 9 15 14 13 9 0 2 9 1 9 1 9 1 9 9 1 9 9 8 2
68 13 9 1 9 0 0 7 9 9 13 1 9 9 13 1 9 9 1 9 1 9 15 13 15 9 9 1 9 1 9 9 8 0 2 7 15 14 13 9 1 9 15 13 0 2 7 13 1 7 9 14 13 1 9 9 1 9 9 9 15 13 7 13 15 9 9 0 2
68 7 13 8 8 13 1 9 1 9 1 9 9 9 0 1 9 15 1 9 7 13 9 15 1 15 7 13 7 9 14 13 9 1 9 9 1 9 1 15 2 7 13 9 7 9 13 1 9 9 9 1 9 9 1 9 7 7 13 9 9 1 15 1 9 1 9 9 2
87 7 13 9 9 9 9 1 9 1 9 1 9 15 13 1 15 12 9 1 15 12 9 7 12 9 1 15 12 9 7 15 13 9 12 0 7 9 1 9 13 15 1 9 0 1 12 9 1 12 0 9 2 7 13 9 1 9 0 1 9 9 2 9 9 1 9 9 2 2 7 13 9 13 9 9 0 2 9 10 15 0 1 12 1 8 2 2
91 7 13 9 9 1 9 1 9 1 9 9 13 1 1 15 9 1 9 1 15 2 7 13 7 13 9 0 1 9 9 9 1 9 9 2 7 13 9 1 9 9 9 9 9 1 9 0 0 2 7 13 1 0 3 1 9 1 9 9 2 7 1 9 9 9 13 9 9 0 3 1 9 15 1 9 0 15 13 9 9 15 13 9 1 9 1 9 9 9 0 2
79 7 13 7 13 9 9 1 9 8 9 15 1 9 2 9 0 0 2 0 9 12 9 2 13 2 0 2 7 15 14 13 9 9 1 15 9 9 0 2 7 13 9 0 7 9 9 14 13 1 0 1 9 2 7 7 9 9 14 13 1 9 9 0 1 9 0 1 7 13 9 9 0 0 1 9 9 12 0 2
24 9 0 1 9 9 12 12 1 9 9 2 9 2 2 9 2 13 9 9 9 1 9 9 9
2 8 8
61 13 9 2 9 0 2 9 9 0 1 9 1 9 15 1 9 9 9 0 9 9 0 2 7 13 9 7 9 15 1 9 0 1 9 9 9 8 8 2 13 1 9 0 1 1 9 0 2 2 7 13 7 8 2 0 9 1 9 9 2 2
106 13 9 0 0 7 9 9 0 13 9 0 0 1 9 9 9 9 9 0 9 9 0 2 7 13 1 7 9 0 1 9 9 1 9 7 9 13 1 9 9 9 1 1 9 1 15 1 9 9 14 13 1 9 0 2 7 14 13 0 1 12 12 9 1 9 15 13 1 9 0 1 9 0 1 9 9 9 13 1 9 0 9 0 1 9 0 0 2 7 13 1 9 9 1 9 0 1 7 13 9 1 15 9 9 12 2
134 7 13 9 9 0 9 1 9 9 0 9 9 11 3 7 9 9 14 13 1 9 9 0 1 9 7 9 0 1 9 2 9 1 9 1 9 9 1 9 2 7 13 7 9 13 9 9 15 13 1 9 1 9 1 9 7 9 15 0 13 2 1 9 9 14 13 1 9 9 1 9 15 13 14 13 9 9 2 9 2 0 7 13 1 9 0 1 9 9 1 9 9 9 2 15 13 7 0 1 9 15 13 9 15 0 14 13 9 1 9 9 9 2 2 7 13 9 11 9 9 9 1 9 9 9 1 1 9 9 0 7 9 9 2
39 7 13 9 9 9 0 1 9 9 8 8 8 0 7 13 9 2 9 9 2 3 7 9 15 1 9 2 14 13 0 1 9 9 15 13 9 9 2 2
44 7 13 9 12 1 9 0 1 15 1 9 1 12 9 0 1 9 9 2 1 9 7 2 9 2 13 13 1 9 9 9 0 2 7 13 9 9 9 9 1 9 9 8 8
75 1 2 9 2 7 2 9 2 14 13 9 2 1 9 15 0 9 1 9 9 9 2 2 0 7 9 13 1 9 1 9 9 2 9 2 2 7 13 1 7 9 9 0 2 13 0 13 9 1 9 1 9 9 13 1 9 1 9 7 9 1 9 9 9 9 7 9 9 0 1 9 7 9 2 2
153 7 13 8 9 9 0 1 9 2 9 2 1 9 9 13 15 13 1 9 0 0 2 7 13 2 9 13 9 1 9 2 7 3 9 1 9 1 9 7 9 1 9 13 9 1 15 1 9 1 9 2 7 9 9 9 9 1 9 7 7 0 10 13 1 9 9 1 9 1 1 9 15 9 0 8 8 0 1 9 0 7 1 0 7 7 9 14 13 9 15 1 9 9 1 9 0 1 15 1 14 13 1 9 1 9 1 9 9 9 14 13 1 9 9 7 9 1 9 2 2 7 13 7 9 9 9 1 9 0 0 9 0 8 8 7 9 0 8 8 2 13 0 1 8 8 1 9 9 1 9 9 2 2
11 9 0 2 0 1 9 9 7 9 7 9
2 8 8
33 13 9 0 9 9 1 9 0 7 0 1 9 1 9 7 9 1 9 9 15 13 1 15 9 0 1 9 9 9 9 9 0 2
35 7 14 13 9 1 9 9 2 9 2 0 9 9 7 9 8 0 8 8 8 1 9 9 1 9 9 0 7 9 9 9 9 9 0 2
31 7 13 9 1 12 1 9 0 9 9 7 9 0 8 8 8 8 8 8 1 9 9 1 8 8 8 8 8 8 8 2
43 7 14 13 9 1 9 9 1 9 1 9 9 9 7 9 0 7 0 7 0 7 3 1 9 9 0 2 7 13 9 0 1 12 12 9 1 9 1 9 1 10 9 2
47 7 14 13 9 9 9 0 1 9 1 9 9 1 9 13 0 1 9 12 12 9 1 10 9 2 7 13 9 0 7 13 9 9 0 9 0 1 9 9 9 1 9 1 12 12 9 2
63 13 1 7 9 7 9 13 1 12 9 0 2 9 2 0 1 9 9 9 0 1 9 9 9 0 11 8 8 1 9 2 7 13 9 0 0 13 9 9 7 9 9 8 8 8 8 8 8 9 0 9 1 9 1 9 9 0 13 12 1 9 9 2
19 7 13 9 0 1 9 9 9 0 2 7 14 13 9 0 1 3 9 2
27 7 13 9 1 9 0 9 9 0 1 9 2 9 7 3 12 9 0 13 9 1 9 2 9 2 0 2
18 7 13 9 9 0 9 1 9 0 1 9 9 7 9 9 9 0 2
16 9 0 8 8 13 1 9 1 9 7 13 15 1 9 9 2
2 8 8
204 13 7 9 13 7 13 9 0 9 9 9 1 9 9 1 9 10 15 0 2 7 9 15 13 15 9 14 13 1 2 1 9 9 9 9 1 9 9 15 9 9 0 1 9 9 0 1 9 2 9 1 9 2 13 1 15 1 9 9 1 9 2 9 2 1 9 0 2 7 13 9 1 9 0 7 13 15 9 2 9 1 9 2 1 9 7 13 15 1 9 7 13 15 1 9 1 9 9 7 9 1 9 0 1 9 7 13 1 9 1 1 9 2 7 9 14 13 1 9 15 7 7 13 1 9 15 7 9 15 2 7 9 13 9 9 15 13 15 9 0 7 9 9 9 7 9 1 9 7 9 0 7 0 1 9 15 13 9 1 9 9 7 9 0 9 1 9 9 1 9 2 13 9 7 13 9 9 0 0 15 13 1 9 9 0 0 9 9 0 1 9 9 9 9 9 0 9 1 9 0 1 9 9 2
71 13 9 13 9 2 9 1 9 2 1 9 15 0 1 9 1 9 7 1 9 15 12 9 7 1 13 1 9 1 9 1 9 9 2 7 1 12 9 1 9 9 2 13 1 9 9 1 9 12 9 1 9 9 13 1 15 9 1 9 7 9 9 7 9 13 1 9 1 9 0 2
113 9 1 9 1 9 9 9 13 9 9 9 15 7 9 9 9 1 9 1 9 9 0 1 9 9 2 7 15 13 9 7 8 8 2 8 2 7 14 13 9 15 0 1 0 1 15 2 7 1 15 14 13 9 15 2 1 13 15 1 9 1 9 0 0 0 1 15 9 2 1 7 13 9 13 1 9 1 15 2 7 13 9 7 13 9 0 9 9 0 2 7 13 1 9 15 8 9 9 1 9 9 0 0 0 15 13 13 15 9 9 8 8 2
229 13 9 1 0 1 9 9 7 9 0 1 9 1 9 1 9 2 7 13 9 1 2 9 2 7 15 13 1 9 9 9 1 9 9 7 13 7 9 9 1 9 14 13 9 0 1 9 7 9 9 2 7 13 7 15 13 1 9 9 1 9 12 9 2 7 15 13 12 9 0 0 1 9 2 7 13 12 1 15 1 9 9 15 7 13 0 1 9 0 1 15 2 7 13 7 15 13 9 12 13 9 1 9 9 9 2 7 13 7 15 1 0 1 9 9 13 9 0 0 7 15 14 13 1 9 3 7 13 9 1 9 9 7 13 1 9 2 7 15 13 9 1 9 7 9 15 0 1 9 9 2 7 15 1 9 0 13 1 15 1 14 9 9 15 13 15 1 9 0 1 7 13 15 9 1 9 9 7 13 1 15 9 9 15 2 10 9 14 13 1 9 7 13 7 15 13 9 0 2 7 14 13 2 9 1 9 2 9 9 0 1 9 15 9 0 7 9 15 1 9 7 1 9 15 1 9 1 9 2
11 9 2 9 2 12 2 2 2 7 14 13
2 8 8
65 13 9 2 9 0 2 9 1 9 1 9 1 12 1 9 15 13 9 15 1 9 9 9 9 0 9 9 15 9 1 10 13 1 12 1 9 9 1 9 0 2 7 9 9 3 1 9 9 8 8 1 9 13 9 9 1 9 0 1 9 9 1 10 9 2
86 13 9 9 3 1 9 0 1 9 2 9 0 2 9 8 8 1 9 1 9 1 9 1 9 13 15 2 9 9 9 0 2 7 13 1 9 12 9 1 9 8 1 9 2 1 9 0 0 8 2 2 7 13 8 9 9 1 9 15 1 7 15 2 9 0 2 7 13 1 9 15 1 2 7 13 9 1 9 15 13 1 15 1 9 2 2
75 7 13 7 13 9 9 1 9 12 1 9 9 1 9 0 8 1 3 1 8 8 9 8 8 1 9 9 9 9 2 9 0 7 4 9 0 8 1 9 9 1 9 1 9 2 2 7 13 15 9 0 15 13 1 15 9 9 1 9 1 9 9 1 9 15 9 0 7 13 12 9 1 9 8 2
50 7 13 8 9 9 11 11 1 9 15 1 9 12 9 2 0 1 7 12 1 15 8 9 8 11 8 7 9 8 8 8 8 13 1 9 9 1 9 1 9 13 0 9 9 8 8 1 9 0 2
153 7 13 2 9 2 7 9 13 1 9 12 1 9 15 3 1 9 1 9 2 7 13 9 2 9 2 7 9 9 9 13 9 12 1 9 1 9 0 2 7 7 9 9 14 13 1 9 9 2 7 13 9 7 10 9 2 14 13 9 1 9 7 9 0 0 2 7 13 1 9 15 1 7 14 13 9 0 9 1 9 9 7 9 0 1 9 1 0 1 9 0 1 9 9 2 7 13 9 1 7 1 9 9 9 2 9 2 1 9 0 2 9 2 0 15 13 1 15 12 1 2 9 2 1 9 0 2 7 13 9 7 9 13 1 9 9 1 9 9 9 13 1 2 9 9 9 15 0 1 9 0 2 2
74 7 1 9 7 9 13 1 9 9 9 9 15 1 9 9 1 7 13 9 9 9 9 15 1 9 2 14 7 2 9 2 13 7 9 13 9 9 8 8 1 9 1 9 9 9 2 7 13 9 9 8 8 8 1 9 1 9 2 8 8 8 2 1 9 9 7 15 1 9 9 0 1 9 2
11 9 1 9 0 13 9 1 9 9 8 8
39 13 9 9 0 9 8 8 0 9 1 12 9 13 1 2 9 2 9 1 9 7 13 1 15 9 0 8 8 9 9 15 1 2 9 9 8 8 2 2
59 7 13 8 1 9 9 0 9 13 15 1 12 9 0 1 3 13 1 15 1 9 9 0 7 9 9 9 1 9 9 0 1 9 9 15 0 1 9 9 1 9 0 2 0 7 15 13 15 2 9 9 0 13 15 9 1 9 2 2
113 7 1 9 15 0 0 13 8 1 7 2 9 0 1 9 9 0 1 9 9 9 7 1 9 15 9 9 9 0 0 1 9 9 7 0 1 9 2 2 0 7 2 9 0 0 13 1 9 9 0 1 9 1 9 7 9 9 9 7 9 9 0 2 2 7 13 9 0 9 9 15 1 9 0 1 2 9 9 1 9 9 1 9 0 9 12 9 1 9 9 0 1 9 0 1 9 15 13 1 9 1 9 15 9 9 9 9 9 0 1 9 2 2
36 7 13 8 1 7 2 9 0 1 9 13 1 9 0 1 9 0 7 13 9 0 8 0 7 3 9 0 1 9 9 0 1 8 0 2 2
58 7 13 9 9 0 0 1 9 15 1 9 9 9 8 8 2 7 13 7 13 12 9 1 9 1 9 9 1 9 9 15 1 9 9 12 9 1 8 8 2 8 8 14 13 8 0 1 9 9 9 3 13 9 9 0 1 9 2
31 12 9 1 9 9 9 7 9 9 9 1 9 0 2 9 2 2 9 2 14 13 9 9 15 7 13 9 1 9 9 15
5 9 8 2 9 9
67 14 13 1 9 2 9 0 2 9 1 9 0 1 9 9 0 1 9 9 15 13 9 0 1 9 2 7 13 9 9 1 9 0 13 1 9 9 1 9 15 7 9 10 1 9 9 9 2 1 9 13 9 12 1 2 9 2 1 9 9 7 13 12 0 1 9 2
73 1 9 9 9 9 1 9 9 9 0 9 0 1 9 2 14 7 9 9 2 9 0 2 14 13 1 9 9 9 15 15 13 1 9 9 13 7 15 13 1 9 9 15 1 9 7 13 9 9 15 1 9 9 2 7 13 9 15 1 9 1 9 9 9 9 1 9 9 15 1 9 9 2
118 7 13 9 1 2 9 2 7 14 13 9 9 9 1 12 1 15 12 13 1 9 0 7 13 9 9 1 9 2 7 13 0 7 9 13 9 1 12 1 9 9 1 9 8 9 2 7 13 7 9 1 9 13 1 9 9 9 1 9 1 9 9 15 2 7 13 9 1 9 8 12 1 2 9 2 2 13 9 7 15 13 13 9 9 15 2 7 13 2 9 2 9 3 1 9 2 9 9 0 2 13 1 9 0 13 9 1 9 9 9 1 9 9 0 1 9 15 2
263 7 13 9 2 9 2 15 13 1 0 1 9 15 1 9 1 9 0 2 1 9 13 1 15 9 7 9 13 8 9 0 2 7 7 2 9 0 9 0 2 2 7 13 9 9 15 13 1 9 9 1 9 12 1 9 2 9 2 1 15 12 1 9 1 15 13 9 9 2 7 13 9 9 9 13 1 9 1 9 9 1 9 9 2 9 2 1 9 9 9 15 7 1 15 15 13 1 2 2 8 8 9 8 7 13 8 11 8 1 8 8 8 8 1 9 9 9 15 1 7 13 9 15 9 2 14 7 9 8 8 2 7 1 13 9 2 8 8 8 8 7 11 11 8 8 8 8 8 8 8 8 8 2 7 1 15 9 15 1 9 9 1 9 8 1 9 9 9 13 9 9 9 15 1 9 7 9 9 9 9 9 0 2 7 13 9 1 9 8 0 7 13 9 9 15 13 9 13 1 9 15 9 9 1 9 9 15 7 9 1 9 1 9 9 7 9 15 1 9 0 1 9 14 7 15 13 9 15 1 9 1 0 9 7 1 9 9 9 9 2 7 13 8 8 13 15 8 9 9 1 9 0 0 1 7 13 9 9 15 1 9 2 2
88 7 13 7 2 9 2 13 1 9 9 0 1 9 15 1 9 0 12 2 9 7 9 7 9 2 7 13 1 15 15 13 1 9 9 1 9 0 2 7 13 8 11 11 7 9 8 8 13 1 9 9 9 1 9 1 9 1 9 8 8 15 13 9 13 9 1 9 15 1 9 8 8 13 1 9 1 12 1 15 13 0 1 9 15 13 9 15 2
58 7 13 9 9 1 9 9 9 12 9 2 7 13 9 9 12 9 0 1 9 1 15 9 9 0 2 9 1 9 9 9 9 1 9 0 0 2 7 13 9 0 1 9 0 0 1 9 9 15 1 9 9 1 9 9 9 0 2
48 7 1 9 9 9 2 9 0 2 1 9 9 1 9 2 1 9 15 1 9 2 14 7 15 14 13 9 9 9 15 13 9 0 1 9 0 0 2 7 13 12 1 12 1 9 15 0 2
65 7 13 9 0 9 1 9 1 9 0 9 8 8 8 1 9 2 9 9 2 9 8 8 1 9 13 9 2 9 9 2 7 13 9 9 0 1 9 8 8 1 9 9 0 1 9 9 8 8 1 9 8 2 7 13 9 9 7 9 9 13 1 9 9 2
77 7 13 12 9 1 9 0 15 13 13 1 9 1 9 0 3 2 7 13 12 1 9 9 2 9 2 7 13 12 1 9 9 2 9 2 7 12 1 2 9 2 7 12 1 2 0 2 7 12 1 2 0 2 1 15 9 2 7 13 9 12 1 9 2 9 2 7 13 9 9 1 9 9 1 12 9 2
22 7 1 9 15 13 1 9 9 9 9 14 7 9 15 1 9 0 13 9 9 9 2
13 9 2 12 12 9 9 8 9 1 9 9 9 0
2 8 8
46 13 7 13 9 9 0 1 9 9 0 1 9 0 1 9 9 9 0 2 1 9 15 1 1 12 12 9 1 9 9 13 7 9 9 14 13 0 9 1 9 9 9 1 9 0 2
52 13 9 9 0 1 9 0 1 9 9 9 9 7 9 9 1 9 9 9 1 9 12 1 12 2 7 13 9 1 9 9 9 0 7 15 13 0 1 9 0 7 0 1 1 1 0 7 0 2 0 2 2
99 7 13 1 9 9 9 9 9 9 1 9 9 0 0 7 13 0 1 9 9 1 9 0 2 15 13 1 9 9 9 15 9 9 1 9 0 2 7 13 9 15 9 9 9 1 9 9 1 9 7 13 0 13 12 1 12 1 9 9 1 9 0 13 15 9 9 2 1 9 7 13 9 0 1 9 13 1 12 7 12 9 7 1 9 0 0 13 1 9 0 1 9 9 15 13 1 9 9 2
46 7 13 9 7 9 9 0 7 14 13 9 9 1 9 9 0 0 2 1 9 7 9 9 9 9 15 0 1 9 1 9 0 1 9 0 7 9 9 1 9 9 1 9 9 9 2
76 13 15 1 9 9 9 0 1 9 9 9 2 9 2 9 0 9 9 0 15 14 13 9 1 0 1 9 9 15 1 0 9 2 7 13 0 1 9 9 9 15 14 13 9 1 9 0 0 9 1 9 0 2 7 9 1 9 9 7 9 2 7 1 9 9 0 1 9 9 7 9 9 7 9 0 2
38 7 9 9 0 13 0 1 9 15 15 13 0 9 2 3 13 14 13 15 1 9 2 7 3 9 0 1 9 0 13 9 9 13 9 15 9 12 2
110 7 13 9 9 9 0 1 9 9 9 1 9 0 9 2 7 13 9 7 15 14 13 1 9 9 7 13 1 9 1 9 9 2 7 13 9 7 15 14 13 1 9 9 0 9 1 9 0 7 13 9 9 1 9 15 1 9 9 9 7 9 9 2 15 13 7 15 2 9 2 0 1 9 0 7 1 9 15 13 9 9 7 9 9 3 2 7 13 9 0 0 1 9 1 9 1 0 1 9 9 0 9 9 7 13 1 15 10 9 2
52 7 13 1 9 9 7 14 13 9 9 0 1 9 9 0 7 4 9 9 9 9 15 2 7 13 9 9 9 9 12 12 9 0 7 7 13 9 15 1 9 0 15 13 9 15 1 9 0 12 12 9 2
43 7 1 9 12 13 9 0 1 9 0 7 0 1 9 0 1 9 0 1 9 0 7 0 9 1 9 9 1 9 9 9 0 1 9 9 15 14 13 9 1 9 15 2
71 7 1 9 9 9 0 9 1 9 9 13 1 9 9 0 1 9 0 0 15 13 1 9 0 1 0 9 0 1 9 9 1 9 0 7 0 2 7 13 9 9 0 0 15 13 15 9 1 12 9 13 12 9 7 12 9 0 1 9 7 9 13 1 9 12 12 9 0 9 12 2
51 7 13 9 9 9 0 9 1 7 15 1 9 0 1 9 0 7 9 12 1 12 1 9 9 3 13 9 9 0 0 7 1 3 13 9 9 1 1 15 9 9 9 0 15 13 9 1 0 1 15 2
79 7 13 9 7 13 9 9 0 1 9 9 0 1 9 0 1 9 9 9 0 1 12 12 9 1 9 9 7 9 9 14 13 0 9 1 9 9 9 1 9 0 7 14 13 1 9 9 2 9 1 7 15 14 13 9 1 9 9 0 1 0 9 15 13 7 9 9 14 13 0 7 1 9 0 1 9 0 9 2
173 7 13 9 0 1 9 0 1 9 0 12 12 9 9 12 2 13 9 9 7 9 0 7 9 9 7 9 7 9 7 13 9 9 9 9 0 1 9 12 12 9 0 7 15 0 1 9 1 9 9 8 7 1 9 9 15 13 15 9 9 1 9 9 15 13 9 15 1 9 9 0 2 1 13 9 9 0 1 15 7 13 9 0 1 9 7 0 1 9 8 8 1 9 0 7 13 0 9 9 1 10 9 1 12 9 7 13 0 9 9 1 9 8 1 9 12 12 9 7 9 0 12 12 9 7 9 1 12 7 12 12 9 1 9 9 1 9 9 15 2 14 9 8 8 8 7 14 13 9 0 9 9 7 9 9 9 0 2 7 1 9 9 9 1 9 13 9 1 9 12 12 9 2
136 1 9 0 13 9 1 9 9 0 13 1 9 15 13 0 7 13 1 15 9 9 9 2 7 3 9 0 0 0 2 7 13 9 9 9 1 9 8 8 9 7 9 13 9 0 13 1 12 12 9 1 15 12 12 1 9 2 0 1 7 15 14 13 1 9 0 1 9 7 9 9 0 2 7 13 7 9 13 1 9 0 1 9 9 0 7 9 15 1 9 7 13 9 15 1 12 9 7 13 9 1 9 9 15 7 14 13 9 15 1 9 9 7 1 9 9 15 13 9 9 9 9 9 9 9 0 7 9 9 9 1 9 0 1 9 2
22 9 14 13 9 15 7 9 13 9 2 9 2 9 0 1 9 2 9 9 7 9 2
2 8 8
38 13 9 0 2 1 9 0 2 1 9 9 0 9 1 2 9 9 7 9 2 1 9 9 0 1 9 7 15 13 12 12 9 2 12 12 9 2 2
36 13 9 0 7 15 14 13 9 2 9 9 7 9 2 9 1 9 15 0 2 7 13 1 12 9 0 15 2 9 8 2 15 13 9 8 2
35 7 13 9 1 9 9 1 9 9 1 9 9 9 1 9 9 9 15 13 15 2 0 1 9 0 2 7 13 1 15 9 0 1 9 2
29 7 13 9 9 8 8 7 9 10 9 14 13 1 9 13 1 15 9 9 9 15 13 0 1 9 9 9 0 2
88 7 13 9 0 1 9 2 1 9 2 9 2 7 2 9 2 7 2 9 0 2 2 9 9 1 9 9 1 9 1 9 9 7 9 9 1 9 7 9 9 9 1 9 2 7 10 9 14 13 9 13 9 9 9 1 9 9 1 9 9 9 15 2 7 13 9 9 1 9 7 13 12 12 9 2 15 13 7 15 14 13 1 0 9 13 15 9 2
58 7 13 9 9 0 9 12 12 9 1 9 1 9 0 1 9 9 9 2 7 13 0 1 12 12 9 9 9 2 7 14 13 15 9 0 9 9 0 7 13 9 9 15 14 13 1 9 1 12 12 1 12 12 13 0 1 9 2
47 7 13 7 13 9 1 9 0 9 9 1 9 15 13 1 9 9 9 1 15 2 1 9 1 7 9 13 0 1 9 9 2 15 13 7 9 0 14 13 9 0 1 9 9 7 9 2
59 7 13 9 0 1 9 1 2 9 2 1 9 9 1 9 1 9 2 0 1 7 15 13 9 1 9 2 7 9 13 9 0 9 1 9 0 13 1 12 12 9 2 7 10 9 13 1 12 12 1 9 7 9 9 15 1 12 9 2
46 7 13 9 7 15 1 9 9 10 7 14 9 1 9 9 9 9 0 15 13 1 12 12 9 7 1 3 14 9 1 9 0 0 9 7 7 15 14 13 9 0 1 9 9 0 2
51 7 13 8 7 9 13 9 0 1 9 9 9 0 0 15 13 1 12 9 1 9 9 7 9 1 9 0 1 9 9 1 12 12 9 0 1 9 1 9 2 1 12 12 13 9 15 0 1 0 9 2
22 7 14 13 9 15 1 9 0 9 1 9 9 9 0 0 1 9 9 9 0 0 2
10 9 2 9 9 1 9 0 9 1 11
57 13 1 9 0 7 15 13 9 1 9 9 0 1 9 9 0 2 8 8 2 2 7 0 2 8 2 2 7 0 2 8 2 13 9 7 9 9 1 0 9 0 1 9 9 7 8 8 8 8 1 9 9 1 9 11 0 2
48 7 13 9 10 14 13 15 9 0 1 12 12 9 2 7 13 9 12 12 9 1 9 1 9 0 2 8 2 7 12 12 9 0 1 8 0 13 1 9 1 9 1 12 9 0 1 9 2
78 1 9 0 2 13 9 9 8 8 9 9 9 2 9 0 1 9 0 2 2 8 2 2 7 15 9 9 0 13 9 12 1 9 9 1 9 9 9 1 9 2 8 2 2 1 9 1 9 1 9 0 1 9 2 8 2 13 9 15 12 12 9 2 1 9 9 2 8 2 1 9 0 1 9 9 9 0 2
31 9 2 9 2 1 9 8 8 13 9 15 9 1 9 9 2 9 1 9 13 9 9 7 9 13 9 1 2 9 9 2
67 13 9 0 1 9 9 3 1 9 9 9 1 9 2 9 9 0 2 7 2 9 9 0 2 2 9 2 7 1 9 1 9 0 7 9 9 0 15 13 15 9 8 8 2 7 13 9 0 9 15 1 7 13 9 15 13 9 9 1 9 2 9 0 0 1 9 2
41 7 13 9 0 0 9 9 1 2 9 9 0 2 2 0 2 9 2 1 9 9 1 9 1 9 0 2 7 0 1 7 9 2 14 13 1 9 1 9 2 2
71 7 13 9 8 8 1 9 3 1 9 0 8 1 9 7 9 2 7 13 9 1 9 1 9 9 1 9 0 2 1 9 15 13 0 2 7 13 9 0 1 11 1 2 9 2 7 8 0 9 1 9 0 2 0 2 7 13 7 15 13 9 15 7 13 1 9 1 9 9 9 2
73 7 13 9 9 1 9 0 7 0 1 9 9 0 0 1 9 1 9 2 7 13 2 9 8 8 9 2 2 7 13 9 8 8 8 2 9 0 1 9 9 7 2 9 1 9 15 1 9 2 7 7 9 9 2 13 9 2 2 7 13 7 8 13 2 9 1 9 9 1 0 9 2 2
2 9 9
51 7 13 9 7 9 9 13 1 9 9 7 9 9 1 9 2 1 9 2 9 9 2 9 7 13 3 1 9 2 9 2 7 2 9 0 2 7 1 9 9 9 7 9 9 2 7 13 0 1 9 2
99 7 13 9 2 8 8 2 1 9 0 0 0 9 15 2 8 2 1 9 1 9 2 7 13 7 2 9 9 13 1 10 9 15 13 15 9 9 9 15 7 9 14 13 2 9 2 7 13 15 2 2 7 13 7 2 8 9 13 1 9 9 8 8 9 9 0 7 13 9 8 9 2 7 13 1 15 9 9 9 7 13 9 7 13 9 15 1 9 2 7 13 7 8 13 1 10 9 2 2
56 7 13 9 15 13 9 9 15 1 2 9 9 1 9 10 13 9 9 0 2 2 7 13 2 7 9 13 1 9 9 7 14 13 1 0 9 1 9 7 14 1 9 9 7 13 1 9 0 1 9 9 7 9 9 2 2
31 7 13 2 8 2 1 2 9 9 1 9 9 1 9 9 7 9 2 7 13 9 15 9 9 7 13 15 1 9 2 2
70 7 13 7 2 9 13 9 1 9 7 13 9 1 9 2 15 13 1 9 15 2 2 0 1 7 2 9 13 1 9 9 1 9 0 2 2 7 13 7 9 2 13 2 1 9 9 9 2 9 7 9 1 9 2 2 0 1 7 2 9 14 13 1 9 1 1 10 9 2 2
64 7 13 9 0 7 9 1 2 8 2 13 3 9 9 1 9 9 7 13 12 1 9 1 9 1 9 9 1 9 7 9 0 13 9 1 9 1 9 2 7 13 7 8 2 13 9 1 9 1 9 7 13 9 1 15 7 9 9 8 8 8 0 2 2
69 7 2 8 2 13 10 9 2 7 13 8 8 2 9 9 9 1 9 9 1 9 2 8 8 2 7 2 9 8 0 2 2 0 1 9 15 2 9 1 9 0 2 2 7 13 9 9 9 9 9 8 8 7 2 9 14 13 1 1 15 2 2 1 15 14 13 9 9 2
64 7 13 9 2 8 2 1 9 0 9 1 2 9 9 0 9 15 9 9 9 2 7 13 7 9 9 9 13 9 1 9 0 1 9 15 2 1 1 13 9 1 9 7 2 1 9 9 9 0 7 9 9 1 9 1 9 2 14 7 13 9 9 2 2
49 7 13 2 9 8 8 8 2 9 0 1 2 9 2 7 2 9 9 0 2 13 1 9 0 9 0 9 0 7 9 0 1 9 9 1 9 9 8 8 1 9 15 9 1 9 9 9 9 2
48 7 13 2 8 2 1 9 0 9 15 7 13 9 13 9 0 2 7 15 13 7 9 9 13 1 9 9 2 2 7 13 9 1 9 9 1 9 1 1 2 9 9 1 9 9 9 2 2
24 8 2 8 1 9 9 9 12 2 0 13 9 1 9 7 9 13 1 9 15 1 0 0 9
9 8 8 2 8 8 2 8 8 8
49 13 8 3 9 9 9 0 1 0 1 9 13 1 9 0 2 7 14 13 9 9 0 11 8 9 0 13 9 15 2 7 15 8 1 7 2 0 9 14 13 9 0 1 15 8 8 8 2 2
81 7 7 13 9 7 9 0 7 0 1 9 9 0 1 9 0 2 13 9 0 1 9 0 8 8 9 1 9 1 2 9 2 7 9 0 13 1 9 9 9 9 12 1 8 0 1 9 9 1 2 9 0 2 2 7 13 9 9 0 8 8 9 9 9 9 1 9 1 9 9 9 8 8 1 9 9 0 1 9 9 2
139 7 13 8 1 9 3 7 9 14 13 0 1 9 7 15 14 13 1 9 9 15 2 7 13 9 8 8 9 1 9 8 8 2 13 7 15 13 1 2 9 0 1 9 2 2 7 13 9 0 15 13 15 9 0 1 9 0 8 8 1 9 15 8 2 7 13 9 1 9 1 2 9 2 7 9 0 1 0 2 14 13 9 0 2 7 13 15 9 2 0 1 7 9 15 14 13 2 9 1 10 13 15 8 8 2 0 2 7 15 15 1 8 8 2 2 7 13 7 9 2 13 7 14 13 13 1 9 0 7 9 7 9 2 7 13 9 0 2 2
76 7 13 9 0 7 0 1 9 8 1 9 2 9 9 0 0 1 9 2 7 13 8 7 2 0 9 0 7 9 0 1 9 0 2 14 13 15 1 9 15 2 2 7 13 7 9 15 2 14 13 1 9 0 7 9 0 2 7 9 9 0 14 13 9 9 2 2 7 13 1 9 9 1 9 9 2
125 7 1 9 15 1 9 14 13 8 9 0 13 0 2 7 13 2 2 9 9 0 2 2 7 13 1 7 2 9 1 9 0 2 7 9 1 15 13 0 2 7 13 9 7 0 9 14 13 15 0 2 7 14 13 15 0 2 2 7 1 9 15 9 0 2 13 9 9 0 7 9 14 13 1 9 2 7 7 1 9 9 15 2 14 13 1 9 15 7 13 2 2 7 13 1 9 9 0 0 1 9 9 9 0 8 8 9 9 0 15 2 13 3 1 9 9 1 9 9 1 9 9 0 2 2
52 7 13 1 9 15 7 9 7 9 14 13 1 9 8 8 9 2 0 2 8 8 1 9 9 2 1 7 15 2 0 9 2 2 7 13 7 9 2 13 9 0 1 9 9 1 9 7 9 9 0 2 2
69 1 9 15 13 9 7 9 1 9 9 0 1 9 0 7 13 9 0 1 9 0 1 9 9 1 9 9 0 1 9 9 1 9 7 9 7 13 1 2 9 0 2 15 13 1 9 9 0 12 7 2 13 1 9 1 7 9 9 0 2 9 9 1 9 0 2 0 2 2
84 7 13 9 8 9 1 9 1 2 9 2 1 9 15 1 9 9 0 1 9 15 1 9 8 2 7 13 9 1 9 9 0 15 13 1 9 9 1 9 9 0 2 8 2 8 2 8 2 9 1 9 0 2 7 13 2 2 9 7 14 13 9 12 9 15 8 8 7 8 1 15 8 8 7 8 15 7 15 8 8 9 15 2 2
72 7 13 9 9 0 8 8 13 3 1 9 15 1 9 0 1 9 0 7 0 1 9 0 8 8 7 9 9 8 14 13 14 1 2 9 0 1 9 2 2 7 1 9 0 13 9 9 0 9 8 8 7 9 0 2 14 13 9 9 9 2 2 7 7 15 13 1 2 9 0 2 2
274 1 9 9 15 13 9 8 8 1 9 15 1 9 2 1 9 9 9 9 0 1 9 0 0 2 7 13 9 9 0 8 8 15 13 15 9 8 8 9 3 1 9 8 1 2 9 2 7 9 9 8 8 7 14 8 1 9 1 8 13 2 7 14 8 1 8 7 13 1 9 15 0 2 2 7 13 7 2 9 0 0 1 9 0 1 9 9 7 9 7 9 0 7 0 7 0 2 2 7 1 9 8 9 9 9 15 13 15 9 8 1 9 9 0 7 0 13 8 2 2 3 9 0 13 0 9 0 1 9 9 1 9 1 9 0 2 7 1 9 15 9 9 9 7 9 1 9 0 2 2 7 13 2 2 8 13 8 8 7 13 9 0 1 9 9 9 2 0 7 8 13 1 10 9 9 9 9 2 8 8 13 1 9 0 2 7 10 9 2 7 1 9 9 10 8 8 1 9 2 14 13 7 3 9 1 9 7 9 0 1 9 9 9 1 9 9 8 2 2 7 13 2 2 8 9 14 13 7 13 1 15 9 1 8 1 9 9 0 13 1 15 9 0 9 0 1 9 9 8 2 2 7 13 9 9 0 1 9 0 1 2 9 9 9 0 1 9 9 0 1 9 9 2 2
17 9 2 9 13 2 0 1 9 2 1 9 9 9 9 0 1 9
2 8 8
49 13 9 0 3 9 15 13 0 1 9 9 15 13 1 2 9 0 1 9 2 13 15 1 9 1 9 1 9 9 9 0 1 9 0 7 9 15 9 1 9 2 8 8 2 7 2 8 2 2
95 7 13 9 9 9 9 9 9 1 9 1 9 9 9 7 9 8 8 9 9 0 1 9 1 9 12 12 9 2 12 12 9 2 1 9 9 0 15 14 13 1 9 2 8 2 8 2 8 2 2 9 1 0 9 0 2 9 2 9 12 2 7 13 8 2 2 14 9 14 13 9 9 0 1 9 7 1 9 9 7 9 15 14 13 1 0 1 9 13 15 9 1 9 0 2
78 7 1 0 9 9 13 9 1 9 9 1 2 9 2 7 9 15 13 15 2 0 1 9 2 14 13 15 13 15 9 7 7 15 1 15 13 12 12 9 9 12 1 15 13 12 12 9 9 15 7 13 9 9 12 9 7 14 13 9 3 12 12 9 0 1 9 9 12 9 3 7 0 7 13 9 9 15 2
42 7 13 9 1 7 9 8 8 9 0 8 8 8 9 0 2 7 15 13 9 1 9 2 0 7 9 9 1 13 0 1 9 9 9 15 1 9 9 15 9 0 2
21 7 13 9 13 9 0 1 9 9 9 0 1 9 0 1 9 9 9 9 0 2
19 7 13 9 9 1 15 1 9 9 9 9 9 0 9 9 9 9 9 2
86 7 13 7 13 9 0 9 1 9 7 9 9 9 0 13 1 9 12 1 12 0 2 7 13 9 12 1 12 12 13 9 12 1 12 12 7 13 1 12 9 12 7 13 0 1 12 12 9 2 7 1 9 9 9 7 9 14 13 9 1 12 12 9 9 12 7 12 12 9 12 15 13 7 9 1 9 9 14 13 12 12 9 1 12 9 2
17 9 1 9 9 9 2 9 13 9 9 0 1 9 15 13 9 15
2 8 8
26 13 9 9 9 0 0 8 8 7 9 13 9 0 1 9 9 1 9 0 1 9 1 9 9 9 2
19 7 13 1 9 1 9 3 7 9 13 9 1 9 1 9 1 0 9 2
36 7 13 7 9 9 0 1 9 9 9 15 13 9 15 0 1 9 7 7 9 0 9 1 10 9 0 1 9 9 9 1 9 7 9 9 2
37 7 13 9 9 0 1 9 1 9 1 9 9 1 9 0 2 9 7 9 13 1 9 7 9 9 7 9 7 9 7 9 7 9 0 7 0 2
57 7 13 1 7 2 0 1 9 2 13 1 9 12 9 2 7 13 2 0 1 9 0 2 9 0 7 2 0 1 9 0 7 0 2 12 9 7 2 0 1 9 9 2 12 9 7 13 2 0 1 9 0 7 0 9 2 2
57 7 13 2 0 1 9 0 2 1 9 0 1 9 0 1 9 2 7 13 12 9 1 1 15 12 9 1 9 9 2 7 13 2 9 1 9 7 9 2 12 9 1 9 7 13 2 0 1 9 7 9 7 9 2 12 9 2
40 7 13 8 7 15 13 0 9 9 15 14 13 1 9 9 2 9 0 1 9 7 9 7 9 2 1 9 9 0 1 2 9 9 1 9 2 2 8 2 2
25 7 13 7 9 1 9 9 0 0 1 9 9 0 1 9 2 9 8 8 2 13 9 15 0 2
53 1 15 14 13 0 9 0 1 9 2 9 8 2 1 9 1 9 0 1 9 2 8 2 0 7 1 9 9 9 15 13 9 1 15 1 9 9 9 7 9 9 1 9 0 1 9 7 9 1 9 9 9 2
92 7 13 10 9 1 9 15 13 1 15 9 9 1 9 9 2 1 0 15 9 9 9 1 9 9 9 9 0 15 13 9 15 1 9 13 9 7 1 9 1 9 2 9 1 7 9 13 9 1 9 9 0 0 13 15 9 2 7 7 9 15 13 15 9 0 1 9 9 9 0 13 14 13 0 7 0 1 9 9 0 2 7 1 7 13 1 9 9 9 0 0 2
52 7 13 9 1 9 9 2 1 9 7 9 13 1 9 9 0 2 15 13 7 9 9 1 9 0 1 9 9 9 9 14 13 1 9 9 15 7 1 7 13 9 0 1 9 7 7 3 9 9 1 9 2
12 9 2 12 12 9 9 9 9 9 9 7 9
71 9 2 2 9 2 2 13 0 0 0 1 7 13 9 9 15 0 1 9 9 7 9 7 13 9 9 9 9 1 9 9 9 2 7 13 9 0 1 2 9 2 7 9 14 13 0 1 0 7 9 9 8 8 1 9 1 9 10 9 15 13 9 15 9 12 1 12 1 9 9 2
49 7 13 9 13 1 9 2 9 2 9 1 9 2 8 7 9 13 1 7 9 13 2 7 13 9 7 9 9 13 1 9 9 0 1 9 9 9 15 13 9 15 1 9 12 12 9 1 0 2
52 7 13 9 9 9 8 8 1 9 1 2 9 2 1 9 9 0 1 9 8 7 9 15 1 9 9 9 2 7 13 1 9 9 0 1 9 9 7 9 1 9 15 13 1 15 7 9 15 13 9 15 2
49 7 13 0 1 9 1 9 9 0 9 1 12 9 0 13 1 9 10 9 7 9 9 0 9 1 9 9 0 1 9 12 0 2 0 1 9 9 9 9 9 1 9 9 9 9 7 9 0 2
34 7 13 8 9 9 9 1 9 9 0 7 9 9 0 1 9 0 1 9 9 7 9 9 1 9 7 9 9 0 7 9 9 9 2
77 1 9 9 15 13 9 0 1 9 9 7 9 9 9 7 1 12 1 12 1 9 13 9 7 9 0 1 9 15 13 9 9 9 1 9 1 9 9 7 9 9 1 12 1 12 1 0 7 9 9 9 1 9 2 7 3 9 9 0 0 1 15 13 9 15 1 9 0 7 13 12 1 12 9 1 12 2
13 9 2 9 2 8 2 1 9 9 0 1 9 0
34 13 2 9 1 9 2 9 9 2 8 2 0 1 9 0 1 9 9 0 1 9 0 15 14 13 9 1 9 0 2 9 2 12 2
40 7 13 9 9 9 9 8 8 2 1 9 0 7 2 8 14 13 1 9 1 9 9 0 1 8 7 1 15 7 13 1 9 9 7 9 0 1 9 2 2
36 7 13 7 9 0 1 9 0 14 13 7 13 1 15 9 13 9 1 15 1 9 9 7 9 7 9 9 1 9 13 1 9 0 1 9 2
13 9 2 2 9 2 13 9 12 1 12 1 9 9
84 9 2 2 9 2 2 13 9 2 9 2 1 9 0 1 9 13 13 9 15 13 9 9 0 9 9 1 9 9 2 7 13 10 9 13 1 9 9 12 1 9 9 9 0 2 7 13 9 1 9 9 1 7 9 2 9 2 13 12 1 12 1 9 9 9 7 15 1 9 15 1 9 9 1 9 13 1 12 7 12 1 12 0 2
79 7 13 9 9 0 1 9 1 9 9 9 0 1 9 0 1 1 9 9 1 9 2 7 13 10 9 9 0 1 9 9 9 0 1 9 9 0 9 13 9 1 0 9 1 9 9 1 9 7 9 9 15 1 9 9 0 1 10 9 2 7 13 9 0 1 9 9 9 0 0 1 9 9 9 15 1 9 0 2
10 9 13 9 9 9 1 9 12 12 9
2 8 8
52 13 9 0 9 12 9 0 0 1 9 9 9 1 9 9 9 13 9 15 1 9 0 7 0 7 0 1 9 9 0 1 7 13 9 15 1 9 2 7 13 9 10 9 12 12 9 2 12 12 9 2 2
76 7 13 9 9 8 8 1 2 9 2 7 9 15 9 13 1 9 1 9 9 8 8 7 13 1 9 1 7 13 9 15 1 9 8 7 8 1 9 9 9 1 9 2 7 9 13 9 9 1 9 8 8 8 1 9 8 2 9 1 9 9 2 11 2 8 2 8 2 14 13 1 9 9 0 0 2
38 7 13 8 7 15 13 9 9 9 0 1 9 8 8 8 1 9 9 0 2 14 13 15 2 7 13 9 9 8 2 8 8 8 2 8 1 9 2
85 7 13 1 7 15 13 0 9 9 9 7 9 0 1 9 9 8 9 9 1 9 9 0 1 15 2 7 13 7 15 14 13 9 9 12 9 0 8 8 9 1 9 9 9 9 0 2 7 13 7 9 9 9 0 9 1 9 8 8 14 13 1 9 1 9 0 7 7 9 0 1 15 14 13 0 7 14 13 9 1 9 0 7 0 2
72 7 1 9 1 9 2 13 8 7 9 13 1 9 9 1 9 9 12 9 1 9 9 9 9 7 9 9 7 9 9 2 0 7 15 14 13 9 9 9 1 9 0 0 1 9 0 7 0 7 7 15 14 0 1 9 1 9 9 1 10 9 9 7 9 13 1 9 9 1 9 0 2
3 9 8 8
15 8 8 2 8 8 0 1 8 13 8 3 1 12 9 2
53 9 1 9 8 0 8 2 8 1 0 8 8 8 7 9 0 2 8 13 1 15 9 15 0 1 9 9 0 1 9 0 1 8 2 7 1 7 13 1 8 8 8 13 0 8 8 8 8 2 9 7 9 2
41 9 15 0 0 15 13 1 9 12 13 9 15 2 9 9 2 8 8 2 7 13 1 9 9 0 15 14 13 8 8 1 15 1 0 8 2 0 13 9 15 2
100 8 8 8 8 8 8 8 8 8 1 9 1 9 2 8 8 1 9 2 13 15 1 9 0 2 15 13 8 8 8 2 7 13 13 9 1 9 8 8 8 1 9 8 8 2 7 9 8 8 9 8 8 2 9 15 0 2 0 7 0 7 1 1 2 13 8 1 9 0 1 15 13 1 9 12 2 7 13 10 9 8 8 0 13 9 13 1 1 15 8 13 8 7 14 13 1 9 8 8 2
32 7 1 15 1 8 8 9 9 1 0 15 9 9 0 8 2 8 8 2 7 13 7 15 1 0 8 8 13 15 10 9 2
52 13 8 8 0 1 9 0 8 8 8 7 13 9 2 9 2 1 9 12 2 9 8 8 1 9 7 9 7 9 1 0 7 9 2 7 1 15 11 8 2 8 2 9 8 8 8 7 1 15 2 2 2
38 7 7 13 8 1 9 15 13 1 9 2 8 2 9 1 9 7 15 13 7 13 1 9 0 2 0 1 9 8 7 9 0 2 9 1 9 0 0
16 1 9 0 1 9 8 2 1 9 0 1 2 9 9 2 0
3 8 8 8
127 1 13 9 9 9 1 9 0 7 15 13 9 1 9 15 7 9 9 15 7 9 0 1 15 7 9 15 1 9 0 2 7 3 9 15 7 9 15 1 9 1 9 15 0 2 7 14 9 7 10 9 13 9 1 9 9 1 9 10 9 7 9 9 15 1 9 0 7 0 2 7 1 9 15 13 9 9 1 9 0 1 9 9 2 9 0 0 1 9 0 1 8 1 9 8 15 13 1 9 9 2 9 2 0 2 7 13 10 9 9 0 1 9 15 1 9 9 0 7 15 9 0 7 9 0 0 2
99 7 14 8 0 7 8 7 9 1 9 8 0 1 9 9 8 8 0 2 8 8 0 13 1 9 9 0 1 9 9 0 1 9 9 1 9 0 8 8 9 0 1 9 2 9 1 9 0 7 1 9 0 7 3 9 1 9 9 1 9 8 8 7 9 9 7 9 9 7 9 9 0 8 8 8 8 1 9 0 8 9 2 7 7 13 1 9 0 2 9 0 1 9 0 8 8 8 8 2
23 1 9 13 8 0 1 9 10 9 8 8 9 1 8 9 7 7 1 0 1 9 8 2
107 7 1 8 9 9 9 9 9 0 1 9 1 9 2 14 8 8 8 1 9 1 9 9 8 8 1 9 2 8 8 9 9 9 8 8 9 1 9 8 8 1 9 0 2 7 14 8 15 13 1 9 9 15 13 7 15 14 13 2 7 7 9 1 10 9 8 8 8 8 8 1 9 1 15 0 1 9 10 13 1 1 2 8 2 2 7 9 14 13 9 1 9 2 7 7 9 9 7 9 1 9 15 14 13 13 9 2
55 7 1 0 3 9 9 0 1 15 8 2 14 7 9 15 8 1 10 9 10 1 9 9 1 9 8 1 9 9 15 13 9 12 8 8 8 8 8 8 8 1 9 9 0 8 8 8 8 8 9 15 1 9 0 2
165 8 8 8 13 9 0 1 9 8 0 2 9 15 13 1 9 1 9 15 7 9 15 0 2 7 1 9 1 9 9 0 1 10 9 2 8 7 9 7 9 0 0 13 0 1 9 8 2 7 13 9 9 0 1 8 1 9 0 7 0 2 7 13 1 9 1 9 1 9 9 1 9 9 9 9 0 0 0 1 9 0 1 9 1 9 9 12 9 0 7 0 7 0 7 0 2 7 13 1 9 15 9 9 15 13 1 9 15 9 0 15 13 9 0 1 9 1 9 9 15 13 1 9 2 7 13 1 9 9 8 0 7 9 0 2 8 0 2 13 1 9 0 1 9 9 9 2 7 13 10 9 0 1 9 15 1 9 9 0 0 0 1 9 0 2
34 7 13 9 9 1 9 0 0 1 9 8 0 8 8 8 8 2 7 9 9 9 7 9 1 9 8 7 9 9 0 1 10 9 2
49 7 13 9 9 9 9 0 8 8 8 1 9 15 8 9 1 9 9 0 1 9 1 9 0 1 9 9 7 3 1 9 9 15 13 1 15 9 0 1 9 0 7 9 9 0 1 9 0 2
45 7 1 9 9 0 0 1 9 13 9 0 1 9 0 12 1 8 1 8 7 13 10 9 8 8 9 0 8 8 9 9 0 1 9 0 9 9 0 0 7 15 13 1 15 2
19 12 2 9 9 0 1 9 0 7 9 15 9 1 9 9 0 1 9 2
15 12 2 9 1 9 8 0 7 0 1 9 9 0 0 2
21 12 2 9 1 9 9 1 9 0 8 8 7 9 8 8 8 8 8 1 15 2
23 12 2 9 1 9 9 0 1 9 9 9 9 1 9 9 8 0 7 1 9 9 9 2
42 12 2 9 9 9 0 1 9 15 1 9 7 9 0 8 9 0 1 9 8 8 8 8 8 1 9 0 7 13 8 8 1 9 1 9 2 8 2 1 9 8 2
24 8 1 9 1 9 2 8 0 2 1 9 12 12 9 1 9 7 9 1 8 9 1 8 2
22 1 9 7 14 9 9 0 1 9 9 13 0 1 15 1 9 7 15 1 9 9 2
26 8 2 9 7 9 0 1 9 9 7 9 0 1 9 9 8 8 9 1 9 0 8 8 0 0 2
45 0 2 8 9 9 0 0 2 13 9 0 1 9 9 1 9 0 7 9 9 15 2 7 13 3 8 2 7 1 0 7 15 0 1 8 8 8 7 9 9 8 8 0 8 2
24 0 2 8 9 9 0 8 8 8 1 9 1 9 9 0 8 8 9 1 15 1 10 9 2
130 3 15 13 9 15 1 9 13 7 9 0 1 9 9 9 12 13 9 1 9 0 9 12 2 7 9 10 9 13 1 9 15 1 9 8 1 9 9 9 0 2 14 9 1 9 9 8 8 8 8 8 13 9 15 1 9 7 9 7 9 1 8 8 1 8 0 2 7 15 13 15 1 9 8 8 7 9 1 9 9 9 0 2 8 8 7 15 1 0 9 1 9 1 9 9 7 9 1 9 10 9 1 9 0 1 9 3 1 8 8 8 8 1 9 9 15 14 13 1 15 8 1 9 8 8 1 0 9 0 2
18 8 9 0 1 9 0 1 9 9 2 9 9 8 0 1 9 9 2
5 0 9 2 9 2
2 9 8
83 13 9 12 1 9 2 9 2 0 9 0 1 9 15 9 9 8 8 2 7 13 9 9 1 11 8 1 2 9 9 1 9 2 8 8 0 8 8 9 0 2 7 13 8 9 9 9 1 15 13 9 9 0 2 7 13 9 9 1 9 8 8 1 9 8 2 7 13 8 8 9 2 7 13 8 8 8 7 13 1 8 9 2
51 7 1 9 9 15 13 8 8 9 9 1 9 9 9 8 11 8 2 7 13 1 7 15 13 1 9 10 9 1 9 7 9 13 15 13 9 0 9 1 15 1 9 15 1 9 9 1 9 8 8 2
72 7 1 9 9 13 8 9 9 0 8 8 8 13 15 2 8 8 0 1 9 7 15 13 1 15 9 0 1 15 9 0 2 1 15 9 9 1 9 15 8 8 8 0 1 15 7 15 15 13 9 9 1 15 2 7 9 8 9 9 1 9 9 7 9 8 0 1 9 0 9 15 2
116 7 13 9 1 9 9 7 9 12 8 0 15 2 9 9 1 9 0 2 1 9 8 8 1 9 9 2 9 9 2 1 9 0 8 8 2 7 13 9 8 1 10 9 9 9 0 1 8 0 1 1 9 0 7 9 9 7 9 2 7 13 8 8 9 1 9 8 8 7 15 7 13 13 1 9 9 2 7 13 8 1 9 9 9 8 8 1 9 9 0 0 8 8 9 0 8 2 7 1 9 15 13 8 8 8 8 8 1 9 2 8 8 8 1 9 2
47 7 13 8 8 9 1 9 0 8 13 1 15 8 9 9 1 9 8 2 7 9 9 8 0 1 9 1 9 2 7 13 8 9 1 9 9 9 8 8 8 1 9 13 15 8 8 2
2 9 9
31 9 13 8 9 1 9 1 9 9 2 13 9 0 1 9 7 15 13 9 8 8 7 15 0 1 9 0 2 8 8 2
18 2 13 9 0 0 13 9 9 1 9 8 1 9 7 13 1 9 2
29 2 13 9 9 0 12 9 1 9 8 1 9 2 7 13 7 15 13 1 9 8 8 0 2 7 14 13 9 2
40 2 13 1 9 0 1 1 9 2 7 13 9 9 0 7 9 14 13 0 1 9 1 9 7 13 9 1 0 2 7 7 1 9 1 9 0 1 9 15 2
49 2 13 9 0 1 9 12 9 1 9 1 8 8 2 7 14 13 9 9 7 9 9 13 1 15 8 2 8 2 9 1 9 1 9 12 15 13 1 9 0 1 9 15 1 15 13 8 8 2
108 8 8 7 8 1 9 9 8 8 2 7 9 9 13 2 8 8 9 0 2 7 14 8 9 3 1 10 9 2 8 8 0 13 9 0 1 9 0 2 1 9 15 1 9 9 1 9 12 9 0 1 7 13 8 8 1 9 8 8 2 9 7 9 9 15 13 1 9 8 8 2 0 2 1 9 0 2 1 8 8 0 13 12 8 0 8 8 8 8 2 1 7 13 9 2 7 9 2 8 2 0 13 9 9 1 8 8 2
45 14 8 8 8 9 15 0 2 8 8 9 0 1 15 13 0 3 2 7 9 13 9 9 0 0 2 15 13 9 2 8 2 13 1 7 9 0 13 8 9 1 9 8 8 2
56 8 1 9 9 0 7 9 9 0 2 0 7 0 2 1 9 0 0 1 0 2 8 8 0 0 8 1 9 2 8 8 8 7 3 9 7 14 13 3 9 1 9 0 7 1 9 9 15 2 7 9 9 9 10 8 2
80 7 7 9 7 13 9 0 9 0 2 7 14 0 2 8 8 9 0 2 13 8 13 9 7 9 9 8 8 7 9 9 8 8 13 9 0 1 9 9 8 8 2 7 13 9 9 9 8 1 9 9 1 9 9 7 9 9 1 9 8 9 2 7 13 9 9 9 1 9 7 8 13 9 9 0 9 9 9 0 2
27 9 14 13 0 7 8 7 8 13 7 8 9 7 9 9 14 13 9 9 2 7 14 13 1 9 0 2
81 1 15 8 8 14 13 1 9 1 9 7 9 2 8 8 0 14 13 9 0 9 2 8 8 1 9 15 10 9 0 1 9 0 15 13 9 15 1 9 9 8 2 7 7 13 8 14 13 9 1 9 9 2 7 1 9 8 13 8 9 1 0 7 12 1 9 15 13 9 7 15 13 8 8 7 13 7 15 9 0 2
53 1 9 14 13 3 9 0 0 1 9 9 15 1 9 2 7 1 9 7 9 0 0 1 10 9 13 15 9 0 8 1 9 8 2 8 8 3 12 9 8 8 2 8 8 1 0 2 14 7 9 15 0 2
79 9 9 15 13 10 9 15 13 1 15 9 15 7 15 13 1 9 15 2 7 9 0 8 8 1 9 2 1 9 2 7 1 9 0 9 15 2 7 9 0 1 9 13 15 1 8 9 15 2 7 13 1 9 15 9 7 13 15 2 7 0 1 15 7 15 13 9 1 9 9 13 9 1 15 9 0 1 9 2
95 14 13 10 9 1 7 13 9 10 2 1 9 9 9 0 13 15 1 9 2 8 8 2 1 8 0 2 13 1 8 9 9 2 7 3 9 9 8 8 2 7 14 13 9 0 1 9 2 9 7 8 1 9 0 1 9 2 7 14 13 9 7 12 2 7 12 2 14 7 15 14 13 9 9 9 2 7 14 13 9 0 1 9 13 9 0 1 15 1 9 8 0 1 0 2
77 9 13 1 9 0 2 7 13 0 1 9 9 15 1 9 1 9 7 15 1 9 2 7 9 9 0 7 13 15 1 9 9 15 7 9 7 9 0 2 9 7 15 14 13 2 7 13 7 13 7 13 9 9 9 13 9 9 0 1 9 9 0 2 7 15 9 0 15 13 9 9 0 0 0 7 0 2
4 9 9 9 9
33 8 2 2 9 2 2 13 9 2 8 2 0 3 2 9 9 1 9 13 15 1 9 0 1 9 2 7 13 7 15 9 0 2
49 7 13 1 9 7 1 15 8 9 0 2 7 7 15 8 1 9 15 2 7 13 9 7 9 0 15 7 9 9 13 9 8 2 8 8 13 7 12 12 1 15 13 9 12 9 13 9 9 2
27 7 13 9 1 15 13 15 9 1 7 9 15 13 15 13 1 9 15 0 2 7 13 7 15 0 9 2
33 7 13 3 7 9 13 0 1 9 0 1 8 2 7 7 0 13 1 15 7 13 1 15 9 2 7 13 7 13 9 9 15 2
21 7 13 9 0 7 9 1 9 7 9 1 9 9 2 1 9 15 13 9 0 2
22 7 13 9 15 13 15 9 7 9 15 1 9 0 1 9 9 15 7 9 9 15 2
27 7 13 8 9 7 15 13 7 9 14 13 9 2 7 14 13 1 15 9 1 9 1 9 1 10 9 2
6 8 8 8 8 8 8
2 0 11
45 13 9 9 9 1 9 8 9 8 2 12 9 2 15 13 9 2 1 15 13 9 9 15 9 8 11 2 12 9 2 7 13 15 1 9 1 15 1 9 15 1 9 1 15 2
63 7 13 9 9 13 9 1 9 9 8 8 9 2 12 9 2 1 9 15 1 9 15 1 9 9 2 7 13 0 1 9 15 2 7 7 9 13 7 8 0 0 1 9 9 2 13 15 0 7 13 1 15 1 9 7 13 9 15 1 9 1 15 2
5 8 1 9 1 9
48 8 2 8 2 13 9 0 1 9 2 8 2 9 0 1 9 1 15 8 2 1 9 0 8 13 15 1 15 2 7 13 9 9 8 1 9 15 13 1 9 8 2 8 8 1 8 8 2
36 7 14 13 9 1 9 0 1 9 9 9 10 9 2 7 9 9 1 9 9 0 1 15 2 7 14 13 1 9 9 0 7 13 9 15 2
52 8 8 8 8 1 1 8 1 9 2 7 15 13 1 9 8 0 1 8 9 13 8 8 8 1 9 1 9 2 7 13 8 8 9 0 1 9 2 8 2 1 9 8 15 14 13 15 8 1 9 9 2
30 8 8 0 8 8 12 2 8 8 8 8 8 8 8 8 1 2 8 2 8 8 8 2 2 2 8 8 13 8 8
10 2 9 2 9 2 2 9 2 2 9
56 13 9 1 8 9 8 0 8 8 8 1 9 8 0 9 0 1 9 8 1 9 8 8 0 8 8 12 2 7 14 13 1 9 15 8 8 8 8 14 13 8 8 1 9 9 12 9 1 9 15 1 8 8 8 8 2
43 1 9 0 2 13 8 8 8 8 8 8 8 8 8 8 8 8 1 9 2 1 9 13 9 0 1 9 1 9 8 8 8 8 8 8 8 1 15 13 13 1 9 2
65 7 13 8 7 2 8 2 13 9 0 7 0 0 2 7 13 1 7 15 13 9 0 1 9 1 8 1 9 12 7 9 1 9 9 0 1 9 9 0 9 2 7 13 2 2 8 0 9 9 9 8 2 8 8 8 9 1 9 1 9 9 9 15 2 2
76 13 7 8 0 13 12 9 1 9 1 9 12 2 12 7 9 1 9 8 2 12 2 8 8 1 9 12 2 8 2 7 15 13 1 9 1 8 7 13 8 8 1 12 9 7 13 1 9 15 13 8 9 15 14 7 15 14 13 9 1 9 15 2 7 1 9 8 8 14 13 8 8 1 12 9 2
1 9
74 7 1 9 9 15 2 13 8 9 9 0 8 8 9 8 9 8 8 8 2 1 9 13 12 1 9 8 8 1 9 1 9 9 0 8 0 9 0 1 9 2 1 15 13 9 0 13 8 8 2 15 8 9 8 8 8 8 8 9 2 7 14 13 8 8 2 8 9 8 0 2 1 9 2
33 7 13 9 12 9 1 12 8 1 9 1 8 12 2 8 7 9 1 9 8 2 12 7 9 8 2 12 8 8 12 2 12 2
1 9
79 7 1 9 0 2 13 9 9 15 1 15 14 13 9 8 8 1 9 15 14 13 15 1 9 9 0 1 9 0 1 9 2 1 15 13 8 1 15 14 13 8 8 1 8 9 9 0 1 9 12 2 7 13 9 1 9 12 2 9 7 9 12 2 8 2 1 9 8 8 8 1 9 15 1 8 12 2 12 2
28 7 14 13 8 9 7 9 9 9 13 2 7 15 8 13 1 9 0 14 13 1 9 0 15 13 1 15 2
2 8 9
49 7 1 9 8 8 2 13 9 0 1 9 9 8 11 8 8 8 8 8 8 2 7 13 0 8 8 3 1 15 2 7 13 8 8 0 1 9 0 8 8 1 8 8 2 12 1 9 0 2
58 7 13 8 1 7 8 13 1 9 9 1 15 9 9 7 9 2 2 7 8 13 13 1 9 0 1 9 0 2 7 14 13 8 8 1 9 8 8 2 7 14 13 8 8 8 1 9 1 9 9 0 1 9 1 0 9 2 2
27 7 13 8 7 8 0 13 0 9 1 9 8 8 8 2 7 7 9 13 3 9 1 9 9 0 2 2
34 7 13 1 9 7 13 8 8 0 7 15 8 9 9 15 13 1 15 8 8 1 9 1 8 9 0 2 7 15 13 9 8 0 2
1 9
33 7 1 9 15 2 13 9 0 1 9 8 8 8 8 8 2 8 9 8 2 9 1 9 9 1 9 8 8 0 1 9 15 2
52 7 13 8 7 8 13 13 1 9 15 1 9 1 8 1 9 12 2 12 2 2 7 9 13 8 1 9 10 9 2 7 1 9 1 9 12 2 12 1 9 2 13 9 9 9 9 7 13 1 9 2 2
68 8 8 8 0 1 9 0 9 8 8 9 2 7 15 13 9 8 8 9 9 8 8 9 12 2 7 13 9 9 1 9 1 12 9 9 12 2 7 1 9 0 2 13 8 8 9 9 0 7 13 1 15 9 1 9 15 1 8 9 9 9 1 9 0 1 9 15 2
61 7 13 8 1 9 9 1 9 0 9 12 7 13 15 1 9 8 9 14 12 15 13 1 9 2 7 15 8 1 9 15 1 15 13 9 1 9 0 2 7 13 1 15 1 9 7 13 1 9 8 7 9 0 8 8 8 1 9 0 0 2
28 8 8 8 9 0 8 8 12 9 1 12 8 2 1 9 2 12 1 12 2 8 8 2 12 1 12 2 2
5 1 9 8 8 0
2 8 0
52 9 9 13 9 1 9 7 9 2 9 15 0 13 1 9 8 8 2 8 8 1 9 9 9 8 8 8 8 1 9 2 7 15 0 1 9 0 1 15 1 0 7 15 0 1 9 9 8 8 8 8 2
52 14 9 1 9 7 9 7 13 1 9 0 1 9 1 9 8 8 8 2 7 1 9 1 9 1 9 15 9 0 2 7 1 9 9 1 9 9 0 0 1 9 9 0 2 0 10 13 9 9 0 0 2
56 7 3 13 9 8 8 8 8 8 1 9 0 2 8 8 8 1 9 0 14 13 1 9 1 15 13 1 15 9 0 2 7 1 9 9 9 1 9 2 13 8 9 1 9 9 2 1 9 9 2 1 8 9 7 9 2
73 9 10 8 1 9 15 2 1 15 1 15 1 9 9 13 9 8 8 9 1 9 7 13 8 8 8 15 2 14 15 13 1 9 8 0 1 9 8 8 13 13 15 8 0 2 7 15 9 15 13 7 8 1 9 0 2 13 2 9 9 1 15 7 0 8 1 15 9 1 9 7 9 2
73 9 1 9 8 8 13 1 9 0 7 2 2 2 0 2 0 9 9 9 9 2 9 9 15 13 15 13 9 15 2 7 9 0 1 9 9 1 15 8 8 8 1 9 2 9 1 0 9 0 1 9 0 7 9 8 9 8 8 2 8 1 9 9 7 9 8 8 7 9 1 9 15 2
16 9 9 3 9 7 9 8 8 8 2 9 9 9 7 9 2
93 1 9 13 1 9 9 9 0 2 14 8 8 3 3 8 9 2 8 8 9 13 1 8 9 1 0 2 8 8 9 13 1 8 0 1 9 2 14 8 0 8 8 1 9 8 8 7 14 9 0 8 8 1 9 9 2 3 9 9 15 9 2 3 8 9 15 9 2 8 8 14 8 1 15 9 7 13 9 1 15 8 8 8 8 2 9 1 9 2 1 8 0 2
21 0 1 9 2 2 2 1 9 15 2 9 13 8 9 9 7 8 13 1 9 15
2 8 11
49 13 9 7 8 0 13 9 2 9 2 8 1 1 9 2 1 9 9 2 1 9 15 0 1 9 2 7 13 9 0 9 8 8 9 2 7 13 9 0 2 8 2 9 9 8 1 9 9 2
57 7 13 9 0 1 9 0 1 9 7 9 1 9 2 8 8 2 8 2 12 8 2 0 1 9 9 0 2 7 13 1 1 9 2 13 9 9 2 3 2 1 15 13 1 9 0 2 1 9 9 9 9 0 9 9 2 2
32 7 13 7 2 9 14 13 13 7 8 2 2 7 13 7 8 14 13 9 1 9 8 2 0 7 9 9 14 13 8 0 2
43 7 13 9 0 13 9 9 8 8 7 9 1 9 13 1 15 13 13 1 9 9 2 7 13 8 8 8 9 1 9 8 7 2 9 8 3 1 15 13 1 9 2 2
75 7 13 2 9 9 0 2 13 1 9 0 1 9 9 15 2 8 9 9 8 0 9 8 8 9 0 7 9 0 2 2 7 13 7 15 2 13 8 1 9 2 7 13 9 0 13 15 1 9 9 1 9 15 1 8 8 8 8 8 0 8 8 8 8 0 2 7 15 13 9 9 0 3 2 2
33 7 1 9 13 9 0 1 2 9 9 1 9 8 2 1 1 12 9 1 9 15 1 9 9 0 2 8 8 2 1 9 9 2
68 7 13 9 13 1 12 9 2 9 2 0 9 9 9 0 1 9 2 7 13 9 9 0 8 8 9 1 1 9 1 9 2 1 1 7 13 9 15 2 7 13 9 9 3 1 9 0 7 9 13 15 9 2 1 9 8 0 2 9 9 0 7 0 2 1 9 2 2
81 7 13 9 9 0 1 9 0 1 9 0 1 9 0 0 7 0 1 9 8 0 0 2 1 9 9 1 9 15 2 7 13 1 9 1 9 9 0 7 0 9 0 1 9 9 9 1 9 8 2 12 8 9 9 2 2 7 15 9 9 15 15 13 15 12 9 0 1 9 2 9 2 0 2 1 9 9 0 1 9 2
81 7 13 9 0 0 1 9 7 9 13 1 9 8 0 7 9 9 9 15 0 1 9 2 7 13 9 9 0 1 9 9 9 2 8 12 2 7 2 8 12 2 0 9 2 7 13 7 9 9 0 13 8 7 9 0 13 15 9 1 9 0 0 2 13 1 9 9 9 9 15 13 1 9 9 1 9 9 7 9 15 2
20 7 13 8 9 0 1 7 9 9 0 13 1 9 9 9 0 2 8 2 2
20 9 0 13 9 9 8 2 0 7 8 13 9 1 2 9 0 1 9 9 2
5 8 8 2 8 8
53 13 9 0 2 0 9 0 2 7 1 9 9 0 1 9 7 9 2 13 9 9 1 9 9 7 9 0 7 9 9 2 7 13 9 1 15 2 9 9 0 1 9 9 0 1 9 9 0 7 9 15 2 2
66 13 1 9 3 9 9 1 0 7 8 1 9 1 9 9 7 9 9 7 9 9 9 1 9 15 0 2 7 15 1 9 9 9 1 9 2 1 7 13 1 9 9 8 8 9 2 1 9 14 13 15 9 9 0 8 8 1 9 15 0 8 8 1 9 0 2
105 7 13 1 9 0 13 1 9 7 9 0 0 8 8 7 0 8 8 8 13 9 9 9 1 9 0 2 7 13 7 9 0 13 1 9 1 9 9 9 0 7 9 7 9 2 7 9 9 9 0 7 0 0 7 9 9 1 9 7 9 15 7 9 15 2 7 13 1 2 9 9 9 9 0 1 9 9 0 0 1 9 9 0 7 9 15 2 9 1 9 9 9 0 15 13 15 9 9 9 1 9 9 12 2 2
48 7 13 9 0 0 7 9 0 13 1 2 9 1 9 9 1 9 9 0 2 9 1 9 9 1 9 9 1 15 1 9 9 1 9 15 0 2 7 9 9 9 0 1 9 1 9 2 2
29 7 13 9 1 9 2 9 9 2 2 13 9 15 13 9 1 15 2 1 10 1 10 9 9 7 9 7 9 2
55 7 13 9 0 0 1 9 8 15 13 15 9 7 9 9 12 2 7 13 9 0 0 7 9 0 1 9 14 13 2 9 9 9 3 1 12 9 2 7 13 9 1 9 9 1 9 9 1 9 1 15 1 1 9 2
72 7 13 1 8 7 9 0 0 14 13 9 1 9 1 9 15 9 9 14 13 1 0 2 7 2 9 9 9 0 2 2 7 13 9 1 9 2 9 9 2 9 1 9 9 2 7 13 7 10 9 13 9 1 9 15 2 7 14 13 9 0 13 1 9 9 9 9 9 1 9 9 2
25 13 9 1 9 0 8 1 9 8 2 9 8 8 2 2 8 2 14 8 9 7 8 13 9 9
7 8 2 8 2 9 0 2
79 13 9 9 0 11 8 8 3 7 9 15 14 13 1 9 15 9 9 9 2 1 0 9 2 2 0 9 9 15 1 9 0 9 0 1 9 2 7 0 8 1 7 15 2 13 9 1 9 9 2 2 7 13 9 0 9 1 9 0 2 0 9 1 9 9 0 8 8 8 1 7 15 9 2 9 8 8 2 2
132 13 9 9 0 11 8 8 3 7 9 14 13 2 1 0 9 2 1 9 15 9 9 9 0 2 7 13 9 9 0 15 13 15 8 0 1 7 15 2 9 2 2 7 13 1 9 0 13 15 9 2 9 2 0 3 2 2 8 8 8 8 2 9 9 2 7 14 13 3 9 1 0 9 1 0 9 1 9 15 8 9 1 8 8 8 8 8 2 2 7 13 7 9 9 2 9 9 1 9 9 8 8 8 8 9 1 9 0 2 2 7 13 7 15 8 9 0 15 2 9 9 8 8 1 8 9 8 8 8 8 2 2
24 7 13 8 2 2 13 7 13 9 9 1 9 9 2 9 1 9 2 0 1 9 9 2 2
94 7 9 1 9 1 9 9 15 13 1 15 10 9 2 13 9 9 0 2 2 14 8 8 8 8 2 2 2 2 2 14 15 9 7 14 13 7 8 1 15 9 1 8 8 2 0 3 7 15 9 13 8 8 8 8 8 2 7 1 8 8 7 8 9 0 9 8 7 15 13 8 8 8 2 8 2 9 2 13 8 1 8 8 7 13 1 0 15 7 13 9 15 2 2
95 7 13 7 13 9 0 2 0 1 9 9 0 1 9 1 9 9 9 0 7 9 9 0 2 7 13 7 2 9 9 0 13 9 8 8 1 9 9 9 9 15 8 1 15 8 8 1 9 2 2 7 13 0 7 9 2 14 13 1 0 9 13 7 13 1 9 9 14 13 1 9 9 1 9 0 2 2 7 13 1 7 15 2 1 1 15 14 13 7 8 1 0 9 2 2
62 7 13 13 0 1 3 1 9 15 2 9 9 0 0 2 1 9 7 9 15 8 1 9 0 9 0 1 9 2 7 13 7 2 9 0 9 0 8 8 0 14 13 14 0 1 15 13 1 15 9 9 0 2 15 13 1 9 2 9 0 2 2
86 1 15 2 13 8 8 1 7 15 2 14 13 13 9 1 9 9 2 0 1 9 15 2 1 9 9 2 2 7 13 7 9 9 1 9 7 9 2 9 8 2 2 0 7 9 2 14 13 13 9 9 0 1 9 15 9 1 9 2 7 13 9 0 1 9 9 9 0 1 8 7 9 0 2 7 13 9 9 0 7 0 1 9 15 2 2
151 7 13 9 8 0 9 1 9 0 2 15 13 15 9 0 2 2 7 13 2 2 14 8 7 14 8 9 1 9 9 7 9 10 13 1 9 15 7 13 1 9 8 7 8 7 9 2 8 8 9 0 2 2 7 13 9 1 9 9 15 1 7 15 2 9 0 13 9 1 9 0 1 9 2 8 8 9 9 9 1 9 15 1 9 10 9 2 7 7 8 9 1 9 8 9 8 8 8 1 8 0 8 8 2 2 7 13 1 9 15 13 1 9 0 1 9 0 1 9 2 0 14 15 9 8 8 2 2 0 7 9 14 13 1 9 9 15 2 13 1 9 8 1 1 9 15 13 15 0 2 2
7 9 2 8 9 13 8 0
2 8 8
86 13 3 8 8 1 8 9 9 2 9 2 0 1 9 9 0 8 8 0 1 9 9 8 8 2 15 13 9 7 9 14 13 15 15 8 1 9 15 2 7 13 8 8 9 8 8 7 15 14 13 9 9 1 9 1 9 9 7 14 13 9 9 8 1 9 15 8 0 2 1 7 13 9 8 8 13 15 1 0 1 9 8 8 1 15 2
90 7 1 9 1 15 7 13 9 0 0 1 9 9 1 9 9 8 15 14 13 0 1 9 8 8 2 7 13 7 9 2 15 14 13 8 2 8 1 9 0 8 8 1 9 2 7 13 9 9 0 7 0 1 9 15 2 1 1 7 9 0 8 13 9 9 8 8 8 0 7 9 1 9 15 9 2 7 14 13 9 9 15 14 13 9 1 15 10 9 2
72 7 13 7 13 9 9 0 9 1 8 2 9 9 2 2 7 13 9 9 2 1 9 15 1 9 2 7 13 9 9 9 8 8 9 0 1 9 1 9 2 8 0 2 2 9 1 9 8 8 8 8 8 2 7 3 13 9 9 9 8 8 7 9 9 8 8 1 9 1 9 9 2
49 7 13 9 9 1 9 3 7 15 14 13 9 9 0 1 10 9 1 9 9 0 9 0 2 13 9 0 0 2 1 8 9 9 9 0 1 9 0 2 8 8 1 9 2 7 13 8 9 2
26 7 13 0 0 1 9 0 9 1 9 3 2 8 8 1 9 8 8 2 7 9 0 1 10 9 2
10 9 13 1 9 9 8 8 1 9 15
1 8
33 13 9 0 3 7 9 13 9 13 15 12 8 1 9 1 15 1 9 9 8 2 1 8 9 0 2 1 9 9 1 9 9 2
63 7 13 8 8 8 2 9 9 9 1 8 2 1 9 2 8 8 2 7 9 15 13 8 13 1 8 8 2 14 13 3 8 8 2 2 7 13 9 0 9 9 1 9 9 9 12 9 1 9 9 9 8 0 2 7 14 8 8 9 1 9 9 2
86 7 13 9 13 1 9 9 1 9 2 9 2 2 1 1 9 0 2 7 13 7 9 9 15 13 13 1 9 1 9 7 9 2 7 13 9 15 1 9 9 0 2 7 13 9 0 9 8 1 9 2 7 13 8 7 9 13 1 9 9 15 9 1 9 15 2 7 10 9 13 1 1 9 0 1 9 9 1 9 9 8 1 9 7 9 2
9 9 8 8 8 8 13 8 8 8
53 13 2 9 2 1 8 3 9 1 9 8 8 13 15 1 9 8 8 8 1 8 7 8 7 8 8 8 7 8 7 8 7 8 7 9 2 13 1 15 9 8 8 8 8 11 8 8 8 8 2 8 2 2
18 7 13 7 8 2 8 8 1 9 7 9 0 1 1 10 9 2 2
60 7 13 9 8 1 8 1 9 2 9 2 0 1 9 2 8 8 8 1 9 2 13 7 15 2 13 8 9 8 11 8 8 8 8 0 1 9 2 9 1 9 2 2 7 13 9 10 9 1 9 1 2 8 9 9 1 9 9 2 2
11 9 2 9 7 12 9 1 9 1 9 9
30 9 2 8 2 2 9 2 2 8 2 13 9 0 7 9 1 9 9 1 9 1 9 0 9 13 9 7 12 9 2
48 7 13 1 9 9 0 1 8 8 1 9 1 9 1 9 8 2 9 2 2 0 7 9 13 9 0 2 1 9 8 9 1 9 9 1 9 0 2 7 13 9 9 1 9 1 10 9 2
40 7 1 8 13 2 9 2 9 1 9 2 9 8 2 0 0 2 13 1 9 9 0 1 9 3 9 9 9 2 8 2 1 9 2 8 0 2 9 8 2
9 8 8 2 8 13 9 1 9 0
79 13 9 0 8 8 8 0 1 9 0 1 9 0 8 8 8 2 7 9 13 7 9 9 0 13 1 9 13 9 0 13 1 9 8 9 0 1 9 9 9 0 7 0 2 1 9 15 13 15 9 8 2 7 9 9 0 9 9 2 2 7 13 8 13 8 1 9 0 1 9 9 9 0 1 9 8 8 8 2
42 7 13 8 1 9 2 9 8 9 15 13 9 0 1 9 2 9 9 0 8 15 13 9 1 9 9 1 9 0 13 9 15 1 9 1 9 7 0 7 9 2 2
63 7 13 8 7 15 13 9 8 1 9 8 8 2 1 9 9 9 0 1 9 0 1 9 0 1 9 2 7 9 1 9 15 14 13 1 8 1 9 9 9 0 1 9 0 2 7 13 1 7 15 14 13 9 1 9 1 9 9 0 1 9 0 2
36 7 13 8 9 9 0 8 8 15 13 1 15 2 8 1 9 8 9 9 0 7 9 9 9 15 7 10 9 0 1 9 0 1 9 2 2
20 7 13 8 1 15 9 9 8 8 1 9 9 9 9 1 9 0 8 8 2
57 7 13 9 9 13 9 0 1 9 8 8 15 13 15 9 9 8 8 2 0 1 9 0 1 8 2 7 7 8 14 13 15 1 9 15 8 8 10 9 2 1 1 9 0 13 1 9 15 13 15 9 0 1 10 9 2 2
40 7 13 9 9 9 8 8 1 9 9 0 7 13 1 9 8 2 0 2 7 9 9 15 15 9 8 8 1 9 2 2 9 1 2 9 1 8 9 2 2
14 9 1 9 7 0 1 9 9 9 0 1 12 12 9
2 8 8
56 13 9 0 7 0 2 7 9 0 1 9 1 15 7 9 0 1 9 9 14 13 2 2 7 13 1 2 9 9 9 0 1 15 1 12 12 9 0 7 9 9 0 1 9 1 9 9 9 1 9 1 9 9 7 9 2
25 13 15 1 9 9 2 9 0 2 0 0 2 1 9 9 9 0 8 8 8 7 0 8 8 2
75 7 13 9 0 2 7 9 13 1 9 9 0 1 9 8 8 9 9 0 8 8 9 9 9 8 8 9 9 1 9 8 8 0 9 0 13 9 9 0 7 9 0 7 0 7 0 7 9 8 7 9 9 1 9 9 7 9 7 9 7 9 7 9 7 9 8 8 7 9 0 2 0 0 2 2
115 8 8 9 2 9 0 1 9 8 9 7 9 8 8 0 8 8 9 9 7 9 9 7 9 9 0 2 2 7 13 8 2 7 9 0 13 1 9 9 13 7 13 9 1 9 9 2 2 7 13 2 2 13 9 1 9 9 1 9 0 7 15 13 13 9 1 9 0 1 0 2 2 7 13 8 2 7 10 9 13 9 9 8 8 0 1 8 9 9 8 0 8 8 9 0 2 0 2 2 7 13 8 8 1 7 8 14 13 8 8 8 8 9 15 2
6 9 9 9 13 9 9
41 13 9 9 9 9 0 0 9 8 11 8 8 8 1 9 8 3 9 9 0 8 9 1 9 9 9 8 8 0 9 11 11 8 7 9 8 1 9 8 8 2
40 7 1 9 1 9 7 9 13 9 0 1 9 7 9 15 13 15 9 9 1 9 1 9 9 9 7 9 1 9 0 0 0 1 9 1 9 2 9 2 2
9 2 8 2 13 7 13 9 8 8
35 8 2 8 2 8 8 8 2 13 9 1 9 9 2 8 2 0 1 8 7 15 14 13 7 13 8 11 8 0 1 9 1 9 0 2
96 7 13 11 8 1 9 2 8 2 1 9 8 1 9 8 2 2 15 13 1 9 0 13 9 13 1 15 8 0 2 14 13 1 9 9 2 2 8 11 8 14 13 15 9 15 2 2 7 14 8 2 2 2 8 14 8 9 2 2 8 8 14 13 9 2 2 8 8 8 8 2 2 14 13 8 1 9 8 0 1 9 0 7 9 15 0 2 2 8 14 13 15 9 15 2 2
39 7 1 8 8 13 9 9 2 8 2 9 2 7 13 2 9 9 0 2 8 0 1 9 8 1 8 8 2 14 15 9 0 8 8 8 8 8 2 2
21 7 13 8 7 15 13 9 1 9 0 1 10 9 7 13 8 9 1 9 15 2
16 8 13 9 1 2 9 0 2 8 7 13 8 8 0 12 9
67 9 0 2 8 2 8 2 2 9 2 2 8 2 8 8 8 2 13 8 0 7 0 8 8 8 1 9 1 9 0 2 7 13 0 9 1 15 1 9 9 0 1 9 9 8 7 8 2 7 13 9 1 9 9 0 1 9 1 9 1 10 9 8 8 8 9 2
25 7 13 9 9 0 1 9 7 8 13 8 3 8 8 0 1 9 12 9 1 9 9 9 0 2
98 7 13 9 9 0 8 8 8 3 9 0 8 8 9 7 9 9 0 1 9 9 2 7 13 9 9 0 8 11 8 1 8 1 9 15 13 15 2 8 8 0 2 2 7 13 7 2 9 13 9 15 8 1 15 0 1 7 9 0 15 9 0 1 9 0 2 2 7 13 9 9 8 8 7 15 13 2 8 1 9 9 15 2 2 7 13 2 9 9 0 1 9 1 9 9 9 2 2
34 7 13 9 1 9 9 9 0 7 9 0 0 1 9 9 1 8 1 9 15 13 15 9 0 2 8 1 9 15 8 1 9 2 2
63 7 13 8 8 2 2 8 1 9 8 1 9 7 7 13 7 15 13 1 9 0 15 9 0 7 7 8 13 9 8 8 7 13 1 9 15 1 9 10 9 2 2 7 13 9 9 7 9 0 8 8 7 13 1 1 8 8 9 15 13 9 0 2
57 7 13 8 8 0 1 9 1 9 0 9 9 15 1 9 2 7 13 9 0 0 2 7 13 9 1 9 9 9 0 1 9 8 8 8 9 2 7 13 9 0 7 15 14 13 1 8 8 8 1 9 15 13 9 15 0 2
53 7 1 8 2 13 9 7 9 0 1 8 8 1 9 1 9 9 13 8 8 1 7 15 9 0 2 7 13 8 1 9 9 9 7 9 13 9 9 1 9 9 9 1 9 0 8 8 8 1 9 1 8 2
5 8 8 1 9 9
32 1 9 13 15 9 0 2 13 9 9 0 8 8 7 9 9 0 13 1 9 12 0 1 9 12 9 0 13 1 9 0 2
26 7 2 9 9 0 2 2 8 8 8 2 7 9 0 0 9 9 14 13 15 9 0 1 9 15 2
5 2 8 8 8 2
87 7 13 2 9 9 0 2 1 9 9 9 0 0 8 8 9 9 8 8 1 9 9 0 1 9 0 7 12 2 7 13 9 1 8 8 13 15 8 1 8 0 7 1 9 13 1 9 9 2 8 8 9 7 10 9 13 9 8 9 0 7 14 3 9 8 8 1 15 1 9 0 8 8 2 7 13 1 9 9 8 1 9 0 1 9 0 2
6 8 2 8 2 8 2
41 13 2 9 9 0 2 2 8 8 8 2 9 12 1 9 9 8 8 2 7 13 1 9 9 9 9 1 0 8 0 8 8 9 7 9 9 0 1 9 0 2
13 7 1 9 9 9 9 1 9 0 7 1 15 2
3 9 9 0
52 13 2 9 9 0 2 2 8 8 8 2 9 0 8 0 15 8 1 9 8 2 7 15 9 0 9 7 13 1 9 9 9 1 9 0 2 7 9 9 1 9 8 1 9 0 1 9 13 8 8 0 2
21 9 9 0 2 14 8 0 9 14 13 8 8 1 9 8 8 2 9 8 13 8
6 8 8 2 8 8 8
44 13 9 9 0 9 8 11 11 9 0 8 8 8 15 13 9 1 9 9 0 9 1 9 0 1 9 0 1 9 9 9 0 7 9 0 7 9 0 7 0 9 9 0 2
34 7 13 9 8 9 1 9 0 1 9 9 9 9 11 11 11 7 9 0 1 9 9 9 9 9 7 9 9 0 9 8 11 11 2
19 7 13 8 0 7 9 15 13 0 7 13 9 13 8 8 1 9 9 2
60 7 1 9 13 9 0 1 9 0 8 8 9 11 9 8 8 9 15 0 9 1 9 9 9 1 8 7 9 9 0 1 9 1 9 8 2 8 2 7 9 0 0 7 13 15 1 2 9 9 9 0 2 7 15 9 9 8 8 9 2
51 7 13 11 1 9 0 9 1 9 9 0 0 1 9 7 9 1 9 13 9 0 1 9 9 0 2 7 13 7 9 2 14 13 9 15 8 8 9 9 15 7 14 13 1 9 15 8 8 8 2 2
88 7 13 9 0 1 9 1 9 0 8 8 1 3 1 9 8 1 9 9 7 9 15 2 14 13 0 9 8 8 9 9 1 8 7 2 8 2 7 9 0 14 13 9 9 0 0 1 9 9 0 7 7 13 1 15 8 8 8 8 8 8 8 8 8 8 8 9 8 8 8 8 2 2 7 13 2 2 8 8 14 8 8 1 9 7 9 2 2
58 7 13 2 2 8 8 14 13 1 9 7 6 1 9 7 9 7 9 7 9 0 7 0 1 9 9 7 9 9 2 8 8 13 1 9 8 8 7 14 13 8 8 9 7 8 1 9 7 9 8 1 9 8 8 8 8 2 2
45 7 13 1 9 1 9 9 0 15 13 15 9 8 8 7 13 9 9 1 9 7 2 9 0 1 9 9 2 8 1 9 8 8 9 1 7 15 13 8 9 1 9 7 9 2
59 7 14 13 9 0 1 9 1 9 13 15 1 9 15 1 9 9 9 15 9 0 1 9 0 9 0 2 9 7 15 13 1 7 9 9 15 15 13 15 2 7 13 9 15 1 9 1 9 0 2 0 0 7 15 14 13 1 15 2
10 9 0 0 1 9 9 9 2 9 2
43 13 9 0 0 1 9 9 0 1 9 9 0 0 1 9 1 9 0 2 9 2 0 1 9 1 9 9 9 0 0 1 9 0 1 9 0 0 1 2 9 9 2 2
43 7 13 9 9 9 0 7 0 7 9 9 0 9 0 1 9 1 9 1 12 9 0 8 8 8 8 2 7 13 9 1 9 7 9 0 13 1 9 9 0 1 9 2
59 7 13 9 9 9 0 9 8 8 1 2 9 2 7 2 9 0 9 0 13 0 1 15 7 13 9 15 15 13 1 9 8 8 0 1 9 8 8 8 8 0 1 9 0 0 2 9 7 9 0 0 1 9 8 0 13 0 2 2
66 7 13 9 9 0 0 1 9 1 7 2 9 9 9 0 1 8 8 9 0 8 7 9 8 0 7 9 0 0 1 8 9 9 14 13 1 9 7 9 9 9 1 10 9 2 7 1 10 9 13 9 1 9 9 15 0 1 9 0 7 0 1 0 9 2 2
86 7 1 1 7 8 1 2 9 9 0 2 13 7 2 9 9 0 8 8 2 2 7 15 14 13 7 2 13 8 8 1 9 0 0 1 9 9 0 8 8 9 9 0 2 2 7 13 1 7 2 9 1 9 14 13 1 9 9 9 13 9 9 9 0 0 2 7 13 9 9 0 1 9 8 8 9 9 0 7 9 9 9 1 9 2 2
62 7 13 8 7 9 15 13 9 1 9 9 0 1 9 8 7 8 8 13 1 9 2 9 0 8 8 1 9 9 9 9 0 1 9 1 9 7 15 15 13 9 10 9 7 9 15 1 9 9 9 7 9 8 8 1 9 8 8 8 8 2 2
64 7 14 13 9 15 14 13 1 9 2 9 9 0 8 8 9 9 2 1 12 9 0 0 15 2 9 9 9 0 2 7 9 1 9 7 8 1 9 7 9 0 2 2 2 7 0 2 9 0 1 9 9 9 2 7 0 2 9 0 7 9 9 2 2
12 9 0 2 9 2 8 2 14 13 13 1 8
1 8
61 13 9 2 8 8 2 0 3 1 7 9 15 13 1 9 9 2 8 2 0 1 9 2 8 2 1 9 0 2 9 2 12 1 9 8 0 14 13 13 1 8 2 0 1 15 9 1 9 9 0 15 13 1 9 9 1 9 9 8 8 2
43 7 13 9 7 9 1 9 8 1 8 8 8 8 13 1 8 1 9 7 9 1 8 9 0 8 8 9 9 0 14 13 1 9 1 12 9 1 8 8 12 1 8 2
48 7 13 9 7 15 13 7 13 9 13 1 10 9 1 9 15 13 8 1 15 7 13 1 9 9 15 1 8 9 2 7 13 9 1 9 15 8 8 1 8 2 7 13 1 9 12 9 2
37 7 1 12 9 0 2 9 2 0 13 9 0 13 1 8 8 2 8 2 1 9 2 12 9 2 1 9 0 7 13 0 0 0 8 8 8 2
87 7 1 1 8 9 0 2 13 9 9 1 9 7 9 15 13 9 13 1 9 9 1 8 2 8 2 2 7 13 7 8 13 1 9 0 1 8 7 13 15 8 8 8 1 15 1 9 0 8 1 1 9 15 1 9 0 9 2 7 13 8 1 9 0 9 1 15 1 10 9 2 7 13 1 15 9 0 9 0 1 9 9 0 1 9 15 2
47 7 13 9 0 13 8 8 1 9 8 13 1 9 9 15 14 13 15 9 8 2 7 15 13 15 9 0 1 9 1 9 9 0 1 12 9 0 2 9 2 0 1 8 8 1 8 2
47 7 13 8 7 15 13 1 9 8 1 9 1 9 0 1 9 15 7 7 9 13 15 1 9 2 7 13 9 7 8 8 13 8 8 0 13 2 7 0 14 8 1 9 15 1 9 2
10 9 2 9 9 13 1 9 9 9 0
2 9 8
74 13 9 9 9 1 9 3 9 1 9 9 9 0 9 8 9 9 7 12 1 0 9 7 9 9 1 15 12 13 9 9 0 1 12 1 9 0 2 1 9 9 9 9 9 0 1 9 13 1 9 2 7 13 9 0 7 9 9 1 9 13 1 9 9 8 8 0 8 8 8 8 1 15 2
79 7 13 9 0 9 8 11 13 9 7 9 9 9 0 8 11 7 12 1 9 1 9 8 8 9 9 1 9 2 9 2 0 1 9 1 15 13 1 0 2 9 1 8 8 8 1 9 9 15 8 8 8 8 1 9 9 8 8 8 9 2 2 7 13 9 1 0 0 2 8 1 9 9 9 8 8 8 2 2
90 7 13 9 1 12 9 1 15 12 9 0 1 9 7 9 9 9 7 9 9 9 9 8 9 11 2 7 1 9 9 9 13 9 9 9 9 0 7 12 0 1 9 0 1 9 8 1 9 8 0 2 7 13 12 8 9 8 1 9 7 13 12 9 7 15 14 13 0 9 7 14 13 1 15 0 9 2 7 13 0 8 1 9 0 9 8 1 12 8 2
15 9 2 9 1 9 12 9 9 1 12 12 9 1 9 0
2 8 8
174 13 9 0 1 9 9 0 0 1 9 0 0 12 9 9 1 9 15 1 9 15 0 12 15 13 15 9 0 2 7 13 9 0 1 9 0 7 9 13 9 0 1 9 1 9 12 0 0 1 9 0 1 7 13 9 9 0 0 1 12 12 9 7 12 12 2 12 1 12 12 9 2 2 7 13 9 9 15 14 13 1 9 1 1 12 9 0 2 1 9 1 7 13 9 9 0 1 0 1 12 12 9 2 7 13 1 9 9 9 9 0 1 0 1 12 12 9 7 14 9 14 13 9 1 9 0 0 9 0 1 9 9 2 9 0 2 15 13 9 1 9 1 9 9 0 1 9 15 1 9 9 12 9 9 15 13 0 1 0 0 0 1 9 0 2 7 15 9 0 15 14 13 9 2
137 7 13 9 7 9 8 1 9 0 1 9 0 13 1 9 9 0 7 9 9 0 13 9 0 2 13 1 15 7 9 13 1 9 0 13 9 0 1 9 1 15 8 8 8 9 0 8 0 1 9 0 0 13 1 12 7 9 12 9 0 15 13 9 15 1 9 1 9 9 15 9 0 1 9 1 9 0 0 15 8 1 15 9 0 2 7 13 9 0 7 9 9 1 9 15 0 1 9 9 0 9 9 1 8 1 9 8 8 8 1 8 9 9 14 13 1 9 9 0 1 9 1 9 9 0 7 1 9 8 9 1 9 8 14 1 12 2
19 13 8 8 9 15 12 12 9 2 13 8 9 0 1 9 9 8 8 0
104 13 9 9 0 1 9 9 0 7 15 13 1 8 9 1 9 8 8 13 15 9 2 8 8 2 7 2 8 2 0 1 9 0 0 1 9 9 8 8 2 7 13 9 8 8 2 9 0 1 15 1 9 12 7 12 12 9 15 8 9 0 0 1 9 7 9 9 1 0 9 1 10 9 1 9 9 9 9 9 2 2 7 13 9 0 13 1 9 12 12 9 0 8 1 9 9 9 0 7 9 9 8 8 2
84 7 9 9 7 9 13 9 1 9 2 9 2 12 1 9 1 9 0 7 9 0 8 8 8 9 1 9 7 9 7 9 8 0 0 1 9 9 1 9 8 8 8 2 8 2 8 2 1 9 2 8 8 8 2 2 2 7 13 9 1 9 1 9 9 13 9 0 1 9 9 8 8 9 2 15 13 9 1 9 9 1 9 0 2
132 7 13 9 9 8 8 1 9 9 11 0 8 8 8 0 8 8 8 8 2 7 13 9 0 1 9 7 9 9 2 13 1 15 9 9 1 9 0 7 9 9 0 15 8 1 9 0 2 7 1 9 9 13 9 1 0 15 8 8 8 8 12 9 1 9 0 7 12 8 1 9 0 2 7 13 9 9 8 8 8 7 13 9 1 9 1 9 0 13 15 8 9 8 1 9 0 8 8 8 8 8 1 9 0 2 7 13 9 1 9 13 12 9 13 1 15 9 0 7 9 0 9 2 7 13 9 0 12 7 9 15 2
71 7 13 9 0 8 8 1 9 1 9 9 9 0 1 9 2 0 1 9 9 0 1 9 8 8 12 12 9 1 12 12 2 8 8 13 9 0 9 9 9 1 9 7 9 0 7 13 1 8 9 8 13 7 9 0 13 1 15 9 9 7 9 7 13 9 9 1 9 15 0 2
76 7 13 9 0 8 8 9 0 2 0 7 9 9 9 2 9 0 9 7 7 9 8 1 15 13 1 9 7 13 1 15 1 9 1 9 8 2 2 7 13 9 8 8 9 2 7 13 9 0 1 9 0 8 9 9 1 9 8 8 8 8 8 8 0 8 8 8 8 8 0 8 1 8 8 8 2
9 2 8 8 2 13 9 0 1 8
51 8 2 2 9 2 2 13 2 9 0 0 1 9 2 2 8 8 2 9 9 9 8 1 9 15 8 8 9 15 2 0 8 8 8 8 1 8 2 8 8 1 9 8 0 2 1 9 12 12 0 2
46 7 13 9 13 15 9 2 1 9 9 9 9 0 9 15 2 2 14 13 9 12 9 8 8 0 0 8 8 0 1 12 8 9 0 1 9 0 13 1 1 12 12 0 2 2 8
49 7 13 1 7 9 0 1 9 7 9 0 13 1 9 12 12 0 2 7 13 9 1 9 2 8 8 2 1 9 10 9 15 12 12 0 1 9 7 1 7 9 9 15 7 8 8 1 9 2
9 9 9 0 2 0 1 9 7 9
117 9 2 2 9 2 2 13 9 7 9 0 1 3 8 1 9 1 9 9 7 9 13 9 9 7 9 0 7 0 2 7 13 9 1 9 9 0 1 9 1 9 9 7 9 9 9 13 9 9 9 13 1 9 9 0 9 15 1 9 2 7 13 9 15 13 15 1 9 0 9 9 9 8 11 9 8 8 7 1 9 0 9 9 7 9 9 11 11 9 8 9 9 7 9 7 9 7 9 9 9 0 1 9 1 9 9 8 7 9 9 1 9 0 0 1 9 2
13 9 1 2 9 1 9 2 1 9 1 9 8 8
73 9 2 2 9 2 2 13 9 9 0 1 9 15 15 13 15 0 1 3 1 9 9 9 0 9 8 11 11 1 9 2 9 9 1 9 0 2 9 9 1 9 8 8 8 8 8 1 9 9 0 8 8 8 9 0 1 8 8 8 8 12 9 0 1 9 8 9 9 8 8 9 9 2
9 9 13 8 8 1 9 12 12 9
35 8 2 8 2 13 2 9 8 9 2 3 7 9 13 9 0 8 8 8 12 9 1 9 12 12 9 1 9 8 9 7 9 0 0 2
57 7 13 8 1 9 9 7 15 9 0 1 9 7 8 8 2 9 9 2 13 0 1 3 8 8 0 13 12 1 12 0 9 1 12 1 12 1 8 9 0 2 7 13 7 9 0 1 9 7 13 9 9 9 12 12 9 2
62 8 8 0 1 9 0 7 9 0 0 1 9 1 14 13 9 0 1 9 1 12 12 9 2 7 13 8 1 9 12 9 2 9 2 7 13 1 12 9 0 2 9 2 0 2 8 8 1 8 8 13 8 8 1 9 1 9 8 9 0 9 2
68 7 1 9 0 1 9 0 13 9 9 0 1 9 12 12 9 13 15 9 0 7 1 1 0 9 2 7 13 9 1 10 9 0 12 1 12 13 9 12 9 1 9 2 9 2 7 9 2 7 13 1 9 12 9 0 0 7 12 9 0 7 12 9 0 1 9 0 2
12 9 9 0 13 9 9 15 12 12 9 1 8
1 8
28 13 9 9 0 1 9 7 15 13 0 1 3 9 9 1 9 12 12 9 1 9 9 9 0 1 9 0 2
46 7 13 9 7 10 9 13 1 9 9 8 9 15 12 9 7 9 15 0 12 12 9 2 7 13 9 1 7 2 10 9 0 1 9 9 9 0 0 1 9 9 7 9 9 2 2
26 7 13 9 9 0 7 8 14 13 2 0 1 9 9 9 7 9 2 1 9 13 1 9 9 15 0
17 9 1 9 9 9 9 7 9 2 9 13 9 1 9 12 12 9
2 8 8
50 13 9 0 9 1 9 0 0 15 13 9 9 1 9 9 9 2 1 9 12 12 9 2 1 9 0 1 9 9 7 9 0 7 9 9 2 7 13 9 1 9 9 9 9 9 7 9 1 9 2
24 13 9 0 1 9 9 9 9 9 7 9 1 9 1 9 9 0 15 13 1 9 9 0 2
40 7 13 0 9 1 9 9 10 9 1 9 1 9 9 9 0 7 9 13 1 15 1 9 9 0 7 9 9 1 9 15 0 0 1 9 9 15 0 0 2
36 13 1 7 9 13 1 9 0 12 9 1 9 9 10 9 1 9 9 9 9 7 1 7 13 9 9 1 9 9 0 1 0 7 13 9 2
65 1 9 9 15 13 2 9 2 7 9 9 7 9 13 9 9 1 9 0 9 1 9 9 0 1 9 9 7 9 0 7 9 9 2 7 13 9 10 9 1 12 12 9 2 7 13 9 9 1 8 7 9 2 8 8 8 2 13 9 1 9 9 10 9 2
33 7 13 9 7 13 9 9 0 9 9 1 9 0 1 9 9 9 1 7 9 14 13 9 15 13 1 9 9 0 13 9 12 2
48 7 13 9 1 9 9 0 9 1 9 9 7 9 1 9 1 9 9 9 0 9 7 9 13 1 9 9 0 15 13 7 9 9 1 9 0 1 9 9 9 9 14 13 1 9 9 15 2
42 7 13 9 9 0 2 7 1 13 9 9 14 13 9 14 12 9 1 9 12 13 1 15 2 7 13 9 15 14 13 9 1 9 12 1 9 9 0 9 9 9 2
17 9 1 9 9 1 9 9 2 9 2 12 12 9 9 1 9 12
2 8 8
51 13 7 13 9 9 0 1 9 9 0 1 8 7 8 7 9 0 0 1 12 12 9 9 9 2 7 12 12 9 9 9 0 2 1 9 15 13 9 13 9 9 1 9 9 1 9 0 7 13 9 2
59 13 9 0 9 1 9 14 13 1 9 9 0 1 9 9 9 0 0 14 13 9 15 1 12 12 9 9 9 0 7 1 12 12 9 2 1 0 9 2 1 9 9 0 7 15 9 15 13 15 9 0 1 9 15 1 9 9 0 2
44 7 13 9 2 1 9 13 9 1 12 9 2 9 2 0 7 1 9 2 7 9 1 9 0 7 14 13 1 9 7 14 13 9 9 0 1 9 1 9 9 1 9 0 2
33 7 13 9 9 9 1 9 1 2 9 2 15 13 15 9 9 8 8 8 1 3 1 9 9 0 1 9 1 9 7 9 3 2
55 7 13 9 2 7 9 0 13 9 7 9 1 9 2 0 1 7 9 9 15 0 15 13 7 14 13 1 9 0 15 13 9 9 9 1 9 7 9 9 9 15 1 9 7 9 9 15 1 9 9 1 0 1 9 2
34 7 13 9 1 9 0 7 10 9 15 0 8 2 1 9 1 9 15 9 0 3 12 12 9 1 9 9 1 9 0 13 9 15 2
101 7 13 9 9 9 1 9 9 0 8 8 1 2 9 2 7 15 13 15 9 13 1 9 9 2 7 9 9 13 7 9 9 14 13 9 9 1 1 12 12 9 1 0 2 12 8 1 12 12 9 2 1 9 9 0 2 7 14 13 9 9 0 12 1 12 1 0 7 15 0 12 12 9 2 7 13 7 9 7 9 13 0 13 9 9 1 9 9 1 9 9 1 9 9 7 9 9 9 9 0 2
35 7 13 7 13 9 1 9 9 0 0 1 9 9 9 7 9 0 7 0 9 7 9 10 9 13 1 12 12 9 2 12 12 9 2 2
64 7 13 9 0 9 9 1 9 9 10 13 0 7 13 1 9 0 1 9 15 9 9 9 9 1 9 0 7 9 9 9 9 15 13 1 15 9 7 13 9 9 9 1 15 1 9 2 1 9 1 9 9 1 9 0 1 9 9 15 1 9 9 0 2
68 7 13 9 9 1 9 9 0 1 3 7 9 13 9 0 1 9 9 1 9 1 9 7 9 9 1 9 15 1 9 1 9 0 1 1 15 9 9 7 9 8 2 7 13 9 1 15 9 9 0 7 0 2 9 9 2 1 9 0 7 9 9 0 1 9 1 9 2
33 7 13 7 14 13 3 9 1 9 9 1 9 15 13 9 9 9 1 9 12 1 12 14 13 1 12 1 12 1 9 9 9 2
26 8 13 1 9 15 0 1 8 1 9 9 15 2 8 13 1 9 9 9 7 13 9 15 1 9 0
2 8 8
71 13 9 9 0 8 8 1 9 9 9 1 8 1 9 13 9 9 2 0 2 1 9 9 0 2 7 13 8 1 9 13 1 15 1 9 2 8 2 9 1 9 1 9 9 0 8 8 8 1 7 8 14 13 1 9 9 0 7 0 1 10 13 9 0 7 7 13 9 15 0 2
42 7 15 9 0 15 13 9 9 1 9 1 9 9 9 1 8 2 7 13 13 1 9 1 9 1 15 1 9 9 15 9 1 9 15 1 9 0 1 9 9 0 2
45 7 13 9 9 0 1 7 13 1 9 15 14 13 1 1 15 9 9 7 9 7 15 1 1 9 9 9 9 0 1 9 15 0 2 7 13 1 8 1 9 15 0 7 9 2
55 7 13 8 7 15 13 10 9 1 9 9 9 9 0 0 2 7 13 9 9 9 0 7 9 9 9 0 8 8 13 15 0 1 7 8 0 1 9 1 0 9 1 9 9 8 8 1 9 0 13 15 8 1 3 2
90 7 13 9 9 9 1 9 9 9 0 1 9 0 15 13 1 9 9 15 9 9 0 9 0 2 1 9 9 9 9 0 2 7 15 9 15 13 9 7 15 13 1 9 9 0 7 13 15 9 1 9 15 1 9 9 9 1 9 9 2 7 13 9 1 9 0 1 9 9 9 0 0 2 7 1 7 9 1 9 1 9 9 9 0 1 9 0 7 0 2
196 7 13 9 7 9 15 13 1 9 9 14 13 1 9 15 1 9 0 1 9 0 1 15 13 9 9 7 9 9 0 0 7 9 9 2 13 9 1 9 0 1 9 15 1 9 0 1 9 9 9 1 9 1 7 9 0 14 13 9 1 15 7 14 13 9 0 1 9 9 1 9 9 1 9 13 1 9 2 15 14 13 9 0 7 14 0 1 8 2 7 13 10 9 1 9 13 15 9 0 1 10 9 7 9 1 15 1 9 0 1 9 0 7 0 1 9 9 9 1 9 7 9 2 9 7 8 13 9 15 9 1 9 8 1 9 1 9 2 9 2 2 9 1 15 1 7 13 1 9 0 0 1 15 1 1 9 9 7 9 1 9 9 0 7 0 0 2 9 7 9 13 0 7 8 14 13 1 7 13 9 9 0 0 1 9 9 15 0 1 9 1 9 0 1 9 2
1 9
41 7 1 9 2 13 9 9 0 8 8 1 9 1 9 2 8 8 2 13 3 2 7 8 8 8 14 8 8 1 9 9 9 1 8 13 8 8 1 9 9 2
54 7 13 9 0 7 2 9 0 15 8 8 9 15 1 9 8 15 7 15 13 9 0 9 1 9 9 1 9 0 2 7 13 8 7 13 1 15 1 9 9 9 1 9 1 9 9 7 9 1 9 7 13 2 2
52 7 13 1 9 0 1 9 9 0 8 8 15 13 7 9 15 1 0 9 15 14 13 1 9 0 1 9 9 9 1 9 1 9 9 9 2 7 13 9 0 7 10 9 2 13 0 1 9 9 0 2 2
10 9 1 9 9 13 0 1 9 1 9
2 8 8
49 13 9 9 0 9 11 11 11 9 0 1 9 9 2 1 9 13 15 0 1 3 7 9 0 1 9 9 9 9 9 9 8 11 11 2 1 9 1 9 1 9 9 7 9 1 9 7 9 2
106 13 10 9 2 7 15 0 1 9 15 1 9 2 1 9 13 1 15 9 11 9 9 9 9 9 2 7 13 13 1 9 13 15 9 1 9 9 1 9 7 9 1 10 13 9 2 13 9 9 1 9 9 0 1 9 9 9 9 1 9 7 9 2 7 13 7 9 9 9 0 1 9 9 9 7 9 15 9 13 9 2 0 1 9 2 7 9 13 1 9 9 7 15 13 1 9 13 2 8 8 7 13 8 0 2 2
51 7 13 9 9 9 9 1 9 9 9 9 8 1 9 9 15 14 13 1 9 15 1 9 1 10 13 9 15 1 9 15 0 1 9 9 15 2 1 9 1 9 8 8 9 9 9 1 9 9 8 2
39 7 13 7 9 9 9 9 1 9 13 1 9 0 9 8 11 11 7 2 13 8 8 2 8 9 8 0 1 9 9 9 7 7 13 8 0 1 15 2
79 7 13 1 9 1 9 8 8 2 9 9 9 9 1 9 9 8 11 8 0 2 1 7 13 9 0 1 9 0 7 9 0 7 9 9 7 13 2 2 8 1 15 14 8 2 9 13 1 9 7 13 1 9 9 1 9 15 1 9 7 9 15 2 9 1 15 1 9 8 8 9 7 7 13 8 13 0 2 2
56 7 13 9 9 11 1 9 9 0 7 1 15 13 1 9 9 0 7 13 1 15 1 9 0 2 9 7 15 9 0 7 0 13 9 1 9 1 0 7 9 2 7 13 10 9 9 9 9 9 1 9 0 1 9 0 2
81 7 13 9 9 9 1 9 0 2 7 9 0 13 1 9 9 1 9 0 2 7 13 9 0 1 15 1 9 13 1 9 9 9 8 1 9 9 0 0 9 7 9 0 1 9 1 9 7 9 1 9 14 13 9 1 9 1 9 9 0 2 7 15 13 9 15 1 9 7 9 7 9 1 9 1 9 0 1 15 2 2
109 7 13 9 9 9 0 9 11 11 11 9 1 9 9 0 1 9 9 12 13 1 15 9 0 0 9 1 9 0 2 7 9 13 1 9 9 9 7 9 1 9 2 2 9 1 2 9 9 0 1 9 13 1 15 9 1 9 9 15 9 7 15 13 1 9 0 0 7 13 9 0 1 9 0 0 1 15 0 7 0 2 7 13 1 7 9 2 14 13 8 1 9 9 2 7 0 1 7 2 9 1 9 9 14 13 9 15 2 2
92 7 13 1 10 9 9 1 9 0 1 9 9 9 9 9 9 9 11 11 1 2 9 9 2 1 9 1 9 2 9 2 9 0 2 7 13 1 9 9 0 1 9 9 9 9 1 9 1 9 0 1 9 9 7 9 2 9 1 9 12 1 12 1 9 9 9 1 9 0 1 9 9 2 9 0 1 15 9 1 9 9 2 7 9 9 9 9 9 1 9 0 2
48 7 13 1 9 9 0 7 13 1 9 0 1 9 9 11 1 9 0 2 7 9 13 9 1 9 1 9 9 2 7 9 9 0 1 9 7 14 13 1 9 1 7 13 1 9 15 2 2
19 13 7 0 9 0 1 0 13 7 9 8 12 1 12 1 9 9 9 2
24 9 0 1 2 9 2 1 12 9 1 9 1 9 2 9 2 9 12 1 0 9 2 9 2
2 8 8
97 13 9 0 0 1 12 1 0 9 9 2 9 0 2 1 9 15 9 0 1 9 9 2 7 15 0 9 1 9 2 9 8 8 7 13 15 1 9 9 9 15 13 1 15 9 1 9 2 9 1 9 0 13 1 9 9 9 0 1 9 7 9 9 13 1 9 15 7 9 9 1 9 0 1 9 9 1 9 2 2 7 13 2 9 2 9 7 13 15 1 7 15 2 9 0 2 2
68 7 13 9 15 13 9 0 1 2 9 2 1 9 12 9 13 1 15 9 9 1 9 1 9 9 2 9 2 7 9 15 1 9 9 1 1 9 9 15 13 15 9 15 9 1 9 7 9 1 9 15 13 1 15 9 0 1 9 9 0 0 7 9 0 1 9 0 2
103 7 13 9 9 9 9 1 9 9 9 7 9 9 0 1 9 9 15 9 8 8 2 7 1 15 12 0 1 9 2 9 2 13 9 13 15 1 12 9 1 9 9 9 1 9 9 9 1 9 2 7 13 9 0 1 9 9 0 1 9 9 9 0 1 12 9 2 7 3 12 0 1 9 2 9 2 1 9 15 9 8 8 8 13 9 9 0 1 9 9 0 2 13 1 9 9 15 1 8 1 12 9 2
156 7 13 9 1 2 9 2 7 9 9 13 9 3 9 9 1 9 2 9 2 1 9 9 7 9 7 9 7 13 9 1 15 7 13 9 7 9 8 8 7 15 13 9 0 1 15 13 7 15 13 1 9 9 0 0 1 9 9 1 9 2 7 13 9 9 9 1 9 9 8 8 8 8 8 8 7 9 8 8 7 9 9 8 11 7 9 8 8 8 7 9 8 8 7 11 8 7 9 8 8 2 7 9 8 8 8 8 8 8 7 9 8 8 9 7 9 8 8 7 9 8 8 8 7 9 8 8 8 8 2 7 13 9 2 9 2 1 2 9 2 2 7 2 9 8 13 0 13 9 1 9 0 1 15 2 2
42 7 13 2 9 2 1 9 9 7 13 9 0 2 1 9 10 13 15 9 1 9 9 2 2 7 13 7 15 13 2 14 13 9 7 13 1 9 9 9 0 2 2
82 7 13 9 0 1 2 9 2 9 8 8 9 0 2 7 13 7 9 15 2 13 9 1 15 7 13 9 14 13 9 0 1 2 9 2 1 9 9 0 7 9 1 9 2 2 7 13 1 2 9 2 2 2 0 7 9 0 13 1 9 9 9 9 1 9 15 13 15 1 9 1 9 1 8 7 8 1 9 9 0 2 2
30 9 0 2 0 1 9 9 1 9 1 0 9 2 9 1 9 0 2 0 1 9 9 2 9 9 2 7 9 9 15
48 13 9 9 13 1 9 0 2 0 1 9 8 9 9 0 15 13 2 9 9 2 7 9 0 0 1 9 9 15 2 7 13 9 9 1 9 0 9 9 1 9 0 2 2 13 8 12 2
75 7 7 13 9 0 1 9 8 8 3 1 9 15 9 9 0 8 8 7 2 3 9 0 1 9 9 2 1 9 2 0 1 9 9 1 9 2 13 9 7 0 1 9 1 9 0 9 8 8 7 9 9 0 8 8 2 1 2 9 9 1 9 1 0 9 13 2 1 10 1 15 9 9 2 2
42 7 13 9 0 1 9 2 7 9 7 9 13 1 9 9 1 9 1 9 1 9 7 9 2 7 9 9 10 9 1 9 9 1 9 9 7 0 1 9 0 2 2
84 7 13 9 2 2 13 9 1 9 1 9 0 1 9 1 9 1 9 15 1 9 9 9 0 12 7 12 7 12 7 9 1 9 0 1 9 1 9 0 1 9 9 10 9 7 9 9 8 0 1 9 9 1 9 2 2 7 9 1 9 0 0 7 9 9 7 9 9 7 1 0 9 1 9 10 1 0 1 9 2 9 2 12 2
106 7 7 13 9 9 0 1 9 9 9 0 7 0 1 9 1 9 0 1 9 9 15 9 1 9 0 1 9 9 2 9 9 2 7 9 15 9 2 7 14 9 0 13 1 7 9 0 1 9 2 13 1 9 1 9 9 9 9 9 0 2 14 3 8 2 1 9 0 1 10 13 1 2 9 9 2 2 7 13 9 0 1 9 1 9 0 0 1 9 9 0 2 7 13 1 9 0 1 9 9 0 1 8 1 9 2
51 7 13 9 9 3 9 0 1 9 8 8 15 13 15 9 1 9 0 7 13 2 2 7 15 0 7 15 13 9 15 2 2 0 1 7 15 14 13 9 1 9 2 7 13 1 15 9 1 9 2 2
65 7 13 9 9 8 8 13 1 9 3 8 8 8 1 9 0 13 9 0 1 9 1 15 7 2 9 0 13 15 7 13 9 1 9 9 1 9 9 0 14 3 1 15 13 1 9 9 0 2 7 1 9 15 13 1 9 7 13 15 1 9 10 9 2 2
64 7 13 9 0 7 9 0 14 13 9 2 13 9 0 9 9 2 9 9 2 2 7 9 0 2 0 1 10 9 7 15 13 1 9 0 7 1 9 9 9 0 9 1 9 9 9 2 9 9 0 9 1 9 0 15 14 13 9 0 2 7 9 2 2
100 7 13 8 13 9 0 1 9 7 15 13 1 9 0 2 9 1 9 0 2 2 2 7 9 1 9 7 9 7 13 9 2 2 7 13 2 2 13 9 0 2 2 7 13 8 7 9 0 13 2 1 0 2 9 10 13 15 9 2 7 13 2 2 15 14 13 9 15 2 1 2 9 9 2 7 9 0 2 15 9 9 10 9 2 2 7 15 13 1 7 15 14 13 9 0 1 9 1 9 2
118 7 13 8 1 9 15 9 9 2 7 9 9 0 13 1 9 1 9 7 9 2 7 15 0 1 9 7 9 15 13 0 7 13 1 9 15 15 9 0 9 1 10 9 2 2 15 13 1 7 15 9 0 1 9 9 9 9 9 2 7 1 9 9 1 9 10 9 1 9 0 0 1 9 9 2 13 8 1 7 9 9 0 13 9 1 15 9 0 2 7 13 2 2 13 3 9 1 9 10 1 9 2 7 7 9 14 13 1 9 0 7 14 13 1 9 15 2 2
18 9 1 9 9 1 9 7 9 9 2 8 8 13 9 9 9 9 9
2 8 8
67 9 13 1 9 0 13 1 7 9 9 0 1 0 13 1 9 2 9 1 9 9 9 0 1 9 1 9 0 2 7 13 9 1 9 9 9 0 1 9 0 2 1 9 9 8 8 2 7 1 9 2 9 0 2 15 13 0 1 9 15 1 9 9 2 9 2 2
99 7 1 8 2 8 13 15 2 7 1 9 15 1 9 9 0 2 9 9 8 8 2 13 9 9 1 9 9 9 9 8 8 8 1 3 7 9 2 9 1 15 13 1 15 0 2 14 13 9 9 1 9 9 9 1 9 13 9 9 0 0 1 9 9 8 8 7 9 9 7 9 15 2 7 14 13 9 0 0 13 15 0 2 7 13 8 8 1 7 10 9 2 14 13 1 15 9 2 2
65 7 13 10 9 9 1 0 1 9 2 7 13 9 9 8 8 2 9 2 9 9 2 2 3 2 1 9 9 8 9 2 2 8 8 0 1 8 8 9 0 2 2 0 1 7 2 9 9 0 1 9 9 15 15 1 15 9 0 1 9 9 9 0 2 2
96 7 13 1 9 0 7 2 9 0 1 9 13 10 9 7 13 15 1 9 9 9 9 0 1 9 9 1 9 2 2 7 13 8 13 1 9 8 8 2 7 15 0 0 2 9 9 9 9 1 9 13 9 9 9 7 9 7 9 7 1 9 0 2 7 15 15 13 0 1 9 9 15 1 9 2 7 13 9 0 1 9 10 9 2 7 14 13 9 15 1 15 1 9 9 9 2
1 9
91 1 9 0 2 13 9 2 8 2 3 9 0 1 9 13 1 15 9 0 1 9 2 8 2 2 9 9 0 2 8 8 1 9 9 1 10 13 15 9 0 7 9 0 1 9 8 8 2 15 13 9 9 1 9 9 1 9 1 9 15 1 9 9 8 8 1 9 2 7 13 7 14 9 1 0 0 1 9 2 7 7 9 15 0 0 1 9 7 9 9 2
99 7 13 9 1 9 7 15 14 13 1 9 0 0 1 9 15 13 1 15 9 9 1 8 8 2 8 13 1 9 7 9 1 9 15 1 9 1 9 14 13 15 2 7 13 1 9 9 9 1 9 7 9 1 9 13 12 0 0 7 12 0 1 9 2 13 0 1 15 1 9 1 1 9 2 7 15 9 13 1 9 2 8 0 1 9 10 15 0 2 2 7 13 9 0 1 2 9 2 2
30 7 13 8 8 2 12 9 2 8 13 1 9 0 13 1 9 15 7 15 14 13 8 1 9 9 15 13 9 15 2
10 9 2 9 9 0 13 1 12 12 9
83 13 9 0 9 1 9 9 9 0 1 9 12 1 12 1 12 12 9 2 12 12 9 2 9 1 12 12 9 2 12 12 9 2 1 9 0 2 7 13 9 9 8 8 1 9 1 2 9 2 1 9 7 13 9 9 1 2 9 9 7 9 7 9 7 4 9 9 2 0 1 7 9 13 1 9 9 9 7 9 9 9 0 2
95 7 13 7 9 15 9 1 9 0 7 0 13 1 9 7 9 7 9 2 0 1 9 9 0 0 15 13 9 0 12 12 9 2 7 13 9 0 1 9 1 9 9 0 15 13 9 15 12 9 7 14 13 0 9 2 7 13 8 2 2 14 9 12 9 2 9 2 0 14 13 1 9 0 1 9 9 7 9 9 2 0 7 15 14 13 9 9 0 1 10 9 1 9 0 2
41 7 13 7 9 9 0 1 9 1 9 14 13 1 9 1 9 1 9 7 15 14 13 9 1 9 9 0 1 9 15 13 7 13 12 12 9 1 9 9 9 2
64 7 13 1 7 3 9 1 9 9 9 1 9 9 15 13 9 15 1 9 2 0 1 7 9 0 7 0 1 9 14 13 1 9 0 9 9 9 0 0 1 2 8 2 7 9 0 8 8 7 9 0 0 2 9 15 14 13 9 0 1 9 9 0 2
23 2 9 2 1 9 0 7 9 0 2 0 2 0 2 8 13 9 9 2 7 13 9 2
5 8 8 2 8 8
66 9 1 9 7 9 1 9 0 1 9 9 7 9 9 13 1 9 0 2 7 1 1 13 9 1 8 9 9 0 2 13 9 9 1 9 1 9 2 7 13 1 9 1 9 9 9 14 13 15 9 0 2 0 1 9 9 1 9 9 1 1 9 2 0 2 2
34 7 13 9 9 7 8 1 10 9 1 9 2 7 13 8 9 9 7 0 9 0 2 9 9 0 2 2 8 8 8 2 8 2 2
32 7 7 13 9 9 0 8 8 1 9 9 0 9 9 13 9 9 8 8 9 1 9 1 9 8 1 9 9 9 1 9 2
111 7 13 8 1 7 9 1 9 2 14 13 1 8 8 2 2 7 13 7 2 9 0 14 13 1 1 9 1 9 0 8 1 15 9 2 2 7 13 9 9 1 9 9 15 1 9 13 9 9 0 7 0 1 9 1 9 9 1 9 2 7 13 1 9 7 13 2 2 7 9 15 9 9 9 0 1 9 9 7 9 1 9 9 14 13 1 9 7 13 2 2 7 13 0 7 15 2 14 13 9 1 9 7 1 9 7 9 7 9 2 2
112 7 1 9 1 9 1 9 1 9 9 0 13 9 9 9 8 8 7 9 15 2 0 2 1 9 9 9 7 13 7 13 8 7 14 13 2 9 0 7 9 0 2 2 7 13 7 9 0 8 1 9 13 0 1 2 9 9 0 9 1 9 9 2 1 9 0 1 8 7 8 2 7 13 0 1 7 2 9 0 9 14 8 9 1 15 2 2 7 13 8 1 9 0 7 0 7 13 1 7 9 9 2 14 13 1 9 0 2 9 10 9 2
66 7 13 8 1 7 2 9 9 0 2 1 9 14 13 9 0 1 9 1 15 2 8 2 9 0 1 9 0 7 9 1 9 9 0 1 9 0 7 9 9 1 9 9 2 7 13 9 0 1 7 1 10 9 14 13 2 9 1 9 9 0 0 1 9 2 2
47 7 13 1 2 9 2 9 0 1 9 0 7 8 13 7 9 1 9 0 1 9 9 1 9 2 9 1 9 2 14 13 1 2 9 9 2 7 13 1 9 2 9 2 1 9 0 2
86 7 13 7 8 13 2 9 13 9 2 1 9 15 13 15 9 9 0 8 8 2 7 13 9 0 13 1 15 2 9 2 7 9 14 13 1 9 0 9 0 1 9 9 13 1 15 9 9 0 1 9 9 7 13 9 1 9 9 7 13 9 1 9 9 1 9 0 9 7 13 9 15 0 1 0 13 9 1 15 1 9 0 1 9 0 2
1 8
30 1 8 2 13 9 9 8 8 8 8 7 9 15 14 13 1 9 9 15 1 9 7 13 1 9 9 0 1 15 2
39 7 13 7 9 1 9 9 13 0 7 8 2 14 13 7 14 13 9 9 0 1 9 2 7 9 7 9 0 14 8 8 1 9 9 1 8 8 2 2
66 7 13 9 1 10 9 7 9 0 2 8 7 9 13 1 9 0 1 9 9 0 8 8 1 9 9 0 2 7 9 0 1 9 0 1 9 9 9 0 1 9 8 0 1 9 9 15 12 12 9 7 13 0 10 13 1 15 9 8 10 9 1 12 12 9 2
73 7 13 9 0 9 9 0 1 9 0 0 2 8 8 8 2 8 8 13 1 15 1 9 9 8 1 9 1 9 0 1 9 9 0 2 7 1 15 9 9 9 9 9 1 9 9 9 2 7 9 1 9 9 1 9 9 0 7 9 9 9 0 0 2 1 9 1 9 0 1 9 9 2
33 7 9 9 9 9 0 0 13 8 9 15 1 9 0 1 9 1 9 9 15 1 9 15 7 9 9 9 9 9 0 1 15 2
3 8 8 8
43 1 8 13 9 8 8 1 9 9 9 7 13 9 0 1 9 7 9 2 7 13 1 9 0 2 2 8 8 7 8 8 1 9 1 9 0 2 9 1 9 0 2 2
39 7 1 8 2 13 9 9 0 3 7 9 15 0 9 9 9 0 1 9 2 7 15 13 9 9 0 1 9 8 7 13 9 0 1 9 0 1 9 2
21 7 13 9 8 8 7 8 14 13 9 0 1 7 13 9 1 9 9 1 9 2
31 7 13 2 2 8 7 8 7 13 9 0 14 13 9 1 9 7 7 13 9 0 13 8 2 1 7 8 8 8 2 2
58 7 7 13 9 0 13 0 1 3 9 15 9 9 8 8 1 9 9 7 14 13 1 9 0 1 9 1 9 15 7 13 15 9 2 1 9 0 2 13 9 9 3 2 0 7 0 9 0 1 9 7 9 0 2 9 0 2 2
51 7 1 8 2 13 8 8 0 9 9 0 1 9 9 8 1 7 13 0 9 1 9 15 9 2 9 7 1 9 9 1 9 0 2 7 13 7 1 9 0 9 0 9 1 10 9 13 0 9 0 2
6 9 13 9 9 9 0
2 8 8
43 13 9 0 9 1 9 9 14 2 8 8 8 2 1 9 9 1 7 9 9 0 0 13 9 7 13 9 9 9 9 0 7 9 9 15 1 9 0 1 9 9 0 2
30 13 9 0 1 9 9 0 9 9 9 9 0 1 9 0 1 9 9 9 0 9 15 1 9 9 2 9 2 0 2
37 7 13 2 9 2 7 9 9 8 8 13 1 9 1 9 0 9 0 9 1 9 1 9 8 8 2 7 13 9 9 9 1 9 9 9 0 2
34 7 13 9 0 1 9 12 12 9 2 12 12 9 2 7 0 12 12 9 2 12 12 9 2 7 15 0 9 0 13 1 10 9 2
46 7 13 0 9 9 1 9 0 2 9 2 12 7 13 1 9 2 9 2 7 1 9 2 9 2 1 9 9 15 2 7 1 9 0 7 13 9 9 2 9 2 7 13 9 0 2
56 7 13 9 1 9 1 9 3 7 9 9 13 0 7 13 8 8 9 1 9 10 7 0 13 9 15 2 7 13 9 9 1 7 9 9 9 9 0 1 9 9 0 2 7 7 7 9 13 1 9 9 0 7 9 0 2
60 7 13 9 9 9 9 1 9 9 9 9 9 9 7 9 9 9 1 9 9 7 13 9 13 1 1 9 15 1 9 9 15 1 9 7 9 1 9 9 15 1 9 15 13 12 12 9 2 7 13 7 13 9 10 9 1 12 12 9 2
95 1 9 8 13 2 9 2 7 9 14 13 9 1 9 14 2 8 8 8 2 15 13 15 1 9 0 7 0 7 13 9 9 1 9 15 1 9 9 9 9 0 0 1 9 9 1 9 0 1 9 0 15 13 9 1 9 9 2 7 13 9 0 9 1 9 8 8 8 13 9 1 9 9 1 9 15 2 7 15 15 14 13 1 9 9 8 8 15 13 15 9 0 7 0 2
16 12 12 9 9 9 2 9 0 13 9 9 0 1 9 15 0
2 8 8
44 13 9 0 0 9 9 0 1 9 15 0 9 7 9 15 13 12 12 9 2 12 12 9 2 9 9 9 7 9 13 1 9 9 14 13 0 9 1 15 1 9 9 9 2
114 13 9 9 9 1 9 0 1 9 9 9 0 1 9 1 9 9 1 9 9 0 15 13 0 1 9 2 7 1 9 9 9 0 1 9 9 9 0 1 9 7 1 9 9 14 7 9 13 0 9 9 0 1 9 9 15 0 15 13 9 0 13 9 9 2 1 9 9 0 1 9 9 0 0 7 13 1 9 13 9 1 9 0 2 7 3 0 1 12 12 9 0 1 9 9 7 9 13 1 9 9 7 14 13 0 9 1 9 15 1 9 9 9 2
63 7 13 9 9 0 9 0 1 9 1 9 15 1 0 7 7 13 1 9 9 9 1 9 15 1 15 2 7 13 15 1 9 9 0 1 9 1 9 9 0 1 9 9 9 0 1 9 0 7 9 9 1 9 0 15 13 9 14 13 1 9 9 2
68 7 13 9 0 1 9 1 9 15 9 0 15 13 1 9 0 1 9 1 9 1 10 9 1 1 12 1 12 2 1 9 1 9 0 1 9 9 0 15 13 0 1 9 2 7 13 9 1 15 1 9 15 13 9 1 9 7 13 15 9 0 1 9 9 0 1 9 2
81 7 1 9 12 7 1 9 9 1 9 0 1 9 0 7 0 1 9 0 1 9 0 1 9 0 7 0 9 1 9 9 1 9 9 9 0 1 9 9 15 14 13 9 1 9 15 2 7 13 1 9 9 9 0 7 9 9 7 9 7 0 1 9 7 9 7 14 13 0 0 7 9 1 9 7 0 9 1 9 9 2
2 9 0
72 7 1 9 9 9 0 1 9 1 9 9 13 1 9 9 0 1 9 0 0 15 13 1 9 0 1 0 9 0 1 9 9 1 9 0 7 0 2 7 13 9 9 0 0 15 13 15 9 1 12 9 13 12 9 7 12 9 0 1 9 7 9 13 1 9 12 12 9 0 9 12 2
50 7 13 9 9 9 0 9 1 7 15 1 9 0 0 7 12 1 12 1 9 9 3 15 0 1 9 9 0 0 7 1 3 13 9 9 1 1 15 9 9 9 0 15 13 9 1 0 1 15 2
79 7 13 9 0 12 12 9 1 9 0 1 9 0 7 13 9 9 7 9 0 7 9 9 7 9 7 9 7 13 9 9 9 9 0 1 9 12 12 9 0 7 15 0 1 9 1 9 9 7 9 7 3 1 9 9 15 13 15 9 9 1 9 9 15 13 9 15 1 9 9 0 15 13 9 9 0 1 15 2
128 7 13 9 1 9 9 0 13 1 9 15 13 0 7 13 1 15 9 9 9 2 7 3 9 0 0 0 1 9 9 9 1 9 9 2 7 13 9 9 0 13 1 9 12 12 9 1 15 12 12 1 9 2 7 14 13 1 9 0 1 9 7 9 9 0 2 7 13 9 1 9 0 1 9 9 0 7 9 15 1 9 7 13 9 15 1 12 9 7 13 9 1 9 9 15 7 14 13 9 15 1 9 9 2 7 1 9 9 15 13 9 9 0 9 9 9 9 0 7 9 9 9 1 9 0 1 9 2
25 8 8 13 8 9 8 2 9 2 1 9 15 2 9 0 13 9 0 1 9 9 0 0 1 9
3 8 8 8
59 13 9 0 0 1 2 9 2 7 9 8 8 14 13 9 0 1 9 0 8 8 8 7 9 9 0 8 8 7 9 9 9 0 9 9 2 8 8 1 9 9 9 0 7 0 1 9 1 9 9 0 0 7 9 1 2 9 2 2
54 7 13 9 7 9 0 0 13 15 9 9 0 0 2 8 2 8 2 8 2 2 8 8 1 9 0 2 1 9 9 1 9 9 0 0 7 3 9 0 15 13 9 9 1 2 9 2 7 9 0 0 1 9 2
54 7 13 7 9 13 1 9 9 13 9 9 7 9 1 9 9 9 9 13 9 0 1 9 2 1 7 13 15 9 2 7 14 13 9 9 9 9 0 0 9 0 7 9 9 9 15 13 1 15 9 0 1 9 2
33 7 13 7 13 9 9 9 9 0 0 1 9 9 9 7 13 2 9 9 2 2 7 7 13 1 9 9 0 1 9 9 0 2
74 7 13 8 1 9 9 9 0 9 9 1 9 9 9 0 0 15 13 15 9 0 2 7 1 1 9 0 1 9 0 2 3 9 1 12 12 9 0 1 9 0 1 8 9 0 7 15 13 15 9 0 2 7 14 13 10 9 1 9 9 8 0 9 0 7 3 1 8 7 8 0 1 9 2
55 7 1 1 9 0 2 13 9 0 7 9 9 0 7 3 9 0 9 9 0 0 1 9 9 9 2 9 2 0 1 9 0 0 1 9 2 1 9 10 9 0 0 2 7 13 7 9 0 0 13 0 1 12 9 2
90 7 13 9 7 9 0 13 1 9 9 9 7 9 15 13 1 15 9 0 2 9 9 1 2 9 2 1 9 9 0 2 7 9 10 9 9 15 7 9 9 15 1 9 0 2 7 9 9 15 1 9 9 0 9 1 9 9 0 2 7 14 13 0 0 1 10 9 1 9 9 15 9 2 9 9 2 1 9 9 1 8 8 8 8 8 8 8 8 8 2
45 7 13 9 0 0 2 1 9 15 9 1 8 2 1 9 9 9 1 9 9 0 2 0 7 9 15 13 9 0 7 13 1 15 9 15 15 14 13 1 15 1 9 7 9 2
10 9 2 9 9 9 9 13 1 9 9
55 13 9 0 1 9 9 9 9 9 1 9 9 0 2 7 1 9 0 15 13 15 9 9 0 1 9 1 9 9 9 9 0 2 9 2 0 2 7 13 9 1 9 2 9 2 0 1 9 9 0 1 9 9 9 2
33 9 2 2 9 2 13 9 0 0 9 9 9 9 15 13 15 9 0 1 9 0 0 3 9 1 9 15 1 9 1 9 15 2
32 7 13 9 9 13 15 9 9 0 8 8 8 13 1 15 9 9 9 0 7 15 9 0 7 14 13 1 9 9 1 9 2
82 7 13 1 7 9 9 9 14 13 1 9 9 15 13 1 9 9 7 9 0 7 9 7 9 0 2 7 7 9 0 14 13 9 15 1 9 0 2 7 13 9 9 1 9 9 0 1 9 9 9 7 9 15 13 1 15 1 10 14 13 9 1 9 9 1 9 9 2 7 13 9 7 9 1 9 15 13 1 9 9 0 2
64 7 13 2 9 2 7 9 14 13 1 9 0 7 0 7 9 0 7 9 0 7 1 9 9 7 9 7 9 9 7 9 0 2 7 13 9 3 1 9 9 7 9 7 13 9 15 1 9 9 15 13 9 15 1 9 9 7 15 1 9 9 9 9 2
37 7 13 9 9 9 9 1 9 9 9 7 13 15 7 0 0 7 9 15 7 9 15 7 9 1 15 7 9 9 1 9 9 7 9 8 9 2
73 7 13 9 13 15 9 9 12 0 1 9 9 9 0 9 15 8 13 9 1 12 9 0 1 9 9 9 0 1 9 9 9 9 7 13 9 9 0 1 9 9 1 9 9 15 1 9 0 2 9 2 0 2 15 13 9 7 13 9 0 9 9 0 7 14 13 9 1 9 7 9 9 2
62 7 13 9 13 15 9 9 1 9 9 7 3 12 12 9 9 9 0 7 0 1 9 0 1 9 0 1 9 1 15 15 15 0 1 9 9 7 9 9 7 9 7 9 7 9 0 7 9 2 7 3 0 1 9 9 9 7 9 7 9 15 2
20 9 1 9 0 1 9 0 9 0 2 9 0 1 9 12 12 9 1 12 9
27 13 9 9 0 1 9 1 9 0 1 9 0 1 12 12 9 1 12 12 1 9 9 15 1 9 0 2
60 7 1 9 15 9 9 0 8 8 8 2 13 9 9 9 0 0 9 8 8 2 1 9 0 13 15 3 7 9 0 13 9 0 1 15 1 9 0 2 9 15 13 1 9 9 9 7 9 0 1 9 9 0 15 13 9 15 1 9 2
38 7 13 7 3 9 0 1 9 0 1 9 1 9 9 2 9 1 9 7 9 2 2 1 9 9 9 0 1 9 15 13 1 9 2 9 2 0 2
60 7 13 8 7 15 13 1 9 0 9 9 0 1 9 1 9 0 1 9 0 1 9 2 14 3 15 13 1 9 8 7 9 9 9 9 1 9 9 7 9 9 0 1 9 9 0 1 9 1 9 9 0 0 15 13 15 9 9 0 2
64 7 13 7 15 14 13 9 0 1 10 9 7 9 9 9 0 2 0 1 7 9 9 0 1 9 13 13 9 9 0 1 9 15 1 9 2 9 2 0 7 7 10 9 13 9 9 0 1 9 7 9 9 15 13 9 0 0 1 9 15 1 9 9 2
75 7 1 15 13 1 9 9 0 1 9 0 15 13 1 9 2 9 1 9 2 2 13 7 3 9 13 0 1 9 9 1 9 9 15 14 13 9 1 9 0 1 9 0 2 0 1 7 15 1 1 10 9 9 9 0 1 9 0 0 14 3 9 7 9 9 1 9 7 9 9 9 1 9 9 2
27 7 13 9 9 1 9 9 9 0 0 1 9 9 9 0 1 9 9 0 1 9 2 9 1 9 2 2
81 7 13 9 0 13 9 1 9 9 0 1 9 0 15 13 1 9 0 1 9 9 2 7 13 9 0 1 2 9 1 9 7 9 2 13 0 9 15 1 9 0 2 9 2 12 7 13 9 9 9 15 0 12 0 7 13 9 1 9 9 1 9 0 7 9 7 9 9 1 9 15 0 1 9 12 12 9 9 12 9 2
7 9 2 9 0 1 9 9
2 8 8
25 13 9 0 9 0 1 9 9 1 9 9 9 1 9 9 1 9 9 1 9 9 1 9 0 2
53 7 13 9 0 1 2 9 2 7 9 13 9 1 9 9 0 1 9 9 9 9 2 0 1 7 9 0 13 9 1 9 9 0 7 0 7 9 1 9 9 9 9 1 9 0 9 1 9 9 1 9 9 2
21 7 0 1 9 7 15 14 13 9 9 0 1 9 0 0 0 13 7 9 9 2
45 7 3 9 1 9 9 9 9 0 7 9 9 7 14 13 9 7 9 9 9 9 1 9 9 0 2 9 1 9 9 9 9 10 9 7 9 9 9 1 9 8 7 4 0 2
42 7 13 9 1 9 12 0 1 9 9 9 15 14 13 9 15 0 0 7 0 1 9 9 15 0 7 9 15 1 9 1 0 1 9 15 1 9 7 1 9 0 2
85 7 13 2 9 2 7 9 0 1 9 9 0 2 12 9 2 13 9 15 1 9 9 9 1 9 1 9 9 0 15 13 7 9 14 13 9 1 9 1 9 12 12 9 1 9 0 15 13 9 14 13 15 9 1 9 9 15 13 1 15 9 0 2 13 1 7 9 13 9 0 1 9 12 12 9 2 12 12 9 2 1 9 9 0 2
20 7 1 13 9 9 9 12 14 13 9 1 12 9 1 12 9 13 1 15 2
2 9 9
90 1 9 0 2 13 9 9 1 9 9 9 1 9 9 1 0 15 9 9 9 1 9 9 9 9 0 15 13 9 15 1 9 13 9 7 1 9 1 9 2 9 1 7 9 13 9 1 9 9 0 0 13 15 9 2 7 7 9 15 13 15 9 0 1 9 9 9 0 13 14 13 0 7 0 1 9 9 0 2 7 1 7 13 1 9 9 9 0 0 2
48 7 13 9 7 9 9 13 1 9 0 1 9 9 0 1 9 0 0 1 9 13 1 9 9 2 7 7 9 9 1 9 15 15 9 1 9 0 7 9 15 13 9 7 14 13 1 9 2
13 9 0 13 1 9 1 9 9 1 9 9 1 9
2 8 8
47 13 9 0 1 9 1 9 9 1 9 9 9 1 9 1 10 9 0 1 9 9 2 9 2 2 7 9 9 1 9 1 9 1 9 1 9 9 1 9 0 1 9 9 9 1 9 2
148 7 9 0 1 15 2 7 13 9 0 0 9 1 9 2 15 9 0 1 9 1 9 9 1 9 2 7 15 9 15 13 1 15 9 9 1 9 15 1 9 9 9 8 8 2 7 13 9 0 1 9 2 9 0 2 8 8 1 2 9 2 7 15 13 9 9 9 9 0 2 9 1 9 9 9 9 1 9 2 2 7 7 0 9 9 13 1 9 13 9 9 9 9 1 9 9 9 2 2 7 13 9 9 1 9 1 9 0 1 9 9 15 1 9 7 13 1 9 2 7 15 10 13 9 1 9 9 0 1 15 1 9 9 9 1 9 9 2 1 9 1 9 9 0 1 9 0 2
9 9 0 0 1 9 12 9 1 9
64 2 13 2 9 2 1 9 0 0 7 9 13 1 12 9 2 9 2 7 1 9 0 1 9 2 9 2 0 1 9 12 9 9 0 2 1 9 0 7 0 2 7 13 9 7 9 9 9 0 15 14 13 15 9 0 1 10 9 14 13 12 12 9 2
96 7 13 7 9 0 13 9 1 9 9 0 13 9 0 9 1 9 9 0 1 9 2 7 1 15 9 0 1 9 9 9 1 9 0 2 7 13 7 9 0 1 9 13 9 9 9 2 9 7 15 13 1 12 9 9 0 13 9 0 1 9 0 2 7 13 1 7 10 9 13 1 15 13 1 12 12 9 7 12 9 2 1 9 7 9 0 1 9 13 9 12 1 12 12 9 2
29 7 13 7 8 13 1 9 9 1 9 2 0 2 7 0 2 13 9 1 9 9 7 1 9 9 0 1 15 2
64 7 13 7 9 0 13 9 0 1 12 9 7 13 9 0 7 0 2 7 13 9 1 9 9 0 2 7 13 1 7 9 0 0 15 13 1 15 9 9 13 1 9 12 12 9 2 0 1 7 9 0 13 1 9 9 15 1 9 9 1 9 9 0 2
100 7 13 9 0 7 9 0 13 12 9 2 9 9 0 13 9 0 9 15 1 9 9 0 2 1 9 9 15 13 9 0 2 7 1 7 9 15 1 9 0 2 7 13 9 1 7 9 0 13 9 10 9 1 9 2 7 13 9 0 1 12 9 1 9 15 1 12 12 9 1 12 12 7 13 8 9 9 0 2 7 13 1 7 3 9 0 14 13 1 15 9 2 1 9 9 15 1 9 0 2
70 7 13 1 7 9 0 13 9 12 7 12 9 0 1 9 9 2 9 1 9 0 0 8 13 9 9 9 2 7 2 13 9 0 1 9 9 12 9 0 1 9 9 9 2 13 15 9 0 15 13 15 9 8 8 2 7 13 1 9 9 15 13 15 9 9 0 1 9 0 2
118 7 13 9 7 9 0 1 9 0 13 1 9 0 2 7 7 9 9 9 1 9 12 1 12 13 2 9 0 2 2 7 13 9 13 1 9 9 9 1 9 0 9 15 12 12 9 2 13 9 15 1 9 9 2 7 15 13 1 9 0 1 9 9 9 15 1 9 9 2 7 13 9 9 12 9 2 7 13 9 1 9 7 3 9 1 9 1 9 2 7 13 9 0 0 7 9 9 9 13 9 0 14 13 15 1 9 9 15 7 13 15 1 9 0 1 9 9 2
25 9 0 1 9 9 9 0 1 9 2 9 0 0 1 9 7 9 7 9 0 1 9 9 7 9
46 2 13 9 9 0 7 0 2 3 1 9 2 9 7 9 0 1 9 15 13 9 9 0 1 9 7 9 2 1 9 1 9 13 1 15 9 0 7 1 9 15 9 1 9 9 2
72 7 1 9 8 9 9 9 0 2 1 9 15 1 9 9 7 9 0 0 8 8 2 1 7 9 9 0 14 13 9 15 13 1 15 1 9 0 2 13 9 2 7 7 1 9 0 2 1 9 9 9 0 15 13 9 0 2 1 1 9 0 1 9 9 8 8 0 15 13 9 0 2
67 7 13 0 8 0 3 7 9 0 1 9 13 1 9 15 0 1 9 1 9 12 9 2 1 9 9 9 2 9 9 0 0 2 9 8 8 8 2 7 9 9 9 0 1 12 9 1 9 7 9 10 9 1 9 9 0 13 1 9 0 13 9 15 1 9 15 2
44 7 1 9 15 13 9 1 7 9 0 13 0 7 15 8 1 9 0 1 9 2 7 1 9 7 9 0 14 13 1 12 12 9 13 9 0 1 9 1 0 1 12 9 2
72 7 14 13 9 8 8 9 1 9 1 9 9 0 0 9 15 1 9 7 9 2 7 15 13 7 9 15 13 9 15 1 9 12 9 13 1 9 9 9 1 2 9 9 0 2 9 12 2 9 1 7 9 0 1 9 0 2 0 13 1 9 9 1 9 1 9 9 0 0 1 9 2
53 7 13 3 1 7 9 9 0 1 9 9 9 0 0 13 1 9 0 0 2 0 1 15 9 9 0 1 9 12 1 12 0 1 9 0 0 2 7 13 1 7 15 13 9 9 9 1 9 9 9 0 0 2
56 7 13 9 0 2 1 9 9 15 2 1 9 9 1 9 0 1 9 7 9 2 0 2 1 9 2 9 1 9 0 7 0 13 1 9 9 0 2 7 13 1 9 9 15 1 7 14 13 9 9 0 1 9 9 8 2
60 7 13 1 7 9 0 13 1 9 0 1 9 0 7 9 15 13 1 9 9 0 2 0 7 14 13 9 0 0 2 2 14 3 7 13 9 0 1 9 9 9 0 1 9 9 9 1 9 1 9 9 9 1 9 1 9 15 13 15 2
69 7 13 7 15 4 3 9 1 9 9 9 9 0 2 0 7 9 9 9 15 9 2 7 7 9 0 14 13 9 1 9 9 7 9 7 13 1 9 9 0 2 7 13 1 7 3 0 9 0 1 9 1 9 9 13 1 12 9 1 9 15 13 12 1 12 9 7 9 2
77 1 9 15 2 13 2 9 0 1 9 2 1 9 13 15 7 0 9 9 0 1 9 13 1 9 0 1 9 0 7 9 9 9 0 1 9 9 9 9 0 2 9 9 9 7 9 9 0 0 2 7 9 9 9 0 1 9 15 0 1 9 8 2 9 1 9 9 9 9 1 9 7 9 15 1 9 2
44 7 13 9 9 9 0 1 9 1 0 9 2 8 2 8 0 2 8 0 2 7 9 1 9 0 1 9 15 13 9 15 1 1 9 9 0 1 9 7 9 15 1 9 2
28 9 0 14 13 9 9 0 7 13 1 9 9 9 9 2 8 13 9 9 7 8 1 9 15 1 9 9 0
83 2 13 9 0 1 9 0 1 9 9 1 9 9 2 9 2 7 8 13 1 9 8 9 0 1 9 9 15 7 9 9 1 10 9 1 9 9 15 1 9 9 1 9 9 2 7 13 7 9 0 13 1 9 9 0 1 9 0 1 9 1 9 8 2 8 2 15 13 9 1 9 0 0 7 9 1 9 9 1 9 13 9 2
109 7 13 9 0 0 8 8 3 9 1 0 9 0 13 1 9 9 0 1 9 0 9 1 9 0 7 2 9 0 1 9 9 2 1 8 1 9 0 2 2 13 8 12 2 2 7 13 9 0 9 9 9 7 9 9 9 1 15 2 7 13 2 9 2 7 9 9 9 9 8 8 13 9 9 15 13 8 8 8 8 11 7 9 8 8 8 2 7 13 9 2 9 0 2 11 8 7 13 1 15 8 8 8 8 8 8 8 8 2
90 7 13 9 8 7 9 8 1 9 9 9 9 1 9 9 9 9 9 15 13 9 0 12 9 1 9 9 1 15 2 1 9 13 1 15 1 9 0 9 1 9 9 9 2 7 13 9 9 9 0 0 0 9 1 9 9 9 12 2 7 13 9 1 9 10 9 1 9 1 9 7 15 9 0 1 9 9 9 9 15 13 7 13 15 9 1 9 9 0 2
82 7 13 9 0 1 9 7 8 13 1 9 15 1 9 9 7 13 15 1 9 2 7 13 7 9 0 1 9 13 1 9 0 0 2 7 13 0 1 15 1 9 9 9 1 9 9 7 9 9 2 9 0 2 1 9 13 12 9 2 7 13 8 9 8 8 1 9 1 9 9 8 8 13 9 1 15 9 0 8 8 8 2
182 7 13 7 9 0 15 13 9 15 1 9 0 13 1 9 9 0 13 9 9 0 7 9 9 0 0 7 9 9 2 7 13 7 15 13 9 1 8 9 9 0 1 9 9 1 9 9 2 7 13 1 9 1 9 9 9 1 9 15 13 1 15 9 9 15 0 7 9 15 0 15 9 2 14 13 9 9 1 10 9 2 2 7 13 9 13 15 1 9 15 1 8 1 9 1 15 9 15 7 15 13 9 9 9 0 1 9 0 2 7 13 2 2 14 9 13 8 7 13 9 9 1 9 15 2 15 9 14 13 0 9 1 8 2 2 7 13 1 9 9 9 15 9 9 0 7 13 2 2 7 8 1 8 8 8 7 2 3 9 1 9 9 2 7 1 9 9 14 13 1 9 9 0 7 14 8 8 14 13 0 2 2
14 0 2 14 13 2 1 9 2 9 2 7 2 9 2
53 2 13 0 7 15 2 14 13 2 1 9 2 9 9 0 2 2 8 2 7 9 2 9 0 2 9 8 11 8 2 7 15 2 0 2 1 9 15 0 7 2 13 1 9 9 9 15 7 9 9 15 2 2
64 7 13 9 1 9 0 0 0 1 9 9 1 15 9 9 0 8 8 8 2 7 0 2 13 1 9 7 9 9 2 0 7 13 0 1 9 1 0 1 9 15 7 9 15 0 1 9 9 9 15 7 9 9 15 2 7 15 1 9 9 9 0 2 2
57 7 13 8 7 9 8 8 13 9 0 7 0 9 9 15 1 9 1 9 7 2 0 13 13 9 7 13 15 1 9 15 1 9 15 13 9 0 7 9 13 1 9 9 1 9 9 2 9 15 13 7 13 0 1 9 2 2
37 7 13 7 9 9 0 8 8 2 13 9 0 1 9 15 1 9 15 0 7 9 15 0 2 15 7 10 9 13 8 1 9 1 10 9 2 2
37 7 13 9 9 9 0 1 9 2 9 2 8 8 1 9 2 9 0 2 8 11 8 2 7 13 9 9 11 8 7 13 1 15 1 9 0 2
14 9 1 9 9 0 7 9 9 9 0 1 9 9 9
77 2 13 9 0 1 9 1 9 12 1 9 1 9 1 9 9 0 15 9 1 9 2 9 9 2 7 13 9 9 7 9 0 2 7 13 9 0 7 1 9 9 9 1 9 9 0 1 9 9 15 1 9 9 0 7 13 1 9 9 0 1 9 9 0 7 9 9 0 1 9 0 1 9 0 1 9 2
137 2 13 9 9 9 9 0 0 1 3 1 9 1 12 1 12 9 2 9 9 9 0 1 9 9 9 0 1 9 1 9 0 0 2 7 7 13 9 0 9 9 0 1 9 13 1 0 1 9 1 9 9 0 1 1 7 13 1 15 9 1 9 0 1 9 9 15 13 15 1 9 9 9 2 7 14 10 9 3 15 13 9 15 1 9 0 1 9 9 15 13 1 8 7 9 9 13 9 1 9 7 13 9 0 7 0 15 9 9 9 9 1 9 7 15 10 13 3 2 7 13 9 9 9 1 9 9 0 1 12 9 1 9 0 1 9 2
46 7 13 9 0 1 2 9 2 1 9 9 0 1 9 0 1 9 0 1 9 15 9 0 1 9 9 0 15 13 9 1 9 9 0 1 9 12 12 9 1 9 2 9 2 0 2
5 9 9 1 9 9
149 7 13 9 9 2 9 2 1 9 1 9 9 0 1 9 7 13 9 15 1 9 0 7 9 9 7 9 9 1 9 9 2 9 1 9 9 9 0 1 9 1 9 15 13 1 15 9 0 1 9 1 9 9 9 7 15 2 15 13 1 9 9 2 0 2 1 9 0 2 7 9 9 9 9 0 1 9 1 9 1 9 9 7 9 9 0 2 15 13 9 1 9 1 9 9 1 9 9 9 1 9 9 0 7 9 1 9 1 9 0 1 9 12 12 9 1 9 9 0 2 7 15 10 13 9 1 9 15 1 8 7 13 9 1 9 9 0 1 9 2 9 2 0 15 13 9 9 9 2
2 9 9
125 14 7 9 1 9 9 13 9 0 1 9 15 13 1 9 1 9 7 9 0 2 7 14 13 9 0 7 14 13 1 9 9 15 13 1 15 9 15 9 1 9 9 2 7 2 9 2 9 1 9 0 7 9 9 9 15 1 9 9 7 9 2 7 9 9 15 1 9 9 0 7 13 1 9 9 0 1 9 9 0 7 9 9 0 1 9 0 1 9 0 1 9 2 1 9 9 9 9 1 9 0 1 9 14 12 1 12 7 14 13 9 9 1 9 0 2 7 9 0 13 1 9 0 9 2
90 1 10 9 13 9 1 7 9 0 1 9 9 0 13 1 9 1 9 9 9 9 14 13 15 9 0 7 9 0 13 9 1 9 13 1 9 1 9 0 9 0 2 9 7 9 9 15 13 2 0 2 1 9 15 1 9 1 9 9 9 0 1 15 1 9 12 1 12 2 14 13 0 9 1 9 9 9 0 15 13 0 9 1 9 9 7 0 1 9 2
18 15 13 14 9 1 8 7 8 1 9 14 13 7 13 9 1 8 2
64 14 0 7 9 2 8 8 2 2 8 9 0 1 9 1 9 0 9 1 9 9 0 13 8 8 9 8 1 9 1 9 9 7 7 10 9 15 8 13 9 7 9 1 15 7 13 15 1 9 1 9 1 2 8 8 2 1 9 8 8 8 8 8 2
133 8 10 9 1 2 8 8 2 9 15 13 1 9 8 8 7 9 0 13 9 15 1 9 9 1 9 9 8 8 9 0 1 9 2 7 13 9 9 0 0 1 2 9 9 2 1 7 13 1 9 9 8 8 8 9 8 7 13 1 7 8 0 14 13 1 7 13 1 15 8 0 2 7 13 8 9 10 9 1 9 9 7 9 9 9 0 1 9 9 0 8 8 15 13 9 0 15 8 13 1 2 8 8 2 1 9 1 8 8 14 13 0 1 9 7 7 8 0 8 1 9 7 7 1 2 8 2 7 13 9 15 0 2
130 3 7 9 9 8 8 14 13 8 8 9 0 1 2 8 8 2 7 13 1 9 0 1 15 2 2 8 8 8 9 8 8 1 9 10 9 2 7 13 8 8 1 2 9 2 15 8 1 8 0 1 9 8 8 8 8 1 9 9 1 9 2 7 13 2 8 8 9 9 15 13 1 9 1 8 2 8 8 2 1 9 8 8 2 9 9 8 8 8 8 0 7 7 13 7 13 1 10 9 1 15 7 13 8 8 2 7 7 9 1 8 2 8 2 13 1 9 9 2 7 15 14 13 8 8 1 7 13 2 2
14 9 2 8 8 2 13 1 10 9 8 8 1 0 2
36 0 2 7 8 8 14 13 9 1 8 2 8 8 2 7 14 2 8 2 15 1 0 8 8 7 2 9 2 1 8 7 9 8 1 15 2
169 0 2 7 8 8 15 1 8 8 13 1 15 7 15 9 0 1 15 2 7 15 13 7 15 8 0 7 1 9 0 0 1 8 1 15 2 8 7 9 1 8 7 8 7 13 9 9 8 8 7 7 15 13 1 9 1 9 9 2 7 3 0 1 9 1 10 9 1 9 9 0 1 8 9 12 7 9 1 9 9 2 7 7 13 9 9 9 9 0 8 8 9 2 1 9 13 9 1 2 8 2 7 13 1 9 1 8 7 9 1 15 7 13 9 15 7 9 1 15 2 13 7 8 15 9 9 0 15 13 1 8 1 8 0 7 13 1 15 1 8 0 2 7 14 13 10 9 9 8 8 8 9 9 8 8 1 8 8 7 15 9 13 7 15 14 13 7 13 2
55 7 14 13 9 9 0 8 8 1 9 15 1 9 9 2 0 1 9 9 0 1 8 7 13 9 9 0 1 9 1 9 9 9 1 9 7 13 13 7 9 13 1 9 1 9 9 9 7 9 0 0 1 9 15 2
55 0 2 7 8 9 1 9 1 9 7 1 9 1 9 2 14 13 9 7 14 13 1 9 9 8 8 2 7 13 1 9 9 7 9 15 13 1 9 2 1 15 13 9 9 9 8 7 15 14 13 8 7 14 9 2
58 0 2 7 9 9 8 8 8 13 1 9 1 15 1 9 1 8 2 7 9 8 8 13 7 15 1 8 9 1 9 0 1 9 15 1 8 2 7 15 13 1 7 8 14 13 13 1 15 2 7 1 9 9 15 1 8 2 2
75 7 13 2 7 8 9 14 13 1 9 7 15 13 8 8 2 7 1 9 9 7 8 2 13 7 13 1 9 0 1 9 0 2 8 14 13 1 0 7 14 13 1 9 1 0 2 8 8 1 15 15 8 1 9 1 9 1 15 1 9 0 2 7 8 14 13 1 9 15 1 8 1 9 2 2
101 7 13 9 9 15 2 2 7 13 15 15 9 9 0 2 0 2 7 1 10 9 9 1 9 9 9 1 8 10 13 9 0 2 9 1 9 9 0 2 0 7 1 9 9 9 0 1 9 7 7 13 8 15 9 0 2 7 15 13 8 14 13 15 8 1 15 14 13 1 15 9 1 9 0 2 3 9 9 15 2 7 15 13 1 0 2 7 14 13 9 8 8 8 8 7 15 14 13 1 15 2
116 1 15 13 9 2 8 8 2 9 8 8 1 9 1 15 7 15 14 13 1 9 9 0 1 8 7 7 9 9 0 1 8 7 8 13 9 0 0 8 8 0 1 9 9 0 1 9 9 7 1 15 2 8 8 8 1 9 2 9 2 1 8 7 1 2 9 0 2 7 2 9 2 8 8 0 0 15 1 8 9 15 2 7 14 0 8 8 14 9 1 7 9 7 9 1 15 13 1 8 1 1 9 0 2 7 15 7 1 9 9 7 9 7 8 0 2
109 8 8 9 2 8 8 2 1 15 7 8 0 7 0 8 13 2 8 2 7 9 15 1 9 1 9 0 1 8 2 15 9 15 13 7 9 14 13 1 8 7 7 9 9 8 8 8 8 1 15 1 9 9 8 8 2 7 7 1 9 0 0 8 0 1 15 2 7 14 13 9 0 1 9 7 1 9 2 7 15 15 8 8 13 9 0 7 13 9 15 1 9 2 7 14 13 8 9 9 7 9 1 8 7 15 15 9 0 2
44 7 9 9 9 1 8 9 7 9 9 1 9 9 0 2 15 1 9 2 8 8 2 1 9 9 15 7 9 7 9 1 15 1 9 13 9 7 13 15 1 9 13 14 2
4 9 9 0 2
43 13 9 0 9 9 1 9 7 9 1 9 10 2 13 1 9 15 1 9 7 13 9 1 9 2 7 7 15 14 13 0 15 14 13 9 15 14 1 9 9 0 0 2
76 7 7 13 9 9 0 1 9 13 1 9 1 9 9 15 8 8 8 9 1 9 1 9 9 15 1 9 0 2 7 14 9 0 1 9 13 8 1 9 10 9 8 8 1 1 9 15 9 9 0 1 9 0 9 8 8 8 1 9 0 14 13 15 3 8 8 8 8 9 9 1 9 9 7 0 2
60 7 9 0 13 1 9 0 1 9 7 1 9 9 15 2 7 15 9 13 1 15 9 1 9 0 1 9 10 13 1 15 1 9 7 13 1 15 1 9 2 7 3 9 1 9 10 13 1 9 9 15 9 0 7 14 13 1 9 9 2
114 1 9 0 1 9 2 13 9 13 9 0 9 2 13 9 8 8 0 15 7 15 13 9 2 9 2 0 0 9 1 9 9 15 13 8 7 7 8 2 0 1 9 0 9 8 9 1 9 9 0 1 9 2 13 9 0 1 15 1 7 14 13 15 9 2 7 13 8 8 9 7 9 13 1 9 1 9 15 13 15 8 1 8 2 13 8 7 13 9 0 2 8 8 8 8 9 2 9 0 13 9 8 8 2 7 9 8 9 1 2 8 8 2 2
90 13 9 8 0 0 7 14 13 1 9 8 0 8 8 1 9 2 7 7 2 8 2 0 13 9 8 8 1 9 2 7 13 8 2 12 3 1 8 9 1 9 2 7 7 9 0 8 14 14 13 9 10 9 2 7 7 14 13 8 1 9 7 9 9 9 1 9 0 8 8 1 15 13 9 1 8 2 12 7 15 1 9 9 9 12 9 1 9 9 2
97 13 9 0 1 9 9 0 0 2 7 15 13 8 8 1 9 8 8 1 9 2 7 14 13 2 8 2 1 9 7 13 8 8 8 8 0 0 1 9 0 2 13 2 9 2 9 8 8 1 9 9 8 1 9 1 9 9 9 0 8 15 13 8 8 8 9 7 9 1 15 2 13 9 1 9 15 1 8 8 0 8 2 1 9 8 8 8 8 8 1 9 7 15 13 8 8 2
132 14 8 1 9 2 7 15 1 9 15 0 4 1 9 9 9 1 9 8 8 7 1 9 15 8 9 1 9 9 1 9 2 8 8 9 9 13 9 2 8 8 9 9 7 2 8 8 2 13 15 13 1 9 15 7 13 1 8 9 0 1 15 1 0 2 7 13 9 8 8 1 9 9 1 9 7 13 15 1 9 0 1 9 0 8 9 8 1 9 1 9 15 0 2 1 15 13 1 9 9 8 15 9 0 0 2 9 7 9 13 9 1 0 9 1 13 8 1 9 1 9 15 0 1 2 9 9 2 1 9 15 2
31 13 9 13 1 9 7 7 13 1 15 9 9 1 9 9 15 2 7 15 15 9 0 1 9 0 2 7 9 13 9 2
2 8 8
3 8 2 12
74 0 7 8 8 13 1 9 8 1 9 9 9 2 0 7 15 0 7 0 2 7 7 15 13 9 0 14 13 9 9 0 8 8 0 2 8 13 0 1 9 15 9 1 8 2 9 8 2 2 8 8 8 1 9 13 9 1 9 7 3 2 7 1 9 13 9 8 7 13 0 1 8 8 2
50 14 8 1 15 13 9 7 13 8 2 12 1 9 0 1 9 8 8 2 1 9 15 8 8 8 2 7 2 9 2 8 8 8 1 9 1 9 0 2 8 8 9 1 2 9 8 2 12 2 2
82 9 9 9 9 1 9 8 8 2 1 9 7 9 9 9 2 2 2 1 9 9 1 15 13 9 14 1 15 13 15 2 8 8 8 9 7 13 2 9 8 2 12 2 1 8 13 9 1 15 1 7 9 13 9 7 9 2 7 1 7 8 13 1 15 8 14 13 1 9 15 13 8 9 1 9 15 8 8 9 2 2 2
76 13 0 7 8 8 13 15 9 9 8 1 3 2 7 15 14 13 1 9 0 2 14 13 9 15 1 8 8 8 8 8 8 1 9 9 2 9 9 9 1 7 1 9 0 9 15 13 7 13 9 15 1 9 2 7 9 7 9 0 0 13 9 0 8 9 1 8 2 12 7 1 15 1 9 9 2
29 15 13 9 7 13 9 8 9 1 9 7 9 8 2 7 15 14 13 9 2 9 0 1 9 1 9 9 0 2
54 7 15 13 15 7 13 9 8 8 8 8 8 0 2 8 13 9 7 15 13 9 9 9 8 8 2 7 15 13 1 0 9 9 8 8 9 0 1 15 13 9 9 1 9 0 15 15 9 0 1 9 8 8 2
63 9 13 3 15 13 8 1 10 9 2 8 8 14 13 0 3 7 13 15 7 13 3 9 9 0 2 7 13 9 0 9 1 7 1 9 15 7 13 1 8 2 12 8 8 9 8 8 2 9 9 1 9 9 8 0 8 8 8 13 7 13 8 2
92 9 1 9 10 2 14 8 7 8 7 8 13 1 8 8 8 8 8 1 9 2 8 9 1 9 8 8 8 8 2 9 8 2 12 2 7 9 8 9 0 2 8 8 9 1 9 1 9 8 8 1 9 2 1 15 13 2 9 9 9 2 2 7 1 15 13 8 8 9 8 8 8 8 8 8 8 8 8 8 8 8 2 1 7 8 1 0 7 13 1 15 2
144 7 14 8 3 7 8 7 8 9 1 9 9 8 8 8 7 13 0 1 8 9 2 7 14 9 1 8 15 13 15 1 9 9 8 2 12 7 15 13 15 1 9 7 15 14 13 15 7 13 15 2 1 9 7 8 13 1 9 15 0 7 13 9 0 2 1 7 8 2 12 15 0 9 1 9 7 7 13 7 7 8 13 9 2 7 13 7 9 0 13 9 9 1 9 9 9 0 2 7 7 15 13 8 0 2 8 8 8 1 9 9 9 8 8 8 7 9 8 2 15 13 1 1 9 2 8 0 1 9 2 7 15 2 13 0 7 0 8 8 9 8 2 2 12
51 8 13 9 9 1 9 15 8 1 3 1 15 13 9 13 8 8 1 8 13 1 9 7 13 15 8 2 7 1 15 8 9 1 8 8 2 12 1 7 15 1 2 9 2 8 9 7 9 7 9 2
53 7 13 8 8 8 1 9 15 13 15 9 2 1 15 13 9 9 13 9 8 15 9 0 2 7 13 9 1 9 1 9 15 2 7 7 15 13 1 9 8 8 14 13 1 15 9 8 8 8 7 13 13 2
25 14 1 1 8 8 8 14 13 1 8 8 8 2 13 9 9 15 9 1 9 2 9 7 9 2
54 2 8 8 8 1 8 8 8 8 9 7 8 15 8 8 8 8 8 8 8 2 7 1 9 0 7 8 8 8 2 2 2 2 2 8 8 8 8 1 15 7 13 8 8 7 1 9 0 7 13 1 9 15 2
17 2 8 2 13 9 9 2 0 2 2 13 1 8 9 1 8 9
88 13 2 8 2 3 7 13 8 8 1 9 0 1 9 9 1 9 9 9 1 9 13 9 9 0 2 2 9 8 8 2 1 9 8 8 9 1 9 0 15 13 9 15 2 7 0 7 8 2 7 15 1 9 8 8 2 14 13 1 8 9 2 1 9 9 8 8 8 9 9 9 2 8 8 1 9 1 9 9 0 0 1 9 0 8 8 9 2
62 7 13 9 1 7 8 1 9 9 15 2 13 1 9 9 9 9 1 9 15 13 15 9 1 2 8 2 7 2 8 2 2 7 1 9 13 1 7 9 15 14 13 1 9 2 7 14 13 9 9 8 8 2 7 14 13 3 9 1 12 9 2
66 1 9 0 13 2 8 2 9 9 1 9 9 9 2 9 2 1 9 2 7 13 8 8 9 1 9 2 2 9 8 2 13 1 15 2 2 13 9 9 3 9 0 0 1 9 15 2 9 9 0 9 1 15 7 13 15 1 9 15 2 13 3 1 12 9 2
101 7 1 9 7 0 8 15 9 9 14 13 1 9 2 7 1 8 9 9 9 0 8 2 8 8 8 8 9 0 1 9 0 2 8 8 1 9 1 9 8 9 8 8 8 13 8 8 2 9 9 1 15 7 15 13 7 13 1 10 9 14 13 9 9 0 2 8 8 3 15 14 13 1 8 8 3 15 14 13 9 15 1 9 9 0 2 3 7 13 9 9 2 7 14 13 1 15 1 9 15 2
70 8 13 9 9 8 9 0 7 0 2 8 13 8 8 9 15 1 8 1 9 8 8 2 7 13 9 15 13 1 9 2 7 13 9 15 0 9 0 2 7 13 9 15 1 9 1 15 13 9 0 1 8 7 13 9 15 1 9 9 0 2 7 3 1 15 13 9 9 8 2
149 7 14 13 1 9 8 9 9 1 9 15 1 9 2 7 1 9 13 9 9 9 2 7 13 8 8 8 8 1 9 2 1 15 13 1 15 8 8 9 9 2 9 1 9 13 1 9 15 0 2 7 13 8 9 15 8 9 0 1 9 15 0 8 8 8 0 2 3 1 9 13 9 1 9 9 2 7 13 1 8 8 8 1 9 9 2 7 9 15 14 13 9 1 8 8 0 8 8 11 8 8 8 8 8 1 9 9 1 9 0 2 7 8 8 13 1 9 1 9 0 14 13 1 9 7 0 15 14 13 1 15 9 0 1 9 9 7 9 8 8 2 1 1 9 1 9 9 2 2
8 1 13 9 2 2 2 1 9
52 3 2 13 9 7 15 13 2 13 1 9 2 14 2 7 15 1 9 13 2 7 1 9 10 13 9 1 9 15 1 9 2 13 0 7 9 9 13 2 7 7 9 0 1 9 7 0 15 14 13 15 2
152 14 13 1 10 9 0 1 9 13 9 1 9 7 15 13 1 15 2 7 2 7 1 1 8 9 9 1 9 0 2 7 7 13 9 9 8 8 1 0 9 1 15 2 13 9 1 7 9 13 9 8 8 9 9 15 2 9 9 15 1 9 8 8 2 9 8 8 8 8 8 2 7 15 1 9 13 9 1 10 13 8 8 2 7 13 8 8 2 8 14 15 9 0 9 8 8 2 7 7 3 8 1 15 9 2 7 7 13 8 1 9 13 1 9 8 8 8 8 8 8 2 14 7 15 13 1 0 9 1 9 8 9 8 8 2 7 4 13 1 9 9 9 9 2 7 15 8 13 1 15 9 2
124 14 9 9 1 9 2 7 14 9 8 8 8 1 9 1 9 15 2 13 1 15 9 9 7 9 0 15 13 1 9 0 7 9 9 2 1 10 2 2 2 9 1 8 2 9 0 2 15 13 7 15 13 1 9 9 14 1 15 13 1 9 2 7 1 1 7 8 2 8 8 2 8 2 7 1 15 8 13 4 3 8 8 8 13 9 9 0 2 7 13 1 9 8 8 10 9 1 0 9 1 9 0 2 14 1 0 15 14 9 7 13 9 0 1 9 13 1 9 15 9 9 7 9 2
127 8 8 9 1 9 9 0 8 8 2 13 8 8 9 0 8 2 7 13 8 9 15 13 1 9 1 9 2 1 9 7 9 13 1 2 9 0 2 2 7 13 1 8 8 9 0 2 0 1 9 9 9 1 9 7 0 8 9 9 1 15 8 0 1 8 8 13 1 15 9 9 2 7 13 8 1 7 13 9 1 9 15 13 14 13 1 15 15 9 15 8 15 14 13 1 15 1 9 1 9 9 2 9 1 9 9 2 8 8 8 1 8 8 7 13 14 13 15 1 9 1 9 1 10 9 0 2
160 14 8 8 14 13 0 2 7 9 1 15 13 1 15 13 8 8 8 2 7 14 13 8 1 8 0 15 1 15 8 8 2 8 13 9 8 8 8 15 13 13 9 0 2 9 14 13 10 9 9 1 2 9 9 2 8 8 2 9 0 0 2 0 2 2 7 9 8 9 0 8 13 7 14 9 0 1 15 9 7 13 9 9 15 8 1 9 15 2 14 9 9 13 1 15 9 0 1 15 8 8 8 1 9 15 2 7 14 9 2 7 15 13 2 9 14 13 8 8 14 9 9 2 7 14 8 8 8 1 15 9 2 8 8 14 13 15 14 0 2 7 15 13 1 15 8 9 2 14 13 1 15 9 1 9 7 14 15 13 2
21 13 1 9 9 9 8 9 9 8 8 2 13 9 9 0 1 9 9 9 0 9
50 13 9 9 8 8 7 9 9 14 13 9 1 9 1 8 8 0 2 0 7 9 9 8 2 12 13 1 9 9 9 9 0 7 1 1 0 9 1 9 0 2 0 7 8 13 9 1 15 8 2
45 7 13 9 15 7 9 15 13 1 15 8 14 13 0 9 0 1 9 7 2 15 9 9 8 8 0 1 9 0 8 8 8 0 8 8 0 1 9 0 8 8 8 0 2 2
68 7 13 8 1 9 13 3 8 1 9 9 9 1 9 0 7 13 1 15 9 0 1 9 8 8 2 7 9 9 0 1 9 8 8 2 7 9 0 1 9 9 8 8 2 7 9 1 9 7 9 9 7 9 1 9 0 1 9 2 7 13 9 1 9 9 9 8 2
88 13 8 8 1 2 9 0 15 13 1 9 7 9 15 8 8 9 2 2 7 13 7 15 2 9 0 15 13 1 15 9 1 9 9 1 9 2 7 15 9 0 15 13 1 15 9 9 0 0 1 9 9 1 9 9 9 7 9 9 15 2 1 1 7 13 1 8 0 9 0 1 0 9 2 7 1 0 13 8 14 13 9 0 1 15 8 2 2
85 7 13 7 9 9 13 1 8 9 1 15 2 8 8 13 15 8 1 9 8 0 7 0 7 9 9 1 9 2 7 13 8 9 7 9 1 10 9 2 7 14 13 1 15 9 15 13 7 1 15 9 9 1 8 1 8 0 2 1 7 3 9 7 8 13 1 9 0 1 9 9 0 1 9 0 7 9 2 7 14 13 10 9 1 2
7 2 9 9 8 8 8 2
16 2 9 9 1 9 0 1 10 13 9 0 0 0 1 9 2
15 2 9 9 8 8 9 0 9 15 8 1 9 1 0 2
5 2 8 9 0 2
7 2 9 1 9 9 2 2
35 7 13 1 2 9 8 8 13 1 9 7 4 8 2 7 8 8 0 1 9 1 9 0 1 10 8 8 1 9 8 8 0 8 8 2
30 7 13 2 2 8 8 1 9 8 8 7 14 8 1 9 9 0 2 8 8 10 9 8 8 8 8 8 8 2 2
31 7 13 2 2 14 8 8 9 9 9 15 9 9 1 10 9 1 10 13 9 1 9 1 9 8 8 8 9 13 2 2
35 7 13 8 2 7 8 13 1 9 9 7 10 9 15 9 1 9 1 9 2 7 13 7 13 8 8 1 9 10 13 8 8 8 2 2
18 7 13 3 9 1 2 9 0 7 9 0 9 1 9 8 0 2 2
293 7 13 7 2 9 15 13 1 15 8 1 9 0 8 8 13 15 9 0 1 9 9 2 7 1 9 8 8 1 9 8 9 7 9 9 9 9 7 9 9 9 1 9 8 0 0 2 8 8 13 8 8 1 9 8 1 9 1 9 9 15 13 1 9 1 10 9 2 8 8 13 9 1 9 9 1 9 9 14 13 1 8 9 2 7 3 9 9 13 7 8 9 15 8 1 15 8 8 1 9 9 7 9 7 9 1 1 9 9 9 0 8 8 9 9 7 13 9 13 2 7 9 9 13 13 7 9 8 8 0 8 8 13 8 8 9 1 9 2 7 9 0 1 9 9 9 9 9 2 13 2 0 7 9 8 0 7 7 1 15 9 1 1 15 13 1 15 1 9 1 9 1 9 15 1 0 7 13 8 8 2 7 10 9 13 1 15 13 8 1 9 9 7 15 13 1 15 2 8 8 13 8 1 9 9 8 2 12 15 13 1 9 8 2 12 15 13 1 9 8 1 15 2 1 3 2 7 1 8 8 1 9 9 1 9 0 2 13 9 9 1 8 13 8 8 1 9 15 13 2 7 15 13 1 8 2 12 13 14 9 1 15 8 2 8 8 8 13 13 8 7 15 0 1 9 9 7 13 1 9 7 13 1 9 8 9 0 8 13 10 9 2 2
398 7 13 2 7 9 15 13 1 15 8 1 9 12 12 7 12 12 12 9 14 13 0 9 0 8 1 8 8 2 7 15 9 9 8 8 0 1 9 0 8 8 8 0 8 8 0 1 9 0 9 8 8 8 0 2 7 3 9 1 9 1 9 1 15 13 8 10 9 1 15 9 15 12 7 12 1 12 1 9 2 1 7 9 13 7 13 1 15 1 9 15 8 8 8 1 9 0 7 0 1 9 15 2 8 8 15 8 8 1 1 9 8 9 2 7 0 9 0 1 9 13 1 9 10 9 1 7 13 13 9 1 9 0 1 15 13 8 13 9 1 15 2 14 9 9 14 13 9 1 9 0 1 9 8 0 1 15 13 1 9 0 15 13 7 13 1 9 8 9 0 2 7 9 15 1 9 8 8 8 8 1 9 7 1 15 8 8 7 4 8 8 8 1 9 15 2 1 9 1 7 9 8 0 13 0 1 9 1 12 1 12 1 15 13 13 1 9 12 7 12 1 12 1 9 0 2 8 8 8 9 9 1 9 15 1 9 7 9 1 9 15 8 8 2 7 13 7 8 0 9 8 8 8 7 13 3 9 8 8 10 9 15 13 8 8 2 7 7 8 8 8 8 8 8 9 0 1 9 14 13 8 8 8 2 8 8 13 1 9 8 8 9 0 2 8 8 8 1 8 8 1 9 1 9 8 8 7 9 15 1 7 8 9 9 7 9 8 8 9 8 8 8 8 8 8 8 1 9 9 1 9 8 8 8 1 15 1 8 9 2 7 3 9 1 9 9 8 8 1 9 0 8 8 13 8 8 3 7 8 8 8 2 8 8 8 8 1 9 9 0 1 9 0 1 9 8 8 8 2 7 8 8 9 1 9 9 9 1 9 7 4 1 9 7 1 9 2 2
79 7 9 1 9 13 8 2 2 0 7 9 9 0 13 1 9 9 14 7 15 14 13 1 15 9 1 9 1 10 13 15 1 9 0 0 3 2 7 1 9 8 8 8 9 0 7 14 8 9 1 8 8 2 8 8 8 8 9 1 9 8 8 1 15 13 15 8 8 3 8 8 15 9 1 9 8 8 2 2
9 8 14 0 7 14 0 7 14 0
72 9 12 13 9 9 9 0 2 0 1 0 9 0 2 7 13 9 0 1 9 8 8 8 8 2 1 9 0 8 2 7 13 1 9 9 9 9 9 8 8 9 2 7 14 13 1 8 8 0 8 8 7 14 1 8 8 7 14 1 8 8 2 7 0 8 2 7 14 8 1 15 2
19 13 1 9 9 8 12 1 9 2 12 2 9 9 0 2 2 2 2 2
13 8 2 2 10 9 13 1 9 1 9 9 2 2
55 8 2 2 8 8 8 8 8 8 8 2 2 8 2 2 8 8 3 2 2 8 8 2 2 14 9 0 8 8 13 0 2 2 2 2 2 9 9 12 15 2 8 7 8 8 8 8 8 8 8 7 8 8 2 2
145 13 8 9 8 8 2 7 13 15 9 9 9 0 2 1 9 9 1 9 8 8 7 9 2 7 13 8 1 7 8 1 15 9 2 9 0 2 9 9 2 9 0 2 2 2 7 15 1 9 9 2 7 7 15 9 0 14 14 13 1 9 7 9 8 8 8 8 2 7 7 15 9 0 14 13 9 1 9 9 0 2 7 14 14 13 15 15 9 1 9 8 8 7 13 9 0 8 8 7 1 9 9 1 9 0 9 2 7 13 9 7 15 13 1 9 7 8 8 1 9 8 8 13 9 2 7 13 8 1 8 8 2 7 13 9 8 8 9 7 9 1 9 15 0 2
33 13 9 9 8 1 0 1 15 2 8 8 1 15 8 7 15 13 2 14 13 1 9 0 2 7 15 13 1 9 1 8 9 2
26 7 15 13 8 1 15 14 8 2 7 13 9 9 2 2 9 13 8 8 8 2 2 9 8 2 2
71 7 13 8 7 13 9 9 8 1 9 8 9 9 0 2 12 9 8 0 2 7 13 8 8 1 0 9 0 2 7 13 1 9 15 1 9 7 13 9 2 7 9 9 13 2 13 7 13 9 1 9 9 9 2 14 7 13 15 1 9 15 2 7 13 9 8 2 8 2 9 9
14 2 8 8 8 2 8 8 14 8 8 8 7 8 2
20 8 8 2 2 8 1 9 2 2 9 8 2 8 1 9 0 8 8 8 2
4 2 2 2 2
26 9 9 1 9 0 1 9 9 0 0 1 0 8 8 2 9 0 2 9 8 8 2 1 9 9 2
30 7 15 13 0 8 0 1 8 9 9 8 1 9 15 0 9 2 12 8 8 1 9 9 9 9 9 8 8 2 2
2 2 2
11 2 9 0 2 7 9 0 1 9 0 8
62 13 1 9 9 0 1 9 0 9 1 2 9 0 8 8 8 2 2 13 1 9 10 9 1 9 9 2 9 7 15 13 9 0 1 9 0 2 7 14 13 1 15 9 9 8 7 9 9 8 8 2 9 9 0 1 9 9 1 9 0 2 2
90 1 9 0 1 9 8 13 15 8 8 2 13 8 1 2 9 0 2 9 8 0 2 7 13 2 2 9 0 13 1 9 15 13 9 7 9 8 8 8 0 1 9 15 1 9 0 8 8 2 7 3 9 8 1 9 9 15 2 7 15 1 8 9 1 12 7 12 12 1 9 0 2 7 7 13 10 9 0 7 15 13 0 1 12 8 0 1 15 2 2
16 14 1 9 0 1 9 0 7 13 8 8 0 1 9 0 2
17 12 2 2 9 9 0 0 2 8 8 8 8 1 15 1 15 2
11 12 2 13 8 1 0 8 8 9 8 2
11 12 2 8 14 13 13 1 15 8 8 2
40 12 2 8 8 9 9 0 1 9 1 8 9 9 10 9 9 12 8 2 8 2 7 9 9 13 7 8 8 8 0 1 9 0 1 8 8 1 9 2 12
17 12 2 14 9 1 9 9 12 13 9 1 9 0 1 9 2 2
153 7 13 8 2 2 14 10 9 13 1 9 9 2 7 13 8 8 8 9 2 8 8 8 8 1 9 0 7 1 0 8 8 2 7 13 10 9 9 0 1 9 0 12 7 0 12 2 14 7 9 0 2 8 8 1 10 9 15 13 1 9 0 12 1 8 2 7 15 13 15 8 8 8 13 9 12 8 2 8 9 1 9 0 1 9 8 8 9 9 9 12 9 0 1 15 15 13 9 0 8 8 7 15 14 13 1 9 0 1 9 7 9 15 1 9 2 7 13 10 9 1 9 8 15 13 9 15 1 8 8 2 7 13 1 15 1 12 9 1 9 9 2 7 1 9 0 14 13 1 9 0 8 2
27 7 13 8 2 2 14 9 9 1 9 0 15 9 15 13 1 15 8 2 7 13 8 8 1 9 0 2
13 12 2 2 13 1 9 7 13 9 0 9 0 2
18 12 2 0 15 14 13 8 8 2 8 2 13 9 9 8 8 8 2
14 12 2 9 8 8 8 1 8 8 9 8 8 8 2
25 12 2 9 0 1 9 1 9 12 2 12 14 13 9 15 1 7 15 8 0 8 8 9 0 2
30 12 2 9 0 14 8 8 9 0 1 9 9 9 2 1 9 7 13 1 8 9 7 9 1 7 13 1 9 2 2
103 7 13 8 1 2 9 9 0 1 9 0 2 2 7 13 7 9 13 9 1 15 2 1 9 7 14 8 9 0 1 9 0 2 1 9 7 10 9 0 0 9 1 9 9 0 15 8 8 8 0 1 9 9 15 13 7 3 8 0 0 13 1 15 8 8 0 3 1 9 9 15 0 2 1 1 7 13 0 1 10 9 2 8 8 8 7 9 0 1 15 13 7 13 9 15 13 7 13 1 9 0 2 2
60 7 13 2 7 9 0 2 13 1 9 0 1 9 2 7 13 1 9 0 1 9 8 8 9 8 0 1 15 2 8 9 1 9 15 0 2 8 8 8 9 15 8 9 2 7 9 0 1 8 9 0 8 8 9 1 9 9 0 2 2
30 7 13 1 7 2 9 0 14 13 9 9 15 0 0 7 0 2 7 1 9 9 9 7 13 1 9 9 0 2 2
8 1 9 15 2 9 9 9 0
36 7 8 7 8 9 1 8 8 2 1 9 9 0 2 14 14 8 7 8 8 8 8 2 7 7 8 8 2 1 8 0 1 10 9 0 2
44 9 8 8 8 13 9 9 2 1 9 8 1 15 2 9 0 13 7 9 15 2 8 8 8 9 0 15 8 1 15 2 7 15 13 8 8 1 8 8 9 8 8 8 2
76 13 9 0 8 9 7 9 7 9 2 7 0 1 0 9 9 0 8 2 1 9 9 2 0 8 8 8 8 2 0 8 8 8 8 2 7 10 9 14 13 2 9 8 2 8 1 15 9 1 9 8 8 8 8 2 1 14 8 7 14 8 2 8 8 8 1 9 10 2 7 9 9 0 8 9 2
52 7 13 0 2 1 9 15 8 2 1 7 13 15 2 1 9 0 0 2 9 9 15 13 1 9 2 7 9 15 13 15 9 0 1 9 15 0 0 1 10 9 0 0 7 0 2 2 2 7 15 13 2
59 1 9 2 13 9 9 0 2 1 9 0 0 2 13 7 1 9 7 9 1 12 0 2 15 1 0 1 9 2 1 7 13 0 0 9 15 2 7 1 9 15 13 9 15 2 7 1 9 7 9 15 13 1 9 7 14 13 9 2
51 7 1 9 0 1 9 0 1 9 9 0 7 0 7 0 2 13 9 9 10 2 7 13 7 9 9 13 2 1 10 9 2 13 1 15 9 7 0 7 0 2 0 7 0 2 9 13 7 9 0 2
132 14 9 1 7 3 15 13 1 10 9 1 9 2 7 9 15 13 1 9 9 13 9 2 7 14 15 13 8 8 1 0 1 9 7 9 0 15 13 15 1 9 7 0 7 0 2 8 8 1 15 1 7 9 9 2 7 13 7 13 1 9 15 2 1 10 9 0 2 8 7 8 2 7 14 13 9 1 15 2 7 14 15 1 8 1 2 9 9 2 2 10 2 7 2 13 9 15 15 14 13 1 15 9 15 2 2 9 7 15 14 13 2 1 0 9 1 9 0 8 2 7 9 13 2 1 9 2 15 8 8 9 2
114 8 8 9 7 8 8 8 14 13 0 2 8 8 7 13 9 8 8 9 15 2 7 13 1 9 15 2 1 10 9 0 2 14 13 7 1 15 8 8 0 9 0 2 1 15 8 8 0 2 7 1 15 8 13 15 7 15 13 1 15 2 1 9 1 7 15 13 1 15 8 2 1 8 0 2 13 7 13 9 0 1 15 13 2 1 9 0 2 1 7 13 9 9 2 7 9 9 2 8 8 8 2 7 8 2 1 9 7 8 2 13 8 8 2
62 7 7 13 9 14 13 1 9 15 2 1 7 8 8 8 2 8 8 2 1 9 2 7 7 9 14 13 1 2 7 14 9 2 9 2 1 9 1 9 9 13 7 13 1 15 0 0 7 0 7 13 15 2 1 10 9 0 2 1 9 9 2
51 7 13 13 9 1 2 9 8 8 2 8 2 7 13 1 0 1 9 2 7 13 1 9 15 9 9 1 12 0 2 1 9 0 7 9 2 8 8 14 8 1 9 1 9 9 7 14 1 9 8 2
10 8 8 13 9 7 3 1 15 8 8
18 9 9 12 2 12 2 12 13 8 8 8 9 15 1 9 9 0 2
22 7 13 14 13 15 1 9 0 1 9 2 9 9 0 2 9 9 9 1 9 2 12
143 14 13 1 8 9 15 1 9 2 9 15 13 15 1 9 2 7 13 8 0 8 0 2 8 2 1 9 1 9 2 0 9 9 0 8 8 9 9 1 9 0 7 13 14 13 0 1 9 8 2 8 2 7 13 9 2 12 9 9 15 13 1 8 0 1 9 8 8 1 8 8 8 2 7 13 8 0 9 8 7 8 2 8 8 8 8 8 1 8 9 2 7 9 15 0 2 8 9 8 8 8 8 1 9 2 8 8 1 15 1 9 9 14 9 2 0 8 8 8 9 0 8 8 2 8 8 8 2 8 8 8 8 0 9 0 9 7 9 2 7 1 15 2
113 13 2 8 2 8 8 2 7 13 13 1 9 8 8 7 13 15 2 9 0 8 8 8 1 9 7 9 8 8 2 2 9 9 9 1 9 9 15 2 2 9 8 8 13 15 7 13 15 1 9 8 8 2 2 9 9 0 8 8 1 9 7 9 1 7 13 9 2 2 7 14 13 8 8 8 8 8 2 0 0 1 9 0 2 7 15 14 13 7 13 1 9 9 0 2 8 13 2 8 2 0 1 0 9 7 9 1 9 7 9 7 9 2
146 9 9 1 9 9 0 2 13 9 15 13 8 0 9 9 1 8 2 7 13 9 0 1 9 0 13 8 1 9 0 8 2 7 13 8 13 0 8 8 8 8 15 13 9 9 9 9 7 13 14 13 1 0 1 9 15 7 13 8 8 0 1 9 15 8 8 8 8 8 8 8 2 13 15 9 2 2 2 7 13 13 3 15 13 8 8 1 9 15 7 13 1 8 8 7 13 9 15 1 9 9 0 2 7 14 13 1 9 0 8 2 8 8 8 8 8 2 15 13 2 7 1 9 0 13 8 8 8 9 0 1 8 0 8 8 15 9 1 8 9 1 9 9 0 8 2
69 7 0 15 8 9 15 1 10 9 7 9 0 8 8 8 15 13 15 8 8 1 9 9 9 2 9 12 7 14 13 0 1 9 0 8 2 13 13 1 9 15 9 0 1 9 2 15 9 8 8 8 8 0 8 8 8 13 0 8 8 1 8 1 9 1 9 9 0 2
7 13 15 7 13 13 15 12
193 1 9 1 9 8 8 2 0 0 9 2 7 14 15 13 1 15 9 2 2 8 1 9 1 8 1 9 15 1 9 2 13 8 2 12 2 9 0 13 1 15 2 2 13 15 7 13 13 9 1 9 2 9 13 7 13 1 8 8 8 2 2 2 8 9 9 1 9 1 9 2 1 8 8 2 1 8 8 2 1 8 8 8 8 13 1 15 8 2 1 8 1 9 9 7 8 8 8 8 8 8 1 9 15 2 2 2 2 8 8 2 14 8 2 7 8 1 9 2 1 8 8 2 7 14 8 9 3 0 1 8 8 2 7 14 13 9 1 8 8 3 7 13 8 9 8 8 1 9 8 8 2 8 8 14 8 2 8 8 8 0 2 8 8 8 9 7 13 9 8 8 2 2 8 12 2 12 2 1 8 2 8 8 8 8 2 8 8 2 8 12 2 2
152 7 9 9 8 8 1 8 2 12 2 1 9 9 1 9 2 13 15 9 1 9 2 9 9 2 0 2 2 15 9 15 1 9 9 1 9 0 2 14 13 9 0 7 13 1 9 2 2 7 13 8 2 2 14 2 9 0 13 0 7 13 8 8 1 9 2 8 9 8 2 7 8 1 15 12 9 2 7 13 9 15 0 7 14 13 1 15 13 1 15 1 15 1 8 0 7 0 8 2 7 7 13 1 15 9 0 1 9 8 8 1 9 9 9 2 7 7 13 1 15 9 8 1 15 7 13 15 8 8 13 15 8 2 2 1 2 8 2 2 9 2 8 2 2 9 12 2 12 2 12 2 2
131 15 15 13 0 15 1 9 0 13 1 10 9 1 9 2 7 15 15 13 1 9 2 8 13 13 2 8 2 9 12 7 13 8 9 8 8 2 8 8 13 1 9 9 2 7 1 9 0 1 9 15 9 12 2 2 7 1 9 9 1 15 9 9 1 9 2 8 14 8 9 1 9 8 8 8 2 8 8 13 0 1 2 9 9 2 9 8 8 2 2 7 15 15 13 1 9 0 2 7 2 13 15 2 9 7 9 8 8 7 9 7 9 7 9 7 9 8 8 1 9 14 8 8 9 7 1 9 9 14 8 2
12 7 15 15 13 1 15 1 9 15 13 15 2
129 1 8 8 1 9 0 2 12 9 1 2 9 9 2 8 8 0 8 8 9 7 9 2 8 9 15 8 9 0 8 8 8 2 8 8 2 2 1 15 14 13 1 8 8 1 10 9 8 8 8 8 1 8 8 7 8 7 0 7 0 7 8 2 2 8 8 9 9 8 8 9 15 2 2 7 9 1 8 8 13 1 9 2 7 1 9 8 8 8 8 2 2 1 15 13 8 8 1 9 13 8 8 1 9 2 1 0 8 8 8 8 8 7 8 8 14 13 1 15 13 8 8 1 8 8 1 9 0 2
58 7 7 9 9 8 2 8 8 8 9 15 2 9 2 1 9 15 8 8 8 2 14 13 13 1 8 9 0 15 13 15 8 2 7 15 1 9 2 1 9 15 1 15 14 2 8 2 8 8 2 14 15 13 15 15 2 2 2
46 8 8 1 9 2 1 9 9 0 0 2 7 8 13 9 8 2 7 13 8 8 8 8 8 8 8 8 2 7 13 1 15 9 2 7 7 7 15 15 2 14 13 8 8 9 2
44 8 8 2 13 8 8 8 2 7 13 8 8 8 8 8 0 1 9 2 8 0 2 2 8 8 8 1 15 8 2 8 8 7 13 1 8 15 13 13 15 1 9 9 2
7 2 9 8 2 1 9 0
62 1 9 9 0 1 9 8 8 8 8 9 0 15 13 1 0 1 9 0 0 8 8 8 2 8 7 9 2 2 13 9 0 1 9 8 2 8 2 1 9 1 9 0 8 8 7 9 9 0 0 2 9 8 2 1 9 8 9 1 8 8 2
63 7 13 9 9 3 1 9 9 9 9 0 9 8 8 8 8 9 9 0 9 8 8 8 8 9 9 9 8 8 7 9 9 0 1 9 8 1 9 9 8 9 8 8 9 0 8 8 8 7 9 0 1 9 0 7 9 7 9 8 0 7 0 2
17 7 13 9 8 8 9 1 9 0 1 9 7 1 9 1 0 2
30 2 1 9 2 12 12 9 2 12 12 9 9 2 12 12 12 9 9 2 12 12 1 12 9 7 12 1 12 9 2
35 1 9 2 9 8 12 0 2 12 8 9 2 12 12 9 7 12 9 2 9 0 12 1 12 2 9 12 1 12 7 9 12 1 12 2
81 7 13 8 9 0 1 9 9 9 8 2 7 13 8 9 9 0 1 9 9 0 8 8 9 0 2 7 13 1 9 0 13 1 9 10 9 2 1 15 9 9 1 9 9 7 9 9 9 2 9 9 0 1 9 2 8 9 1 9 8 1 9 1 9 9 0 0 8 8 9 9 0 1 9 8 7 9 9 15 0 2
35 7 13 9 8 9 9 9 7 13 8 8 9 8 8 8 8 2 7 1 9 1 9 9 0 8 8 7 9 0 8 8 8 8 8 2
127 7 13 9 1 9 15 13 1 8 9 13 1 9 0 2 2 9 0 2 8 8 0 2 9 9 8 2 8 7 9 7 9 9 1 0 2 7 9 1 9 9 0 13 1 9 9 9 0 1 9 9 0 2 7 9 9 0 2 8 2 8 7 9 9 0 1 9 2 7 13 9 0 2 9 9 9 9 2 9 8 0 2 9 8 0 2 9 9 2 9 9 9 1 9 2 8 9 2 9 9 0 2 8 2 9 9 0 2 9 8 2 8 1 9 2 8 0 2 9 0 0 8 2 9 0 0 2
6 9 9 9 8 8 0
48 9 9 8 9 8 2 8 2 2 8 2 2 1 9 8 8 0 8 8 13 9 1 9 13 1 15 1 0 0 7 15 8 8 8 1 9 15 9 0 2 0 13 1 8 9 1 9 2
77 7 13 9 8 8 1 9 1 9 9 7 1 9 9 12 9 2 7 13 1 9 9 9 9 8 8 1 8 9 8 8 8 8 8 8 2 7 13 1 9 0 1 9 9 0 15 13 9 1 15 7 14 13 9 1 9 15 9 9 0 2 7 14 13 9 9 0 8 11 2 9 9 9 1 9 9 2
81 1 9 0 2 13 8 1 8 9 15 13 1 9 8 8 9 8 0 2 9 15 13 9 0 1 9 7 12 9 0 1 9 8 2 15 9 9 0 8 8 8 8 8 8 8 8 8 8 8 8 0 2 7 13 10 9 1 9 9 0 0 1 0 9 8 9 8 8 8 2 8 8 8 8 9 8 1 9 12 9 2
97 1 9 0 2 13 9 9 8 0 0 8 8 8 1 9 9 8 8 1 9 8 8 1 9 1 12 9 0 2 7 13 9 9 12 9 9 1 9 9 2 13 15 9 9 9 8 8 9 12 1 9 2 8 8 12 9 9 13 8 8 2 8 8 12 8 8 12 9 0 9 8 8 8 1 2 9 8 0 8 8 9 2 2 9 12 9 9 12 9 0 8 8 8 8 8 8 2
7 8 13 9 15 1 9 8
38 13 9 0 1 9 0 9 9 12 2 12 0 7 9 9 0 1 9 13 1 9 9 15 1 9 0 1 9 0 13 1 9 9 1 9 1 9 2
36 7 13 9 0 7 9 0 13 1 9 9 7 9 9 9 0 9 1 9 0 1 9 1 8 7 8 1 9 9 9 9 9 1 9 9 2
54 7 13 9 7 15 13 9 10 9 1 9 1 9 7 9 7 13 1 9 1 9 9 0 1 9 0 1 9 1 9 0 1 9 9 9 0 7 0 15 13 1 9 1 9 1 9 1 9 9 0 1 9 0 2
64 7 13 9 1 9 1 9 9 9 9 0 1 9 9 7 9 0 13 1 9 0 9 12 1 9 7 9 9 9 9 0 0 1 9 0 1 9 8 7 15 13 7 10 9 15 13 9 15 13 1 9 8 0 0 1 9 8 8 7 14 13 9 8 2
75 7 13 1 7 9 0 13 1 1 9 10 9 1 9 9 9 0 0 9 15 1 9 0 1 9 1 8 7 9 7 8 7 15 13 9 8 9 13 1 15 9 15 1 9 1 9 9 0 1 9 9 1 9 7 9 10 9 1 9 0 7 15 13 15 10 9 1 9 9 0 9 1 10 9 2
13 8 13 1 9 0 9 1 9 7 9 1 9 0
30 13 9 1 8 9 12 2 12 0 7 9 9 1 9 7 9 7 9 1 9 13 9 15 1 9 0 1 9 0 2
41 7 13 8 8 8 2 9 0 1 9 9 7 9 2 7 9 13 1 9 1 0 9 1 9 0 1 9 1 9 0 7 0 2 9 1 9 7 9 0 0 2
43 7 14 13 9 9 1 9 9 1 9 12 2 7 13 9 12 2 12 1 9 9 15 13 9 15 1 7 15 14 13 9 1 9 9 1 15 7 14 13 1 12 9 2
23 7 9 8 8 8 7 1 0 9 1 9 9 1 9 9 12 1 9 14 13 1 15 2
25 7 13 8 1 7 13 9 0 1 9 9 0 1 7 13 9 15 1 9 0 1 9 9 0 2
22 7 13 9 9 1 8 1 8 0 1 9 8 0 2 7 13 12 9 0 1 9 2
25 7 13 8 8 1 7 12 9 0 7 0 13 1 9 1 9 15 13 7 9 15 9 12 9 2
22 7 13 2 2 3 9 0 1 9 1 10 9 7 9 7 7 14 13 1 15 9 2
29 7 13 9 0 1 9 9 7 9 7 9 9 1 9 13 1 9 8 1 9 1 9 9 15 1 8 7 8 2
56 7 13 8 8 9 0 1 9 1 2 9 0 2 2 7 9 15 14 13 15 8 1 9 9 14 13 1 9 8 1 8 7 7 9 1 9 2 0 2 13 9 15 13 1 9 2 14 7 15 14 13 9 9 10 9 2
41 7 13 8 15 13 9 9 1 9 9 9 9 1 9 15 13 9 15 1 9 9 9 0 15 1 12 12 9 7 12 12 9 2 12 1 12 12 9 0 2 2
16 9 0 0 2 8 8 14 13 9 9 15 7 9 9 9 0
19 13 9 0 0 9 7 8 9 9 8 8 14 13 9 15 1 9 9 2
28 7 13 1 7 9 13 9 9 0 13 0 0 0 1 7 9 0 0 0 13 1 9 0 0 1 12 9 2
64 7 1 9 0 1 9 9 8 8 0 1 9 15 13 9 0 9 7 14 8 1 9 9 1 9 9 9 1 9 1 9 15 7 13 1 7 9 8 1 9 0 7 14 13 8 1 9 15 2 7 13 1 7 9 0 14 13 1 9 9 9 1 9 2
76 7 13 9 9 15 7 9 9 0 13 1 9 0 0 7 1 15 2 7 13 1 7 9 1 9 9 13 1 0 0 7 7 9 0 13 1 9 9 12 15 13 1 9 9 0 2 7 13 1 7 9 9 13 9 9 7 0 15 7 9 9 7 9 0 9 1 9 9 7 9 9 0 1 9 0 2
24 7 13 1 7 9 9 0 7 0 0 1 9 9 1 15 2 7 14 13 1 9 9 0 2
21 7 13 1 9 9 9 1 0 9 0 1 9 9 15 1 9 1 9 9 0 2
5 9 9 9 12 9
16 13 9 0 1 9 9 9 1 9 9 7 9 9 0 2 2
28 13 9 0 1 9 0 7 9 9 9 1 9 9 12 13 12 12 9 1 9 9 9 9 9 7 9 9 2
38 13 9 7 9 12 14 13 9 1 9 9 9 1 9 9 13 12 12 9 1 9 12 1 15 13 9 9 15 13 1 15 9 7 9 7 9 0 2
80 13 1 9 7 9 0 1 9 12 13 1 9 12 12 7 12 9 1 12 12 7 12 9 1 9 12 13 0 15 1 9 9 7 9 7 9 7 0 7 13 1 15 9 12 9 1 9 1 9 0 7 7 9 0 13 12 12 7 12 9 7 13 1 9 1 9 9 7 9 1 15 7 9 1 9 7 9 9 0 2
51 7 13 9 0 15 13 1 9 1 9 12 12 7 12 9 0 15 13 12 9 9 9 0 7 12 9 9 7 12 9 9 7 9 0 0 7 12 12 7 12 9 7 12 9 9 0 7 12 9 0 2
56 13 9 7 3 9 0 1 9 9 7 9 7 15 14 13 1 9 9 0 7 7 10 9 1 15 9 13 9 15 1 9 1 15 1 9 9 15 7 9 15 1 9 9 15 7 7 1 10 9 13 9 9 0 1 9 2
6 9 0 0 1 9 0
70 13 9 0 0 1 9 0 0 13 9 15 1 9 1 9 0 1 15 2 7 13 9 7 7 9 9 0 14 13 9 15 1 9 9 1 7 13 9 0 8 8 1 9 9 1 9 9 9 9 1 9 12 9 0 1 9 1 9 7 13 9 9 0 1 9 1 12 12 9 2
65 7 13 9 9 9 9 1 9 15 10 9 1 12 5 1 9 0 1 9 15 13 1 1 12 12 9 7 13 9 9 7 9 9 0 14 13 1 9 15 13 1 15 9 0 1 15 7 13 15 1 15 9 9 9 9 0 1 15 7 15 13 12 12 9 2
171 7 13 9 0 1 9 1 9 7 8 1 9 7 9 1 9 0 1 9 9 9 1 9 9 7 14 13 9 9 15 1 9 9 12 7 13 9 8 12 12 7 12 12 9 7 9 12 12 7 12 12 9 7 13 1 12 5 1 9 9 7 1 9 1 9 9 9 1 9 15 0 1 9 1 10 9 14 7 15 13 9 0 1 9 9 9 0 9 9 9 1 9 9 9 0 9 1 9 0 7 0 1 9 0 0 1 9 9 0 14 7 9 13 7 9 9 1 9 0 14 13 1 9 9 0 1 9 9 9 9 0 0 2 7 13 9 0 9 15 13 1 0 7 13 1 9 9 0 1 9 9 0 1 9 9 0 7 15 13 1 9 15 0 1 12 9 1 0 9 0 2
12 9 0 13 9 0 1 12 1 2 9 0 2
61 13 9 0 0 7 9 0 14 13 9 0 9 1 12 1 9 7 9 1 2 9 0 2 1 9 9 9 9 12 2 7 14 13 9 7 13 1 0 1 15 9 1 9 9 9 9 13 1 9 9 9 8 8 7 13 1 12 9 1 9 2
27 7 13 9 13 9 0 9 9 9 8 8 7 12 1 9 2 9 9 2 8 8 8 8 8 8 8 2
74 7 13 9 1 7 9 1 9 1 9 2 9 0 2 13 1 9 1 9 0 1 9 9 2 7 13 9 0 8 8 8 7 15 13 9 7 13 0 9 1 9 0 15 13 1 15 9 1 9 12 7 14 13 1 9 15 14 13 9 15 9 15 15 13 15 8 2 7 7 15 13 9 0 2
21 7 9 13 7 13 9 1 9 9 9 9 1 0 1 9 0 1 9 9 0 2
151 7 1 9 9 9 2 9 0 2 9 0 1 9 0 7 9 13 1 9 0 7 9 15 13 15 9 0 0 1 9 15 0 2 7 1 15 9 9 0 7 0 7 0 9 0 1 9 9 2 7 3 9 1 7 2 9 0 2 14 13 1 9 9 15 1 9 2 7 15 15 13 15 9 9 9 15 7 13 9 15 9 9 7 9 0 1 9 0 2 1 9 9 9 15 13 1 9 7 9 14 13 0 2 7 7 9 9 0 13 7 13 15 9 7 14 13 1 15 9 2 7 13 7 9 2 13 1 0 9 0 9 7 9 2 7 13 1 7 15 2 14 13 9 0 9 0 0 9 15 2 2
70 7 13 8 7 9 1 9 9 8 8 0 1 9 1 9 0 2 9 9 13 1 9 1 0 2 7 13 1 9 9 9 0 7 13 2 2 14 9 0 13 8 8 9 9 0 0 13 1 9 9 15 1 9 0 7 9 15 1 9 7 9 15 13 15 1 9 0 7 0 2
15 9 2 9 2 1 0 15 7 0 15 9 1 9 9 9
146 13 9 1 9 9 1 9 9 9 9 0 1 9 2 9 2 1 9 2 0 2 9 9 9 0 9 1 9 9 7 9 1 9 1 9 7 9 8 7 13 10 9 9 1 2 9 7 9 1 9 1 9 7 9 0 1 9 1 9 0 1 9 7 9 9 9 1 9 15 0 3 1 0 9 1 15 7 1 9 9 7 9 1 9 1 9 9 0 2 7 13 9 10 9 9 9 0 13 2 8 2 8 8 1 12 9 7 7 14 13 3 9 8 8 7 9 1 9 1 9 12 9 7 9 9 9 1 9 7 9 9 7 9 2 2 7 13 9 9 7 9 13 9 9 9 2
92 7 13 9 0 0 9 15 1 9 1 9 7 9 2 8 2 1 9 9 1 9 9 1 10 13 2 7 13 9 0 7 10 9 0 13 1 8 7 9 9 7 13 1 9 0 7 15 13 1 9 1 9 1 8 1 12 8 9 7 13 9 9 15 13 1 9 15 1 9 8 9 1 2 9 0 7 9 1 9 7 9 9 7 9 1 9 7 13 9 0 2 2
9 9 9 0 1 9 12 12 9 0
98 13 9 13 15 9 9 1 9 9 7 9 9 1 9 0 13 1 12 7 12 12 9 0 7 13 10 9 1 9 9 9 0 7 13 9 0 1 9 15 2 7 13 9 9 9 1 9 9 0 2 7 9 9 0 9 1 9 15 2 7 9 9 1 9 9 1 1 9 2 7 9 1 9 9 1 9 1 15 13 1 9 9 9 9 7 15 13 15 1 0 7 9 13 9 0 1 9 2
39 7 13 9 0 1 9 0 7 9 7 9 10 13 15 9 0 1 9 7 9 0 13 1 12 12 9 13 9 9 1 9 1 9 7 9 7 9 0 2
40 7 13 9 9 9 7 9 9 0 13 1 12 12 9 0 14 13 9 9 1 15 1 9 12 9 1 9 9 9 7 9 9 9 0 1 9 9 9 9 2
15 9 0 2 12 5 1 9 13 9 0 7 9 0 13 9
132 13 9 7 9 1 9 9 0 9 15 7 13 1 8 1 9 1 9 0 1 9 9 0 7 9 9 2 7 1 13 1 9 13 7 1 15 9 0 1 9 9 1 9 0 7 9 9 15 7 9 0 15 1 9 15 1 9 15 13 1 15 9 7 9 9 15 13 1 15 9 7 13 7 12 5 1 9 1 9 13 1 9 0 7 7 9 13 1 9 7 13 1 12 5 1 9 15 2 7 9 15 1 7 9 9 0 3 1 9 1 9 7 9 1 7 9 13 7 13 1 9 0 7 13 1 9 9 0 1 9 8 2
69 7 13 1 2 9 2 9 9 0 1 9 0 9 8 8 7 9 9 13 1 9 1 9 0 1 10 9 0 7 0 1 7 9 15 13 15 9 0 0 7 0 7 0 7 9 9 7 9 7 9 9 7 9 7 9 9 13 1 9 9 15 14 13 9 1 9 9 15 2
72 14 8 8 8 7 15 9 9 9 1 9 8 8 7 13 1 9 1 9 15 13 9 9 7 9 15 13 1 9 1 9 9 9 1 9 9 9 9 7 9 9 15 1 9 0 2 7 3 9 1 9 9 9 0 7 9 9 9 14 13 1 9 0 7 15 14 13 1 9 9 0 2
45 7 14 13 9 7 13 1 1 9 1 8 8 7 13 9 8 8 9 9 0 1 9 9 8 9 13 1 15 7 8 0 13 9 1 9 0 1 9 9 0 8 8 8 9 2
52 7 7 13 9 9 9 9 1 10 9 2 7 13 8 8 13 1 7 9 9 9 1 9 0 15 12 9 9 9 14 7 15 8 9 15 15 13 1 7 9 0 7 0 13 9 9 7 1 0 9 0 2
7 9 9 0 8 9 8 8
61 13 9 0 9 12 2 12 0 9 2 9 0 2 8 8 7 9 15 8 8 8 7 12 0 1 9 9 2 1 9 13 15 9 1 9 9 8 8 1 9 15 2 1 9 9 9 0 0 9 12 2 12 0 2 7 0 1 9 9 0 2
40 3 7 9 9 8 1 2 9 0 0 2 13 15 9 15 7 15 9 1 15 8 14 13 1 9 0 13 1 15 7 14 13 1 15 9 1 9 7 9 2
19 7 2 9 0 2 13 9 1 9 7 13 8 7 14 13 13 9 0 2
57 7 13 9 15 3 3 1 9 9 0 15 13 15 1 9 9 9 8 8 3 13 15 9 15 1 9 9 9 2 7 13 1 0 9 1 9 0 7 9 0 1 9 7 9 1 9 1 9 9 9 0 13 9 9 1 9 2
15 7 7 15 14 13 9 9 0 1 0 9 15 1 9 2
33 7 15 13 13 1 9 14 13 15 1 9 8 7 9 15 9 15 7 9 13 7 13 15 2 3 8 14 13 9 0 7 0 2
28 7 14 14 15 13 9 15 13 9 1 9 9 2 9 0 2 1 1 9 15 13 9 9 0 7 9 9 2
25 7 7 9 0 13 0 9 1 9 8 8 12 1 9 10 9 15 13 9 8 1 9 9 0 2
39 7 0 7 9 15 14 13 9 1 9 1 9 0 0 2 7 2 9 2 2 7 15 9 9 0 9 7 14 9 2 13 15 7 7 13 13 1 15 2
53 7 9 1 9 9 8 8 13 7 9 8 2 9 0 2 2 7 15 13 7 9 0 15 13 1 15 9 2 9 0 2 7 14 13 9 9 2 0 2 7 13 2 2 15 14 13 9 9 1 9 15 2 2
73 7 13 9 7 9 0 14 13 2 9 9 2 1 9 9 2 9 0 15 8 9 8 8 1 15 1 9 1 1 9 2 9 0 2 2 7 9 15 13 1 9 9 7 9 15 2 7 3 0 15 13 1 0 9 13 1 15 9 15 2 9 1 9 15 13 7 13 1 9 9 15 0 2
66 7 13 9 7 9 8 9 0 9 8 8 0 1 9 9 7 9 7 9 13 1 9 0 2 7 9 1 9 15 9 2 1 9 8 9 12 2 13 9 15 1 9 13 9 9 7 9 15 7 13 9 9 9 0 0 7 13 9 9 9 0 1 9 7 9 2
46 9 9 0 13 15 9 9 0 9 0 0 9 8 8 7 13 7 15 13 1 9 2 9 9 7 4 9 2 2 0 1 7 2 9 13 1 9 1 9 7 15 14 13 1 2 2
24 8 7 8 13 7 9 8 2 13 8 8 1 9 0 1 9 15 8 8 13 9 9 2 2
15 7 13 2 2 9 0 14 13 1 9 7 15 9 9 2
15 7 14 13 9 1 9 1 9 7 13 1 9 15 2 2
10 0 1 9 13 1 9 9 0 1 9
30 13 9 0 1 9 1 9 9 0 1 9 1 9 8 2 1 12 12 7 12 12 9 13 1 15 1 9 9 0 2
37 13 9 8 8 9 9 0 1 9 9 9 12 8 1 9 1 9 15 13 9 15 2 7 15 9 0 1 9 1 9 9 1 9 9 9 9 2
35 7 13 8 1 9 9 8 8 9 1 9 1 9 9 0 1 0 9 2 7 15 9 15 13 13 15 8 1 9 1 9 9 1 0 2
5 12 12 9 2 2
5 9 9 0 1 8
41 13 9 0 0 1 8 9 9 9 0 1 9 0 0 1 9 1 9 1 9 0 13 12 12 9 1 12 1 9 9 1 9 12 7 1 9 9 15 12 5 2
38 7 13 9 1 9 15 13 15 1 9 8 9 9 7 9 0 1 9 0 1 9 9 13 9 15 1 12 12 1 12 12 1 9 9 1 9 0 2
22 13 9 7 9 9 9 0 13 1 12 12 1 12 9 0 1 9 9 15 12 5 2
21 13 9 9 9 15 13 1 9 9 1 14 2 8 8 2 2 8 8 8 9 2
12 8 0 0 2 0 0 1 0 1 12 12 9
196 13 9 0 0 15 1 0 7 13 9 0 0 9 12 2 12 0 7 13 9 0 0 9 9 0 1 9 7 9 9 0 0 1 9 1 9 9 1 9 0 0 1 9 13 12 12 9 13 1 9 9 7 9 7 9 7 9 9 7 9 0 2 7 13 9 0 15 13 9 1 9 9 7 9 9 0 7 9 9 0 2 7 13 9 1 9 9 0 2 9 9 9 13 1 9 1 9 9 7 9 8 7 9 9 0 7 9 9 7 9 7 9 9 9 9 9 0 0 1 9 9 0 1 9 9 9 1 9 1 9 0 7 0 7 0 9 1 9 9 7 9 8 0 2 0 1 9 9 7 9 7 9 0 1 9 9 7 9 1 9 1 9 9 9 9 9 2 7 13 9 9 0 1 9 9 0 7 9 8 7 9 7 9 7 9 9 7 9 9 14 3 1 9 9 9 2
71 7 13 9 1 7 10 9 14 13 0 1 9 0 7 7 3 0 1 9 0 1 9 1 9 7 9 9 7 9 0 13 7 9 9 1 9 0 0 1 0 1 9 15 1 9 0 7 7 9 0 7 0 13 1 9 1 9 7 9 9 9 7 9 9 0 9 1 9 9 9 2
73 7 13 9 9 9 0 9 9 9 9 7 9 13 9 9 9 1 9 9 7 9 0 0 1 9 1 9 1 9 0 0 1 10 9 7 15 1 9 1 9 9 1 9 0 1 9 0 15 13 9 0 1 9 0 7 13 9 7 9 0 1 9 7 9 13 15 1 9 0 7 0 0 2
112 7 13 9 9 9 0 9 9 15 13 9 15 1 9 9 0 1 9 12 12 9 2 12 12 9 2 13 9 15 1 9 0 7 0 7 0 7 9 9 9 0 0 7 9 7 9 7 13 9 15 0 12 12 9 2 12 12 9 2 7 0 1 9 12 12 9 2 12 12 9 2 7 13 1 9 1 9 0 1 9 1 9 7 9 7 9 9 0 0 7 13 9 1 9 0 15 13 1 15 9 1 9 0 7 0 7 9 9 8 7 9 2
87 7 13 9 9 9 0 0 8 8 8 7 15 14 13 1 9 9 9 9 0 1 9 9 0 7 0 7 9 15 14 13 9 15 1 9 7 14 13 9 0 9 9 0 1 9 0 1 9 13 1 9 1 9 9 1 9 0 1 9 2 7 13 8 1 9 9 9 0 9 1 9 1 9 0 7 9 9 9 1 9 9 7 9 9 1 9 2
108 7 1 9 15 13 9 9 9 0 0 8 8 7 9 9 0 13 9 9 1 1 12 9 0 1 9 7 9 0 13 0 1 9 0 7 9 7 9 7 9 7 9 9 0 7 0 7 9 7 9 0 7 9 9 7 9 8 7 9 7 9 9 8 9 2 7 14 13 9 0 1 9 15 0 9 9 9 9 0 15 13 7 13 1 1 9 8 8 8 1 9 9 0 1 9 0 9 0 13 1 9 0 7 9 0 1 9 2
36 7 13 9 9 0 8 8 7 9 0 13 9 1 9 0 13 9 0 0 2 0 1 1 9 1 9 7 9 9 0 1 9 7 9 0 2
8 9 13 9 15 1 9 2 2
13 9 1 9 9 2 8 2 1 9 7 9 7 9
71 13 8 13 9 0 1 9 7 9 1 9 9 0 9 0 1 9 15 7 9 15 2 7 9 9 9 9 15 14 13 0 1 9 9 2 15 1 0 15 9 9 0 1 9 1 9 2 8 2 1 9 8 2 8 8 2 8 8 2 7 9 0 1 9 9 7 9 7 9 0 2
75 7 13 9 9 9 0 8 8 8 1 9 1 9 9 0 9 12 9 0 1 9 0 9 1 9 9 0 0 1 9 9 10 9 0 2 7 14 13 9 0 1 9 9 0 9 8 8 8 8 1 9 7 9 9 1 10 9 1 9 1 9 13 1 12 9 2 7 13 1 9 9 0 1 9 2
123 7 13 9 0 1 2 9 0 2 7 9 0 14 13 1 9 1 9 0 1 9 0 2 8 2 1 9 9 9 9 7 9 1 9 9 15 13 1 15 9 1 9 9 0 1 9 15 7 15 13 1 9 2 8 2 1 9 0 7 15 13 1 9 0 0 1 9 8 7 9 2 8 8 1 15 14 13 15 9 9 0 1 9 0 1 9 1 9 9 1 9 0 0 7 15 1 0 15 9 7 9 9 1 9 7 15 13 9 15 7 9 9 9 1 8 9 8 8 8 9 9 0 2
57 7 13 9 7 9 1 9 0 7 9 0 14 13 9 1 9 0 1 9 9 0 1 9 7 9 7 9 9 9 15 2 8 8 13 9 9 15 14 13 8 1 9 1 9 9 1 9 10 9 0 7 13 0 8 1 9 2
15 9 9 0 2 9 0 13 9 9 1 9 0 2 0 0
48 1 9 9 7 9 15 13 15 9 7 9 0 0 0 1 9 0 2 13 9 0 1 9 9 0 9 9 0 9 9 1 9 0 1 9 9 1 9 7 13 1 9 9 9 0 1 15 2
53 13 9 9 7 9 0 13 9 9 1 9 0 0 1 9 1 9 1 9 9 0 1 9 9 0 1 9 1 9 15 2 9 1 7 9 1 9 7 1 0 9 0 13 9 9 0 1 9 9 0 1 9 2
38 7 13 9 9 7 9 9 9 9 1 9 0 13 9 0 2 0 7 9 0 13 9 9 1 9 9 15 13 1 15 7 9 0 15 13 1 15 2
22 7 13 1 9 9 15 1 12 9 1 7 9 0 9 15 1 9 9 1 9 9 2
38 13 8 8 9 9 2 9 12 9 2 7 9 0 13 1 9 9 1 0 1 9 0 15 13 15 1 9 0 1 9 9 7 9 1 9 8 0 2
28 7 13 7 9 8 0 14 13 1 15 9 9 0 13 9 9 1 1 15 9 9 0 9 0 1 9 0 2
53 7 13 9 8 8 9 0 1 9 9 9 0 1 7 15 0 1 9 0 9 1 9 9 0 0 2 0 9 0 1 9 9 2 7 9 9 0 2 7 9 9 9 0 1 9 9 1 9 0 1 9 9 2
53 7 13 9 8 8 9 9 9 0 1 9 9 7 9 9 1 9 0 9 1 9 0 1 12 12 9 3 0 1 9 7 0 1 9 2 0 7 9 1 9 9 1 9 9 0 2 7 13 9 1 9 0 2
50 7 13 8 7 1 1 9 15 13 9 9 1 9 9 9 8 2 0 7 0 9 9 1 9 0 15 9 9 1 9 0 7 15 15 13 1 15 9 9 2 1 9 1 9 9 7 9 7 9 2
48 7 13 1 7 15 1 1 9 9 7 9 14 13 9 8 1 9 9 3 7 7 13 8 1 9 0 9 8 2 7 13 9 1 9 15 1 9 0 15 13 15 9 7 13 1 9 9 2
47 7 13 8 9 1 9 1 9 9 0 7 0 1 9 1 9 0 0 7 9 8 8 9 0 1 0 9 1 9 1 8 8 9 1 9 9 9 7 9 0 0 1 9 2 8 2 2
13 13 9 9 9 0 1 9 7 8 1 12 12 9
66 13 9 0 0 2 0 0 9 15 1 9 0 2 9 2 2 1 9 9 9 0 1 9 9 9 1 9 1 0 9 2 7 14 13 9 15 13 9 9 9 9 0 2 7 14 13 9 1 10 9 2 9 0 1 9 9 9 0 1 9 1 12 12 9 0 2
79 7 13 9 8 8 8 9 9 1 9 0 2 7 9 9 0 1 9 9 2 1 7 9 0 1 9 9 13 9 0 1 9 9 7 9 9 8 8 2 8 8 8 2 7 9 1 9 9 15 13 1 15 9 9 0 2 7 1 9 15 9 0 1 9 9 1 9 9 1 9 9 0 1 9 0 1 1 9 2
12 9 1 9 9 1 9 1 9 14 2 8 2
55 13 9 1 9 9 1 9 9 7 9 1 9 1 9 1 9 1 9 9 0 0 1 9 8 1 9 7 15 13 9 9 1 9 0 1 9 0 1 9 7 13 9 0 1 10 9 1 12 5 1 8 9 0 2 2
52 9 0 1 9 13 0 9 10 9 7 7 9 14 13 9 0 1 10 9 7 13 9 1 9 7 9 0 7 7 9 0 1 9 9 1 9 1 9 1 9 0 1 9 0 2 1 9 9 2 9 0 2
7 9 9 9 0 0 2 2
58 9 15 13 10 9 9 0 7 9 15 13 9 15 0 7 9 13 1 9 9 0 7 13 15 9 9 10 9 7 14 13 7 13 1 10 9 9 1 9 9 9 0 0 1 9 7 8 1 9 0 1 9 9 9 0 1 9 2
28 7 13 9 0 1 9 9 7 10 9 14 13 1 9 1 15 0 9 7 14 13 1 0 9 1 9 9 2
35 2 8 13 7 15 13 1 9 0 7 13 9 0 8 13 1 15 9 1 9 7 9 7 9 9 13 1 15 9 7 14 9 2 2 2
24 15 13 15 9 0 9 9 0 1 9 0 7 13 1 15 9 9 0 7 9 9 0 2 2
10 7 13 2 2 6 13 8 8 2 2
59 7 6 8 13 1 15 9 2 1 9 9 15 7 9 1 9 15 13 9 9 0 0 2 8 2 13 9 9 15 1 9 9 7 9 9 0 1 12 12 9 1 9 12 9 1 9 9 7 13 9 15 1 15 14 13 12 12 9 2
34 7 13 9 7 9 15 13 15 9 1 8 13 9 13 1 12 5 7 9 9 15 13 15 9 9 2 8 2 14 13 1 9 2 2
52 7 13 7 9 15 13 15 9 1 9 14 13 1 9 7 13 9 9 1 9 0 1 9 0 9 9 10 9 15 12 5 1 8 9 0 1 9 8 7 13 9 0 1 9 12 5 1 9 7 15 9 2
37 7 13 9 1 7 9 13 1 9 12 2 9 9 2 7 14 13 9 9 0 1 9 9 0 7 9 13 1 1 9 15 13 7 13 9 9 2
50 1 9 15 13 8 8 9 9 9 9 9 0 7 3 1 9 9 1 9 8 0 1 9 0 13 9 7 9 0 7 13 1 9 1 7 15 13 3 9 1 9 9 15 13 1 9 1 9 2 2
20 0 7 9 9 1 9 9 15 9 9 1 9 1 9 9 0 1 9 0 2
52 7 13 8 8 8 9 9 9 9 7 9 10 9 14 13 1 9 0 7 15 1 9 13 7 13 15 9 9 9 7 9 0 7 7 9 9 0 1 9 1 9 7 15 9 9 0 9 0 7 9 0 2
25 7 13 9 1 8 8 9 9 9 9 8 8 8 9 9 0 1 9 0 7 13 3 9 2 2
28 7 14 13 7 13 3 9 1 9 9 9 0 0 1 9 9 1 9 9 9 0 1 8 7 13 1 9 2
19 7 13 8 7 13 1 15 0 9 1 10 9 15 13 1 15 9 0 2
45 7 13 8 8 9 9 9 9 0 7 3 9 13 1 9 1 9 9 0 7 0 1 9 9 0 1 9 1 9 9 0 0 0 7 13 3 9 1 9 1 10 9 1 9 2
57 7 13 8 7 9 9 13 9 1 9 9 9 1 9 0 9 9 0 7 13 9 9 1 9 9 1 9 0 1 9 9 0 1 9 0 7 13 7 15 1 7 10 9 9 0 1 9 9 7 15 9 0 1 9 9 9 2
106 7 13 9 1 9 9 14 13 0 1 9 9 1 9 9 9 1 9 9 9 0 0 2 8 2 1 9 9 9 7 9 0 9 9 0 15 13 0 1 9 1 9 9 0 15 13 1 9 0 0 1 9 0 1 9 0 0 7 10 9 14 13 9 9 10 9 1 9 12 12 9 2 7 15 15 13 9 0 1 9 1 9 9 9 8 1 9 10 9 1 9 0 1 9 1 9 9 9 7 9 7 9 1 9 0 2
11 9 13 1 9 8 1 9 9 1 9 0
54 13 9 8 8 8 9 9 0 0 7 9 15 14 13 1 9 9 0 1 9 9 0 1 15 1 9 9 0 1 9 9 9 9 0 1 9 1 9 7 9 1 9 7 10 9 13 9 0 1 9 1 9 0 2
32 7 13 9 8 7 9 13 1 15 7 13 9 0 1 9 0 1 9 0 1 9 9 9 7 15 1 1 9 9 0 9 2
57 7 13 9 9 0 0 14 13 9 13 1 15 7 9 14 13 1 9 0 1 9 9 0 1 9 10 9 0 9 1 7 15 13 9 9 9 0 2 1 10 9 0 7 9 9 15 9 0 1 9 9 9 9 1 9 0 2
44 7 13 9 1 7 15 7 13 9 9 1 9 12 9 13 1 9 0 9 9 9 9 1 9 1 9 15 7 9 15 7 13 9 0 9 1 9 9 9 0 1 9 15 2
14 9 0 2 0 2 0 0 1 9 0 9 1 9 0
39 13 9 0 1 9 7 9 0 1 9 0 1 9 15 1 9 0 9 9 1 9 9 7 9 9 1 9 0 0 1 9 1 9 9 0 7 9 15 2
143 7 13 9 8 8 9 9 9 1 7 9 0 13 9 15 1 9 0 12 12 9 2 7 13 9 15 1 12 12 9 2 7 13 1 9 9 12 5 1 9 7 12 5 9 0 7 12 5 0 2 7 14 13 1 9 9 0 0 1 9 8 1 9 12 12 9 0 2 7 14 13 9 0 9 15 1 9 12 5 1 8 7 8 7 8 0 1 9 9 0 1 9 0 7 1 9 12 12 9 9 0 1 9 12 9 8 1 9 0 2 8 8 1 9 1 12 9 1 9 1 9 9 1 9 7 9 2 7 13 9 12 9 9 1 9 2 7 7 15 0 1 9 2
131 7 13 9 9 9 7 15 14 13 9 9 1 9 1 9 9 0 1 9 9 9 0 9 2 0 1 9 0 0 1 9 1 9 12 9 0 1 9 12 12 9 2 7 1 9 12 9 2 7 13 9 12 9 9 1 9 7 13 12 5 1 9 15 1 1 9 2 7 9 0 13 1 9 0 0 1 9 1 9 12 9 0 2 7 13 1 9 9 0 1 9 9 15 2 7 3 9 9 2 7 13 9 15 1 1 9 7 13 12 9 9 1 9 2 7 13 9 15 12 12 9 2 7 13 9 15 1 12 12 9 2
95 7 13 8 2 8 8 7 9 9 14 13 1 9 9 9 7 9 9 9 0 7 9 0 9 1 9 9 1 9 7 9 9 7 9 9 7 9 7 9 9 0 1 9 2 7 3 9 9 8 0 1 9 10 9 2 8 8 1 9 9 15 1 1 9 1 9 12 5 2 7 13 9 10 9 12 12 9 2 7 13 9 15 1 12 12 9 2 7 13 9 1 12 9 9 2
32 7 13 9 9 9 2 14 15 14 13 9 1 9 9 0 1 9 9 1 9 9 1 9 9 9 0 1 1 12 12 9 2
8 12 12 9 9 9 1 12 9
48 13 8 8 9 9 9 7 9 9 7 9 9 9 9 1 9 0 1 12 9 0 13 12 12 7 12 12 9 1 9 12 12 9 0 8 1 9 12 5 1 9 9 0 0 1 9 0 2
53 7 13 8 7 9 9 0 13 12 8 8 9 1 9 12 5 1 9 9 9 0 1 9 0 0 1 7 9 8 8 1 9 9 1 9 13 12 8 8 8 1 9 12 5 1 9 9 0 1 9 1 9 2
34 13 7 9 0 1 9 0 10 1 9 9 7 9 9 0 13 12 12 9 0 8 1 9 12 5 1 9 9 0 0 1 9 0 2
9 9 13 9 0 0 1 9 9 9
58 13 9 9 2 9 2 0 7 9 0 13 1 0 9 9 1 9 9 9 1 9 9 9 9 0 2 7 1 0 7 13 9 9 9 9 0 1 9 9 0 1 12 12 9 7 13 9 9 0 1 9 9 9 9 1 10 9 2
50 7 13 0 9 0 1 9 2 8 2 0 7 9 9 9 9 15 13 9 15 1 9 0 13 1 12 12 9 2 7 7 9 9 9 0 9 15 1 9 1 9 9 12 14 13 1 12 12 9 2
15 1 9 9 2 9 9 9 7 9 9 9 7 9 7 0
41 13 9 9 9 8 8 9 9 9 12 2 12 0 1 9 9 0 9 1 9 9 15 1 9 0 7 9 1 9 0 9 15 1 9 0 1 9 9 9 0 2
100 7 1 15 13 9 15 13 2 9 9 2 1 9 1 15 9 1 9 9 1 9 0 1 0 9 0 7 0 2 7 14 13 1 9 1 9 0 0 2 13 1 9 15 9 9 9 7 13 1 12 5 9 1 9 12 5 9 0 2 7 13 15 9 9 0 1 9 9 1 1 12 1 12 5 9 0 7 9 9 0 1 9 9 1 1 12 5 7 15 1 9 9 9 9 7 9 9 9 0 2
50 7 13 9 9 7 9 9 15 13 0 1 15 7 13 1 12 5 13 10 9 1 12 5 13 10 9 1 12 5 7 13 9 15 1 9 9 9 1 9 0 1 9 9 10 1 7 1 9 9 2
13 7 13 9 9 9 9 0 7 13 1 12 5 2
38 7 13 9 9 1 9 0 0 1 9 0 12 2 12 13 12 12 9 1 9 15 13 15 0 7 13 9 0 9 0 1 12 12 9 1 9 0 2
48 7 14 13 9 9 9 0 9 9 0 1 9 0 2 12 5 13 15 9 9 7 9 12 5 7 9 9 12 5 7 13 9 9 9 7 9 0 7 14 13 12 5 7 12 5 1 9 2
60 7 1 7 9 14 13 9 0 1 9 9 1 9 0 13 12 12 9 2 7 13 1 12 12 9 2 14 7 15 13 1 9 9 15 9 1 9 9 0 7 9 15 1 9 0 7 13 1 12 5 9 1 12 5 1 9 12 2 12 2
43 14 9 9 7 15 13 1 9 0 1 9 12 5 7 14 13 1 12 5 1 9 0 0 7 13 1 12 5 7 15 14 13 9 0 7 0 1 0 8 8 9 9 2
59 7 13 9 1 9 9 9 0 1 9 12 5 7 13 1 12 12 9 1 9 13 9 0 1 9 9 13 12 12 9 7 13 1 12 12 9 7 13 9 15 1 9 0 1 12 5 9 1 12 5 9 0 9 1 9 9 9 2 2
32 14 9 0 7 14 13 9 7 15 14 13 1 9 12 12 9 1 9 13 0 1 9 9 1 15 7 13 1 12 12 9 2
23 7 13 9 7 9 15 1 9 0 14 13 1 9 0 12 2 12 1 9 12 12 9 2
44 7 7 13 9 1 9 9 9 0 7 0 1 12 12 9 1 9 9 15 12 12 9 1 9 0 7 14 13 9 9 10 9 9 12 12 9 1 9 0 1 9 0 0 2
20 7 13 9 0 9 9 15 12 12 9 7 13 1 12 12 7 12 12 9 2
18 7 1 9 0 13 9 9 1 9 9 9 15 12 5 1 9 0 2
61 7 13 9 1 9 15 7 15 13 1 9 0 12 2 12 9 12 12 9 1 9 0 1 15 7 13 9 10 13 15 1 9 12 1 12 12 9 1 9 13 7 15 13 9 9 9 0 0 1 1 9 9 9 9 0 1 0 9 9 0 2
52 14 1 9 7 14 13 9 7 15 13 12 12 9 2 12 5 1 9 9 2 13 9 9 0 1 9 12 5 1 15 2 1 9 13 9 9 0 12 12 2 12 5 1 9 9 2 7 9 0 12 5 2
7 12 9 9 13 1 9 0
97 13 12 9 9 0 1 9 1 9 9 0 1 9 1 7 13 9 9 0 9 9 8 8 8 9 9 0 0 0 1 9 9 12 9 9 13 9 15 9 1 9 9 9 0 0 9 0 1 9 0 2 1 9 1 9 12 9 0 1 9 9 9 15 9 1 9 9 8 8 13 9 9 0 13 0 9 0 1 9 9 9 0 1 15 13 9 7 9 9 9 1 12 1 12 12 9 2
53 7 1 15 13 0 1 9 9 9 0 1 9 9 1 9 9 0 0 1 9 7 13 12 9 9 15 0 7 13 9 15 1 9 0 7 13 12 9 0 1 9 1 9 1 9 9 1 9 9 15 9 0 2
62 7 13 9 9 0 0 9 9 9 8 8 9 8 8 9 9 0 1 9 9 1 9 9 0 1 9 1 9 9 9 0 15 13 9 12 9 1 9 9 0 1 9 15 7 9 9 15 1 9 7 9 7 15 15 13 9 9 0 1 9 2 2
80 7 13 8 8 8 9 9 9 0 7 9 1 9 9 0 13 9 0 7 9 0 1 9 9 1 7 15 1 9 15 13 15 9 9 9 0 0 9 1 9 2 1 7 3 9 1 9 0 1 9 9 0 0 1 9 9 1 9 9 9 1 9 9 1 9 0 1 9 1 9 9 9 15 7 9 8 9 1 15 2
44 7 13 7 15 9 1 9 9 1 9 9 0 13 9 0 1 9 3 7 0 9 9 9 14 13 1 12 12 9 1 9 2 7 13 13 15 9 0 13 15 1 9 2 2
48 7 9 1 7 13 9 9 0 10 9 0 7 13 9 15 13 1 15 15 13 1 12 9 13 1 9 15 1 9 7 13 9 9 1 9 9 9 0 0 1 9 9 9 1 12 12 9 2
56 7 13 7 3 9 0 14 13 9 15 7 9 9 9 1 10 9 0 1 9 0 2 7 9 1 9 15 0 0 1 12 9 13 9 0 14 13 1 12 12 9 7 7 13 9 9 1 12 12 9 7 7 9 14 13 2
29 7 13 7 9 0 0 0 1 9 13 9 1 9 9 9 9 9 1 9 9 9 9 15 1 12 1 12 9 2
49 7 13 8 8 2 9 9 9 2 1 0 9 9 9 7 9 1 9 0 1 9 0 7 9 9 13 9 1 9 9 7 13 9 15 1 9 10 9 7 9 15 13 1 9 9 1 9 2 2
39 7 13 7 9 0 1 9 9 13 1 9 1 9 0 1 9 9 7 9 7 9 9 1 9 1 9 9 9 0 1 7 15 13 0 1 9 0 9 2
61 7 13 7 9 0 0 7 9 9 13 1 9 9 13 9 15 13 1 15 9 15 1 9 15 13 1 9 9 0 1 7 9 9 1 9 13 9 9 9 1 10 9 1 9 9 9 9 9 0 1 9 1 9 0 7 9 1 9 14 13 2
8 9 13 12 12 9 0 1 12
30 13 9 0 0 7 9 0 15 0 9 1 9 9 0 2 0 1 7 15 13 1 12 12 9 1 9 12 1 9 2
83 7 13 9 15 13 15 2 9 9 9 0 7 9 9 2 2 7 9 0 1 9 15 0 1 9 0 1 7 9 15 15 13 1 12 12 9 2 13 15 9 0 1 9 1 15 13 14 12 12 9 2 7 9 0 1 9 0 1 0 1 12 12 2 13 15 9 9 1 15 13 12 12 9 2 7 9 9 15 14 13 12 9 2
57 7 13 9 1 9 15 13 1 9 15 12 9 12 1 15 0 2 7 9 0 1 9 13 1 9 9 1 9 7 14 13 1 9 9 13 1 9 7 0 2 0 1 7 9 9 0 15 13 9 15 13 15 9 0 1 0 2
11 9 9 9 9 9 1 9 7 9 1 9
52 13 2 9 9 2 7 9 2 9 1 9 2 1 9 0 13 1 9 15 1 9 9 9 1 9 1 9 15 0 7 14 13 1 9 1 9 0 1 7 13 9 1 9 1 9 9 0 7 2 8 2 2
37 7 13 9 14 13 9 9 9 9 0 1 8 0 7 9 1 8 7 9 15 1 9 0 9 1 9 9 7 9 9 1 12 2 12 2 12 2
43 1 9 0 13 9 8 8 9 0 9 0 8 8 0 1 9 9 1 9 1 9 1 9 9 9 0 13 9 15 1 9 9 9 9 1 9 1 0 9 1 9 8 2
34 7 13 8 7 1 1 10 9 9 2 8 2 0 1 9 0 0 7 9 2 8 2 0 7 9 2 8 8 2 7 9 0 0 2
22 7 13 8 7 9 0 13 9 9 9 1 9 9 9 7 9 9 9 1 9 15 2
12 9 9 1 9 0 1 12 7 9 12 9 12
27 13 9 0 1 9 0 7 9 9 9 7 9 7 0 1 9 1 9 13 9 12 12 7 12 12 9 2
21 7 13 9 7 9 9 13 1 9 9 7 9 7 9 7 9 9 7 9 9 2
58 7 13 9 7 9 9 14 13 7 12 5 1 9 9 1 9 14 13 7 0 2 7 15 15 13 1 9 9 0 1 9 0 15 13 9 15 12 5 9 1 7 15 15 1 12 7 12 5 1 9 0 1 9 0 0 7 0 2
58 7 13 9 8 8 2 9 9 0 7 12 5 1 9 15 13 1 9 13 9 9 15 12 9 2 7 13 1 7 3 12 12 9 13 15 9 1 9 2 0 7 0 9 1 9 9 13 1 9 9 9 0 7 9 9 1 9 2
51 7 13 9 8 1 9 7 9 9 1 9 9 2 9 0 13 1 12 12 9 9 12 1 12 12 9 9 12 2 7 13 9 9 1 9 0 1 12 12 9 9 12 1 7 13 12 12 9 9 12 2
26 7 13 7 15 1 12 9 0 13 9 12 12 9 1 9 0 0 9 1 12 9 0 1 9 9 2
29 7 13 9 9 1 9 1 9 1 12 12 9 9 12 1 12 12 9 9 0 2 7 15 15 13 12 9 0 2
5 7 1 9 0 2
35 13 9 1 9 9 9 0 1 9 9 1 9 13 1 9 9 9 1 9 13 9 9 1 10 13 1 9 7 9 9 1 9 9 9 2
18 7 13 3 7 9 9 13 1 9 9 15 9 0 13 12 12 9 2
17 7 13 0 7 3 12 12 15 1 9 7 9 0 9 9 9 2
22 7 13 1 9 9 0 9 0 15 13 9 9 0 1 9 9 1 9 15 9 0 2
10 9 2 8 8 2 1 9 9 9 0
35 13 9 0 0 0 7 9 9 0 14 13 9 9 8 8 1 9 9 9 9 12 0 0 2 7 7 9 0 0 14 13 9 1 15 2
126 7 13 9 9 9 8 1 9 9 1 9 1 9 0 15 13 1 15 9 1 9 0 15 13 9 15 2 7 3 1 9 9 9 15 13 15 9 8 8 9 9 0 1 7 14 13 9 0 9 0 1 9 1 12 12 9 0 2 12 12 9 2 2 7 14 13 9 9 15 13 1 9 0 7 9 9 1 9 9 9 9 9 0 9 9 9 8 8 1 7 13 9 9 9 9 1 9 9 9 0 15 14 13 9 0 9 9 15 14 13 9 1 9 10 13 1 15 9 1 9 9 7 9 9 8 2
96 7 13 9 1 9 9 9 9 13 9 8 1 15 1 9 8 9 0 13 1 15 9 1 15 15 1 15 1 9 13 15 1 9 7 12 9 2 7 13 1 10 9 9 9 9 9 1 9 9 8 8 2 7 14 13 9 9 9 1 9 0 2 7 13 9 1 9 8 8 1 10 9 7 13 0 9 0 7 15 13 0 9 9 9 9 9 8 7 3 9 1 9 9 9 9 2
9 0 0 13 9 9 1 9 9 0
119 13 9 9 0 0 9 9 0 1 9 9 0 1 9 0 7 13 7 9 15 0 1 12 9 1 9 12 9 1 9 15 0 1 9 12 0 9 1 9 9 15 1 9 1 0 12 9 1 9 7 12 9 1 9 8 0 1 9 15 13 9 15 1 9 9 1 9 9 9 9 9 1 9 0 2 7 13 7 9 1 9 9 1 9 9 0 0 1 9 9 9 7 9 15 1 9 12 5 1 9 9 15 1 9 1 0 1 9 7 9 9 7 9 9 1 9 9 8 2
39 7 13 9 1 9 13 15 9 0 0 0 1 9 2 7 3 9 8 9 1 9 0 1 9 15 9 9 9 9 0 1 12 9 7 9 9 8 0 2
20 7 13 7 10 9 14 13 1 9 0 13 9 9 0 1 9 9 0 0 2
36 7 13 9 1 8 9 9 1 9 7 9 0 7 9 8 8 1 9 0 1 9 9 9 0 2 7 13 8 12 9 1 12 9 1 0 2
77 7 13 9 0 1 9 9 7 9 9 9 9 0 9 8 8 7 9 0 1 9 9 13 9 9 0 7 9 9 9 9 9 13 7 9 0 0 1 9 7 1 15 9 0 1 9 7 9 9 7 7 9 9 9 1 9 0 1 9 0 14 13 7 9 0 13 1 15 9 7 9 0 13 15 9 9 2
73 7 13 8 9 0 15 13 9 0 1 9 9 1 7 15 9 0 0 2 0 1 7 9 9 9 1 9 7 9 15 0 1 9 9 9 8 13 7 9 0 1 9 15 1 9 8 0 1 15 15 13 9 9 1 9 7 9 1 1 9 0 0 1 9 9 9 9 8 7 9 9 9 2
76 7 14 13 8 7 9 9 1 9 0 7 9 1 9 9 12 0 1 9 12 5 1 9 9 1 9 0 1 9 7 3 9 9 9 9 7 9 9 7 9 9 13 1 9 9 7 13 0 1 9 9 9 1 9 9 0 1 9 9 15 1 9 0 0 1 9 9 9 0 1 1 12 9 9 0 2
15 7 13 1 7 9 0 1 15 0 1 9 0 9 0 2
88 7 1 9 15 2 13 9 9 0 0 9 8 8 7 8 9 9 9 9 0 1 9 7 9 9 7 3 9 1 8 9 1 9 1 9 0 7 13 1 9 7 13 9 0 1 9 9 9 0 0 1 9 0 15 14 13 1 9 9 7 1 0 9 9 9 9 0 1 9 9 9 1 9 9 13 1 9 9 9 9 8 1 12 9 1 9 15 2
41 7 13 7 9 9 1 9 9 12 0 1 9 12 5 1 9 9 1 9 0 1 9 13 9 9 9 14 13 9 9 0 1 9 0 1 9 9 15 1 9 2
100 7 13 9 9 0 0 8 8 9 9 0 1 7 15 13 0 1 15 1 9 7 9 13 1 0 9 9 9 1 9 1 0 9 7 1 9 9 7 7 0 13 1 0 15 13 9 9 2 7 13 1 7 9 9 0 1 9 15 13 1 9 0 9 1 8 9 1 9 0 1 9 15 8 7 9 0 1 9 9 0 1 9 8 8 7 9 9 8 8 1 9 9 0 1 9 9 1 9 0 2
36 7 13 9 9 0 1 9 1 9 0 7 9 9 9 0 1 9 7 0 2 0 1 9 9 9 0 1 9 1 9 9 1 10 9 9 2
5 12 12 9 2 2
7 9 0 13 1 8 1 9
26 0 9 0 13 1 9 13 7 14 13 9 9 0 1 9 9 7 9 0 1 9 0 0 7 9 2
33 7 9 7 9 9 7 0 12 12 9 14 13 9 1 15 1 1 9 9 7 9 0 1 9 0 1 9 1 9 9 1 9 2
33 7 1 9 0 1 9 9 9 0 0 7 9 9 7 9 0 1 9 9 14 7 9 1 15 1 1 9 9 14 13 0 9 2
20 7 13 15 1 9 9 9 9 1 9 1 9 1 9 9 9 9 0 2 2
41 7 13 9 8 8 9 9 9 0 0 14 13 7 9 9 0 0 1 9 0 14 13 9 1 9 1 9 0 1 9 8 9 1 9 9 9 0 1 9 0 2
11 12 9 0 13 1 9 9 0 0 1 9
92 13 12 9 0 0 9 9 0 9 9 0 7 9 0 1 9 0 1 9 0 1 10 9 12 1 9 9 0 15 13 9 9 0 1 9 9 1 9 9 0 1 9 9 1 9 9 15 13 1 12 5 1 9 9 1 9 0 0 1 12 5 3 9 0 7 3 9 9 1 9 1 9 7 9 9 1 9 7 9 0 0 0 1 9 7 9 0 7 3 9 0 2
59 7 13 9 1 9 9 9 0 7 9 13 1 9 9 0 0 1 9 0 9 9 0 7 1 9 9 0 13 1 9 0 1 9 1 9 7 15 1 9 9 1 9 9 1 9 7 9 0 1 9 1 9 7 9 9 1 9 0 2
85 7 13 9 9 0 1 9 9 9 8 8 7 9 13 1 9 0 1 9 9 15 1 9 0 14 9 15 0 7 0 9 15 14 13 1 9 9 0 0 1 9 9 9 1 9 9 0 7 3 9 15 1 9 9 15 0 1 9 0 1 9 1 9 9 0 0 7 9 13 9 9 9 1 9 0 7 1 0 9 9 15 1 9 0 2
23 7 13 7 9 0 14 13 9 9 0 1 9 12 7 12 9 7 13 1 1 9 9 2
82 7 14 13 9 9 9 9 9 0 8 8 9 9 0 0 9 1 9 0 8 1 9 9 9 9 1 9 7 9 1 9 9 0 1 9 0 0 9 0 7 10 9 14 13 9 9 1 9 9 0 13 9 15 1 9 7 9 0 7 14 13 9 0 1 9 9 9 1 9 9 7 9 1 9 1 9 7 9 15 1 9 2
74 7 13 9 9 0 8 8 7 9 9 9 13 7 13 1 9 0 7 0 0 1 9 0 9 0 0 1 9 9 15 13 9 1 8 9 15 1 9 0 1 9 0 0 7 15 14 13 7 8 9 0 0 1 9 7 9 9 1 9 9 3 9 9 7 9 0 1 9 0 7 9 9 9 2
44 1 9 15 13 9 0 9 9 0 8 8 7 9 13 9 7 9 0 1 9 9 9 0 7 9 13 1 10 9 1 9 0 7 13 1 1 9 9 0 1 9 9 0 2
56 7 13 1 7 9 9 0 14 13 9 0 9 1 9 7 13 1 9 0 7 9 0 1 9 9 7 13 7 9 9 9 0 1 15 13 9 15 0 1 9 0 14 13 0 1 9 9 9 1 9 1 9 1 9 0 2
48 7 13 1 9 9 0 7 13 1 15 1 9 9 9 1 9 0 1 9 9 7 9 0 1 15 1 9 9 7 14 13 9 9 0 15 13 9 0 1 9 9 1 9 0 1 9 13 2
5 12 12 9 2 2
4 9 9 8 8
38 13 9 0 1 9 9 0 1 9 9 9 0 1 9 8 8 1 9 1 9 1 9 0 1 12 12 9 1 12 12 9 1 9 9 1 9 12 2
6 13 9 9 12 5 2
25 13 9 1 9 12 12 9 9 0 1 12 12 9 1 9 9 1 9 12 1 9 13 12 5 2
21 7 13 9 0 12 12 9 1 12 12 1 9 9 1 9 12 1 9 12 5 2
25 13 9 0 1 10 9 9 1 9 9 9 13 12 12 9 1 12 12 1 9 9 1 9 12 2
25 13 9 1 8 1 9 0 7 9 7 9 0 2 7 9 2 7 9 2 7 9 9 7 9 2
10 9 0 1 9 13 12 12 9 1 12
39 13 9 9 0 1 9 12 12 9 2 12 12 9 2 1 9 0 12 7 13 9 10 13 1 12 12 9 1 9 9 0 9 1 9 15 1 9 0 2
63 7 13 9 9 0 14 13 1 9 0 15 13 1 12 12 9 1 0 1 9 0 7 9 9 0 15 1 9 9 7 9 7 9 7 9 1 9 7 9 7 9 9 0 15 13 9 15 1 9 0 7 0 7 14 13 9 0 1 15 1 10 9 2
80 7 13 9 0 1 9 9 0 1 7 9 9 13 1 9 0 9 12 12 9 9 1 9 1 9 9 15 1 9 14 7 9 0 1 15 13 9 7 13 9 9 0 1 15 1 7 13 9 15 1 9 0 9 9 0 7 9 14 7 0 15 13 1 9 0 7 9 0 1 15 13 9 1 15 1 9 9 1 9 2
79 7 13 9 9 8 8 8 8 7 9 9 15 13 9 9 1 9 15 10 9 13 1 12 12 9 13 9 1 9 9 7 7 12 12 15 14 13 9 15 1 9 14 13 9 0 8 8 7 9 0 1 8 13 9 15 7 13 9 1 15 1 9 9 1 9 7 9 0 7 9 0 1 15 13 1 9 9 9 2
9 9 13 1 9 8 0 1 9 9
37 13 0 1 9 1 9 9 9 0 0 1 9 9 9 1 9 0 0 9 15 7 1 9 0 2 7 15 1 9 9 15 13 1 15 9 0 2
65 13 10 9 1 9 15 13 1 15 9 0 9 0 1 9 1 7 15 1 9 1 9 15 13 1 15 9 9 0 2 7 7 15 13 1 9 10 9 0 2 7 13 8 8 9 9 9 9 0 7 9 13 1 9 0 1 9 9 9 7 9 9 1 15 2
34 7 13 8 8 9 0 7 9 9 9 9 0 8 8 7 9 13 9 0 9 9 0 1 9 15 9 1 9 7 9 7 9 15 2
42 7 1 9 15 13 8 8 9 1 9 9 1 9 9 1 9 9 7 9 14 13 1 9 0 1 9 9 9 0 1 9 7 9 1 15 14 13 1 15 9 0 2
20 13 7 9 9 9 9 9 13 1 9 9 1 9 9 0 1 9 9 9 2
54 1 9 15 1 8 9 9 9 8 8 7 9 0 1 9 9 7 14 14 13 9 9 1 9 9 15 13 8 1 7 8 13 1 9 9 1 9 0 7 1 12 5 1 8 1 10 9 8 1 9 9 1 9 2
20 9 9 0 1 9 12 5 1 9 1 9 9 9 7 9 15 1 9 9 9
66 13 9 9 1 9 9 0 1 9 9 9 1 9 7 13 15 0 7 15 9 0 1 9 9 9 15 13 9 0 1 9 0 7 9 9 1 9 9 9 7 9 0 7 0 2 7 13 0 1 9 9 9 9 9 7 9 9 9 15 13 1 9 9 1 9 2
61 7 13 9 0 14 13 9 9 9 1 9 0 7 13 12 12 9 7 15 13 12 12 9 2 7 13 0 9 9 9 1 9 9 7 9 1 0 7 15 13 9 9 0 1 9 9 9 7 3 9 9 1 9 9 9 1 9 1 9 0 2
60 7 13 8 8 9 0 1 9 9 0 2 9 2 9 9 15 13 1 9 9 9 1 9 1 15 2 14 9 10 9 15 9 9 9 1 9 7 14 13 1 15 9 0 13 1 15 9 0 15 13 9 15 1 9 0 2 9 8 2 2
38 7 13 8 8 7 13 9 9 9 1 9 1 9 9 9 9 9 7 9 15 1 9 0 3 1 9 7 9 9 7 9 0 7 13 9 1 9 2
64 7 13 8 1 9 9 9 2 9 2 1 9 9 9 1 9 7 9 15 1 9 15 13 1 15 9 0 2 0 2 7 9 9 15 1 9 7 13 7 9 9 9 1 9 0 13 1 9 2 9 2 7 13 1 9 9 1 9 1 9 9 0 0 2
39 1 9 15 13 8 8 9 0 9 0 1 9 0 0 9 9 12 5 1 9 0 1 9 9 9 1 9 2 7 13 7 13 9 1 9 2 9 2 2
55 7 13 7 9 9 1 9 1 9 13 1 12 5 7 15 13 1 15 7 13 1 9 9 9 1 9 1 9 0 2 9 2 7 15 13 7 9 1 15 9 1 9 1 15 7 15 15 13 15 13 1 9 9 9 2
55 7 13 9 9 1 9 1 1 9 9 9 1 9 2 0 7 9 9 9 13 1 9 9 0 1 9 15 13 15 0 7 13 15 2 7 13 1 7 3 9 1 9 9 9 1 15 9 9 9 1 9 0 7 9 2
63 1 9 15 13 8 8 9 0 7 9 9 9 9 9 7 9 9 9 9 1 9 1 9 14 13 1 9 1 9 9 2 7 15 14 13 1 9 2 7 13 1 9 9 9 1 9 9 0 12 2 0 0 2 9 2 9 2 9 2 1 9 0 2
29 7 13 7 3 9 0 1 9 9 1 9 0 2 7 13 9 9 1 9 9 1 9 1 9 9 9 1 9 2
25 7 13 7 9 9 0 9 1 0 1 9 9 2 7 13 15 1 9 15 1 9 9 1 9 2
35 7 13 1 9 9 1 9 9 0 1 9 9 9 2 9 15 13 1 9 9 7 9 2 7 13 1 9 9 10 9 14 1 9 0 2
77 7 13 8 8 9 0 9 7 9 9 1 9 0 0 9 9 9 1 9 1 9 0 1 9 0 1 9 9 1 9 9 0 1 9 9 9 0 2 9 2 7 13 7 9 14 13 1 9 9 9 0 2 7 9 9 9 2 7 9 1 9 9 7 9 2 14 7 15 13 9 0 1 9 0 1 9 2
37 7 13 7 8 9 9 9 1 9 1 9 14 13 1 9 2 14 13 9 1 9 2 7 13 9 8 0 2 1 9 2 1 12 1 12 5 2
80 7 1 9 0 13 8 8 0 9 9 0 0 7 9 9 9 13 9 1 9 9 9 0 9 12 7 13 9 1 9 0 0 7 13 9 9 9 1 9 1 9 2 0 1 7 9 9 13 0 0 1 9 9 2 7 7 3 8 1 9 9 7 9 1 9 7 9 1 9 0 15 13 9 15 7 13 9 9 9 2
72 7 1 9 0 13 8 8 9 9 0 0 7 9 9 9 9 0 7 9 1 9 9 12 13 1 9 7 7 15 13 13 1 9 9 1 9 0 7 0 1 10 9 13 1 9 9 9 7 9 9 1 9 0 1 9 2 0 1 7 9 9 9 13 1 9 9 9 1 1 12 5 2
79 7 13 9 9 9 9 7 15 1 9 8 9 9 9 1 9 13 1 15 9 0 9 9 9 1 9 1 9 9 9 2 7 7 8 8 1 9 9 9 7 15 15 13 9 0 1 9 9 1 9 1 9 9 9 9 1 15 1 9 9 1 9 9 0 7 13 1 8 9 0 15 15 9 0 1 9 9 0 2
35 7 13 8 8 9 9 9 9 0 0 7 9 9 13 15 0 1 9 15 13 1 9 9 7 9 7 9 1 9 9 1 9 9 9 2
36 9 9 0 1 9 7 9 0 1 9 15 0 13 9 9 15 0 15 14 13 15 1 9 0 1 9 9 9 1 8 1 9 7 9 0 2
24 7 13 9 0 7 9 0 13 1 9 0 1 9 0 9 14 13 1 9 9 9 9 0 2
52 7 13 7 3 9 1 9 9 0 9 1 10 13 1 15 1 9 2 0 1 9 8 1 9 9 0 1 9 9 0 9 0 2 7 15 0 2 1 9 9 9 0 15 13 9 1 9 15 1 9 12 2
22 7 13 9 0 13 9 9 9 0 0 1 9 9 1 9 9 0 7 0 1 9 2
16 7 13 9 9 9 0 13 9 1 9 9 0 2 7 13 2
34 2 14 13 9 2 1 9 2 1 9 0 2 2 0 1 7 8 13 1 9 12 1 15 13 1 9 9 0 15 13 9 9 15 2
15 7 13 2 2 14 13 9 9 9 1 9 1 9 0 2
29 13 9 0 1 9 9 0 0 9 1 15 7 15 14 13 1 9 0 0 7 9 9 9 1 9 9 0 2 2
65 7 13 2 2 7 8 8 9 9 14 14 8 9 2 1 9 9 1 9 1 9 0 1 9 7 9 0 2 0 7 15 2 13 9 2 7 7 15 13 1 9 7 9 0 2 9 0 2 9 1 9 0 1 9 7 9 7 7 9 0 7 14 13 3 2
25 7 13 2 2 13 9 9 0 1 9 1 1 9 9 0 7 0 1 9 7 9 9 1 9 2
17 8 8 1 10 9 2 8 7 8 14 8 9 1 10 9 2 2
54 7 13 9 1 7 9 9 0 1 8 14 13 9 9 9 1 9 1 9 0 0 2 9 7 9 13 9 9 9 1 9 9 9 9 9 2 7 14 13 9 12 9 9 0 1 9 9 0 0 1 9 9 0 2
54 7 13 1 9 9 1 9 1 9 9 9 0 7 9 9 9 0 1 9 15 13 1 9 2 0 1 7 15 1 0 7 13 9 9 0 0 1 9 1 9 1 9 0 1 9 9 1 10 13 15 9 1 9 2
26 1 15 13 9 0 1 9 9 9 9 0 8 8 9 9 0 7 9 9 0 1 9 1 9 0 2
36 7 13 1 9 15 7 13 9 0 9 9 9 0 1 9 7 3 9 9 0 7 15 1 9 15 7 13 9 0 1 9 9 0 1 9 2
26 7 13 9 1 7 3 9 1 9 9 9 0 7 0 1 9 1 9 9 9 7 9 0 1 15 2
10 9 9 9 0 1 9 7 9 9 8
59 13 8 2 8 8 8 9 9 0 9 1 9 8 1 9 9 13 9 9 0 1 9 9 9 9 9 0 7 0 7 0 1 9 13 9 9 9 1 9 9 9 0 1 9 9 0 1 9 8 2 8 2 7 15 13 15 9 8 2
4 7 13 8 2
52 8 1 9 2 8 2 9 0 1 9 9 0 1 9 0 9 7 9 9 9 9 15 13 1 9 0 1 9 9 1 9 9 0 7 9 9 9 9 15 1 9 0 1 10 13 9 9 0 1 10 9 2
30 7 13 9 9 9 1 9 8 8 8 9 9 9 0 9 1 9 15 1 9 8 1 9 9 9 7 9 1 9 2
61 7 13 8 2 8 7 9 13 9 9 0 1 9 7 9 8 0 1 9 0 7 14 13 1 15 9 9 9 1 9 1 9 9 9 1 9 9 7 9 1 9 9 1 9 0 1 9 7 9 8 9 0 7 0 1 9 9 9 1 15 2
8 9 13 1 9 9 9 9 9
79 13 9 12 2 12 0 9 0 8 8 9 1 9 9 9 8 8 1 9 9 15 0 8 8 7 9 9 1 9 0 8 8 8 7 9 9 1 9 8 8 2 7 13 8 1 9 1 9 2 2 13 9 7 9 1 9 2 7 9 0 1 15 2 9 9 0 0 7 9 0 1 9 0 1 8 7 9 2 2
53 7 13 2 2 13 9 3 9 0 1 9 7 9 2 7 13 9 9 9 9 0 2 7 13 9 0 7 9 15 0 1 15 13 1 9 7 13 1 9 1 9 9 1 15 7 13 9 15 9 9 15 2 2
41 7 1 9 15 13 8 1 7 13 1 7 9 0 1 9 7 9 2 13 1 9 0 13 9 15 13 9 8 1 9 9 9 8 8 1 9 1 9 0 2 2
35 7 13 7 9 0 1 9 13 9 0 2 1 9 9 9 0 1 9 9 7 9 9 9 1 9 2 7 9 9 9 9 9 1 9 2
29 7 13 7 3 2 9 0 1 9 7 9 1 9 9 2 1 9 9 0 2 1 9 9 9 1 9 0 2 2
22 7 13 7 9 1 9 2 0 7 0 1 1 2 7 13 9 7 9 7 9 2 2
10 9 9 13 9 0 0 1 9 9 15
68 13 9 9 9 1 9 15 9 12 2 12 0 9 15 9 9 9 9 0 7 13 12 7 2 12 2 12 9 2 13 9 7 9 15 13 1 9 15 9 9 0 7 15 13 1 9 9 2 13 9 14 13 9 9 1 9 12 0 1 9 9 0 0 1 9 12 9 2
14 13 9 7 10 9 14 13 9 0 15 13 15 9 2
24 7 13 9 9 7 9 1 9 1 10 9 2 7 13 15 1 9 7 9 1 9 9 0 2
10 9 0 7 9 0 13 9 0 1 9
42 13 9 1 9 1 9 9 0 15 13 15 9 0 0 1 9 9 2 7 13 9 9 9 1 9 9 0 1 9 13 9 9 0 1 9 1 9 9 9 1 9 2
26 7 13 9 0 1 9 0 9 9 8 8 13 9 9 12 2 12 0 7 9 9 9 9 8 8 2
70 7 13 1 9 13 1 9 7 9 2 13 9 15 1 9 9 0 7 9 1 15 1 9 15 13 9 9 2 2 7 7 15 2 13 9 1 9 9 0 13 9 9 0 1 9 9 7 9 7 9 9 0 2 7 13 9 2 9 0 2 1 9 9 15 9 0 7 9 0 2
41 7 13 9 0 1 9 7 9 13 0 0 1 7 15 2 1 15 9 1 9 9 0 7 9 15 1 9 9 9 0 7 0 7 0 7 9 1 9 0 2 2
27 7 13 9 9 0 13 9 9 9 0 1 9 9 0 2 1 7 8 9 9 0 8 8 8 1 9 2
44 7 13 7 8 14 13 2 1 9 0 2 9 9 0 1 9 0 1 9 9 9 9 1 9 1 9 9 9 0 1 9 1 9 0 1 9 0 9 15 1 9 9 9 2
31 7 1 0 7 13 9 9 9 7 9 7 9 0 2 7 9 0 7 9 9 15 7 9 9 1 9 0 9 7 0 2
18 9 0 1 9 9 13 9 0 1 7 15 13 2 9 0 2 1 9
81 1 9 15 13 1 15 9 0 0 1 9 1 9 9 0 1 10 13 15 2 9 0 2 1 9 0 0 0 2 1 9 0 13 15 1 9 9 0 7 9 0 2 13 9 9 9 1 9 9 8 1 9 2 7 13 15 2 9 9 0 7 9 9 0 1 9 0 0 1 7 9 0 13 1 9 1 9 7 9 2 2
9 9 0 9 0 0 13 15 9 0
55 13 9 9 0 0 9 12 2 12 0 1 9 0 9 0 1 9 7 9 9 2 7 13 9 2 9 0 1 9 7 9 9 2 13 0 15 7 15 13 1 2 9 9 9 9 7 9 1 15 7 9 1 15 2 2
37 7 13 1 9 9 12 1 9 9 0 0 1 9 12 1 0 1 9 13 1 0 9 2 7 13 9 9 1 9 9 9 1 0 7 9 0 2
15 9 13 1 9 9 13 1 9 9 1 9 7 9 1 0
80 13 9 1 9 0 1 9 9 1 9 2 9 9 2 13 1 9 9 1 9 0 7 9 1 15 1 9 15 0 2 1 15 8 8 2 8 8 2 7 9 8 8 2 7 9 8 8 2 8 8 8 8 2 8 8 8 8 13 15 9 0 1 9 8 8 2 12 9 2 9 8 8 8 8 9 7 9 0 0 2
58 7 14 13 8 8 8 7 9 9 0 0 0 1 2 9 0 2 7 15 13 9 0 1 9 9 9 7 14 13 1 9 9 9 1 9 9 15 1 9 0 2 0 1 7 9 0 13 1 9 12 7 15 9 0 1 9 9 2
55 7 13 7 13 9 9 9 9 1 9 9 15 1 9 9 9 0 7 14 13 1 9 2 0 1 7 2 9 0 0 9 1 9 13 1 9 1 9 2 1 9 15 13 1 15 2 9 1 9 7 9 1 15 2 2
56 7 13 7 9 1 9 13 1 9 9 2 7 9 9 2 7 7 15 9 7 13 9 7 14 13 9 1 15 7 9 9 1 9 7 9 2 9 0 2 9 9 2 7 9 9 2 7 9 9 7 15 14 13 0 2 2
23 7 13 7 9 2 13 1 9 9 1 9 2 8 8 8 8 1 9 9 8 8 2 2
6 9 1 9 1 9 9
73 1 9 9 0 0 1 9 9 1 9 9 9 0 2 2 9 9 2 14 7 9 13 9 7 9 0 9 12 2 12 0 1 9 9 12 13 1 9 1 9 9 0 15 13 1 9 9 0 1 8 0 2 7 9 12 0 1 9 9 1 9 9 9 1 9 1 9 15 1 9 9 15 2
36 7 13 9 1 9 9 0 9 9 9 9 1 9 1 9 2 7 7 9 15 13 15 9 1 9 9 8 2 8 2 9 1 9 13 9 2
54 7 13 9 8 8 9 9 0 1 9 0 1 9 7 9 0 13 1 9 9 9 0 15 13 1 9 9 0 2 7 13 9 9 9 0 1 15 1 9 8 9 1 9 2 1 9 9 9 0 1 9 1 15 2
72 7 13 7 9 9 13 9 0 1 9 9 9 1 9 2 1 9 0 1 9 7 9 9 0 1 9 9 8 7 9 15 1 0 2 9 1 9 8 2 8 2 2 0 1 9 12 12 9 1 9 9 8 1 9 2 7 1 7 9 0 13 9 0 1 9 9 9 8 0 1 9 2
59 7 13 9 8 8 9 9 9 9 0 1 9 7 9 9 9 1 9 9 0 7 9 0 8 8 8 9 9 13 9 9 15 1 9 9 9 1 9 15 1 9 0 8 1 9 0 1 9 9 0 15 13 1 12 1 12 9 0 2
19 7 13 9 9 8 8 7 9 15 8 8 1 9 9 9 1 9 9 2
13 9 2 9 9 8 8 1 9 9 7 9 8 9
27 13 9 1 9 9 9 1 9 9 1 9 9 1 9 9 7 0 9 15 13 9 9 9 1 0 0 2
26 13 9 0 1 9 9 9 15 13 15 1 12 7 12 9 8 13 9 9 0 1 9 0 3 2 2
15 7 9 0 7 9 9 9 9 10 1 9 7 0 2 2
24 1 15 1 10 9 9 7 9 9 9 0 3 1 9 9 7 9 7 9 9 7 0 9 2
27 7 13 9 1 9 9 9 0 1 9 9 1 9 9 1 15 1 9 9 9 9 0 1 9 8 2 2
20 7 13 1 9 9 1 9 9 9 8 0 1 9 9 1 9 9 15 2 2
62 7 13 7 15 1 9 9 0 13 7 9 0 1 9 7 9 10 9 1 8 1 9 0 7 9 15 7 9 15 0 1 9 1 9 9 7 15 13 1 15 1 9 9 9 0 0 1 9 14 13 7 15 14 13 9 14 12 5 1 9 0 2
16 7 13 9 7 1 9 15 8 8 8 8 8 8 7 13 2
40 8 8 7 15 1 9 13 7 3 9 13 9 9 9 1 15 10 1 12 7 12 7 9 12 9 9 1 9 9 9 8 0 1 10 13 14 12 12 9 2
9 12 5 1 9 9 1 9 1 9
28 13 9 9 9 0 7 9 9 1 9 9 9 1 9 13 12 5 2 1 15 13 12 12 7 12 12 9 2
31 13 9 7 12 5 1 9 8 1 9 2 7 12 5 1 15 8 1 9 2 7 7 12 5 1 0 1 9 1 9 2
9 13 8 9 8 8 9 1 9 2
5 9 8 3 2 2
4 13 1 9 0
37 1 9 0 2 13 2 9 8 2 15 9 9 9 2 13 1 9 15 9 9 7 9 0 2 7 13 1 9 15 9 1 9 7 9 9 2 2
15 9 10 9 13 9 9 10 9 2 7 9 9 0 15 2
12 7 15 15 13 9 1 9 15 1 10 9 2
12 7 9 9 1 9 0 13 9 0 1 15 2
44 14 14 13 1 15 7 13 1 9 0 1 9 9 12 0 2 7 13 13 1 9 2 9 2 7 13 0 1 15 7 13 13 15 1 9 0 13 1 9 2 9 9 2 2
43 7 13 9 1 15 1 9 0 2 7 13 1 9 0 7 0 0 1 9 9 7 9 7 13 9 13 1 9 1 15 1 9 8 1 9 7 0 7 13 1 9 15 2
25 7 1 9 0 1 9 2 13 9 9 13 9 0 1 9 9 9 1 9 15 7 9 1 15 2
55 7 10 9 13 9 1 9 9 12 7 1 9 9 2 7 9 9 9 0 7 9 9 0 0 13 1 9 9 15 1 9 9 2 13 9 9 1 9 9 9 1 9 0 2 7 13 1 9 2 8 2 7 12 9 2
20 8 8 2 9 9 9 1 9 9 9 2 13 9 9 9 8 10 9 2 2
34 7 13 9 1 9 0 10 9 15 13 13 15 9 9 9 0 2 1 9 9 9 2 7 13 13 1 15 0 15 13 1 12 9 2
13 13 8 8 2 7 10 9 14 13 10 9 2 2
14 7 9 15 13 13 1 15 13 1 15 9 0 0 2
20 13 8 8 10 9 1 9 2 0 9 0 1 9 7 13 9 10 9 0 2
27 14 9 0 7 15 9 0 9 0 10 9 1 9 1 9 1 10 13 13 10 9 2 0 1 9 9 2
6 9 7 9 9 2 2
5 9 0 0 2 2
29 13 0 1 12 9 1 9 0 9 9 9 2 7 13 9 1 0 0 2 7 13 1 15 1 9 13 1 9 2
17 13 12 9 1 9 0 1 9 15 1 9 1 9 7 9 0 2
31 7 13 9 0 1 8 9 2 7 15 2 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 2
32 13 9 14 13 9 1 9 1 9 9 13 1 9 9 1 9 9 9 7 9 9 1 9 9 7 9 1 9 0 7 0 2
22 13 9 9 9 8 8 8 7 10 9 13 9 1 9 0 0 7 13 9 9 0 2
4 9 9 1 9
25 13 9 0 1 9 9 1 9 0 13 1 9 1 9 0 1 9 7 9 7 9 7 9 2 2
28 7 15 15 13 1 9 15 1 9 2 9 2 9 7 9 9 15 0 7 13 9 1 9 14 9 1 15 2
28 13 9 1 7 9 0 13 9 12 15 13 1 12 12 7 12 9 1 8 1 9 12 12 7 12 12 9 2
36 7 7 15 13 9 9 9 9 9 1 9 0 1 9 9 9 1 9 9 12 9 7 7 9 9 9 13 12 7 12 12 7 12 9 2 2
34 7 1 9 9 0 1 9 0 1 9 13 9 0 1 9 9 12 7 13 1 12 12 7 12 9 1 9 12 12 7 12 12 9 2
38 7 7 15 13 9 9 9 1 9 0 7 1 9 9 9 1 9 12 9 7 7 9 13 1 12 7 12 12 7 12 12 9 1 9 7 9 2 2
51 7 0 7 9 0 1 9 0 12 13 1 9 9 9 9 7 13 1 12 12 9 7 15 13 1 9 0 1 9 9 0 7 15 12 9 1 9 15 13 1 12 12 7 12 12 7 12 12 9 2 2
21 8 8 13 7 9 8 1 1 9 13 2 2 8 2 8 1 9 9 2 8 2
23 7 7 8 1 9 9 0 1 9 7 9 7 9 7 9 15 8 8 7 9 0 2 2
31 1 9 0 7 13 9 12 12 9 1 9 10 9 1 9 12 12 9 7 15 13 12 7 12 12 7 12 9 2 2 2
43 7 1 9 9 0 0 1 12 9 0 13 9 9 0 1 9 7 9 7 9 9 7 9 1 10 13 12 12 9 7 15 13 12 12 7 12 12 7 12 12 9 2 2
2 2 2
3 14 9 2
36 7 7 15 13 9 9 9 0 1 9 9 15 13 15 9 0 14 13 15 13 9 0 9 15 15 13 12 7 12 12 7 12 12 9 2 2
16 7 13 1 12 12 7 12 12 7 12 12 9 1 9 0 2
9 8 13 1 9 9 9 0 1 9
21 13 9 8 8 9 9 9 0 2 9 9 0 0 1 9 9 9 0 1 9 2
20 13 2 8 2 1 7 9 14 13 1 9 9 9 9 0 7 9 7 9 2
19 7 13 2 8 2 1 9 0 1 2 9 2 9 9 0 0 1 9 2
14 7 1 0 7 13 1 12 12 9 0 1 9 12 2
20 7 13 9 0 1 9 9 9 9 0 1 9 15 13 1 9 9 1 9 2
26 7 13 7 9 9 14 13 9 1 9 0 1 9 0 1 9 9 2 14 1 1 9 1 9 0 2
26 7 13 2 8 2 1 7 9 15 13 0 1 9 0 1 15 13 1 9 9 1 9 7 9 9 2
33 7 13 9 0 7 9 9 0 1 9 14 13 1 9 0 9 9 9 7 9 0 7 9 7 9 7 15 13 13 15 1 9 2
25 7 13 7 13 9 0 1 9 9 9 9 7 7 15 14 13 0 9 1 9 1 9 10 9 2
20 7 13 9 9 9 0 7 13 1 9 15 0 9 1 9 9 9 1 9 2
16 7 13 7 9 15 14 13 9 9 1 9 9 1 9 0 2
15 2 9 2 13 1 9 9 9 15 7 9 9 15 1 9
28 13 9 15 13 15 9 0 0 1 9 1 9 9 9 1 9 9 0 1 9 1 9 7 2 9 0 2 2
75 7 13 1 9 15 13 15 9 0 1 9 9 9 0 7 9 0 7 9 13 1 9 2 9 2 4 3 1 9 15 1 9 1 9 2 7 7 3 9 9 9 1 15 2 7 9 9 9 9 1 1 9 15 1 9 1 9 1 2 9 2 9 7 9 2 1 9 9 9 15 1 9 7 9 2
28 7 13 7 9 13 1 9 9 0 1 9 9 9 0 1 2 9 2 2 7 9 9 9 1 9 9 15 2
35 7 9 0 1 2 9 2 13 1 2 9 2 7 2 9 13 7 15 14 13 1 0 9 0 1 9 9 9 7 9 9 9 15 2 2
58 7 13 1 7 9 9 13 13 1 2 9 2 1 9 0 9 12 2 7 13 1 2 9 2 1 9 9 9 1 9 15 13 1 15 9 9 1 9 9 0 0 2 0 1 7 9 2 9 2 1 9 9 9 13 9 1 9 2
75 7 13 2 9 2 7 9 9 2 7 15 0 9 1 9 2 13 9 1 9 1 9 9 1 9 9 0 15 13 2 9 2 1 9 9 2 7 7 9 0 14 13 9 0 1 9 9 2 13 1 9 13 9 1 9 1 9 15 1 9 9 0 2 7 0 9 9 0 9 1 9 1 9 0 2
53 7 1 9 9 1 9 2 9 2 14 7 9 13 1 9 7 9 9 7 9 1 9 9 15 14 13 1 9 0 1 9 0 7 9 9 7 13 9 0 0 9 1 9 9 9 9 2 7 3 9 9 0 2
14 9 9 9 13 9 9 1 9 9 1 9 9 2 2
7 7 13 15 1 9 0 2
12 13 9 9 9 0 1 9 9 1 9 0 2
27 13 9 9 1 9 0 1 9 1 9 9 0 1 9 9 9 1 9 9 1 9 1 9 9 1 9 2
52 13 9 7 9 7 9 13 1 9 9 0 1 9 1 9 15 13 9 0 7 13 13 9 9 9 1 9 9 1 9 9 13 1 15 15 9 1 9 0 1 9 9 1 9 9 1 9 7 9 9 0 2
41 7 13 9 9 0 1 9 9 0 1 9 9 7 9 13 1 9 12 9 9 1 9 0 7 14 13 1 12 9 3 1 9 0 1 7 0 13 1 9 9 2
44 7 13 9 7 9 0 15 0 0 1 9 9 0 1 9 9 0 7 13 9 9 0 1 10 9 7 1 9 9 13 9 9 1 9 9 0 1 9 9 1 9 0 2 2
10 12 12 9 13 1 9 9 9 1 9
44 13 0 0 0 9 0 1 9 0 1 9 9 0 1 9 9 1 9 9 7 9 1 12 12 9 13 1 9 1 0 1 12 9 2 7 1 15 13 0 0 9 9 9 2
56 7 13 9 0 0 7 0 1 12 5 1 10 9 15 9 9 0 1 9 0 13 1 9 0 1 9 7 15 13 1 9 1 9 0 8 8 2 8 8 9 1 9 9 7 9 1 9 7 0 0 1 9 0 1 9 2
69 7 13 10 9 7 15 13 1 9 0 1 0 9 0 1 9 0 7 7 0 1 9 15 15 13 14 13 1 15 9 1 9 9 0 2 0 8 2 1 13 0 15 13 1 9 2 9 2 10 1 9 7 0 2 7 13 1 9 0 9 0 7 9 9 1 9 0 3 2
68 7 13 9 7 9 0 13 1 9 9 0 1 7 9 0 1 9 9 1 9 0 7 0 7 13 15 9 9 9 0 1 1 13 9 1 9 10 1 9 2 9 7 0 1 12 5 1 9 9 1 14 12 9 0 13 1 9 0 2 7 3 9 0 7 1 9 0 2
44 7 13 10 9 1 7 15 1 0 7 13 9 1 9 0 1 9 9 1 9 9 0 1 10 15 13 1 9 9 7 9 7 9 7 9 15 1 9 9 1 9 9 0 2
24 7 13 9 0 7 9 9 9 9 14 13 1 9 0 1 9 0 1 9 9 15 0 0 2
13 9 9 1 9 13 1 9 13 9 9 0 1 9
51 13 9 1 9 9 0 2 0 1 8 8 8 8 2 8 8 0 1 9 9 1 9 1 9 0 2 1 9 15 13 15 9 9 9 8 8 0 1 9 9 9 0 7 9 9 9 0 1 9 9 2
124 7 13 9 9 1 9 15 7 2 9 9 13 1 9 9 1 9 0 1 0 2 7 9 15 0 13 1 9 1 9 9 7 13 1 9 15 9 0 2 7 1 9 15 13 9 8 1 9 15 2 7 13 1 2 8 8 2 7 15 13 13 1 1 15 1 9 9 9 15 13 9 9 0 1 9 9 9 15 13 9 9 1 9 2 0 1 9 9 1 15 1 9 9 2 7 1 7 13 9 15 1 9 9 1 9 0 9 1 15 2 7 1 9 10 9 7 9 1 9 0 8 1 9 2
17 8 13 9 1 9 1 9 15 8 8 2 8 8 2 1 9 0
48 13 9 9 0 0 2 8 2 9 0 1 9 1 9 9 0 2 8 8 8 8 9 9 0 1 9 1 2 8 8 2 0 7 14 9 2 9 2 1 9 9 7 1 9 1 9 0 2
40 7 13 9 1 9 9 9 1 9 2 13 10 9 7 9 13 9 0 1 9 1 8 7 8 7 8 7 9 8 8 7 1 10 9 13 9 9 0 0 2
53 7 13 9 9 2 8 8 2 0 7 9 2 9 2 7 15 13 8 8 9 3 1 9 0 1 9 9 9 9 9 1 9 7 2 8 8 2 8 8 7 13 9 1 9 1 9 1 9 15 1 9 9 2
31 7 13 8 1 9 0 9 9 0 1 10 13 15 1 10 9 9 0 2 7 1 9 1 10 13 9 0 1 9 0 2
11 7 9 13 3 9 7 3 9 9 0 2
15 9 0 13 9 0 7 13 15 13 9 15 1 9 2 2
3 9 2 2
51 13 9 0 9 8 8 8 9 1 9 0 8 8 0 7 13 7 15 13 9 15 1 9 1 9 0 7 13 9 9 0 7 14 13 1 15 9 1 9 9 1 9 9 15 15 9 2 9 2 9 2
61 7 13 7 15 13 9 15 1 9 7 9 7 9 2 7 0 2 8 8 14 8 1 15 2 7 13 8 7 13 3 9 1 0 0 7 13 10 9 9 1 9 1 15 8 8 8 1 15 8 13 9 15 1 0 9 1 9 0 1 0 2
151 13 8 9 0 15 13 1 15 9 1 9 2 8 2 9 1 10 13 15 8 0 7 9 0 1 7 9 0 13 9 8 7 13 15 1 0 7 7 9 8 2 8 8 13 15 7 13 9 1 12 9 1 9 15 2 9 15 13 15 9 0 9 7 13 7 9 0 8 8 0 7 14 8 1 8 8 8 8 0 2 7 7 13 1 15 9 7 9 1 10 9 0 7 7 13 15 8 8 2 7 13 9 0 7 15 3 7 8 8 9 0 8 8 9 15 7 7 13 7 13 1 8 8 9 8 8 9 2 9 2 9 2 7 14 8 1 15 7 8 8 9 9 15 2 7 9 15 1 8 8 2
11 9 0 13 1 9 9 0 1 9 9 9
28 13 9 0 9 1 9 1 9 9 1 9 1 9 0 7 9 13 1 15 7 13 1 9 12 9 1 9 2
52 7 13 9 9 0 1 9 9 1 9 9 13 13 7 13 1 9 0 2 7 13 9 9 1 9 9 15 13 0 1 9 0 1 9 9 7 13 9 9 0 9 13 1 9 1 9 9 7 9 9 0 2
32 7 13 9 1 9 13 1 9 8 0 1 9 8 9 9 1 9 1 9 1 9 13 9 9 9 15 1 9 1 9 15 2
46 7 13 9 0 7 9 13 9 15 13 1 9 0 1 9 1 9 9 9 7 13 1 9 1 9 8 0 1 9 9 15 13 9 1 9 7 9 13 1 9 12 9 7 9 0 2
80 7 13 9 9 9 15 1 9 1 9 1 9 9 9 12 2 12 0 7 13 9 1 9 7 12 9 13 1 9 15 2 8 8 8 2 12 9 2 8 8 8 8 2 12 9 2 8 8 8 8 2 12 9 2 7 8 8 2 12 9 2 8 8 8 8 2 12 9 2 7 13 9 0 1 8 8 8 8 9 2
56 7 13 9 7 9 9 9 13 7 9 9 9 0 13 0 7 13 9 1 9 0 9 9 9 1 9 13 15 9 15 1 9 15 1 9 14 7 9 0 13 2 7 13 1 9 9 1 9 7 9 13 1 15 9 12 2
56 13 9 0 1 2 9 2 7 9 9 0 13 9 1 9 9 9 7 13 12 9 1 9 1 15 2 7 13 9 1 9 9 9 1 9 0 7 0 1 9 8 1 9 10 9 7 14 13 1 9 9 1 9 1 9 2
33 7 13 9 7 9 0 9 1 9 9 1 7 13 9 1 9 7 13 9 9 1 9 7 13 1 9 1 9 9 1 9 9 2
8 9 1 9 9 1 2 9 2
28 13 9 0 1 9 9 1 9 1 9 9 9 0 9 1 9 1 9 0 1 9 15 1 9 9 7 9 2
38 13 9 2 8 8 8 2 9 9 7 9 9 13 9 9 1 9 0 1 9 15 1 9 9 0 15 13 1 10 9 9 9 2 7 9 13 9 2
39 7 14 13 9 0 0 9 1 9 1 9 9 9 1 9 2 7 13 1 15 1 9 9 1 9 1 9 7 9 0 15 13 9 7 13 9 1 9 2
14 7 1 9 15 13 1 15 9 3 9 1 9 9 2
28 7 0 7 15 13 9 9 9 0 1 9 1 9 9 2 1 9 9 9 0 13 9 9 1 9 1 9 2
4 9 13 9 8
21 1 9 14 13 1 9 0 2 13 9 9 0 1 9 9 1 9 0 9 2 2
6 9 9 1 9 9 2
4 14 1 9 2
22 7 15 9 13 7 13 1 9 0 2 7 13 1 9 9 0 1 7 9 9 15 2
29 7 13 9 15 13 9 0 1 9 7 9 7 9 2 9 13 9 1 9 15 2 1 9 1 9 9 0 9 2
24 10 9 0 13 15 9 1 9 9 13 1 9 15 1 9 0 13 7 9 9 13 1 9 2
22 7 13 9 15 7 9 9 7 9 15 0 7 9 1 15 14 13 1 9 0 0 2
24 7 13 9 1 9 0 9 0 1 9 9 15 14 13 9 0 1 9 0 7 1 0 0 2
20 7 13 10 9 15 13 1 9 9 9 7 9 9 9 7 9 9 9 15 2
20 7 15 9 0 13 1 9 0 13 1 9 9 15 1 9 1 9 9 9 2
26 7 13 9 15 13 9 0 1 12 12 9 1 9 15 13 9 8 0 1 9 0 7 0 9 9 2
17 8 7 15 13 9 15 1 9 0 2 7 1 0 9 9 0 2
19 7 13 9 15 1 9 1 9 1 9 7 9 9 0 7 9 9 0 2
31 13 9 1 9 1 9 13 9 7 9 13 9 1 9 15 1 9 0 2 9 0 9 2 7 15 0 1 9 0 0 2
9 14 15 9 0 13 8 8 2 2
37 7 1 9 0 13 9 1 9 7 9 9 0 9 15 1 10 9 1 9 9 2 13 7 9 9 1 1 10 9 13 7 13 1 1 12 5 2
27 7 13 9 8 8 9 7 3 9 0 7 0 0 1 9 8 1 15 9 9 9 1 9 7 9 2 2
23 7 13 7 10 9 0 7 13 1 9 9 9 1 9 9 1 9 0 1 9 1 9 2
19 13 8 2 8 13 1 9 2 12 9 2 7 13 9 0 1 9 0 2
16 2 9 0 9 9 7 7 3 9 7 15 9 1 9 9 2
20 0 7 9 14 13 1 10 9 8 7 15 9 1 9 9 7 9 9 2 2
49 7 13 9 9 0 1 9 7 9 7 9 9 9 1 9 9 13 9 12 1 12 12 9 1 9 0 1 9 0 1 9 1 9 9 9 1 12 12 9 1 9 12 1 12 12 9 1 12 2
55 7 13 9 0 1 9 8 1 9 9 8 0 1 9 15 1 9 0 1 9 0 1 1 12 9 13 9 1 9 9 9 1 9 9 0 1 0 9 1 9 12 2 7 13 9 0 1 10 9 1 9 9 1 9 2
16 7 13 9 9 9 0 1 9 8 0 1 1 12 12 9 2
41 7 1 9 14 13 9 0 0 1 7 13 1 15 12 12 9 9 1 9 1 9 14 7 15 13 9 0 13 9 7 13 1 10 9 7 14 13 15 15 0 2
14 7 13 7 9 14 13 9 9 1 13 9 9 9 2
18 7 13 9 1 7 13 9 9 1 9 7 9 0 1 9 9 9 2
18 7 1 3 7 14 9 13 1 9 9 0 7 0 1 9 9 0 2
15 7 15 13 9 1 9 1 9 1 15 7 13 9 0 2
58 7 8 9 1 9 15 1 9 7 13 9 15 0 1 9 1 9 1 9 0 7 1 7 9 13 9 9 9 0 1 9 7 13 1 10 9 0 8 7 9 13 1 7 13 10 9 1 9 9 9 7 9 0 1 9 1 9 2
9 9 9 13 1 9 9 0 1 9
44 13 9 9 9 9 0 1 9 0 8 8 8 1 9 0 1 9 0 8 8 9 1 9 2 1 9 15 9 0 0 2 7 13 15 9 0 1 9 9 9 15 8 8 2
27 7 13 9 0 14 13 9 9 12 2 12 0 1 9 9 0 1 9 9 1 9 0 2 9 8 8 2
46 7 13 9 0 2 2 1 0 7 13 8 9 0 1 9 0 2 7 13 9 0 2 1 9 9 15 1 9 9 0 2 7 9 0 1 15 2 1 9 9 1 9 10 9 2 2
12 9 9 8 9 9 1 9 9 1 9 15 0
51 14 13 9 15 13 1 9 9 9 8 9 9 9 9 0 2 1 9 15 13 9 9 0 13 15 9 12 2 12 0 8 8 0 1 9 9 1 9 12 9 7 0 7 9 7 9 9 7 9 0 2
32 7 13 9 0 1 9 9 0 1 9 1 7 14 13 9 0 1 9 8 1 9 9 0 0 15 13 15 1 1 12 9 2
64 7 13 9 9 0 0 1 9 0 7 13 9 9 1 9 9 9 15 13 1 15 9 2 9 1 9 9 9 9 1 9 2 7 1 9 15 9 9 8 8 2 7 9 9 9 9 8 8 8 2 7 9 9 9 8 8 8 2 8 8 9 8 8 2
16 8 8 0 1 9 8 1 9 2 7 13 1 9 1 9 2
21 7 13 2 2 14 15 9 0 13 9 9 0 1 9 7 9 1 9 0 2 2
22 8 8 9 0 1 9 0 7 1 9 7 9 8 8 7 13 1 9 7 9 2 2
13 0 1 7 2 8 8 8 9 1 9 8 2 2
36 7 13 2 2 14 9 1 9 9 9 7 9 8 8 9 9 0 8 8 8 8 8 8 0 7 9 13 8 8 7 9 7 9 3 2 2
96 7 1 9 15 13 8 0 1 9 2 2 8 8 9 7 9 8 1 9 7 9 1 9 0 1 9 8 11 8 2 7 13 9 7 9 3 1 9 1 0 13 1 9 7 13 0 9 1 9 2 2 0 1 7 2 9 8 8 1 9 15 7 9 15 1 9 13 15 9 1 9 13 8 9 2 7 14 13 1 15 10 9 9 1 15 1 9 1 7 9 13 9 9 0 2 2
50 7 13 2 2 14 9 9 7 9 13 3 1 9 0 7 13 0 1 9 1 9 12 0 7 9 9 12 2 7 13 3 1 9 9 9 9 12 0 15 13 1 15 9 0 1 9 9 0 2 2
9 9 0 1 9 13 9 7 13 9
28 1 9 15 12 15 13 15 2 13 9 0 0 1 9 8 8 13 1 9 15 13 1 9 9 9 1 9 2
20 7 13 2 8 8 2 7 8 13 1 9 12 1 9 13 1 15 9 13 2
35 7 13 1 9 15 9 9 9 1 9 9 0 1 15 7 9 9 9 7 9 1 9 15 13 13 15 1 9 0 1 9 15 1 9 2
100 7 13 9 1 7 9 0 13 1 9 0 0 1 12 9 1 9 9 0 1 9 7 9 0 7 9 9 2 14 7 0 1 10 9 14 13 1 9 1 9 1 9 15 2 7 13 15 13 1 9 1 9 7 9 1 9 9 7 9 15 13 1 15 2 7 15 13 9 15 1 9 1 9 1 9 9 9 15 0 2 9 1 9 9 7 9 15 13 9 15 1 9 9 9 0 0 1 9 9 2
7 9 9 9 1 9 0 0
23 13 9 0 7 9 9 9 0 1 9 0 13 1 12 8 0 9 1 12 8 9 12 2
45 7 13 9 13 15 9 0 1 9 0 7 9 7 9 9 0 1 9 9 13 1 12 8 0 7 1 9 12 8 7 1 8 12 8 7 1 9 12 8 7 1 9 12 8 2
45 7 13 9 1 9 9 9 1 9 0 9 1 9 9 0 0 2 7 13 9 9 1 9 0 9 12 1 12 8 7 1 9 12 8 7 1 9 12 8 7 1 9 12 8 2
14 9 1 2 9 2 13 8 2 15 8 6 1 9 2
53 13 9 13 15 9 1 9 2 9 0 2 1 9 0 8 8 9 1 9 1 9 9 0 1 2 9 2 1 9 7 9 15 1 9 0 2 7 9 7 13 13 1 9 9 15 1 9 9 1 9 9 15 2
33 7 13 9 1 9 15 13 15 9 2 9 2 1 9 1 9 2 1 9 0 1 9 0 2 15 13 9 0 1 9 1 9 2
7 7 15 9 9 2 2 2
17 7 15 9 0 1 9 9 7 9 9 7 9 7 9 2 2 2
10 7 15 13 9 6 1 9 2 2 2
28 7 13 9 1 9 15 1 7 2 9 0 13 2 2 0 9 2 9 2 1 2 9 7 9 9 0 2 2
118 7 13 8 1 9 15 1 9 2 2 9 13 9 1 9 15 1 9 9 7 9 2 9 1 9 0 7 9 1 9 0 7 9 1 1 9 0 2 13 1 9 9 15 7 9 15 15 13 9 15 1 9 9 2 7 1 15 9 15 1 9 0 2 9 13 3 9 1 9 9 13 9 2 7 9 9 0 9 15 9 9 1 9 7 9 2 7 9 1 1 9 13 1 9 9 7 9 9 2 8 9 7 9 2 14 13 9 8 2 7 9 0 2 7 9 0 2 2
66 7 1 9 1 9 2 9 0 2 1 9 2 13 9 7 9 0 0 1 9 9 7 9 15 9 15 9 1 9 9 1 9 9 7 9 7 9 1 9 9 0 2 9 15 13 7 13 9 0 9 13 1 9 9 7 9 1 9 9 13 9 9 7 9 2 2
121 7 13 9 7 9 15 13 1 15 9 1 9 7 9 0 7 0 0 2 13 9 9 7 9 9 2 7 9 9 0 2 7 9 9 7 13 9 1 9 2 7 9 15 13 9 9 7 9 7 13 9 7 9 2 7 9 1 9 9 7 15 9 0 1 9 2 9 7 13 1 9 10 9 1 9 7 9 7 9 1 9 9 15 1 9 7 1 9 9 15 1 9 1 9 2 7 1 9 9 1 9 1 15 9 15 7 9 15 13 9 9 7 13 9 15 7 13 9 15 2 2
29 7 13 9 2 9 2 1 9 2 8 8 7 8 8 8 15 8 1 8 9 7 1 8 9 7 1 8 9 2
35 7 1 0 9 13 2 15 15 9 9 0 15 13 15 9 0 0 1 9 15 0 1 15 2 7 9 1 9 7 9 1 9 15 2 2
7 12 12 9 0 1 9 9
54 13 9 0 13 15 9 0 1 9 7 9 9 7 9 0 1 9 1 9 12 12 9 9 0 1 9 0 15 15 1 9 1 12 1 12 9 2 7 15 13 9 15 1 12 12 9 14 13 1 15 9 1 1 2
14 7 13 9 7 9 9 0 1 9 9 15 12 5 2
58 7 13 9 7 9 9 9 9 0 13 1 7 15 1 1 12 12 9 7 9 1 9 0 10 1 12 1 12 9 14 13 1 15 1 12 12 3 2 12 5 7 13 9 1 9 0 7 15 9 0 1 9 9 0 1 9 0 2
14 7 13 9 1 9 12 9 7 9 1 12 9 0 2
37 7 13 15 13 1 15 9 1 9 9 0 1 15 2 7 13 9 9 7 9 9 7 15 13 7 0 0 10 9 7 15 13 7 13 1 9 2
46 0 15 13 15 9 15 9 1 7 9 7 9 13 9 0 1 9 9 0 2 7 15 1 9 9 1 9 9 9 2 7 13 9 1 9 9 0 1 9 1 9 0 1 10 9 2
8 9 0 1 9 8 2 0 2
58 13 8 2 8 8 8 9 9 2 9 9 13 2 13 9 9 0 1 7 9 9 0 1 9 0 2 8 8 2 14 13 9 1 9 9 0 0 1 9 9 2 9 9 0 0 2 13 9 7 9 7 9 0 1 9 9 0 2
35 7 13 10 9 1 7 9 0 14 13 9 1 1 12 12 9 2 1 9 9 9 0 7 0 2 7 3 9 9 0 0 1 9 9 2
20 7 13 9 9 1 9 2 1 9 0 7 9 0 1 9 9 9 1 9 2
41 7 1 9 1 15 2 13 8 1 9 9 1 9 0 1 8 7 9 7 1 9 9 9 0 0 1 9 9 1 9 15 13 9 0 1 9 0 0 1 9 2
33 7 13 8 7 13 9 9 0 0 10 2 9 9 1 9 0 1 9 7 9 1 9 7 9 14 13 9 9 2 1 15 0 2
40 7 13 9 9 7 9 0 13 13 7 9 1 10 13 2 9 0 0 2 7 13 9 15 13 7 13 1 9 9 0 0 1 9 1 9 2 15 9 0 2
57 7 1 9 9 2 13 9 8 7 13 9 0 8 7 13 9 1 9 0 1 8 1 9 9 2 7 7 9 1 9 2 15 13 8 13 15 0 0 0 0 2 1 9 0 7 9 9 0 2 14 13 9 1 9 1 9 2
58 7 9 1 10 9 2 13 8 7 15 1 0 9 9 0 1 9 0 2 7 7 13 0 0 2 9 1 9 9 0 1 9 0 1 9 15 9 0 2 7 13 7 15 1 9 7 9 7 9 9 13 9 8 0 1 9 0 2
69 7 13 8 1 10 9 13 9 0 1 9 0 0 9 2 1 9 2 7 9 2 7 13 7 15 14 13 10 9 1 9 1 9 7 13 15 1 8 0 7 9 9 0 0 2 7 13 1 15 2 9 2 7 13 9 9 0 0 7 14 3 8 7 8 2 2 9 0 2
91 7 1 10 9 2 7 14 9 10 2 9 9 2 0 0 2 2 15 13 1 2 9 0 2 7 9 7 8 2 7 15 14 13 1 15 9 9 7 9 0 0 2 14 13 1 9 9 2 0 2 0 2 1 9 0 1 9 2 7 9 15 15 9 9 1 9 9 2 9 14 13 0 7 0 7 0 2 0 1 8 7 8 2 9 7 9 2 7 8 0 2
111 7 7 7 14 0 9 15 9 7 9 9 0 1 10 1 9 9 9 0 0 2 7 9 9 7 9 0 0 2 0 2 7 1 0 9 9 15 1 1 2 9 0 2 2 1 9 7 9 0 14 13 9 9 0 0 1 9 2 0 2 7 0 2 7 0 7 13 10 9 1 9 0 2 0 1 9 0 13 1 15 9 1 9 0 2 2 1 9 9 0 0 2 9 9 9 7 9 2 9 0 0 7 9 15 1 9 2 9 0 2 2
41 7 1 9 2 14 9 8 0 0 15 9 9 0 7 0 0 2 0 0 2 8 1 9 9 0 2 0 1 9 2 7 9 9 1 9 9 0 7 9 0 2
26 8 8 8 8 8 9 9 2 9 9 2 1 0 2 8 8 1 9 0 7 0 7 9 0 0 2
25 7 7 10 9 13 1 9 7 9 9 0 1 0 9 9 0 1 9 9 0 2 8 8 9 2
12 8 2 9 7 9 9 1 8 1 9 9 9
34 13 0 9 0 0 3 2 7 9 0 1 9 9 9 7 7 15 13 7 9 7 9 9 9 1 9 0 15 9 0 1 9 2 2
52 7 13 9 9 7 9 0 0 8 8 1 9 1 9 2 8 8 12 8 2 7 15 14 13 1 15 7 13 9 9 9 2 14 13 8 1 9 9 9 9 9 1 9 12 9 0 1 9 0 1 9 2
18 7 13 2 8 0 1 9 9 2 8 8 8 8 3 0 9 2 2
35 7 13 0 2 8 0 1 7 3 9 1 10 9 0 8 9 9 9 1 8 2 7 9 0 1 7 15 14 13 9 1 9 9 2 2
22 7 13 8 1 9 1 15 14 13 1 15 9 8 1 12 9 2 9 2 1 8 2
16 7 13 2 14 9 13 15 9 1 0 9 1 9 0 2 2
31 7 13 2 9 9 13 8 1 9 2 2 14 8 8 7 15 9 8 8 9 0 1 9 9 0 1 9 7 9 2 2
58 7 7 13 9 8 8 8 2 7 9 14 13 1 8 9 2 2 13 8 2 14 8 15 7 13 13 9 15 2 8 8 9 1 9 9 9 1 9 9 1 9 9 2 7 13 9 1 9 13 1 15 0 9 1 9 0 2 2
11 9 9 9 0 2 0 1 9 12 12 9
44 13 9 9 7 9 0 8 8 11 8 8 3 2 1 9 9 9 1 9 2 9 0 1 9 2 1 9 12 12 9 0 2 1 9 1 9 9 0 1 9 7 1 15 2
47 7 13 1 9 13 15 9 9 0 2 7 9 15 14 13 1 9 0 7 0 14 13 0 1 9 12 1 12 1 9 9 1 9 7 12 1 12 1 9 9 0 2 8 8 8 2 2
44 7 13 2 7 9 10 9 13 9 0 1 9 1 9 9 9 7 9 1 9 1 9 9 0 7 9 9 9 1 9 0 1 9 1 9 9 9 9 9 0 1 15 0 2
20 7 13 7 9 14 13 9 15 1 9 9 0 13 9 15 1 9 9 0 2
16 9 0 2 9 9 0 14 13 0 1 9 0 1 9 12 0
34 13 9 0 0 13 0 7 9 9 14 13 1 9 1 9 9 0 1 8 8 0 3 7 13 9 9 0 1 9 9 0 1 9 2
65 7 13 9 15 13 1 0 1 12 9 7 0 1 9 9 0 7 0 15 13 9 15 1 8 1 9 2 9 9 1 9 0 2 7 15 1 9 9 0 2 8 8 2 15 13 1 9 9 2 15 7 9 1 9 9 0 13 1 9 0 1 9 9 0 2
51 7 13 9 0 9 0 1 9 0 1 9 1 9 0 7 9 8 2 7 13 9 9 9 1 9 0 1 9 1 9 0 7 9 0 2 8 8 1 7 9 13 9 0 1 9 0 1 9 9 9 2
20 7 13 9 3 9 9 9 0 0 7 8 7 8 1 9 9 0 1 9 2
55 7 13 9 1 9 9 7 9 0 9 1 9 1 9 9 9 0 7 9 8 1 10 13 1 9 9 7 9 0 7 9 15 14 13 9 9 7 13 0 1 9 0 1 9 9 8 8 9 15 1 9 1 9 9 2
31 7 13 9 3 9 9 15 13 1 9 7 1 1 15 9 15 13 1 9 9 0 1 9 7 9 2 9 9 7 9 2
20 7 13 10 9 0 9 0 7 9 0 9 8 0 1 9 8 7 9 0 2
23 7 0 13 9 9 15 13 9 9 9 9 0 7 9 8 1 9 12 7 1 9 12 2
44 7 13 9 1 10 9 1 7 9 1 9 1 9 9 9 15 0 1 9 9 9 1 9 9 0 7 9 9 1 9 9 0 1 9 0 2 7 9 9 9 1 9 9 2
37 2 9 9 9 0 2 7 13 9 1 7 15 15 14 13 9 0 0 7 9 9 0 1 9 7 14 9 1 9 9 0 14 13 1 9 9 2
85 7 13 9 7 15 1 9 9 0 1 9 15 9 15 2 8 8 2 7 9 9 1 9 9 1 0 0 15 13 9 9 0 1 9 9 9 1 9 0 2 7 1 9 9 9 9 1 9 1 9 9 0 2 14 7 9 10 9 14 13 9 15 7 13 9 0 1 9 9 0 2 7 9 9 9 0 1 9 9 9 0 7 9 8 2
36 7 1 9 2 7 1 9 12 9 13 10 9 1 9 9 0 7 9 8 9 0 1 9 9 2 7 13 1 9 1 9 1 9 10 9 2
94 7 13 9 7 9 15 13 15 9 8 8 2 8 8 2 13 1 10 9 1 9 0 2 7 13 9 9 0 1 9 12 1 12 12 9 1 9 0 2 13 9 9 9 0 7 9 8 1 15 12 12 9 7 15 13 12 5 2 7 13 10 9 9 12 7 13 1 12 12 9 1 9 0 2 14 7 9 9 0 7 9 8 13 15 0 7 13 12 5 7 12 12 9 2
49 7 13 10 9 9 0 9 12 7 13 1 12 2 12 12 9 1 9 2 7 9 0 13 9 9 9 0 7 9 8 7 13 1 12 12 9 1 9 0 7 15 13 12 5 1 9 9 0 2
52 7 1 9 9 12 13 9 9 0 1 9 12 2 12 8 9 1 9 0 2 14 7 0 7 9 9 0 7 9 8 13 1 12 5 7 15 13 12 8 9 1 9 9 1 9 15 13 15 9 8 8 2
78 7 13 9 9 9 0 7 13 9 9 9 8 0 1 7 13 9 9 0 1 9 9 1 9 12 5 2 7 9 9 9 9 0 15 13 1 7 13 9 1 9 1 12 12 9 1 9 0 9 12 7 13 1 12 12 9 0 1 9 9 12 7 1 0 7 13 9 15 1 9 9 0 9 1 9 8 3 2
51 7 9 0 15 13 15 9 15 9 15 1 7 9 14 13 9 0 1 8 9 0 13 1 10 9 2 7 7 14 3 0 1 9 15 13 9 9 9 0 1 9 8 1 9 9 0 1 8 8 0 2
97 7 13 9 3 1 7 9 9 0 7 9 8 14 13 9 0 1 9 9 0 1 9 9 1 9 0 7 0 2 0 15 7 15 13 9 0 2 7 7 9 15 13 2 7 9 0 1 9 0 1 9 7 1 9 14 13 2 3 7 14 9 9 13 0 0 0 1 9 9 9 0 2 15 1 9 1 7 9 0 7 0 14 13 9 0 1 9 0 2 7 13 9 0 1 9 9 2
18 9 9 0 2 14 13 0 1 9 8 9 9 0 1 9 1 9 9
77 13 9 8 11 8 11 8 8 9 9 0 9 9 0 1 9 9 0 1 9 1 9 2 9 9 7 9 2 1 9 0 2 7 7 13 9 9 0 1 9 8 1 9 0 2 0 1 7 9 0 1 8 0 0 1 9 9 1 9 15 13 9 15 1 9 0 2 7 13 9 0 1 0 1 9 0 2
147 7 13 9 8 11 8 8 9 9 7 9 0 1 9 1 9 3 1 9 15 1 9 9 9 9 0 9 9 7 9 14 13 1 1 9 9 15 14 13 1 15 9 0 1 9 9 0 1 9 2 8 2 7 0 9 15 1 12 1 9 9 2 9 2 2 7 13 7 9 9 14 13 15 9 7 14 9 8 2 7 7 9 1 0 1 9 0 1 9 1 15 9 1 9 9 1 9 2 8 8 8 9 9 1 8 9 9 1 1 9 8 9 2 8 8 1 8 7 9 0 1 9 7 9 15 1 9 12 9 1 9 2 7 7 13 9 9 10 1 12 2 12 9 1 9 0 2
24 7 13 7 9 13 15 12 9 0 15 9 9 2 7 7 9 0 15 1 12 9 8 8 2
76 7 1 9 9 0 1 9 9 8 13 8 7 1 0 9 1 9 1 10 14 13 9 1 15 1 9 9 2 7 9 15 13 9 0 1 9 15 13 1 15 9 2 7 1 0 1 9 0 7 3 9 1 9 2 7 13 9 0 0 2 1 1 9 15 13 9 15 1 9 1 9 1 9 9 8 2
15 7 13 8 7 9 1 9 15 9 9 0 1 9 15 2
55 7 1 9 9 9 0 9 1 9 9 9 1 9 0 0 7 13 9 0 1 9 12 9 2 13 9 7 10 9 14 13 1 9 0 1 9 9 1 8 2 7 7 15 14 13 9 15 15 14 13 1 9 9 9 2
35 7 13 8 7 9 9 0 1 9 1 9 9 7 9 1 9 9 9 2 7 13 7 15 1 9 9 9 14 13 9 1 9 9 9 2
115 7 1 0 1 9 9 9 9 13 9 8 7 9 1 9 9 9 13 9 9 9 1 9 2 7 7 15 1 9 9 9 9 15 14 13 8 9 0 1 9 0 1 9 8 8 7 14 9 15 1 9 0 14 13 0 7 9 9 1 0 9 2 7 13 7 9 0 15 9 9 9 1 9 0 1 9 1 9 0 2 7 13 9 1 9 9 9 0 2 7 3 9 1 9 9 9 9 7 13 0 9 15 14 13 9 15 1 9 0 7 13 15 9 0 2
43 7 1 9 13 15 8 1 9 9 9 13 7 9 9 0 1 9 9 15 9 9 9 1 9 9 0 1 9 9 7 9 8 1 9 7 9 9 0 14 13 9 0 2
32 7 13 9 8 9 9 9 0 0 1 9 0 1 9 7 15 9 0 2 7 0 9 2 7 9 8 2 8 2 7 9 2
43 7 13 7 9 0 1 9 0 13 12 1 12 1 0 9 1 9 2 7 13 9 9 1 10 9 12 12 9 2 7 13 9 0 1 9 1 9 12 1 12 12 9 2
50 7 1 9 15 13 8 8 8 9 9 9 9 0 7 9 9 0 1 9 9 0 7 0 1 9 0 0 1 9 9 2 0 7 3 9 1 9 1 10 9 1 9 9 7 9 9 1 9 0 2
14 2 8 2 0 0 9 0 13 9 9 0 1 8 9
36 13 9 1 9 0 3 2 7 9 8 0 13 9 9 9 0 1 9 8 9 0 7 13 0 9 0 13 9 1 0 9 0 1 9 2 2
25 7 13 9 1 9 0 1 9 2 13 9 9 8 8 15 13 9 15 12 9 1 8 9 2 2
26 8 8 15 0 9 3 13 9 15 1 8 9 1 7 8 0 1 9 9 1 9 8 9 0 0 2
16 7 13 9 9 9 0 1 9 9 1 9 9 9 1 9 2
31 7 1 9 14 13 1 8 0 9 1 8 9 1 9 13 9 0 2 7 0 7 15 14 13 8 1 9 0 1 9 2
34 7 13 9 9 9 8 8 8 9 1 0 9 2 9 2 0 0 9 9 1 10 1 12 12 7 12 12 9 1 9 1 9 9 2
20 7 1 9 12 0 9 15 13 1 9 15 13 0 9 12 12 9 1 9 2
15 7 13 12 9 3 9 9 7 9 15 1 9 9 0 2
25 7 13 8 8 9 9 0 1 12 9 1 9 9 0 1 9 1 9 0 13 1 15 1 9 2
28 7 13 9 1 9 12 9 1 9 1 9 9 0 15 13 1 9 0 13 1 12 7 12 12 9 1 9 2
36 7 13 9 9 7 9 8 9 1 9 9 9 0 1 9 9 7 13 9 7 15 13 9 0 1 9 1 9 1 12 12 9 1 9 9 2
37 7 13 9 1 9 9 9 1 9 9 1 9 0 1 9 9 0 14 7 9 0 13 7 9 14 13 9 9 8 9 1 9 15 0 1 9 2
17 7 13 9 1 9 9 0 2 13 7 15 4 1 15 9 9 2
13 9 9 9 13 9 0 7 15 14 13 9 9 0
43 13 9 9 9 7 9 0 1 15 1 9 9 0 0 13 9 9 9 0 1 15 9 9 15 0 1 9 1 9 9 0 7 1 9 9 15 0 1 9 7 9 0 2
33 7 13 10 9 13 9 0 1 9 9 0 0 15 13 0 9 1 9 1 9 0 7 9 9 7 9 0 1 9 9 9 9 2
18 7 13 9 9 1 9 0 0 1 7 13 9 1 9 0 1 9 2
29 7 13 0 9 1 9 1 10 9 2 9 8 8 8 8 13 1 15 8 8 9 0 13 12 9 9 9 0 2
24 7 9 1 9 13 1 9 9 0 9 1 9 1 10 9 7 9 15 1 9 1 9 0 2
32 7 13 9 0 1 9 9 0 0 8 8 1 9 9 9 9 0 1 9 9 10 9 7 9 9 0 0 0 1 9 9 2
72 7 1 9 14 13 9 9 0 2 14 7 9 9 9 2 7 9 9 1 9 9 1 9 9 9 2 1 9 1 9 9 0 1 9 15 13 9 9 1 7 9 15 13 1 0 1 12 12 2 12 12 12 2 9 2 9 9 15 13 9 1 7 13 10 9 1 9 9 15 1 0 2
58 2 9 9 9 0 1 9 2 13 9 0 1 9 0 0 1 9 7 9 1 15 1 9 9 2 7 15 13 0 9 0 1 9 1 9 7 9 15 1 9 9 0 0 14 13 12 1 12 2 7 15 3 0 9 9 1 9 2
38 7 1 1 9 0 0 0 0 7 14 9 0 13 15 13 9 9 9 9 1 9 0 2 7 10 9 14 13 1 15 0 9 0 1 8 8 0 2
49 7 13 9 0 1 9 9 3 2 0 2 9 9 15 1 9 1 9 7 9 13 9 7 9 0 0 2 7 0 2 9 9 9 9 15 1 9 1 9 9 2 8 2 7 9 9 1 9 2
38 7 9 1 10 9 13 9 9 0 1 9 9 9 9 2 7 7 13 9 0 9 0 9 9 1 9 15 13 0 9 15 1 9 9 8 8 0 2
43 7 13 9 9 9 1 12 9 7 0 1 12 8 2 7 13 9 9 15 1 12 9 2 7 13 1 9 8 9 8 7 8 2 9 1 9 8 0 0 1 9 0 2
14 7 14 13 9 10 9 0 0 1 12 12 9 0 2
51 2 9 9 9 2 13 9 9 1 9 9 7 9 9 9 9 1 9 9 14 13 0 2 7 15 1 9 0 1 15 2 7 9 9 0 1 9 13 0 7 15 14 13 12 1 12 1 9 9 0 2
45 7 13 9 9 9 0 0 1 12 9 9 0 2 7 9 1 9 9 9 0 7 14 9 10 9 13 7 13 9 15 1 1 12 7 12 12 9 0 7 15 1 9 9 12 2
136 0 7 1 10 9 14 9 7 13 9 0 1 9 9 0 2 7 9 10 9 14 13 1 0 9 1 9 7 13 9 9 2 7 9 0 1 9 15 13 1 9 9 0 0 1 12 12 9 0 2 7 0 1 9 10 9 13 1 9 1 9 15 2 7 13 9 9 2 8 2 1 9 9 15 0 1 12 12 9 0 2 7 9 2 8 2 0 13 1 12 9 9 9 9 1 9 12 2 14 1 9 9 7 14 9 13 9 0 13 1 12 7 12 12 9 2 15 1 9 1 0 1 12 12 9 1 9 0 14 13 9 0 1 10 9 2
78 1 9 7 9 9 9 0 13 9 9 9 0 0 7 15 13 0 9 1 9 9 7 14 13 9 9 9 0 0 1 9 2 1 9 14 13 1 12 9 1 9 0 1 9 9 2 2 15 1 9 1 7 15 0 1 9 0 2 7 1 1 15 9 7 9 7 3 9 2 15 13 9 15 0 9 1 0 2
49 13 3 7 9 1 9 1 0 7 13 1 0 1 12 12 9 0 0 1 1 12 12 9 0 7 15 1 9 9 12 2 7 1 0 7 13 9 15 1 9 9 0 9 1 9 2 8 2 2
13 9 2 8 13 0 9 9 1 9 9 1 9 0
38 13 9 0 1 9 9 0 1 8 0 9 9 1 9 9 1 9 9 7 9 7 9 0 1 10 9 0 1 9 1 0 7 13 1 15 9 0 2
32 7 13 9 1 9 2 7 9 0 8 8 15 13 9 9 15 1 9 7 9 13 7 1 9 0 8 0 1 9 0 2 2
24 7 13 8 8 1 9 9 1 9 8 1 9 2 8 13 7 9 0 1 9 15 8 2 2
12 7 14 13 9 1 9 0 1 9 0 2 2
32 7 13 8 15 13 1 9 13 9 9 12 1 9 9 9 0 2 14 3 0 1 9 9 1 9 9 7 9 1 9 0 2
20 7 15 13 2 9 0 15 9 0 1 9 7 9 0 15 13 9 0 2 2
44 7 1 9 0 13 9 0 7 9 15 13 1 9 9 9 1 9 12 7 13 9 9 8 8 9 1 8 13 15 9 9 1 9 1 10 9 1 9 0 1 9 9 9 2
40 7 13 9 1 9 2 7 8 8 2 8 8 2 8 8 2 7 15 9 0 1 8 8 2 7 8 8 2 13 9 1 9 9 0 0 1 9 9 2 2
16 7 13 9 0 7 8 0 1 9 9 7 9 9 9 0 2
48 7 13 8 8 9 9 8 8 0 1 9 9 0 1 9 9 8 8 13 9 9 9 0 1 9 9 8 8 2 9 9 0 1 9 0 15 13 8 7 15 13 1 9 7 9 2 2 2
11 15 15 13 8 0 1 9 1 9 2 2
23 7 1 15 13 8 2 7 9 0 13 15 9 1 9 7 7 9 0 14 13 0 2 2
29 7 13 9 8 8 9 0 1 8 1 9 1 9 9 7 13 1 0 7 13 15 1 9 2 9 0 2 0 2
16 7 13 8 1 9 0 0 1 8 1 13 9 15 1 9 2
18 8 1 9 9 0 1 9 1 0 9 14 13 8 1 9 1 8 2
22 7 13 8 9 15 1 8 9 1 9 9 0 1 9 15 13 1 9 9 9 0 2
28 7 13 9 8 8 8 0 7 9 0 8 8 13 9 9 9 7 9 1 9 9 7 9 9 8 1 9 2
17 2 8 2 0 13 1 9 9 9 1 9 1 9 9 9 1 9
41 13 9 9 0 7 9 9 0 7 9 8 2 8 2 0 3 1 9 9 9 1 9 9 0 1 9 9 9 9 0 1 9 1 9 9 15 13 15 9 0 2
34 7 13 9 15 13 12 8 9 1 9 2 9 9 8 8 7 9 0 1 9 8 8 1 9 9 9 7 9 0 0 9 8 8 2
68 7 1 9 9 14 13 9 9 1 9 1 9 1 9 0 1 9 1 9 9 1 9 9 9 9 1 9 7 9 7 9 1 9 9 9 7 9 9 1 7 1 9 9 7 9 9 1 9 9 2 7 13 9 1 9 1 9 15 13 1 15 9 9 9 0 1 9 2
46 7 13 9 1 9 1 9 9 1 9 7 9 9 15 0 1 9 12 1 12 1 9 9 0 1 9 2 1 1 7 9 9 0 0 1 9 9 0 1 9 1 9 9 9 0 2
59 7 13 9 9 1 9 13 15 9 9 0 7 9 1 9 13 8 0 1 9 0 0 13 1 15 9 9 0 9 1 9 9 0 0 0 2 0 1 7 9 1 9 15 9 0 1 9 9 0 14 13 9 15 1 9 9 1 0 2
37 7 13 9 8 7 10 9 1 9 15 0 13 1 0 9 9 0 7 13 1 9 9 1 9 0 1 9 12 9 1 9 13 1 12 12 9 2
24 9 2 9 2 8 2 0 1 9 12 12 9 1 9 9 15 0 1 12 12 9 1 9 12
72 13 9 0 9 9 9 1 9 9 0 1 9 2 8 2 1 12 1 12 1 9 0 1 9 9 12 7 1 12 1 12 1 9 0 9 12 7 15 9 9 0 1 9 0 1 1 8 1 9 9 0 1 9 1 9 1 9 15 13 1 15 9 0 1 9 9 0 1 9 9 8 2
67 7 13 9 15 13 15 9 9 0 1 9 1 9 9 0 7 9 9 0 0 1 9 8 1 9 13 1 12 12 9 1 9 9 0 1 1 12 12 9 0 1 12 2 0 1 7 9 9 0 1 12 12 9 1 9 0 0 0 1 9 9 0 13 12 12 9 2
55 7 13 9 15 13 9 9 2 8 2 7 2 8 2 1 9 9 7 9 9 1 9 14 13 9 0 1 9 9 0 1 9 2 0 7 10 9 13 1 12 1 12 1 9 0 0 1 9 7 13 1 9 9 9 2
94 7 13 9 7 9 9 8 7 8 1 9 1 9 0 7 0 1 9 9 0 1 9 9 15 13 9 9 1 9 15 1 9 9 0 8 1 9 0 7 0 2 7 3 9 9 9 0 2 13 1 9 9 7 9 0 9 9 9 0 1 9 9 0 1 9 13 1 8 8 7 12 0 1 9 13 8 1 9 9 7 13 1 9 9 15 1 9 9 0 1 10 9 0 2
48 7 13 9 9 9 1 9 1 9 0 2 0 7 15 9 0 1 9 1 9 9 0 1 9 1 9 0 7 13 9 0 1 9 15 1 9 0 9 9 0 13 7 13 1 9 0 0 2
59 7 13 9 1 9 9 9 0 1 10 13 9 7 9 9 0 1 9 9 1 9 1 2 8 2 7 2 8 2 7 3 9 9 9 0 1 9 9 9 9 7 9 9 1 9 9 0 7 13 1 9 9 9 7 9 1 9 9 2
83 7 13 9 1 9 0 9 1 9 13 1 9 9 9 0 7 9 9 9 7 9 1 9 0 13 15 9 9 2 0 1 9 9 9 9 9 9 1 9 8 7 8 1 9 0 1 9 1 9 0 1 9 9 7 9 7 9 2 7 13 9 9 1 9 0 15 13 1 8 7 8 0 15 1 9 0 2 1 9 15 9 0 2
13 9 0 2 9 9 9 0 1 9 9 9 2 2
6 7 14 13 2 8 2
27 13 9 1 9 0 1 3 1 9 0 1 9 9 1 9 0 1 9 0 0 0 7 9 9 9 0 2
36 7 13 8 8 9 9 0 1 9 8 8 9 9 0 1 9 9 2 8 2 0 2 2 14 9 0 1 9 0 7 9 1 15 0 2 2
37 7 13 1 9 1 9 2 9 0 2 1 9 2 8 2 8 2 8 2 2 2 1 9 9 13 9 0 7 15 15 9 1 9 8 9 2 2
22 7 13 8 9 9 1 9 9 8 9 1 8 7 15 9 9 0 1 9 9 9 2
15 7 13 2 14 13 9 0 1 8 1 12 9 0 2 2
25 7 1 7 7 7 13 9 0 1 9 0 7 7 14 13 9 15 7 14 13 15 1 9 2 2
40 7 13 8 3 2 2 14 1 0 1 9 9 0 7 9 0 9 9 1 9 0 7 9 0 0 13 9 9 0 1 9 1 9 9 0 1 9 9 2 2
28 7 1 9 9 13 9 1 7 9 9 1 8 1 9 8 14 13 15 9 9 1 9 8 7 9 9 0 2
33 7 13 8 2 2 15 14 13 9 0 1 9 10 9 7 15 14 13 9 0 9 1 9 9 14 13 3 0 9 1 9 2 2
7 14 13 9 9 9 2 2
5 1 9 9 0 2
34 1 10 9 13 9 2 9 2 9 0 13 1 15 2 15 13 9 9 1 9 15 13 15 9 7 9 1 9 0 1 9 9 0 2
41 9 13 15 9 1 9 13 1 15 9 1 9 0 0 13 1 9 0 14 13 15 9 0 7 9 1 9 9 9 0 1 15 1 15 9 1 9 0 8 8 2
31 2 2 9 0 14 13 9 9 9 9 0 0 1 9 9 15 7 13 1 9 7 13 7 13 9 1 15 1 8 9 2
44 14 9 9 15 13 15 9 0 1 9 0 13 9 13 9 9 1 7 9 8 13 13 9 1 9 0 1 9 14 13 15 15 9 7 13 9 9 15 14 13 9 10 9 2
80 7 14 14 0 10 1 9 0 15 7 9 9 0 8 8 1 9 1 9 8 7 15 13 9 15 1 15 2 7 14 9 0 13 7 15 13 13 9 1 9 0 7 0 1 10 9 4 3 1 9 0 1 8 1 8 7 3 1 9 0 13 1 8 7 1 9 9 7 9 0 7 9 0 1 9 1 9 9 0 2
88 7 13 9 9 1 9 9 9 9 7 9 9 9 0 8 8 1 9 9 9 7 9 1 9 9 7 13 8 1 9 9 9 0 1 9 9 10 9 1 7 15 14 13 9 9 9 8 8 2 7 0 9 14 13 1 9 13 9 7 10 9 14 13 9 0 7 14 13 8 9 9 9 0 8 8 7 9 9 9 12 9 0 14 13 1 9 9 2
7 7 7 15 9 2 2 2
58 0 7 9 13 7 13 9 9 9 0 7 9 15 1 9 0 1 9 9 0 15 13 9 9 0 7 15 14 13 7 7 1 9 7 13 1 10 9 0 15 13 15 9 9 0 1 7 15 13 9 0 1 9 1 9 9 0 2
20 2 2 9 0 14 3 9 0 9 1 9 1 9 10 9 9 1 9 0 2
47 12 2 14 9 0 13 1 9 14 13 1 15 9 9 1 0 9 9 1 0 9 9 1 9 9 9 1 8 7 9 7 3 1 9 3 7 9 7 14 1 9 9 0 1 9 0 2
45 12 2 14 9 9 9 13 9 9 0 1 9 1 9 9 15 13 1 15 4 1 9 9 0 7 9 0 7 14 1 9 9 0 0 1 9 0 14 13 13 9 9 1 9 2
69 12 2 14 9 10 13 1 9 13 9 9 1 9 9 0 1 9 0 1 9 9 1 9 7 15 15 14 13 9 0 1 8 8 1 9 10 9 1 9 0 0 1 9 9 0 7 9 9 15 13 15 1 9 9 0 7 13 8 8 7 13 7 13 15 9 7 9 9 2
53 12 2 14 9 14 13 1 9 9 0 1 9 9 0 7 9 0 9 0 7 13 9 9 9 0 1 9 0 7 1 9 7 1 9 1 9 7 9 9 0 9 1 9 9 7 9 0 7 9 15 1 9 2
59 12 2 14 9 0 0 14 13 0 9 1 9 9 9 14 13 15 1 8 15 14 13 9 1 0 9 1 9 9 1 9 1 10 9 7 9 0 15 13 9 0 8 8 9 15 13 1 10 9 0 1 9 7 13 9 9 0 0 2
70 12 2 14 9 13 7 13 9 1 10 9 1 9 9 9 1 9 15 0 7 3 1 9 9 0 0 1 9 9 0 1 9 1 9 0 9 0 1 9 9 13 1 15 9 7 15 13 9 1 9 0 15 13 15 0 1 9 9 15 2 2 9 0 1 15 13 9 7 15 2
112 14 0 1 9 13 7 9 0 1 0 9 14 13 1 9 8 0 8 8 7 7 13 1 9 0 7 1 9 9 13 9 15 13 1 15 9 0 1 9 7 13 1 9 9 8 0 9 7 1 9 0 7 13 8 0 1 9 0 9 1 9 9 1 0 9 0 7 9 9 1 0 1 9 9 10 9 1 9 13 0 9 0 1 15 1 7 9 8 7 2 9 9 2 9 1 10 13 1 9 15 13 1 15 9 7 1 15 8 1 9 9 2
51 2 2 9 9 14 9 15 13 9 9 15 13 15 1 9 9 13 1 9 1 8 13 1 15 1 9 9 7 13 7 1 0 9 7 13 7 8 8 14 13 9 0 1 9 8 1 7 13 9 0 2
32 14 10 9 9 0 2 7 14 3 15 13 15 1 9 9 9 7 1 7 1 9 9 0 1 9 0 1 9 0 8 8 2
34 7 3 7 9 13 1 9 9 1 9 9 1 1 10 9 0 7 7 15 13 13 9 7 15 13 9 1 9 9 1 15 1 9 2
15 2 2 9 0 15 15 9 0 0 2 7 9 0 3 2
65 14 15 13 1 9 9 8 1 9 8 9 7 13 9 10 13 15 9 1 9 9 7 15 13 1 9 9 9 9 7 3 1 9 9 1 9 7 0 1 9 9 8 15 13 7 13 9 1 9 15 0 1 9 0 7 15 13 9 1 9 13 9 0 9 2
140 7 1 9 1 7 9 13 9 9 15 1 8 1 7 15 9 9 0 7 13 7 8 14 13 0 1 0 9 0 7 14 3 15 13 1 7 14 9 0 1 9 1 9 9 1 0 9 0 1 9 9 0 7 15 15 13 7 8 14 13 9 10 1 15 1 9 1 15 13 9 0 9 14 13 15 9 0 1 9 0 7 9 9 9 9 0 9 1 9 9 9 15 14 13 10 9 1 9 9 9 0 7 15 13 9 9 0 1 9 9 0 1 9 0 1 9 14 13 1 9 12 8 1 9 10 13 2 9 9 2 1 9 7 9 2 9 9 2 3 2
77 7 1 9 13 1 10 9 7 14 9 14 13 9 9 0 1 2 9 9 2 1 15 13 9 9 9 0 1 9 1 9 9 7 9 9 1 9 0 9 1 15 1 15 9 0 1 9 7 1 7 9 9 9 1 9 9 0 9 0 1 15 13 7 9 14 13 1 9 8 0 1 9 13 1 10 9 2
37 14 9 9 9 0 13 9 1 9 0 1 9 9 9 1 8 7 1 9 9 9 0 14 13 1 9 9 9 13 9 1 9 1 9 1 9 2
80 7 7 9 15 13 0 1 1 10 9 13 13 1 15 9 1 9 9 0 1 9 0 7 13 9 9 1 10 9 15 9 0 0 1 9 7 7 9 14 13 9 1 1 10 9 7 15 13 9 0 1 9 9 7 7 15 13 9 0 0 1 9 9 7 9 9 1 9 0 1 7 13 3 9 0 1 1 10 9 2
10 9 9 0 13 9 9 1 15 1 9
30 13 9 0 1 9 9 12 2 12 0 7 1 0 9 15 13 15 9 0 2 9 1 9 9 7 9 1 9 0 2
24 7 1 0 7 13 9 0 2 0 9 1 9 1 9 0 0 1 2 9 9 10 9 2 2
61 7 13 9 0 1 2 9 9 0 2 8 8 2 1 2 9 2 7 9 9 0 13 9 9 1 15 1 9 1 9 2 9 0 1 9 0 2 2 0 1 7 9 10 9 2 14 13 1 9 9 7 9 15 1 9 9 0 1 9 2 2
57 7 13 7 8 0 2 8 9 2 1 9 9 15 13 15 9 0 1 9 2 9 8 8 2 14 3 7 7 9 13 1 9 0 7 0 9 9 9 1 9 12 9 1 9 15 1 9 9 15 13 1 15 1 9 15 0 2
31 7 13 1 7 9 9 0 7 0 1 9 9 0 1 9 1 9 9 0 2 2 1 9 9 9 7 9 9 9 2 2
37 7 13 8 7 9 0 1 9 0 7 0 12 12 9 2 1 9 9 9 15 13 15 9 9 0 0 1 8 2 14 13 1 9 1 9 0 2
27 7 13 1 7 9 9 0 13 1 9 9 1 12 9 7 13 9 0 1 9 1 9 0 0 1 9 2
45 7 13 2 1 9 0 2 7 2 9 9 0 2 13 9 1 9 0 0 1 9 9 2 9 1 0 7 9 7 9 9 0 2 0 1 9 9 1 10 9 1 9 10 9 2
31 7 13 7 3 12 9 0 0 2 13 9 15 1 9 2 7 7 15 13 12 9 1 9 1 9 9 9 0 7 0 2
19 7 13 7 9 0 9 1 9 1 9 0 0 1 9 9 9 0 0 2
24 7 15 13 7 9 0 1 8 7 8 7 8 0 1 9 9 7 9 9 1 9 9 0 2
16 9 9 0 13 1 8 9 1 9 9 0 0 1 9 7 9
65 13 9 12 2 12 0 9 9 0 8 8 1 9 0 1 7 13 9 0 1 9 0 9 0 1 9 7 9 1 9 15 2 1 9 9 0 7 1 9 1 9 0 13 7 13 9 8 2 7 13 7 8 13 1 9 7 13 9 0 13 9 1 9 2 2
151 7 13 8 1 9 0 1 9 9 1 9 8 9 8 8 8 8 1 10 13 15 9 2 8 8 2 1 8 9 9 0 1 9 9 1 9 2 8 2 1 9 1 9 12 9 3 1 9 0 2 0 2 2 9 1 15 13 9 8 8 0 1 9 1 9 9 10 9 2 7 13 7 9 9 0 0 8 8 13 9 15 1 9 1 9 9 0 1 9 0 9 0 1 9 15 1 9 9 1 9 8 1 9 12 8 2 7 7 10 9 14 13 0 0 7 9 0 9 15 1 15 13 1 9 9 0 1 9 9 2 7 1 0 7 13 9 9 1 15 9 1 12 1 7 13 9 9 9 12 2 2
8 9 9 9 13 1 9 8 8
20 13 9 0 1 9 9 9 1 9 9 1 9 9 9 9 1 9 9 9 2
51 7 13 9 9 9 1 9 15 1 10 7 13 1 9 9 1 9 9 13 1 15 7 9 9 13 1 9 0 7 0 7 13 1 9 1 10 14 7 9 9 13 10 9 7 14 13 9 1 10 9 2
50 13 9 1 9 9 9 7 9 9 7 9 1 9 14 13 9 15 1 9 9 9 1 9 9 0 1 9 9 7 1 8 13 1 9 9 9 0 1 9 1 9 9 1 9 9 1 9 9 0 2
53 7 13 9 9 9 0 1 9 15 13 9 15 1 9 9 7 15 7 13 7 13 9 9 9 15 1 9 0 7 15 9 9 9 1 9 7 3 0 1 9 0 15 14 13 9 9 1 15 1 9 0 9 2
52 7 13 9 9 9 1 9 10 13 1 7 10 9 13 0 1 9 1 0 1 9 9 0 7 7 9 9 15 1 9 14 13 1 15 7 13 9 1 9 1 9 1 0 0 7 13 9 9 1 9 15 2
24 7 13 9 9 9 1 8 9 10 13 3 1 7 9 14 13 8 13 1 12 1 9 9 2
8 9 2 8 2 2 9 13 9
43 13 9 0 1 9 1 9 9 1 9 9 0 8 8 2 8 8 2 7 0 8 8 2 7 9 1 9 1 9 9 9 1 9 9 1 9 0 1 9 9 0 0 2
49 7 9 9 0 1 9 1 9 10 9 7 9 1 9 2 7 14 9 0 13 7 13 9 8 8 2 8 2 1 9 1 9 0 1 9 0 7 9 0 1 9 0 1 9 9 9 1 9 2
59 7 13 9 0 1 9 9 15 0 9 8 8 2 9 15 1 9 1 1 10 9 1 9 13 15 8 1 9 9 0 0 2 8 2 8 8 1 9 0 1 9 15 1 9 0 8 8 8 8 8 1 8 9 9 12 2 12 0 2
42 7 1 9 0 7 0 7 14 9 13 0 2 7 7 8 13 9 8 1 9 9 1 9 9 1 9 2 8 8 1 9 1 9 1 7 15 0 1 9 9 9 2
32 7 13 7 13 9 1 9 9 9 8 8 9 8 2 1 9 9 1 9 0 1 9 9 1 9 1 9 9 9 9 9 2
33 9 7 9 0 8 14 13 1 9 9 9 9 0 7 9 1 8 8 8 7 15 1 9 8 2 1 9 1 2 9 0 2 2
51 7 13 8 1 9 9 0 2 9 0 1 0 0 2 7 13 2 13 7 14 8 1 9 2 7 15 9 0 1 9 1 10 9 2 7 13 1 15 9 0 1 9 0 1 9 1 9 8 8 0 2
6 9 9 1 9 9 0
45 13 9 9 9 8 1 9 9 9 9 0 8 8 1 9 2 8 2 0 9 12 2 12 0 1 7 15 13 1 9 9 1 9 9 13 9 9 7 13 1 8 8 8 0 2
18 7 13 8 8 8 9 9 9 9 7 9 9 9 7 9 1 15 2
53 2 10 9 0 2 7 14 13 7 13 1 9 9 3 1 9 9 15 2 7 15 13 1 9 0 1 9 9 9 0 7 9 0 1 9 9 2 1 9 9 9 9 0 1 9 15 14 13 9 1 9 15 2
31 7 13 8 14 13 7 15 13 1 9 9 9 1 9 9 1 9 9 1 9 8 9 9 0 7 9 8 1 9 9 2
49 7 13 1 7 9 0 15 13 1 8 0 1 9 7 0 1 9 0 1 8 7 9 0 13 9 1 9 9 8 13 15 1 9 9 1 8 7 9 1 9 7 13 9 0 1 9 1 9 2
65 7 8 13 7 9 0 2 1 9 10 9 2 13 7 9 8 14 13 1 9 8 1 9 0 2 7 13 1 9 9 9 1 9 0 7 13 9 15 9 0 1 9 8 1 9 2 1 9 1 9 15 0 7 13 1 9 9 9 9 7 9 9 8 9 2
35 7 13 2 2 10 9 13 1 9 0 13 1 9 9 9 1 9 9 7 15 13 1 12 12 8 2 7 9 0 9 0 1 10 9 2
13 12 9 7 12 9 9 7 9 1 9 1 9 0
46 13 9 9 9 0 9 0 1 9 9 1 9 1 9 15 13 9 7 9 9 15 1 15 1 9 0 0 2 1 9 9 9 1 9 9 9 0 2 7 9 9 9 9 1 9 2
36 7 13 9 0 2 2 14 13 1 9 9 9 1 9 9 0 1 9 1 9 15 2 9 9 0 9 1 9 1 9 9 1 9 9 2 2
38 7 13 9 0 15 13 15 9 0 1 9 1 9 9 9 7 0 1 9 12 9 1 9 9 8 8 2 7 9 15 8 8 7 9 15 1 9 2
19 7 13 9 3 0 1 12 9 9 7 9 13 9 7 9 9 7 9 2
7 12 12 9 1 9 0 0
39 13 9 0 1 9 9 9 1 15 1 9 9 9 0 1 9 12 5 1 9 9 0 2 7 13 15 1 9 9 9 9 1 9 0 1 12 9 2 2
27 7 13 9 9 0 9 1 10 9 12 12 9 1 0 2 7 12 8 1 0 7 12 12 9 1 0 2
18 7 13 0 9 1 9 9 7 9 9 1 9 9 9 1 9 9 2
9 8 2 8 14 13 1 2 9 2
23 13 9 9 9 9 0 1 9 0 7 13 9 1 9 9 0 2 13 9 1 9 0 2
25 7 13 7 9 8 8 2 14 13 9 0 7 0 9 0 7 13 10 9 1 9 9 7 9 2
23 7 13 1 7 8 2 13 2 1 9 9 9 9 1 9 0 7 13 9 9 0 2 2
110 7 13 8 1 9 0 1 9 9 7 2 9 13 1 15 9 1 9 7 1 9 1 9 15 2 7 14 13 8 1 0 2 7 14 13 1 9 9 12 2 7 14 13 8 9 9 8 1 9 9 2 0 1 2 7 9 13 1 15 7 1 9 0 2 9 0 2 9 2 7 9 9 7 9 13 7 13 1 9 7 9 2 7 9 1 9 8 8 0 2 7 1 10 9 14 13 9 8 1 9 15 7 7 15 0 1 9 9 0 2
9 8 7 9 13 1 9 9 1 9
43 13 7 9 0 0 9 1 15 9 9 9 8 8 13 1 0 9 1 9 9 0 1 9 2 9 0 2 13 0 2 8 8 1 9 0 0 13 1 15 2 9 2 2
43 7 13 0 7 10 9 13 1 9 1 9 9 1 9 0 1 9 13 15 2 9 2 0 2 13 1 15 1 9 1 9 9 15 13 1 15 2 1 9 9 1 15 2
38 7 14 13 0 9 15 13 15 8 7 9 15 1 9 9 2 9 9 2 1 2 9 2 8 8 13 1 9 9 0 15 13 15 9 0 1 9 2
34 7 9 13 9 15 1 1 9 0 1 9 0 2 7 13 9 1 9 1 9 1 9 15 13 1 15 9 0 1 2 9 0 2 2
25 7 0 7 9 0 13 1 9 9 2 9 2 9 9 9 0 7 9 9 9 15 13 1 15 2
51 7 13 9 1 2 9 2 7 15 9 1 9 8 2 13 9 8 0 9 1 9 9 9 9 8 8 8 7 9 9 9 7 9 9 9 8 8 7 9 9 9 8 8 2 7 9 9 9 9 9 8
9 9 0 13 12 9 0 1 9 9
37 13 9 9 0 1 9 9 12 2 12 0 1 9 9 12 9 1 0 1 9 0 1 9 9 1 9 9 9 9 15 14 13 9 9 1 9 2
52 7 13 9 1 9 9 0 1 9 9 1 9 12 9 1 9 1 9 1 1 9 9 1 9 9 7 13 9 9 1 9 9 0 1 9 2 7 7 13 9 1 9 7 13 9 15 9 12 5 12 0 2
6 9 9 9 1 9 0
45 13 12 1 9 0 1 9 9 0 0 2 1 9 0 9 7 9 0 1 9 0 2 0 1 9 9 2 9 1 9 9 9 1 9 1 9 0 15 13 9 12 2 12 0 2
39 7 13 9 9 1 9 9 9 9 0 1 9 9 9 2 1 9 13 1 15 9 15 9 1 9 0 1 9 0 1 9 9 0 1 9 9 9 15 2
14 9 0 13 9 0 1 9 0 1 9 0 7 9 0
41 13 9 0 1 9 9 0 1 9 0 15 13 15 9 0 0 1 9 1 9 0 1 9 7 15 13 9 1 9 0 0 1 9 1 9 0 7 0 1 9 2
18 7 13 9 0 9 9 8 8 2 10 9 0 14 13 9 9 2 2
21 7 15 13 8 0 0 1 9 0 2 7 15 8 0 1 9 7 9 0 2 2
97 7 13 8 2 10 9 15 9 1 9 7 13 9 1 9 7 9 1 9 0 7 9 15 1 9 0 1 15 9 14 13 9 1 9 7 9 0 0 1 9 2 2 0 1 7 9 0 14 13 9 0 1 9 1 15 14 9 0 9 9 8 8 7 13 7 9 0 1 9 13 7 15 13 9 7 9 7 9 0 13 9 0 7 0 7 15 0 9 9 0 1 9 1 9 9 0 2
30 7 13 9 7 2 9 0 13 9 9 3 2 7 7 3 9 0 0 1 15 9 15 7 9 15 0 7 0 2 2
24 0 7 9 1 9 0 13 9 9 9 1 0 9 0 1 9 9 1 9 9 0 1 9 2
28 7 13 7 9 1 0 7 13 13 9 9 9 7 1 9 9 15 1 9 13 9 9 0 1 9 1 0 2
9 9 0 8 12 12 2 12 2 12
15 9 0 8 8 8 8 8 13 1 9 1 9 9 7 13
59 14 9 1 9 0 1 9 10 9 14 1 9 9 9 0 15 13 9 9 1 8 9 0 8 1 9 9 15 1 9 15 13 15 2 7 15 13 9 8 7 9 15 1 9 9 0 2 13 8 3 7 15 1 0 9 1 9 15 2
22 7 9 15 13 15 0 13 1 0 1 9 2 7 7 7 15 13 1 9 9 2 2
71 7 1 12 9 1 9 7 9 7 9 1 9 0 7 0 13 9 8 8 2 0 2 2 8 8 8 8 8 2 0 2 2 1 9 1 9 9 0 15 14 13 1 9 9 15 1 9 0 1 9 1 12 9 2 7 15 13 1 8 12 9 8 8 8 9 0 0 0 1 9 2
35 9 2 8 8 8 8 2 9 15 13 9 1 0 1 9 15 7 9 15 2 7 9 15 0 13 8 2 8 13 9 15 13 9 9 2
22 9 0 1 15 13 15 1 13 15 1 9 15 9 15 1 9 1 9 15 2 8 2
11 8 0 8 8 7 15 13 1 9 2 2
67 13 8 1 2 9 2 2 2 8 1 9 1 9 1 9 8 7 9 1 15 8 9 1 9 12 7 12 1 9 9 0 0 2 7 9 1 9 15 8 8 1 9 1 9 0 7 13 9 9 0 1 9 15 12 1 9 1 7 8 8 9 1 9 1 15 2 2
61 13 8 9 0 1 9 14 12 15 13 15 1 0 1 9 0 7 9 0 2 7 13 9 15 13 1 1 9 1 9 9 2 2 14 8 9 9 15 2 8 8 1 9 8 8 8 1 9 1 7 9 0 1 15 15 8 8 8 3 2 2
157 7 9 1 8 2 0 2 8 13 1 15 2 13 0 2 0 7 9 0 15 13 1 15 1 9 15 13 15 15 7 9 9 9 2 7 15 3 15 13 1 9 2 7 10 9 1 9 2 9 1 9 0 1 9 2 7 15 13 1 9 9 0 9 2 7 13 2 2 3 9 0 0 15 13 13 1 9 9 2 13 9 1 9 8 8 8 7 9 7 9 0 1 9 7 9 0 7 1 9 13 9 1 9 9 8 8 0 1 9 9 2 7 13 15 14 13 1 9 2 13 9 1 9 13 1 15 2 8 8 9 1 9 3 2 8 8 1 9 8 8 8 0 7 13 2 7 14 8 1 9 8 8 0 1 9 2 2
59 7 1 7 13 13 8 1 9 7 9 1 9 9 2 7 9 1 9 15 0 9 2 1 0 15 8 7 9 15 0 2 13 15 2 9 2 1 9 9 0 1 15 2 13 2 2 1 9 8 9 8 2 7 9 13 1 9 2 2
73 7 1 9 9 15 1 9 9 13 2 2 8 8 9 9 1 9 15 2 8 8 1 9 15 2 7 1 8 8 1 8 8 1 9 7 9 8 8 9 0 2 8 1 9 2 7 13 2 15 9 0 2 8 8 7 8 1 15 1 9 8 8 7 13 8 8 0 8 8 8 9 2 2
47 13 9 8 1 9 0 8 1 8 7 14 13 1 9 0 7 9 0 2 7 13 1 9 9 0 13 1 9 9 2 8 8 8 1 9 15 8 13 1 0 7 9 2 7 3 8 2
26 15 13 9 0 2 7 15 14 8 9 2 14 8 8 8 8 2 8 8 8 0 15 9 15 2 2
10 8 8 2 9 1 0 7 9 15 0
64 13 9 12 2 12 0 9 8 8 9 9 1 9 0 9 9 1 9 9 8 2 0 7 9 8 0 1 9 9 9 0 7 9 0 1 9 9 8 8 1 9 9 15 1 9 0 2 7 13 15 9 1 9 9 0 9 2 7 7 13 1 9 0 2
62 7 13 9 8 8 2 13 9 12 2 12 0 15 9 0 15 13 1 15 9 9 15 2 7 14 13 15 9 2 7 13 1 9 9 1 9 0 1 9 9 7 13 9 0 1 9 7 15 13 1 9 1 9 9 1 7 13 9 15 9 0 2
42 13 8 1 9 8 8 1 9 9 0 1 9 9 0 8 15 13 15 9 9 1 9 8 8 7 13 12 1 9 9 7 9 9 7 9 1 9 0 1 8 9 2
53 7 13 9 8 8 1 9 2 8 8 8 1 15 7 13 9 1 9 15 7 9 15 7 9 7 9 8 8 9 7 9 8 8 1 15 9 7 1 15 9 15 2 7 7 9 9 0 7 9 9 8 0 2
94 7 14 13 15 9 9 1 9 15 9 1 9 9 7 9 1 9 9 8 7 13 15 9 1 9 15 2 8 8 1 9 9 8 8 8 9 9 1 9 0 2 1 7 9 1 0 7 7 9 9 15 14 13 9 0 1 9 9 0 13 1 15 1 9 9 0 1 9 2 0 1 7 9 13 9 15 0 2 7 13 8 8 1 9 9 2 7 14 8 1 9 9 9 2
45 7 14 13 9 9 0 1 9 0 1 9 1 9 8 1 9 7 9 2 7 13 7 15 13 1 15 14 13 9 9 0 2 7 7 15 9 0 1 9 9 0 1 9 8 2
13 9 0 13 1 9 1 9 0 1 9 9 9 8
30 13 9 1 9 0 9 12 2 12 0 1 9 9 9 0 1 9 9 8 2 7 15 13 13 2 9 9 0 2 2
31 7 13 9 1 9 0 1 9 1 8 8 9 9 8 8 8 9 9 1 9 8 0 0 1 9 9 0 1 9 15 2
52 7 13 9 1 7 2 1 9 1 9 7 9 15 13 9 10 9 2 7 7 15 13 9 1 9 0 0 0 1 9 1 9 0 1 9 9 15 1 0 9 7 15 13 1 15 9 8 1 9 0 2 2
14 9 9 2 9 8 8 8 9 1 9 9 1 9 2
38 13 9 9 0 12 9 13 9 15 1 9 0 0 1 9 1 9 8 8 1 9 0 2 7 13 15 9 2 9 8 1 9 15 8 8 8 2 2
108 7 13 10 9 1 9 1 9 9 0 15 13 1 15 0 0 1 2 9 9 0 2 7 15 9 15 13 15 9 1 9 9 13 1 15 7 1 9 9 0 9 0 13 1 9 15 9 12 9 13 1 9 0 0 1 9 7 13 1 9 2 11 8 2 7 13 9 1 7 10 9 13 0 1 15 0 7 13 9 9 1 1 9 1 9 1 9 0 13 2 9 10 9 1 9 9 8 8 8 8 1 9 9 9 1 9 2 2
57 7 13 8 7 9 8 8 8 10 9 7 1 10 9 2 13 9 0 0 9 1 9 0 7 0 0 9 15 7 15 13 8 8 14 13 9 15 9 1 9 15 9 1 9 8 1 9 0 15 1 9 1 9 9 9 15 2
5 13 1 0 2 2
4 7 0 0 2
71 13 8 8 13 2 9 15 13 15 9 2 0 1 9 8 8 2 9 9 9 2 1 9 15 1 9 9 2 15 9 9 0 1 9 0 9 0 10 13 1 15 2 7 15 0 2 7 7 15 13 1 9 0 2 1 10 9 2 7 13 9 0 2 1 9 15 13 1 15 0 2
38 13 9 2 1 9 15 0 2 1 8 0 1 9 2 7 15 13 9 9 15 1 9 7 9 7 9 7 9 2 7 9 9 15 1 9 7 9 2
46 7 10 9 2 1 9 9 2 13 1 15 0 2 7 15 9 1 9 0 0 2 7 0 2 13 15 9 2 1 15 2 7 13 15 9 9 2 1 9 9 15 0 2 9 9 2
56 7 7 13 9 2 1 9 9 8 2 7 0 7 13 1 0 2 7 7 13 9 1 7 9 9 2 15 13 15 7 13 1 15 2 9 9 2 1 9 15 1 9 2 7 7 15 13 1 10 9 2 7 7 15 2 2
4 7 7 15 2
9 7 7 9 9 2 15 15 13 2
99 7 13 9 0 2 1 9 9 9 2 15 7 10 9 2 13 9 9 9 15 1 9 9 2 7 9 9 15 1 9 0 2 14 13 2 7 7 15 14 13 2 7 7 9 10 9 2 9 9 0 2 7 9 15 13 9 12 12 9 2 7 9 0 9 2 15 12 12 9 2 7 7 15 7 13 2 7 14 13 15 12 12 9 2 12 12 3 2 7 13 12 12 2 1 0 7 0 9 2
5 15 9 10 9 2
74 9 15 2 1 0 9 2 7 15 14 9 2 7 7 15 14 13 13 1 9 2 9 9 9 15 2 13 15 3 2 7 7 9 15 14 13 2 7 13 2 7 13 2 7 9 9 1 9 9 0 2 7 7 9 2 1 9 2 1 9 9 2 7 14 15 14 13 2 7 13 2 7 13 2
46 1 9 2 7 1 9 0 2 13 9 9 2 1 7 15 7 9 1 1 15 2 0 1 9 9 2 1 10 9 9 2 7 7 9 10 13 15 2 15 9 9 7 9 9 0 2
21 7 3 10 9 0 9 1 7 13 2 7 13 2 7 13 1 9 7 9 2 2
53 7 7 13 9 2 0 9 2 1 1 15 13 1 15 9 9 2 7 15 9 1 9 2 7 9 0 7 0 2 15 7 13 1 9 2 7 13 9 15 2 1 9 0 2 0 1 7 13 2 7 7 13 2
30 9 7 15 0 2 1 0 9 2 14 1 9 2 15 13 1 15 9 2 7 14 13 2 1 7 13 9 15 2 2
14 13 9 9 2 7 13 1 9 2 13 1 0 2 2
5 7 0 0 2 2
6 9 0 13 9 9 9
18 13 9 0 1 9 2 9 9 9 9 2 7 9 1 9 9 0 2
51 7 13 9 8 8 2 9 9 9 9 0 2 9 9 1 9 1 9 15 7 9 9 15 2 7 9 15 9 0 1 9 0 2 8 8 1 9 9 2 7 13 7 15 8 9 9 9 7 9 9 2
96 13 9 8 8 9 9 8 8 7 9 9 9 0 7 0 9 1 9 0 2 9 0 1 9 9 1 9 15 9 0 1 9 2 7 13 8 1 9 15 2 9 9 14 13 9 9 7 14 9 7 14 9 9 9 7 13 1 15 9 2 7 7 13 1 9 7 9 2 7 7 15 14 13 0 9 7 9 13 10 9 1 10 9 0 2 8 8 9 9 9 9 0 7 9 0 2
21 7 9 13 13 2 7 15 13 1 15 1 9 1 9 8 8 1 9 0 2 2
30 8 8 9 9 9 9 9 0 15 8 1 15 12 8 9 7 9 0 2 7 8 2 7 15 0 9 9 9 0 2
48 7 13 8 8 9 9 7 13 1 9 15 2 7 7 13 1 9 15 8 8 9 15 8 8 1 15 8 8 9 2 7 9 9 9 9 7 15 9 0 1 9 0 8 8 1 9 9 2
64 7 13 8 13 8 8 2 8 9 0 2 9 1 9 1 8 8 0 8 1 15 9 8 8 1 15 9 8 8 7 1 9 8 8 2 7 7 7 7 15 1 9 7 8 1 9 9 8 8 8 7 14 13 9 0 1 15 7 13 8 1 15 1 2
36 7 15 3 9 9 0 1 9 0 1 9 9 9 0 7 0 1 0 9 0 13 15 0 9 1 9 0 7 9 1 0 9 1 9 9 2
57 9 9 13 8 8 1 9 0 13 2 9 15 13 1 9 0 1 9 0 2 8 8 2 9 1 7 9 1 9 9 2 14 13 1 9 9 2 9 2 13 9 2 7 13 1 9 1 9 9 0 15 13 1 15 9 0 2
61 7 9 0 1 10 9 2 1 9 9 15 2 15 7 9 0 1 9 15 7 9 1 9 9 2 1 9 9 1 9 15 2 7 1 9 15 13 7 13 1 15 10 9 2 0 7 9 9 0 1 9 1 9 0 2 14 13 1 14 9 2
147 13 0 1 9 0 1 9 2 15 13 1 9 0 15 13 15 1 9 9 0 2 9 9 0 1 9 1 9 9 2 7 15 13 1 9 10 9 7 15 13 9 0 1 9 2 7 7 15 13 1 9 9 13 15 1 9 1 9 9 2 15 13 9 15 0 1 9 0 1 9 0 7 0 2 7 13 1 9 13 9 10 9 1 15 13 1 9 9 1 9 0 2 13 1 15 9 7 13 9 7 7 13 15 2 7 13 9 0 1 9 7 13 1 9 15 2 1 15 13 9 0 1 9 0 1 9 15 13 15 2 7 13 1 15 9 9 9 15 7 9 15 1 1 0 1 9 2
117 14 13 1 15 13 9 0 1 9 9 0 1 9 15 1 10 9 15 13 1 15 9 1 9 9 2 7 13 1 9 9 0 7 0 1 9 0 2 7 13 9 1 9 1 10 13 9 0 9 15 1 9 2 7 1 9 10 9 0 1 9 9 2 9 0 2 1 9 1 9 15 14 13 1 9 0 2 1 7 13 2 8 8 2 1 9 9 9 1 9 9 9 9 9 0 2 9 1 9 1 9 9 0 1 9 9 0 1 9 2 1 9 15 9 1 9 2
102 9 7 9 9 0 2 13 1 1 12 9 1 9 0 7 0 2 1 7 13 9 0 7 0 2 7 9 13 1 9 9 9 7 9 0 1 9 9 15 1 9 14 13 1 0 7 0 1 7 13 10 9 9 0 7 0 7 0 14 9 1 9 1 15 1 9 9 1 9 7 9 1 9 2 13 1 15 9 9 1 9 7 9 2 1 9 9 0 0 2 13 9 0 1 9 1 1 9 9 7 9 2
50 9 0 9 1 9 9 9 0 1 9 1 9 0 15 9 9 1 7 9 0 15 13 1 15 9 9 0 7 0 2 14 13 1 9 0 0 1 9 2 7 15 9 1 9 10 9 7 9 15 2
55 7 7 14 13 9 0 1 9 9 9 0 1 1 15 2 7 1 9 9 7 13 1 9 0 0 1 9 15 2 7 1 9 15 1 9 0 7 0 1 9 1 15 7 13 9 1 9 9 15 1 15 1 9 0 2
5 9 0 8 8 8
38 9 1 9 9 15 13 1 9 1 9 15 9 15 1 9 9 13 8 8 9 9 8 13 2 9 15 13 2 8 8 2 1 9 9 9 9 2 2
18 9 9 15 9 0 2 7 9 0 2 7 9 0 1 9 0 2 2
13 7 9 7 13 2 9 2 7 13 9 9 2 2
14 7 14 15 13 1 15 9 0 2 8 0 0 2 2
12 13 15 7 13 1 9 1 9 9 1 9 2
4 1 3 2 2
8 7 7 2 8 8 2 2 2
9 15 9 9 9 0 0 0 2 2
14 13 2 7 13 1 9 9 9 0 1 9 15 2 2
13 7 13 9 0 7 0 1 9 9 1 9 15 2
5 9 1 15 2 2
15 7 7 9 2 1 9 9 2 13 1 9 15 0 2 2
8 9 0 1 9 9 15 2 2
14 7 9 9 1 10 13 15 1 9 0 7 9 0 2
3 7 2 2
10 7 13 9 9 1 0 9 0 2 2
10 9 14 13 0 2 7 9 15 2 2
9 7 13 9 7 13 9 9 2 2
20 2 7 9 15 13 0 2 7 9 0 7 13 9 2 0 2 1 9 2 2
4 7 9 2 2
16 1 9 9 2 7 13 2 9 0 1 10 9 0 2 0 2
16 8 10 13 9 12 2 12 0 13 9 0 1 9 10 2 2
10 7 14 13 9 2 8 2 0 2 2
24 1 0 0 2 7 9 2 7 9 9 2 7 9 15 13 15 9 1 9 12 9 0 2 2
8 15 13 9 1 9 9 2 2
11 3 13 9 9 1 9 7 13 9 2 2
15 7 13 9 1 9 9 15 7 13 13 1 9 9 2 2
4 9 0 2 2
13 7 7 13 15 7 13 15 1 0 9 7 9 2
9 14 9 9 1 9 9 15 2 2
16 7 9 9 1 0 9 15 7 9 15 2 7 9 15 2 2
9 13 1 0 1 9 15 8 2 2
11 7 8 8 15 9 15 13 8 8 2 2
8 8 8 9 1 9 15 2 2
6 7 9 15 0 2 2
11 7 9 15 7 9 15 2 7 9 15 2
7 9 0 2 9 9 9 8
13 13 9 0 7 9 9 1 9 1 8 9 8 2
25 7 13 9 0 1 9 2 9 0 2 0 7 9 13 1 9 0 1 9 1 7 9 9 0 2
36 7 13 9 15 14 13 9 12 2 12 0 7 9 13 1 9 12 1 7 9 9 0 2 7 14 12 5 1 9 1 15 1 8 9 8 2
21 7 13 9 1 9 13 1 15 1 9 15 9 9 0 0 7 9 15 8 8 2
35 7 13 9 9 7 12 1 9 12 9 0 13 1 7 13 8 9 2 1 1 13 12 5 1 9 7 15 0 1 9 9 1 9 9 2
29 7 13 9 1 7 12 5 1 9 8 1 8 13 1 12 9 7 13 9 1 7 9 9 13 1 9 1 9 2
12 9 13 9 9 0 1 14 9 13 9 9 0
33 13 9 0 0 1 9 0 1 15 1 9 9 9 1 14 9 2 15 10 13 1 2 9 2 9 15 0 9 7 0 1 9 2
64 7 9 0 13 12 2 12 9 2 9 0 0 1 9 12 8 9 2 2 9 15 1 9 9 8 12 13 7 13 12 8 9 7 13 1 9 12 12 9 2 12 9 2 7 13 9 1 9 12 9 2 1 15 13 1 9 9 7 9 9 1 9 0 2
30 7 1 9 9 1 14 9 2 0 0 2 7 7 9 0 13 9 7 9 1 9 0 2 1 1 9 0 1 9 2
16 9 8 12 12 2 12 2 12 9 1 9 0 1 9 0 0
41 13 9 8 7 0 0 1 9 9 0 0 1 9 13 1 9 0 2 9 1 9 1 9 9 15 13 1 9 0 2 1 9 0 7 0 7 0 13 1 9 2
39 7 14 13 9 8 7 0 10 1 9 9 13 1 0 15 9 0 15 13 9 7 13 9 0 0 9 0 13 1 9 15 13 9 0 0 1 9 9 2
40 7 1 9 0 15 13 1 9 2 9 8 0 7 3 9 9 0 0 7 9 1 9 9 7 9 9 0 13 1 1 10 9 0 7 0 15 13 15 9 2
44 7 13 9 1 9 0 7 9 0 0 15 13 9 1 9 13 1 9 0 1 9 9 9 0 1 9 9 7 1 9 15 7 13 9 0 1 9 9 1 9 1 9 0 2
125 8 8 0 10 13 1 10 9 0 1 9 1 9 9 0 9 9 1 9 0 0 1 9 0 1 9 7 3 9 0 0 8 8 7 9 0 2 7 3 13 1 9 15 13 1 9 9 0 0 7 10 9 13 0 1 9 2 7 14 13 13 9 9 8 2 9 9 0 0 1 9 8 2 7 3 1 9 0 1 10 13 1 8 8 9 9 0 0 2 7 7 0 0 8 8 13 9 15 1 0 1 9 7 1 9 9 15 13 1 9 9 7 13 2 0 14 15 1 7 15 9 0 1 9 2
59 7 13 1 8 2 0 0 0 13 1 7 9 15 13 1 15 9 15 9 1 9 7 7 15 14 9 1 7 13 9 0 9 1 9 8 13 13 9 9 0 7 0 1 9 9 9 0 2 7 15 13 1 9 9 9 0 7 3 2
79 7 7 15 13 9 0 8 8 1 9 7 15 13 9 15 13 7 13 1 10 9 1 0 9 0 1 9 1 9 7 13 9 1 9 0 0 2 7 7 15 13 9 0 1 15 15 8 9 1 8 0 2 8 7 0 7 3 9 15 7 9 15 13 1 12 9 12 9 7 9 15 1 9 1 0 0 7 0 2
39 7 13 9 0 0 7 9 1 9 1 9 9 0 13 8 1 9 9 7 9 1 9 13 0 9 0 7 0 1 7 13 1 15 13 1 15 8 0 2
34 7 13 10 9 7 2 9 9 2 7 13 9 1 15 13 9 1 9 9 7 9 0 0 7 15 15 13 9 0 0 1 9 0 2
5 9 0 7 9 0
17 13 8 8 8 9 9 9 13 2 13 9 9 1 9 9 0 2
11 7 14 13 0 1 9 9 0 0 0 2
11 7 13 9 9 15 13 15 0 1 9 2
13 7 9 1 9 14 13 8 8 1 9 1 9 2
20 10 9 0 13 0 1 9 2 7 14 1 9 2 1 9 0 1 9 0 2
25 7 14 13 3 1 0 1 9 9 15 2 7 1 9 9 9 14 13 8 1 9 7 9 15 2
21 9 0 13 9 1 9 9 13 15 15 13 1 15 1 8 1 9 0 1 9 2
34 7 9 1 9 0 15 13 0 1 9 15 1 9 9 9 13 9 1 9 13 1 15 9 0 1 9 0 13 9 9 9 0 9 2
29 7 9 9 8 8 1 9 9 15 1 9 9 0 14 13 0 1 9 1 1 10 9 1 9 0 1 10 9 2
20 7 14 13 0 1 9 9 1 9 9 0 1 9 7 13 1 15 9 0 2
43 7 7 13 8 2 0 1 0 9 15 2 1 10 1 15 9 0 15 13 9 0 1 9 0 9 1 9 1 9 9 2 2 13 9 9 0 7 13 1 9 15 0 2
18 9 0 13 9 7 4 9 0 1 9 7 9 1 9 1 9 15 2
30 9 7 9 10 9 2 7 13 1 9 2 15 9 0 9 12 15 13 9 9 0 1 9 9 0 2 1 9 9 2
19 7 13 9 1 9 10 9 1 15 13 1 9 0 9 15 1 10 9 2
15 9 0 7 9 0 14 13 7 13 2 1 1 9 0 2
19 7 13 9 0 2 9 1 9 2 13 7 10 9 13 13 1 9 15 2
13 7 9 10 9 14 13 9 1 8 7 13 15 2
19 7 8 8 14 13 9 0 1 1 8 8 2 1 9 8 9 9 15 2
23 8 8 9 9 9 0 7 0 0 1 9 0 2 1 15 13 0 1 10 9 9 2 2
51 13 9 10 9 1 15 13 15 8 8 1 9 15 1 9 15 2 8 13 14 13 0 9 13 9 0 1 9 1 2 0 2 7 15 14 13 1 8 2 7 15 9 0 1 9 7 9 7 9 9 2
24 7 9 1 9 0 1 9 14 13 15 13 15 9 12 0 7 9 0 2 1 9 9 8 2
17 13 8 9 1 9 9 7 9 7 9 2 7 13 15 13 15 2
12 15 14 13 7 14 13 1 15 1 9 9 2
31 15 7 13 1 15 0 7 14 13 1 9 15 1 0 15 0 15 13 9 15 1 9 9 15 1 9 9 1 8 0 2
48 10 9 13 8 8 7 13 9 9 9 1 9 9 0 2 1 9 1 9 9 0 1 9 9 2 7 15 13 15 1 9 7 9 2 7 1 9 9 2 7 1 9 9 0 8 7 0 2
24 13 8 1 9 9 9 15 0 9 0 2 9 9 1 9 1 0 0 7 9 8 7 0 2
15 1 10 2 9 2 14 13 0 7 13 9 13 9 9 2
52 7 1 9 8 9 10 2 9 2 1 9 2 13 1 9 15 15 13 1 9 0 1 9 0 0 9 1 9 9 1 9 2 9 2 13 9 15 9 0 0 0 1 9 9 7 0 1 9 9 7 9 2
22 7 1 10 9 2 13 9 9 1 9 0 1 9 1 9 1 9 9 1 9 15 2
19 0 13 9 15 1 9 2 9 9 2 9 1 9 0 7 0 1 9 8
55 13 9 1 9 9 9 0 8 8 8 9 1 9 9 1 7 9 9 9 7 9 9 2 9 9 0 7 9 9 9 2 14 13 15 1 9 0 0 2 7 1 7 15 13 9 0 1 9 0 0 0 1 9 0 2
57 7 7 13 0 9 0 9 8 8 7 9 9 8 8 1 9 9 0 2 13 9 12 2 12 0 1 9 8 8 13 9 15 1 9 0 1 8 7 9 2 7 15 13 7 15 2 14 13 1 9 8 8 1 9 0 2 2
33 7 13 9 9 0 8 8 8 7 12 1 9 9 15 13 9 9 0 1 8 1 9 15 0 9 9 0 13 9 1 12 9 2
27 7 13 9 8 8 9 12 2 12 0 9 9 0 7 13 1 15 9 1 9 0 7 9 7 9 0 2
8 7 13 9 9 1 9 15 2
22 7 1 0 7 13 8 1 9 9 0 2 1 9 9 1 9 1 9 0 7 0 2
70 7 13 9 9 0 1 9 7 9 15 2 0 1 9 9 9 7 9 0 2 7 13 1 9 9 9 0 7 0 7 0 1 1 9 0 1 9 9 9 9 7 9 9 1 9 2 2 0 1 7 9 9 15 1 9 2 14 7 14 13 0 9 1 9 15 1 9 0 2 2
19 7 13 10 9 1 9 1 9 2 9 9 2 15 13 9 0 7 0 2
17 7 13 8 7 9 15 1 0 9 1 2 9 15 1 15 2 2
31 7 7 12 9 14 13 1 9 2 1 15 9 1 9 12 12 9 1 9 9 7 9 15 1 9 0 1 9 1 9 2
76 7 13 9 0 13 1 9 0 9 1 9 2 8 8 2 7 2 8 8 8 2 0 1 9 1 9 7 9 15 7 9 15 1 9 13 1 9 1 9 2 7 13 9 15 12 9 0 1 9 12 9 2 7 13 15 9 0 1 9 0 15 2 8 2 1 9 9 8 1 9 0 0 1 9 0 2
34 7 13 9 2 9 9 2 1 9 9 2 9 0 2 1 0 2 15 13 1 9 9 15 1 1 9 8 8 2 9 9 10 9 2
32 7 13 9 9 0 8 8 2 2 1 9 13 9 0 2 13 9 0 0 2 2 0 1 9 9 1 9 9 13 1 0 2
38 7 13 2 9 0 1 9 2 7 2 8 8 2 9 12 2 12 0 9 1 9 12 12 9 1 9 9 7 9 15 1 9 0 1 9 8 8 2
33 7 13 9 8 7 2 8 8 2 15 9 9 15 13 1 9 1 9 9 1 9 2 13 9 0 1 9 15 1 12 12 9 2
19 7 13 9 0 1 9 8 8 7 9 9 15 14 13 1 9 9 0 2
6 12 5 9 9 1 9
56 13 9 0 0 7 9 9 0 1 9 14 13 12 5 1 0 9 9 0 2 12 9 7 0 2 1 15 1 10 9 0 0 7 15 1 9 15 8 7 9 2 8 8 1 0 8 9 9 0 1 9 9 7 9 0 2
38 7 13 9 1 9 9 7 9 0 0 9 15 13 0 1 9 9 7 15 1 12 7 12 5 1 9 9 7 13 15 13 1 9 7 9 1 9 2
47 7 13 7 9 9 0 1 9 0 1 9 13 7 1 9 9 1 9 1 12 12 9 1 1 9 9 0 0 9 15 12 9 1 9 0 7 13 9 9 0 12 12 9 1 0 0 2
12 9 0 2 0 1 9 9 1 9 0 1 9
56 13 9 0 1 9 9 0 7 9 15 13 9 9 1 9 9 0 1 9 9 1 9 0 1 9 15 13 1 12 12 9 9 0 2 7 9 9 0 15 14 13 12 12 9 1 9 1 9 13 1 15 13 12 12 9 2
34 7 13 9 1 7 10 9 14 13 1 9 9 0 1 9 1 9 1 9 0 2 7 9 9 9 9 1 9 0 7 9 15 0 2
87 7 13 1 2 9 0 2 9 0 7 3 0 1 12 9 13 9 0 7 13 1 9 15 1 9 1 9 1 9 2 1 10 9 2 0 1 7 0 10 9 13 1 9 9 9 7 9 7 9 7 9 7 9 1 9 7 9 0 2 0 1 7 9 0 15 13 1 9 0 14 13 9 15 12 9 9 2 13 1 9 9 7 9 9 7 9 2
26 7 13 9 7 9 13 0 0 9 0 1 9 1 9 0 2 7 7 9 9 1 9 13 1 9 2
39 7 13 9 8 8 8 9 9 1 9 0 0 2 7 3 9 0 0 1 9 7 9 2 1 9 9 1 0 9 2 1 10 1 10 9 0 7 0 2
34 7 13 9 7 9 14 13 8 8 0 1 9 12 2 7 13 1 9 12 9 9 0 13 1 9 15 9 9 1 8 1 9 9 2
8 9 0 9 1 9 0 1 9
64 13 9 9 9 0 9 0 9 9 7 9 0 1 9 0 9 1 9 9 9 1 9 9 0 1 1 9 9 8 8 1 12 9 0 1 9 1 9 0 0 7 0 0 7 0 8 8 1 9 1 12 1 0 9 15 1 15 9 9 0 1 9 0 2
38 13 8 9 8 8 8 9 9 0 1 9 15 13 9 12 2 12 0 1 9 9 9 0 7 9 9 7 9 0 1 9 0 7 9 1 9 0 2
86 7 13 8 7 15 1 0 7 13 1 9 9 0 1 9 0 10 1 9 0 7 9 9 13 1 9 15 9 9 7 9 9 0 1 10 9 1 9 9 0 1 9 1 1 9 0 2 0 1 7 9 14 13 9 0 1 9 9 1 9 7 9 9 9 1 15 13 1 9 0 9 15 7 14 13 9 1 9 0 1 9 1 9 9 9 2
29 7 13 8 9 9 1 9 9 15 0 1 9 10 9 1 9 9 1 15 13 9 9 7 9 15 1 9 0 2
8 9 1 9 9 0 2 9 0
51 13 2 9 9 0 2 9 0 2 9 1 9 2 9 12 2 12 0 2 1 9 9 1 9 7 9 9 9 8 1 9 1 8 2 8 2 8 2 8 2 8 2 8 8 8 2 1 9 1 9 2
57 7 13 9 9 2 8 0 2 7 15 14 13 1 9 2 9 9 9 9 9 0 2 15 13 9 15 1 8 2 7 9 9 9 0 1 9 0 2 9 9 2 7 9 9 9 1 9 0 0 1 8 1 9 1 9 15 2
12 9 13 9 1 9 9 9 1 9 8 7 8
35 13 9 9 0 8 8 8 9 12 2 12 0 9 1 9 8 13 12 9 1 9 9 13 9 1 9 9 1 9 9 9 0 7 0 2
63 7 13 9 1 9 1 2 9 9 9 0 2 7 9 8 7 9 15 9 0 8 8 14 13 1 9 9 0 1 9 9 0 1 9 0 9 2 1 9 1 9 9 0 7 9 9 9 1 9 1 9 15 7 1 15 13 9 9 0 1 10 9 2
23 7 13 1 7 9 7 9 8 9 1 9 9 12 15 13 9 9 0 1 9 9 0 2
71 7 13 9 7 9 8 7 9 0 1 15 13 1 9 9 1 9 0 7 0 0 1 9 0 7 15 13 9 15 0 1 12 12 9 13 9 0 0 13 1 9 0 1 9 7 9 9 7 3 9 9 2 7 15 15 13 1 9 9 0 0 1 9 0 1 9 0 7 0 9 2
102 7 13 9 1 7 10 9 13 1 9 9 12 0 1 9 9 0 1 9 1 1 9 9 0 13 1 9 7 8 7 9 8 2 1 9 7 15 9 0 1 9 9 0 1 15 2 9 1 9 9 15 0 0 7 0 2 7 1 9 9 15 0 2 9 1 9 9 8 7 8 1 9 9 8 7 9 8 1 9 9 0 2 7 1 9 9 0 15 13 1 9 9 0 7 0 1 15 7 1 9 0 2
32 7 13 9 7 15 13 9 9 1 9 9 0 0 1 9 8 1 9 0 2 9 8 2 1 9 9 0 1 9 7 8 2
37 7 13 7 15 1 10 9 7 14 9 13 1 9 1 9 8 7 8 1 9 15 1 9 9 1 9 9 0 9 9 1 15 1 9 7 0 2
37 13 1 7 9 9 8 13 1 9 9 0 0 7 9 0 0 0 1 9 0 2 7 15 15 13 1 9 9 7 9 9 8 0 1 9 0 2
46 7 13 9 7 9 1 9 7 9 8 1 9 9 9 0 14 13 1 9 1 9 0 1 9 9 9 1 9 1 9 7 1 1 9 9 7 9 9 9 13 9 0 0 7 0 2
49 7 13 7 13 9 0 1 9 2 15 14 13 9 9 15 1 9 1 9 0 1 8 7 9 0 2 1 9 9 7 13 9 0 1 9 1 9 9 0 1 9 9 0 1 9 7 9 0 2
31 7 13 9 8 1 9 8 0 0 0 2 14 13 9 0 1 9 15 1 9 9 9 14 13 1 15 1 9 9 8 2
88 7 13 9 9 0 0 1 9 0 1 12 9 0 2 0 9 1 9 9 1 9 15 13 9 15 2 9 7 9 8 7 8 2 7 0 9 0 7 9 1 9 9 0 1 9 0 7 0 1 9 9 8 2 8 2 15 13 12 9 9 1 0 2 7 9 0 9 0 2 7 13 9 0 0 1 9 0 1 9 9 0 13 1 9 2 8 2 2
10 9 0 1 9 9 0 1 9 7 9
48 13 9 0 0 0 1 9 1 9 15 13 15 9 12 2 12 1 9 8 8 8 9 9 0 7 9 8 8 9 9 9 9 9 9 1 9 9 8 15 13 9 7 9 7 9 8 8 2
74 7 13 15 9 15 1 0 9 1 15 1 9 0 1 9 1 12 9 0 1 9 9 1 9 0 1 9 0 0 9 1 9 12 0 1 7 13 9 0 1 9 0 0 0 1 9 9 1 15 13 9 0 1 9 9 9 7 9 1 8 7 14 9 12 7 9 13 15 9 9 1 9 0 2
59 7 13 9 8 8 8 9 9 0 1 9 1 9 15 13 9 1 15 1 9 2 0 7 0 2 1 9 9 0 0 1 9 8 8 1 9 9 0 8 8 0 1 7 1 9 9 0 1 10 9 7 13 9 1 9 1 9 0 2
21 7 13 1 9 15 9 12 2 12 0 1 9 1 8 8 9 9 0 7 13 2
7 8 8 9 9 7 13 2
96 8 8 8 9 9 7 15 13 9 1 9 9 1 9 9 0 1 9 7 9 9 1 9 1 9 0 0 1 9 7 13 9 9 9 9 1 15 9 1 9 9 9 0 0 1 9 0 1 9 1 15 13 1 0 1 9 15 13 9 9 0 1 9 1 9 7 9 7 15 7 13 1 15 9 9 1 9 9 9 15 13 1 9 9 15 1 9 7 9 9 9 15 1 9 0 2
22 7 13 8 1 7 9 10 9 1 9 15 9 1 9 9 9 1 10 9 1 9 2
54 7 13 8 2 8 7 15 1 9 1 9 1 9 9 0 1 9 7 9 8 7 15 1 15 13 10 9 0 1 9 9 15 13 9 9 9 1 9 9 9 0 7 15 13 15 1 9 0 7 9 0 1 9 2
79 7 13 7 15 1 9 1 7 15 14 13 9 9 9 9 9 0 1 9 0 1 9 9 1 0 9 12 8 7 15 13 9 1 9 1 9 9 0 1 7 15 13 9 1 7 15 15 0 1 9 1 9 0 14 13 9 15 0 1 7 7 15 1 0 9 13 9 0 0 1 9 7 1 9 0 1 1 9 2
45 7 13 7 15 13 9 1 7 14 13 3 9 9 0 1 9 0 7 14 13 0 1 9 0 1 9 7 15 14 13 9 9 1 9 7 9 9 10 13 8 10 9 1 9 2
38 7 1 9 15 13 8 2 8 8 8 9 9 0 7 15 13 9 1 9 9 0 1 9 7 9 9 1 9 0 7 15 9 1 9 1 9 0 2
31 7 13 8 2 8 8 9 9 0 1 9 9 1 9 1 9 9 9 0 15 1 0 8 14 9 1 15 1 9 0 2
71 7 1 9 0 13 8 8 9 9 9 0 7 9 0 1 9 1 9 12 14 13 9 0 1 9 1 9 12 7 13 9 9 1 12 12 9 1 9 12 1 1 13 9 0 1 12 8 9 1 12 8 9 0 1 9 9 0 0 1 9 9 13 1 1 12 12 9 1 9 12 2
59 7 14 13 9 9 9 9 0 15 13 1 15 9 0 1 9 1 9 9 12 1 12 8 9 1 15 12 8 9 9 0 7 12 8 9 9 1 9 0 1 1 13 9 9 12 9 1 15 12 9 9 0 7 12 9 9 9 0 2
35 14 1 9 1 0 0 7 13 9 9 0 1 9 9 9 0 1 9 0 1 9 1 9 12 12 9 1 1 9 8 8 7 9 0 2
10 0 9 1 9 0 13 9 15 1 9
54 13 9 8 8 8 9 9 7 9 7 0 0 0 7 9 9 0 14 13 1 9 9 1 9 0 1 9 9 15 0 1 9 9 9 9 1 9 1 9 9 15 9 0 1 9 9 0 1 9 1 9 9 9 2
62 7 13 9 9 1 9 15 13 9 12 2 12 0 1 9 9 9 0 9 1 9 0 1 9 0 1 9 9 1 9 7 9 9 0 15 13 9 0 1 9 0 7 13 9 9 0 1 12 5 1 9 9 7 13 9 0 1 0 1 12 9 2
48 7 13 7 9 9 0 13 1 9 9 15 13 1 9 9 9 7 9 9 9 9 0 0 7 0 1 9 9 7 13 1 9 9 7 9 9 1 9 9 0 1 9 0 1 9 0 9 2
67 7 13 1 7 9 9 7 9 9 9 0 14 13 1 9 9 2 0 1 0 9 7 14 13 9 9 0 1 9 1 1 7 1 9 9 9 7 14 13 9 9 1 0 9 1 7 14 13 9 1 12 5 1 9 7 9 9 9 9 1 9 12 9 9 12 9 2
40 1 9 15 2 13 9 8 8 8 9 9 0 7 9 9 9 0 1 9 0 13 9 1 9 9 0 7 13 9 9 0 9 9 7 9 1 9 9 9 2
55 7 13 7 15 13 9 12 9 1 9 1 12 9 7 7 3 9 1 9 1 9 1 9 13 15 1 12 2 12 5 0 7 14 13 9 1 9 9 1 9 9 15 13 15 9 0 9 0 7 0 7 0 9 0 2
49 7 13 1 7 9 9 0 9 14 13 9 15 1 9 9 13 9 15 1 12 12 9 0 7 9 9 15 13 9 15 1 12 12 9 0 7 13 7 10 9 14 13 12 5 1 9 9 0 2
59 7 13 9 8 8 9 9 9 0 7 9 9 0 13 9 0 0 13 1 9 9 7 13 10 9 13 3 1 9 0 1 9 0 7 3 1 9 0 7 14 13 10 9 1 0 7 0 9 9 9 0 7 14 13 9 9 7 9 2
13 13 12 9 0 1 9 0 1 9 1 9 7 9
86 13 9 8 0 2 9 9 9 0 1 7 9 9 1 9 9 9 0 15 13 15 9 9 7 9 1 9 8 13 1 9 9 9 0 0 9 9 7 9 9 8 1 9 1 9 9 9 9 0 1 9 9 1 9 0 1 9 1 9 7 9 9 7 9 7 9 9 9 2 8 2 1 10 13 1 9 9 1 9 7 9 9 9 0 0 2
34 7 13 7 15 13 9 1 9 9 1 12 9 1 9 12 9 7 13 9 1 12 9 13 9 0 1 9 7 12 9 13 9 15 2
60 7 13 9 1 12 9 1 9 1 9 0 1 9 9 0 1 9 0 1 9 7 9 8 7 13 9 7 15 13 1 9 9 1 9 8 9 15 13 15 9 9 0 1 9 0 7 0 1 9 1 9 7 9 1 12 9 1 9 0 2
28 7 13 7 9 13 1 9 1 9 0 1 9 0 1 9 9 9 9 1 9 0 7 9 9 0 1 15 2
9 9 9 9 0 1 12 9 1 9
13 13 9 9 0 9 15 1 9 1 9 9 0 2
13 13 9 9 1 12 9 1 9 12 9 1 9 2
11 7 13 9 14 13 12 9 1 9 0 2
52 7 13 9 0 7 9 14 13 9 0 1 9 9 9 0 0 2 7 15 14 13 1 9 0 1 9 9 9 9 15 13 15 1 9 7 14 13 12 9 1 9 7 13 9 0 1 9 1 12 9 9 2
27 13 9 9 1 9 9 9 9 1 9 9 7 8 1 9 1 9 9 1 9 0 15 13 1 9 8 2
18 13 7 9 15 13 9 15 9 0 1 9 0 14 13 12 12 9 2
12 7 13 0 15 13 15 9 15 12 12 9 2
14 7 14 13 9 9 9 0 12 5 1 9 0 2 2
4 9 9 9 9
21 13 9 9 1 9 9 9 7 9 9 0 1 9 9 1 9 0 12 12 9 2
36 7 13 9 8 9 9 9 9 0 7 9 9 13 9 7 13 9 0 1 1 12 12 9 1 1 13 9 9 0 9 15 13 12 12 9 2
35 7 13 8 8 7 9 13 1 9 15 12 9 0 1 9 15 9 9 0 7 9 9 1 9 9 7 9 9 8 7 9 9 0 2 2
12 7 13 7 10 9 13 1 1 9 0 13 2
50 7 14 13 9 0 9 9 1 9 9 7 9 0 7 9 7 13 9 9 1 9 8 13 1 9 1 8 7 13 9 15 9 12 1 1 13 9 9 0 1 9 12 7 13 9 1 8 1 8 2
7 0 9 8 0 0 8 9
53 13 9 0 1 9 8 8 9 9 15 1 9 0 9 12 2 12 0 7 13 8 2 8 9 9 7 9 9 9 0 1 9 0 0 9 1 9 1 9 0 1 9 9 7 9 0 0 7 9 9 0 0 2
65 7 14 13 8 2 8 8 9 9 0 1 9 7 15 14 13 9 1 9 7 9 9 0 1 9 1 9 9 9 8 8 9 1 9 0 7 9 0 7 9 7 13 9 9 9 9 0 1 9 0 1 9 1 9 9 8 13 9 1 15 9 9 0 0 2
34 13 9 9 0 12 12 9 13 1 15 9 0 12 12 9 1 9 9 9 9 9 0 1 15 7 13 9 9 9 7 9 7 9 2
25 13 8 2 8 7 9 14 13 1 9 9 1 9 7 9 7 15 9 9 9 9 1 9 0 2
85 7 13 8 2 8 9 9 1 9 0 15 13 15 9 8 8 1 15 1 9 9 0 7 9 15 2 8 13 9 9 9 7 9 0 0 14 13 1 9 9 1 9 15 1 9 9 0 2 7 13 9 1 15 9 9 9 0 1 9 0 7 15 13 9 9 0 1 15 2 12 9 2 9 9 0 7 13 1 9 12 9 1 9 0 2
22 1 9 0 13 1 9 9 9 0 9 1 0 9 9 7 9 0 7 13 12 9 2
55 7 13 8 8 9 9 0 0 7 9 13 1 9 1 10 9 7 9 9 15 1 0 1 9 8 8 14 9 8 0 0 8 13 9 9 9 0 1 9 7 13 7 13 9 1 9 9 9 7 9 0 8 8 0 2
57 7 13 9 0 1 9 9 0 0 1 8 14 13 1 9 0 1 9 9 0 1 9 8 8 0 1 8 1 9 13 1 12 5 1 9 9 15 1 1 13 9 15 0 7 1 0 8 0 1 9 13 1 12 5 9 0 2
20 7 1 0 7 13 9 0 1 9 9 9 7 9 9 9 0 1 9 0 2
24 7 13 8 7 9 14 13 1 15 9 1 9 9 7 9 0 7 9 7 1 1 15 9 2
26 13 15 1 9 9 9 9 0 1 9 9 0 0 7 15 13 1 9 9 9 0 1 8 9 1 9
6 8 13 9 1 9 9
58 13 9 0 1 9 9 7 15 13 9 1 9 9 1 9 7 8 13 9 9 0 1 9 7 9 0 13 9 1 15 7 15 9 1 9 7 9 0 1 9 9 0 7 9 1 9 9 1 9 9 1 9 7 9 0 0 2 2
23 8 8 1 9 15 13 15 9 8 8 9 9 7 9 0 0 1 9 9 0 1 9 2
33 7 13 1 7 9 1 9 0 7 9 0 0 1 9 7 14 13 9 0 9 12 12 9 9 1 9 1 9 9 0 1 9 2
25 7 13 9 0 9 9 1 9 0 1 9 15 13 9 15 7 9 1 15 9 9 7 9 0 2
23 7 13 9 9 0 1 9 9 9 0 1 9 9 1 9 7 9 0 13 1 9 0 2
100 1 9 1 9 8 15 13 9 9 9 0 1 9 9 9 0 1 9 0 1 9 9 7 3 9 9 0 1 9 1 9 0 7 9 9 0 1 9 9 0 1 9 0 7 15 13 13 15 1 12 7 12 9 1 9 7 13 9 9 1 9 1 9 0 0 7 15 15 13 13 9 9 1 9 9 1 9 7 9 13 9 0 15 13 1 12 12 9 7 14 13 9 9 15 9 15 0 1 9 2
9 9 9 0 7 0 1 9 9 9
63 13 12 9 0 7 0 9 9 0 1 9 0 9 0 9 9 1 15 13 9 9 9 1 9 0 7 15 1 9 9 0 0 1 9 9 9 0 1 9 0 1 9 0 1 9 9 9 9 9 9 1 9 9 15 1 9 7 9 9 0 1 15 2
63 7 13 9 1 9 0 0 7 9 15 13 0 1 15 13 9 1 9 8 0 1 9 9 7 13 9 9 12 12 9 0 1 9 7 13 9 9 0 7 0 1 9 9 0 0 1 1 12 12 9 0 1 9 9 1 15 1 9 9 0 7 9 2
50 7 13 7 9 2 9 0 2 13 15 0 1 9 9 1 9 9 1 9 12 12 9 0 2 7 7 15 13 9 9 9 9 15 12 12 9 0 1 9 9 9 1 9 9 1 15 1 9 9 2
30 7 13 9 8 1 9 0 9 15 12 12 9 0 1 9 9 9 7 9 1 9 14 7 15 14 13 9 1 9 2
92 7 13 9 0 0 14 13 1 9 9 9 0 1 1 12 9 0 1 9 0 1 9 1 9 13 12 12 9 0 7 13 1 9 15 9 9 0 15 13 1 15 9 1 9 7 13 9 9 9 0 7 9 9 9 7 9 0 1 9 2 7 13 9 9 1 1 12 12 9 13 1 15 9 9 7 9 0 1 9 12 5 1 15 13 9 8 0 1 1 12 5 2
27 13 7 9 13 14 13 9 12 9 0 0 7 0 9 9 0 0 7 15 13 9 15 12 8 9 0 2
11 9 1 9 7 9 9 0 1 8 1 8
37 13 9 8 8 9 9 9 1 9 0 7 9 13 9 1 9 0 1 8 0 1 9 9 7 9 7 9 7 13 9 9 9 0 1 9 2 2
57 7 13 7 9 9 13 9 7 13 1 9 9 0 1 9 1 9 9 0 1 8 7 1 9 0 9 9 9 2 8 2 1 9 1 9 7 9 0 1 9 0 1 15 7 1 9 9 9 9 7 9 9 0 1 9 0 2
70 7 13 1 9 15 1 9 9 9 9 0 2 9 0 7 9 0 15 13 15 9 9 0 1 9 1 9 0 7 1 9 15 9 9 0 7 9 9 1 9 7 9 0 0 1 9 15 0 9 9 7 9 9 1 9 9 1 9 9 9 2 9 0 2 7 9 9 0 0 2
62 7 13 8 8 9 9 9 9 0 0 1 9 8 7 15 13 0 9 9 9 1 9 9 0 1 8 1 9 9 9 0 7 9 0 0 1 7 9 9 0 1 8 13 7 13 1 12 12 9 1 9 0 9 1 12 12 9 1 9 12 2 2
39 7 13 9 9 9 9 1 9 15 13 9 0 1 9 1 9 0 7 9 9 15 7 15 2 9 9 9 0 0 1 9 1 9 0 1 9 1 15 2
9 12 12 9 9 9 1 8 1 9
27 13 9 8 1 9 7 9 8 1 1 9 9 1 15 1 9 9 0 1 9 13 9 15 12 8 9 2
50 13 9 15 13 1 15 8 9 9 1 9 0 7 9 1 9 1 9 9 0 1 9 1 12 9 9 0 1 9 8 7 8 7 8 7 9 9 1 9 7 9 9 9 1 9 8 8 2 8 2
12 7 9 7 9 9 0 8 1 9 9 0 2
47 7 13 8 8 9 0 9 8 2 8 7 9 13 9 1 9 1 9 9 1 9 7 13 9 9 1 15 0 1 12 9 7 9 0 7 0 1 9 1 9 9 13 12 9 1 9 2
6 9 9 9 9 7 9
73 13 9 0 7 0 1 9 7 9 9 0 7 0 9 1 9 0 0 15 13 9 1 0 9 2 7 13 1 9 9 0 0 0 0 9 0 1 9 9 1 9 7 13 1 1 15 12 9 1 9 1 9 7 9 13 1 9 0 1 9 7 9 1 9 9 0 7 0 7 0 7 0 2
100 7 9 1 15 13 9 9 9 0 1 9 7 9 1 9 12 5 1 9 9 1 9 12 7 13 9 9 0 1 9 15 13 12 12 9 1 15 9 9 1 9 9 15 12 12 9 2 7 9 0 1 9 9 15 12 12 9 9 12 7 1 15 7 7 9 9 0 1 9 14 13 9 12 5 1 0 1 9 9 0 1 9 7 13 9 9 1 9 1 9 0 1 15 1 9 9 0 1 15 2
72 13 1 15 8 8 9 9 0 1 9 0 1 9 0 7 9 0 3 1 9 9 0 1 9 1 9 0 1 10 14 3 1 9 9 9 9 0 0 9 12 1 9 9 15 0 1 9 9 1 9 0 13 1 9 0 12 5 2 7 14 13 1 15 9 0 1 9 9 9 1 9 2
11 9 0 1 9 1 9 9 9 9 1 8
82 1 9 15 13 1 15 9 9 7 9 0 0 7 9 9 9 7 9 0 1 9 0 1 9 2 9 1 9 9 9 9 1 9 8 1 9 9 12 2 13 9 1 9 9 7 9 2 0 0 2 1 9 9 9 0 1 9 8 2 7 15 13 1 9 9 15 1 9 7 13 9 0 9 0 1 9 9 0 1 9 9 2
45 7 13 9 9 9 2 9 9 0 1 9 9 7 9 2 14 13 14 7 13 1 10 9 1 9 15 9 13 9 7 9 0 15 13 9 14 13 1 12 1 9 7 9 2 2
31 7 13 9 15 13 13 1 2 9 0 2 0 2 2 9 9 9 14 13 9 15 14 13 9 7 13 1 9 1 9 2
23 7 7 10 9 0 1 9 0 7 0 1 9 13 1 15 9 8 9 9 7 9 2 2
5 9 0 7 9 8
32 13 8 8 13 2 14 13 9 9 1 10 9 1 9 2 9 0 7 0 0 2 9 0 7 0 0 2 9 9 1 9 2
5 9 13 1 9 2
12 13 9 0 9 0 15 13 15 9 9 8 2
10 14 13 9 15 1 9 9 9 0 2
16 13 9 15 1 9 1 9 13 1 9 9 7 13 7 13 2
4 7 15 13 2
13 13 8 13 7 9 12 9 9 0 1 9 0 2
16 1 9 9 8 8 13 1 9 9 0 9 9 7 9 9 2
8 9 1 9 7 9 1 8 2
6 9 9 7 9 0 2
6 9 9 7 9 9 2
11 9 1 9 1 9 7 9 9 1 9 2
20 13 0 7 8 9 0 1 9 8 8 7 9 8 8 7 9 8 11 8 2
16 8 1 1 7 8 9 9 15 13 9 1 15 8 1 15 2
23 9 9 9 1 9 9 7 9 0 7 9 9 9 1 0 7 9 1 9 15 1 9 2
8 9 1 9 14 13 1 9 2
16 13 9 9 1 9 9 9 0 0 1 9 9 0 1 9 2
6 13 1 9 0 0 2
7 14 13 15 13 1 15 2
10 1 15 9 7 13 1 9 0 3 2
10 7 9 14 13 0 14 1 9 0 2
12 9 0 14 13 9 9 7 9 9 9 9 2
10 1 8 8 13 8 8 1 9 0 2
21 14 13 9 2 1 9 7 1 15 2 1 9 7 8 8 13 0 1 9 15 2
12 13 9 7 13 9 7 13 9 1 8 8 2
7 13 7 15 13 9 9 2
11 1 15 13 9 9 0 0 7 9 0 2
11 9 14 13 1 9 7 14 13 9 15 2
14 9 8 13 1 12 7 9 1 8 13 9 1 9 2
13 14 13 9 9 9 9 8 1 9 9 15 0 2
8 13 8 8 0 1 9 15 2
48 14 13 9 2 8 2 1 9 7 9 0 0 15 0 9 1 9 9 1 9 15 9 12 2 8 8 8 7 8 8 7 8 9 9 8 8 9 0 9 1 9 15 13 1 9 0 0 2
7 14 13 8 11 8 9 2
21 13 13 1 9 1 9 7 14 15 0 1 9 9 0 7 9 9 0 7 0 2
12 14 15 9 9 9 0 7 9 9 1 15 2
8 9 0 7 9 9 9 3 2
17 7 1 9 9 9 13 0 9 1 9 15 7 13 9 1 9 2
6 9 2 9 9 2 2
6 9 1 2 9 0 2
28 1 9 9 0 0 2 13 9 9 0 1 9 9 1 9 9 9 9 1 9 0 9 0 1 9 15 0 2
55 7 13 9 9 1 15 1 9 1 9 9 9 15 13 1 9 0 1 9 0 1 9 9 9 12 2 9 2 9 9 2 7 13 13 1 9 0 9 9 0 1 9 0 7 0 2 15 0 15 13 13 9 7 9 2
66 7 13 9 9 9 9 8 8 8 1 2 9 2 7 9 9 13 0 1 12 9 7 15 14 13 1 9 2 0 1 7 15 2 13 3 1 9 9 0 1 9 15 9 7 9 1 9 1 10 2 7 13 1 9 1 9 9 7 9 1 15 1 9 15 2 2
38 7 13 2 2 0 10 13 1 15 15 9 9 2 9 1 7 15 14 13 9 9 7 9 1 1 9 9 15 2 9 1 9 9 0 1 9 2 2
12 9 9 0 13 1 9 2 9 9 1 9 2
44 13 9 8 8 9 12 2 12 0 9 9 0 2 9 8 8 2 12 9 2 1 7 13 9 9 1 15 13 1 7 15 13 0 15 13 1 15 2 9 9 1 9 2 2
26 7 13 9 10 9 2 9 2 1 9 0 1 9 0 1 9 0 0 1 9 1 9 9 7 9 2
27 7 13 9 9 1 9 0 7 15 0 1 9 2 13 9 15 7 13 1 15 9 1 9 0 1 15 2
56 7 13 0 9 9 1 9 0 13 7 9 15 13 0 2 7 7 15 13 1 9 1 9 2 7 13 1 15 8 7 13 9 15 1 9 1 9 2 7 13 1 15 13 9 15 7 13 2 7 13 1 15 12 12 9 2
104 7 13 7 9 8 13 7 13 0 1 15 1 9 0 1 9 9 7 13 1 15 9 0 1 9 9 9 1 8 2 7 13 9 15 13 9 9 1 9 7 13 9 1 15 1 9 9 7 9 2 7 13 9 2 2 8 13 1 9 15 9 0 2 2 7 13 9 8 8 1 10 9 7 13 1 15 2 2 1 15 14 13 1 15 1 9 1 9 12 9 2 7 7 8 8 1 9 13 7 13 12 9 2 2
12 9 0 13 1 9 2 9 9 1 9 0 2
34 13 9 0 1 2 9 2 1 0 9 1 9 1 9 0 13 1 9 0 1 9 0 1 9 2 9 13 1 9 0 1 9 2 2
28 7 13 9 7 9 0 14 13 0 9 0 7 15 1 9 2 9 0 2 15 13 9 15 1 9 1 9 2
24 7 9 2 9 2 0 13 9 1 2 9 0 7 9 1 9 7 9 0 7 9 9 2 2
65 7 13 9 1 2 9 2 1 9 13 15 2 9 9 0 2 15 13 1 1 9 8 11 8 2 2 14 9 9 1 9 2 13 1 9 9 7 9 9 7 9 8 7 1 9 10 1 9 0 1 9 1 7 13 1 9 0 2 9 9 1 9 0 2 2
21 7 13 9 2 2 7 9 9 13 1 9 7 9 7 9 7 9 9 7 9 2
15 7 13 9 9 1 9 9 7 1 9 15 8 11 8 2
4 9 13 1 9
17 2 2 13 8 8 13 2 1 9 9 9 0 1 9 0 2 2
75 13 9 8 0 13 1 9 9 9 9 2 7 13 9 15 13 15 9 0 1 9 9 9 0 13 0 1 9 0 1 9 2 1 9 7 0 1 9 0 13 7 9 0 13 1 9 9 1 9 0 7 1 9 9 9 1 9 9 2 7 7 15 13 1 9 9 0 9 15 15 13 15 1 9 2
61 2 2 7 13 9 0 7 15 13 9 9 9 13 9 0 1 9 8 15 13 9 0 1 9 9 0 2 7 7 10 9 13 9 9 9 0 1 9 7 1 9 15 9 9 7 9 9 8 0 7 9 9 0 7 9 0 1 9 1 9 2
44 2 2 7 1 9 9 2 13 9 9 9 1 9 9 0 1 9 1 9 2 7 7 9 15 13 1 9 1 9 7 9 1 9 0 0 1 9 9 9 0 1 9 0 2
49 7 14 13 10 9 0 8 8 2 7 13 9 1 9 9 9 1 9 7 15 13 1 9 15 9 9 9 9 2 8 1 9 9 0 1 9 2 9 1 9 0 9 15 13 15 1 8 2 2
20 7 9 9 0 15 13 13 9 0 1 15 9 1 9 9 7 9 1 9 2
46 1 9 1 9 9 0 13 9 9 0 7 15 9 9 1 9 7 9 0 0 1 9 2 7 15 13 9 9 8 2 15 9 2 7 9 8 7 9 1 9 15 7 9 15 0 2
40 2 2 7 7 13 0 1 9 0 7 0 7 0 13 1 9 9 0 0 1 9 2 7 14 9 0 14 13 1 9 9 0 1 9 15 1 9 9 2 2
44 1 7 13 0 9 0 0 2 1 7 10 9 13 9 15 4 1 9 9 3 7 7 3 9 1 9 9 0 15 13 9 7 8 9 1 15 2 7 9 15 1 9 15 2
9 12 12 9 9 9 1 9 9 9
27 13 9 9 9 9 0 0 1 1 9 9 9 9 1 9 0 1 9 0 7 0 1 1 12 12 9 2
30 7 13 9 13 1 9 9 12 9 12 1 12 1 9 9 15 1 8 7 13 9 0 2 7 15 0 2 1 8 2
40 7 13 9 0 1 9 9 9 0 1 9 9 0 1 9 15 13 9 15 13 15 9 0 1 9 0 1 9 1 9 9 1 9 0 7 1 9 9 15 2
51 7 13 9 9 7 9 0 0 8 8 13 1 9 0 1 9 2 8 2 1 8 2 7 9 9 9 1 9 7 9 0 1 9 13 1 9 9 0 1 9 2 8 2 15 13 9 9 15 1 9 2
41 7 13 9 0 12 12 9 1 9 9 9 12 7 13 9 15 1 1 12 12 9 9 0 14 7 9 0 1 10 9 13 1 9 9 9 9 1 9 9 0 2
16 8 13 9 9 1 9 0 2 8 15 13 1 9 1 10 9
17 13 9 8 8 9 9 1 0 9 13 1 9 7 1 9 9 2
33 7 13 2 2 8 14 8 0 9 2 2 0 1 7 9 13 1 9 9 1 9 0 7 2 14 13 0 9 1 10 9 2 2
3 7 13 2
20 2 14 1 9 1 9 7 15 9 15 13 1 9 1 10 9 1 9 2 2
54 7 13 8 1 9 0 1 9 8 8 8 8 1 9 9 12 2 12 0 7 9 14 13 9 15 1 9 9 7 12 9 7 15 13 9 0 7 2 9 13 1 15 1 9 0 3 1 9 9 12 2 2 2 2
11 2 7 15 0 1 10 9 2 2 2 2
20 2 8 8 1 9 1 0 9 1 0 9 7 9 1 9 7 8 9 2 2
74 7 9 1 9 1 15 13 9 9 9 9 9 9 0 7 9 15 1 9 2 13 8 2 2 8 8 8 8 1 9 7 9 3 1 9 9 9 1 9 9 7 9 1 9 7 9 9 1 9 14 13 1 9 1 9 2 8 8 8 7 8 1 9 9 0 1 9 9 9 1 10 9 2 2
22 7 13 7 15 14 13 9 9 9 1 9 9 7 14 13 9 1 1 9 15 10 2
45 1 9 0 2 13 9 0 1 9 0 8 8 9 12 2 12 1 8 9 0 1 9 9 7 0 0 1 9 0 1 9 15 9 1 9 15 1 9 0 1 8 1 9 0 2
11 9 0 13 9 12 1 9 15 1 12 9
79 13 9 0 1 9 9 0 9 12 2 12 0 1 9 9 9 9 1 9 1 9 9 9 9 9 15 13 1 12 9 1 9 12 0 2 7 9 0 1 12 9 13 0 1 9 1 9 9 2 7 9 9 0 1 0 1 9 7 9 0 15 1 9 9 7 9 7 9 9 2 7 13 1 9 9 9 9 0 2
68 7 13 9 8 8 1 9 0 0 1 9 14 13 10 9 7 13 15 9 8 8 9 9 9 1 9 7 9 9 0 1 9 9 9 9 7 13 8 8 1 9 9 9 9 9 0 0 1 7 13 9 9 8 8 1 9 1 9 13 1 15 9 9 9 1 9 9 2
43 7 13 0 0 1 9 9 1 7 9 0 7 0 1 9 9 13 9 9 0 9 12 9 0 9 9 0 1 9 9 9 7 9 9 0 1 9 7 15 13 9 9 2
7 9 0 13 9 9 9 0
22 13 9 0 0 7 9 13 1 9 9 7 13 9 0 13 12 12 9 1 9 0 2
34 7 13 9 1 9 0 0 10 9 1 9 9 0 15 9 9 1 9 0 1 9 12 5 1 9 1 9 9 7 9 9 1 9 2
34 7 13 9 1 9 9 9 1 9 1 9 9 0 1 9 9 0 1 9 12 12 9 0 7 13 1 12 12 9 1 9 9 0 2
28 7 13 7 9 9 0 0 1 9 13 1 9 12 9 7 13 1 1 12 12 7 12 12 9 1 9 0 2
16 9 9 9 0 7 9 15 14 13 1 9 9 7 9 7 9
3 0 2 2
46 13 9 9 8 8 7 15 14 13 2 9 0 2 15 13 15 9 9 0 9 0 1 9 9 15 7 7 9 9 15 1 0 9 0 7 0 13 9 7 9 9 15 7 9 15 2
59 7 13 9 8 7 0 0 1 9 9 9 0 15 8 8 8 13 9 2 7 7 0 2 1 9 9 15 1 9 9 7 13 9 1 9 15 1 9 15 9 15 1 9 1 9 8 9 1 9 9 7 9 9 8 8 9 9 0 2
31 7 13 9 9 0 2 15 13 1 9 1 9 8 8 8 2 9 8 8 9 1 9 9 7 9 9 8 1 9 15 2
94 7 13 9 9 8 8 1 9 15 9 9 9 9 0 1 1 8 9 9 1 15 7 9 9 15 7 9 7 9 9 15 13 9 15 1 12 9 0 14 13 9 0 7 13 9 12 1 15 9 12 2 12 0 7 15 8 8 8 9 2 8 8 8 8 2 8 8 8 9 9 8 8 8 9 0 9 7 3 9 1 9 8 8 7 9 15 9 1 9 0 7 9 0 2
40 2 2 9 9 9 9 9 2 1 9 15 2 13 8 9 9 9 9 9 15 13 1 12 9 0 2 0 1 7 3 9 0 14 13 9 15 1 9 0 2
13 7 13 2 2 14 9 0 0 7 14 13 2 2
15 0 1 7 1 9 9 1 9 9 7 9 0 7 0 2
25 2 2 0 0 9 2 7 13 8 1 9 0 15 13 9 0 1 9 0 15 13 1 9 0 2
34 2 2 9 9 9 2 7 14 13 9 9 1 9 7 9 9 9 0 1 9 9 0 1 1 9 13 9 1 9 0 7 9 0 2
8 8 8 2 9 9 9 9 0
35 13 8 8 9 0 1 9 9 0 7 9 2 9 9 2 13 1 9 1 9 7 9 0 1 9 9 0 9 1 9 0 1 9 0 2
65 13 8 1 9 8 8 1 9 9 15 13 1 15 8 1 9 9 7 0 1 9 9 2 7 13 9 0 1 9 0 7 0 9 13 1 9 0 1 9 10 9 15 13 1 9 9 9 14 13 1 9 1 9 0 2 7 13 9 9 0 1 9 9 9 2
16 0 1 7 15 1 9 9 9 7 14 15 14 13 1 15 2
13 9 9 9 9 2 9 9 1 9 8 8 1 9
14 13 9 9 9 9 1 9 9 8 8 1 9 2 2
8 1 9 9 0 1 9 2 2
27 7 9 9 9 9 1 9 9 9 8 8 7 9 0 1 15 1 9 8 1 9 1 9 0 7 0 2
17 7 13 9 9 9 0 0 1 9 12 1 9 9 9 9 2 2
19 7 13 1 9 9 0 1 9 9 9 7 9 9 1 9 9 0 2 2
25 9 0 1 9 0 8 2 9 9 9 2 7 15 14 13 9 15 1 9 1 9 12 9 0 2
15 13 9 7 9 9 8 8 8 9 9 1 9 0 2 2
15 7 14 13 0 9 0 7 0 7 0 1 9 0 2 2
15 7 14 13 9 9 7 9 1 15 1 9 9 0 2 2
10 1 9 8 9 15 1 9 0 2 2
19 7 1 0 7 15 9 9 9 1 9 0 14 9 7 9 1 15 2 2
12 7 13 9 7 15 13 9 0 7 0 2 2
18 7 9 0 1 9 9 13 7 9 9 8 8 8 7 9 0 2 2
10 7 15 14 13 1 9 7 9 2 2
14 7 14 13 8 9 9 0 7 0 1 10 9 2 2
6 7 1 15 9 0 2
9 9 9 2 15 1 9 9 2 2
9 7 0 1 9 0 7 9 2 2
63 13 8 2 8 8 8 9 9 9 0 1 9 1 9 0 1 7 15 0 7 9 7 13 9 15 9 9 8 0 1 9 9 7 9 9 1 9 1 9 14 1 9 15 2 7 13 2 14 15 13 1 9 9 15 7 15 9 2 9 2 9 2 2
64 7 13 9 8 1 9 13 1 15 1 9 2 9 9 2 1 9 0 13 9 9 0 9 15 1 9 1 9 0 2 7 13 2 7 13 9 13 7 9 9 1 9 2 7 10 9 0 7 0 7 13 8 8 0 9 7 8 15 15 9 10 9 2 2
24 0 1 7 9 13 8 1 15 7 13 13 13 1 9 1 9 9 7 8 1 9 15 2 2
90 7 14 13 9 9 9 1 9 15 1 9 0 0 2 8 2 1 9 0 2 7 13 2 7 8 8 8 8 9 13 0 7 9 0 7 8 8 7 8 8 7 13 1 9 7 0 8 1 15 2 7 13 9 0 0 7 0 7 7 13 9 15 8 8 8 1 15 8 8 8 2 0 1 7 9 13 8 1 15 7 13 13 13 9 0 7 13 1 15 2
15 7 13 9 9 9 15 1 9 9 0 1 9 7 13 2
14 7 8 8 1 9 7 14 13 7 8 7 15 0 2
43 7 13 8 2 8 7 13 14 13 1 9 8 1 9 7 9 7 13 7 8 13 15 9 7 9 9 15 2 14 8 8 8 7 8 0 7 13 9 1 9 1 9 2
36 7 13 9 8 9 15 0 1 8 8 7 9 15 15 13 15 1 9 1 7 13 9 9 0 1 0 0 7 9 15 15 13 1 9 9 2
25 7 13 9 9 1 9 15 1 9 1 9 0 7 7 15 13 9 0 1 8 8 7 13 9 2
39 7 13 8 2 8 1 9 9 15 13 15 9 9 9 9 0 7 13 1 15 9 0 15 13 1 9 1 0 7 13 2 14 8 13 1 9 8 8 2
56 7 13 9 9 9 15 1 10 13 7 15 14 13 1 9 0 7 13 2 14 8 8 0 13 15 9 7 9 8 8 8 8 8 8 8 2 14 8 9 1 9 2 7 13 0 1 15 2 14 3 9 9 0 1 15 2
16 7 13 1 9 1 9 9 2 14 13 8 8 7 14 8 2
57 7 13 9 9 1 15 13 1 9 9 9 7 13 1 9 0 2 2 6 1 9 2 2 7 7 13 15 9 1 9 0 9 1 9 7 13 9 15 1 10 9 13 9 9 2 2 7 9 9 0 8 1 9 8 2 2 2
6 12 5 1 9 9 9
35 9 9 15 13 1 9 9 0 2 14 9 7 13 1 9 15 9 0 7 0 2 7 0 15 9 2 9 2 15 13 13 9 0 0 2
129 7 14 13 9 0 1 9 9 9 7 9 7 9 9 9 1 9 13 1 12 5 1 9 9 2 7 7 13 9 0 9 9 9 9 2 7 14 15 13 1 9 12 9 9 9 2 7 13 9 9 1 9 1 12 12 9 2 1 9 12 12 9 1 9 0 2 7 1 0 7 15 1 9 0 13 9 12 9 1 9 2 7 13 0 12 9 1 9 2 7 0 13 12 9 1 0 2 1 9 13 1 9 1 9 9 9 1 9 2 7 15 10 13 15 9 1 9 9 8 7 9 9 15 2 9 1 9 0 2
41 7 13 9 7 12 5 1 9 9 1 9 0 1 12 5 3 9 9 0 2 7 7 13 9 1 9 7 14 13 9 15 13 1 15 9 9 9 15 1 9 2
12 9 0 13 1 2 9 2 13 1 9 9 15
71 13 9 0 9 12 2 12 0 1 2 9 2 14 13 15 9 0 1 9 0 2 7 13 1 9 9 9 9 7 9 9 9 2 7 9 9 1 9 1 9 9 2 7 9 9 0 2 7 9 9 2 2 1 9 9 0 2 1 9 9 1 8 7 9 9 0 0 1 9 0 2
41 13 1 9 2 9 12 2 12 0 9 2 9 9 1 9 12 2 1 9 9 0 1 9 7 9 9 0 7 0 7 0 7 9 7 9 9 9 0 7 0 2
17 7 13 9 9 1 9 1 2 9 9 9 0 2 7 13 9 2
28 7 13 9 9 9 1 9 0 2 8 8 2 1 9 15 13 15 9 2 1 9 9 9 2 1 9 0 2
50 7 13 1 9 13 15 1 9 7 9 13 0 1 9 1 9 1 9 9 9 0 7 0 7 9 9 9 1 9 0 2 1 9 1 9 9 9 0 1 9 2 9 1 9 9 0 0 1 9 2
35 7 13 8 7 9 9 9 7 9 7 9 7 9 0 2 7 9 9 1 9 8 8 2 14 13 1 9 9 1 9 0 1 9 0 2
105 7 13 7 9 2 13 1 9 9 2 1 9 9 2 9 0 2 1 9 9 0 2 1 9 0 7 0 7 9 9 0 13 12 12 9 13 1 9 0 1 9 0 2 9 1 9 9 9 2 7 9 0 1 9 7 9 14 13 1 15 14 9 0 0 2 9 1 9 0 0 1 9 2 10 13 9 1 9 1 9 1 9 9 0 7 8 7 9 0 2 1 9 1 9 9 9 2 15 13 9 9 0 1 9 2
43 7 13 1 9 9 15 13 15 9 1 9 12 1 9 0 2 15 13 1 9 9 9 1 12 1 12 1 12 7 9 1 12 1 12 5 2 9 1 9 9 9 9 2
54 7 13 7 3 9 0 1 9 0 15 13 1 9 9 0 2 4 1 9 3 7 7 1 9 9 0 2 2 1 15 9 15 13 15 9 9 0 7 9 9 7 9 1 9 2 1 9 1 9 12 2 9 2 2
40 1 9 15 2 13 9 9 9 0 1 9 2 8 8 2 7 9 13 0 9 0 1 9 2 7 7 15 13 1 15 13 1 12 5 1 9 0 1 9 2
35 7 13 7 9 12 5 1 9 0 0 1 9 9 0 13 1 9 2 2 7 15 9 14 13 0 14 13 1 9 9 1 9 9 2 2
10 9 7 0 13 1 9 0 1 9 0
18 1 9 1 9 0 8 1 9 9 2 13 9 0 8 8 7 13 2
14 8 8 9 9 9 1 9 2 1 9 9 1 8 2
44 8 8 1 15 13 15 9 0 0 0 13 9 9 0 1 9 12 12 9 1 9 9 1 9 7 9 9 1 12 9 0 1 1 15 9 13 9 7 9 0 1 9 0 2
68 7 13 9 9 9 1 9 9 0 1 9 9 1 10 13 15 10 9 0 7 14 13 15 9 0 1 10 9 7 9 9 9 1 9 0 7 9 0 7 13 9 9 9 9 1 9 9 9 1 9 0 1 9 9 9 7 9 9 1 9 9 0 1 9 1 9 0 2
21 7 13 9 1 9 1 1 10 9 15 13 9 9 0 1 9 0 1 9 0 2
15 7 13 9 0 7 9 9 9 1 9 9 0 1 8 2
42 8 8 1 9 9 9 0 1 9 0 1 9 0 1 9 9 9 1 9 1 9 0 7 9 9 1 9 0 13 9 0 1 9 9 0 13 9 0 1 9 9 2
59 7 13 9 9 9 7 9 0 0 13 1 9 9 13 9 0 1 9 7 13 9 15 0 1 9 0 0 1 9 9 1 9 7 9 0 7 9 9 9 1 9 0 2 0 9 0 2 1 9 15 1 9 9 7 9 7 9 0 2
10 8 8 2 9 13 9 13 1 9 15
31 13 9 9 0 8 8 7 9 15 13 9 13 1 9 9 13 0 7 0 2 0 1 2 9 10 13 9 9 9 2 2
20 7 13 8 1 9 0 1 9 0 2 7 9 9 8 15 1 9 15 2 2
22 7 15 13 1 7 9 9 7 9 0 7 9 0 2 1 9 9 9 9 0 2 2
35 7 13 1 2 9 1 8 9 7 9 15 1 9 0 2 2 0 7 2 9 9 0 15 9 0 7 0 7 0 7 4 0 3 2 2
34 7 13 7 9 9 2 15 9 0 1 9 2 2 0 1 7 0 1 9 1 9 7 9 9 7 9 2 13 1 9 9 9 2 2
19 7 13 7 9 13 1 1 12 12 9 1 8 9 8 8 9 9 12 2
13 9 0 13 9 0 1 9 9 0 7 9 9 0
39 13 9 0 1 9 9 9 0 1 9 9 9 0 0 15 13 15 1 9 0 7 13 9 15 2 7 13 1 9 9 15 1 9 13 9 9 1 15 2
33 7 13 9 9 0 1 9 9 0 2 7 13 7 13 1 0 7 13 1 9 0 2 7 15 14 13 9 0 9 1 9 9 2
18 7 13 9 0 9 15 1 9 9 1 9 7 9 9 0 1 9 2
24 7 13 1 9 10 1 7 8 7 13 1 9 0 9 0 1 9 10 9 7 15 1 9 2
59 7 13 9 1 9 9 9 2 8 8 0 9 9 1 10 9 1 9 8 9 1 9 0 1 15 7 15 9 9 1 9 12 1 12 1 0 1 9 0 7 13 10 9 1 12 5 1 9 15 13 1 15 1 9 0 1 9 0 2
112 7 13 10 9 1 9 9 1 9 0 2 7 13 8 9 9 0 0 9 8 8 8 2 7 9 9 0 13 9 15 1 9 9 1 9 0 1 9 2 7 7 14 13 7 14 9 13 9 1 9 1 9 2 7 7 13 13 1 9 15 0 9 7 14 13 1 15 1 9 9 0 2 15 1 9 0 9 1 9 9 9 9 7 9 9 7 9 0 1 9 9 0 7 15 10 13 1 15 9 1 9 0 2 7 13 9 0 1 9 9 9 2
64 2 2 9 0 7 13 8 1 7 15 1 0 1 9 10 9 7 14 13 9 1 9 0 9 15 7 9 0 1 10 9 7 7 1 15 7 13 9 0 1 9 9 1 9 0 1 10 13 1 15 1 9 1 9 9 9 7 9 9 7 9 9 0 2
54 7 15 13 15 9 1 9 15 7 13 2 1 9 9 9 9 10 13 1 15 1 9 2 1 9 9 0 9 7 15 13 1 15 1 9 0 1 9 12 7 13 1 8 9 9 0 1 10 13 9 15 12 9 2
23 7 1 9 7 9 14 13 2 8 7 9 14 13 9 7 9 14 13 1 9 1 15 2
95 7 13 7 13 9 9 1 9 9 9 0 7 14 13 1 9 9 0 2 9 7 9 15 1 9 9 9 0 0 14 13 1 9 1 9 0 1 9 2 7 7 15 14 13 1 9 0 1 9 9 0 7 7 3 14 13 1 9 9 1 9 0 1 9 9 1 9 9 0 0 2 7 14 9 15 1 9 0 9 0 1 9 9 1 9 0 0 1 9 1 9 1 10 9 2
19 7 1 15 13 9 1 9 9 9 0 15 9 0 9 2 7 0 9 2
9 0 9 1 9 0 1 9 7 8
26 13 9 0 0 0 0 9 1 9 9 9 0 1 9 9 9 1 9 0 0 7 0 9 1 8 2
22 13 9 0 1 9 0 9 2 8 2 1 12 9 1 9 9 0 0 9 1 8 2
17 13 8 9 13 9 9 9 9 3 9 9 0 15 13 9 15 2
19 13 9 0 0 9 9 9 9 7 9 0 1 9 9 1 9 9 0 2
28 13 9 1 7 9 0 13 9 1 9 1 8 2 9 2 0 1 9 1 9 9 15 1 9 0 1 9 2
19 7 1 0 7 13 9 0 1 9 9 0 9 1 9 8 0 1 15 2
33 7 13 9 9 9 1 9 9 9 7 9 0 14 13 9 2 8 8 2 1 8 0 0 1 9 7 15 13 9 0 1 9 2
25 7 13 9 9 1 9 9 9 0 1 9 9 0 2 8 8 2 7 8 1 9 1 9 0 2
6 8 13 9 0 1 9
17 13 9 9 0 1 9 7 8 1 9 0 1 9 1 9 9 2
47 13 9 8 8 9 9 9 1 9 9 0 15 13 9 9 12 2 12 0 1 9 9 1 9 9 1 9 9 1 9 9 1 9 1 9 9 1 9 9 8 1 9 15 1 9 0 2
14 9 9 0 13 1 9 0 7 0 1 9 9 15 0
97 13 9 9 0 0 7 0 15 13 9 15 1 9 0 1 9 0 1 1 12 12 9 1 9 9 15 1 9 0 14 3 9 9 9 0 7 8 7 8 7 3 8 0 1 9 1 9 0 1 9 9 15 0 7 9 9 0 7 9 1 8 9 7 15 13 1 9 9 7 9 0 1 12 9 7 13 8 1 9 0 0 1 9 0 1 9 9 9 9 8 9 9 7 9 7 9 2
45 7 13 9 9 9 0 9 8 8 7 9 9 15 13 15 9 0 1 9 9 7 0 12 5 13 1 9 9 9 9 0 9 7 9 9 9 9 9 13 1 9 10 9 0 2
55 7 13 1 7 9 0 9 0 1 9 9 7 9 9 1 9 9 1 9 0 8 8 1 9 0 1 9 9 9 7 1 15 9 13 1 9 9 0 9 8 9 9 0 0 1 9 9 9 0 7 9 0 7 0 2
65 7 13 7 9 0 0 1 9 0 1 9 7 9 13 1 9 9 0 1 8 8 7 9 7 9 7 9 7 9 7 8 1 9 1 12 12 9 2 12 8 9 2 7 1 0 7 13 9 9 0 1 9 0 0 1 1 12 8 9 2 12 8 9 2 2
51 7 13 7 9 1 9 9 9 14 13 1 9 9 9 0 7 13 7 9 0 1 9 13 9 1 9 9 0 1 9 0 1 9 1 9 0 1 7 9 13 1 9 0 9 15 13 9 1 10 9 2
60 7 1 9 0 13 9 0 0 1 9 0 0 1 9 12 12 9 1 15 9 1 9 9 1 9 0 1 9 9 15 12 12 9 7 9 1 9 8 0 1 9 1 9 1 9 12 5 12 9 1 9 0 7 12 12 9 1 9 0 2
12 7 13 9 0 1 9 9 0 1 9 9 2
39 1 15 13 9 9 7 9 0 1 9 9 15 15 13 1 1 9 1 9 1 9 0 0 1 15 13 1 9 9 9 1 9 0 0 1 9 9 0 2
44 7 13 9 9 9 1 9 0 0 0 1 9 9 7 9 7 9 7 9 1 9 9 9 0 0 9 7 9 7 9 1 9 7 3 9 0 1 10 9 1 9 9 0 2
57 7 13 9 1 9 9 7 9 7 9 9 1 9 1 9 0 1 9 9 0 13 9 0 7 0 13 9 0 1 9 9 0 7 9 9 9 0 1 10 9 7 9 9 9 9 7 9 0 1 9 9 7 9 0 1 15 2
76 7 13 9 9 9 9 9 9 1 9 9 0 9 8 8 1 7 9 0 9 14 13 1 12 9 0 9 1 9 9 9 7 9 0 1 9 9 9 10 9 1 9 9 0 14 3 7 10 9 0 1 9 0 0 0 1 9 9 7 9 9 0 7 9 15 1 0 7 13 15 9 9 0 9 0 2
38 7 13 8 1 9 14 13 8 8 1 9 9 0 7 9 0 1 9 9 7 9 14 13 8 8 9 0 1 9 0 1 9 9 0 1 9 0 2
10 9 9 9 9 9 13 9 9 1 9
16 13 9 1 9 7 9 9 9 1 9 9 9 9 9 9 2
32 13 9 9 9 9 9 9 9 0 1 9 9 7 9 7 13 9 0 1 9 13 1 9 9 9 9 0 9 1 0 9 2
23 13 10 9 1 9 9 9 7 9 7 9 9 1 9 0 1 9 1 9 7 9 0 2
39 1 9 0 13 9 0 1 9 9 9 9 0 1 9 1 9 9 9 9 9 9 9 7 9 9 9 9 0 1 9 1 9 9 15 13 15 9 0 2
27 7 13 9 1 9 9 9 0 1 9 9 9 15 13 9 7 9 9 9 0 1 9 1 9 9 9 2
33 7 13 1 9 9 9 0 15 13 1 9 8 1 9 9 0 7 9 9 13 1 9 9 9 7 9 9 9 1 9 9 0 2
32 13 7 9 8 8 9 9 14 13 1 9 9 1 9 1 9 9 0 7 15 14 13 9 13 9 1 9 9 1 9 9 2
36 7 13 9 9 1 9 9 9 9 9 1 9 7 0 9 1 9 1 9 9 9 15 13 9 9 1 9 9 9 0 1 9 9 9 0 2
5 9 0 1 9 0
62 13 9 8 8 9 9 7 9 0 7 9 13 9 9 1 9 9 0 9 7 0 0 7 15 13 15 13 1 12 5 1 9 9 0 1 10 9 7 9 0 0 15 13 1 12 5 8 8 9 9 12 5 9 1 9 9 0 0 1 9 8 2
58 13 8 2 8 1 9 0 9 12 2 12 7 9 0 13 9 0 1 9 0 1 15 13 1 15 1 9 0 0 1 7 15 1 9 9 0 1 9 9 7 9 9 1 9 9 7 15 13 9 0 1 9 1 9 7 9 9 2
9 8 2 9 0 1 9 0 7 0
68 13 8 2 8 8 8 9 9 0 7 15 13 9 12 2 12 0 9 1 9 1 9 9 8 1 9 9 0 1 9 13 9 0 9 1 9 1 9 7 9 7 9 0 1 10 13 1 9 0 7 9 0 7 9 9 7 9 1 9 1 9 9 0 1 9 7 9 2
27 13 8 1 9 8 2 8 1 8 8 8 9 0 1 9 8 7 15 13 0 9 1 9 0 1 8 2
62 7 13 7 9 9 10 9 13 1 9 0 9 1 9 1 9 0 15 13 15 7 9 9 7 9 7 9 9 7 13 7 15 13 9 1 9 9 1 9 9 0 1 9 9 0 1 9 9 9 1 9 9 0 1 9 9 1 9 1 10 9 2
81 7 13 8 2 8 7 9 1 9 9 7 9 8 1 10 9 14 13 9 0 1 9 9 0 1 9 8 7 9 15 0 7 15 7 13 9 8 0 9 1 8 9 0 7 13 9 15 1 9 0 7 14 15 1 9 13 9 0 9 0 1 8 9 0 7 13 1 9 9 1 9 1 9 0 7 13 9 0 1 9 2
43 7 13 8 2 8 7 15 13 15 9 1 9 0 1 9 9 15 9 9 0 1 9 1 9 7 9 7 9 9 1 9 13 1 15 13 15 9 0 1 9 9 0 2
39 7 13 9 1 9 9 1 9 1 9 9 7 9 8 13 1 9 15 9 9 7 9 1 9 0 7 9 9 0 1 9 1 9 1 9 9 1 15 2
58 1 9 0 13 8 7 15 13 0 9 9 1 9 0 7 0 1 9 10 9 1 9 9 9 0 7 0 0 1 7 1 0 9 10 9 15 9 1 9 9 7 9 1 10 13 1 9 9 0 1 0 9 1 9 1 9 0 2
57 7 13 8 2 8 1 7 15 13 0 9 1 9 9 9 0 0 1 9 9 8 1 9 9 0 1 9 0 1 10 9 7 9 9 0 1 9 1 9 0 1 10 9 7 9 7 9 0 15 13 7 13 9 1 10 9 2
9 9 9 13 1 9 0 1 9 9
49 13 9 9 7 9 1 9 9 1 9 0 1 9 12 12 7 12 12 8 1 9 9 9 9 8 1 9 9 7 13 9 8 8 9 9 7 9 7 9 13 1 9 9 1 9 9 1 9 2
51 7 13 9 7 9 9 14 13 1 12 5 1 9 0 1 9 0 7 15 9 13 0 7 14 15 0 9 1 10 15 0 1 9 9 2 7 7 0 15 7 13 10 9 1 12 5 1 9 9 12 2
28 7 13 9 8 8 1 9 7 9 14 13 1 9 9 0 1 9 1 12 8 0 1 12 8 1 9 12 2
74 7 13 9 8 1 7 13 9 9 1 9 0 1 9 8 1 9 9 0 7 0 2 7 13 9 9 12 9 1 9 9 12 9 7 13 9 9 1 12 5 0 7 9 9 8 9 1 9 9 9 9 9 9 2 7 13 9 0 9 9 9 0 7 3 9 9 7 0 9 0 0 1 15 2
24 7 13 9 0 9 9 1 9 9 0 7 9 0 1 9 1 10 13 1 9 7 9 15 2
12 12 12 9 1 9 12 9 1 9 0 1 9
44 13 8 2 8 8 9 9 0 1 9 9 7 15 13 0 9 9 0 1 9 12 9 1 9 0 1 9 1 9 12 12 7 12 12 9 2 1 15 12 12 9 9 0 2
20 13 15 1 9 9 9 0 7 9 1 9 8 2 9 8 9 9 7 9 2
42 13 8 1 7 9 0 1 9 12 9 2 7 13 9 15 12 12 7 12 12 9 2 7 1 0 9 9 15 0 1 9 0 2 7 9 15 0 1 0 9 0 2
32 7 13 8 7 9 9 13 1 9 9 0 0 1 9 12 12 7 12 8 1 9 12 12 9 1 15 12 12 9 9 0 2
4 9 9 9 9
20 13 9 9 9 1 9 9 9 0 1 9 9 7 9 1 9 7 9 0 2
50 13 9 8 8 9 9 9 7 15 13 9 2 12 2 12 9 9 7 9 0 1 9 1 9 9 7 9 9 9 7 9 7 13 7 9 9 15 13 9 1 9 15 13 0 8 8 9 1 9 2
50 7 13 7 15 13 9 9 0 1 9 2 12 2 12 9 9 1 9 1 9 9 9 0 7 9 9 9 1 9 7 13 1 9 2 12 2 12 9 1 9 9 7 9 0 0 1 9 7 9 2
19 7 13 7 9 0 13 9 15 0 1 9 1 9 9 9 1 9 0 2
33 7 13 9 1 9 1 2 9 2 7 9 13 1 15 0 2 12 2 12 9 9 13 9 1 15 1 9 9 8 9 1 9 2
17 9 0 13 9 9 9 9 0 1 9 0 7 13 1 9 9 15
20 13 9 0 9 9 9 1 9 0 1 9 0 1 9 9 9 9 12 9 2
59 7 13 9 15 13 15 9 9 9 9 0 7 9 1 9 2 9 7 9 0 1 9 12 2 9 9 1 9 7 9 0 7 13 9 1 9 15 0 15 13 1 9 15 7 9 15 7 3 9 9 15 0 1 9 9 7 9 0 2
42 7 13 9 10 9 1 9 1 9 9 9 0 0 15 13 9 0 1 9 0 1 9 7 9 0 1 9 15 1 9 9 0 0 15 13 9 9 0 1 10 9 2
136 7 13 9 1 7 9 9 1 9 9 0 1 9 0 0 14 13 9 0 2 9 15 13 9 9 1 9 9 9 0 0 1 9 9 9 15 13 15 8 1 10 9 2 7 13 9 7 13 0 1 9 9 1 9 7 9 0 1 9 9 1 9 8 0 1 9 9 0 9 9 0 2 7 3 7 13 10 9 1 9 0 1 9 9 9 0 8 7 9 0 1 9 9 9 15 13 15 1 9 9 15 0 2 0 7 9 9 9 9 0 0 1 9 1 9 0 13 15 9 1 10 9 2 7 13 9 15 1 9 9 9 0 1 9 0 2
103 7 13 9 7 15 1 0 7 13 9 9 7 9 0 1 9 7 9 0 9 0 9 9 0 12 1 9 10 13 1 9 9 15 13 13 9 0 1 9 1 9 9 9 0 7 8 2 0 7 10 9 14 13 9 9 0 1 10 9 0 12 9 1 1 12 5 7 13 15 1 0 9 7 9 0 2 9 15 13 9 15 1 9 14 9 15 1 9 9 15 13 9 9 9 1 9 0 9 1 9 9 0 2
109 7 13 9 7 9 9 9 0 1 9 9 7 9 0 14 13 9 9 9 0 1 9 0 1 10 9 7 14 13 9 9 0 14 3 9 1 9 9 0 1 15 9 0 7 9 15 14 13 1 9 9 9 15 15 13 9 0 1 9 7 9 7 9 7 9 7 9 0 0 1 9 9 0 2 9 15 13 1 9 9 9 9 9 0 7 9 15 1 9 0 7 0 1 9 9 9 7 9 0 1 9 0 1 9 7 0 1 9 2
58 7 13 9 7 9 9 0 0 1 10 9 0 0 13 3 9 9 1 9 15 13 9 0 7 0 1 10 9 1 9 7 9 9 0 7 3 8 0 7 10 9 14 13 9 0 1 9 0 7 13 1 15 9 0 1 9 0 2
58 7 13 9 1 9 9 9 7 9 0 7 9 9 0 1 9 0 7 9 9 1 9 9 8 1 9 8 9 0 1 9 9 15 0 2 0 7 9 9 9 0 7 9 1 9 9 0 1 9 0 12 5 9 0 1 10 9 2
7 9 0 1 9 1 9 9
34 13 9 9 9 0 7 0 0 9 9 0 1 9 9 1 9 9 7 9 1 9 9 9 0 1 9 0 13 1 1 12 12 9 2
32 13 9 8 8 9 9 7 9 9 1 9 9 9 0 13 1 1 12 5 7 13 14 12 5 0 1 12 9 1 9 9 2
23 13 8 1 7 9 1 9 9 0 15 9 9 1 9 9 7 9 9 0 1 9 0 2
70 13 8 1 7 9 0 1 9 0 14 13 9 1 9 12 1 9 12 12 9 1 9 9 0 7 13 9 1 9 9 0 1 9 9 9 9 1 9 8 1 9 12 7 1 9 0 12 12 9 1 9 1 9 9 0 2 7 13 9 9 0 1 9 9 1 9 9 15 0 2
27 7 13 7 9 0 1 9 7 15 0 1 9 9 0 14 13 9 1 9 0 1 9 12 12 9 0 2
31 13 8 7 9 0 14 13 9 15 1 9 9 9 7 9 9 9 12 1 9 12 2 7 15 13 9 12 9 9 0 2
27 7 13 8 9 0 1 9 12 9 0 1 9 1 9 2 0 7 12 9 13 3 1 9 0 7 9 2
29 0 7 7 3 9 1 9 9 13 9 15 1 0 1 9 1 9 0 7 15 15 13 9 9 0 1 9 2 2
12 7 9 9 15 14 13 9 15 1 9 0 2
14 12 12 9 1 9 9 9 0 1 9 0 1 9 9
45 13 9 9 9 0 9 9 9 9 0 9 1 9 9 8 8 9 9 2 7 13 9 9 9 9 1 9 0 12 2 12 7 9 9 12 12 9 1 9 9 1 9 0 0 2
35 7 14 13 9 9 9 9 9 9 0 0 1 9 1 9 0 7 13 1 9 0 9 0 1 9 9 0 1 9 9 1 9 9 0 2
68 7 13 9 8 8 7 15 13 9 9 0 0 1 9 9 13 1 9 1 9 1 9 9 1 9 15 1 9 9 0 15 13 9 15 0 1 9 9 2 7 13 9 9 1 9 1 9 9 1 9 1 9 9 1 9 1 10 13 15 9 0 1 9 7 9 1 9 2
43 7 13 9 9 9 1 9 0 1 9 9 1 0 9 7 7 13 9 9 9 1 9 1 9 9 13 1 10 9 1 9 0 1 9 1 9 15 13 9 1 10 9 2
44 13 9 1 7 9 9 15 13 9 9 15 1 9 8 8 9 9 9 9 0 8 8 1 9 7 9 9 7 9 2 1 9 1 9 12 9 0 1 9 9 0 7 0 2
10 9 2 8 0 2 13 9 8 1 9
53 13 9 9 9 9 0 9 12 2 12 0 1 9 9 1 9 9 15 13 9 8 7 13 15 1 9 9 9 9 9 9 1 9 9 0 1 9 9 1 8 8 0 8 13 12 5 1 9 0 0 1 9 2
69 7 1 9 15 13 9 8 8 9 9 9 9 9 7 9 9 1 9 0 2 1 9 9 2 7 15 14 13 9 9 8 8 9 9 0 1 9 0 1 9 1 8 9 9 7 9 1 9 1 9 0 1 7 15 13 1 9 0 1 9 15 1 9 9 9 9 8 8 2
65 7 13 8 8 8 9 9 9 9 9 8 7 9 13 1 9 15 14 13 15 9 7 13 15 1 7 15 13 9 0 1 9 9 8 1 9 0 8 8 0 15 13 9 1 9 9 0 2 1 9 9 10 9 1 9 9 0 15 13 1 9 9 15 2 2
23 7 15 9 15 13 9 7 1 9 1 9 15 13 15 10 9 7 9 1 9 1 9 2
101 7 13 1 7 9 8 1 9 0 1 9 9 0 9 9 1 9 8 8 8 1 9 12 9 12 1 9 12 2 12 0 1 9 1 9 9 0 0 0 1 9 8 0 1 9 9 7 14 13 9 1 15 1 9 7 15 15 13 15 1 9 0 2 7 13 0 1 9 9 1 9 14 13 9 1 15 7 13 15 1 9 9 7 13 7 15 13 9 9 1 9 9 7 9 9 9 0 7 9 0 2
52 7 7 13 9 8 8 7 13 0 1 9 0 8 8 14 13 1 9 13 1 9 1 7 15 13 9 13 7 13 9 15 1 9 7 1 1 9 0 1 7 9 14 13 2 1 9 9 15 2 1 9 2
12 12 5 9 1 9 9 1 9 0 1 12 9
45 13 9 1 9 9 0 1 9 9 1 9 7 9 0 7 9 1 9 9 0 1 9 9 1 9 9 1 9 9 0 1 9 7 15 13 1 9 12 5 1 12 9 0 2 2
13 1 9 9 9 0 1 9 7 9 0 1 8 2
40 13 9 0 1 7 9 8 8 9 9 9 14 13 1 9 9 9 0 1 9 9 12 2 12 0 1 9 9 9 0 7 9 0 1 9 1 9 9 9 2
66 13 9 7 8 2 8 14 13 1 9 9 0 9 9 1 9 0 1 9 9 9 1 9 9 9 7 9 9 7 9 15 13 15 9 1 9 9 1 9 9 0 0 7 0 1 9 9 9 9 9 7 9 9 0 7 9 9 7 9 1 9 9 7 9 9 2
46 13 9 8 1 9 15 1 9 9 9 0 9 9 9 1 9 7 9 15 7 9 0 0 1 9 7 9 9 1 9 9 1 9 0 15 13 12 5 1 9 9 0 1 9 2 2
16 7 9 9 1 9 0 7 9 1 9 0 1 9 0 0 2
31 13 8 2 8 14 13 1 8 8 9 9 0 1 9 15 1 9 1 9 0 9 9 9 0 1 9 9 15 1 9 2
52 13 9 7 15 13 0 9 9 1 9 9 9 7 9 0 1 9 13 9 0 12 5 1 15 1 9 0 1 12 5 1 9 1 9 0 1 9 1 9 0 1 9 0 1 9 0 1 9 12 12 9 2
50 7 1 9 9 9 9 13 9 9 9 0 1 9 9 1 15 12 9 1 9 9 9 7 9 1 9 0 1 12 9 0 1 9 9 7 9 7 9 7 9 0 7 9 1 9 9 0 1 8 2
12 9 0 0 1 9 0 7 9 9 0 1 8
39 13 9 12 2 12 0 9 8 8 9 9 7 9 0 1 8 8 9 9 9 7 9 0 9 9 0 1 9 7 9 9 1 9 9 0 1 9 0 2
42 7 13 8 7 10 9 13 1 9 9 9 1 9 7 9 0 7 9 9 1 9 0 7 13 9 0 1 9 1 9 0 1 9 9 9 0 1 9 9 9 0 2
106 7 1 9 15 13 9 9 9 7 9 0 7 10 9 1 9 10 13 9 15 7 9 1 15 1 9 9 9 7 9 9 9 1 9 15 0 1 9 2 0 1 7 9 13 4 3 9 9 1 9 9 0 1 9 2 7 7 3 1 9 1 9 0 1 9 1 9 13 1 0 0 7 13 9 9 2 7 13 1 9 9 15 1 9 1 9 1 9 7 9 9 0 9 7 9 0 7 9 9 7 9 7 9 7 9 2
109 7 13 9 8 7 9 13 8 9 0 1 9 2 8 8 13 1 9 9 9 7 9 15 1 8 8 7 9 9 0 1 9 0 2 7 9 9 9 9 1 9 9 9 13 0 7 0 2 1 9 1 9 9 9 8 8 9 9 7 9 9 1 9 9 9 0 1 9 1 9 7 9 7 9 0 7 9 1 9 8 7 9 7 9 0 1 15 7 9 9 7 9 9 7 9 0 1 15 7 9 9 9 7 9 0 7 9 15 2
69 7 13 1 7 15 13 9 1 9 0 1 9 9 1 9 9 8 8 2 0 1 9 9 9 7 9 9 0 8 0 7 9 9 7 9 7 9 9 0 2 3 1 9 9 0 1 10 1 9 9 1 9 0 1 10 9 2 7 13 9 1 15 1 9 9 0 1 9 2
11 9 0 2 0 1 9 9 9 7 9 9
24 13 9 8 8 9 9 1 8 8 8 9 9 7 9 0 9 9 9 1 9 1 9 9 2
36 13 9 7 3 9 0 1 9 9 7 14 13 9 0 9 1 9 9 9 9 0 7 9 0 0 2 7 9 1 9 9 7 9 9 9 2
44 13 9 0 7 9 9 0 1 9 9 9 7 9 9 7 9 9 9 7 9 9 13 9 0 2 7 13 1 9 15 1 9 9 0 1 9 0 0 1 9 9 1 9 2
15 9 9 1 8 0 1 12 9 7 9 9 1 12 12 9
34 13 9 9 0 1 9 0 7 9 1 9 9 0 1 8 1 0 1 12 9 7 13 12 12 9 3 1 12 9 1 9 9 0 2
54 7 13 9 1 9 9 1 9 0 13 12 12 9 7 13 9 15 1 12 12 9 1 9 1 9 1 9 9 12 9 1 9 0 1 9 12 7 15 13 1 15 9 9 12 12 9 7 13 9 12 12 9 3 2
130 13 7 9 0 13 9 1 9 1 8 1 7 9 0 13 1 9 9 2 7 13 9 9 8 8 9 9 9 9 9 0 1 8 1 9 0 9 1 9 9 7 9 0 1 9 0 7 15 10 13 15 9 9 1 9 0 7 15 13 1 9 9 0 7 9 9 9 0 1 9 9 15 13 1 9 9 9 1 9 9 9 9 1 9 1 9 9 1 9 7 9 9 0 0 2 7 13 9 9 0 9 1 9 7 1 9 9 9 0 2 0 2 9 1 7 9 0 1 9 14 13 1 9 9 1 9 0 1 9 2
18 9 8 0 1 9 2 9 9 9 0 1 9 1 12 12 9 9 12
40 13 9 8 8 8 9 8 0 1 9 7 9 9 0 1 9 15 7 9 13 1 12 12 9 1 9 12 1 9 13 9 15 12 5 1 15 1 9 0 2
27 7 13 1 9 1 2 9 2 7 9 9 0 1 9 7 8 14 13 1 1 12 12 9 1 9 0 2
43 7 13 7 9 9 9 7 9 0 8 8 8 1 9 7 9 15 1 9 8 8 7 9 15 1 9 0 13 9 0 1 9 9 0 1 9 9 7 9 9 9 15 2
31 7 13 1 10 9 1 7 9 9 13 1 9 0 1 9 9 8 8 1 8 0 9 12 7 13 9 9 0 1 9 2
53 7 13 1 9 0 1 9 0 1 9 7 15 13 1 9 0 0 1 12 12 9 7 15 9 9 1 9 1 9 0 1 9 0 15 13 1 9 0 0 7 9 1 9 9 1 9 7 9 1 9 9 0 2
53 7 13 9 0 7 3 9 1 9 9 0 1 9 1 9 2 7 9 1 9 0 1 9 15 7 13 9 9 0 12 9 0 9 1 9 15 13 1 15 12 1 9 9 1 9 9 9 0 7 0 1 9 2
45 7 13 7 9 0 14 13 8 1 9 1 12 2 12 9 0 1 9 9 0 0 1 8 7 15 14 13 1 9 9 0 1 0 7 9 15 1 9 0 7 9 9 1 9 2
77 7 13 7 9 9 13 9 0 1 9 1 9 7 8 15 13 9 9 15 7 9 15 0 7 0 7 13 9 9 9 1 10 9 2 0 1 7 9 1 9 15 9 8 0 1 15 9 9 1 9 0 1 9 9 9 9 9 2 7 7 8 1 9 0 1 9 9 15 1 9 1 9 9 0 1 9 2
47 7 13 1 10 9 1 7 9 9 7 9 0 9 8 8 8 14 13 9 9 12 7 12 9 0 1 9 9 9 9 1 9 1 9 8 9 7 9 9 9 15 13 15 8 1 9 2
7 9 9 9 0 0 9 0
40 13 9 8 8 8 9 9 0 7 9 0 1 9 15 7 9 14 13 9 2 0 2 1 1 9 1 9 0 2 1 9 2 7 9 9 0 1 10 9 2
46 7 13 1 9 0 1 9 15 1 9 8 8 9 9 9 7 9 9 1 9 0 7 9 0 7 9 7 15 13 9 1 9 1 9 7 9 1 9 9 7 9 7 9 7 9 2
60 7 13 7 9 9 0 13 1 9 0 9 1 9 0 1 9 0 0 8 7 13 9 1 9 0 2 0 1 9 9 1 1 9 1 9 9 8 1 9 1 9 2 0 1 7 9 14 13 1 15 9 15 12 12 9 9 1 9 0 2
44 7 13 7 9 7 9 14 13 1 9 9 0 1 9 9 1 9 7 9 9 1 9 1 1 9 0 1 8 8 7 9 0 2 9 1 9 9 1 9 9 9 7 9 2
46 7 13 9 0 7 8 8 9 9 0 14 13 9 9 9 0 1 9 9 9 1 9 7 9 1 9 9 9 0 2 0 1 9 9 0 1 9 1 9 9 9 7 9 9 0 2
10 9 1 9 9 7 9 1 9 7 9
64 13 8 8 9 9 9 0 1 9 9 9 8 13 9 0 7 9 15 13 9 0 1 9 9 9 0 1 9 1 9 9 7 9 15 13 13 1 1 15 9 9 1 9 2 7 13 7 15 14 13 9 1 9 0 7 9 15 1 9 1 10 9 9 2
56 7 13 8 1 9 0 1 9 0 1 9 1 9 7 9 1 9 9 1 1 15 9 9 9 7 13 9 9 1 0 0 0 1 9 2 7 7 13 9 0 1 9 7 9 1 9 9 0 1 9 9 0 1 9 0 2
50 7 13 8 7 9 9 9 1 9 9 13 12 12 9 7 12 5 1 15 1 9 9 7 13 9 0 1 12 5 1 9 9 8 0 7 12 5 1 9 7 12 5 1 9 9 9 0 1 9 2
88 7 13 9 9 1 9 7 9 9 9 0 1 9 9 12 7 12 7 15 9 0 1 9 0 7 9 1 15 9 1 9 10 9 1 9 7 0 0 1 9 9 9 0 1 9 9 1 9 9 1 9 1 9 1 9 0 9 9 9 0 1 7 9 9 9 0 9 8 8 8 0 1 9 0 0 1 9 9 0 1 9 1 9 1 9 12 9 2
37 7 13 9 9 0 9 1 9 9 9 0 1 9 8 8 1 9 1 9 9 0 1 9 0 9 15 1 9 1 9 1 12 1 12 9 0 2
11 9 9 0 13 1 9 9 1 9 9 9
70 13 9 9 0 0 2 8 2 9 12 2 12 0 1 9 9 15 15 13 1 8 9 15 1 9 9 9 1 9 9 9 0 1 9 9 9 9 7 13 9 0 1 9 15 0 15 13 9 12 2 12 0 9 0 15 13 15 9 1 9 0 7 1 9 0 9 1 10 9 2
37 7 13 9 8 8 2 9 9 9 9 9 9 9 2 15 13 9 0 1 9 2 8 2 1 8 7 9 14 13 9 0 1 9 9 9 9 2
150 7 13 7 10 9 13 1 9 9 9 0 15 13 1 9 9 0 15 13 9 9 0 7 9 0 13 9 0 7 15 0 9 0 1 9 9 2 7 13 10 9 9 9 0 1 9 9 0 2 7 13 9 8 7 9 0 13 7 13 9 9 0 1 9 9 0 9 9 2 7 0 13 9 0 1 9 0 1 9 0 7 9 9 1 9 1 9 1 9 9 0 13 9 9 9 9 7 9 0 0 7 9 1 9 0 7 9 0 7 9 0 0 2 13 1 15 9 15 0 7 13 9 8 7 9 9 0 14 13 9 9 0 1 9 9 14 12 9 1 9 0 9 1 9 15 1 9 0 0 2
23 7 13 9 2 8 2 14 13 9 1 9 9 9 0 1 9 9 9 1 9 9 12 2
17 7 1 10 9 13 9 9 0 1 9 9 9 15 1 1 9 2
39 7 1 9 9 13 9 8 1 7 9 13 9 1 9 9 9 0 1 9 9 9 2 13 9 9 0 7 9 8 2 7 13 7 9 13 0 9 0 2
8 0 9 0 0 2 1 9 9
36 13 9 9 9 15 13 9 12 9 0 1 9 9 9 9 0 1 9 0 7 0 1 9 7 9 9 9 0 1 15 1 9 12 12 9 2
48 13 1 15 2 1 9 9 2 8 8 9 9 9 7 13 7 15 14 13 9 9 0 1 9 9 0 7 0 7 9 7 9 7 9 0 7 0 1 9 15 14 13 1 10 9 1 9 2
37 7 13 8 8 7 3 12 9 9 0 14 13 1 9 2 7 13 1 9 15 9 1 9 0 1 9 2 3 1 9 9 2 1 9 9 9 2
100 7 1 0 15 14 13 9 9 0 1 9 0 1 9 7 9 9 9 9 9 0 7 9 9 9 0 7 9 9 8 1 9 7 9 0 9 9 0 7 9 9 9 0 8 8 7 9 9 9 8 2 7 14 13 3 1 9 9 0 9 0 1 9 7 15 8 8 7 15 13 1 9 1 9 9 0 0 2 12 9 2 7 3 9 7 9 7 9 7 9 0 7 9 9 0 7 9 7 9 2
27 1 9 0 14 13 12 9 0 3 1 15 9 9 0 7 9 7 9 7 9 7 9 7 9 7 9 2
18 7 13 8 8 7 3 0 1 12 9 1 9 14 13 1 9 9 2
8 9 0 1 9 9 1 8 0
82 13 9 0 1 9 9 0 0 1 9 0 1 9 9 9 0 0 1 9 1 8 8 8 0 7 0 12 5 7 13 7 13 10 9 1 9 1 9 0 1 9 9 0 1 9 9 7 9 15 13 9 1 15 1 9 9 9 0 0 9 8 8 8 1 9 9 0 7 13 9 9 9 9 0 7 0 1 9 1 12 9 2
53 7 13 9 7 9 9 0 13 1 9 0 0 1 9 9 0 1 9 0 7 0 7 0 1 9 7 9 13 9 1 9 0 1 9 9 1 9 2 1 1 9 0 1 9 9 7 9 7 9 9 7 9 2
36 7 13 7 9 9 0 0 13 1 9 9 9 13 1 9 9 0 0 1 9 1 9 9 1 9 9 7 9 7 9 7 9 7 9 15 2
58 7 13 7 9 0 1 9 9 9 0 1 8 8 8 0 1 9 13 9 0 1 9 8 1 9 15 13 15 7 9 1 9 9 1 9 9 0 1 9 9 9 0 1 8 8 7 9 9 15 1 9 0 1 12 9 1 9 2
8 9 0 1 9 9 1 9 9
47 13 9 9 9 0 0 1 9 9 9 9 1 9 15 0 1 9 8 8 9 9 9 9 0 1 9 2 9 1 9 9 0 0 1 9 1 9 1 9 7 9 9 1 9 1 9 2
96 7 13 2 9 9 2 7 9 9 9 0 15 13 9 9 13 9 9 1 9 1 9 2 7 13 9 9 9 1 9 9 10 9 7 1 15 9 1 9 9 0 7 13 15 9 0 2 7 9 1 9 9 9 9 1 9 15 1 9 7 13 15 9 9 1 9 1 9 1 9 1 9 9 8 1 9 12 12 9 7 13 1 9 0 9 15 1 9 7 13 9 15 1 9 0 2
86 1 9 0 13 9 8 0 15 13 1 15 9 1 9 9 0 1 9 7 13 9 9 9 9 7 9 9 1 9 9 0 7 13 9 9 1 9 0 1 9 13 1 15 9 1 9 12 5 7 9 0 0 0 1 9 13 1 12 7 12 5 7 9 0 1 9 13 1 12 7 12 5 7 9 0 0 7 9 9 1 9 1 9 12 5 2
10 9 0 1 9 12 9 1 9 9 0
79 13 9 7 8 2 8 8 14 13 9 9 9 1 9 9 0 0 1 9 9 8 1 9 9 1 9 9 0 7 9 15 1 9 0 0 0 0 1 9 9 7 7 8 2 8 14 13 9 0 1 9 0 1 9 8 7 15 13 9 15 1 9 9 15 14 13 1 9 0 1 12 9 0 7 12 1 9 9 2
100 13 9 9 9 0 1 9 9 1 9 8 2 8 8 8 9 9 9 9 7 9 9 8 8 9 9 9 9 9 0 7 9 0 1 9 9 9 7 9 9 7 9 0 7 9 9 7 9 7 13 9 0 1 9 8 2 8 8 7 15 0 9 7 13 9 9 0 0 1 9 9 9 1 9 1 12 9 7 13 15 9 9 0 0 1 9 1 9 1 9 9 15 14 13 9 15 1 9 0 2
118 13 8 2 8 8 1 7 9 9 14 13 13 9 9 7 9 9 1 9 1 1 7 7 9 0 9 15 14 13 8 9 7 15 15 13 15 9 0 15 13 8 0 9 1 9 9 1 9 9 0 7 9 15 1 9 0 1 9 15 7 9 15 1 9 1 9 12 9 0 14 13 9 15 1 0 1 9 0 0 8 8 8 1 9 7 9 8 8 0 1 9 9 7 1 15 0 15 8 9 1 9 9 15 0 0 1 9 9 15 13 15 0 1 9 7 9 15 2
53 14 1 9 0 7 15 13 1 9 0 1 9 1 9 8 8 7 15 10 13 9 15 1 9 9 9 7 9 1 0 0 7 9 15 1 9 1 9 7 9 9 7 9 9 0 0 1 9 9 0 1 9 2
69 13 8 2 8 8 7 15 13 1 9 9 9 7 9 9 9 9 9 0 1 9 0 1 9 0 8 8 9 7 15 13 1 15 0 0 1 12 12 9 0 1 9 9 9 7 15 13 1 12 5 3 1 9 0 15 13 1 9 7 13 7 13 8 0 1 8 9 0 2
49 13 8 2 8 8 9 15 1 9 15 1 9 0 0 1 9 1 9 9 15 13 1 9 7 15 13 0 9 1 9 0 7 0 1 15 9 9 1 9 9 1 1 9 9 1 9 15 0 2
5 9 13 9 9 0
48 13 9 9 7 9 1 9 9 0 2 7 15 8 9 1 9 9 9 9 13 15 9 1 9 1 9 9 1 9 0 2 1 9 13 1 15 9 9 1 9 9 1 8 0 8 13 9 2
38 7 14 13 9 13 15 9 8 8 1 9 9 0 0 1 9 0 15 13 9 9 9 7 9 1 9 1 9 13 1 0 1 9 7 9 1 9 2
46 7 9 1 9 13 7 9 2 13 1 9 9 0 7 9 9 15 13 0 1 9 7 9 2 7 13 9 0 1 7 15 13 0 9 7 7 15 9 9 0 1 9 9 15 2 2
18 7 1 0 10 13 1 9 0 9 9 0 9 8 8 8 8 8 2
18 9 13 9 0 8 8 8 8 1 9 15 1 2 9 1 0 9 2
42 13 9 0 9 8 8 8 8 1 9 9 0 2 1 0 1 12 9 1 9 9 0 1 9 15 7 9 15 1 9 15 7 13 15 13 1 9 7 13 1 8 2
39 7 13 2 9 9 0 2 7 15 8 9 1 9 2 9 13 1 9 9 9 8 8 2 9 7 9 2 1 9 7 9 15 13 1 9 15 1 9 2
44 7 13 9 2 9 1 15 13 15 9 2 8 2 1 9 15 0 9 2 1 9 13 15 9 13 15 9 8 8 8 13 1 15 9 1 9 13 15 9 9 9 8 8 2
40 7 1 15 13 1 9 7 8 8 2 13 1 0 1 9 9 0 2 8 8 9 7 9 9 0 2 9 15 13 9 15 1 9 15 1 0 9 0 2 2
35 7 13 9 9 9 8 8 8 7 9 2 14 13 9 9 7 9 2 7 7 13 9 9 1 0 9 0 13 9 9 7 9 15 2 2
38 7 13 8 1 2 9 2 2 2 9 14 13 1 9 9 15 13 1 9 9 15 1 9 13 15 9 15 13 1 7 9 0 9 9 15 0 2 2
33 7 13 9 1 2 9 9 9 15 13 15 9 1 9 9 9 15 1 15 9 0 2 7 15 9 1 9 15 1 9 9 2 2
35 7 13 1 9 9 2 9 9 9 9 1 0 0 15 13 15 1 9 7 9 0 9 13 1 15 9 9 1 9 15 7 9 15 2 2
45 7 13 8 15 13 1 9 9 9 7 9 15 1 9 9 15 1 7 15 13 9 9 2 0 7 1 9 0 7 13 1 9 2 7 13 7 3 0 9 7 9 1 9 2 2
49 7 1 9 9 0 1 9 8 8 7 9 15 1 9 15 13 9 0 1 9 9 8 2 7 13 9 9 1 9 1 9 8 8 7 13 9 1 9 0 15 13 1 8 8 1 9 9 9 2
10 8 8 13 9 1 9 9 7 9 0
24 13 9 8 8 9 9 9 9 1 12 8 1 9 9 9 0 0 7 9 9 1 9 0 2
51 13 8 1 9 15 1 9 0 1 9 2 9 9 7 9 9 0 0 2 15 13 1 15 12 9 7 9 1 12 9 0 7 13 15 9 9 9 1 9 1 9 8 8 1 9 1 9 0 1 9 2
58 13 8 8 7 15 1 12 8 1 9 0 0 7 14 8 0 0 1 9 9 1 9 7 9 7 7 15 13 1 9 14 13 1 9 0 1 9 7 0 9 1 15 7 9 0 0 14 13 12 5 1 9 9 0 1 9 0 2
36 13 7 9 0 15 9 9 0 1 9 0 1 9 9 1 9 0 7 0 1 9 9 9 7 9 9 0 7 0 7 9 9 7 9 9 2
31 7 13 9 8 8 1 7 9 0 13 9 9 0 1 9 7 9 7 9 1 9 8 0 1 9 9 0 1 9 0 2
26 14 9 0 7 13 9 1 9 9 0 1 9 9 0 1 0 15 1 1 9 1 9 9 0 0 2
28 7 13 8 8 1 9 0 1 9 1 9 9 0 0 1 9 1 9 9 0 7 9 9 9 1 9 9 2
11 2 9 0 2 2 12 12 9 0 1 9
50 13 0 1 12 9 1 9 0 1 9 9 9 1 9 9 9 0 7 0 9 0 1 9 9 9 9 0 1 9 1 9 12 0 15 13 9 15 12 12 9 0 2 7 9 9 15 13 1 15 2
49 7 13 9 1 9 9 9 1 9 1 9 0 1 9 1 9 9 9 1 9 9 0 15 13 1 7 9 9 0 1 9 15 12 12 9 2 7 15 9 13 1 9 9 9 0 1 10 9 2
68 7 13 9 2 7 1 15 9 8 8 8 7 9 8 8 2 9 9 9 9 8 8 8 8 8 7 9 8 8 8 8 8 8 8 8 8 2 1 9 9 1 9 8 8 9 9 7 9 8 8 8 9 9 9 7 3 9 0 1 9 9 9 0 7 9 0 0 2
74 7 13 9 2 15 13 1 9 2 9 9 10 9 1 9 9 15 13 2 9 1 0 0 15 13 15 9 8 8 8 9 9 9 0 1 9 9 1 9 9 2 1 12 8 9 2 7 13 9 1 9 9 9 1 9 9 7 9 8 1 9 9 9 0 10 1 9 9 7 9 9 1 9 2
68 7 13 9 1 9 9 1 9 10 9 2 7 1 9 9 10 9 9 15 1 9 9 0 15 14 13 7 9 9 15 7 15 13 1 9 9 2 7 1 9 10 9 9 1 10 9 1 9 9 9 15 1 9 15 13 1 15 0 1 9 9 1 9 15 1 9 0 2
33 7 13 9 9 15 1 9 9 8 1 9 9 9 9 1 9 7 9 9 0 1 9 1 7 0 1 9 9 13 15 9 9 2
57 7 13 9 10 9 2 15 13 15 9 0 13 7 9 0 15 12 5 1 9 9 7 9 10 14 13 1 15 9 12 5 7 9 8 7 9 1 9 12 5 2 1 9 0 7 9 9 9 1 9 9 9 1 9 9 0 2
12 9 0 1 9 9 9 13 9 0 9 1 9
81 7 13 9 9 1 9 2 9 2 7 9 2 7 9 0 2 1 9 2 13 9 9 0 8 8 9 9 1 9 9 1 9 1 9 2 7 13 9 0 9 12 2 12 0 9 0 0 9 0 9 0 7 9 15 13 1 9 12 9 0 1 9 9 0 1 9 9 7 13 1 9 9 9 9 7 9 0 9 1 15 2
28 13 8 1 9 13 9 0 1 9 0 8 8 7 9 14 13 1 9 9 0 1 9 9 2 9 0 2 2
21 7 13 9 15 9 1 9 9 1 9 0 1 9 9 9 1 9 14 9 0 2
56 7 1 7 8 13 2 1 9 9 7 9 15 1 7 13 9 15 1 9 2 2 14 7 15 13 7 9 13 9 0 7 13 9 9 2 7 7 15 13 1 9 1 9 1 1 9 9 7 9 0 0 1 9 0 9 2
49 7 1 9 9 0 0 2 13 9 2 8 8 2 0 0 1 7 9 0 1 9 7 9 9 7 9 13 9 0 1 9 1 12 12 9 0 1 9 13 9 9 15 1 9 13 1 8 8 2
41 7 13 10 9 1 9 2 8 8 2 15 13 15 9 1 1 9 15 15 13 1 15 9 9 0 9 1 15 15 13 15 9 9 7 15 13 15 1 9 9 2
43 7 13 9 0 0 0 9 7 9 1 9 9 7 9 8 1 9 2 7 13 9 1 9 1 10 9 2 10 13 9 1 0 9 0 1 9 7 7 9 1 9 0 2
34 7 13 9 0 1 9 9 0 1 9 9 2 8 2 0 1 9 9 8 8 9 9 2 7 15 13 9 1 9 9 7 9 8 2
14 7 15 13 9 0 1 9 0 1 12 1 12 9 2
21 7 13 9 1 9 10 9 1 9 0 1 9 8 8 8 8 7 9 8 8 2
83 7 13 9 1 9 0 9 15 7 9 14 13 9 15 9 9 12 2 0 7 15 13 9 9 1 2 9 2 9 10 9 15 13 15 9 2 9 0 2 0 1 9 2 9 9 0 0 2 1 2 9 2 9 15 0 7 9 15 1 15 2 7 1 7 9 15 1 2 9 9 1 9 9 9 2 9 1 9 9 9 1 15 2
21 8 14 13 9 2 9 0 0 2 1 9 1 14 2 8 2 1 9 9 1 0
29 13 2 9 2 7 9 0 13 1 9 13 15 2 9 0 0 2 2 7 13 7 13 1 15 9 8 8 0 2
44 7 13 9 9 0 1 9 9 0 8 8 9 9 15 0 1 9 10 2 9 2 2 7 13 15 1 15 1 9 9 13 15 0 1 8 2 1 9 9 9 8 1 8 2
17 7 13 7 9 15 8 8 0 1 9 10 9 7 9 1 15 2
45 7 9 7 13 15 8 15 1 9 2 9 9 2 1 9 1 9 1 9 2 2 1 9 9 7 9 9 9 7 9 2 2 7 13 9 1 2 8 2 9 15 7 9 15 2
33 7 13 9 0 0 9 9 9 0 1 2 9 0 1 9 7 9 2 7 9 8 15 13 1 9 9 9 9 0 0 1 9 2
35 7 13 8 9 7 9 0 1 9 15 0 15 13 1 9 1 9 0 2 7 13 9 15 1 2 9 0 2 14 13 10 9 1 15 2
25 7 13 9 0 1 7 9 8 13 1 9 9 9 8 7 13 9 9 7 9 1 9 1 9 2
35 7 13 9 0 1 2 9 2 7 9 0 13 8 2 14 9 15 9 10 9 1 9 2 2 7 13 0 7 9 0 2 13 9 2 2
73 7 7 13 15 13 9 0 2 0 1 9 10 9 2 13 8 7 10 9 2 9 9 13 15 9 9 1 9 1 9 1 9 0 2 7 7 13 10 9 13 9 1 9 10 9 14 13 13 9 2 2 7 13 15 1 9 1 9 0 13 1 9 0 1 9 0 9 1 9 1 9 0 2
52 7 13 9 7 9 9 0 13 8 1 9 0 2 7 13 7 9 2 14 13 9 7 3 9 1 9 1 9 0 7 0 2 14 13 15 9 0 2 14 7 15 14 13 9 9 1 9 13 7 13 2 2
25 7 1 9 9 9 9 0 2 13 9 0 0 15 13 15 9 15 2 14 9 7 13 9 8 2
43 7 1 9 15 1 2 9 2 13 8 7 2 9 9 0 9 15 1 9 9 0 1 0 1 9 0 2 7 1 9 9 8 8 1 9 9 7 13 9 10 9 2 2
21 7 9 9 13 1 9 2 9 9 0 2 9 0 1 9 8 1 10 9 2 2
12 12 12 9 1 8 1 9 9 9 0 1 9
43 13 9 9 9 0 0 8 2 9 2 1 9 15 0 1 9 9 1 9 9 0 9 15 12 8 9 1 9 9 0 1 9 0 15 13 8 7 9 7 9 1 9 2
57 13 1 15 1 2 9 9 2 8 8 8 9 0 1 9 2 7 13 7 10 9 13 1 15 9 0 2 7 13 8 9 1 8 8 7 13 7 9 1 9 9 1 9 9 0 1 10 9 1 9 9 9 9 0 1 9 2
54 7 13 1 7 3 9 0 14 13 9 1 9 15 1 15 9 9 0 1 9 1 8 7 9 7 1 9 9 9 0 7 14 13 1 9 9 1 9 0 7 0 1 9 9 9 0 1 9 7 15 9 9 9 2
45 7 0 1 9 7 9 9 9 0 0 13 1 9 9 0 2 12 12 9 2 7 9 9 0 1 15 12 12 9 2 7 9 9 0 12 9 7 0 9 9 13 12 12 9 2
22 7 13 7 8 13 1 0 1 12 12 9 7 7 9 9 13 12 12 7 12 9 2
68 7 13 1 7 8 2 8 2 8 14 13 1 9 9 15 1 9 7 14 13 12 9 0 1 15 1 9 9 12 7 13 9 9 1 9 1 12 9 1 9 10 9 2 7 7 9 0 0 0 1 9 9 9 7 14 13 0 7 0 1 9 12 0 1 9 1 9 2
58 7 9 1 9 1 9 9 1 9 9 0 0 1 9 1 9 13 8 8 7 9 13 9 0 1 9 15 1 9 9 9 0 1 9 0 14 13 9 15 1 8 8 9 1 9 15 7 13 7 10 9 13 9 15 12 12 9 2
58 13 7 9 13 9 9 0 7 1 15 9 0 9 7 9 9 13 13 1 9 0 1 9 0 7 1 0 13 1 15 9 1 9 9 9 1 9 1 9 9 0 0 1 9 1 9 9 1 9 9 0 7 0 7 3 9 0 2
44 7 13 7 15 14 13 1 9 0 9 0 1 9 1 9 1 9 9 15 1 9 1 9 7 7 15 14 13 9 1 10 9 14 1 9 9 0 1 0 7 8 1 0 2
31 7 13 8 8 8 7 15 13 9 1 9 1 9 0 1 9 9 7 13 9 15 1 9 0 1 15 1 9 0 0 2
12 13 7 10 9 0 1 9 0 0 7 0 2
13 0 1 12 12 9 9 9 0 0 1 9 9 0
58 13 12 1 9 9 0 1 9 9 9 7 9 1 9 9 0 1 9 9 9 0 0 1 7 13 9 0 1 9 7 9 1 9 9 7 9 0 7 9 7 9 8 7 9 0 13 9 15 12 12 9 2 12 12 9 0 2 2
43 7 13 9 1 7 10 9 0 13 12 5 1 9 9 2 7 13 9 0 9 9 1 9 9 9 9 0 1 9 10 13 1 9 2 7 9 9 9 7 9 9 15 2
23 7 13 9 8 8 9 9 14 13 9 9 12 1 9 9 9 0 0 1 9 12 9 2
13 12 9 9 9 0 9 9 9 0 7 0 1 9
89 13 0 7 9 9 0 9 9 9 9 0 1 9 0 7 0 1 9 0 9 7 9 7 9 1 1 12 9 2 7 13 1 9 0 0 9 9 9 9 1 9 9 0 8 7 9 0 9 8 1 9 0 1 9 9 1 9 15 0 1 9 9 15 7 9 0 15 1 9 9 15 1 12 12 9 7 3 9 9 9 15 0 1 9 9 9 1 15 2
48 7 13 9 7 9 9 0 13 1 15 9 0 1 9 0 1 9 9 9 0 7 8 7 9 2 7 9 15 9 13 9 1 9 9 15 1 9 9 15 13 1 9 9 0 1 9 0 2
65 7 13 7 9 0 0 0 12 12 9 7 3 9 9 0 0 1 9 7 1 0 7 14 9 9 1 9 0 7 0 14 13 1 9 10 9 2 7 14 13 9 1 9 9 0 1 9 9 15 1 9 9 9 7 9 7 8 15 13 9 9 15 1 9 2
93 7 13 9 9 0 1 9 1 9 9 0 0 8 8 7 9 9 9 8 1 9 9 1 15 13 9 1 9 0 1 9 9 0 15 14 13 13 9 0 1 9 9 0 7 13 1 12 5 1 15 1 9 0 1 9 0 0 12 2 12 1 9 12 8 9 1 12 8 9 1 8 7 12 8 9 1 9 0 7 12 8 9 1 9 0 7 1 12 12 9 1 8 2
45 7 13 7 12 5 1 9 9 0 1 9 0 7 0 1 12 12 9 13 1 9 13 9 9 15 1 9 1 9 14 13 1 12 5 9 15 13 9 0 9 0 13 12 9 2
61 7 13 8 8 1 9 9 9 9 9 1 9 1 9 0 2 7 13 9 9 9 9 0 8 8 9 1 9 0 1 9 7 9 0 7 9 9 7 9 0 0 15 13 9 15 1 9 7 13 1 9 0 0 1 9 0 1 15 9 0 2
8 9 0 1 9 1 12 9 0
260 13 9 9 0 1 12 9 0 15 9 7 9 7 9 7 9 8 8 7 9 7 9 7 8 7 9 9 0 7 9 7 13 9 1 12 9 0 15 9 7 9 7 9 7 9 7 9 7 8 7 8 7 13 9 0 1 9 0 1 9 0 1 9 1 9 1 9 12 8 8 9 1 9 8 1 9 12 7 13 9 0 1 8 1 9 12 5 7 13 0 9 1 15 15 9 7 9 8 7 13 9 0 1 9 1 9 12 5 7 13 0 9 1 8 7 9 7 1 9 1 9 12 5 13 1 9 7 9 0 7 9 0 7 1 9 12 5 7 13 1 9 0 7 9 9 8 8 8 7 1 9 12 5 7 13 1 9 8 8 0 7 9 7 9 7 1 8 12 5 7 13 1 9 7 9 7 9 0 7 9 7 9 0 7 14 13 9 0 1 9 0 1 9 9 7 13 8 8 1 8 7 13 9 7 9 7 9 9 7 13 8 8 1 9 7 13 9 1 9 9 8 1 1 13 8 8 1 9 1 9 12 5 7 13 1 9 9 9 7 13 8 8 1 9 1 9 12 5 7 13 1 9 0 7 9 8 8 8 9 2
15 9 13 1 12 9 1 9 2 9 2 1 0 9 0 0
17 13 9 0 1 9 1 9 9 9 0 1 0 9 0 1 8 2
38 13 8 9 0 0 9 1 1 9 0 1 12 9 0 1 12 9 15 8 7 8 7 8 7 9 7 9 7 9 7 15 1 9 1 9 0 0 2
20 13 1 15 1 2 8 2 8 8 9 9 9 9 7 9 1 9 9 0 2
11 7 13 7 9 9 13 12 12 9 0 2
48 7 13 9 0 1 9 9 1 0 1 9 9 0 9 1 9 1 10 9 1 9 12 1 9 1 9 9 1 9 9 7 9 7 13 1 9 9 0 9 1 9 9 0 7 9 9 15 2
47 7 13 8 8 7 9 1 9 0 7 0 13 1 9 12 9 0 1 9 1 9 0 1 9 7 9 9 0 7 0 1 9 0 1 0 9 0 7 13 1 9 0 1 9 9 0 2
18 7 13 7 10 9 13 9 9 1 9 1 9 0 7 9 15 2 2
16 7 13 0 1 9 0 1 9 9 9 0 1 9 9 15 2
29 7 13 8 8 7 9 9 13 1 9 1 9 0 7 1 1 9 7 13 9 1 9 0 0 1 9 13 9 2
22 7 13 7 9 0 14 13 0 9 0 1 9 9 9 9 0 0 1 9 1 9 15
6 9 8 8 1 8 0
70 1 9 9 9 0 1 9 9 9 1 9 9 2 9 1 9 0 8 9 9 1 8 0 1 9 12 5 7 13 1 12 12 9 2 1 9 9 9 9 0 2 7 9 2 7 9 9 9 0 1 9 12 5 7 13 1 12 12 9 1 12 12 9 1 9 9 1 9 12 2
39 7 13 9 1 9 9 7 9 7 9 0 1 9 12 5 7 13 1 12 12 9 2 9 9 9 1 8 7 9 0 2 7 9 9 0 7 9 0 2
27 7 13 3 9 9 0 1 9 12 5 7 13 1 12 12 9 2 1 12 12 9 1 9 9 2 9 2
111 1 1 13 9 9 9 7 9 1 9 12 5 7 13 1 12 12 9 1 9 9 2 9 12 1 12 12 9 1 9 9 1 9 7 1 9 1 9 9 1 9 9 7 1 15 9 0 13 0 1 7 9 9 9 13 12 5 1 9 9 0 1 9 1 9 0 7 9 0 7 0 7 9 0 2 9 9 2 2 1 1 13 10 9 1 12 5 8 8 0 2 7 12 5 1 9 0 2 7 12 5 1 9 0 2 7 12 5 1 9 2
65 1 9 0 2 13 9 9 1 9 9 9 12 5 2 7 9 0 12 5 7 13 9 9 1 9 2 8 8 2 1 12 12 7 12 12 9 2 7 1 9 1 12 9 2 7 9 10 9 14 13 1 9 9 0 7 7 15 13 1 9 3 1 9 0 2
15 12 5 9 1 8 8 0 7 12 5 9 1 9 9 0
17 1 9 9 9 1 1 9 9 1 9 9 2 9 1 9 0 2
79 13 9 3 9 9 1 9 12 5 7 13 1 12 12 7 12 12 9 9 9 9 9 9 0 1 9 12 5 7 13 1 12 8 7 12 12 9 2 1 9 9 0 7 13 1 12 8 2 7 9 9 0 1 12 12 9 2 7 9 0 1 12 12 9 2 1 1 13 9 9 8 8 1 12 7 12 12 9 2
17 7 13 9 0 1 9 12 5 7 13 1 12 7 12 12 9 2
17 7 1 9 1 9 9 0 1 9 9 2 9 1 9 0 2 2
123 7 14 13 9 9 15 1 12 8 7 12 12 9 2 1 15 12 12 9 1 9 8 2 8 8 1 9 0 1 9 12 5 1 9 12 2 7 13 12 8 7 12 12 9 2 7 13 9 9 0 1 9 9 2 1 1 9 2 1 9 12 5 7 13 1 12 7 12 12 9 2 7 13 1 9 9 0 1 10 9 1 0 9 9 1 1 12 5 1 12 12 9 1 12 12 9 2 1 1 13 9 10 9 1 12 8 7 12 12 9 1 15 12 12 9 1 9 0 8 8 1 9 2
71 14 9 9 0 0 2 7 14 13 9 15 1 12 12 9 1 9 9 2 9 1 9 0 2 1 15 1 12 12 9 9 1 9 9 0 8 8 1 9 8 2 1 1 13 9 9 1 10 9 1 12 7 12 12 9 2 1 15 12 12 9 1 9 9 0 8 8 1 9 8 2
10 9 9 0 1 9 8 1 1 9 0
28 13 9 1 9 9 0 9 0 1 9 9 0 0 1 9 1 9 9 0 1 9 9 8 1 1 9 0 2
58 7 13 9 15 13 1 9 15 13 9 12 2 12 0 1 9 0 0 0 1 9 0 1 9 7 13 9 9 0 0 1 9 1 9 0 0 7 9 0 1 9 1 9 1 9 0 1 9 0 7 9 0 0 7 9 0 9 2
53 7 13 8 8 9 9 9 0 0 1 7 9 10 9 15 9 9 0 1 9 9 0 15 13 9 15 1 9 9 8 2 1 7 13 9 9 9 0 1 9 0 1 1 9 9 15 13 15 9 0 1 9 2
37 7 1 0 7 13 9 0 1 9 1 10 9 1 1 9 9 0 1 9 9 15 1 9 1 9 0 7 9 9 0 1 9 9 1 9 0 2
11 9 1 8 0 7 9 9 13 12 12 9
74 13 9 1 9 9 8 8 9 9 15 13 15 0 1 0 7 0 1 9 9 15 13 15 9 8 0 1 9 0 1 9 9 1 9 9 15 1 9 2 8 8 2 7 13 9 15 12 5 1 9 8 8 9 0 1 0 9 9 0 15 13 9 15 0 1 12 12 9 2 12 8 9 2 2
55 7 13 9 0 0 9 1 9 9 13 9 9 9 15 7 9 9 9 14 13 1 9 2 8 2 9 2 7 13 7 9 0 13 9 9 7 13 9 0 1 9 9 15 1 9 9 15 14 13 9 9 9 1 15 2
40 14 7 9 13 9 1 9 9 1 9 7 9 15 7 9 0 15 13 9 1 15 1 9 7 13 1 9 7 3 9 13 1 9 0 1 9 7 9 9 2
13 7 13 2 8 7 13 9 10 9 1 9 2 2
35 7 1 9 9 2 8 8 2 13 8 8 9 9 0 1 9 0 7 2 8 8 2 13 9 9 9 1 9 9 7 9 0 1 15 2
49 7 13 9 9 0 2 8 8 2 1 9 1 9 0 1 9 0 7 15 13 9 1 9 7 9 15 2 0 1 7 9 13 1 8 1 2 9 2 9 0 14 7 15 14 13 9 1 15 2
46 7 13 9 14 13 1 9 0 1 9 8 0 1 9 2 8 2 1 9 8 8 0 1 9 9 9 9 12 5 1 8 8 8 8 8 3 14 7 9 14 13 10 9 1 9 2
13 9 0 9 1 9 2 9 0 2 8 1 10 9
64 13 9 1 9 9 0 7 15 14 13 9 1 9 9 9 8 8 1 9 1 7 13 9 1 9 8 9 1 9 9 9 13 1 2 9 9 2 7 13 9 1 2 9 0 7 9 13 7 13 9 9 9 1 9 9 7 7 15 14 13 0 9 0 2
46 7 13 9 9 15 13 15 9 0 8 8 7 9 8 2 13 7 13 9 1 7 9 13 1 9 9 7 13 1 9 0 1 9 15 1 9 7 14 13 9 9 1 9 0 2 2
40 7 14 13 12 1 9 9 9 0 1 8 1 9 15 1 9 9 7 1 15 2 1 8 15 15 0 1 9 15 1 9 0 7 9 0 0 1 9 0 2
19 7 1 9 9 8 13 9 0 8 8 9 15 9 9 0 1 9 9 2
37 7 13 8 8 8 1 8 7 13 15 0 0 1 9 9 0 1 9 9 0 7 0 13 13 1 15 9 9 15 1 9 0 1 9 9 0 2
13 9 2 9 0 13 1 9 9 0 9 1 9 0
75 13 9 0 1 9 0 1 7 9 2 9 9 2 7 9 0 15 0 0 1 9 9 0 1 9 9 7 9 1 9 9 13 7 9 9 0 1 9 9 15 9 1 9 0 1 9 10 9 1 9 0 2 1 1 7 9 0 1 9 9 13 7 13 9 0 1 9 0 1 9 1 9 9 0 2
33 7 13 9 1 2 9 9 7 0 0 2 1 9 1 2 9 2 7 9 13 9 9 0 1 9 8 8 8 8 8 1 9 2
35 0 1 15 2 7 9 9 1 2 9 8 2 7 9 0 7 0 1 9 1 9 0 7 9 9 0 0 13 1 9 1 9 1 9 2
47 7 13 7 9 0 1 9 2 13 7 9 9 0 0 0 15 9 0 1 9 1 9 15 7 1 9 9 9 9 15 0 2 1 9 7 13 9 9 0 1 9 0 9 1 9 2 2
28 7 13 1 7 0 15 13 9 9 15 9 9 1 9 0 0 1 15 9 1 9 1 9 0 1 9 0 2
21 1 9 0 2 7 14 9 1 9 9 1 9 13 13 9 9 1 9 9 9 2
43 7 1 9 13 9 9 9 9 0 0 1 9 9 1 9 9 9 0 2 7 13 9 0 9 1 10 9 2 0 1 9 15 0 1 9 0 7 9 9 0 1 9 2
40 1 9 0 2 7 7 9 9 9 0 1 9 9 14 13 1 9 9 9 0 1 9 10 9 1 9 9 0 2 7 14 13 9 1 9 9 0 1 9 2
63 7 1 9 9 0 1 9 0 2 13 9 1 9 9 1 7 9 9 15 13 1 7 13 9 10 9 0 7 13 1 9 9 9 1 9 0 14 13 15 9 9 0 1 9 15 2 13 9 2 2 1 1 13 9 1 9 15 1 9 1 9 0 2
15 9 0 2 9 8 8 13 1 9 1 9 0 1 9 8
62 13 9 0 0 1 9 9 9 8 1 2 9 0 2 1 9 0 1 9 9 9 0 8 8 1 9 1 9 9 15 0 1 12 9 0 9 1 9 9 0 0 13 9 2 9 1 9 2 1 9 1 9 0 1 9 0 7 0 1 9 8 2
97 7 13 9 9 15 15 13 1 9 9 1 9 15 2 7 9 9 8 8 13 1 9 0 1 9 9 0 8 8 8 8 15 13 9 12 2 12 0 2 7 3 1 12 9 1 9 9 9 9 0 2 12 0 12 2 1 8 2 13 7 9 9 8 1 8 9 12 2 12 0 14 13 1 9 9 7 7 9 0 14 13 1 9 9 1 9 8 8 9 1 9 9 8 7 9 8 2
8 8 9 0 0 1 9 7 9
10 13 9 9 0 1 8 1 12 9 2
6 12 2 9 9 0 2
35 7 15 9 0 2 0 2 13 1 9 7 13 9 0 1 9 15 1 9 0 1 8 7 13 1 9 9 7 9 9 0 0 1 9 2
35 7 13 9 10 9 2 1 9 9 0 1 8 2 9 0 1 9 0 2 9 9 8 0 2 9 9 0 1 8 2 9 9 9 0 2
6 7 0 10 9 12 2
51 9 8 0 15 13 1 9 2 1 9 9 0 9 15 1 9 9 9 9 0 2 7 1 9 8 8 8 2 8 8 9 0 1 9 2 13 9 1 9 8 7 13 1 15 9 9 0 14 13 1 2
48 7 13 3 2 9 9 7 9 0 2 1 9 9 8 8 8 2 15 13 9 12 2 7 13 15 1 9 15 9 15 8 7 9 9 15 1 8 2 7 13 1 9 9 9 0 1 8 2
20 7 3 9 9 0 2 15 13 1 9 0 7 15 14 13 9 1 9 15 2
8 7 3 2 9 9 0 2 2
57 14 7 9 0 9 1 9 0 15 13 9 1 9 0 1 8 9 12 2 12 0 2 15 2 9 9 9 0 0 2 2 7 13 9 15 9 12 2 7 13 3 1 2 8 2 8 2 2 7 13 1 9 0 0 1 8 2
6 12 2 9 9 0 2
31 7 15 15 13 15 9 0 1 8 7 13 1 0 15 7 9 15 1 9 1 9 0 1 9 0 1 9 7 1 9 2
25 7 13 10 9 2 9 1 9 15 0 7 0 7 1 9 15 0 0 8 8 8 8 0 2 2
12 8 7 15 1 9 8 2 9 1 9 0 2
22 7 9 0 2 0 2 15 13 1 9 0 1 9 9 1 9 8 8 7 9 15 2
81 7 0 10 9 2 8 2 9 1 8 8 8 8 2 2 7 15 9 9 0 15 9 8 8 8 9 9 1 9 7 9 7 9 7 9 9 1 8 7 1 15 7 15 13 9 0 1 9 0 2 7 9 2 8 8 2 7 0 15 8 8 2 7 1 10 9 8 7 15 0 9 1 9 15 7 9 8 7 9 8 2
6 12 2 9 9 0 2
35 13 1 9 12 1 9 9 9 0 15 14 13 7 13 9 12 2 7 13 15 9 9 0 9 12 7 15 13 1 13 1 9 12 0 2
14 7 1 9 12 13 9 9 15 13 1 9 9 12 2
32 7 9 10 9 13 15 2 9 9 0 2 1 8 9 9 8 15 13 9 9 9 9 9 9 1 9 7 9 9 9 12 2
47 9 7 9 9 8 1 9 12 2 13 9 0 1 9 0 1 0 2 7 13 9 9 1 9 9 12 7 13 1 9 9 15 1 9 7 1 9 9 9 7 1 1 15 8 9 15 2
38 7 1 9 1 9 9 15 13 9 9 1 9 1 9 9 0 2 1 9 8 8 7 13 9 9 1 9 9 12 1 12 5 9 12 1 12 5 2
38 7 13 8 9 9 0 1 9 13 1 9 9 2 8 1 9 8 8 8 2 1 9 1 8 8 8 2 7 0 1 9 8 2 1 9 8 2 2
51 7 13 9 9 9 1 9 12 9 1 9 9 0 1 9 0 1 8 1 9 2 9 9 15 13 1 9 1 9 9 15 1 9 8 7 9 9 7 9 1 9 8 7 13 1 9 1 9 9 15 2
50 7 1 9 0 15 13 1 12 9 12 2 13 9 7 9 9 0 7 13 12 5 1 9 15 13 15 9 1 9 7 9 9 0 1 0 15 14 9 9 7 14 13 1 12 5 7 13 1 9 2
31 7 1 9 9 1 8 1 9 9 0 2 13 9 9 1 9 0 9 0 13 1 15 8 9 1 9 9 1 8 8 2
15 9 1 9 1 8 7 8 1 2 9 2 0 2 0 2
52 13 9 2 8 2 0 9 12 2 12 0 7 9 0 1 9 9 9 0 9 8 1 9 8 8 1 8 2 8 9 9 1 8 7 9 9 0 8 8 2 2 7 7 2 9 1 9 10 9 13 2 2
36 7 13 9 1 9 0 0 0 9 9 15 7 9 2 13 9 1 9 15 1 9 0 7 13 9 1 9 0 7 9 9 15 1 15 2 2
22 7 13 9 1 9 7 13 9 9 0 8 8 1 9 1 9 2 1 9 0 2 2
23 7 13 7 15 13 2 9 0 1 9 9 1 9 7 9 9 1 9 1 9 0 2 2
21 7 13 9 8 2 8 1 8 1 7 15 2 9 9 0 2 1 9 7 9 2
18 7 13 9 1 9 9 0 9 12 2 12 0 9 1 8 9 0 2
7 9 0 13 1 2 8 2
2 8 2
4 8 2 9 9
17 13 9 0 7 9 9 0 8 8 13 9 9 9 0 1 9 2
25 7 14 13 9 9 0 2 8 8 8 2 9 7 9 7 9 9 0 1 9 1 9 1 9 2
37 7 14 13 9 0 2 1 9 2 9 0 0 8 8 2 7 15 9 1 9 8 0 0 15 13 9 1 9 0 7 0 0 1 9 8 0 2
31 7 13 8 8 8 8 9 9 8 0 9 10 9 1 9 2 8 8 8 2 1 8 1 9 8 1 9 9 9 0 2
32 7 13 9 7 9 0 7 1 9 9 9 9 0 1 9 0 1 15 1 9 1 9 0 7 9 1 10 9 8 1 15 2
10 12 1 9 9 1 9 13 9 1 9
30 13 1 12 9 1 15 9 9 7 9 9 9 9 0 1 9 1 9 9 9 2 7 15 1 9 0 1 9 8 2
48 7 13 9 9 7 15 1 9 15 1 9 9 7 9 7 0 0 2 9 1 12 1 9 8 0 2 1 9 2 9 2 13 15 9 0 15 8 8 1 9 9 7 9 0 1 9 9 2
24 7 13 10 9 9 1 9 9 0 0 0 1 9 7 9 9 13 7 13 9 8 9 12 2
14 9 0 0 13 2 9 8 14 13 9 1 2 8 2
63 13 9 13 15 9 1 9 9 9 0 0 7 9 9 8 8 14 13 9 1 9 2 9 9 0 2 2 8 2 1 9 9 0 7 14 13 1 9 1 9 9 0 9 1 9 2 7 7 13 9 8 7 7 9 14 13 2 0 7 9 0 2 2
38 7 13 9 15 13 9 2 8 2 0 9 1 15 1 9 15 1 2 9 8 2 2 1 7 3 2 9 0 7 13 8 1 9 1 9 8 2 2
67 7 13 9 9 0 1 9 0 1 9 9 0 2 8 2 7 0 2 8 2 7 9 9 0 2 8 2 1 9 9 9 9 1 10 9 0 9 9 8 8 2 1 9 1 9 1 9 0 1 9 9 0 7 2 9 0 2 13 9 7 15 13 9 9 9 15 2
31 7 13 8 9 9 0 1 9 0 0 0 7 15 13 1 2 9 9 9 0 1 9 10 1 8 1 9 9 9 2 2
17 7 13 9 1 7 9 9 0 1 9 15 7 2 13 9 15 2
28 7 7 13 9 0 7 13 1 9 1 9 9 7 9 7 14 15 14 13 9 7 9 9 2 15 13 15 2
35 7 13 9 2 2 7 14 13 9 2 1 9 9 2 9 0 7 14 8 14 13 9 0 0 15 14 13 1 15 9 1 9 0 2 2
44 7 13 9 7 15 0 1 7 9 0 14 13 1 9 9 0 2 7 9 9 13 1 2 9 9 0 7 0 1 9 0 1 9 7 13 9 1 9 9 1 9 9 2 2
51 7 13 9 7 9 7 9 9 15 13 15 9 9 1 9 0 2 13 9 0 15 13 1 15 9 9 1 9 8 7 13 9 9 0 1 9 2 8 13 1 9 1 10 9 9 9 1 9 0 2 2
18 8 9 13 1 9 2 9 8 2 7 13 1 2 8 13 9 8 2
54 13 9 9 7 9 0 9 8 8 1 9 2 9 8 2 7 0 1 15 2 9 1 15 13 1 9 9 2 9 2 1 9 0 1 9 9 0 2 0 1 9 9 2 7 15 13 1 15 9 2 9 9 2 2
14 7 13 8 9 1 2 0 7 0 1 9 0 2 2
37 7 13 2 8 2 9 8 1 9 9 9 9 15 13 15 1 9 9 0 7 13 1 15 1 9 1 9 2 15 13 9 8 1 9 9 2 2
33 7 13 8 2 15 13 8 8 13 1 9 0 9 1 9 9 8 1 9 9 2 2 0 7 2 9 9 14 13 1 9 0 2
16 7 9 9 9 1 9 9 7 15 9 0 1 9 0 2 2
50 7 13 1 7 2 9 9 0 13 1 1 12 9 1 9 9 9 1 9 1 9 15 9 0 7 9 1 9 2 7 13 15 7 13 15 1 0 7 13 1 15 9 7 9 9 9 9 2 2 2
14 7 13 2 2 10 9 0 7 0 1 9 0 2 2
20 7 13 7 2 9 8 9 0 7 14 8 1 15 14 0 7 14 0 2 2
24 7 13 7 2 9 13 0 9 15 13 9 9 1 9 0 7 13 1 9 7 9 15 2 2
13 7 14 13 9 9 7 9 0 1 9 15 2 2
10 7 13 9 9 7 9 7 9 2 2
25 7 13 9 8 13 1 9 9 15 13 9 9 1 2 9 8 2 7 13 15 13 1 15 2 2
10 14 13 9 9 0 1 9 7 9 2
51 13 9 2 9 2 0 9 1 10 9 13 1 15 2 1 9 0 13 9 9 8 1 9 7 9 7 13 9 0 9 1 9 9 8 8 1 9 1 9 0 7 13 1 15 9 0 9 9 9 9 2
30 7 13 9 9 9 1 9 0 2 7 14 13 9 0 1 9 9 0 0 1 9 9 9 1 9 7 0 7 9 2
24 2 2 9 0 7 0 9 0 1 9 15 9 9 1 9 9 1 9 0 1 9 9 0 2
94 13 10 9 1 9 0 0 0 1 9 9 0 2 7 13 9 9 9 0 2 7 15 15 13 9 0 13 9 0 0 2 7 13 1 15 9 7 0 2 7 13 9 0 1 9 9 15 2 7 14 13 10 9 7 14 13 0 1 9 9 2 7 15 14 13 9 9 7 13 0 9 0 2 7 14 1 0 7 13 9 9 1 9 1 9 9 9 1 0 1 0 9 0 2
74 9 8 8 9 9 0 0 1 9 9 0 13 7 9 7 9 0 1 9 7 0 14 13 1 13 9 9 9 9 0 1 9 9 1 9 9 0 2 7 13 9 0 1 9 0 1 9 0 1 9 0 1 9 9 9 0 1 9 9 9 7 9 0 9 0 1 9 0 0 7 1 9 0 2
24 7 13 9 0 1 0 1 9 0 1 9 0 15 13 9 15 1 9 0 7 9 9 0 2
56 7 1 9 0 7 14 9 0 13 1 9 9 9 1 9 9 9 0 1 9 2 7 1 0 7 13 9 0 1 9 9 1 9 0 9 9 1 7 13 15 9 1 9 9 0 0 1 9 9 7 9 1 9 9 0 2
133 2 2 0 9 0 7 13 9 8 8 1 9 0 0 1 9 0 0 1 9 9 1 9 0 7 0 0 13 0 1 1 9 0 7 9 0 0 7 13 9 0 1 9 15 13 1 15 8 1 9 9 2 7 13 1 9 0 0 1 9 9 9 1 9 0 2 7 3 13 9 1 9 9 0 7 1 15 9 0 0 7 9 0 0 0 1 9 9 15 13 15 9 1 9 2 8 2 9 9 9 0 1 9 7 9 2 7 13 9 9 0 0 7 14 13 10 9 0 9 7 9 7 9 7 0 3 7 13 1 9 9 0 2
73 7 14 13 9 10 9 0 1 9 0 1 9 2 7 1 0 1 13 9 1 9 9 9 2 7 9 9 9 2 7 13 9 7 9 8 0 14 13 9 15 1 9 9 7 9 15 2 7 1 9 9 15 13 9 15 1 9 1 9 9 1 9 15 2 7 9 15 13 1 9 9 0 2
23 7 13 7 9 0 14 13 0 7 13 9 1 9 15 1 9 1 9 7 0 7 9 2
50 7 13 9 8 8 7 9 0 0 14 13 9 9 0 15 13 9 9 9 9 1 9 2 7 1 0 1 9 9 1 9 9 0 2 7 9 9 9 0 1 9 9 0 1 9 7 9 7 9 2
29 2 2 9 9 7 7 14 13 7 13 9 1 9 9 1 9 1 9 9 0 1 15 7 9 9 0 1 9 2
64 13 9 8 8 8 9 1 9 9 0 7 0 1 9 7 9 9 9 9 0 0 7 15 1 0 7 13 9 9 1 9 1 9 10 7 13 9 1 0 1 0 9 0 2 7 9 10 13 9 0 9 7 15 13 7 13 9 1 7 14 13 1 0 2
43 7 9 9 7 13 0 14 13 0 2 8 8 8 1 9 7 13 9 7 13 9 15 2 7 9 9 0 7 14 13 9 0 7 1 15 8 1 9 9 0 1 9 2
18 14 1 9 9 9 15 13 15 9 1 9 1 10 9 7 13 8 2
106 8 8 8 7 3 9 13 15 9 1 9 7 1 9 10 13 1 9 8 8 2 8 7 9 13 10 9 2 7 8 7 8 7 8 7 0 8 14 13 9 1 10 9 2 9 9 1 9 0 7 15 13 1 9 13 15 7 15 13 7 9 15 1 9 0 2 7 15 14 13 7 13 1 9 2 7 9 9 9 0 1 9 0 2 7 7 15 13 1 9 0 1 9 0 7 0 9 7 0 1 15 9 1 9 8 2
151 2 2 9 9 0 7 1 9 0 7 9 9 1 9 1 0 9 1 9 10 7 13 9 1 0 9 0 2 13 9 8 8 7 9 0 13 0 7 15 0 1 9 1 9 15 2 7 1 9 9 7 13 1 15 9 0 2 7 7 14 13 9 9 0 0 2 7 14 13 3 9 1 9 7 1 0 14 13 3 9 2 8 1 14 9 7 13 9 9 2 14 13 9 1 9 9 9 1 10 9 2 7 14 13 9 15 0 2 7 13 8 7 13 3 9 0 1 8 9 0 0 7 9 9 9 0 2 7 7 9 14 13 9 8 8 0 1 9 2 7 8 8 8 7 13 9 0 1 0 9 2
154 7 13 9 0 0 1 9 9 0 8 8 8 8 7 9 0 1 9 14 13 1 9 2 7 0 7 9 0 13 13 9 0 9 0 8 1 9 9 9 0 1 9 0 2 15 13 1 9 9 8 8 8 8 3 2 7 7 7 13 1 9 9 7 9 9 9 0 1 9 7 9 9 0 1 9 9 13 9 9 0 1 15 2 7 1 9 0 1 9 12 2 12 2 12 2 12 2 7 1 9 9 0 2 1 9 1 9 12 2 7 9 1 9 0 9 12 7 1 9 0 1 9 15 0 1 9 0 0 1 15 2 7 9 0 0 1 9 9 9 0 7 15 13 15 1 9 13 7 13 1 9 9 2 2
61 2 2 9 0 7 9 0 7 13 8 8 8 7 15 1 9 9 0 7 14 9 0 0 0 9 1 9 0 0 2 7 1 0 0 7 9 1 0 13 13 9 0 9 1 9 0 0 1 9 0 8 8 13 9 0 1 9 0 1 9 2
45 7 1 3 13 9 0 9 15 1 9 0 0 2 7 15 14 13 9 9 0 1 0 2 9 1 9 9 9 7 15 13 15 1 9 1 0 1 9 9 9 0 7 9 0 2
36 7 1 9 9 7 15 0 1 9 8 8 7 9 15 2 7 1 9 15 0 1 9 0 15 13 1 15 9 0 0 13 1 12 9 0 2
88 7 7 15 1 9 0 14 13 9 9 9 0 7 9 15 1 9 0 7 1 9 15 1 9 0 0 1 9 9 7 0 9 2 7 9 9 0 8 0 1 9 0 2 7 9 8 7 9 15 9 9 9 0 7 9 2 9 0 2 2 7 13 1 9 0 9 8 8 1 7 15 14 13 9 9 0 1 9 0 0 1 9 15 13 1 9 12 2
40 7 13 8 7 15 14 13 15 9 8 8 1 9 14 13 14 13 1 9 9 2 7 3 9 8 8 8 8 8 8 8 14 8 7 13 7 8 1 9 2
51 2 2 9 1 9 8 8 2 7 13 8 8 8 7 3 9 1 9 0 7 9 7 9 1 9 1 9 9 9 0 7 9 9 1 9 2 8 9 9 0 1 9 0 1 9 0 0 1 9 0 2
46 7 13 9 0 0 1 10 9 2 7 1 15 9 15 2 1 9 9 9 9 0 1 9 9 0 1 9 0 7 9 9 7 9 9 2 7 3 9 0 1 10 9 2 1 15 2
10 2 9 1 9 9 7 9 15 0 2
15 2 9 1 9 9 1 9 7 9 9 1 15 1 15 2
25 2 9 1 9 9 1 9 15 1 9 9 1 9 0 1 9 9 0 1 9 0 7 9 0 2
25 2 9 1 7 9 9 0 13 1 9 9 1 9 0 7 9 9 0 1 9 1 9 10 9 2
53 7 1 9 9 9 15 13 15 9 0 2 7 9 9 9 9 9 7 9 0 2 13 9 1 7 9 9 9 0 2 7 0 1 9 9 0 2 7 7 13 0 7 14 9 9 1 9 14 13 0 1 9 2
24 14 9 9 1 9 9 9 7 13 8 2 8 8 7 15 14 13 15 1 9 1 9 0 2
11 14 9 9 1 9 9 9 7 13 8 2
13 8 8 7 15 14 13 15 1 9 1 9 0 2
39 14 8 8 9 9 0 7 14 13 9 9 0 1 9 0 8 1 9 0 7 0 1 13 7 9 0 1 9 1 9 15 7 9 9 15 1 0 9 2
12 9 13 9 0 1 12 12 9 1 9 1 15
25 13 9 8 8 9 9 9 1 9 9 7 15 13 9 12 12 9 1 9 9 0 1 9 9 2
33 13 1 9 9 9 0 12 2 12 7 9 13 9 0 9 15 1 12 12 9 13 1 9 10 9 7 14 13 3 9 1 15 2
19 1 9 15 13 9 8 8 9 9 1 9 9 9 0 1 9 9 0 2
20 13 9 1 9 9 9 9 9 0 1 9 0 7 0 0 1 9 9 0 2
34 7 13 1 9 9 0 1 9 9 0 0 9 1 9 9 0 1 9 9 0 1 10 9 7 9 15 1 9 0 7 0 1 9 2
7 9 1 9 0 1 9 0
33 13 8 8 8 8 9 9 9 0 0 7 15 14 13 1 9 0 1 9 9 9 0 1 9 9 0 1 9 9 0 1 9 2
48 7 13 9 7 15 13 1 9 9 9 9 1 13 15 13 9 1 9 9 7 9 1 9 0 7 9 13 7 9 0 13 0 9 7 13 1 9 9 0 0 9 1 9 9 1 9 0 2
40 7 13 8 8 7 15 3 9 9 0 1 9 0 0 0 1 9 8 1 9 0 1 9 7 15 14 13 1 2 15 8 8 15 9 0 7 13 9 0 2
45 7 13 1 9 1 9 2 1 15 12 9 9 7 15 9 9 9 0 7 13 1 9 9 1 9 1 9 9 1 9 7 9 9 0 1 9 9 0 7 9 9 1 9 0 2
24 7 13 2 8 9 10 9 1 9 0 2 7 15 8 8 1 9 15 9 9 13 9 15 2
46 7 13 9 1 9 8 9 2 7 15 13 7 15 7 13 1 10 9 0 7 7 15 1 9 0 1 15 15 9 15 13 1 15 9 0 7 9 0 0 1 15 13 1 9 9 2
8 9 0 1 9 1 9 9 0
17 13 9 0 9 0 1 9 9 1 9 1 9 7 9 9 0 2
23 0 13 9 1 15 1 9 9 9 9 7 9 9 0 1 9 9 9 0 1 10 9 2
38 7 13 7 9 9 9 0 1 8 0 13 9 1 9 1 9 9 1 9 2 1 9 10 13 1 9 9 0 1 9 2 1 9 0 1 9 15 2
36 7 13 0 1 9 9 9 9 0 1 9 2 7 9 9 0 1 9 9 2 7 14 13 9 1 9 0 1 9 7 13 9 1 9 0 2
76 1 9 13 8 8 8 9 9 9 7 9 1 9 0 7 9 9 0 13 1 0 9 9 1 9 0 2 0 1 7 15 7 13 9 0 0 1 9 9 1 9 9 0 13 1 12 5 1 9 9 0 0 1 0 9 0 2 7 14 10 9 0 1 9 0 2 7 8 1 9 9 9 0 9 0 2
56 7 13 8 8 7 9 9 0 13 9 9 9 15 9 13 0 7 9 0 8 13 13 7 13 1 10 9 9 9 0 1 9 9 0 7 9 9 2 9 1 15 13 1 15 1 9 9 8 7 9 0 1 9 9 0 2
90 7 1 9 9 0 1 9 9 0 0 9 13 8 8 8 7 15 14 9 1 9 1 9 1 9 2 0 15 9 9 0 1 9 7 9 7 9 8 8 13 8 8 0 7 0 9 2 7 0 15 9 9 9 0 8 8 13 1 9 0 0 9 2 0 1 7 9 3 13 9 0 2 7 1 7 7 9 14 9 7 13 1 9 9 0 1 9 9 15 2
17 7 1 9 15 13 8 8 8 9 9 9 0 1 9 9 0 2
61 14 9 9 8 0 1 9 9 0 13 1 0 9 2 7 13 8 1 9 9 1 0 15 7 9 9 9 9 0 1 9 15 0 2 13 1 9 9 7 9 0 1 9 0 1 15 2 7 13 1 9 9 1 9 9 15 13 9 8 0 2
76 7 1 9 9 9 9 0 1 9 0 13 8 8 8 7 9 9 0 1 9 9 9 15 7 14 13 14 9 0 0 7 14 13 1 9 1 9 0 2 7 1 3 13 9 0 1 9 9 15 0 0 1 9 1 9 10 9 1 9 15 13 8 8 0 9 1 9 9 15 14 13 1 9 10 9 2
15 14 8 8 8 9 9 9 9 8 1 9 9 9 2 2
57 7 13 7 8 0 14 13 0 8 8 1 9 0 2 7 9 1 15 9 9 0 15 13 1 15 9 0 1 9 0 2 7 15 13 1 15 1 9 9 0 7 9 1 9 0 1 9 0 7 1 7 9 9 9 0 0 2
17 7 13 1 9 0 8 8 8 9 9 9 8 1 9 9 0 2
34 0 7 9 9 8 8 0 1 9 9 0 14 13 2 7 7 9 10 1 9 7 9 9 13 2 9 1 9 9 9 1 9 9 2
71 7 13 0 2 7 13 15 1 9 9 9 0 1 9 0 2 7 13 9 0 9 2 0 0 2 15 14 13 1 12 12 9 2 7 1 0 7 9 9 13 0 1 9 0 1 9 1 9 0 2 1 1 7 15 1 9 9 13 9 9 0 0 13 1 12 1 12 12 9 3 2
54 7 13 8 8 8 7 15 1 9 0 2 13 3 9 1 9 0 1 9 7 9 9 7 9 9 15 1 9 1 9 9 9 0 1 9 9 2 8 8 0 9 13 2 7 9 1 15 13 9 9 1 9 9 2
48 7 13 8 8 7 15 14 13 9 9 9 0 1 9 1 9 15 2 7 9 1 10 9 1 9 9 9 0 1 9 0 2 15 13 7 9 1 15 9 0 1 9 0 9 1 9 0 2
8 9 13 1 9 9 0 1 9
63 13 9 9 0 0 1 9 15 9 9 0 1 9 1 9 9 1 9 9 0 1 9 9 3 7 13 9 1 0 9 9 0 9 15 1 9 1 9 1 9 0 7 0 1 9 9 1 9 9 2 0 1 9 0 7 0 7 0 7 9 7 9 2
48 7 13 8 8 9 9 7 9 9 9 0 0 7 3 9 0 13 1 9 1 9 9 2 0 7 9 0 1 9 9 7 7 9 14 13 9 9 0 1 1 9 9 0 1 9 15 0 2
40 7 1 9 15 13 8 2 8 8 9 9 9 9 0 7 9 9 1 9 9 14 9 1 15 2 0 1 7 3 12 12 9 1 9 13 1 15 13 15 2
36 13 15 1 9 15 13 9 9 0 9 9 9 1 9 9 0 0 1 9 7 9 1 9 9 1 9 9 9 0 1 9 0 7 9 0 2
46 7 13 9 9 1 9 0 1 9 0 7 9 9 0 7 9 9 0 7 9 9 7 9 0 1 9 9 7 9 7 9 1 9 0 7 9 0 1 9 9 7 9 9 0 0 2
46 7 13 9 9 1 9 0 1 9 9 7 9 7 9 9 0 9 9 1 9 0 0 1 9 9 0 9 9 1 15 1 9 9 7 15 1 9 1 9 9 9 0 7 9 0 2
99 7 13 9 9 0 14 13 9 12 2 12 9 0 0 1 9 7 9 1 9 9 7 15 13 9 1 15 9 9 0 0 7 9 9 1 9 9 0 1 9 1 9 9 9 1 9 0 2 7 7 9 9 0 1 9 9 1 9 9 15 1 9 9 9 1 9 0 1 9 9 1 9 0 1 9 9 7 9 0 7 9 9 7 9 0 1 7 13 9 0 1 9 9 9 7 9 10 9 2
11 9 0 1 9 9 9 0 13 1 12 9
31 13 9 8 8 2 9 9 7 9 0 0 2 7 15 13 0 9 9 1 9 0 1 9 9 0 1 8 9 12 0 2
38 7 13 9 1 9 15 1 9 9 9 1 9 0 1 9 0 0 9 12 2 12 0 7 15 14 13 9 1 9 7 9 10 9 1 9 9 0 2
44 7 13 0 7 9 9 0 0 1 9 13 9 0 14 9 1 15 2 0 1 7 15 13 9 9 7 9 0 7 0 13 9 0 7 9 0 7 9 1 9 7 9 0 2
51 7 13 9 9 7 9 0 7 3 9 1 9 13 9 1 9 15 1 9 9 9 9 1 9 0 0 7 9 9 9 1 9 0 7 0 1 1 9 9 0 0 1 9 13 9 9 0 1 9 0 2
51 7 13 7 15 13 9 1 9 0 7 0 7 9 9 9 0 1 9 7 9 9 0 7 9 9 9 0 7 9 9 7 9 15 7 9 9 0 1 9 1 9 0 1 9 9 9 0 1 9 0 2
54 7 13 7 9 0 15 9 9 7 13 9 0 1 9 0 0 1 9 12 5 7 7 15 13 7 13 9 0 1 9 0 0 1 7 15 1 0 7 13 10 9 7 13 1 15 1 12 1 12 5 1 9 0 2
28 7 13 7 9 0 15 13 15 9 13 9 0 1 9 1 9 0 0 1 1 9 9 7 9 1 9 9 2
73 7 13 8 1 7 9 13 1 9 9 9 1 9 7 9 0 13 8 0 0 7 9 0 7 9 9 7 9 0 7 9 7 9 15 7 0 9 9 7 9 0 1 9 9 8 8 1 1 9 0 7 0 0 0 13 15 9 9 1 9 1 9 1 9 9 9 0 1 9 0 1 9 2
7 12 9 0 1 9 9 9
14 13 9 0 0 9 0 1 9 9 9 9 9 2 2
70 1 0 10 9 9 10 13 9 1 9 0 7 0 1 9 9 9 7 13 9 0 0 1 9 0 1 9 0 1 9 9 9 1 9 9 0 9 7 15 13 9 15 1 9 1 9 7 9 1 1 2 0 2 7 13 9 1 0 9 13 9 15 9 12 2 12 0 12 5 2
44 7 13 14 13 1 9 0 9 9 1 9 0 7 0 1 9 9 9 14 7 9 0 13 1 9 9 9 1 9 0 1 9 1 9 9 9 1 9 9 7 9 9 9 2
63 1 0 9 15 13 15 9 3 9 9 9 9 0 1 9 9 0 13 1 12 9 9 12 2 12 0 1 9 0 1 9 9 1 9 15 0 1 9 9 7 9 9 7 9 9 9 9 0 9 10 1 9 15 1 9 0 9 1 9 1 9 0 2
37 7 13 8 8 9 0 1 9 0 0 9 9 1 9 9 1 9 15 2 9 9 7 0 9 1 9 9 9 0 9 1 9 9 15 1 9 2
35 7 13 8 2 7 9 1 9 9 1 9 13 1 10 9 3 7 7 9 9 9 7 9 13 9 0 1 9 9 9 1 9 9 0 2
45 7 1 9 15 13 15 9 1 9 0 3 9 9 9 1 9 9 0 1 9 9 9 2 7 13 9 9 1 9 9 1 15 1 1 13 9 0 1 9 9 1 9 0 9 2
97 7 1 9 9 0 7 14 13 1 9 0 1 9 9 9 9 9 1 15 1 9 15 13 15 1 9 9 7 13 9 0 9 9 12 2 12 2 12 0 1 0 9 9 12 5 1 12 5 1 9 15 13 15 9 12 2 12 0 7 1 9 9 15 12 9 7 13 0 9 1 10 9 9 9 0 1 12 5 14 7 15 13 7 13 9 9 9 1 9 12 9 7 13 1 12 5 2
87 7 13 2 0 2 14 13 9 0 9 15 1 9 0 1 9 7 13 1 9 1 12 12 7 12 12 9 1 15 12 7 12 12 9 1 9 9 9 15 13 15 1 9 9 12 2 12 0 7 13 15 1 9 9 9 12 2 12 0 7 13 9 10 9 0 9 15 12 9 1 0 9 9 12 5 7 13 0 9 12 5 7 0 9 12 5 2
31 14 9 0 7 0 9 15 12 12 7 12 12 9 7 13 2 0 2 1 9 15 1 9 12 9 13 13 15 1 9 2
6 9 9 0 1 9 0
16 13 9 0 7 15 14 13 9 1 9 0 0 1 9 0 2
72 7 13 9 9 0 0 8 8 8 7 9 0 9 15 14 13 1 9 9 9 0 7 1 15 9 1 9 9 8 8 7 1 9 9 15 0 1 9 0 2 0 1 7 9 9 7 9 0 13 7 13 1 10 9 1 9 15 8 8 7 13 1 15 9 1 9 9 15 1 9 0 2
78 7 13 1 9 15 1 9 9 9 9 0 9 12 2 12 0 7 15 13 0 9 9 10 9 7 9 9 15 0 7 9 9 15 13 1 9 15 1 10 9 14 9 7 13 1 15 9 1 7 13 1 9 0 7 7 13 1 15 9 9 0 2 7 7 0 1 15 14 9 7 13 7 15 9 9 9 0 2
34 7 13 8 7 15 13 9 1 9 9 1 9 7 7 13 9 1 9 8 1 10 9 7 14 13 9 0 1 3 1 9 9 0 2
7 12 5 9 1 9 9 0
42 13 9 9 9 0 0 1 9 15 13 15 9 0 1 9 7 0 1 9 9 0 15 13 15 9 1 9 12 5 1 9 0 7 13 9 1 15 9 1 9 0 2
17 7 13 7 9 13 1 9 0 9 9 9 0 1 9 12 5 2
20 7 13 9 9 9 8 8 9 1 7 15 1 9 9 9 9 7 9 15 2
48 7 10 9 13 9 9 9 9 0 1 9 9 9 15 1 9 9 1 9 0 1 9 9 7 9 9 1 9 7 9 9 0 1 9 2 1 9 9 9 0 1 9 9 15 13 15 9 2
66 7 13 9 8 7 9 13 1 9 0 1 9 7 9 9 0 7 13 1 9 0 15 13 1 9 15 7 1 9 9 15 13 9 2 0 1 7 9 9 7 9 15 13 1 9 0 13 1 9 0 2 7 9 9 13 10 9 1 9 15 7 13 1 9 9 2
9 12 9 1 9 9 9 1 9 0
14 13 9 9 9 2 9 0 1 9 0 1 9 0 2
15 13 9 1 12 9 1 7 13 12 9 1 0 9 0 2
18 7 13 9 9 1 9 1 12 9 1 9 9 7 12 9 1 9 2
51 13 9 8 9 9 0 0 1 7 15 1 0 9 1 9 13 9 9 1 9 1 9 0 2 7 13 8 9 9 1 12 9 2 0 15 9 9 1 9 9 8 1 9 0 7 13 9 1 9 0 2
32 7 13 9 9 9 9 0 7 9 9 0 7 9 9 9 1 9 7 9 9 0 2 7 9 9 9 0 2 9 9 9 2
34 7 13 9 3 9 9 1 9 9 1 9 9 2 1 9 9 7 13 0 1 9 7 9 9 9 2 7 9 9 1 9 0 9 2
18 7 13 9 0 1 9 0 1 9 2 7 13 1 9 9 9 9 2
27 7 13 9 0 9 1 9 9 13 1 9 9 2 1 9 1 9 9 0 1 9 9 9 1 9 0 2
32 7 13 8 7 9 0 1 9 0 15 9 1 9 0 0 1 9 7 9 0 2 7 9 9 1 9 7 9 1 8 9 2
16 7 13 9 1 9 9 1 9 1 13 9 7 13 9 9 2
7 0 9 1 9 0 1 9
22 9 9 0 0 13 13 9 9 0 7 13 1 15 0 7 0 1 9 9 0 2 2
32 7 15 1 9 7 9 0 0 9 1 9 13 9 1 9 9 7 1 9 15 13 0 1 9 1 9 9 9 15 0 2 2
33 7 7 13 9 14 13 1 9 12 5 1 9 0 0 7 0 9 7 0 7 14 9 15 13 9 15 9 10 9 1 9 0 2
15 7 14 14 13 10 9 1 9 0 0 1 9 0 0 2
28 1 9 13 9 8 8 8 9 9 9 1 9 0 2 7 9 9 1 9 0 0 7 0 9 8 8 0 2
44 13 1 7 9 0 1 9 0 0 0 9 1 9 9 15 0 0 1 9 1 9 1 9 9 9 2 1 9 7 9 9 0 13 7 9 0 1 9 0 13 1 9 0 2
17 7 1 9 9 0 1 9 0 7 9 0 0 1 9 7 9 2
5 8 3 9 0 2
15 9 13 1 9 9 7 8 7 15 13 1 9 9 0 2
46 13 1 15 7 9 0 0 0 9 0 1 9 2 7 1 15 12 12 9 9 1 9 15 2 13 9 15 1 9 9 1 9 0 7 9 7 1 9 9 10 9 1 9 1 9 2
31 8 8 1 9 0 13 9 8 8 8 7 9 9 13 1 9 9 1 9 7 9 7 15 15 13 9 1 9 9 0 2
8 7 7 8 1 9 0 0 2
28 8 8 7 15 1 9 1 9 9 1 9 0 7 14 9 7 1 9 9 0 7 15 9 0 1 9 0 2
21 8 8 1 9 8 8 9 0 7 15 7 9 9 0 1 0 1 9 1 15 2
72 7 9 9 1 9 9 1 9 9 7 9 0 1 0 9 1 0 1 9 9 1 9 0 7 9 9 9 0 1 9 7 9 10 9 13 1 9 0 3 1 9 9 9 0 2 7 1 15 13 8 8 1 9 9 0 1 9 2 8 1 15 7 9 0 9 9 9 0 1 9 0 2
44 9 15 13 9 0 1 9 0 9 1 9 0 2 7 9 0 13 1 15 12 9 0 1 9 2 7 1 15 9 9 0 7 9 9 9 7 9 9 1 9 9 9 0 2
79 1 9 15 13 8 8 2 9 9 9 9 2 7 9 0 0 13 0 1 9 0 9 2 0 7 9 9 1 9 0 9 1 9 1 9 1 15 2 8 8 7 9 0 13 9 1 9 9 1 9 1 1 12 9 7 12 12 9 7 12 9 7 12 9 2 14 1 9 7 14 13 9 1 12 9 1 9 0 2
9 7 13 7 9 9 1 9 9 2
48 7 15 13 9 1 9 9 15 0 2 14 1 9 1 9 9 7 15 0 9 9 1 9 9 9 7 13 7 15 14 13 9 9 9 0 1 0 9 1 9 1 9 9 1 9 9 0 2
25 14 8 8 2 9 0 2 7 13 7 9 9 1 10 9 1 9 7 9 0 0 2 9 9 2
63 0 7 3 9 0 0 7 3 9 1 9 0 2 7 13 9 15 9 9 0 1 9 0 9 2 7 7 10 9 13 9 0 1 9 0 2 1 9 1 7 9 9 0 9 0 1 9 9 1 9 0 7 7 9 0 0 13 9 7 9 9 0 2
26 7 13 9 7 13 9 9 15 3 7 15 14 13 1 12 1 9 7 7 14 13 7 15 14 13 2
40 14 1 9 1 9 0 7 13 8 8 7 9 0 1 15 9 0 1 9 2 7 7 13 9 7 13 1 9 0 9 2 7 14 9 13 7 13 1 15 2
19 7 7 13 7 15 1 9 0 2 12 9 0 2 13 9 1 9 0 2
31 7 13 13 9 0 7 13 7 9 1 9 0 13 13 2 7 13 15 1 9 9 1 9 0 7 3 9 9 1 9 2
38 15 1 9 9 0 7 0 1 9 9 7 15 9 0 2 7 1 9 15 13 1 9 7 9 9 9 9 0 2 13 15 1 9 9 1 9 0 2
24 9 9 9 7 13 9 1 9 3 7 15 13 0 1 9 9 9 9 7 15 13 9 15 2
9 12 12 9 9 1 0 9 1 9
98 13 9 8 13 1 15 2 9 9 2 7 9 0 0 9 9 1 9 13 1 12 5 1 9 9 13 1 12 8 9 1 9 9 0 12 0 1 9 12 8 9 1 9 8 8 7 12 8 9 1 9 12 9 0 1 9 0 1 9 7 9 2 0 2 0 1 9 12 8 9 1 9 7 12 8 9 9 7 12 8 9 9 9 7 12 8 9 1 9 7 12 8 9 1 9 9 0 2
44 7 1 9 15 13 9 9 9 15 1 9 9 0 15 1 9 0 15 13 1 15 10 9 9 9 1 9 1 9 7 9 9 1 9 9 1 8 1 10 9 1 9 0 2
47 13 9 2 8 0 1 9 2 1 9 9 1 7 9 0 0 1 9 0 1 0 1 9 1 9 9 0 1 9 13 12 9 0 1 2 9 0 2 7 2 8 1 9 7 9 8 2
11 12 12 9 9 15 1 8 7 8 7 8
63 13 8 8 9 9 9 0 0 7 9 0 1 9 7 9 1 8 7 8 7 8 13 9 0 1 9 0 0 7 9 9 0 1 9 12 1 9 0 12 13 1 12 8 8 1 9 1 12 5 1 9 9 1 9 0 7 13 9 1 12 8 8 2
45 13 7 3 0 1 12 8 7 9 0 1 9 7 9 12 1 9 9 9 0 7 9 9 9 0 7 0 7 9 0 7 0 7 9 9 1 9 1 9 9 0 1 8 2 2
46 7 13 8 7 9 13 1 9 9 9 1 9 9 0 1 9 9 9 0 1 9 0 7 3 9 9 0 1 9 0 7 9 9 1 9 12 13 1 9 9 0 1 12 9 3 2
33 7 13 8 1 7 8 15 0 9 0 1 9 1 9 0 7 8 1 0 9 0 1 9 7 8 13 1 0 1 9 0 0 2
10 9 9 0 2 9 9 13 1 9 0
25 13 9 8 8 9 9 0 9 9 1 9 9 0 1 9 12 5 1 9 0 0 1 9 0 2
41 13 8 7 9 9 13 1 9 0 9 1 9 9 7 9 1 9 2 7 13 1 9 0 9 12 2 12 0 1 7 9 1 9 9 14 13 1 9 9 9 2
43 13 9 7 9 9 1 9 9 15 1 9 0 1 9 9 2 14 13 1 9 9 1 9 0 0 1 9 0 2 7 7 15 14 13 9 1 9 9 15 9 1 9 2
24 7 13 8 7 15 13 0 9 9 1 9 9 0 1 9 1 9 8 7 9 0 1 9 2
47 7 13 9 8 8 9 9 9 9 9 1 9 0 2 7 9 14 13 0 1 9 0 1 9 9 9 9 2 7 13 9 9 12 1 9 2 7 14 13 9 9 0 1 9 9 9 2
25 7 13 8 9 9 0 1 9 9 9 9 1 9 9 2 0 1 7 10 9 0 1 9 9 2
8 9 9 9 9 0 1 9 0
68 13 9 9 0 1 9 0 12 1 9 1 9 0 8 1 9 9 2 7 1 9 15 13 1 15 9 9 0 8 2 1 9 12 5 1 9 0 1 9 9 7 14 13 9 9 1 9 12 12 9 2 12 12 9 2 9 1 12 12 9 12 12 9 1 9 0 12 2
44 14 1 8 9 1 9 7 14 13 9 9 9 2 9 0 2 9 0 1 8 9 15 13 9 15 12 5 7 13 12 12 9 9 1 12 8 9 1 9 0 12 2 12 2
51 7 13 10 9 0 1 9 1 9 8 9 0 1 9 1 12 8 9 1 9 9 15 12 5 0 1 9 0 8 8 7 9 9 0 1 12 8 9 1 1 13 9 9 0 1 9 1 12 8 9 2
25 1 9 0 13 9 9 0 1 9 12 12 9 1 9 1 9 9 9 9 0 1 12 12 9 2
35 7 1 8 9 0 1 9 9 0 7 14 13 9 9 0 1 15 1 9 9 0 1 12 8 9 9 1 1 12 8 9 1 9 12 2
119 7 13 9 9 9 2 0 0 2 9 9 9 15 1 9 12 5 7 13 12 12 9 2 12 12 9 2 9 1 1 12 12 9 1 9 0 2 13 10 9 1 9 1 9 1 9 0 1 9 9 0 1 12 12 9 2 12 12 9 2 1 9 12 5 0 1 9 8 7 9 9 0 1 12 12 9 1 9 9 12 5 7 13 9 9 9 1 9 9 1 15 9 9 9 9 0 1 12 12 9 1 12 9 7 9 1 9 9 1 9 15 1 12 12 9 1 12 9 2
92 1 9 0 7 14 13 9 15 14 13 1 9 12 9 7 9 9 12 12 9 2 1 8 9 0 1 9 0 7 14 13 9 9 15 0 1 12 12 9 1 9 9 12 1 12 12 9 1 9 8 8 9 1 9 12 5 7 13 8 9 9 9 1 9 12 5 1 9 0 12 2 12 7 13 12 12 9 9 1 1 12 12 9 1 9 0 2 9 13 12 2 2
48 7 13 10 9 1 9 9 9 8 9 0 1 9 12 5 7 13 12 12 9 2 9 8 7 9 9 0 1 9 12 5 7 13 1 12 12 9 2 13 9 9 1 12 12 9 1 12 2
25 7 1 9 9 0 1 9 7 14 13 9 9 0 1 12 12 9 1 12 12 9 1 9 0 2
218 7 1 8 9 9 2 9 9 2 7 14 13 8 9 15 1 9 12 5 7 13 12 12 9 9 1 1 12 12 9 1 12 2 7 13 10 9 1 9 1 9 8 9 0 1 9 12 5 7 13 12 12 9 7 15 10 13 9 1 8 7 9 9 0 1 12 12 9 1 9 9 13 12 5 1 1 14 13 9 9 0 1 9 12 12 9 7 13 9 0 1 9 1 12 12 9 1 12 12 9 2 13 9 9 9 0 1 12 12 9 1 12 1 12 12 9 1 7 1 9 13 9 9 2 8 8 2 0 13 9 9 15 1 12 9 0 1 9 0 12 9 8 9 1 9 12 12 9 12 12 9 2 7 13 9 9 15 14 13 9 0 1 9 9 1 9 1 8 7 9 1 9 13 12 8 9 2 7 9 1 9 9 7 9 9 15 12 8 9 7 13 9 9 1 12 8 9 1 1 13 9 9 7 9 12 12 9 7 13 1 9 9 1 9 0 1 9 2
102 7 13 9 9 9 1 9 15 9 0 1 15 9 9 15 1 9 9 9 15 13 9 1 15 1 9 9 12 7 12 12 9 2 9 15 13 1 9 0 1 9 1 9 9 9 1 9 12 7 9 9 9 1 9 0 1 10 9 2 7 3 9 9 1 12 1 9 9 12 12 9 1 9 9 0 1 9 0 7 9 9 0 13 1 9 9 13 9 14 13 1 15 1 9 12 9 1 9 9 9 15 2
34 7 13 9 3 7 9 8 8 1 9 12 13 12 12 9 1 9 9 1 0 8 7 9 9 0 1 9 15 13 9 15 1 9 2
35 1 9 0 13 9 2 0 8 8 2 8 0 1 8 9 15 1 9 12 5 2 7 13 12 12 9 9 1 12 8 9 1 9 12 2
36 7 13 9 9 2 9 8 8 8 8 8 2 1 9 0 12 9 9 0 1 8 9 15 7 13 12 12 9 1 12 9 1 9 0 12 2
6 0 0 13 12 9 0
84 13 8 8 8 9 9 0 0 8 2 9 2 1 9 9 9 9 13 9 0 7 0 2 7 13 9 12 2 12 0 1 9 9 0 1 9 15 13 1 15 9 9 0 0 1 9 12 7 1 0 9 9 9 9 9 1 9 9 9 0 2 0 1 7 15 13 9 1 10 9 1 7 13 1 9 1 15 9 9 1 9 9 0 2
37 13 8 8 7 8 8 13 1 9 9 9 1 9 9 1 9 9 9 0 15 14 13 1 9 15 9 2 7 14 10 9 0 1 9 8 3 2
24 13 1 7 9 13 3 9 9 9 1 9 8 8 7 9 2 1 9 9 9 1 9 9 2
36 7 13 7 9 13 1 1 9 15 0 7 0 1 9 9 0 1 9 0 7 9 9 1 9 2 1 9 9 0 0 1 9 1 9 0 2
20 9 2 9 9 13 15 9 9 1 9 9 7 9 9 0 1 9 9 15 0
48 13 9 9 7 9 0 1 9 9 9 9 0 0 1 9 0 9 1 0 9 7 9 13 2 7 1 9 9 9 0 1 9 0 0 7 9 9 9 9 9 15 14 13 1 1 12 9 2
108 7 1 9 9 0 1 0 0 8 8 1 9 1 7 9 1 9 15 0 0 1 9 9 9 9 7 14 13 1 9 15 1 9 0 7 9 15 9 9 0 0 1 9 15 9 9 0 7 9 1 9 9 9 0 0 14 3 9 7 9 7 9 14 7 9 13 7 9 9 9 0 0 1 9 15 1 9 1 9 9 15 0 7 7 9 9 1 9 0 1 9 9 9 1 9 9 1 9 9 9 15 13 1 15 9 9 0 2
18 7 13 1 9 9 9 1 1 12 1 12 1 9 1 9 12 0 2
80 1 9 0 13 9 1 7 9 9 7 0 9 9 9 9 0 7 9 9 1 9 0 14 13 1 15 9 15 0 1 9 0 0 1 9 9 0 7 8 15 13 1 1 12 5 1 9 9 9 0 2 7 7 9 15 13 9 8 1 9 9 0 1 9 0 15 13 1 0 9 1 9 0 0 1 1 12 12 9 2
25 7 13 0 0 8 8 7 13 9 1 9 7 9 0 1 9 0 7 7 13 9 9 8 8 2
53 7 13 7 9 9 0 1 9 9 1 9 1 9 0 1 9 9 15 8 9 9 9 1 9 0 15 13 8 9 1 15 1 9 0 1 12 9 2 7 13 9 15 1 12 9 1 9 7 12 9 1 9 2
73 1 9 0 13 9 0 1 9 0 1 9 9 0 1 9 9 1 9 9 1 9 0 1 9 1 9 9 0 13 9 9 9 1 9 9 15 0 1 9 1 9 9 0 1 9 1 9 7 9 9 9 0 1 9 9 9 7 3 9 9 1 9 0 7 9 1 9 15 0 1 9 0 2
41 7 13 9 9 0 0 0 8 8 7 9 9 9 1 9 9 9 0 0 1 9 7 9 1 9 9 1 9 9 9 9 7 0 2 14 13 9 1 9 9 2
61 7 13 8 7 13 0 0 1 9 9 1 9 1 9 1 9 12 12 9 2 7 3 7 13 1 9 10 1 15 1 9 2 0 7 13 8 0 1 9 9 8 0 1 9 9 0 0 1 9 9 2 7 1 0 13 9 1 9 9 0 2
57 7 13 9 0 1 9 9 7 9 9 9 9 0 9 8 8 7 9 0 9 15 14 13 7 13 9 0 7 9 13 1 9 9 9 0 1 9 7 9 1 9 0 1 9 9 9 9 1 9 9 9 1 9 9 7 9 2
33 7 13 8 7 13 9 9 0 1 9 0 1 9 9 0 1 12 12 9 2 9 7 10 9 14 13 9 7 14 13 3 9 2
41 7 13 8 7 9 9 8 0 14 13 9 0 15 14 13 9 1 1 9 0 1 9 12 15 13 1 9 12 1 12 1 9 9 7 9 1 9 0 1 9 2
77 7 13 9 9 9 7 9 14 13 9 0 1 9 0 2 7 14 13 9 1 9 15 1 9 9 2 7 13 7 9 1 9 7 9 13 1 9 0 7 14 13 0 1 9 1 9 2 7 13 1 7 9 9 13 1 12 9 1 9 7 12 9 1 9 7 7 9 15 1 9 9 0 14 13 12 9 2
12 8 13 8 9 9 9 1 9 1 1 9 0
64 13 9 9 0 8 8 9 15 9 0 8 8 1 8 9 12 2 12 0 1 7 15 2 0 9 2 0 1 7 15 13 9 1 9 9 8 1 9 15 1 9 1 9 0 1 9 0 0 1 9 9 1 9 7 9 0 7 1 9 9 9 8 8 2
62 7 13 8 1 9 1 9 0 7 9 13 9 9 9 0 2 0 1 1 9 0 2 8 8 0 8 8 8 8 0 1 9 13 2 9 9 8 8 2 7 9 15 0 8 8 2 8 8 2 2 8 1 9 9 1 15 0 1 9 9 15 2
101 7 13 8 1 7 9 1 9 9 1 9 14 13 9 1 9 9 9 15 1 8 8 2 8 8 8 0 7 13 8 2 2 0 7 9 0 2 0 1 15 2 7 0 13 9 10 9 8 8 7 13 0 9 2 2 0 8 2 9 0 2 2 0 7 9 1 9 0 7 0 14 13 0 2 0 1 9 15 1 7 13 1 9 1 9 8 7 8 2 0 1 15 13 15 9 9 1 9 1 9 2
93 7 13 7 15 13 1 9 15 7 1 9 15 0 1 9 8 9 9 0 8 8 15 13 8 9 1 9 2 7 7 15 13 9 1 9 1 9 15 13 15 9 8 0 1 9 15 1 7 13 9 9 1 15 2 1 9 0 7 0 7 1 9 0 2 2 0 9 0 1 10 9 2 9 9 9 2 1 15 8 13 9 9 15 1 9 1 9 2 9 15 0 2 2
8 9 13 9 9 2 9 9 2
21 13 9 1 9 9 0 9 9 13 2 9 9 2 13 15 9 0 1 9 9 2
41 7 13 9 9 0 1 2 9 0 2 9 8 8 7 9 14 13 15 9 0 7 0 13 1 9 9 7 14 13 1 9 9 15 14 13 9 12 2 12 0 2
58 7 13 9 0 1 9 8 8 8 9 0 9 12 2 12 0 13 15 2 1 9 9 8 2 9 15 9 0 8 8 7 0 0 8 8 2 7 13 9 9 0 2 7 13 7 9 15 13 1 15 13 1 9 0 1 9 9 2
15 9 0 0 7 12 12 9 1 9 7 9 12 0 1 8
46 13 9 0 13 1 9 9 12 2 12 0 1 7 1 12 12 9 0 2 14 13 1 9 2 7 7 0 1 9 9 1 9 0 0 2 7 7 12 5 1 0 9 0 1 9 2
55 7 13 9 2 9 0 1 9 0 2 15 13 15 9 9 0 0 1 9 1 9 9 0 2 7 13 2 8 8 2 1 9 1 15 2 0 1 9 12 9 8 1 9 0 1 9 2 13 9 12 5 1 10 9 2
24 7 13 9 3 1 7 9 0 15 13 15 9 1 9 0 0 14 13 12 5 1 9 15 2
17 7 13 9 2 8 13 1 9 8 8 9 0 1 9 9 0 2
31 7 12 5 1 9 13 1 9 1 9 7 9 2 7 12 5 1 9 7 9 2 7 12 5 1 9 12 5 1 8 2
38 7 13 1 7 9 0 13 9 0 1 9 0 1 9 2 7 13 9 9 12 5 1 9 9 1 9 12 5 1 9 7 9 7 12 5 1 9 2
35 7 13 9 1 9 9 9 1 9 1 9 0 1 9 9 9 1 9 1 8 0 7 9 9 9 1 9 7 9 9 0 7 9 9 2
26 7 13 9 9 9 0 0 9 0 1 9 9 0 7 9 9 7 9 0 0 9 7 9 9 9 2
13 9 9 13 9 2 9 0 9 2 1 9 2 2
2 1 9
40 1 9 15 0 1 9 15 1 9 9 15 9 0 2 13 9 9 2 9 9 2 9 0 9 2 2 15 13 15 9 0 0 1 9 7 13 1 9 0 2
20 7 13 9 9 1 9 15 1 9 2 9 2 9 0 1 9 0 7 0 2
33 7 13 9 9 12 9 0 13 15 9 7 9 0 13 1 9 15 9 0 1 9 9 15 13 1 15 1 9 9 8 8 8 2
98 7 13 7 9 0 15 13 15 9 9 13 9 1 9 0 13 1 15 9 8 0 1 9 0 7 0 1 9 0 2 1 9 0 0 9 13 1 15 9 9 0 0 1 9 0 2 7 13 9 8 8 0 1 8 10 9 2 7 13 1 9 15 7 9 15 1 9 0 0 7 9 1 9 0 1 9 8 1 9 8 8 9 9 1 9 9 0 1 9 1 9 9 7 9 1 9 0 2
30 7 13 9 9 1 9 7 15 13 9 9 1 9 9 1 9 7 9 15 13 9 9 0 2 7 13 1 9 0 2
18 7 1 9 1 9 9 8 7 9 13 0 1 9 9 1 9 9 2
24 7 13 9 9 9 0 1 9 2 9 0 2 7 15 14 13 9 10 9 3 1 9 0 2
9 9 1 9 9 9 1 9 13 9
36 13 9 1 9 1 9 9 1 9 9 9 9 9 1 9 15 1 9 9 0 1 9 15 1 9 13 9 1 9 9 0 7 9 15 0 2
54 13 9 1 9 1 9 9 9 9 1 9 9 9 0 1 15 9 1 9 15 1 9 0 2 1 1 15 9 13 1 9 9 0 1 9 7 9 1 9 0 2 1 9 1 9 0 1 15 1 8 1 9 0 2
119 7 13 2 8 2 7 15 13 0 9 9 9 1 9 9 7 9 2 9 15 9 9 0 7 9 2 2 1 10 13 9 1 9 0 15 13 1 9 12 2 8 9 1 15 1 9 9 9 15 13 15 9 0 1 9 9 0 2 7 1 9 15 9 9 9 7 9 7 9 7 9 9 0 8 8 7 9 0 1 9 14 7 13 8 2 8 8 2 9 9 9 2 13 1 9 9 9 9 1 9 1 9 9 2 7 13 7 15 14 13 1 9 1 9 0 7 9 0 2
45 7 13 2 8 2 1 2 9 2 0 1 9 9 1 9 0 2 13 1 15 9 9 0 2 7 13 9 9 9 15 1 9 2 7 9 9 0 2 7 9 9 0 2 0 2
45 7 7 9 15 13 9 0 7 2 0 0 2 1 9 0 7 9 2 1 9 1 9 9 1 15 1 9 15 2 0 2 1 9 9 1 9 9 9 0 7 0 7 9 0 2
38 7 13 9 0 7 9 1 9 9 1 9 13 1 9 1 9 9 9 9 1 9 7 13 1 9 9 15 1 9 0 1 15 1 9 1 9 0 2
34 7 13 7 2 9 15 13 1 9 1 9 15 1 9 0 2 7 13 1 9 1 9 9 7 9 15 13 15 9 1 9 0 2 2
33 7 13 1 9 1 9 9 2 7 9 0 15 13 1 9 0 1 9 0 2 7 13 9 9 15 1 9 1 9 9 0 0 2
77 1 9 0 2 13 9 8 8 8 2 9 9 2 1 9 0 1 9 9 8 2 8 8 1 9 9 9 8 8 1 9 9 0 9 7 9 2 1 9 1 9 1 9 0 1 9 0 7 9 9 7 13 8 8 9 9 9 1 9 2 7 9 9 9 7 9 1 9 9 2 7 9 9 9 0 0 2
13 7 13 9 1 9 9 9 1 9 9 1 9 2
38 13 7 8 8 1 8 1 9 9 7 9 9 0 2 0 2 2 7 9 15 1 9 9 9 0 1 9 9 7 9 0 2 7 9 9 0 0 2
13 9 13 9 1 9 0 13 1 9 7 9 7 9
33 13 9 9 0 1 9 1 9 0 2 13 1 9 9 9 7 9 7 9 1 9 0 0 1 7 13 15 13 1 15 9 2 2
74 7 13 7 13 9 0 2 15 9 9 0 1 9 9 2 2 9 9 1 9 9 0 7 9 9 13 8 1 15 7 13 2 2 7 13 9 9 1 9 13 15 2 9 9 0 2 2 0 9 1 9 2 13 9 9 15 1 9 9 9 9 0 8 8 2 9 1 9 9 2 7 9 15 2
26 7 13 2 9 2 1 9 1 9 15 13 1 9 9 13 15 9 7 9 1 9 9 1 9 0 2
28 7 13 12 9 13 1 9 9 8 2 13 9 1 9 1 9 9 9 0 1 9 1 9 9 15 1 15 2
24 7 1 15 13 1 9 9 7 9 8 2 13 1 9 9 15 0 1 9 13 15 1 2 2
20 7 13 9 15 7 9 15 1 9 9 7 14 13 1 9 9 1 15 2 2
1 2
51 7 13 9 9 9 9 8 8 13 9 0 9 1 9 9 1 9 7 9 1 15 2 7 13 9 9 1 2 9 0 2 8 8 9 9 1 9 9 13 1 15 9 13 1 9 13 15 0 1 9 2
35 7 13 8 1 9 0 7 13 1 9 9 1 9 7 13 7 9 0 1 9 13 15 7 13 15 7 14 13 1 15 15 13 1 9 2
18 7 13 8 9 9 9 1 9 9 7 13 1 9 9 1 9 15 2
23 7 7 13 9 1 9 9 13 15 8 9 15 13 7 1 9 2 9 1 9 0 2 2
52 1 9 9 1 9 0 2 7 2 13 9 9 1 9 9 15 7 13 1 15 1 9 9 7 9 8 8 2 8 9 9 13 8 1 15 7 13 7 9 15 1 9 15 7 13 1 9 9 1 9 2 2
21 7 9 9 8 13 1 9 9 7 9 9 8 1 15 15 13 13 9 0 2 2
22 7 9 1 9 9 9 7 9 8 8 1 10 13 1 15 1 9 9 8 8 2 2
11 7 9 0 1 9 7 9 1 9 2 2
10 7 9 8 9 7 15 0 0 2 2
75 7 13 9 2 14 13 0 9 7 9 0 7 9 1 9 1 10 9 7 9 15 2 7 14 1 10 9 13 9 7 13 9 15 1 9 7 9 2 7 7 15 13 9 9 7 9 7 9 1 9 0 2 0 1 7 13 15 13 1 15 9 1 15 9 7 1 15 9 7 13 9 9 9 2 2
106 7 13 2 7 13 9 1 9 9 9 1 10 9 15 14 0 1 15 7 15 13 9 1 9 2 7 14 13 9 15 13 1 15 2 2 7 13 9 1 2 7 10 13 1 15 9 1 9 1 9 9 0 2 7 9 9 0 7 9 1 9 9 7 9 15 1 0 9 7 9 9 1 9 7 9 9 15 1 9 10 13 15 2 9 15 13 0 15 13 1 9 10 9 1 9 15 1 9 9 10 9 7 9 15 2 2
3 9 8 8
20 13 8 8 9 9 9 13 2 14 9 1 7 13 9 9 0 1 9 0 2
19 7 14 9 1 9 7 9 9 0 9 8 8 13 1 9 0 7 0 2
28 7 1 9 9 1 9 7 9 15 0 9 1 9 7 9 0 9 7 1 9 9 0 7 9 9 1 15 2
21 13 8 8 7 9 9 1 9 0 9 2 7 7 9 15 1 9 7 9 0 2
18 1 9 15 13 1 9 9 9 9 9 9 15 13 15 0 7 0 2
32 7 1 9 15 14 13 9 1 9 9 7 13 1 15 9 1 9 7 13 15 9 1 9 1 9 13 9 15 1 9 0 2
50 7 13 9 8 2 1 9 9 7 9 2 7 1 9 1 9 15 13 1 9 9 0 1 9 15 13 15 9 1 12 7 1 15 13 13 10 9 1 9 15 1 9 1 9 0 7 9 7 9 2
66 7 13 7 1 9 15 14 13 9 1 1 10 9 2 7 14 13 1 15 2 1 9 9 15 14 9 1 9 9 10 13 1 9 2 7 7 9 9 13 1 9 13 1 9 9 2 1 9 7 9 0 1 9 0 15 9 9 9 7 15 9 14 13 15 15 2
10 1 9 2 13 8 8 9 9 15 2
18 7 9 9 8 8 13 9 0 9 1 9 9 1 9 1 9 0 2
20 9 15 0 1 9 1 9 12 9 14 13 9 9 1 15 7 9 1 15 2
39 7 13 7 10 9 14 13 1 0 1 9 9 9 2 7 7 8 13 2 8 2 7 2 8 2 0 1 9 9 9 15 14 13 15 2 9 9 2 2
30 7 1 9 9 15 13 8 8 7 8 8 13 0 9 9 0 1 9 9 1 9 7 9 7 9 2 9 0 2 2
94 13 8 8 7 8 15 13 9 1 15 1 8 2 7 1 9 9 8 2 15 0 1 0 1 10 13 7 13 8 8 8 8 8 8 8 8 8 8 8 8 8 7 9 15 2 7 15 13 1 9 7 9 10 1 12 9 14 13 2 7 7 9 0 0 1 9 14 13 1 9 0 2 7 7 9 9 1 10 9 14 13 0 1 9 2 7 14 1 9 0 0 1 9 2
39 13 8 8 9 15 2 1 15 13 9 1 9 9 8 7 9 1 9 9 1 9 1 9 9 13 9 7 13 9 0 2 9 7 9 10 13 1 9 2
6 9 1 9 2 14 8
78 9 9 9 9 0 1 9 1 9 9 0 1 9 0 1 7 1 9 0 2 13 9 9 9 1 9 8 14 13 1 9 1 9 0 1 8 2 1 9 9 15 13 9 0 1 9 0 13 1 9 9 9 15 15 13 8 8 2 9 9 9 0 7 13 15 1 9 9 0 1 9 9 0 1 9 9 0 2
97 7 9 7 15 14 9 0 1 9 2 8 8 8 13 2 7 0 0 14 13 2 7 9 0 13 9 9 7 15 14 13 7 13 9 0 1 10 9 1 9 8 8 1 9 9 1 9 9 2 13 3 1 9 9 1 9 7 0 1 9 9 9 2 7 15 1 13 14 13 7 1 13 9 1 9 9 1 8 13 0 10 13 1 15 1 9 0 14 3 7 13 9 9 8 9 9 2
60 14 9 15 13 1 9 7 14 13 1 9 9 2 7 9 9 14 13 1 9 9 1 9 9 9 13 9 7 13 9 9 7 13 9 9 1 9 2 8 8 14 13 7 13 9 14 15 13 15 15 2 7 13 1 9 14 1 9 15 2
42 7 9 7 9 13 9 9 2 7 15 9 9 1 9 7 9 7 9 7 13 10 9 14 13 1 9 0 1 10 15 0 1 9 9 7 9 7 9 9 1 9 2
47 9 1 9 13 9 3 2 7 9 9 7 9 9 0 1 9 7 9 1 9 0 2 7 1 9 0 7 9 7 1 8 7 9 15 7 9 15 15 9 15 13 7 13 1 15 9 2
52 7 8 1 9 14 13 7 13 0 8 8 9 9 1 9 15 2 7 14 13 1 15 7 13 1 8 9 0 1 9 7 13 0 1 15 13 9 9 15 1 1 2 7 0 1 15 13 9 9 15 0 2
36 7 9 0 13 1 15 15 13 1 9 2 7 9 14 14 13 15 13 15 1 9 1 9 9 7 9 1 9 9 9 1 14 9 9 0 2
44 7 7 8 14 8 1 9 0 7 13 1 10 9 2 7 14 9 8 12 13 1 15 1 9 1 9 9 0 3 15 2 15 13 9 9 9 0 1 9 0 1 9 9 2
16 9 0 13 9 15 1 9 1 9 15 13 15 9 9 1 8
60 13 9 0 9 15 7 9 15 1 9 15 13 9 1 9 9 1 8 2 7 13 9 1 9 1 9 9 0 1 9 9 12 2 12 1 9 8 8 8 7 9 13 9 0 7 0 0 2 7 7 9 15 15 9 1 9 7 1 9 2
17 7 13 9 8 9 9 9 0 0 1 9 8 0 1 9 9 2
107 7 13 8 8 8 9 9 0 7 9 0 13 1 9 9 15 9 2 0 1 9 9 1 9 0 2 0 2 8 14 13 3 9 0 0 0 7 14 13 3 9 0 2 7 1 3 13 9 9 1 9 9 0 0 1 9 9 0 7 0 1 9 0 2 2 7 13 9 8 8 1 9 7 9 9 9 9 0 1 9 9 0 0 7 9 15 7 9 9 0 1 0 0 1 9 9 0 0 1 9 0 2 1 9 10 9 2
26 7 13 8 9 8 9 9 9 9 9 0 7 0 1 9 9 9 1 9 0 7 9 9 0 0 2
50 7 13 1 9 9 9 0 1 9 9 9 7 9 9 0 1 9 0 15 13 1 15 7 3 9 9 0 1 9 9 9 1 15 2 7 9 9 9 0 0 7 0 1 15 9 15 1 9 0 2
6 9 13 1 9 0 9
20 13 9 0 1 7 9 13 1 9 2 9 9 0 1 9 2 1 8 9 2
9 7 13 8 9 1 9 9 9 2
12 9 13 7 9 13 1 9 9 1 9 9 2
40 7 13 9 0 7 8 13 9 2 0 2 1 9 1 0 9 2 7 15 1 9 9 15 13 1 7 9 13 1 9 9 9 9 0 1 9 1 9 9 2
20 7 13 9 9 0 14 13 2 1 9 0 2 9 1 9 0 1 9 9 2
24 7 13 7 9 1 9 0 13 1 9 9 1 9 9 0 1 9 1 9 2 1 9 9 2
29 7 1 9 13 9 9 1 9 9 0 2 15 13 9 9 2 0 15 13 1 9 9 15 1 8 7 1 9 2
9 7 1 9 2 9 13 9 9 2
24 9 0 1 9 2 2 13 9 0 7 9 0 0 1 9 13 9 13 1 9 0 9 9 2
16 7 13 8 1 9 1 9 7 9 1 9 9 1 0 9 2
41 7 13 9 0 1 8 2 1 9 9 1 9 2 13 1 15 7 9 1 9 1 8 13 9 1 9 8 9 13 9 1 9 9 0 1 9 9 9 9 0 2
32 7 1 10 9 2 13 9 0 0 9 1 9 9 0 2 7 13 9 9 0 1 15 1 9 8 1 9 0 1 9 9 2
58 2 2 9 0 7 13 9 0 8 0 1 15 7 13 13 9 15 13 15 9 1 9 9 2 7 13 9 0 7 15 13 15 2 3 2 9 1 9 0 0 1 9 0 13 1 9 9 1 9 1 9 13 1 15 9 1 8 2
28 7 1 10 9 2 13 9 1 9 0 1 8 2 9 9 9 9 0 2 7 15 14 13 8 8 9 0 2
28 7 1 9 0 1 9 2 13 9 9 9 1 9 7 9 9 0 0 2 1 9 9 2 15 13 1 9 2
30 7 1 9 9 9 9 13 9 1 8 7 15 14 13 15 0 9 1 9 2 7 7 15 14 13 1 15 0 9 2
25 7 13 9 0 7 15 14 13 9 1 9 9 0 1 9 1 0 9 2 1 9 9 1 9 2
34 7 1 15 13 15 10 9 2 7 14 15 7 13 3 0 9 1 10 2 7 14 9 7 0 9 0 14 13 1 9 1 9 0 2
14 9 9 12 9 0 14 13 1 12 12 9 1 9 9
24 13 9 13 1 9 9 0 1 9 7 9 9 9 0 13 13 12 1 12 1 9 9 9 2
40 7 13 9 15 13 1 9 7 13 1 9 9 0 1 9 9 0 0 1 9 7 9 15 13 1 9 9 0 2 7 0 9 12 9 0 13 12 12 9 2
19 7 13 9 9 0 12 12 9 1 0 9 0 7 13 12 12 9 12 2
59 7 13 9 7 13 9 9 0 12 12 9 1 9 12 7 12 12 9 9 12 7 13 9 1 9 9 0 0 1 9 12 5 0 1 9 0 1 9 0 7 12 2 7 1 9 9 9 0 1 12 12 9 1 9 0 1 9 0 2
19 7 13 9 0 9 1 9 0 1 12 9 1 9 7 12 8 1 9 2
53 7 1 9 9 0 0 1 9 9 12 14 13 9 1 9 0 1 1 12 12 9 2 13 15 9 1 12 12 7 9 1 12 12 7 9 12 12 7 9 1 12 12 7 9 1 12 12 7 9 1 12 12 2
52 7 13 7 13 9 9 0 12 12 9 7 9 12 12 7 8 12 12 7 8 12 8 7 9 12 8 3 8 8 12 12 7 9 12 12 7 9 12 12 7 9 12 8 9 7 9 12 7 9 12 12 2
53 7 1 9 9 2 7 14 9 15 13 13 12 5 1 0 9 0 9 12 2 14 13 12 5 9 12 7 12 5 9 12 2 7 14 13 9 15 13 0 9 9 0 1 8 0 1 9 12 5 1 12 5 2
25 7 14 13 9 12 1 12 1 0 9 9 0 7 9 12 5 7 9 7 9 1 12 1 12 2
39 7 13 9 7 9 9 0 14 13 9 1 9 9 0 2 7 14 13 9 1 9 9 7 9 7 9 9 7 9 9 9 0 7 9 8 2 9 2 2
51 7 9 1 9 7 14 9 9 8 15 13 9 15 12 5 1 0 9 0 2 1 9 9 12 2 14 13 12 5 9 12 2 7 14 13 9 9 0 7 9 9 0 7 9 1 12 5 1 0 9 2
39 7 13 9 7 9 1 9 0 7 9 9 0 7 0 13 1 9 9 9 0 1 9 0 9 2 7 3 1 9 9 9 9 7 9 1 9 9 0 2
37 7 13 0 9 0 1 9 1 9 9 9 7 13 8 0 7 9 0 1 9 1 9 9 0 1 9 7 9 7 9 7 9 7 9 7 9 2
40 7 13 9 1 9 8 1 9 9 0 9 1 9 9 0 2 7 13 9 0 9 0 1 9 0 1 9 9 2 7 14 13 1 12 1 12 1 9 9 2
13 9 1 9 0 0 7 9 9 0 1 0 1 9
51 13 9 9 8 8 1 9 0 9 12 2 12 0 2 9 9 15 9 15 9 9 1 9 15 8 2 0 1 9 1 9 9 7 9 9 9 0 2 7 3 9 9 1 9 7 13 9 14 13 0 2
19 7 1 9 0 13 7 9 0 13 9 12 2 12 0 9 1 9 9 2
19 7 13 7 9 15 13 9 13 9 0 1 9 9 9 0 1 9 0 2
39 7 13 9 7 9 1 7 8 14 13 9 1 9 13 1 7 15 13 9 9 1 9 15 2 7 13 7 1 10 9 14 13 0 1 9 0 1 15 2
25 7 13 7 9 0 13 7 9 13 9 9 0 2 9 1 9 0 15 13 1 15 1 9 0 2
18 7 0 7 15 9 0 15 13 1 15 8 9 9 1 9 9 0 2
43 7 7 9 15 1 10 9 13 1 9 1 9 0 1 8 2 7 13 7 15 13 3 7 13 10 9 1 9 1 9 13 9 1 1 9 0 0 1 9 0 7 0 2
45 7 13 9 0 1 9 9 9 8 8 8 7 9 13 15 9 0 9 15 7 9 9 1 9 9 7 9 13 8 0 2 1 1 9 9 9 0 1 8 8 8 9 1 9 2
195 7 13 9 9 9 0 1 9 9 9 8 8 1 9 15 1 7 15 13 1 9 1 9 0 9 8 8 7 9 1 9 1 9 9 1 8 7 9 15 1 9 15 8 9 13 8 1 9 7 9 13 8 2 7 13 8 7 8 2 13 9 9 0 1 9 15 7 7 13 9 1 10 9 2 2 7 0 7 9 13 0 3 1 9 2 2 1 9 7 9 9 9 1 10 9 2 1 0 7 13 1 15 9 0 2 7 13 0 2 2 7 13 9 13 7 8 13 0 1 9 9 1 9 15 7 15 14 13 15 1 9 2 2 2 7 13 2 2 13 0 7 9 9 1 9 13 0 1 9 9 15 9 9 9 1 9 1 1 9 9 0 13 7 14 13 9 15 9 15 9 0 2 1 9 7 8 15 9 1 9 14 14 13 1 9 8 8 1 15 13 9 9 9 2 2
64 7 13 8 7 13 8 1 9 9 0 0 1 9 9 9 15 0 1 9 12 13 1 9 15 9 9 1 9 9 0 1 9 1 9 7 7 13 9 1 9 1 9 0 1 9 2 7 14 13 9 0 9 9 1 9 9 7 7 0 1 9 0 2 2
52 14 0 7 13 7 8 2 13 1 9 14 0 8 8 2 7 7 13 9 1 9 7 13 9 9 2 7 7 13 9 0 2 1 9 9 15 7 13 9 9 7 9 15 1 9 0 1 9 1 9 2 2
14 9 2 1 9 1 9 1 9 9 9 1 9 1 9
40 13 9 9 1 9 7 9 2 1 9 9 13 15 9 0 1 9 1 9 9 13 9 13 9 1 15 13 1 9 13 1 9 9 15 13 15 9 1 9 2
39 7 13 9 1 9 7 9 8 7 13 1 9 9 0 2 7 13 7 13 9 2 14 13 14 9 9 0 1 9 1 9 7 9 9 9 0 0 2 2
59 7 13 9 9 0 0 9 9 2 7 13 9 0 1 2 9 9 1 9 1 10 9 2 7 13 9 9 9 1 7 15 2 9 0 2 2 9 2 7 15 9 0 1 9 13 9 15 9 0 15 2 15 13 9 9 1 9 2 2
56 7 13 1 9 0 9 1 9 1 15 2 2 2 2 2 7 9 1 15 13 1 9 2 13 9 9 0 2 2 1 0 9 13 9 0 0 9 1 9 2 15 9 9 15 13 1 15 9 1 9 0 1 12 9 0 2
38 15 13 9 9 1 9 0 0 1 9 1 12 9 0 2 7 15 9 9 1 9 9 0 15 13 9 0 1 9 15 1 9 13 9 15 9 12 2
18 7 1 8 9 13 9 0 9 1 9 9 9 1 9 9 0 2 2
30 7 13 9 1 9 9 0 13 9 0 2 2 15 9 9 0 15 13 1 9 9 9 0 1 9 9 7 1 15 2
25 7 15 9 9 0 15 13 1 9 9 7 9 15 7 13 1 9 0 1 15 15 1 15 9 2
12 7 15 9 9 9 0 15 13 1 9 9 2
18 7 15 9 9 0 15 13 9 15 1 9 9 1 9 9 9 2 2
17 8 8 2 9 9 13 1 9 1 9 15 8 9 0 1 9 9
64 13 9 8 8 8 8 1 9 9 8 8 8 7 15 2 13 1 9 7 9 7 13 9 0 9 0 0 1 9 9 2 9 9 9 2 1 9 8 9 2 0 14 15 1 2 9 2 1 9 7 9 0 1 9 9 9 1 9 9 1 9 7 9 2
73 7 13 8 8 1 9 9 2 8 1 9 9 9 15 13 1 15 9 0 0 2 8 8 2 1 9 9 0 2 1 1 9 15 0 0 2 1 8 1 9 9 0 1 9 9 2 1 9 9 15 1 7 9 9 9 2 7 13 15 1 9 10 9 2 7 7 13 2 1 9 9 2 2
46 7 13 2 2 8 8 9 9 2 1 1 10 9 2 13 1 9 9 9 0 7 3 0 9 0 1 9 2 8 1 9 9 9 7 13 8 9 1 15 1 9 1 9 15 0 2
60 7 1 7 15 13 1 9 1 8 7 9 2 13 1 9 15 9 3 1 9 9 0 0 1 9 0 7 9 15 7 9 1 9 1 9 15 0 2 7 1 15 9 1 9 0 3 7 13 15 1 9 1 9 7 9 1 9 9 2 2
41 7 13 8 8 7 2 8 15 9 9 1 9 7 1 9 9 7 13 9 15 1 9 0 7 9 0 1 9 1 8 7 1 9 9 13 0 9 1 15 2 2
45 7 13 2 14 13 15 14 13 9 9 1 9 7 0 0 15 13 1 9 2 13 15 1 9 15 2 7 7 13 1 8 7 8 7 9 15 1 9 0 15 13 10 9 2 2
10 9 1 9 0 1 9 0 1 9 15
30 13 9 9 9 0 1 9 9 8 8 9 9 1 9 15 1 9 9 9 12 2 12 0 1 9 0 1 9 0 2
34 13 9 9 9 9 1 9 0 2 7 9 15 1 12 12 9 1 9 9 1 9 12 1 12 12 9 1 9 0 1 1 9 0 2
19 13 9 1 9 15 1 9 9 1 9 1 9 0 1 9 9 9 2 2
15 7 13 9 1 9 0 1 9 0 7 9 1 9 15 2
16 7 13 9 1 9 9 1 9 1 9 10 9 1 1 9 2
18 7 13 7 9 1 10 9 14 13 1 9 0 7 9 1 9 9 2
20 7 13 9 8 1 9 9 0 7 9 0 13 9 9 15 13 15 8 8 2
22 7 13 13 1 9 0 7 14 13 1 9 9 0 1 9 1 9 1 9 9 0 2
31 7 13 9 1 9 15 1 9 9 1 9 9 15 1 1 9 9 9 0 7 15 14 13 9 0 1 9 0 1 9 2
12 9 8 13 9 1 9 9 0 1 9 1 9
51 1 0 9 0 1 9 9 1 9 9 0 1 9 1 9 9 15 7 9 15 0 1 9 0 2 13 12 9 9 12 2 12 0 9 1 9 9 0 1 9 1 9 9 0 1 9 9 9 9 0 2
47 7 13 9 9 9 9 8 0 8 8 15 13 12 9 0 1 9 9 0 2 0 7 9 1 9 10 9 13 9 1 9 9 9 0 1 9 15 1 9 2 7 15 8 1 9 0 2
85 7 13 9 1 2 9 0 2 1 9 1 9 9 0 0 1 9 15 9 12 2 12 0 2 15 14 13 7 9 0 0 1 9 2 15 9 0 0 2 7 7 3 0 1 9 7 9 7 9 0 15 13 1 9 9 2 7 7 14 13 1 9 7 7 1 15 13 7 15 1 9 9 1 7 13 9 9 1 9 9 7 4 9 2 2
53 7 13 8 7 2 9 0 1 9 8 1 9 9 0 15 9 1 9 7 9 0 2 7 9 9 9 9 15 2 7 3 1 9 9 0 7 9 9 9 9 1 9 2 0 7 15 9 9 13 9 9 0 2
65 7 13 9 7 9 15 13 9 15 1 9 14 13 0 1 9 9 2 7 9 15 9 9 9 7 9 9 1 9 9 7 9 9 7 9 9 0 2 0 1 7 9 14 13 0 1 0 9 0 7 7 9 15 13 3 1 15 13 1 9 7 13 1 9 2
77 7 13 9 9 1 9 9 0 7 0 1 9 7 3 9 7 9 7 13 1 9 8 8 8 8 8 8 8 8 2 7 1 0 8 8 8 8 8 8 8 8 2 7 1 0 0 8 8 8 8 8 8 8 8 7 1 9 8 8 8 8 8 8 8 8 7 1 9 8 8 8 8 2 8 8 8 2
19 9 9 2 2 1 9 8 9 9 7 13 1 9 9 9 1 9 9 2
21 13 9 9 9 8 8 8 9 9 0 2 7 1 9 8 9 9 13 9 9 2
39 7 13 9 9 2 7 13 9 0 13 1 9 9 0 13 9 15 1 9 2 7 14 15 1 9 15 1 10 9 13 1 9 0 0 1 9 0 2 2
46 7 13 9 9 1 9 0 1 9 15 9 12 2 12 0 1 8 8 9 0 0 2 1 7 9 15 14 13 1 9 9 1 9 15 14 13 7 13 15 3 1 9 9 9 2 2
5 7 13 9 9 2
17 8 8 14 8 8 8 8 1 7 8 1 8 8 1 9 0 2
8 8 9 0 13 1 9 9 0
34 13 8 9 9 8 8 1 9 0 9 15 1 7 13 10 9 0 9 1 9 0 1 9 9 0 1 8 7 13 0 9 1 9 2
37 7 13 0 7 9 9 13 7 13 9 15 1 9 9 0 7 8 9 15 1 1 0 9 7 0 2 8 8 7 13 9 1 8 13 8 8 2
38 7 9 1 9 9 2 9 9 0 2 1 9 2 13 9 9 7 9 1 9 9 0 7 13 9 0 1 9 2 1 9 15 9 0 0 1 9 2
11 9 1 9 13 7 8 13 1 9 15 0
61 1 9 9 0 1 9 0 0 13 9 1 9 9 9 15 0 1 9 9 9 8 8 8 1 9 9 0 9 9 7 7 8 13 9 0 7 9 9 9 1 9 9 15 13 1 15 2 0 8 9 8 13 9 15 0 7 14 13 9 9 2
46 7 13 9 1 9 9 1 9 15 13 15 9 0 0 8 8 8 8 7 9 0 1 9 9 0 1 9 9 12 2 12 0 1 9 9 9 9 13 9 9 0 0 1 9 0 2
26 7 13 9 9 8 8 9 9 0 1 9 0 7 8 13 9 1 9 15 0 14 1 9 9 9 2
20 7 13 9 8 8 8 9 0 8 9 9 1 9 9 1 9 9 9 15 2
15 9 0 1 8 2 9 8 8 7 14 13 8 9 1 15
28 13 8 1 9 9 0 1 9 9 8 8 8 13 1 15 2 9 2 9 0 1 9 9 13 9 9 9 2
47 7 13 8 1 9 15 9 0 0 8 8 2 7 13 9 0 1 9 9 9 2 1 9 8 9 2 7 13 9 1 15 7 13 9 13 1 9 9 1 9 0 7 15 9 15 2 2
5 15 9 15 2 2
18 15 9 15 2 7 13 15 9 15 15 14 13 7 13 1 15 2 2
25 7 13 9 0 1 9 1 2 9 2 7 9 0 13 1 9 7 9 9 2 7 14 13 0 2
34 7 13 1 9 0 9 15 7 8 13 9 1 7 15 13 9 1 9 10 9 1 8 2 7 13 9 1 9 0 1 9 8 8 2
11 7 14 13 9 9 9 9 0 1 8 2
36 7 13 7 9 1 9 0 3 1 9 0 0 1 8 1 9 15 13 9 0 9 15 1 9 1 9 0 1 9 9 9 0 1 9 0 2
16 7 7 9 9 15 14 13 9 9 1 9 0 7 9 0 2
42 7 13 9 9 0 1 2 9 2 7 9 0 13 1 9 9 1 9 15 9 0 1 9 1 9 1 9 2 1 9 7 9 9 0 14 13 1 15 1 10 9 2
39 7 13 7 8 2 13 9 9 14 0 7 14 0 2 7 9 9 14 13 9 0 1 9 15 1 8 7 1 9 9 9 15 7 9 15 1 9 2 2
42 7 13 7 9 0 14 13 1 9 9 2 9 7 9 15 13 9 1 2 9 9 9 9 0 1 9 0 2 7 15 7 13 10 9 14 13 1 9 9 0 2 2
12 9 9 13 9 9 1 9 9 9 9 1 9
37 13 9 8 8 8 9 9 0 7 9 9 9 1 9 9 9 9 1 9 9 9 9 1 9 2 7 13 1 7 9 0 7 0 13 1 15 2
42 7 13 9 8 8 2 7 9 13 1 9 9 0 15 13 15 9 9 2 7 9 9 0 1 1 9 9 9 9 9 8 2 7 9 0 1 9 9 9 12 0 2
30 7 13 10 9 14 13 9 9 9 7 9 9 9 9 1 9 9 9 1 9 2 7 9 15 1 15 1 9 0 2
35 7 13 9 2 1 9 13 15 9 9 1 9 0 2 7 9 13 0 9 1 9 0 1 9 1 9 0 7 9 0 1 9 9 9 2
12 9 9 9 2 8 2 9 0 1 9 1 9
21 13 2 8 8 2 1 9 0 1 9 0 1 9 1 9 0 1 0 1 9 2
78 7 14 13 9 0 2 7 13 2 8 8 14 13 10 9 1 9 9 13 12 9 1 9 7 13 1 9 1 9 8 8 8 8 8 1 9 9 9 9 1 8 2 9 9 0 2 7 13 8 1 9 9 0 9 1 9 1 9 9 9 15 13 8 8 0 2 8 8 1 9 14 13 15 9 1 9 12 2
24 7 13 9 9 8 8 7 2 8 8 2 13 9 0 2 7 15 13 1 9 9 0 2 2
53 7 13 9 1 7 9 2 8 8 2 1 10 9 1 9 9 0 13 9 15 1 9 1 9 0 1 0 2 7 1 9 7 9 9 9 13 12 12 2 8 7 9 9 1 9 0 15 13 15 9 0 0 2
12 9 0 13 2 12 12 9 9 9 1 9 0
23 13 9 0 7 9 9 9 1 9 9 0 13 1 12 12 7 12 12 9 1 9 0 2
44 13 9 15 13 15 9 8 8 9 9 9 1 9 9 8 8 9 9 0 1 9 1 9 9 1 9 9 9 1 9 9 7 9 8 0 7 0 1 9 9 1 9 0 2
75 13 9 1 9 9 9 1 9 1 9 9 15 1 10 13 1 9 9 9 1 9 1 9 9 7 9 1 9 9 7 9 0 1 9 9 7 9 7 9 1 9 9 9 9 9 1 9 0 1 9 0 9 1 9 9 9 7 9 7 9 1 9 15 7 9 9 15 1 10 13 9 0 7 0 2
53 7 13 1 9 1 9 9 0 7 9 9 1 9 1 9 0 9 1 9 1 9 1 9 9 1 9 9 7 9 9 7 9 1 9 15 7 9 9 9 9 8 9 1 7 9 9 7 9 8 7 9 9 2
9 8 13 9 9 1 9 1 9 0
33 13 9 2 9 0 2 1 9 8 8 2 1 9 9 9 7 9 9 0 1 9 9 1 9 1 9 9 0 9 7 0 9 2
30 7 13 2 2 15 9 8 9 1 9 9 1 9 7 9 9 15 9 9 1 15 7 9 9 7 9 1 15 2 2
20 0 1 7 10 9 2 13 1 9 15 13 9 15 1 9 7 9 15 2 2
31 7 13 2 2 13 8 13 1 9 0 2 1 9 7 9 2 7 9 7 9 2 7 9 7 9 7 9 7 9 2 2
17 7 15 15 9 15 7 13 15 9 9 1 8 7 9 2 2 2
36 7 1 9 7 13 1 9 10 9 9 1 10 13 9 1 9 7 9 15 2 1 8 7 8 15 13 9 9 7 9 7 9 0 2 2 2
4 9 9 9 0
34 13 9 0 7 0 1 9 1 9 9 9 0 0 1 9 9 15 13 9 9 2 9 9 9 7 9 9 7 15 13 1 9 0 2
66 7 13 9 0 1 9 7 9 0 1 9 9 0 1 9 2 1 9 9 0 1 9 2 7 9 15 1 9 9 15 1 9 1 9 15 9 1 9 9 15 2 1 9 9 9 15 1 9 9 0 2 7 9 9 7 9 0 1 10 9 1 9 1 9 9 2
41 13 9 9 1 9 0 1 9 0 1 12 9 2 7 13 1 9 1 9 9 0 7 0 2 7 9 1 9 7 9 2 7 9 9 2 7 9 0 1 9 2
15 7 13 9 9 0 13 1 9 0 1 9 0 1 9 2
43 7 13 9 0 9 9 8 8 7 15 14 13 9 9 7 13 1 9 1 15 8 2 7 9 9 1 9 2 7 9 1 9 9 1 9 7 9 7 9 9 9 9 2
12 8 2 0 13 9 0 1 9 7 9 9 13
102 1 9 1 9 9 9 0 8 8 9 9 1 0 2 1 9 9 2 9 1 9 15 1 9 15 1 9 1 9 0 2 13 9 0 1 8 7 15 14 13 1 9 0 1 9 0 0 1 9 0 9 0 1 9 2 7 3 1 9 0 2 2 9 13 8 13 1 9 15 0 7 15 14 13 7 13 9 1 9 1 7 13 1 9 9 15 8 8 2 7 14 13 9 9 7 9 1 9 9 1 0 2
55 7 13 9 1 9 8 2 1 9 9 9 15 2 9 0 13 9 2 1 9 7 9 2 15 13 1 15 9 0 0 15 13 9 7 1 7 8 7 9 0 0 8 8 13 1 0 1 12 5 1 9 0 1 15 2
76 13 7 8 8 13 7 9 15 13 1 9 1 9 13 1 9 15 7 13 0 1 9 2 7 15 15 13 15 9 9 8 8 1 9 15 7 9 13 9 0 1 9 8 8 7 7 0 13 2 9 0 2 1 10 9 2 7 14 13 9 15 2 7 13 9 9 2 15 13 9 9 10 9 1 9 2
36 7 13 9 0 9 1 7 1 9 9 0 8 8 9 9 1 9 2 9 2 15 13 15 9 15 1 9 9 8 0 9 2 9 0 2 2
66 7 13 1 9 7 8 13 1 9 15 9 9 7 15 9 0 1 9 9 0 7 7 9 15 9 2 9 0 7 0 2 1 9 9 13 9 1 9 1 8 2 1 9 9 15 1 7 2 9 2 14 13 1 0 9 1 9 9 1 9 1 9 0 2 0 2
55 7 1 9 9 9 0 8 8 9 7 9 14 13 1 9 8 2 7 13 1 15 7 13 0 0 9 1 9 9 9 2 2 0 7 9 0 0 13 7 9 1 15 9 2 9 9 9 15 13 15 1 15 9 0 2
8 8 13 1 8 9 0 1 9
33 13 9 0 0 1 9 0 1 7 9 0 8 8 15 14 13 8 1 9 0 0 2 14 13 1 15 9 0 0 1 9 9 2
48 7 13 10 9 9 0 1 7 15 13 1 9 0 14 13 9 0 1 9 0 1 9 9 2 7 9 10 1 9 0 2 7 9 1 9 0 2 7 9 0 1 9 7 9 9 9 0 2
127 7 13 2 9 2 7 9 0 14 13 1 9 0 8 8 1 9 8 9 0 1 7 13 8 1 15 9 9 9 0 13 1 9 9 0 15 13 1 9 2 7 7 9 0 13 9 0 1 9 0 0 1 9 9 0 1 9 9 10 9 15 13 1 15 9 9 9 1 9 9 7 1 9 0 7 0 1 9 9 9 0 13 2 9 7 15 13 9 1 7 13 10 9 7 13 9 9 9 2 7 7 9 0 0 1 10 9 1 9 1 9 9 0 7 15 13 8 9 1 7 8 14 13 1 9 3 2
13 9 0 0 13 1 9 9 2 1 9 9 9 0
71 13 9 0 0 0 1 9 9 0 9 2 1 9 9 9 0 1 9 2 7 13 10 9 1 9 9 0 0 0 9 9 0 1 9 1 9 15 1 9 12 2 7 15 13 1 9 15 7 13 9 1 9 9 15 13 15 9 0 8 8 1 9 1 9 2 8 8 2 9 0 2
39 7 13 9 0 1 9 9 8 8 15 13 9 9 9 9 0 7 13 1 8 9 9 1 9 9 15 9 9 9 1 0 15 2 7 13 9 15 0 2
30 7 13 8 1 9 1 9 8 8 9 1 0 2 7 9 0 0 1 9 9 1 9 9 9 9 0 1 9 2 2
29 7 13 9 8 1 2 9 0 2 1 9 0 8 8 7 9 15 13 1 9 9 15 0 1 9 9 9 9 2
28 7 13 2 7 8 8 7 7 8 8 13 7 13 10 9 4 3 9 0 7 9 9 9 1 9 15 2 2
18 9 1 9 9 9 0 1 9 9 1 9 2 9 0 1 9 9 9
36 13 9 7 9 8 9 9 9 1 9 0 1 9 0 0 1 9 9 9 0 2 8 2 13 9 9 1 9 9 9 0 1 9 9 9 2
23 7 13 9 7 9 2 8 2 14 13 1 9 9 9 1 9 1 9 9 1 9 0 2
43 7 13 9 1 7 9 14 13 0 1 9 0 1 9 9 1 7 13 9 1 9 9 9 0 1 9 9 9 9 8 0 0 7 15 15 13 0 1 9 9 7 9 2
42 7 13 9 1 7 9 9 0 1 9 9 9 1 9 9 9 13 1 9 9 0 1 9 0 2 0 1 7 9 14 13 1 9 9 9 0 7 9 9 0 9 2
51 7 13 8 8 9 9 9 9 9 1 9 9 0 7 9 9 9 1 9 9 9 0 1 9 9 9 14 13 1 9 9 7 9 9 9 0 7 9 14 13 0 1 9 9 0 1 9 1 9 0 2
42 7 13 7 9 9 9 1 9 9 9 14 13 1 9 7 14 13 1 9 1 9 9 1 9 0 0 15 14 13 8 9 0 1 9 9 1 9 0 7 9 0 2
62 7 13 9 8 8 9 0 1 9 8 1 9 9 9 7 9 9 9 1 9 9 9 0 1 9 9 9 9 1 9 15 7 13 9 0 9 0 1 9 0 7 14 13 1 9 9 9 0 1 9 2 9 15 13 0 1 9 9 1 9 0 2
60 7 13 8 8 9 0 1 9 0 1 9 7 9 9 13 1 9 0 9 0 1 7 13 9 3 7 13 3 1 9 0 2 13 9 9 15 15 9 1 9 9 7 13 9 9 1 9 9 13 1 15 9 7 7 1 9 1 9 15 2
24 7 13 7 15 13 1 9 0 8 7 9 7 9 1 9 9 7 1 9 9 1 9 0 2
60 7 13 7 9 13 13 0 9 0 7 13 1 9 2 0 1 7 9 9 9 9 1 9 9 9 13 1 9 9 9 1 9 1 9 0 7 13 9 15 8 0 1 9 1 9 9 9 1 9 15 7 14 13 9 15 1 9 9 0 2
54 7 13 9 8 9 9 9 1 9 8 1 9 9 0 7 13 9 9 9 0 1 9 0 0 1 9 0 15 13 1 9 0 0 1 9 9 7 9 9 1 9 9 0 15 1 0 1 15 7 13 9 0 0 2
10 9 9 1 9 13 1 12 5 1 9
38 13 2 9 9 7 9 9 9 2 0 1 9 9 0 2 9 12 2 12 0 7 9 9 0 1 9 13 1 12 5 1 9 12 1 12 1 9 2
10 7 13 9 9 12 5 1 9 12 2
19 7 13 9 9 1 9 15 1 9 2 9 0 1 9 9 7 9 2 2
4 9 9 13 9
65 9 9 9 1 9 2 13 9 9 0 13 1 9 0 7 13 9 15 1 9 13 1 12 2 12 5 2 7 0 7 9 15 14 13 1 10 9 9 9 9 9 1 9 2 7 9 9 15 1 9 0 8 8 0 2 7 14 14 13 2 9 2 9 9 2
72 9 8 0 9 0 9 9 9 2 13 9 9 9 9 1 9 0 0 2 2 13 3 9 1 9 9 1 9 9 9 9 7 7 3 9 1 9 9 9 0 1 8 7 1 9 9 1 9 9 9 1 8 8 8 7 13 7 9 9 9 1 9 9 9 0 1 9 1 9 1 9 2
10 13 7 14 13 7 13 1 9 0 2
13 1 0 13 3 15 13 9 1 7 13 9 0 2
91 14 9 8 9 8 9 9 9 9 2 7 13 1 9 0 15 9 9 9 9 0 1 9 0 2 7 13 0 9 1 9 9 9 8 7 14 13 8 1 9 0 7 15 13 7 9 13 7 14 13 1 12 5 1 9 9 14 13 1 15 9 9 1 9 10 9 7 1 0 7 13 9 1 9 9 0 7 9 9 9 9 1 9 0 9 1 9 1 9 9 2
35 14 8 8 9 9 9 1 9 0 9 0 7 13 7 13 9 9 0 1 9 0 9 1 9 0 13 1 9 0 7 9 1 9 9 2
87 7 13 0 2 9 13 0 1 9 9 9 9 0 15 13 9 15 12 12 7 13 1 12 12 7 7 13 1 9 9 1 9 15 9 9 7 15 7 13 9 9 1 0 9 7 14 13 15 13 7 1 9 0 7 9 0 7 14 13 7 7 13 9 9 1 9 7 15 1 9 12 12 9 9 9 1 9 9 0 13 9 9 9 15 12 12 2
9 8 13 1 9 9 15 0 1 9
18 1 9 13 9 1 9 0 1 9 13 7 13 1 15 1 9 2 2
62 13 2 9 9 2 7 9 9 0 13 9 1 9 0 2 13 1 15 1 9 0 9 9 1 15 1 0 1 9 0 1 9 9 9 1 9 9 9 0 1 9 9 1 9 7 9 0 12 15 1 0 9 15 1 9 9 0 1 9 9 0 2
45 7 13 9 9 7 9 0 0 7 13 9 9 1 9 0 13 1 9 1 9 9 0 0 1 9 9 0 15 14 13 1 9 1 9 9 1 9 0 7 13 1 15 9 0 2
19 7 1 9 15 13 9 8 8 9 9 9 0 2 0 8 9 0 0 2
33 7 13 1 7 9 13 10 9 1 9 12 7 15 9 0 15 13 1 9 1 9 0 1 9 9 1 10 9 1 9 1 15 2
21 7 13 9 8 1 9 1 8 9 9 1 9 2 9 1 8 9 0 0 2 2
31 7 13 7 9 0 1 9 7 9 9 8 7 9 9 0 0 14 13 1 12 5 1 9 9 0 7 13 13 12 5 2
46 7 13 9 9 0 14 13 1 9 0 1 2 9 9 2 1 7 15 1 0 9 9 1 9 7 9 0 1 9 9 0 0 2 13 1 9 1 9 9 1 9 9 9 0 2 2
15 7 15 1 9 9 12 0 1 9 9 1 9 9 0 2
33 7 13 7 9 9 8 8 13 10 9 1 9 1 9 0 0 0 2 7 13 9 1 10 9 1 8 8 9 0 1 9 0 2
73 7 13 8 8 7 9 0 0 14 13 1 9 0 1 9 9 0 2 8 8 0 9 0 1 7 13 9 1 9 9 13 1 9 9 9 0 1 15 1 9 9 0 0 1 9 9 0 1 9 0 2 1 7 13 9 0 0 0 1 9 9 1 9 10 9 2 0 9 1 9 0 2 2
57 7 13 9 9 9 0 1 9 9 0 2 0 1 7 15 1 9 9 1 9 0 1 9 9 10 9 0 1 10 13 1 9 9 12 9 0 1 15 2 0 7 9 9 0 0 13 1 9 9 0 1 10 9 9 12 9 2
61 7 9 1 9 1 9 9 0 1 9 0 1 9 0 2 13 8 8 1 9 1 9 2 0 9 0 1 9 2 7 14 13 9 10 9 9 1 9 9 10 9 1 9 0 1 9 9 0 2 7 13 10 9 1 9 9 1 10 9 2 2
51 7 9 0 13 1 9 0 2 1 10 0 1 9 9 0 1 9 0 1 9 9 9 0 7 9 9 7 9 9 7 9 0 8 0 1 9 9 1 9 9 7 9 0 2 7 9 0 1 9 0 2
50 7 13 7 9 0 1 9 13 1 9 9 1 9 0 14 13 15 9 1 9 9 0 1 9 2 7 1 3 14 13 9 1 10 9 7 14 13 9 0 0 1 9 0 1 9 9 1 15 2 2
27 7 15 9 9 0 9 15 2 1 9 10 9 0 13 9 0 1 9 0 9 14 13 1 9 7 3 2
38 7 13 9 9 0 7 9 15 1 9 9 1 9 9 0 14 13 13 9 9 1 9 9 9 0 1 9 0 2 7 7 13 10 9 0 1 9 2
60 7 13 8 8 9 9 9 0 1 7 15 14 13 1 9 9 1 0 9 9 0 8 1 15 13 15 8 1 9 9 0 1 9 0 13 9 1 9 15 7 9 1 15 7 9 1 9 2 7 9 1 9 1 9 9 7 1 9 0 2
9 8 13 9 12 12 9 1 12 9
20 13 8 9 0 1 9 0 9 9 1 9 7 0 9 0 1 9 0 0 2
44 13 9 0 1 9 9 1 9 1 9 1 9 1 9 0 2 12 2 12 7 2 12 2 12 9 1 15 2 12 2 12 9 9 0 7 12 7 2 12 2 12 9 2 2
77 7 13 9 0 1 9 9 0 7 9 9 15 13 15 8 1 9 1 9 9 7 9 1 9 1 9 12 1 12 13 12 12 9 2 1 15 12 12 1 9 9 7 12 12 9 0 13 9 10 9 1 9 9 9 7 9 9 0 7 9 9 7 9 9 0 7 0 7 9 9 0 7 0 1 9 0 2
41 7 13 9 7 9 9 8 1 9 9 9 1 12 9 12 1 9 1 9 0 13 1 2 12 2 12 9 1 9 9 0 1 9 7 13 2 12 2 12 9 2
76 7 13 9 8 1 9 9 9 1 9 9 0 2 12 2 9 1 2 12 2 12 9 1 9 9 0 0 2 12 2 12 9 7 13 9 7 15 13 1 9 0 9 9 1 9 7 8 13 1 9 15 9 9 0 1 9 9 0 1 9 9 9 0 1 9 0 1 9 9 9 7 9 0 1 9 2
35 7 13 9 1 7 15 8 9 9 0 0 1 9 0 1 9 1 9 0 1 9 0 7 13 1 15 9 0 1 9 8 2 8 2 2
30 7 13 9 1 9 9 1 9 9 1 9 0 1 9 9 1 9 1 1 9 0 15 14 13 1 15 9 9 0 2
8 9 0 1 9 9 9 9 9
26 13 9 1 9 0 1 9 9 7 9 9 7 9 0 1 9 9 9 9 9 9 9 7 9 9 2
21 13 9 7 9 9 9 9 1 9 1 9 9 7 9 7 9 9 1 9 0 2
22 7 13 1 7 9 0 13 9 1 9 15 1 9 0 1 9 9 0 1 9 15 2
28 13 9 0 9 9 0 1 9 9 9 12 1 9 12 13 1 9 9 1 0 15 7 9 0 1 9 15 2
41 7 13 9 9 0 1 9 9 9 9 12 9 1 15 9 12 15 13 9 1 9 9 7 13 1 7 15 13 1 9 9 9 9 0 1 9 0 9 9 0 2
23 7 13 9 9 1 9 0 1 9 0 15 1 15 9 0 7 13 1 0 1 9 0 2
21 13 9 9 7 1 10 9 14 13 9 9 0 1 9 0 7 0 1 9 0 2
19 7 13 7 9 1 9 13 9 0 1 9 9 0 1 9 0 9 12 2
43 7 13 7 9 9 0 13 1 9 9 7 9 7 13 7 13 9 0 15 15 0 7 9 15 14 13 1 15 1 9 7 13 9 1 15 14 13 1 15 1 9 0 2
26 7 7 15 1 9 0 7 13 9 0 7 13 9 1 9 1 9 9 0 15 13 1 15 9 0 2
31 7 13 9 9 7 9 9 9 9 0 15 9 2 9 2 7 14 13 9 15 1 9 1 9 9 15 14 13 9 0 2
40 7 13 1 9 9 9 0 1 9 1 14 9 7 1 9 9 9 0 1 9 9 9 1 9 0 7 9 9 0 1 9 7 9 9 0 7 8 0 9 2
9 9 9 9 13 12 9 1 9 0
37 13 9 9 9 9 1 9 0 7 0 7 9 9 7 9 9 7 9 9 7 13 1 12 9 1 9 1 9 9 0 1 12 5 1 9 0 2
27 7 13 0 9 9 9 0 1 9 9 0 1 9 12 9 9 9 9 9 0 7 9 9 1 9 0 2
67 13 8 8 8 9 9 9 0 1 9 9 12 9 1 9 0 1 9 9 7 9 9 15 1 9 0 9 15 0 9 8 0 7 9 0 1 9 7 13 9 9 15 9 12 2 12 0 13 15 9 8 9 9 9 0 1 9 0 7 9 9 0 0 1 9 9 2
50 7 13 9 8 8 9 9 9 15 13 9 0 14 7 15 13 1 9 9 0 1 10 9 7 13 9 0 1 9 0 1 9 9 7 13 1 9 9 9 8 0 1 9 1 9 15 1 9 9 2
39 14 9 0 0 1 9 7 15 9 9 7 0 1 9 7 13 9 12 9 0 1 9 9 7 9 9 7 7 12 8 8 8 7 0 13 1 9 0 2
40 7 13 7 9 0 1 12 9 1 9 1 9 7 13 9 9 9 1 9 9 1 9 9 8 0 1 9 9 1 9 1 9 1 9 9 7 9 1 9 2
36 7 12 9 9 1 9 9 13 9 9 1 9 9 12 2 12 0 9 15 7 13 9 9 15 12 9 9 0 7 13 0 9 1 12 9 2
34 13 9 7 9 9 1 9 9 0 1 15 13 1 9 9 9 9 9 7 13 9 9 0 1 9 0 1 9 7 13 1 9 9 2
44 7 13 9 7 9 15 13 15 9 9 1 9 9 7 15 13 1 9 8 0 1 9 9 9 13 9 0 1 9 9 9 9 1 7 15 13 1 9 9 0 1 9 9 2
39 7 13 1 9 9 1 9 9 9 0 1 9 1 9 0 7 13 9 9 9 7 1 0 13 9 9 1 9 0 7 9 9 9 14 13 12 9 3 2
9 9 9 9 9 0 13 9 9 9
110 13 9 9 9 9 0 1 9 0 1 9 14 13 9 9 1 9 0 2 7 14 13 9 9 1 12 9 2 12 9 2 1 9 13 12 9 2 1 12 9 2 1 9 12 0 9 15 13 9 9 0 1 9 9 0 0 1 9 1 9 9 9 9 2 7 9 9 9 1 9 9 0 1 9 1 9 9 9 2 7 3 9 15 13 15 9 1 9 9 0 1 9 2 9 1 9 10 9 1 9 9 0 2 7 9 9 1 9 0 2
38 7 13 9 7 9 14 13 9 9 9 9 0 7 9 9 9 1 9 10 9 1 1 9 9 9 0 1 9 9 9 13 9 9 7 13 9 9 2
46 7 13 9 9 9 9 0 1 9 9 1 9 9 2 7 3 9 9 1 9 9 7 9 9 9 15 13 9 1 15 1 9 9 7 9 9 7 9 0 9 1 9 9 7 9 2
38 7 13 9 1 7 9 9 9 1 9 9 14 13 0 8 1 9 9 0 1 9 9 1 9 9 0 7 9 15 1 1 12 9 1 0 1 9 2
90 9 15 13 15 9 0 0 1 9 13 7 9 9 9 9 0 1 9 9 1 9 0 7 15 13 1 9 0 0 1 12 9 1 12 9 3 9 12 2 7 7 9 9 9 1 10 9 1 9 1 9 9 1 9 9 2 13 1 9 9 9 0 1 9 9 0 7 0 9 15 13 0 7 1 9 1 9 1 9 9 0 13 1 9 9 1 10 9 0 2
31 7 13 9 7 9 9 9 8 0 13 1 9 9 7 9 1 9 9 1 9 9 9 0 1 9 9 0 1 9 9 2
31 7 13 9 7 3 9 13 1 9 9 1 15 9 9 9 1 9 9 0 1 9 1 9 9 1 9 9 1 9 9 2
27 7 13 9 0 9 0 1 9 9 15 13 1 0 9 7 0 1 9 9 1 9 9 1 9 1 9 2
100 7 1 15 13 9 9 9 2 9 9 9 2 7 14 9 0 1 9 13 0 1 9 1 9 0 9 0 1 9 7 9 9 9 1 9 1 9 9 0 15 1 7 9 1 9 1 9 0 1 9 1 9 12 9 0 1 9 0 13 9 9 0 7 13 1 12 9 1 0 1 12 9 1 9 0 2 7 15 1 9 9 9 9 1 9 1 9 15 1 9 9 15 13 0 1 9 9 9 2 2
28 7 13 9 1 9 1 7 15 9 1 9 1 9 0 7 9 9 14 13 7 7 9 13 1 9 9 15 2
91 7 1 9 0 14 13 9 9 0 1 9 9 7 15 13 15 1 9 9 0 1 9 9 15 2 7 13 9 8 8 9 9 9 2 9 11 0 1 9 2 7 9 9 9 13 9 0 7 13 9 7 13 7 1 15 9 15 0 1 9 9 7 1 15 9 9 0 8 0 1 0 1 12 9 0 1 7 9 9 9 1 9 0 1 0 1 1 12 9 3 2
46 7 13 8 1 7 9 13 9 9 9 7 9 0 1 9 9 7 9 9 0 0 1 9 9 1 9 15 1 9 9 7 13 1 9 9 9 9 0 1 8 7 9 9 0 0 2
24 9 1 9 9 0 1 9 0 7 0 7 9 1 9 0 1 9 9 9 1 9 9 9 2
56 7 13 8 7 9 0 14 13 0 1 9 9 7 9 9 15 1 9 2 7 14 13 9 9 9 9 0 2 0 7 9 1 10 9 15 13 1 9 0 1 15 13 1 12 5 7 12 5 1 9 0 0 13 12 5 2
9 9 0 1 9 9 9 9 1 9
52 13 8 8 9 0 1 9 0 1 9 8 8 8 7 15 7 1 0 9 1 9 0 13 9 0 9 0 1 9 1 9 0 9 1 9 15 1 9 0 1 9 9 9 9 1 9 13 1 12 12 9 2
35 7 13 8 7 9 15 7 15 9 0 1 10 9 2 15 13 9 9 1 9 15 0 2 13 1 9 9 0 1 9 7 9 1 15 2
32 7 13 8 7 9 0 14 13 1 9 0 1 0 7 9 0 1 9 7 14 13 1 9 9 9 9 0 7 0 7 0 2
28 7 13 8 7 9 14 13 1 12 5 1 9 15 1 9 7 9 0 7 1 0 7 13 0 1 12 9 2
37 7 13 7 9 14 13 1 9 0 1 9 0 7 12 5 1 9 9 14 13 1 9 1 8 7 9 0 7 1 9 9 1 9 9 9 0 2
12 9 9 0 1 9 12 12 9 1 12 9 2
32 13 9 0 1 9 9 0 1 9 9 7 9 9 1 9 9 9 15 12 12 9 1 14 2 12 2 9 0 1 9 0 2
33 13 9 7 9 15 13 9 15 13 9 0 9 1 9 15 13 9 15 1 9 9 1 9 12 7 13 9 9 1 12 12 9 2
36 7 13 9 7 9 0 7 9 0 13 9 0 1 9 9 1 8 7 13 9 9 1 10 9 12 12 9 7 13 9 12 1 12 12 9 2
44 7 13 9 7 9 9 0 1 8 13 1 9 1 9 1 9 1 9 0 1 12 12 9 1 12 12 9 1 9 9 1 9 12 1 9 9 15 12 12 13 9 12 5 2
7 9 9 7 9 13 12 9
23 13 9 1 9 15 1 0 9 0 1 9 1 9 9 0 1 9 8 7 9 7 8 2
37 7 14 13 9 9 0 1 9 7 9 1 9 0 9 12 9 0 1 9 9 0 12 7 12 12 9 1 9 9 15 12 5 9 1 9 0 2
39 7 14 13 9 9 0 1 9 1 12 12 9 9 0 1 12 12 9 1 9 12 1 1 13 8 8 1 9 1 12 12 9 1 9 9 15 12 5 2
113 7 13 9 0 1 7 9 9 0 13 1 9 15 13 15 9 0 1 9 0 7 0 15 9 9 7 9 15 13 9 15 1 12 12 9 1 9 0 1 1 12 12 9 1 9 12 7 9 7 9 1 9 7 9 0 15 13 9 15 1 12 12 9 1 9 0 1 12 12 9 1 9 12 7 13 9 15 1 9 7 9 1 12 12 9 1 1 12 12 9 7 13 9 9 15 1 9 7 9 15 1 1 12 12 9 1 1 12 9 1 9 12 2
32 1 9 9 9 0 1 9 0 8 8 9 7 9 9 15 1 9 1 12 12 9 7 9 7 9 8 1 9 12 9 9 2
11 9 0 2 0 1 9 9 9 1 9 0
49 13 9 9 0 0 1 9 9 9 9 9 1 9 0 0 13 1 9 9 9 0 1 9 0 13 9 0 9 1 15 1 9 7 13 9 15 0 7 1 9 15 13 1 15 9 1 10 9 2
66 7 13 9 8 9 8 9 9 2 8 2 1 9 9 2 7 9 0 15 13 9 1 15 2 9 8 2 13 14 13 0 9 0 0 1 9 9 15 2 8 8 2 1 9 1 9 12 12 9 7 13 8 8 9 0 1 9 9 7 9 7 9 1 9 0 2
43 7 13 1 7 10 9 13 0 1 9 1 9 0 1 1 15 9 0 1 9 7 9 9 7 9 7 9 1 9 9 9 1 9 0 7 9 0 7 9 7 9 15 2
15 9 1 0 9 9 7 9 7 9 1 9 9 1 9 8
79 13 9 9 8 8 9 9 0 9 8 1 9 0 1 9 9 0 1 9 9 1 9 0 1 9 7 9 9 9 0 7 15 13 1 15 1 9 9 1 9 1 9 1 0 1 9 7 1 9 0 13 9 9 8 8 9 9 0 9 15 1 0 9 1 9 1 9 9 1 9 0 1 9 0 1 9 9 0 2
91 7 13 8 2 8 8 9 9 9 0 1 9 0 7 8 2 8 13 1 7 9 9 1 9 9 8 1 9 0 14 13 1 12 9 13 1 9 15 9 1 8 9 9 1 9 8 8 8 15 1 9 7 9 0 7 0 1 9 9 9 0 0 9 15 1 9 7 9 1 9 9 9 0 1 0 9 0 1 9 7 9 1 9 8 1 9 15 1 9 9 2
79 7 0 9 9 1 0 12 9 1 9 1 9 8 1 9 9 0 9 1 9 7 9 15 13 15 9 9 7 13 9 9 0 1 10 9 1 9 9 15 1 9 9 7 9 7 9 0 7 13 10 9 9 9 9 1 9 9 15 1 9 0 1 1 9 0 13 1 9 15 9 1 9 9 15 13 15 9 9 2
76 7 13 9 0 1 9 1 9 0 1 9 9 15 0 7 0 0 1 9 9 0 9 1 8 7 8 7 8 8 1 9 0 7 1 15 13 1 9 0 9 1 9 9 1 9 0 1 10 9 1 9 9 0 1 9 7 9 9 0 1 15 1 1 9 9 0 1 9 0 1 10 9 1 9 0 2
50 7 14 13 10 9 1 9 1 9 1 9 9 9 0 7 9 0 15 14 13 1 15 9 7 14 13 1 9 0 9 0 1 9 7 9 0 1 9 1 9 1 10 9 1 9 1 9 15 0 2
97 7 9 0 9 1 9 0 7 0 7 9 9 0 1 1 9 9 7 9 9 1 15 1 9 9 0 2 7 13 9 1 9 9 0 7 9 9 0 1 8 1 9 1 9 1 9 9 0 1 15 1 15 1 9 9 7 9 1 9 7 9 7 9 9 15 13 15 9 8 7 7 9 9 7 9 9 9 9 7 13 1 9 0 1 9 9 9 9 8 0 10 9 0 1 9 9 2
54 7 0 14 13 9 9 9 7 9 0 1 9 9 1 9 15 7 9 15 7 13 10 9 2 9 0 13 1 9 9 0 7 9 9 9 7 9 7 9 9 7 9 9 1 9 0 7 0 1 9 9 7 9 2
12 0 1 12 9 9 0 1 9 9 0 1 9
51 13 9 0 1 9 9 9 0 1 9 0 15 13 1 9 9 0 1 9 1 0 9 0 2 1 1 12 12 9 0 2 12 12 9 2 0 1 0 2 7 8 0 1 15 14 13 12 12 9 3 2
90 7 13 9 15 13 15 1 9 9 9 9 7 9 0 1 9 0 2 7 9 9 0 1 9 0 13 15 1 12 1 12 12 9 0 2 7 7 9 9 0 7 15 13 1 9 9 0 13 1 12 12 9 2 12 12 9 2 7 15 15 13 15 9 8 8 8 9 9 9 0 15 13 9 15 1 9 0 2 13 7 9 10 9 13 1 9 9 1 9 2
41 7 13 9 7 1 12 12 9 0 1 1 12 12 9 3 2 15 15 13 9 9 1 9 15 1 9 0 2 7 1 15 9 1 9 9 2 7 9 9 3 2
32 7 14 13 3 9 0 1 9 9 15 0 7 7 13 13 9 1 9 7 13 9 15 1 10 9 1 9 9 0 1 9 2
22 7 13 1 7 10 9 13 1 12 12 9 2 7 13 1 1 12 12 9 7 9 2
48 7 13 9 7 0 1 12 5 1 9 13 1 9 9 0 7 0 1 0 0 2 7 15 9 15 13 9 0 1 9 7 1 9 0 0 7 15 13 9 1 9 0 1 9 10 9 9 2
88 7 13 9 9 9 9 0 1 9 0 2 7 13 9 1 9 1 8 9 1 10 9 1 9 8 1 0 8 2 0 7 15 9 0 7 13 9 9 0 2 7 13 9 8 0 15 1 12 7 13 1 12 12 9 0 2 7 13 9 0 1 9 0 7 13 9 0 0 1 9 0 1 9 9 0 1 15 14 13 1 9 1 9 1 9 9 0 2
9 12 9 7 12 9 9 1 9 0
39 13 9 9 1 9 15 9 0 9 9 9 12 9 1 9 9 0 7 9 9 9 7 9 7 9 1 9 1 9 1 12 9 9 1 9 9 9 9 2
41 13 9 8 8 9 0 1 9 9 15 13 1 15 7 13 1 12 9 1 9 9 7 9 9 7 9 7 9 0 7 9 7 9 7 9 7 9 7 9 0 2
63 13 9 9 1 9 9 1 9 9 9 7 9 9 9 7 13 1 9 9 7 9 7 9 2 7 9 9 7 9 9 9 1 9 9 9 0 1 9 0 7 9 9 12 9 1 9 7 9 1 9 0 7 9 9 0 7 13 1 9 9 9 9 2
32 7 13 9 0 1 9 9 0 7 9 1 9 9 1 9 9 1 9 0 1 9 7 13 1 9 9 9 7 9 8 8 2
52 7 13 9 0 1 9 9 1 9 9 0 15 13 9 15 12 12 9 7 15 13 9 1 9 12 7 15 13 1 9 9 9 0 0 7 9 9 9 0 1 9 2 8 8 2 1 9 7 9 10 9 2
70 7 13 9 8 8 9 1 9 9 1 9 9 9 9 9 7 9 0 0 1 9 1 9 7 9 9 1 9 9 0 0 1 9 1 9 9 9 0 1 9 0 7 9 9 9 9 0 1 9 0 1 9 0 7 9 9 9 1 9 10 9 1 9 9 0 1 15 1 9 2
21 7 13 9 9 9 9 1 9 9 0 7 9 10 9 0 1 9 9 7 9 2
40 7 13 1 9 0 1 9 9 0 7 9 7 9 9 13 1 9 0 1 9 9 7 9 10 1 9 9 1 9 9 1 9 9 9 9 1 1 10 9 2
35 7 13 9 0 0 1 8 2 8 8 7 9 8 8 8 9 9 9 9 9 0 1 9 7 9 9 2 7 9 9 9 1 9 15 2
39 7 13 9 2 8 8 2 1 9 1 9 9 1 9 9 1 9 0 7 9 0 1 9 9 0 0 0 7 1 9 0 1 9 9 1 9 9 0 2
36 7 13 9 12 9 9 1 9 9 9 9 1 1 9 2 7 9 9 0 1 9 9 9 1 9 9 7 9 9 9 1 9 9 1 9 2
11 9 0 1 9 9 1 9 1 9 9 0
113 13 9 12 2 12 0 8 0 0 1 9 9 9 0 8 8 2 7 1 9 15 13 1 15 9 9 0 8 8 8 7 2 9 7 9 13 9 8 8 0 0 2 2 7 7 8 14 13 1 9 0 0 2 13 9 9 0 8 8 7 9 14 13 9 1 1 9 9 1 9 7 0 1 0 1 12 9 2 9 7 8 13 1 9 9 1 9 9 9 9 12 2 12 0 9 9 8 8 9 9 1 9 9 9 7 9 15 1 9 2 9 2 2
77 7 1 7 13 9 0 9 12 2 12 0 0 7 9 13 1 9 9 0 1 9 13 8 7 9 7 9 13 9 9 8 8 7 7 9 0 1 10 9 14 13 9 15 1 9 0 2 7 13 8 1 2 9 0 0 2 2 0 2 8 7 9 1 9 7 9 14 13 8 1 9 0 7 9 0 2 2
36 7 9 0 13 9 1 9 0 1 9 9 0 7 14 13 9 9 0 8 8 7 15 2 14 13 1 9 9 1 9 2 9 0 1 9 2
13 7 13 1 9 9 7 9 9 9 0 1 9 2
23 7 13 9 0 7 0 7 9 9 8 13 9 1 9 0 1 9 0 8 8 1 9 2
42 7 13 9 0 1 7 2 9 7 9 0 1 9 1 0 1 9 7 13 1 9 0 9 1 9 9 0 8 8 7 0 8 8 1 8 1 0 1 9 0 2 2
19 12 12 0 1 9 0 13 1 9 7 13 9 2 8 2 1 9 1 8
58 13 1 9 1 12 12 0 1 9 8 7 0 15 7 15 13 9 0 9 7 9 7 0 1 9 9 9 2 1 9 9 0 0 1 15 2 13 1 12 12 13 1 9 8 2 12 8 9 9 8 8 2 1 9 9 0 0 2
29 7 13 10 9 1 9 0 1 9 7 13 1 15 9 0 1 9 2 9 0 1 0 0 1 8 1 9 2 2
34 7 14 13 10 9 2 0 2 1 9 2 9 15 13 9 1 9 15 13 1 9 7 13 9 1 9 0 0 2 9 8 7 8 2
94 7 1 9 10 9 2 8 8 2 7 14 9 0 13 9 1 9 9 2 9 2 1 12 9 1 9 2 12 2 2 7 7 15 13 15 1 9 0 7 1 9 9 0 2 1 9 9 2 7 13 0 0 0 9 0 1 9 7 13 13 0 2 7 1 9 9 7 9 1 9 12 2 7 13 9 0 1 9 15 0 1 9 0 1 9 0 9 7 9 8 1 9 0 2
21 14 13 1 10 9 0 9 1 9 0 7 14 13 1 15 9 14 1 15 13 2
53 7 9 0 15 13 9 15 1 9 0 2 13 1 12 9 7 13 10 9 1 8 7 13 9 2 8 2 1 9 1 9 2 7 13 9 7 9 13 13 15 1 10 9 7 14 13 13 1 15 9 9 15 2
42 7 9 15 15 8 8 2 7 15 9 9 0 7 0 2 13 8 1 9 2 7 9 0 13 1 9 7 13 9 0 2 0 9 7 0 9 0 2 1 15 2 2
29 7 13 2 7 9 0 9 1 10 13 7 15 13 0 9 7 13 2 14 15 9 8 2 9 9 0 1 9 2
42 1 15 9 0 0 1 9 7 9 8 8 8 8 7 13 2 7 15 13 9 0 1 9 2 7 15 13 9 15 7 9 15 1 9 7 13 9 9 1 9 2 2
28 7 13 8 9 0 1 9 1 9 1 0 9 7 9 2 8 8 7 15 9 15 13 9 0 1 9 0 2
34 8 7 13 9 1 9 0 2 0 7 13 9 0 13 1 8 1 9 9 12 9 1 9 9 0 1 9 7 12 9 1 9 15 2
48 7 1 9 8 8 2 7 14 9 13 9 7 14 13 9 8 1 9 10 9 1 9 9 8 2 8 8 2 7 15 1 9 8 7 13 0 9 0 1 9 1 7 9 15 3 15 9 2
11 9 13 9 0 1 9 9 9 15 1 8
38 13 9 9 0 1 9 15 13 1 15 9 9 15 8 8 1 8 7 13 15 9 1 9 0 15 14 13 9 9 0 0 1 9 15 1 12 9 2
51 7 1 9 9 8 8 8 9 13 1 9 9 1 9 9 8 1 9 1 9 0 8 1 9 2 7 13 9 15 1 1 12 12 2 13 9 0 1 9 7 8 13 1 9 0 9 9 1 9 0 2
34 7 9 1 9 9 9 15 1 9 7 14 8 13 9 12 9 13 9 9 0 1 9 0 9 9 9 0 1 9 9 0 1 8 2
32 7 13 9 1 9 9 9 0 1 8 7 1 9 9 9 0 9 9 0 0 7 15 14 13 9 0 1 9 0 2 0 2
43 7 13 1 2 9 0 0 2 1 9 8 15 13 15 9 13 9 9 13 9 1 9 9 7 9 7 9 1 9 9 9 0 0 1 9 0 1 9 9 0 1 8 2
13 0 1 8 13 8 1 9 1 9 9 15 1 8
69 13 9 2 8 2 7 9 1 2 9 0 8 1 9 0 2 13 1 9 8 0 0 1 9 0 8 8 1 9 9 15 1 9 15 15 13 15 1 8 1 9 15 7 9 15 1 9 15 2 0 7 9 10 9 15 13 9 15 1 12 12 9 13 1 15 8 9 15 2
55 7 13 7 9 1 9 0 14 13 10 9 1 9 0 13 1 8 0 1 9 9 12 9 1 9 9 0 1 9 0 8 2 7 12 9 1 9 0 1 8 1 9 2 7 14 13 9 1 15 1 9 0 1 8 2
32 7 13 8 7 15 1 9 9 1 9 1 9 9 1 8 13 9 9 1 8 1 9 0 0 1 9 15 13 15 1 8 2
13 7 13 8 1 9 1 9 0 1 9 8 8 2
19 9 1 9 0 0 2 8 13 9 15 1 9 1 9 9 7 9 9 15
69 13 9 0 0 8 8 1 9 15 1 9 8 9 9 15 1 9 1 9 9 0 2 7 13 9 9 15 0 1 9 7 9 9 15 15 8 1 15 9 9 15 9 8 7 13 7 9 9 9 15 9 1 9 0 1 9 8 8 0 2 9 1 9 1 9 0 8 8 2
87 13 1 15 9 0 1 9 0 0 15 13 15 9 8 8 2 7 13 2 8 13 9 8 8 1 9 8 15 13 12 1 8 9 9 1 9 9 9 0 0 7 13 8 1 15 9 7 15 13 2 9 15 2 1 9 9 0 8 2 2 0 1 7 9 13 1 9 1 9 8 8 1 9 8 2 7 15 9 15 13 8 1 15 1 9 15 2
76 7 13 9 0 15 13 9 9 9 15 1 9 1 2 9 0 2 1 9 9 12 2 12 0 1 7 9 0 1 15 13 7 9 0 0 13 1 12 12 9 0 1 9 9 0 1 9 9 0 2 7 7 10 9 13 15 1 9 0 1 9 7 13 1 15 1 9 1 9 9 9 0 7 9 0 2
82 7 13 9 2 7 8 8 13 1 9 9 15 15 13 1 15 9 0 1 9 15 7 14 13 1 9 15 9 1 9 15 1 7 15 9 7 7 15 14 13 9 7 13 15 1 15 7 3 1 9 1 0 15 2 2 0 2 7 1 9 0 1 15 7 8 8 13 0 9 1 9 15 7 7 15 13 1 15 1 9 0 2
45 7 14 13 9 15 7 13 9 0 0 13 9 9 7 9 15 0 7 15 13 1 7 15 1 0 2 13 9 9 9 9 9 0 9 9 0 13 15 9 9 0 1 9 0 2
104 7 13 9 0 1 9 0 0 7 9 9 9 0 0 13 1 9 9 1 9 0 1 9 8 8 0 7 13 9 1 9 0 1 9 0 2 0 1 7 9 10 13 15 9 0 1 9 13 1 9 15 1 9 7 9 1 9 0 13 9 1 9 9 15 15 13 13 1 15 9 9 0 7 7 15 13 13 1 1 11 8 8 8 8 8 8 8 8 7 9 15 1 9 7 13 1 9 1 15 7 9 1 15 2
47 7 13 7 9 9 13 9 1 9 7 9 15 13 1 9 9 8 8 0 7 11 13 1 9 9 2 7 7 10 9 13 1 9 9 9 9 7 13 9 15 1 9 0 1 9 9 2
57 1 9 0 13 8 8 8 9 9 8 8 7 15 14 13 1 9 9 9 1 9 0 0 1 7 13 9 0 1 9 8 8 8 8 1 9 7 9 9 0 7 0 1 9 9 15 9 1 9 0 1 0 12 1 9 0 2
10 9 8 8 1 9 0 1 12 12 9
28 13 9 0 1 9 9 0 1 9 0 1 9 0 1 12 12 9 1 12 12 9 1 9 9 1 9 0 2
32 7 13 9 0 13 1 9 0 0 7 9 8 8 1 9 0 13 9 7 13 1 9 9 15 9 0 1 9 9 9 0 2
97 7 13 9 7 8 8 1 9 9 0 1 9 9 15 13 1 12 12 9 1 12 12 9 2 7 9 0 0 1 12 12 9 1 12 12 9 2 8 0 7 9 8 0 1 12 12 9 1 12 12 9 2 9 0 0 1 12 12 9 1 12 12 9 2 9 0 1 12 12 9 1 12 12 9 2 9 0 1 12 12 9 1 12 12 9 2 7 8 1 12 12 9 1 12 12 9 2
8 12 12 9 1 9 12 9 0
36 1 0 7 13 9 9 0 15 13 15 9 0 1 9 0 1 12 9 8 8 0 12 12 7 12 12 9 1 9 1 9 15 13 15 9 2
38 13 9 8 8 9 9 0 1 9 2 7 10 9 13 12 9 1 9 0 7 12 9 1 9 8 7 12 9 1 9 8 7 12 9 1 9 9 2
38 0 7 9 9 8 1 10 9 13 12 12 7 12 9 8 8 0 12 12 9 7 7 9 9 1 9 12 12 7 12 9 8 8 0 12 12 9 2
55 13 1 7 9 9 0 13 1 9 0 1 9 15 9 0 13 1 15 9 9 0 2 0 7 9 0 13 9 0 13 1 15 9 9 9 7 13 9 1 9 7 9 0 1 9 7 9 0 7 0 7 9 7 9 2
85 7 13 7 9 13 1 9 12 8 0 1 9 8 1 9 12 9 7 15 13 0 8 1 9 1 9 0 2 7 1 8 9 1 9 0 7 9 8 8 8 9 7 1 15 13 9 8 1 12 8 8 8 0 12 12 9 2 0 1 7 9 13 9 0 13 12 12 9 1 9 0 1 9 9 9 1 9 7 13 9 9 1 9 0 2
10 12 9 9 0 1 9 9 1 14 9
56 13 9 12 2 12 0 0 9 9 1 9 9 1 9 8 8 12 9 1 9 7 13 9 9 1 12 1 12 9 7 13 10 9 9 1 9 9 0 1 9 9 1 9 0 1 9 9 9 0 7 9 9 1 9 0 2
21 7 13 9 9 9 14 13 3 1 1 9 9 0 7 13 1 12 9 1 9 2
51 13 7 9 9 0 1 9 9 7 9 9 14 13 1 9 1 9 9 9 1 9 9 0 1 9 9 7 9 1 15 13 1 9 12 9 15 13 1 15 1 9 9 7 9 7 9 9 7 9 15 2
49 7 13 9 9 9 0 1 9 9 7 9 7 0 1 9 9 1 9 9 1 9 1 12 5 1 12 5 1 9 9 9 9 0 7 13 9 1 9 9 9 0 1 9 9 7 9 1 9 2
4 9 9 13 0
48 13 9 8 8 1 9 9 9 9 0 1 9 2 8 2 8 2 1 1 12 9 10 9 1 9 8 13 9 9 13 9 9 1 9 0 2 7 9 1 9 13 1 1 12 9 1 9 2
63 7 13 7 9 8 8 13 1 9 1 9 8 9 9 9 1 9 1 15 1 9 9 9 9 1 9 9 1 9 9 0 9 15 13 0 1 1 12 9 1 9 1 12 9 1 9 1 9 2 9 1 9 9 9 8 9 7 9 15 1 9 0 2
70 7 7 9 0 1 9 9 13 1 9 0 9 9 10 2 7 7 9 9 14 13 0 9 1 9 8 8 1 9 9 9 9 9 2 7 7 8 8 13 9 9 9 1 9 8 8 9 1 9 15 7 9 0 2 7 1 3 14 13 1 0 9 0 7 13 1 9 9 9 2
58 7 13 9 9 9 14 13 1 9 9 8 1 9 9 1 9 1 9 9 2 7 15 0 0 2 9 1 7 15 14 13 9 9 1 9 1 9 7 9 1 15 0 1 9 1 9 0 9 2 1 7 13 9 15 1 15 1 2
60 1 9 0 2 13 9 9 8 9 9 8 8 1 9 1 9 9 9 0 9 2 8 2 10 9 1 1 12 9 1 9 2 7 13 9 9 9 1 1 12 9 0 9 9 7 9 7 9 7 9 7 9 9 1 9 12 9 1 9 2
52 7 9 9 13 7 9 9 14 13 1 10 9 9 1 15 1 15 1 9 0 1 0 9 1 9 13 1 9 0 0 2 7 1 7 7 14 9 9 13 1 12 1 9 2 13 1 1 12 9 1 9 2
44 7 13 9 9 8 7 13 9 1 9 1 10 9 1 9 9 9 1 9 9 0 1 0 9 2 7 13 1 9 0 1 9 1 9 1 9 12 9 7 15 13 9 0 2
95 7 1 9 10 9 14 13 9 0 13 9 9 8 8 9 9 0 1 9 9 9 9 1 9 0 1 8 7 8 8 8 8 2 7 13 1 9 10 1 9 0 2 7 1 9 13 9 0 0 9 1 9 10 9 2 1 9 9 9 9 2 7 13 9 15 1 9 1 9 9 9 2 7 1 0 7 13 9 1 9 15 2 9 1 9 9 9 9 1 9 0 1 9 0 2
59 7 13 9 0 7 13 8 1 9 9 9 0 1 9 9 10 9 1 9 0 2 0 15 13 1 9 9 15 7 1 15 8 0 1 9 2 7 13 9 7 8 14 13 9 0 0 1 9 9 9 1 9 0 15 13 8 0 0 2
7 9 9 0 1 9 0 9
24 13 9 9 9 0 10 9 9 9 0 1 9 9 1 9 12 8 1 9 12 9 1 9 2
23 13 9 1 9 0 1 9 7 15 9 1 9 9 0 9 0 15 13 9 10 9 0 2
27 7 13 9 0 1 9 9 7 9 0 13 9 0 0 0 7 9 9 15 13 1 10 9 1 9 0 2
98 7 13 7 9 10 9 14 13 1 9 0 1 9 0 1 9 7 15 12 8 1 9 12 9 1 9 1 9 0 15 14 13 15 9 0 1 10 9 12 8 8 13 15 1 12 5 1 9 7 12 8 8 8 13 15 9 0 7 9 9 8 8 1 9 0 1 12 12 9 9 1 9 1 9 0 7 14 9 1 9 12 8 13 7 1 15 7 14 15 14 13 0 7 14 13 9 15 2
11 14 9 1 9 9 12 7 12 7 12 8
86 13 9 0 1 9 0 0 1 9 7 15 14 9 1 9 9 12 8 15 13 1 9 12 9 1 9 2 7 9 12 8 1 9 12 9 1 9 2 7 9 12 8 1 9 12 9 1 9 2 8 8 1 7 13 9 9 9 0 9 12 2 12 0 1 9 9 0 1 9 12 8 1 9 12 9 1 9 0 1 9 1 9 9 9 0 2
7 9 0 1 9 9 9 9
20 13 9 0 9 9 0 1 9 9 9 9 1 9 0 0 1 9 9 9 2
82 7 13 9 8 8 9 9 9 7 9 13 1 9 9 9 9 7 13 15 9 2 8 8 1 9 9 2 7 15 9 9 0 2 0 1 7 9 9 1 0 0 1 9 2 14 7 15 14 13 1 9 15 14 13 9 1 15 2 7 14 13 1 9 12 9 0 7 1 9 0 13 12 7 9 12 9 7 9 15 12 9 2
28 7 13 7 9 14 13 15 1 12 1 12 9 9 0 1 9 7 13 15 1 12 1 12 9 9 1 9 2
17 7 13 7 15 1 0 7 13 9 9 1 9 0 1 9 0 2
7 9 1 9 8 1 9 9
63 13 9 0 9 1 9 9 0 1 9 8 8 9 9 9 0 1 9 8 1 9 9 1 9 1 9 1 9 9 1 9 15 9 9 9 9 7 9 9 1 9 10 1 9 9 8 8 7 9 1 9 9 0 1 9 9 9 1 9 7 9 0 2
38 7 14 13 9 9 1 9 0 1 9 7 9 0 1 9 1 9 0 1 9 9 1 9 0 0 1 9 8 1 9 9 9 0 7 9 15 0 2
83 7 1 0 9 1 9 9 1 9 1 9 8 1 9 12 9 1 9 1 9 9 9 7 9 0 0 1 9 9 1 9 7 9 1 9 0 1 10 13 9 0 1 9 9 9 1 9 7 1 9 2 7 7 9 9 9 9 0 0 1 9 0 1 9 15 13 1 9 1 9 0 1 9 9 0 1 9 9 9 9 1 9 2
8 9 0 1 9 9 9 1 8
33 13 9 8 8 9 9 0 0 1 9 9 0 9 9 1 9 9 0 1 9 9 1 9 8 1 9 1 12 1 12 9 8 2
59 7 13 8 1 7 9 14 13 9 0 1 9 9 1 9 8 9 1 9 7 13 1 9 15 9 15 13 15 9 9 0 0 1 2 9 0 0 1 9 9 1 8 2 7 15 13 1 9 0 1 9 0 1 9 9 7 9 15 2
33 7 13 9 15 13 1 9 9 9 9 1 9 9 13 1 9 0 7 0 7 0 1 9 9 9 9 0 1 9 1 9 0 2
65 7 13 8 8 0 9 9 7 9 9 0 1 9 9 7 9 9 0 15 13 0 1 12 9 1 9 9 13 9 0 1 9 7 9 7 9 9 9 0 7 0 1 9 9 9 9 9 7 9 15 0 1 9 0 9 0 7 1 9 9 0 1 9 0 2
47 7 13 7 9 14 13 9 9 1 9 0 7 9 9 9 0 1 9 1 9 1 9 7 9 0 1 9 9 9 9 1 8 15 13 9 1 9 15 9 12 1 9 9 0 1 9 2
13 9 2 9 0 1 9 0 7 13 1 9 9 15
103 13 9 0 7 9 0 0 1 9 14 13 1 9 9 15 13 1 9 15 7 14 13 9 9 0 1 9 9 7 13 9 1 9 9 7 13 9 0 1 9 15 1 9 0 7 14 13 9 9 0 1 9 9 0 7 0 2 0 1 7 15 1 9 9 0 1 9 1 10 9 1 10 13 1 15 1 9 14 7 9 9 9 1 10 9 1 9 0 13 0 9 1 7 9 10 9 1 9 13 0 1 9 2
35 7 13 9 0 9 1 9 0 15 1 9 0 9 1 9 9 1 9 0 7 0 2 9 15 13 1 9 10 9 1 9 1 9 0 2
81 7 13 9 0 1 9 1 9 1 9 9 1 9 9 7 9 15 1 9 7 9 9 0 2 1 9 1 7 9 0 0 9 0 7 13 9 9 0 7 0 1 9 9 0 1 9 12 9 2 7 13 1 9 9 9 0 1 9 0 1 9 7 9 9 1 9 13 9 0 13 9 15 9 12 2 12 1 9 12 5 2
98 7 13 9 1 7 15 1 9 1 9 15 13 1 9 9 9 0 14 7 9 0 1 10 9 14 13 9 0 7 13 9 0 2 0 7 0 1 9 10 9 13 9 9 15 1 9 0 9 1 9 7 9 9 1 9 7 1 9 9 0 1 9 0 7 1 9 9 1 9 1 15 1 9 0 2 7 15 9 15 14 13 1 9 9 0 7 13 15 1 0 9 9 0 1 9 9 0 2
73 7 1 9 9 2 13 9 9 9 9 0 7 0 1 9 0 1 9 7 13 1 12 5 1 9 2 7 12 5 1 9 12 1 12 5 1 9 2 7 12 5 1 9 9 12 1 1 13 9 9 0 1 9 0 1 10 9 1 12 5 1 9 12 7 13 1 12 5 1 9 9 12 2
44 7 13 9 9 9 9 0 7 0 1 9 9 10 9 1 9 1 9 0 9 7 0 1 9 0 9 9 9 9 0 1 9 9 7 9 9 9 1 15 1 9 9 0 2
66 7 13 9 7 15 1 9 9 9 9 0 1 9 0 7 13 9 15 1 1 12 5 1 12 5 1 9 9 12 8 7 9 10 9 13 0 1 9 1 9 9 1 9 0 7 13 9 9 0 1 9 0 1 8 0 7 8 1 12 5 7 12 5 1 9 2
90 7 13 9 1 9 9 9 15 13 1 9 9 0 7 9 9 15 1 9 0 7 0 7 15 9 10 13 1 9 9 0 2 0 1 7 1 1 12 9 0 13 12 9 1 9 12 5 13 1 9 9 0 15 13 1 9 0 1 9 0 1 12 9 1 9 9 2 12 9 1 9 7 9 2 12 9 1 9 9 2 7 15 9 14 13 1 9 0 0 2
99 7 13 9 7 9 0 13 9 9 15 13 9 1 15 1 9 9 9 1 15 13 15 1 9 0 1 9 9 1 9 15 13 1 9 9 0 2 7 1 15 7 14 9 9 9 1 9 9 0 0 13 9 9 9 15 13 15 9 1 12 12 9 1 9 9 12 1 12 12 9 1 9 9 12 7 15 9 15 13 1 9 9 0 1 10 9 1 12 9 9 12 1 12 9 1 9 9 12 2
8 9 0 9 0 1 8 1 8
86 13 9 0 0 9 9 0 1 9 1 7 13 9 9 0 1 9 9 1 1 9 0 15 13 9 15 1 8 7 13 9 0 1 9 9 0 1 8 9 8 8 7 9 13 1 9 9 1 1 15 8 7 8 8 8 1 9 9 0 1 15 1 7 13 7 13 10 9 9 0 1 8 1 1 9 0 15 13 1 15 1 0 1 12 9 2
60 7 13 7 1 10 9 13 9 0 1 9 1 9 7 10 9 0 1 9 9 15 13 9 1 9 0 1 15 0 1 7 10 9 13 1 9 9 1 15 1 9 7 9 7 9 7 13 9 0 9 0 1 9 1 7 13 9 1 9 2
28 7 1 10 9 13 1 8 1 9 0 0 9 0 13 1 8 1 7 13 9 9 1 9 1 10 9 0 2
39 7 13 9 9 0 1 8 8 1 8 2 8 9 8 8 9 9 1 9 9 0 1 9 9 1 9 10 9 15 13 1 8 1 9 1 15 7 13 2
16 8 9 8 9 1 9 9 9 1 9 9 1 9 1 9 2
32 7 13 9 8 8 9 0 1 9 7 9 9 1 9 7 13 9 15 9 1 9 1 9 9 1 9 7 8 1 0 9 2
40 7 13 9 0 1 8 1 9 8 1 9 0 0 1 9 8 7 13 9 15 12 8 13 9 1 9 12 8 1 9 0 13 15 9 9 9 1 9 0 2
34 7 1 0 9 15 14 13 15 10 9 9 2 9 9 2 9 2 9 9 2 9 2 9 9 7 13 1 15 9 0 1 9 0 2
8 9 0 0 1 9 7 9 9
65 13 9 0 0 1 9 1 9 12 9 0 0 9 0 0 1 9 7 9 9 15 13 1 15 9 0 1 9 10 13 1 12 9 0 13 1 9 2 8 2 7 15 13 9 1 9 1 9 9 0 7 9 9 15 1 9 9 0 8 1 9 0 9 0 2
57 7 13 9 0 9 7 9 9 1 9 13 12 5 9 1 9 9 9 7 9 7 9 15 13 9 13 15 1 9 9 9 1 9 7 9 1 9 0 2 1 9 1 9 1 9 1 9 0 1 9 14 13 12 7 12 9 2
57 7 13 9 9 8 2 9 9 9 2 7 10 9 9 1 9 12 9 0 0 1 9 0 1 9 7 9 8 8 1 9 9 7 9 1 9 2 8 2 1 9 9 9 15 1 9 0 7 9 15 1 9 9 0 1 9 2
77 7 13 2 7 9 0 0 1 9 0 15 13 15 9 0 1 9 9 7 9 9 7 15 1 9 15 9 9 0 0 2 7 9 9 1 9 0 1 9 9 1 9 15 1 9 0 7 9 9 9 15 0 1 9 0 1 9 7 15 10 13 0 1 9 0 7 14 13 10 9 9 1 9 9 9 9 2
31 7 13 7 15 14 13 9 9 0 1 9 9 1 9 9 0 13 9 9 0 1 9 9 7 9 9 1 9 9 9 2
60 7 13 8 9 9 0 0 9 15 1 9 1 9 1 9 9 0 0 9 1 9 9 0 7 9 0 1 9 1 9 0 7 1 9 9 0 7 1 14 9 0 2 7 9 1 9 15 13 15 9 1 15 13 9 9 0 7 9 9 2
72 7 13 9 0 2 9 9 9 12 9 2 7 9 9 0 1 9 13 9 1 9 7 13 15 0 9 9 0 9 1 7 9 9 0 7 9 9 0 0 1 9 9 1 9 1 9 7 9 10 9 1 9 0 14 13 1 9 9 1 0 9 15 0 7 9 9 9 9 1 9 0 2
91 7 13 1 9 10 9 1 9 0 9 1 9 9 9 1 9 1 9 9 7 9 9 9 7 15 10 13 9 0 1 9 9 0 7 0 2 7 7 9 1 9 10 9 14 13 9 0 15 13 1 9 9 0 7 9 9 0 13 1 9 9 0 1 9 1 10 9 1 9 9 9 9 0 7 9 9 15 1 9 1 9 0 7 13 9 9 0 1 9 0 2
42 7 13 9 9 8 2 9 9 9 9 12 9 2 1 9 9 9 8 1 9 10 9 7 0 15 9 1 9 9 9 8 1 9 7 9 9 7 15 13 9 0 2
51 7 13 1 7 9 0 0 14 13 9 0 1 9 0 15 13 15 9 9 0 2 7 7 13 9 1 9 1 9 0 7 14 15 14 13 9 1 0 15 13 1 0 9 1 15 1 9 9 0 0 2
44 7 13 1 9 9 0 1 0 9 1 9 0 1 10 9 1 9 1 9 0 1 9 7 9 9 15 7 9 9 15 9 1 9 9 0 1 9 0 1 15 1 9 0 2
9 9 9 0 1 9 0 1 1 9
45 13 9 8 8 9 9 9 0 1 9 7 9 13 9 9 9 9 9 7 9 0 1 9 9 9 9 0 1 1 0 9 0 7 15 9 1 9 9 0 1 9 9 0 0 2
64 7 13 8 1 9 15 9 12 2 12 0 1 9 9 0 0 1 9 1 9 9 9 8 7 9 9 0 0 14 13 9 9 1 0 1 9 9 0 0 1 7 15 14 13 3 9 9 0 0 15 13 1 15 9 7 9 9 0 1 9 9 9 9 2
34 7 13 7 9 9 10 9 14 13 1 9 9 9 0 1 9 7 9 0 7 14 13 9 9 0 1 9 0 0 1 9 0 2 2
30 7 7 9 9 1 9 9 0 7 0 9 1 9 14 13 1 9 9 0 1 9 0 7 9 9 0 0 1 9 2
46 7 13 9 9 9 0 7 9 9 13 1 9 9 0 1 9 9 0 0 7 9 9 0 9 1 9 9 0 7 9 7 9 13 9 0 1 7 14 13 9 10 9 1 12 9 2
6 9 0 1 8 2 2
2 1 8
28 13 9 8 8 9 9 9 12 2 12 0 1 8 8 9 9 0 9 9 9 1 9 9 0 7 9 2 2
20 13 9 9 0 1 9 9 9 0 15 13 1 15 9 8 1 8 9 0 2
19 7 13 1 15 9 9 1 9 9 0 7 9 15 1 8 1 9 8 2
15 7 1 9 9 0 1 9 0 1 9 0 1 9 2 2
39 13 9 8 8 9 12 2 12 0 1 9 15 0 8 8 9 9 1 9 1 9 1 9 9 9 7 9 7 9 1 9 9 9 13 1 9 10 9 2
52 13 9 9 9 9 0 1 9 9 0 1 9 9 1 9 15 13 9 9 7 9 7 9 7 9 9 7 9 7 9 7 9 9 0 7 9 7 9 1 9 9 9 15 13 1 9 9 7 9 9 0 2
35 13 9 9 0 7 0 1 9 9 9 7 9 1 0 8 9 9 9 7 9 7 9 7 9 9 0 7 9 9 7 9 9 7 9 2
14 13 9 1 9 9 13 9 0 1 9 9 9 0 2
73 1 9 0 13 8 9 0 1 9 1 9 15 0 0 1 9 1 9 12 9 1 15 12 1 9 1 9 9 9 0 7 9 9 0 7 9 15 1 9 1 9 7 13 9 9 0 0 1 9 0 8 7 13 9 9 9 8 1 9 1 9 1 9 1 9 1 9 7 9 1 9 2 2
30 13 9 9 1 9 1 9 1 9 0 1 9 1 9 0 1 9 0 2 8 2 1 9 0 1 9 2 8 2 2
8 9 9 9 0 1 9 7 9
21 13 9 1 9 0 9 9 9 0 1 9 7 9 1 12 9 0 1 9 0 2
57 13 9 9 1 9 1 12 12 9 1 12 12 9 1 9 9 1 9 12 2 1 9 1 12 5 13 9 0 1 9 9 9 15 12 12 9 7 13 9 9 0 1 12 12 9 2 7 13 9 9 1 9 1 12 12 9 2
46 13 9 0 9 0 2 7 9 7 9 0 2 7 9 2 7 9 2 7 15 8 2 7 9 0 7 9 7 9 7 9 2 7 9 0 8 8 2 7 9 7 9 7 9 0 2
44 7 13 9 9 1 9 9 9 2 0 7 9 0 7 9 9 9 7 9 0 2 7 9 0 9 1 9 2 7 9 2 7 9 9 2 7 9 0 2 7 9 9 0 2
24 1 9 1 9 9 2 7 9 9 9 2 7 9 7 0 2 7 9 0 2 7 9 9 2
11 9 1 9 0 1 9 7 9 7 9 8
60 13 8 2 9 8 8 9 9 0 1 7 15 13 0 9 9 9 1 9 0 1 9 7 9 7 9 8 13 9 1 9 0 0 13 9 0 7 8 2 7 13 9 1 9 0 2 8 8 1 9 9 9 7 9 7 9 7 9 9 2
27 13 8 7 9 9 0 14 13 9 0 0 7 0 7 0 0 1 7 13 0 9 1 9 1 9 15 2
26 7 13 8 1 7 9 0 14 13 1 9 9 9 7 9 0 15 13 9 9 9 0 7 8 0 2
13 9 7 9 13 9 9 0 0 1 9 0 7 8
40 13 9 0 7 0 1 9 1 9 9 9 9 0 0 13 9 0 7 8 7 13 9 1 9 0 1 10 9 1 9 9 7 9 7 9 9 7 9 9 2
39 13 10 9 1 9 9 8 8 9 9 0 0 7 9 8 9 8 8 9 9 7 9 0 15 13 9 0 1 9 15 13 8 8 9 12 2 12 0 2
28 7 14 13 9 10 9 0 1 9 0 0 1 9 0 7 0 15 13 1 9 1 9 0 1 9 9 0 2
48 13 15 9 1 9 0 0 1 9 15 1 9 9 9 0 1 9 1 9 1 9 9 0 2 7 15 9 15 13 0 1 9 13 1 15 9 0 1 9 0 1 9 9 0 0 1 9 2
23 7 13 9 1 9 1 9 9 0 1 9 9 0 7 9 9 9 0 1 9 9 0 2
36 7 13 9 8 8 1 7 9 15 1 9 8 13 1 9 0 9 8 8 9 0 1 9 1 9 0 7 9 0 1 9 9 0 1 9 2
50 7 9 1 9 1 9 9 0 1 9 9 1 9 7 9 0 2 13 9 1 7 9 15 13 15 9 0 1 9 15 14 13 1 9 1 0 1 9 0 0 1 9 1 0 9 1 10 9 0 2
43 1 9 15 2 13 9 8 7 9 0 1 7 13 9 15 1 9 1 9 9 15 13 15 1 9 15 0 7 15 1 1 9 0 13 9 9 7 9 0 1 10 9 2
63 7 9 1 9 0 1 9 9 9 15 13 15 9 1 9 9 0 2 13 9 8 7 15 13 9 9 1 9 9 1 9 1 10 9 7 7 3 9 9 15 14 13 0 1 10 9 13 1 15 1 7 13 9 1 9 9 7 9 15 13 1 9 2
65 1 9 0 2 13 9 9 0 1 9 9 9 0 9 12 2 12 0 1 7 9 0 1 9 7 9 0 1 9 9 7 9 1 9 15 1 9 9 1 9 7 9 15 13 9 1 15 1 9 9 0 0 9 9 8 8 1 9 15 1 9 1 9 0 2
32 7 13 7 10 9 13 9 9 0 9 7 7 15 9 0 2 0 7 9 0 7 0 13 1 15 15 0 9 1 9 0 2
16 12 9 0 13 9 9 15 1 9 0 1 9 1 9 9 0
53 13 1 12 9 0 2 13 0 9 0 7 0 7 0 2 1 9 9 15 7 9 9 1 9 1 9 0 1 1 9 15 1 9 0 1 9 9 0 15 13 0 15 9 12 2 12 0 7 1 9 12 9 2
88 7 13 9 0 0 1 9 9 9 0 0 1 9 1 9 0 7 0 15 13 15 9 7 9 0 1 0 9 2 7 13 9 1 9 9 9 1 9 9 7 9 0 1 9 15 1 9 2 7 13 9 0 10 9 1 9 7 13 9 9 1 9 0 9 9 7 9 7 9 7 9 7 9 7 9 0 7 9 9 7 9 8 7 9 9 7 9 2
96 7 13 9 9 1 9 0 2 15 1 0 7 13 15 9 9 9 0 9 8 8 2 1 9 9 9 7 9 0 9 8 8 8 8 9 1 9 0 1 9 9 9 0 1 9 7 9 7 15 9 9 7 9 7 9 9 7 9 0 9 1 9 9 9 0 15 13 1 9 1 9 9 15 15 13 15 1 9 0 7 9 0 1 9 9 1 1 9 9 0 1 15 1 0 9 2
82 7 13 9 9 9 9 1 9 9 9 0 7 9 1 9 0 1 9 9 0 9 9 8 7 9 0 1 9 0 0 1 9 9 0 13 9 7 9 9 0 2 0 7 13 9 0 1 9 9 9 0 1 9 7 9 9 9 7 9 0 1 9 0 1 9 9 9 9 0 0 0 9 15 0 7 9 9 1 9 12 5 2
149 7 13 7 9 9 7 9 0 9 1 9 9 0 13 2 9 0 1 9 2 9 9 9 2 9 8 1 9 2 9 9 0 1 9 2 9 9 0 2 9 9 0 2 9 9 1 9 2 9 8 8 8 0 2 9 8 1 9 0 2 9 9 0 2 9 9 8 8 0 2 9 8 1 9 7 9 9 2 9 0 1 9 9 7 9 0 7 9 8 2 9 9 1 9 7 9 0 2 9 9 9 8 2 9 8 1 9 0 2 9 0 1 9 9 9 2 9 8 1 9 2 9 9 0 2 9 8 1 9 2 9 0 1 9 0 2 9 0 1 9 2 9 0 1 9 7 9 9 2
32 7 13 8 7 13 9 7 9 7 9 0 1 9 9 9 7 9 9 7 9 0 7 7 13 15 1 9 9 0 1 9 2
62 7 1 9 0 1 0 7 13 9 15 14 13 15 9 9 7 9 0 9 8 9 8 8 1 9 9 0 2 7 9 9 0 9 9 8 8 15 13 1 9 0 1 9 9 7 9 1 9 7 9 9 1 9 9 0 7 9 1 9 1 9 2
12 9 13 9 0 0 1 9 9 15 1 9 0
38 13 9 9 0 1 9 9 8 8 1 9 9 9 0 0 1 9 9 0 1 9 0 7 9 15 9 7 9 7 13 9 15 1 9 0 1 9 2
93 7 13 8 8 9 0 2 15 13 15 8 1 9 9 0 0 1 9 8 8 2 1 9 9 9 1 9 0 7 9 9 9 1 9 1 9 9 0 1 9 9 9 9 15 13 15 9 0 7 13 1 15 1 12 1 9 9 0 2 13 9 9 9 0 7 13 9 15 1 9 9 0 0 1 9 1 9 1 9 9 0 0 7 9 9 7 9 9 9 7 9 9 2
63 7 13 9 0 1 9 1 9 9 1 9 9 1 9 7 9 1 9 9 1 0 0 1 9 13 1 1 15 9 9 9 0 13 9 9 9 0 9 1 9 0 1 9 2 10 13 1 15 1 9 1 9 9 9 0 1 9 0 7 1 9 0 2
77 7 13 9 0 7 13 9 9 0 0 1 9 1 9 0 0 0 9 9 1 9 0 1 9 0 1 9 1 9 1 9 0 0 0 7 9 15 13 1 15 9 1 9 7 9 0 2 7 1 1 15 9 1 9 7 9 9 7 9 9 7 9 9 7 9 7 9 7 9 9 1 9 1 9 9 0 2
52 14 9 0 7 13 1 9 7 9 0 1 9 9 0 0 1 9 0 1 9 9 0 2 0 9 15 1 9 0 1 9 12 1 9 2 1 9 0 9 9 0 15 1 15 9 9 1 9 9 1 9 2
25 7 13 9 0 1 9 9 1 9 9 0 1 9 0 1 9 1 9 9 0 0 1 9 0 2
39 7 13 8 1 9 9 1 9 9 9 0 15 13 9 1 9 1 9 1 9 0 13 1 9 9 9 9 0 2 0 0 7 9 0 9 15 1 9 2
34 7 13 7 9 13 1 9 0 14 13 9 15 0 9 13 1 9 9 0 1 9 0 1 9 7 9 1 9 9 0 1 9 9 2
65 7 13 8 7 13 0 9 1 9 9 1 9 0 1 9 1 9 0 13 9 9 0 1 9 9 3 1 9 9 0 9 0 1 9 9 0 7 9 9 9 7 9 7 9 9 0 1 9 9 0 1 9 7 9 9 7 9 0 1 9 9 0 7 0 2
33 7 13 7 15 13 0 9 1 7 14 13 9 9 0 0 1 9 7 3 7 7 13 1 9 0 1 9 1 9 1 15 3 2
8 9 13 1 9 0 1 9 0
3 8 12 9
32 13 9 9 1 9 15 13 15 12 9 1 9 0 1 9 9 9 9 0 0 1 9 0 2 0 7 10 9 0 7 0 2
47 13 8 8 9 9 0 1 9 1 9 13 15 1 9 2 9 12 2 0 15 13 1 8 7 8 7 9 8 1 9 0 1 7 9 13 9 9 9 1 9 0 1 9 9 0 0 2
20 7 13 7 9 13 9 0 7 0 2 7 15 9 13 1 9 9 0 0 2
44 7 13 9 0 7 15 7 15 13 8 7 13 1 15 9 1 1 9 0 7 14 13 1 9 0 0 1 15 1 9 9 7 9 1 9 1 9 0 1 9 9 0 0 2
4 13 2 13 2
3 12 2 12
18 13 9 1 9 9 15 1 15 7 13 1 15 9 7 9 7 9 2
8 9 9 8 2 8 0 9 12
6 9 9 1 9 9 0
6 8 0 9 12 2 12
32 13 9 8 9 15 1 9 1 7 9 8 9 9 7 9 0 0 2 9 7 10 9 9 9 8 7 15 3 9 9 0 2
65 13 9 1 9 9 0 1 9 8 7 9 14 13 12 9 1 9 9 7 13 12 1 9 9 2 8 8 13 12 7 12 1 12 1 9 1 9 12 2 7 13 9 1 9 9 1 9 9 0 2 7 13 8 9 15 1 9 1 10 9 1 12 9 0 2
29 9 1 0 9 12 13 9 12 9 0 0 7 15 13 0 1 9 9 0 2 7 1 15 13 12 9 0 0 2
20 14 14 13 8 0 1 9 9 7 9 7 13 1 12 1 9 0 1 9 2
7 9 9 0 0 1 9 9
6 8 0 9 12 2 12
33 13 9 8 1 9 8 2 9 9 2 13 9 1 9 9 0 0 13 1 9 9 0 0 1 9 1 9 9 9 1 9 0 2
30 13 9 1 9 9 8 9 9 0 7 0 1 12 12 9 0 1 9 9 0 14 13 1 10 9 15 13 12 9 2
24 7 1 9 1 10 9 14 13 9 9 1 9 9 8 1 9 1 9 0 0 2 2 13 2
10 9 9 0 0 7 9 9 0 1 9
6 8 0 9 12 2 12
32 13 9 0 1 9 0 1 9 8 8 0 1 9 9 0 1 9 1 9 0 1 9 1 9 9 9 2 9 9 2 0 2
59 1 9 0 0 1 9 13 9 8 8 0 0 9 1 9 9 0 1 9 7 15 9 0 13 1 9 12 1 9 9 9 1 9 9 7 9 9 0 2 8 2 2 7 9 0 8 12 12 8 2 12 12 9 0 2 2 2 13 2
16 9 9 0 0 7 9 9 0 1 9 2 9 0 7 0 2
3 12 2 12
50 7 1 9 9 9 8 8 0 13 9 9 9 0 1 9 1 12 12 8 2 12 12 9 0 2 2 7 13 9 9 8 7 8 8 12 1 12 7 12 1 12 7 12 1 12 1 9 1 9 2
58 7 1 9 9 9 1 9 7 15 0 9 0 1 9 1 9 0 9 1 12 9 1 9 8 8 2 12 7 13 1 9 9 8 2 12 1 9 1 9 9 0 2 7 15 13 9 9 9 1 9 7 9 7 8 7 9 0 2
10 8 13 9 9 0 0 1 9 9 0
6 8 12 9 12 2 12
28 13 9 9 0 1 9 0 8 8 9 9 7 15 13 9 9 0 1 9 8 9 1 9 9 9 9 0 2
85 7 13 8 15 13 1 9 1 9 9 0 1 9 13 9 0 9 9 1 9 9 0 1 9 2 2 13 1 9 9 9 0 7 13 1 15 9 7 9 0 0 2 2 7 13 10 9 0 1 12 9 0 13 0 9 0 7 0 1 9 9 7 9 15 2 7 13 9 1 9 9 13 1 9 9 0 1 9 12 9 1 9 9 0 2
33 7 13 8 1 9 1 7 9 15 13 15 8 1 9 13 7 13 9 9 1 9 0 1 9 12 9 1 9 9 0 1 9 2
36 7 13 8 7 9 0 15 13 15 9 0 1 9 2 9 9 8 8 7 9 15 0 8 8 2 13 7 13 1 8 8 3 1 10 9 2
38 7 13 8 2 8 8 14 13 1 10 9 1 9 9 9 9 2 2 0 7 9 0 15 13 15 0 9 0 2 14 13 1 9 1 9 9 9 2
10 9 9 13 1 9 15 1 9 1 9
7 8 8 12 9 12 2 12
19 13 9 9 9 0 12 9 13 1 9 15 1 9 9 1 8 9 9 2
48 7 13 9 1 9 9 5 2 8 8 5 2 0 13 1 3 7 15 13 1 9 9 9 0 1 9 7 9 7 9 15 13 7 15 13 14 13 1 9 1 9 0 1 9 0 1 15 2
12 7 13 9 7 15 13 0 9 1 10 9 2
11 9 9 9 13 9 1 9 9 0 1 9
6 9 12 9 12 2 12
111 13 9 8 8 9 9 9 0 7 9 1 9 9 9 1 9 9 9 15 9 9 9 9 0 0 13 1 9 1 9 1 9 15 0 1 9 0 1 9 2 7 13 8 1 9 1 9 0 0 7 10 9 13 1 9 9 1 9 0 1 9 10 13 9 1 15 1 9 1 9 9 0 7 0 1 10 9 2 2 7 7 9 0 1 0 9 1 9 0 13 1 1 9 2 7 13 1 7 9 13 9 1 9 9 9 0 1 9 15 0 2
22 13 7 11 8 15 9 9 9 8 9 9 0 1 9 0 1 9 7 9 15 9 2
37 1 9 15 13 8 8 9 9 0 0 7 9 15 13 9 1 9 13 1 9 9 0 0 13 9 0 7 0 1 9 1 9 9 9 9 0 2
7 9 0 1 9 7 9 0
6 9 12 9 12 2 12
129 13 8 8 11 8 8 9 9 7 9 0 9 0 1 9 8 9 15 1 8 8 9 9 0 1 7 15 13 0 7 9 9 1 9 1 9 0 1 9 0 0 1 9 9 0 1 9 9 0 1 9 7 1 9 9 9 0 7 1 0 10 13 1 9 9 7 9 1 9 9 0 2 7 13 8 1 9 0 0 13 15 1 9 0 9 7 13 15 9 9 0 9 15 1 0 9 13 1 15 9 1 9 9 0 0 7 9 15 0 7 9 13 1 9 0 1 0 9 1 9 9 1 9 7 9 1 9 0 2
39 7 13 7 8 13 9 1 0 9 13 7 13 0 1 9 0 7 9 9 1 9 9 0 1 9 15 1 9 9 9 0 1 9 0 7 9 1 9 2
67 7 1 9 15 13 8 8 9 9 0 7 9 15 1 9 0 13 9 9 9 9 1 9 1 9 0 7 15 13 1 9 1 9 0 0 7 9 15 1 9 13 1 9 1 9 9 1 9 9 9 1 9 1 9 9 9 1 9 9 1 9 7 9 1 9 0 2
28 7 1 15 13 1 9 0 1 9 9 0 13 9 0 7 9 9 15 15 13 1 15 7 13 9 9 15 2
8 9 0 0 1 9 1 9 0
6 9 12 9 12 2 12
52 13 1 8 9 1 9 7 15 13 1 9 0 8 9 1 9 1 9 1 9 0 1 9 0 7 9 13 15 1 9 0 8 8 8 9 9 1 9 9 1 9 0 0 7 1 9 0 9 9 8 8 2
55 7 13 9 9 1 9 1 9 9 9 7 9 1 1 9 9 1 9 0 1 9 7 9 7 9 9 7 9 7 9 1 9 7 9 9 0 7 9 9 9 0 7 0 1 9 9 9 9 9 0 7 9 9 0 2
60 7 13 9 9 1 9 0 0 1 9 9 9 0 7 9 9 9 9 7 9 9 9 1 9 0 7 9 1 9 9 7 9 9 8 1 9 7 9 9 1 9 9 9 9 7 9 9 9 0 1 9 9 0 7 9 7 0 7 0 2
10 8 8 8 13 9 9 0 1 9 9
6 8 12 9 12 2 12
22 13 9 9 0 0 2 8 8 8 2 9 9 0 1 9 1 9 9 1 9 9 2
52 7 13 9 13 15 8 8 8 9 9 1 1 12 12 9 0 7 0 1 9 9 2 7 9 9 0 0 1 9 9 9 1 15 2 1 15 1 15 9 9 1 9 9 7 9 9 1 9 0 1 9 2
25 7 13 9 1 7 15 13 1 9 9 9 9 9 0 1 9 0 9 13 1 9 0 1 9 2
32 7 1 9 1 15 2 13 1 8 8 8 9 0 1 9 0 9 0 1 0 1 9 9 0 0 9 15 12 9 1 9 2
19 7 1 9 12 9 2 13 9 0 9 0 1 9 9 9 0 1 9 2
20 7 13 9 9 2 9 9 2 1 9 9 9 0 0 1 9 0 1 9 2
7 9 8 9 9 0 1 8
6 9 12 9 12 2 12
67 13 1 9 0 1 9 7 9 9 0 13 1 9 7 13 9 0 9 7 9 15 1 9 15 7 13 9 1 9 0 7 9 9 0 7 13 1 9 9 0 7 9 9 0 1 9 9 1 9 9 1 9 9 9 9 9 1 9 0 1 9 8 1 9 1 10 2
60 7 13 9 1 9 0 0 1 9 9 9 9 1 9 9 0 1 9 9 9 1 9 9 1 9 9 9 0 1 9 0 1 9 7 9 9 9 1 9 0 1 9 0 0 7 13 1 9 9 0 1 9 0 9 7 9 1 10 9 2
61 7 13 1 9 9 0 0 1 9 0 1 9 12 1 12 1 9 0 8 7 9 1 9 1 9 1 10 9 0 9 9 9 9 7 9 15 1 9 9 1 9 9 0 1 9 8 7 9 8 8 7 9 9 0 1 9 9 1 9 0 2
10 0 9 9 0 9 1 9 8 1 9
6 8 0 9 12 2 12
35 13 9 8 0 1 9 8 9 9 8 0 9 9 9 1 13 9 9 0 9 1 9 8 9 9 2 7 15 0 1 9 15 1 9 2
24 13 7 10 9 0 9 1 9 9 0 7 1 9 15 7 13 9 0 1 9 8 7 0 2
44 13 9 1 10 9 7 10 9 13 9 15 1 9 9 7 13 9 9 8 7 0 1 9 1 10 9 9 1 9 15 1 9 7 9 9 1 9 0 0 2 2 9 9 2
13 9 0 13 9 12 12 1 9 1 9 9 1 9
6 8 12 9 12 2 12
25 13 9 0 9 0 9 9 1 9 0 1 12 12 1 9 1 9 9 1 9 1 9 9 9 2
22 7 13 10 9 1 9 15 13 1 15 9 1 9 0 0 9 1 15 1 9 0 2
47 7 13 10 9 2 1 9 1 12 12 0 1 9 0 2 9 12 1 12 1 0 9 9 1 9 9 7 0 12 9 2 7 1 0 7 13 9 9 9 9 13 1 12 12 9 0 2
30 7 13 9 9 9 7 9 0 0 9 15 12 12 9 14 13 9 15 1 9 12 9 7 9 1 9 12 9 0 2
73 7 13 9 0 8 8 8 1 9 0 1 10 9 9 9 0 0 1 9 0 15 14 13 1 12 9 0 2 1 12 12 9 0 2 7 15 0 1 9 9 0 2 7 1 9 1 15 2 13 9 7 9 9 0 14 13 1 12 12 9 0 1 9 0 7 15 13 9 9 9 1 9 2
8 9 9 0 0 13 9 9 9
6 8 0 9 12 2 12
44 13 9 9 1 9 0 9 0 0 1 9 1 9 8 7 9 8 1 9 9 13 12 12 8 2 1 15 1 12 12 8 13 15 9 9 0 0 1 9 0 9 1 9 2
46 7 13 9 9 7 9 9 9 0 8 8 9 4 3 13 9 9 0 1 9 9 7 13 3 9 0 1 9 9 9 1 9 8 9 1 9 9 7 9 8 9 1 9 0 9 2
62 7 13 10 9 0 1 12 9 15 9 8 2 8 0 7 9 0 0 1 9 8 7 9 0 1 9 8 8 2 7 9 15 0 12 8 2 7 1 0 7 13 9 9 9 1 15 12 12 9 0 1 9 12 2 7 12 12 9 1 9 12 2
7 9 0 0 1 9 0 0
6 8 0 9 12 2 12
60 13 9 1 9 8 0 1 9 8 2 9 0 9 2 9 1 9 9 0 1 9 9 0 0 13 8 8 1 0 1 12 9 8 8 1 9 8 12 9 2 12 8 2 1 9 2 8 8 15 0 9 13 1 15 0 0 1 10 9 2
89 7 13 9 7 9 0 1 9 9 8 1 9 8 2 8 9 9 2 14 13 1 9 8 1 9 8 0 9 2 8 9 9 2 2 8 8 8 1 9 9 15 1 12 9 7 15 9 9 7 9 7 9 7 9 2 14 0 7 15 1 9 0 0 9 14 13 9 15 7 9 9 15 7 9 15 7 9 15 0 0 7 9 15 0 1 9 9 0 2
3 2 13 2
11 9 0 0 1 9 0 0 2 9 0 2
3 12 2 12
72 9 0 0 1 9 0 0 2 9 0 2 7 13 9 8 14 13 9 8 1 9 9 0 1 9 2 7 13 7 13 10 9 1 8 9 1 9 9 0 0 1 9 1 9 1 9 15 15 13 1 9 8 8 9 8 13 9 15 1 9 9 8 2 12 1 9 1 12 1 9 2 2
41 13 8 8 8 1 9 7 9 9 9 0 1 9 9 0 0 0 1 9 9 0 1 9 7 15 13 0 9 9 9 9 0 9 0 9 0 0 7 9 0 2
3 2 13 2
13 9 0 0 1 9 0 0 2 9 0 7 0 2
3 12 2 12
37 9 0 0 1 9 0 0 2 9 0 7 0 2 7 13 8 8 7 9 13 9 1 9 9 9 13 1 9 9 9 0 1 9 1 9 9 2
50 9 1 15 13 9 9 8 8 0 1 9 9 7 9 9 15 1 9 15 13 1 9 9 5 2 8 8 5 2 0 1 9 8 2 8 0 9 2 7 13 1 0 9 9 0 13 9 0 3 2
50 0 1 9 7 12 9 0 0 13 1 9 0 1 9 1 9 0 1 9 8 1 8 7 13 9 0 1 9 2 7 14 13 1 9 0 1 9 0 3 13 9 9 7 9 9 1 9 9 0 2
11 9 0 2 9 9 0 1 9 9 9 0
6 9 12 9 12 2 12
72 13 9 0 7 0 0 7 9 9 9 9 0 7 9 9 9 9 7 9 9 7 9 7 9 9 9 1 9 13 9 9 9 0 7 9 9 9 0 1 9 7 9 7 9 9 0 7 15 13 1 9 15 1 9 0 7 1 9 9 9 7 9 9 7 9 0 1 9 0 1 15 2
36 7 13 10 9 1 7 9 13 9 9 0 1 9 7 9 9 0 1 9 9 1 9 1 9 15 13 9 15 7 9 15 7 9 9 15 2
170 7 13 7 9 0 13 1 9 9 15 13 1 15 9 0 1 9 9 8 11 8 8 9 0 1 9 9 9 9 7 9 7 13 9 0 8 8 13 1 9 9 9 9 0 7 9 9 9 9 2 7 13 9 7 9 9 1 9 1 9 7 9 1 9 1 9 13 1 9 9 15 13 1 15 10 9 7 1 9 9 15 1 9 7 9 0 7 7 9 9 1 9 1 9 9 9 9 7 9 15 1 9 9 7 1 9 1 8 8 7 1 9 9 9 9 9 15 13 1 9 0 1 10 9 2 7 13 9 9 1 9 0 7 9 15 1 9 1 9 0 1 9 7 1 9 1 9 9 7 9 7 1 9 9 9 7 9 1 9 7 9 9 0 1 9 0 1 9 0 2
25 7 13 9 7 9 0 7 0 0 13 9 9 0 0 1 9 10 9 7 13 1 9 9 9 2
45 7 13 9 9 1 9 0 9 9 1 9 8 8 7 9 9 0 1 8 0 13 9 9 9 8 8 9 9 7 9 7 9 9 0 1 9 7 9 7 9 7 9 7 9 2
29 7 1 0 7 13 9 9 0 0 9 15 1 9 9 15 9 9 0 7 14 13 9 9 9 0 1 9 0 2
5 9 0 0 7 0
6 8 12 9 12 2 12
42 1 15 13 9 1 9 0 0 7 0 2 9 2 2 13 9 2 9 2 1 9 1 9 9 0 2 0 0 1 9 9 1 9 12 1 9 7 0 9 1 9 2
39 7 13 9 15 13 15 9 9 9 1 9 9 1 9 7 13 12 9 2 1 9 9 0 1 9 9 7 9 1 9 0 7 0 1 9 9 9 9 2
32 9 2 2 13 9 9 9 0 0 2 0 2 8 2 15 13 13 1 9 9 7 9 0 1 9 9 9 1 9 0 9 2
34 7 13 8 2 2 8 8 8 2 2 0 7 15 13 3 9 1 9 9 9 0 1 9 1 9 14 13 1 9 9 0 7 0 2
49 7 13 7 10 9 15 15 13 9 9 0 1 9 9 1 12 9 13 1 9 9 1 15 8 7 8 7 8 7 9 8 0 1 9 9 15 1 9 9 9 9 0 1 9 9 15 1 9 2
34 8 2 2 13 9 9 0 0 1 9 0 8 9 1 9 8 7 9 13 9 1 9 9 9 0 8 8 8 15 13 1 9 0 2
31 13 9 9 0 1 9 13 1 12 9 13 8 8 1 9 9 7 9 8 8 8 1 9 1 9 8 15 13 9 15 2
41 7 13 9 15 13 1 0 7 12 1 9 0 2 1 9 0 9 8 1 9 9 7 8 1 9 9 0 8 8 8 9 1 9 15 15 13 15 1 9 0 2
3 2 13 2
5 9 0 0 7 0
3 12 2 12
42 2 9 0 7 0 2 8 2 2 13 9 8 8 1 8 9 13 1 15 9 1 9 0 1 1 15 9 13 9 0 1 9 0 8 8 8 13 15 1 9 0 2
12 7 1 0 7 13 9 1 12 12 9 0 2
28 7 13 7 8 8 8 13 1 9 12 7 13 1 9 12 2 7 14 13 1 15 9 15 1 9 9 0 2
33 8 2 2 13 8 9 9 0 8 8 0 9 1 15 1 9 2 8 9 8 8 2 15 13 1 15 1 9 0 12 12 9 2
38 7 13 9 15 13 1 9 12 7 13 9 7 15 1 0 7 12 1 9 15 1 9 15 9 9 7 9 7 9 7 9 0 1 9 1 9 0 2
39 13 7 10 9 0 13 1 15 12 8 13 9 15 0 1 12 9 2 7 14 13 9 8 9 0 13 1 15 1 9 1 12 12 9 7 8 12 9 2
11 9 9 0 1 9 9 1 9 9 9 12
6 8 0 9 12 2 12
17 13 9 9 9 0 1 9 9 1 9 9 9 12 1 9 8 2
51 7 1 9 1 9 12 14 13 9 9 9 12 12 12 8 1 9 0 1 9 7 9 9 12 12 9 1 12 9 7 9 0 7 9 0 1 12 9 0 7 0 7 9 9 12 12 9 0 1 9 2
56 9 9 12 1 9 8 15 0 9 9 1 9 2 7 1 3 14 13 0 1 12 9 1 15 0 2 7 15 13 1 12 9 7 9 0 1 9 8 7 9 8 2 7 1 9 13 9 9 12 12 9 1 9 9 10 2
10 9 9 9 0 0 1 9 9 1 9
6 9 12 9 12 2 12
64 13 1 9 9 9 2 9 2 9 9 0 0 15 13 13 9 9 9 2 7 13 9 0 0 7 9 0 13 9 0 1 9 7 1 1 15 8 8 9 9 0 0 8 8 8 9 9 0 0 8 8 8 9 9 9 9 0 7 9 15 1 9 9 2
44 7 13 9 1 7 9 0 13 9 1 9 9 7 9 1 8 8 9 9 9 0 7 9 9 8 9 7 9 9 9 8 9 9 0 1 9 0 1 9 7 9 15 9 2
8 9 1 9 0 1 9 9 9
6 9 12 9 12 2 12
96 13 9 0 0 9 2 9 2 7 15 14 13 9 1 9 0 13 9 15 1 15 13 1 12 12 9 1 9 9 9 0 9 2 7 13 8 2 8 8 8 2 0 7 9 0 0 13 7 9 13 1 12 12 7 12 12 9 1 12 9 0 2 7 13 9 7 9 13 9 1 9 9 1 9 9 1 9 1 9 9 7 1 9 14 13 9 15 1 9 1 9 1 9 9 9 2
67 7 13 7 9 0 1 9 0 13 1 15 1 9 10 1 12 7 12 9 0 1 9 1 9 13 1 9 15 9 9 0 9 0 1 9 0 2 7 13 1 7 9 0 13 1 9 0 1 12 12 9 1 9 9 15 1 9 0 7 13 9 9 1 9 9 0 2
8 9 9 0 7 0 0 1 8
6 8 0 9 12 2 12
25 13 8 8 8 8 9 0 1 9 8 0 0 1 9 1 9 9 9 0 7 0 0 1 8 2
7 7 14 13 10 9 0 2
31 7 13 9 9 9 1 9 9 7 9 14 13 8 9 1 9 1 9 9 9 1 0 1 1 8 8 8 7 8 0 2
18 15 7 14 13 9 0 7 0 0 9 1 9 9 9 7 8 8 2
11 9 0 2 9 14 13 1 9 0 1 9
6 9 12 9 12 2 12
73 13 9 8 8 9 9 0 7 9 15 14 13 1 9 0 1 9 2 7 13 8 1 9 1 9 9 0 7 9 15 14 13 1 9 9 9 0 1 9 2 2 7 13 9 9 0 7 0 1 9 9 1 9 0 2 7 13 7 15 14 13 7 9 1 9 7 9 0 14 13 1 9 0
8 0 2 9 0 13 9 0 8
6 8 12 9 12 2 12
30 13 9 0 9 0 0 9 0 8 1 9 0 1 9 2 9 5 2 1 7 13 9 0 1 9 1 9 7 9 2
24 7 13 9 15 13 9 0 1 9 15 1 12 2 12 9 2 1 1 9 0 7 9 9 2
11 9 9 1 8 0 1 9 15 1 9 0
6 8 0 9 12 2 12
32 13 9 0 7 9 9 8 0 7 13 15 9 9 2 7 1 9 7 7 9 9 1 8 0 1 9 15 1 9 9 0 2
34 15 15 13 1 15 8 8 9 0 1 9 9 0 1 9 0 0 1 9 7 9 1 9 1 9 0 13 15 1 15 9 8 0 2
30 7 13 10 9 7 9 1 12 9 0 7 9 9 1 8 13 12 1 12 1 9 1 12 1 12 1 9 9 15 2
49 7 1 9 15 13 15 9 9 0 1 12 9 12 7 14 9 9 1 9 0 1 9 9 13 1 12 7 12 1 12 0 2 7 13 1 15 7 9 9 1 9 0 0 1 9 15 1 8 2
10 9 0 13 9 7 9 0 1 9 9
6 9 12 9 12 2 12
158 13 9 9 0 9 0 1 9 0 7 0 1 9 0 0 2 7 13 9 9 9 8 8 1 9 1 15 9 9 7 9 15 13 1 0 1 9 13 12 9 0 0 9 7 9 7 12 9 0 0 7 9 1 9 0 7 12 9 0 1 9 0 0 0 1 15 9 9 7 9 7 9 9 7 9 9 2 7 13 9 12 9 0 1 9 0 7 9 9 9 0 7 9 0 0 1 15 2 9 9 9 2 7 9 8 8 9 1 9 8 0 7 12 9 0 7 12 9 0 7 12 9 0 8 8 8 7 9 15 7 9 0 2 7 13 9 0 7 9 13 3 1 9 9 1 9 8 7 9 0 7 9 0 1 9 9 0 2
32 7 13 8 7 0 9 0 7 9 13 13 9 15 1 9 9 9 7 13 9 1 15 7 9 15 7 9 15 1 9 0 2
65 7 13 9 9 0 14 13 7 1 9 0 1 9 9 7 9 0 0 1 9 9 15 0 1 9 9 1 9 10 13 1 9 9 1 9 15 0 1 0 9 0 7 9 7 9 13 9 15 1 9 0 1 9 7 1 0 13 1 9 15 7 13 9 15 2
8 9 9 8 12 1 9 9 0
6 8 0 9 12 2 12
18 13 9 9 0 14 12 9 9 1 9 8 9 9 8 1 9 9 2
32 7 1 9 1 9 9 0 7 9 8 13 9 9 9 9 15 12 12 9 0 1 10 9 15 13 12 9 7 13 9 0 2
49 7 13 9 9 0 1 9 9 9 7 0 7 9 9 7 9 7 9 0 1 12 12 7 12 12 7 12 12 9 0 1 9 0 12 1 12 7 12 1 12 7 12 1 12 1 9 9 9 2
43 7 14 13 10 9 12 9 1 12 9 7 9 1 9 7 1 1 15 12 9 0 2 7 0 1 9 7 15 14 13 0 9 8 1 9 9 7 9 9 9 1 15 2
13 0 2 9 13 1 9 1 2 9 9 2 9 0
6 8 0 9 12 2 12
27 13 9 0 9 9 9 1 9 15 7 9 15 1 9 1 5 2 9 9 5 2 1 9 1 9 0 2
28 7 9 1 9 13 8 8 8 9 1 9 9 9 0 7 9 13 1 9 0 1 2 9 9 2 9 0 2
54 7 13 9 7 9 13 1 7 13 9 0 7 0 1 10 9 0 7 13 9 0 1 9 0 1 9 15 13 15 9 0 7 9 10 9 7 9 9 9 7 9 9 7 9 0 1 9 9 0 1 0 9 0 2
8 8 13 1 9 9 1 9 8
6 8 12 9 12 2 12
27 13 9 9 0 8 8 1 9 1 9 15 0 13 1 15 1 9 9 7 9 1 9 1 9 9 8 2
37 7 13 8 1 9 15 15 13 15 1 8 8 8 9 9 7 9 0 13 1 9 1 10 9 0 15 13 1 15 9 9 0 0 2 8 2 2
34 7 13 8 1 9 9 1 9 8 7 9 15 1 9 9 0 2 0 1 13 15 1 7 13 9 1 9 1 8 1 0 9 0 2
17 7 13 9 7 8 14 13 9 7 9 1 9 9 1 9 8 2
10 8 13 1 9 0 9 2 9 9 2
6 8 12 9 12 2 12
35 13 9 9 0 8 8 8 9 9 7 8 14 13 9 9 2 9 9 2 0 1 9 2 9 1 9 9 0 2 0 1 9 9 0 2
18 7 13 8 8 1 15 1 9 9 1 15 13 12 9 1 9 0 2
33 7 13 1 7 9 2 9 9 2 1 9 13 1 9 9 1 9 1 8 7 8 7 15 13 1 9 0 13 1 15 9 0 2
37 7 13 9 9 1 10 9 0 1 9 2 9 9 2 7 15 13 1 9 0 1 9 9 0 1 9 9 12 2 1 9 1 9 0 7 0 2
73 7 13 9 9 0 2 7 15 7 1 0 9 1 12 2 13 8 0 1 9 12 13 1 9 9 0 0 1 9 7 9 9 2 1 9 9 9 8 13 9 0 1 9 15 7 9 9 15 2 2 7 1 9 9 15 2 13 8 8 9 1 9 1 9 9 0 1 9 7 9 9 0 2
21 7 13 9 3 9 1 9 9 15 1 8 0 7 9 9 9 0 1 15 8 2
43 7 13 9 2 9 9 2 15 13 15 9 1 9 0 7 8 7 9 0 7 9 0 2 1 9 9 0 1 12 9 1 9 7 9 7 9 9 0 1 9 12 9 2
5 9 1 9 9 8
6 8 0 9 12 2 12
131 13 9 2 9 0 2 0 9 9 3 1 9 15 0 9 1 9 9 9 0 0 0 9 2 13 9 1 9 7 9 7 9 7 9 9 1 9 9 9 9 0 7 0 1 15 15 13 1 9 0 1 9 8 2 7 13 9 7 9 9 9 0 8 8 8 13 8 0 1 9 9 9 1 9 15 9 9 9 7 9 0 1 9 8 2 7 13 9 2 8 8 8 2 7 9 9 9 0 8 8 8 13 1 9 9 7 9 9 1 9 8 7 15 1 9 13 15 1 9 0 1 9 7 9 1 9 8 2 2 13 2
11 9 1 9 9 8 2 9 0 7 0 2
3 12 2 12
31 7 13 9 2 9 0 2 7 9 9 8 1 9 0 0 13 1 12 12 1 9 9 12 1 9 12 12 1 9 0 2
20 13 9 2 8 0 2 1 9 9 0 0 1 9 8 1 9 9 9 9 2
45 7 13 8 8 1 9 8 0 7 1 15 0 1 12 9 2 13 9 2 8 0 2 7 9 9 0 2 8 8 8 8 2 14 13 9 0 1 9 9 0 15 13 12 9 2
46 7 13 3 7 9 9 0 13 9 0 1 9 7 9 1 9 8 1 9 8 0 9 0 9 9 9 1 9 9 0 1 9 10 9 1 9 7 8 14 13 0 1 0 9 8 2
6 9 9 1 9 1 8
3 9 0 9
24 13 9 0 7 9 0 13 9 9 1 9 9 0 1 9 8 0 1 9 8 9 9 0 2
45 7 13 9 7 8 8 8 2 12 9 2 13 13 9 15 1 9 1 9 13 1 9 0 7 9 8 1 8 0 1 9 15 7 13 9 0 9 1 9 15 7 13 15 9 2
7 9 0 13 9 8 9 8
3 9 0 9
19 13 9 0 1 9 0 1 9 9 9 8 9 9 8 1 9 9 9 2
28 7 13 9 9 7 9 0 7 9 0 1 9 0 13 9 1 9 0 1 9 9 1 9 9 9 0 0 2
24 7 13 1 9 0 13 1 9 9 1 9 0 7 9 9 0 7 13 1 9 9 1 9 2
10 8 13 1 9 9 1 9 9 15 0
3 9 0 9
40 13 9 9 0 8 8 9 15 0 9 9 1 9 1 9 9 9 8 8 8 1 9 15 1 9 9 15 13 15 9 0 1 9 1 9 1 9 8 8 2
30 7 13 8 1 9 9 9 8 11 8 8 7 9 0 1 9 9 9 9 9 8 8 8 7 9 15 1 9 0 2
33 7 13 9 8 1 9 1 9 15 1 9 0 1 9 3 9 7 9 15 0 1 9 9 1 9 9 0 1 9 1 9 9 2
30 7 13 9 9 0 15 13 1 9 0 9 12 9 9 9 13 1 9 0 1 9 9 12 7 9 9 15 13 15 2
17 7 1 10 9 13 9 0 1 9 9 0 0 0 1 9 0 2
27 7 13 9 0 7 0 13 8 8 1 9 8 7 9 8 8 1 9 1 9 9 9 1 9 9 9 2
12 7 13 9 0 1 9 7 9 0 1 9 2
44 7 13 0 1 12 12 1 9 0 7 0 14 13 1 9 0 0 1 12 9 1 9 13 15 8 3 1 9 1 7 15 2 14 13 0 9 1 9 1 9 0 0 2 2
15 7 1 0 7 13 9 9 0 9 1 9 0 1 9 2
13 9 12 9 1 9 0 7 9 2 2 8 2 2
3 9 0 9
45 13 12 9 1 1 15 9 1 0 1 9 15 7 13 12 1 9 9 9 1 9 9 0 9 13 1 15 9 0 1 9 9 9 9 9 7 9 8 9 9 8 1 9 0 2
34 7 13 9 9 0 7 12 9 9 1 9 0 1 9 0 13 1 9 0 1 9 0 1 9 9 7 1 9 0 1 9 8 0 2
9 7 13 9 1 0 0 12 9 2
28 7 13 9 1 9 9 9 0 7 0 1 12 9 7 9 0 0 13 1 9 9 9 1 9 9 8 8 2
39 7 13 9 8 8 9 0 9 7 9 1 8 9 1 9 7 2 9 9 9 0 1 9 9 0 1 9 9 9 9 13 1 12 1 15 9 0 2 2
28 7 13 1 7 0 9 15 8 8 8 7 14 13 9 15 9 7 14 13 1 9 1 9 13 15 9 0 2
55 7 14 13 9 0 7 9 8 8 2 12 9 2 8 8 8 8 8 8 8 2 12 9 2 8 8 8 8 2 12 9 2 13 1 9 15 1 9 9 0 1 9 9 1 9 9 7 14 13 9 1 9 0 9 2
21 7 13 9 1 9 9 0 7 12 1 9 15 13 1 9 1 9 9 9 9 2
38 7 13 9 9 9 0 1 9 8 1 9 1 15 7 2 9 1 9 9 0 1 9 9 13 1 9 7 9 1 9 15 1 9 0 1 9 2 2
50 7 13 9 0 1 10 9 9 9 13 1 9 0 0 2 7 13 9 9 0 1 9 0 8 8 8 7 9 0 13 9 15 7 9 0 1 12 9 7 13 1 9 7 0 1 9 7 9 0 2
39 1 9 0 13 9 0 7 0 1 12 9 7 9 0 0 13 15 9 9 13 1 9 9 1 9 0 0 1 9 9 7 9 0 1 9 1 9 8 2
22 7 13 9 7 9 0 13 12 9 9 0 9 1 12 9 0 1 9 0 1 9 2
40 7 1 9 8 9 8 13 9 0 7 9 13 1 9 9 0 1 9 9 0 1 9 1 9 0 1 9 9 9 2 9 7 9 9 13 9 9 1 0 2
36 7 13 9 0 1 9 0 1 9 0 15 13 1 8 8 7 13 15 9 1 9 9 8 8 8 7 9 9 9 9 0 0 1 9 8 2
33 7 13 9 1 9 1 13 8 8 2 8 8 2 9 15 1 0 9 1 9 1 9 0 7 13 9 0 7 0 9 9 9 2
16 9 0 13 1 9 9 1 9 9 9 1 9 0 1 9 9
60 9 0 13 1 9 9 1 9 9 9 1 9 0 1 9 9 9 0 12 9 2 8 2 13 9 0 9 1 9 0 1 9 9 1 9 1 9 9 1 9 9 9 2 0 9 1 9 9 7 9 9 0 1 9 1 9 0 0 9 2
57 7 13 9 9 0 1 9 0 8 8 1 9 1 9 9 0 1 8 8 1 9 9 0 15 13 12 9 7 15 14 9 1 9 9 9 2 1 9 15 2 9 9 2 7 2 9 9 2 1 9 1 9 7 9 7 9 2
35 7 13 1 9 9 1 0 1 9 9 2 0 1 7 0 15 13 1 9 15 1 9 15 14 13 1 9 7 13 13 1 9 9 0 2
63 7 9 1 9 9 0 7 14 12 9 13 1 9 1 12 1 12 2 7 1 1 15 12 13 13 2 7 13 12 0 1 9 9 15 0 2 7 13 12 1 9 9 15 1 9 9 9 2 7 13 12 1 9 9 1 7 15 13 9 15 1 9 2
38 13 10 9 15 13 15 9 9 0 1 9 0 1 9 9 9 9 2 7 15 9 0 1 9 0 1 9 0 0 1 9 0 1 9 0 1 9 2
6 9 9 0 0 1 9
3 9 12 9
36 13 9 0 7 9 9 9 9 9 7 9 0 0 13 1 9 0 1 9 9 0 1 9 1 9 0 0 1 9 9 7 9 0 1 9 2
44 7 13 9 7 9 0 13 9 1 8 8 2 12 9 2 7 15 9 0 13 1 9 9 0 1 9 9 0 2 8 8 8 2 7 13 1 9 15 1 9 2 0 2 2
37 7 13 8 1 8 1 9 9 1 9 7 9 9 0 1 2 9 9 2 15 13 15 9 0 1 9 15 9 15 13 9 0 1 9 7 9 2
43 7 13 9 9 13 1 9 1 15 7 9 0 13 9 1 8 7 9 1 9 15 1 8 0 1 9 15 2 1 7 15 13 9 0 7 13 9 13 1 9 15 2 2
28 7 13 2 8 9 9 1 9 7 9 13 8 9 15 1 9 15 7 13 13 9 1 9 7 15 13 2 2
31 7 13 9 1 7 9 0 13 1 15 1 9 9 2 7 13 9 2 7 13 9 9 13 9 1 9 9 0 0 2 2
25 7 1 9 13 9 0 9 9 0 13 9 9 0 13 1 9 15 1 9 9 9 9 1 9 2
17 7 1 15 1 9 13 9 0 0 1 9 9 0 1 9 15 2
74 7 13 9 0 0 9 9 7 8 13 1 9 9 15 1 9 9 0 9 1 9 7 14 13 9 9 15 1 9 2 1 9 7 9 0 15 13 9 15 9 9 1 9 0 1 8 8 7 9 0 13 7 13 1 7 15 9 1 15 13 8 8 8 1 9 9 7 13 9 1 8 8 8 2
7 9 0 13 9 9 0 0
3 8 12 9
32 13 9 0 8 8 8 3 9 9 1 9 9 0 0 9 8 8 9 0 1 9 1 9 9 0 8 8 9 9 1 9 2
21 7 13 1 9 9 9 1 9 0 7 9 0 1 9 0 7 9 8 1 15 2
52 7 13 9 0 0 1 9 7 9 8 13 1 9 0 0 7 15 3 0 9 9 0 0 1 8 2 9 9 8 1 10 9 8 9 0 1 9 0 7 0 7 0 1 9 9 0 9 1 9 9 0 2
6 8 13 9 0 1 8
3 8 12 9
42 13 9 9 9 0 8 8 3 9 9 9 0 1 8 8 8 1 9 9 9 0 8 8 1 9 9 9 7 13 9 0 1 9 9 0 9 1 9 0 1 9 2
65 7 13 9 0 0 1 9 7 8 13 1 9 2 13 9 0 7 1 8 8 8 7 8 9 9 8 8 9 0 7 9 9 1 9 9 7 14 8 10 9 1 9 9 1 15 1 15 9 7 8 8 8 8 1 9 9 9 0 8 8 9 1 9 2 2
14 13 9 15 9 12 9 12 9 9 9 0 2 8 2
14 13 9 15 9 12 9 12 9 9 9 0 2 8 2
8 9 7 9 2 0 0 1 8
6 8 12 9 12 2 12
66 1 15 13 0 9 7 9 1 0 0 1 8 1 9 9 5 9 12 7 13 1 9 0 1 9 2 2 9 2 12 9 0 2 9 0 7 9 12 8 9 7 9 0 7 9 7 9 9 12 9 9 12 9 7 9 7 9 12 9 7 9 0 12 9 0 12
8 9 7 9 2 9 8 1 8
6 8 12 9 12 2 12
27 1 15 13 9 7 9 1 9 9 0 1 8 1 9 9 2 9 9 12 7 13 1 9 0 1 9 2
80 9 7 9 0 7 9 0 7 0 7 9 9 7 9 0 2 12 8 9 0 0 7 9 7 9 0 2 12 8 9 0 9 9 7 9 0 2 12 8 9 0 9 0 7 9 7 9 0 2 12 8 9 0 9 0 7 9 2 12 8 9 0 9 0 7 0 2 12 8 9 0 9 0 7 0 2 12 8 9 0
7 8 9 9 8 13 9 8
6 8 12 9 12 2 12
36 13 12 12 9 0 15 13 9 9 8 13 1 9 9 8 0 1 8 8 8 8 1 9 1 9 10 9 0 1 9 8 1 9 9 0 2
13 13 7 8 15 9 9 8 1 9 13 9 0 2
20 1 9 0 1 8 12 9 0 7 12 7 12 1 12 1 15 9 1 9 2
24 1 0 7 13 12 9 0 13 9 9 8 1 9 10 9 0 0 1 9 0 1 10 9 2
8 9 0 1 9 8 1 9 9
6 8 12 9 12 2 12
36 13 9 9 8 0 0 9 1 9 9 0 9 9 0 0 1 9 0 1 8 1 9 0 1 9 8 9 9 1 9 9 8 7 9 15 2
60 13 8 8 9 9 9 7 1 9 2 2 9 9 9 2 2 15 13 12 9 2 7 15 13 9 0 0 1 9 12 9 2 7 13 1 12 9 7 15 9 9 0 7 9 0 7 9 8 7 9 0 1 9 9 7 9 7 9 0 2
33 7 13 8 7 1 9 12 13 1 0 1 9 1 9 7 9 7 9 0 2 7 13 9 9 9 1 9 12 1 12 1 9 2
40 7 1 0 7 13 0 1 12 9 1 12 9 9 1 9 9 1 9 9 0 1 9 15 13 9 1 12 9 7 1 15 13 9 0 1 8 1 9 15 2
9 12 9 1 9 8 8 1 9 0
7 8 8 12 9 12 2 12
29 13 0 1 12 12 9 1 9 9 1 9 8 8 1 9 0 7 9 15 13 9 9 0 1 7 13 12 9 2
15 7 13 0 9 1 7 10 9 14 13 7 13 9 0 2
53 13 9 1 9 9 9 0 1 8 8 7 15 13 1 10 9 1 9 8 3 7 10 9 1 15 9 2 0 15 7 9 13 9 0 7 9 0 0 7 13 1 9 0 7 13 1 7 9 9 9 9 0 2
9 7 9 0 7 9 9 0 0 2
35 13 9 8 8 8 1 9 0 0 7 9 0 1 10 9 0 1 0 2 7 1 9 15 7 13 1 9 9 1 9 0 1 10 9 2
3 2 13 2
7 9 9 0 1 9 0 0
6 8 12 9 12 2 12
39 13 9 9 0 9 9 9 9 12 8 1 9 0 0 1 9 8 1 8 1 9 8 0 0 1 9 8 1 9 7 9 1 9 8 0 9 0 9 2
34 7 13 9 9 10 14 13 9 15 1 9 12 2 7 9 15 0 8 12 12 9 0 2 7 9 15 13 9 9 7 9 9 0 2
34 7 1 10 9 0 9 9 1 9 0 1 9 7 10 9 13 1 15 9 9 9 12 1 9 0 0 15 13 9 15 1 9 0 2
29 13 1 7 9 8 1 9 7 9 15 0 0 1 9 7 9 1 9 7 13 9 0 1 9 9 7 9 0 2
5 9 9 0 1 8
3 12 2 12
54 9 9 13 1 8 8 12 9 2 8 2 13 9 9 9 1 9 9 8 1 8 7 13 1 9 9 0 7 13 1 7 9 9 9 0 7 15 9 1 2 2 9 9 0 2 2 14 13 1 9 0 1 9 2
42 13 1 9 7 10 9 15 0 9 13 1 2 2 9 9 0 2 2 15 13 15 8 1 0 9 1 9 9 9 7 13 0 1 8 7 0 1 9 1 10 9 2
38 7 9 10 9 12 9 7 9 9 9 0 1 15 12 9 7 1 9 12 8 7 0 9 1 15 12 9 7 9 9 1 15 12 8 9 2 9 2
8 0 0 1 9 8 1 9 8
6 8 12 9 12 2 12
26 13 9 8 0 9 9 1 9 12 0 0 1 9 9 8 13 9 15 12 1 12 1 0 9 9 2
42 1 10 9 12 12 9 0 1 9 8 0 12 1 12 1 0 9 15 0 12 12 9 0 2 7 13 8 8 8 9 0 1 9 9 8 1 9 8 8 0 0 2
23 8 8 1 9 0 13 9 0 0 7 9 0 1 9 9 9 8 7 13 9 9 8 2
28 7 1 9 9 13 9 0 7 9 7 9 1 9 9 9 8 8 8 0 9 1 9 9 7 9 9 0 2
47 7 1 9 9 9 8 8 8 0 1 9 8 13 10 9 0 9 15 12 9 0 13 9 1 9 1 12 9 1 9 0 7 12 9 1 9 7 12 9 1 9 7 12 9 1 9 2
22 0 1 9 7 1 9 0 1 12 8 9 1 9 8 8 12 1 12 1 0 9 2
11 9 0 13 9 0 1 9 9 1 9 9
6 8 12 9 12 2 12
31 13 9 9 0 9 9 1 9 8 0 9 0 7 0 1 9 9 1 9 9 9 1 9 7 9 7 15 1 9 9 2
42 13 9 0 12 12 8 2 1 12 12 8 0 2 1 9 1 9 9 0 0 1 9 0 8 0 2 7 13 8 3 12 8 8 1 15 3 1 9 1 12 9 2
20 1 1 12 9 1 9 9 13 12 9 0 8 1 15 12 9 9 7 9 2
8 9 2 2 9 9 2 2 0
6 8 12 9 12 2 12
38 13 9 9 1 9 9 3 9 9 1 9 9 9 1 12 9 0 1 9 2 2 8 8 8 2 2 1 9 8 0 1 9 8 1 9 8 0 2
22 9 2 2 8 8 8 2 2 12 8 8 7 13 1 9 2 2 9 9 2 2 2
12 9 0 2 9 9 0 7 9 0 1 9 0
6 8 12 9 12 2 12
24 13 9 8 11 9 9 0 8 8 9 9 0 0 7 9 0 0 1 7 15 1 9 0 2
47 7 13 9 8 0 9 1 11 9 15 1 9 1 15 9 7 15 1 0 7 13 9 9 9 0 8 8 1 9 9 0 9 0 1 9 9 9 7 9 1 9 9 0 1 9 0 2
33 7 13 11 1 9 9 9 1 9 9 0 1 7 9 0 14 13 9 0 0 1 1 9 0 1 9 1 9 9 0 7 0 2
5 9 0 1 9 0
6 8 12 9 12 2 12
16 1 15 13 0 9 0 1 9 0 1 9 0 0 9 9 2
105 9 2 2 9 0 2 2 2 2 8 13 1 9 9 0 0 1 9 2 9 0 13 9 0 0 1 9 9 9 2 2 9 0 2 9 0 2 2 2 2 8 13 1 9 9 0 0 1 9 9 2 2 8 8 8 2 2 2 2 8 13 1 9 9 0 0 1 9 2 9 0 13 9 0 0 1 9 9 9 2 2 8 8 2 2 2 2 9 2 2 13 2 2 9 9 2 8 13 2 2 2 9 1 9 15
6 9 9 9 9 9 9
6 9 12 9 12 2 12
42 13 12 9 9 9 9 9 9 15 13 1 9 15 13 1 9 9 9 3 9 0 1 9 1 0 9 1 9 1 9 15 1 9 9 1 9 0 1 15 9 9 2
27 7 14 13 1 9 9 9 9 9 1 9 9 0 9 9 1 9 0 7 9 1 9 0 8 8 8 2
44 13 9 0 14 13 9 9 1 9 1 9 1 7 13 9 15 7 13 15 1 9 15 7 15 13 1 9 1 9 9 15 7 13 1 9 9 9 7 9 12 0 1 9 2
26 13 9 0 1 9 15 1 8 9 9 1 9 1 9 0 7 13 1 9 9 12 15 13 1 9 2
47 7 13 9 9 0 0 9 9 8 8 1 9 13 15 1 9 8 8 7 9 12 1 0 0 7 14 13 8 1 9 0 14 0 0 7 14 13 1 15 9 0 7 9 15 9 8 2
45 7 14 13 8 8 8 1 9 9 9 7 9 15 13 1 9 9 7 13 9 1 9 1 9 0 1 9 9 1 9 7 1 9 15 9 9 15 13 13 15 1 9 1 9 2
15 9 0 2 9 0 7 8 7 8 13 9 9 9 1 9
6 8 12 9 12 2 12
38 14 13 9 0 7 8 7 8 9 0 1 9 1 9 1 9 1 9 10 1 9 2 2 2 7 13 9 9 1 9 0 0 9 9 15 9 9 2
26 7 13 9 15 13 9 9 9 15 2 7 9 14 13 1 12 9 13 15 10 9 12 1 9 0 2
32 7 13 7 10 9 12 15 14 13 9 9 0 1 9 9 1 9 1 9 9 9 2 14 13 1 9 1 9 1 9 0 2
29 7 13 9 9 15 7 3 9 1 8 1 9 9 9 9 0 1 9 10 1 9 1 9 9 0 7 9 9 2
30 7 13 1 7 9 9 14 13 1 9 0 7 0 0 1 9 1 9 7 14 13 1 8 9 9 0 0 8 8 2
12 9 0 13 9 9 1 0 9 1 9 9 0
6 8 12 9 12 2 12
40 13 9 9 0 8 8 1 9 0 1 9 9 7 13 9 9 15 13 15 15 0 15 12 9 1 9 0 1 9 9 1 0 9 1 9 0 1 12 9 2
63 7 13 9 0 1 9 0 1 9 9 7 9 9 0 13 9 0 9 1 9 0 1 8 1 1 9 15 1 12 1 12 1 9 1 9 0 1 8 7 8 8 2 9 1 12 1 12 1 9 1 9 9 7 9 0 0 2 0 0 9 0 0 2
66 7 1 1 12 9 13 9 1 15 1 12 9 9 0 2 13 9 9 12 9 7 13 9 9 15 1 12 9 2 7 13 9 1 12 9 0 7 13 13 12 9 2 1 9 15 13 1 15 0 0 15 13 9 1 9 9 15 0 1 1 9 1 12 9 0 2
30 7 13 9 9 1 0 9 0 1 9 9 0 2 1 9 15 13 1 15 1 9 9 9 0 1 8 0 12 9 2
28 7 13 9 0 0 0 0 1 15 0 15 12 9 1 9 0 8 2 7 13 8 0 9 13 15 1 9 2
55 7 13 9 0 0 3 0 0 9 1 9 9 1 9 0 1 9 8 15 13 15 9 9 0 1 9 2 7 13 8 8 8 9 9 9 9 9 1 2 9 0 2 15 13 15 9 15 1 9 0 15 13 9 9 2
71 7 13 9 9 9 9 8 8 2 7 8 8 1 9 7 12 0 13 1 7 8 1 9 15 8 8 7 8 10 9 1 9 0 2 2 7 13 9 9 9 9 9 1 9 1 9 8 9 1 0 0 1 9 9 0 1 9 2 9 15 13 9 0 1 9 9 0 1 9 9 2
42 7 13 9 7 0 1 9 13 9 15 1 9 0 1 9 1 9 7 9 9 15 13 1 9 0 2 7 9 8 1 9 9 9 7 9 7 9 0 14 13 0 2
43 7 1 9 1 15 2 13 7 8 7 1 9 0 2 13 1 9 0 3 7 7 3 9 0 1 9 9 1 9 15 2 7 14 13 1 9 9 0 1 9 9 12 2
97 7 1 9 1 9 2 2 8 8 8 2 5 2 13 9 9 9 9 8 8 9 2 13 3 9 1 9 14 13 1 15 9 0 1 9 9 0 2 1 7 13 0 1 8 8 2 2 13 9 1 7 12 12 9 0 1 9 8 13 13 1 15 9 1 9 2 7 1 9 1 15 2 13 9 9 1 12 1 12 1 8 7 12 1 12 1 8 7 1 0 1 12 1 12 1 8 2
36 7 13 9 9 0 7 9 9 9 1 9 15 13 9 1 9 9 14 13 12 1 12 2 7 0 1 12 1 12 1 9 0 1 10 9 2
7 9 0 1 9 9 9 0
6 8 12 9 12 2 12
13 13 9 1 7 13 9 9 0 1 9 1 9 2
48 7 13 2 2 8 8 8 2 2 9 9 9 14 13 9 1 9 9 0 7 0 1 9 9 9 9 9 1 9 7 9 9 7 1 0 9 9 1 9 0 7 0 7 0 1 9 0 2
28 13 9 9 1 9 12 1 12 1 9 0 7 13 1 12 12 9 0 1 9 0 1 10 9 7 13 9 2
17 13 9 9 9 9 0 0 1 9 9 0 1 9 9 7 0 2
18 13 9 1 9 9 7 9 9 9 1 9 12 9 0 1 10 9 2
12 9 0 1 9 10 1 9 13 1 9 9 0
6 8 12 9 12 2 12
29 14 13 9 1 9 9 9 1 9 0 1 9 0 1 9 9 15 1 9 9 9 9 7 9 1 9 2 2 2
12 7 13 9 1 9 9 9 8 8 9 9 2
28 7 13 9 2 8 8 12 9 0 2 12 1 9 8 0 0 7 12 1 9 9 7 0 1 9 9 0 2
27 7 14 13 9 0 1 8 1 9 1 9 0 1 8 7 8 7 9 1 9 15 1 8 9 9 0 2
29 7 13 9 0 1 9 10 9 0 1 9 1 9 9 9 9 7 1 0 7 13 9 1 9 1 9 9 12 2
23 7 13 9 2 7 9 0 13 1 9 9 0 1 9 9 2 7 9 7 9 7 9 2
6 8 13 9 15 1 9
6 8 12 9 12 2 12
20 13 9 8 0 1 9 12 1 12 1 9 9 9 1 9 1 9 9 12 2
22 1 9 0 13 8 7 15 13 9 12 1 12 1 9 9 1 9 1 9 9 12 2
33 13 7 8 13 0 1 9 1 9 9 9 9 1 9 9 0 7 0 7 13 9 0 1 0 9 1 9 0 1 9 1 9 2
28 9 0 13 1 15 8 8 0 8 8 8 0 8 0 8 8 1 15 9 0 7 0 1 9 9 1 9 2
42 13 2 2 8 8 2 2 0 9 8 1 9 1 8 13 1 9 2 8 2 7 8 13 7 13 12 12 9 1 9 10 9 1 15 1 15 9 0 0 7 0 2
7 9 0 1 9 8 1 8
6 8 12 9 12 2 12
35 13 9 8 0 1 9 9 15 13 1 15 9 9 8 1 9 9 8 0 7 9 14 13 9 0 1 9 1 10 9 1 9 10 9 2
47 13 9 1 9 7 1 8 0 1 12 12 9 1 9 7 9 15 13 1 8 7 0 15 2 7 1 9 14 13 7 7 9 8 0 1 9 2 7 13 9 9 9 0 1 15 13 2
20 7 13 9 7 9 9 0 9 1 10 8 9 0 9 1 15 1 15 8 2
21 7 14 13 8 1 9 9 8 9 0 7 12 9 0 1 9 1 8 1 9 2
34 7 13 8 14 13 12 9 9 7 12 9 0 7 9 15 0 12 12 8 2 1 12 8 9 0 2 1 9 1 8 1 9 9 2
12 9 0 0 13 1 12 9 0 0 1 9 8
6 8 12 9 12 2 12
54 13 9 0 0 0 0 2 8 2 7 15 14 13 12 9 9 0 13 1 8 1 9 1 9 9 9 9 9 0 0 2 8 2 2 1 9 15 13 1 15 1 9 9 9 0 1 9 9 9 1 9 15 0 2
46 7 13 9 2 8 2 8 8 7 15 14 13 9 1 9 0 1 12 9 9 0 2 1 15 1 15 9 0 7 0 7 0 1 9 9 0 1 9 9 8 1 9 9 9 9 2
12 2 2 7 13 9 1 9 9 0 9 9 2
47 7 13 8 9 9 0 1 9 9 0 1 9 9 2 9 14 15 1 9 9 0 0 1 9 9 15 13 1 7 1 15 8 9 8 1 9 1 9 7 9 9 1 9 1 9 9 2
21 7 13 3 9 0 1 9 1 9 1 7 9 1 8 14 13 15 1 9 9 2
48 7 13 7 15 14 13 13 1 9 9 0 9 1 9 15 13 7 13 1 15 1 9 9 1 8 2 0 1 7 0 2 8 2 13 9 15 1 9 9 9 7 13 9 9 9 1 9 2
9 9 0 13 9 9 1 9 9 0
6 8 12 9 12 2 12
39 13 9 0 7 15 14 13 1 9 9 9 0 1 9 9 0 1 9 9 0 1 9 9 1 9 9 8 3 7 15 13 9 15 12 1 9 8 8 2
40 7 13 9 8 0 9 9 9 1 8 8 8 9 9 0 9 15 1 9 1 15 9 7 9 0 13 9 0 1 9 9 0 1 9 9 1 10 9 0 2
36 7 13 9 0 9 9 0 1 9 9 0 1 9 9 0 15 13 1 9 1 9 9 9 0 7 1 9 1 9 9 0 1 9 9 0 2
7 9 9 0 1 9 9 9
6 8 12 9 12 2 12
34 13 9 0 1 9 9 1 9 7 9 0 13 1 9 12 9 8 8 8 9 9 8 2 9 9 9 2 14 13 9 15 9 9 2
21 13 0 1 12 9 1 9 1 10 9 14 7 15 14 13 9 1 9 7 9 2
22 7 14 13 0 1 12 1 9 9 0 7 9 9 9 0 7 0 1 9 10 9 2
11 7 14 13 9 9 7 9 9 1 9 2
5 9 1 9 9 8
6 8 12 9 12 2 12
32 13 9 0 9 9 1 8 7 1 9 15 0 9 0 15 13 9 9 1 9 0 8 8 8 7 9 0 0 8 8 8 2
34 7 13 9 7 1 9 15 0 3 9 9 9 0 1 9 9 9 0 1 9 9 0 7 1 9 15 12 9 7 9 13 9 15 2
41 7 13 9 2 9 0 2 1 9 9 1 9 9 0 1 9 8 7 8 8 7 3 1 9 8 9 9 8 1 1 9 8 8 1 7 13 9 7 9 0 2
25 7 13 9 9 0 13 1 15 7 15 1 0 9 9 7 9 9 9 1 0 9 9 9 9 2
33 7 13 9 2 8 8 8 2 7 9 0 13 12 9 8 0 7 12 9 0 1 9 0 9 0 9 7 9 0 9 12 9 2
40 7 13 9 2 9 0 2 7 9 9 0 1 9 7 9 8 13 7 13 9 9 0 9 7 13 9 9 9 9 8 8 7 15 13 9 1 8 9 9 2
40 7 13 9 2 8 0 2 7 9 9 1 9 14 13 9 0 1 9 0 8 9 9 1 9 1 9 9 9 1 9 0 7 0 1 9 1 9 8 8 2
5 9 9 9 1 9
6 9 12 9 12 2 12
25 13 9 9 1 9 1 1 12 1 12 7 13 9 0 1 9 1 9 7 9 0 1 9 9 2
83 7 13 9 1 9 13 9 15 3 9 7 0 1 9 7 9 15 13 9 1 9 2 9 2 13 15 1 9 9 15 15 13 10 9 7 13 1 9 1 9 15 0 1 9 9 7 1 15 14 13 1 12 9 0 1 15 13 9 1 15 7 9 1 9 7 1 9 9 7 3 15 13 9 1 7 15 13 9 1 9 9 0 2
73 7 13 9 1 9 9 9 1 9 9 15 7 1 12 1 12 1 9 15 1 9 13 2 9 2 1 9 0 7 7 9 0 13 9 1 9 15 13 9 15 1 12 7 12 9 7 15 1 10 1 9 0 1 15 13 9 9 9 7 13 0 9 2 0 2 1 9 1 12 1 12 9 2
8 9 0 1 9 1 8 1 8
6 8 12 9 12 2 12
19 13 9 9 0 1 9 7 9 1 8 1 0 9 0 0 2 8 2 2
29 1 9 8 13 9 0 1 9 1 15 9 8 9 0 2 7 9 0 1 9 0 1 9 8 7 13 9 0 2
62 7 1 9 9 13 0 9 9 9 7 9 15 12 7 9 9 7 9 15 12 12 7 9 9 9 7 9 15 12 7 15 9 1 12 9 2 7 13 9 1 9 9 13 1 15 9 2 14 10 9 7 15 1 12 9 9 9 13 9 1 9 2
18 13 9 9 9 9 1 8 9 0 1 13 9 9 1 0 9 0 2
27 15 7 7 9 15 13 9 9 9 9 0 13 7 15 1 1 9 1 9 0 7 1 8 13 9 15 2
10 9 9 1 9 8 0 7 9 8 0
6 9 12 9 12 2 12
39 13 3 8 9 1 9 8 0 7 9 8 0 1 9 1 9 0 7 0 7 0 7 0 7 0 7 0 1 9 12 2 12 2 7 13 9 9 0 2
43 7 13 0 9 1 9 0 1 8 0 1 9 9 8 0 7 13 9 1 9 0 7 9 9 1 9 1 9 1 9 0 1 9 9 13 1 15 1 9 0 1 9 2
26 7 13 9 1 9 1 9 0 0 1 9 7 9 9 0 7 0 7 9 8 7 0 7 9 15 2
47 7 13 9 9 1 8 8 9 9 1 9 9 0 7 0 7 0 7 9 9 0 7 9 9 1 8 1 10 15 0 1 9 0 1 9 7 9 1 9 7 9 9 0 7 9 15 2
24 13 7 9 1 9 8 13 1 9 8 1 9 9 8 7 13 9 9 0 1 9 1 9 2
7 9 0 13 9 8 1 8
6 8 12 9 12 2 12
23 13 8 8 9 9 7 9 0 9 9 9 9 9 9 0 0 2 8 2 1 9 15 2
51 7 13 8 1 9 8 13 15 1 9 9 9 0 1 0 1 9 0 1 9 1 9 9 2 1 7 8 14 13 9 15 0 1 9 15 1 8 1 9 9 9 9 0 0 13 15 9 12 9 8 2
35 7 13 7 9 15 14 13 1 9 9 9 9 0 9 1 9 0 13 9 15 9 9 1 9 9 2 1 9 1 9 1 9 9 9 2
36 7 13 8 7 12 7 12 1 9 0 1 9 14 13 9 15 0 1 9 1 9 9 9 0 1 8 7 1 9 9 1 9 8 7 9 2
45 7 13 1 7 9 0 1 9 1 9 1 9 15 7 13 1 9 0 1 9 9 2 1 7 15 13 1 7 15 2 4 3 15 13 1 9 9 9 1 9 2 1 9 9 2
7 9 9 9 0 0 1 9
6 9 12 9 12 2 12
33 13 9 9 9 0 0 1 9 15 0 9 12 7 12 9 0 1 9 8 8 1 9 8 8 8 2 1 15 13 9 0 0 2
52 7 13 9 9 9 1 9 7 9 1 9 9 9 9 8 8 1 9 1 9 8 7 9 0 0 1 9 1 9 15 7 0 15 1 9 9 0 1 9 1 9 9 7 9 0 7 9 9 1 9 0 2
45 7 14 8 9 0 1 9 9 8 0 7 0 8 8 1 1 9 9 0 1 9 1 9 0 1 9 0 8 8 13 1 15 9 1 9 7 0 1 9 7 9 7 0 0 2
22 7 14 13 9 0 13 1 15 9 1 9 8 8 8 8 8 1 9 9 8 8 2
31 13 7 9 13 1 9 9 0 1 9 9 0 7 13 9 1 9 0 1 9 9 1 9 9 9 1 9 9 1 9 2
12 9 9 9 8 1 0 1 12 9 1 9 12
6 8 12 9 12 2 12
40 13 9 9 0 0 1 15 1 9 9 9 0 1 9 2 8 2 7 13 1 9 12 9 1 9 0 1 9 12 0 2 2 2 7 13 0 15 13 3 2
65 7 13 9 8 15 13 1 8 9 1 15 2 1 9 1 15 7 9 9 9 12 1 9 9 15 14 13 1 12 9 1 9 0 9 9 2 7 1 9 1 9 15 12 9 9 1 9 9 14 7 15 10 13 0 1 9 0 1 1 9 7 0 12 9 2
23 7 13 10 9 1 7 13 8 1 9 0 9 15 1 9 9 9 1 0 1 9 0 2
32 7 13 8 1 9 15 15 13 3 9 12 9 8 1 9 9 15 0 1 12 12 9 1 9 1 9 1 9 9 9 9 2
25 7 13 9 9 1 9 9 1 9 15 13 15 1 9 12 0 7 15 14 13 0 1 9 8 2
42 7 1 9 9 2 13 9 9 0 0 1 12 9 1 9 0 1 9 1 9 9 0 2 7 1 8 13 9 0 8 0 12 9 7 13 1 12 9 1 9 0 2
55 7 13 9 9 9 1 8 1 0 15 1 9 9 1 9 0 1 14 12 9 0 1 1 8 2 7 13 9 9 11 8 9 9 0 7 8 0 1 9 9 7 7 9 13 1 9 9 1 9 9 9 1 9 0 2
18 7 9 0 13 1 7 13 9 0 1 9 9 1 13 9 0 8 2
24 7 13 9 9 7 9 0 1 1 8 7 0 12 9 1 9 0 13 9 7 9 1 9 2
10 9 8 8 8 13 1 9 9 1 9
6 8 12 9 12 2 12
27 13 9 8 8 8 9 9 7 8 7 8 14 13 9 0 8 8 1 9 9 9 0 1 8 9 0 2
35 7 13 8 1 9 0 0 9 15 1 9 15 0 8 8 1 9 8 1 9 9 0 2 7 9 15 1 8 14 13 8 9 1 9 2
29 7 13 7 15 13 1 8 7 8 9 9 1 9 1 9 9 0 7 8 8 13 1 8 8 9 1 9 0 2
34 7 1 9 15 2 13 8 8 13 1 8 9 9 1 9 8 8 13 12 9 2 7 15 13 9 9 1 9 9 1 8 8 8 2
29 7 13 8 1 9 15 1 8 2 7 8 13 1 9 9 1 8 1 9 9 9 0 1 8 1 10 9 2 2
46 7 1 9 9 15 2 13 7 15 7 1 9 1 9 9 9 1 8 7 8 1 9 9 9 1 9 9 0 2 14 13 9 9 9 9 9 0 1 8 8 8 7 8 0 8 2
8 8 13 1 9 1 9 1 8
6 8 12 9 12 2 12
36 13 9 0 8 8 9 1 9 9 0 1 9 8 8 1 9 0 1 9 1 9 9 9 7 9 7 9 7 9 0 1 9 9 8 8 2
19 7 13 9 8 0 9 9 7 9 13 9 8 1 9 7 9 9 9 2
24 7 13 8 1 9 1 9 9 9 9 7 9 0 7 13 1 9 9 15 7 9 15 0 2
13 8 13 1 9 9 9 0 1 9 1 9 9 9
7 8 8 12 9 12 2 12
43 13 8 9 9 1 9 15 1 9 9 1 0 9 1 9 9 0 1 9 9 9 1 9 9 15 9 9 9 0 2 0 9 1 2 9 9 2 1 9 15 10 9 2
45 7 13 9 0 1 9 0 8 8 1 9 3 1 7 9 0 1 8 1 9 15 1 9 9 1 9 0 13 1 9 15 1 2 9 2 1 9 0 1 9 9 1 9 9 2
34 7 1 9 1 15 2 13 9 1 7 15 13 13 1 9 9 1 10 9 9 1 9 1 9 9 9 9 9 9 8 15 1 9 2
38 7 13 8 9 1 9 9 1 9 9 1 9 1 9 9 9 9 2 9 14 15 1 9 9 13 1 8 7 9 15 8 13 9 15 1 9 15 2
94 7 13 2 7 15 1 10 9 14 13 9 0 1 9 9 8 9 0 1 9 9 0 7 9 9 14 13 0 9 1 9 9 2 2 7 13 9 2 7 15 7 1 9 1 9 9 9 0 1 9 0 7 8 15 13 8 8 9 2 1 9 8 8 2 13 8 8 9 15 1 12 9 0 1 9 9 0 1 9 0 1 9 0 8 8 1 9 9 2 9 1 9 2 2
12 9 9 13 9 1 9 9 1 9 2 8 2
3 9 12 9
27 13 9 8 9 8 2 9 0 1 9 9 0 9 2 9 9 9 15 1 9 9 1 9 0 1 9 2
46 7 13 9 1 9 1 15 7 9 9 15 2 13 9 1 9 2 8 12 2 1 9 9 8 8 2 12 9 0 1 9 9 2 9 8 2 7 2 8 8 2 9 9 9 9 2
31 7 13 9 1 7 9 13 1 9 9 9 1 2 9 7 9 9 2 1 9 9 9 9 8 7 13 9 15 12 9 2
25 7 13 9 2 7 9 9 10 13 9 1 9 9 7 9 1 9 0 2 7 9 1 9 2 2
57 13 9 0 0 14 13 7 9 13 9 9 9 1 9 8 8 9 9 9 2 0 7 9 14 13 1 9 7 9 2 1 10 9 13 9 0 1 9 9 9 8 1 9 0 1 9 13 15 9 1 9 0 1 9 0 0 2
23 7 13 9 0 7 9 0 13 9 13 9 1 9 1 9 9 7 13 9 9 1 9 2
14 7 13 9 0 9 9 1 9 9 8 9 9 9 2
34 7 13 9 1 9 7 9 0 1 9 0 13 9 1 9 0 7 13 1 9 1 9 0 7 13 0 1 9 9 1 2 0 2 2
6 9 9 9 0 1 9
3 9 12 9
28 13 9 9 0 8 8 1 9 9 9 1 9 0 1 8 2 1 9 9 1 9 0 13 1 9 9 0 2
60 7 13 1 9 8 1 9 9 0 9 9 0 8 8 7 13 9 0 1 9 13 12 9 1 7 13 2 1 9 0 1 9 0 1 8 1 9 7 13 1 8 9 1 9 0 8 8 1 9 9 9 8 8 7 9 9 0 8 8 2
13 7 13 9 0 9 0 0 1 9 8 1 9 2
26 7 13 8 14 13 1 9 1 9 9 9 0 1 9 0 1 9 2 0 9 15 1 2 9 2 2
11 8 2 9 0 1 9 9 15 1 9 15
3 9 12 9
20 13 8 8 9 9 0 0 9 9 7 9 0 1 9 9 15 1 9 15 2
47 13 8 8 1 9 0 0 13 15 3 1 9 9 9 1 9 15 0 8 8 1 9 13 15 8 1 9 0 8 8 1 9 8 1 9 8 8 9 9 9 8 8 9 9 9 9 2
26 7 13 8 7 9 0 13 1 9 9 1 9 9 9 0 0 1 7 15 13 7 13 9 1 9 2
36 7 13 8 7 9 0 13 15 1 9 15 1 15 1 9 7 15 13 9 1 9 1 9 0 1 9 2 7 15 15 13 1 15 9 0 2
29 7 13 7 9 1 9 0 7 0 0 7 14 13 9 0 1 9 9 1 9 7 13 7 13 9 9 1 9 2
24 7 1 9 15 13 8 8 9 9 0 7 9 13 9 7 13 7 15 1 0 9 9 0 2
21 7 13 8 9 9 0 1 9 9 9 9 0 1 9 1 9 1 8 13 9 2
14 7 1 0 7 13 9 1 9 9 10 9 0 0 2
4 9 8 13 8
3 9 12 9
26 13 9 0 9 9 9 9 9 8 8 9 9 0 8 8 1 15 9 1 9 7 9 9 1 9 2
34 7 13 9 0 0 1 9 7 9 1 9 13 1 0 9 15 13 9 7 1 9 15 9 1 9 7 9 9 7 9 0 1 9 2
41 7 14 13 8 1 9 9 15 1 9 9 0 7 0 9 14 13 1 9 13 7 13 9 9 9 0 7 7 15 14 13 1 9 0 1 9 9 7 0 0 2
51 7 13 8 1 9 9 1 9 1 9 0 1 9 0 0 7 15 14 13 0 7 9 0 9 9 0 1 9 9 0 7 0 1 9 7 9 9 0 1 15 1 15 9 0 0 1 9 9 9 12 2
43 7 13 9 9 1 9 0 7 9 9 0 1 7 15 2 0 8 8 8 8 2 7 13 9 1 9 9 7 9 9 1 10 13 9 9 7 13 8 7 9 1 9 2
59 13 8 14 13 1 9 0 0 13 15 9 9 1 9 1 9 15 1 9 0 7 9 9 9 0 1 0 14 13 0 9 1 7 9 9 0 0 15 9 9 9 0 9 0 7 0 0 1 9 15 1 9 9 0 1 9 7 8 2
32 7 13 8 1 9 0 7 15 14 13 1 9 0 9 9 0 15 13 1 9 9 1 15 7 9 0 0 8 8 9 0 2
48 7 13 9 1 9 0 8 8 9 9 9 9 9 9 0 7 1 9 0 8 8 9 0 1 9 8 8 8 9 9 9 0 1 9 9 0 7 8 8 9 9 8 0 1 9 9 0 2
34 15 7 14 13 8 1 9 9 3 9 1 9 1 0 13 7 13 15 1 9 9 9 0 1 9 0 9 9 0 1 15 1 9 2
9 8 13 1 8 9 0 1 9 9
42 9 12 9 2 8 13 9 9 0 8 8 9 0 1 9 9 0 8 8 9 9 13 9 0 15 13 15 9 9 0 0 1 1 8 1 9 9 1 9 9 0 2
56 7 13 9 9 0 7 8 13 1 9 1 9 0 0 1 9 0 1 9 9 0 7 9 9 0 0 1 12 9 0 1 8 9 8 8 9 1 9 9 9 7 9 9 15 0 1 9 9 0 1 15 1 15 9 0 2
24 7 13 8 9 9 15 15 13 9 0 7 8 7 9 15 1 9 0 1 9 0 8 8 2
24 1 9 15 13 8 9 0 15 13 1 15 8 0 1 9 9 0 0 8 8 1 9 9 2
55 7 13 8 8 0 1 9 1 9 9 0 8 8 7 9 9 1 9 9 1 9 0 0 8 8 13 8 8 8 9 9 9 8 8 0 1 9 15 1 9 15 0 1 9 9 8 8 8 8 9 9 8 8 8 2
7 9 1 9 0 1 9 9
3 11 12 9
39 13 8 8 11 8 8 8 9 9 9 0 0 9 9 9 1 9 15 0 9 8 13 1 9 8 1 9 7 9 0 1 9 2 7 13 9 8 9 2
24 7 13 9 9 9 8 9 9 0 1 9 0 0 10 9 1 9 0 1 9 15 3 9 2
6 0 8 1 8 9 0
3 8 12 9
13 8 8 13 0 8 8 13 15 8 9 0 9 2
30 2 2 8 8 2 2 2 2 2 13 8 9 0 8 8 8 8 9 0 1 15 13 15 1 9 1 9 9 0 2
29 2 2 8 8 8 2 2 2 2 2 13 9 9 9 0 0 8 8 2 9 0 0 2 1 9 9 9 0 2
40 2 2 8 8 2 2 2 2 2 13 9 9 0 9 15 1 9 9 1 9 9 0 2 1 9 8 8 2 0 0 7 14 13 9 9 15 1 9 0 2
11 8 8 8 13 9 15 1 9 8 8 8
3 8 12 9
35 13 9 0 8 8 0 1 9 0 1 9 0 0 8 8 8 8 8 8 9 1 9 8 9 8 13 8 8 1 9 9 13 3 9 2
35 7 13 7 9 8 9 12 13 9 0 8 8 9 9 0 0 8 8 8 8 12 9 8 13 1 9 8 8 13 8 8 9 15 0 2
35 7 13 7 15 13 1 9 7 13 8 8 1 9 1 9 8 8 1 9 1 9 1 9 9 9 0 1 9 9 8 8 9 9 9 2
24 13 9 0 7 8 13 1 9 9 1 15 13 13 1 9 9 9 8 0 1 9 0 8 2
10 9 12 9 9 0 1 8 1 8 8
4 8 8 12 9
38 13 9 12 9 1 9 9 0 0 2 8 2 1 15 13 12 0 1 9 1 8 8 9 1 9 0 1 9 9 7 9 9 1 8 8 9 9 2
27 7 1 9 0 1 9 9 9 13 9 1 9 12 9 0 1 9 1 9 15 1 9 0 1 9 0 2
30 7 14 13 15 9 15 12 9 1 8 7 13 1 9 0 2 7 3 12 9 1 9 9 7 13 1 9 1 9 2
23 8 8 8 0 1 9 0 13 1 9 9 0 2 8 8 12 9 8 1 9 9 0 2
21 13 8 1 9 12 9 7 13 1 15 9 0 1 8 1 15 8 1 12 9 2
23 7 14 13 9 8 1 9 15 13 9 0 1 9 9 1 9 1 12 9 1 12 9 2
10 8 13 9 1 9 9 0 7 9 8
3 9 12 9
38 13 9 9 0 8 8 1 9 9 9 9 0 1 8 2 1 9 9 13 15 9 7 13 8 7 8 7 8 7 9 2 1 15 13 9 0 0 2
34 13 8 14 13 1 9 9 0 8 8 2 7 1 8 9 0 8 8 2 7 13 8 8 9 13 1 9 1 9 8 8 9 0 2
39 7 13 8 1 9 0 0 1 9 9 0 8 8 1 9 9 2 8 13 9 8 8 9 0 1 9 9 2 1 9 0 8 8 7 13 9 9 0 2
49 8 1 9 7 9 0 13 9 9 15 1 9 1 9 2 8 8 14 13 8 9 15 1 9 8 0 1 8 9 7 8 8 8 2 7 13 9 1 7 8 9 9 9 1 9 1 10 9 2
40 7 13 8 1 9 0 7 9 0 13 15 1 9 15 1 15 1 9 2 7 15 13 9 1 9 1 9 0 8 8 2 1 1 7 13 15 15 10 9 2
7 9 8 13 9 1 9 8
3 8 12 9
28 13 9 0 1 9 9 9 8 1 9 9 1 9 9 1 9 8 13 1 9 9 9 0 0 2 8 2 2
30 13 9 2 7 15 0 9 0 13 15 8 1 9 9 1 8 2 1 9 9 0 1 9 12 9 1 9 1 8 2
41 13 9 12 9 15 8 8 8 1 9 9 0 2 7 8 8 1 9 9 0 1 9 0 2 7 8 8 8 1 9 9 2 8 8 8 1 9 9 7 9 2
29 13 9 1 9 9 7 9 1 8 0 1 9 9 1 9 0 2 7 15 9 9 0 0 1 9 8 1 9 2
42 7 13 9 1 9 9 0 7 9 9 1 9 0 1 9 0 1 9 15 13 8 2 7 13 9 1 9 9 7 9 1 9 7 9 2 9 9 2 15 13 9 2
6 9 8 13 9 1 9
3 9 12 9
49 13 9 0 1 9 0 1 9 9 0 1 9 2 8 2 1 9 9 9 7 9 9 13 9 1 9 1 9 9 0 1 15 13 8 8 1 9 0 15 8 8 1 9 0 1 9 8 8 2
36 7 13 9 1 9 8 1 9 9 8 8 8 9 15 7 9 9 0 0 1 9 9 15 13 15 1 12 9 7 7 1 9 15 9 0 2
36 7 13 9 7 8 9 8 9 9 1 9 0 14 13 8 8 9 9 1 15 0 7 13 9 0 0 1 9 0 0 1 9 9 1 9 2
84 13 9 8 0 14 13 8 8 1 0 8 9 1 9 9 7 15 13 15 1 8 9 2 9 8 8 8 13 1 15 1 9 15 2 7 14 13 13 1 9 8 9 0 1 9 8 8 0 1 9 0 1 9 7 13 8 8 0 1 9 15 13 1 0 0 0 1 9 7 9 0 9 1 9 1 9 9 9 0 1 9 1 0 2
39 7 13 10 9 9 1 9 8 8 8 8 9 9 9 1 9 15 13 8 8 1 12 9 1 15 13 1 9 8 8 13 1 9 9 9 8 8 0 2
11 9 9 8 13 8 1 9 8 8 9 0
3 8 12 9
41 13 9 9 0 9 9 7 9 9 8 8 8 14 13 1 9 0 1 8 1 9 0 1 9 8 8 9 9 0 8 8 9 9 0 1 9 0 1 9 0 2
41 7 13 1 9 9 8 8 9 15 9 9 2 1 9 1 9 0 1 8 8 8 8 2 7 9 1 9 0 14 13 1 9 8 1 9 1 12 1 12 9 2
44 7 13 7 9 9 14 13 9 1 9 9 0 0 1 9 0 1 9 0 2 7 9 8 9 1 9 9 8 8 8 2 7 13 7 9 0 14 13 9 9 9 1 9 2
31 7 13 9 0 1 9 9 0 8 8 8 2 0 1 9 15 1 7 8 14 13 9 0 1 9 8 8 13 8 0 2
31 7 13 7 8 13 9 0 1 9 8 0 1 9 0 2 7 7 9 9 1 9 14 13 1 8 9 9 8 1 9 2
25 7 14 13 8 1 9 1 9 8 7 9 0 2 7 13 1 9 15 1 9 8 1 9 0 2
7 8 13 9 8 8 1 9
3 9 12 9
28 13 8 8 8 9 9 0 15 13 9 1 9 13 15 9 9 8 9 9 9 0 1 9 9 8 8 0 2
13 7 13 8 7 8 13 3 9 9 9 1 9 2
56 13 10 9 1 9 15 13 1 15 9 9 1 9 8 9 8 8 9 0 1 9 1 9 9 7 9 1 12 9 1 9 1 9 9 9 8 8 8 15 13 1 15 9 9 0 1 9 9 1 9 15 13 13 8 9 2
19 7 14 13 0 9 0 1 9 1 9 9 15 0 9 9 9 12 9 2
43 1 9 0 13 8 8 9 9 9 9 9 7 9 0 8 8 8 8 9 7 13 8 1 9 15 1 7 13 8 8 9 9 8 8 1 9 1 9 9 9 8 8 2
4 2 8 9 2
9 8 13 8 8 9 9 9 1 9
3 8 12 9
32 13 8 9 8 8 9 9 0 8 8 8 1 9 9 15 8 8 9 1 9 2 7 13 8 8 1 9 1 9 0 9 2
66 7 13 9 9 0 1 9 1 15 2 8 8 8 9 15 13 15 8 8 8 1 9 0 9 0 1 9 9 1 9 8 2 8 8 1 7 13 9 9 0 9 2 2 13 8 1 9 9 7 9 13 9 8 8 1 9 2 7 9 9 9 0 1 9 8 2
49 13 9 9 0 8 8 0 1 9 7 9 1 9 9 0 1 9 9 0 1 9 12 2 7 14 13 9 0 0 9 9 0 7 15 13 1 9 8 8 2 7 7 9 13 8 8 1 9 2
10 8 13 8 8 9 9 9 1 9 9
3 9 12 9
21 13 8 8 9 9 0 8 8 9 9 9 1 9 9 7 9 9 0 1 9 2
34 7 13 8 1 9 0 0 13 15 3 9 9 1 9 15 0 8 8 7 8 1 9 0 8 8 13 1 9 9 9 1 9 9 2
91 7 1 9 1 9 0 2 13 8 1 7 15 1 9 9 0 0 2 14 13 9 0 1 9 9 0 1 9 0 7 9 0 13 1 9 1 9 0 1 9 7 13 9 9 9 0 7 13 1 9 1 9 15 1 9 9 15 7 9 1 9 7 13 7 9 9 10 13 9 7 9 1 9 9 7 14 9 1 9 9 1 9 7 13 1 9 9 9 9 0 2
26 7 13 8 1 9 9 9 0 9 1 7 15 13 7 9 0 14 13 1 9 9 9 0 7 0 2
38 7 9 1 9 8 7 13 14 13 8 9 9 9 0 0 13 8 7 8 14 13 1 9 10 0 1 9 15 1 7 13 8 9 15 1 10 9 2
55 7 13 8 7 9 15 1 9 0 8 8 13 1 9 9 0 1 9 9 1 8 7 9 7 9 9 9 9 0 1 8 7 9 9 0 7 9 9 9 7 9 0 7 13 1 15 1 9 8 7 13 1 10 9 2
37 13 8 9 9 0 14 13 1 9 9 9 0 1 9 1 9 0 13 1 15 9 1 9 0 8 8 7 13 15 8 1 9 9 15 1 9 2
9 8 1 9 7 8 1 9 9 9
3 9 12 9
37 13 9 9 0 0 8 9 0 1 9 8 8 3 9 9 7 13 9 1 9 9 0 1 9 9 15 13 15 9 0 1 9 9 9 0 0 2
44 7 13 8 1 9 0 13 1 15 1 8 9 15 1 8 7 9 15 13 1 9 15 13 15 9 1 9 1 8 9 1 15 13 1 9 9 9 1 9 8 8 9 9 2
17 7 13 9 1 9 8 1 9 9 9 0 1 9 9 10 9 2
68 7 1 9 0 13 9 0 7 15 13 9 15 7 9 9 13 9 1 9 9 1 9 7 14 13 3 9 9 13 1 9 7 15 9 1 9 1 9 9 0 1 9 9 1 12 9 13 1 9 1 15 9 9 0 1 9 9 7 9 1 9 9 0 7 8 7 8 2
54 7 13 7 9 9 0 0 0 14 13 1 9 9 1 9 0 1 7 10 9 15 8 8 9 8 7 14 8 13 1 9 9 0 7 9 9 0 8 15 9 13 9 9 15 7 14 13 9 15 1 9 9 0 2
48 13 9 0 1 9 8 8 14 13 3 1 9 0 9 1 9 15 1 0 8 1 9 9 15 1 9 9 1 9 9 9 9 0 8 8 9 9 1 9 7 9 7 9 9 0 9 12 2
10 9 13 1 9 9 0 1 9 9 0
3 9 12 9
19 13 8 9 9 9 0 7 9 15 13 1 9 9 0 1 9 9 0 2
48 13 9 1 9 0 0 13 15 3 9 9 1 9 15 0 8 8 7 9 13 1 9 9 0 1 9 7 15 9 1 9 7 9 7 3 9 1 9 9 1 15 1 15 0 9 7 9 2
46 7 13 9 1 7 15 4 3 9 0 7 9 1 9 0 7 13 9 9 0 0 1 7 9 14 13 7 13 14 1 9 9 7 7 9 14 13 9 15 14 1 9 9 7 9 2
19 7 13 9 0 1 9 1 10 1 9 7 9 7 9 7 0 7 9 2
27 7 13 1 9 9 9 0 0 7 9 13 9 15 1 9 10 2 7 13 9 1 8 7 9 13 9 2
29 15 7 14 13 9 9 0 9 1 9 9 0 1 9 15 1 9 9 15 15 13 8 7 8 7 8 7 9 2
10 9 0 1 8 8 13 9 0 1 8
4 8 8 12 9
42 13 8 8 8 9 0 1 9 8 8 0 0 9 1 9 9 1 9 0 7 9 9 0 7 9 9 0 0 1 9 9 9 0 1 9 9 0 0 2 8 2 2
23 7 13 8 9 9 1 9 0 1 9 9 9 1 9 9 9 1 9 1 9 1 9 2
46 7 13 9 1 9 9 7 15 8 3 1 9 0 1 0 9 0 2 8 8 7 8 8 8 8 8 0 9 2 2 7 1 9 1 9 9 13 8 1 9 9 8 9 9 9 2
17 7 13 8 1 15 1 8 9 8 8 9 9 9 8 8 9 2
36 7 13 9 8 1 9 0 9 9 1 9 9 9 0 8 1 0 9 1 1 15 9 0 8 8 9 1 9 8 8 8 8 8 1 9 2
25 7 13 1 9 9 9 9 1 9 9 1 9 8 8 9 0 8 8 1 9 15 7 1 9 2
60 7 13 8 7 2 8 8 0 8 15 9 9 9 9 0 1 8 1 12 2 7 14 8 7 8 0 1 9 7 9 1 9 0 0 1 9 2 2 7 13 7 15 13 7 13 9 9 0 7 1 8 8 7 13 9 9 9 9 0 2
7 9 0 1 15 1 8 8
3 8 12 9
50 13 9 0 8 8 8 1 8 8 8 8 9 7 9 0 1 15 1 9 1 8 15 13 1 9 9 9 0 14 13 8 8 1 8 9 9 8 1 9 9 1 9 15 13 9 1 15 1 15 2
20 7 13 9 9 8 0 1 15 9 15 2 7 15 13 8 8 1 8 2 2
26 9 7 15 13 7 15 1 1 0 1 15 14 12 2 7 7 9 8 9 15 15 15 13 1 9 2
19 1 0 7 8 15 9 0 1 9 2 7 14 13 8 8 1 12 9 2
18 7 13 2 8 8 9 1 7 8 8 14 13 1 9 9 0 2 2
27 7 13 8 7 9 8 8 8 1 10 9 14 13 8 8 1 8 7 13 1 0 1 15 8 9 9 2
34 13 7 9 0 15 13 1 9 0 1 9 1 9 8 13 1 9 10 14 13 1 12 9 8 8 1 9 0 8 8 1 12 0 2
14 9 9 0 1 9 1 9 0 1 9 0 12 2 12
61 9 9 0 1 9 1 9 0 1 9 0 12 2 12 9 12 9 2 8 2 13 9 9 0 1 9 1 9 0 1 9 0 12 2 12 1 9 0 1 12 12 9 0 1 9 0 1 9 9 7 13 9 0 0 1 9 0 0 9 9 2
27 7 13 9 9 9 9 9 0 0 1 9 0 15 13 15 9 0 7 8 7 3 9 0 15 13 9 2
72 7 13 1 7 15 1 9 9 15 13 9 9 0 1 9 1 8 7 8 7 8 8 8 7 8 7 8 1 9 0 8 8 8 13 1 9 0 1 9 0 13 9 9 0 1 9 0 1 12 12 9 7 13 9 0 12 12 9 3 1 1 13 9 9 0 1 9 1 9 7 9 2
45 7 13 9 7 9 9 0 7 0 1 9 1 10 9 14 13 7 13 9 9 0 12 12 9 1 12 12 9 1 9 0 7 13 9 9 0 1 12 12 9 1 12 12 9 2
54 7 13 9 0 9 9 14 13 1 9 13 15 9 9 0 1 9 9 1 9 9 1 7 0 9 13 9 0 1 9 7 13 9 9 9 1 1 9 1 9 9 7 9 9 1 9 0 1 9 9 1 9 9 2
34 13 7 9 1 9 0 13 13 0 0 1 9 0 1 9 9 0 7 13 13 0 1 12 9 0 1 9 0 1 9 0 7 0 2
7 9 9 9 8 13 1 8
3 8 12 9
47 13 8 8 8 9 9 0 7 9 0 9 7 15 1 0 7 13 9 9 9 9 9 9 9 8 2 8 2 1 8 1 9 8 8 9 8 9 0 8 8 9 1 8 1 9 9 2
25 7 13 9 7 15 1 0 7 13 9 8 9 0 1 9 12 9 8 8 9 9 9 1 0 2
30 7 13 9 8 1 7 15 14 13 9 9 1 9 1 9 1 8 0 9 8 8 1 9 1 12 1 12 9 8 2
59 7 13 9 9 8 0 7 9 1 9 1 8 9 0 2 14 13 9 9 0 8 8 8 9 7 9 1 15 2 7 9 9 2 7 9 7 9 0 2 7 9 0 2 7 9 1 9 9 0 2 7 9 8 1 12 1 9 15 2
58 7 13 9 7 15 1 0 7 13 9 7 9 7 8 0 2 9 1 8 2 1 9 15 14 13 1 15 9 8 8 13 12 9 8 8 9 1 9 9 8 0 1 9 2 7 9 0 1 9 2 7 9 9 0 1 8 0 2
45 7 14 13 9 0 12 1 9 9 9 8 2 15 13 9 1 9 0 12 15 13 1 8 8 9 12 7 12 9 1 9 0 2 9 8 8 9 9 9 12 7 12 9 8 2
11 8 1 9 1 9 9 9 8 1 9 0
3 8 12 9
32 13 9 9 9 9 0 8 8 8 7 15 13 9 9 1 9 1 9 9 9 9 0 0 2 8 2 1 9 0 1 9 2
31 13 8 2 7 15 3 9 9 0 1 9 0 1 9 0 0 2 1 15 1 9 9 1 9 0 1 9 8 9 9 2
16 7 13 8 9 0 1 9 9 0 1 9 9 8 1 9 2
23 7 13 8 7 9 0 9 9 15 9 9 15 13 1 9 1 9 1 9 1 9 15 2
41 7 13 9 9 9 9 7 15 1 9 8 13 7 13 10 9 1 9 15 7 9 15 1 9 15 7 9 15 1 9 0 2 7 7 13 1 9 1 9 0 2
28 1 9 0 13 1 0 0 7 9 0 15 13 9 1 9 9 9 0 1 9 10 9 1 9 15 1 9 2
25 7 13 8 7 15 13 1 9 15 13 9 1 9 9 9 9 8 8 8 8 8 1 9 0 2
18 7 13 7 9 15 13 1 8 13 7 13 1 0 1 9 9 15 2
33 7 13 7 15 13 1 9 9 7 9 9 9 9 9 15 15 13 1 9 0 1 8 7 9 1 9 9 8 7 9 1 15 2
19 7 13 8 9 0 1 9 1 9 9 9 0 1 9 1 9 9 9 2
33 7 13 1 8 8 0 8 8 8 8 0 2 7 9 8 8 8 2 8 8 8 8 1 9 2 7 9 1 9 8 8 8 0
9 9 2 9 9 9 7 9 13 0
3 9 12 9
31 13 9 0 7 0 8 8 8 1 9 9 9 8 8 7 9 9 0 0 8 8 2 9 1 15 13 8 8 9 9 2
16 7 13 8 1 8 0 1 9 7 9 1 0 9 15 0 2
36 7 14 13 9 8 2 8 2 0 3 8 8 8 2 9 0 1 9 9 9 0 1 9 1 7 13 8 9 15 9 0 2 9 1 9 2
26 7 1 9 14 12 0 1 9 9 0 1 9 12 2 14 13 14 9 0 1 8 7 9 0 0 2
39 7 13 9 2 15 14 4 13 9 0 8 8 1 9 1 15 2 1 9 9 9 0 8 1 9 8 9 8 8 8 8 8 9 15 8 8 9 9 2
30 7 13 8 1 9 0 14 13 15 9 15 7 9 0 1 9 0 0 8 8 13 8 8 10 9 1 9 1 9 2
12 9 9 13 1 9 15 8 8 9 1 9 9
3 8 12 9
37 13 9 8 7 9 7 8 7 8 1 9 15 8 8 9 9 1 9 9 15 13 1 9 12 9 1 9 0 13 1 9 15 7 13 9 9 2
29 13 9 0 8 8 7 9 9 0 8 8 1 9 9 1 9 0 8 8 8 7 9 9 0 0 8 8 8 2
22 7 13 9 0 8 8 7 9 0 8 8 9 8 1 9 8 8 8 1 9 9 2
29 7 1 9 15 13 9 1 9 15 8 8 8 8 0 2 7 13 8 8 8 1 1 9 9 8 8 9 9 2
27 13 12 9 1 8 8 9 12 0 1 9 0 14 13 1 9 1 9 1 9 8 1 9 9 8 0 2
8 9 9 0 13 1 9 9 0
3 8 12 9
27 13 9 9 0 8 8 8 8 8 0 0 8 8 9 2 7 13 1 9 15 1 9 9 0 1 9 2
35 13 8 8 1 9 1 8 7 13 1 9 1 15 7 13 8 12 0 2 9 1 15 13 8 8 8 1 9 9 9 1 9 9 3 2
35 7 13 9 9 0 8 8 8 14 13 9 9 7 8 14 13 8 8 8 1 8 8 2 7 7 9 9 9 0 2 1 9 8 2 2
25 7 13 1 9 1 8 8 7 9 9 9 8 8 9 8 8 13 9 0 1 8 1 9 9 2
48 7 14 13 9 9 15 13 9 8 1 8 1 0 8 8 9 8 8 2 8 2 8 2 8 1 9 0 1 8 0 1 8 7 8 9 9 2 7 13 9 9 8 8 8 1 8 8 2
15 7 13 8 0 7 8 13 1 9 15 0 8 8 8 2
27 7 13 8 1 9 9 0 8 8 2 7 9 9 0 8 8 1 9 0 1 9 8 1 9 3 9 2
10 9 12 1 9 9 9 1 9 9 8
3 8 12 9
37 13 9 0 0 9 7 12 9 2 1 1 15 12 1 9 9 2 13 1 9 9 1 9 0 1 9 8 2 8 0 1 9 8 9 9 8 2
22 7 13 9 7 9 0 13 0 1 12 12 8 2 1 12 9 0 2 7 13 0 2
54 13 9 1 9 9 1 9 0 13 13 9 9 1 9 0 8 2 7 13 9 1 7 13 9 9 15 13 13 1 9 15 2 7 1 15 13 9 9 7 13 1 7 13 3 1 9 12 15 13 1 9 9 9 2
24 7 13 9 9 0 9 9 2 7 13 1 9 1 7 15 13 9 1 9 1 9 1 9 2
59 0 1 9 7 9 9 13 1 0 9 0 9 1 9 7 13 12 12 9 2 1 9 9 9 0 1 9 1 9 0 2 7 10 9 13 9 0 1 9 9 1 9 7 9 9 1 9 9 7 9 9 1 9 9 1 9 15 9 2
39 7 1 9 9 9 0 1 9 0 13 8 2 9 9 1 9 2 1 0 9 12 1 9 9 2 7 15 13 1 9 12 9 0 7 9 12 1 15 2
7 8 7 8 13 0 9 9
3 9 12 9
35 13 9 0 8 8 9 0 9 9 1 9 0 8 8 7 13 9 9 9 0 8 8 9 9 1 9 7 9 7 9 9 0 9 12 2
56 7 13 9 9 9 8 0 7 15 13 1 9 2 9 9 9 1 9 9 9 1 9 7 9 8 8 8 13 8 8 9 9 15 13 15 9 0 1 9 9 9 0 1 9 9 9 1 15 13 8 7 9 1 9 2 2
25 7 13 1 2 7 8 13 1 9 15 1 9 8 8 8 1 9 9 9 1 9 9 0 2 2
20 7 13 9 7 9 2 13 3 9 9 1 9 7 9 0 1 10 9 2 2
11 8 12 9 1 9 1 8 1 9 9 9
3 8 12 9
32 13 12 9 8 8 1 9 13 1 9 9 1 9 8 1 9 8 1 9 8 9 9 9 1 0 8 8 1 8 3 9 2
12 13 9 1 8 8 8 7 13 13 9 12 2
9 7 14 13 9 0 1 9 9 2
10 9 9 8 8 0 1 8 1 9 0
3 8 12 9
16 13 9 0 8 8 0 1 9 0 1 9 8 9 1 8 2
38 13 9 8 2 8 8 2 8 8 2 7 9 2 8 8 9 2 8 8 0 1 9 0 1 9 0 8 1 9 1 9 1 9 9 1 9 0 2
45 13 9 8 0 2 7 13 9 8 2 0 9 8 1 9 2 1 9 12 12 9 1 8 1 9 9 9 1 9 8 9 1 9 12 1 12 9 1 9 9 15 1 9 0 2
51 7 1 9 9 9 1 9 8 2 13 9 8 0 1 9 8 9 1 9 0 2 7 9 1 0 1 9 9 2 13 9 0 12 12 1 9 0 7 12 12 9 8 7 12 12 9 8 8 1 8 2
21 7 1 9 2 13 9 0 1 8 1 8 8 8 9 1 9 9 9 1 9 2
10 8 8 8 13 1 9 0 1 9 0
3 9 12 9
44 13 9 9 9 8 8 8 9 8 1 9 0 1 9 0 1 8 1 9 1 9 0 1 9 9 9 9 0 8 8 2 9 1 15 13 1 9 1 9 9 9 9 9 2
62 7 1 9 15 1 8 1 9 1 12 1 12 9 9 12 2 13 8 1 9 0 8 8 8 7 9 9 0 8 8 8 8 8 0 8 8 7 9 9 8 8 7 9 9 8 8 7 9 9 8 8 8 8 0 0 8 8 2 9 1 9 2
33 7 13 9 1 7 8 7 8 14 13 8 1 8 8 1 9 0 1 12 9 7 13 8 9 0 1 9 9 8 8 9 0 2
17 7 13 9 7 8 14 13 1 8 8 8 9 9 0 0 8 2
22 7 1 9 15 0 1 8 2 13 8 9 0 1 9 15 1 9 1 12 9 12 2
8 9 13 1 9 9 1 9 15
3 9 12 9
25 13 9 0 9 8 9 9 7 9 9 0 1 9 15 14 13 9 7 9 9 7 9 8 8 2
41 7 1 8 0 1 9 9 8 8 8 8 1 9 9 0 1 9 2 13 8 1 9 9 9 1 9 9 0 1 9 2 9 1 15 13 9 9 8 0 8 2
17 7 13 0 9 9 0 1 9 9 1 1 9 7 9 7 9 2
39 7 13 7 2 9 9 0 8 1 9 14 13 1 15 0 1 9 2 7 7 9 13 7 9 9 1 9 13 7 13 1 9 9 0 8 7 0 2 2
19 7 13 8 7 15 2 13 9 8 1 1 9 9 9 0 8 8 2 2
31 7 1 9 1 9 0 8 1 9 2 13 7 9 8 1 9 0 0 8 8 1 9 13 9 1 10 9 0 1 9 2
16 7 13 9 0 1 9 9 7 9 1 9 9 8 8 8 2
16 7 13 8 8 9 9 15 13 7 13 8 8 0 1 9 2
21 7 13 8 1 7 2 9 0 14 8 15 14 8 9 0 9 9 15 0 2 2
11 12 9 1 9 8 13 1 9 1 9 8
3 8 12 9
40 13 12 9 1 9 9 8 15 8 8 8 2 8 8 2 8 8 8 2 8 8 8 1 9 9 1 9 9 0 1 9 9 13 9 0 0 2 8 2 2
24 13 10 9 1 9 9 1 15 1 9 1 9 0 1 9 8 1 9 1 9 9 9 8 2
37 7 14 13 9 1 9 15 1 9 0 2 7 13 9 15 9 1 9 9 1 9 1 9 9 1 8 7 9 15 0 1 9 0 1 9 0 2
34 7 14 13 9 12 1 9 0 1 9 0 1 9 1 9 1 9 0 1 1 9 2 7 9 9 9 0 7 9 1 9 9 8 2
8 8 9 8 9 0 1 9 8
3 9 12 9
38 13 9 9 9 9 9 0 9 0 9 9 1 9 0 8 8 13 1 15 9 9 0 0 1 9 9 9 1 9 0 1 9 1 9 9 1 9 2
46 7 13 9 9 0 7 9 8 13 1 9 1 9 9 0 1 9 1 9 9 0 8 8 9 9 9 1 9 15 13 1 9 9 7 15 13 9 15 1 9 0 8 8 8 8 2
34 7 13 9 9 9 7 9 8 1 9 1 9 8 8 0 8 8 8 9 1 9 9 0 8 8 9 0 8 8 9 9 1 9 2
8 8 13 9 9 1 9 9 0
3 8 12 9
40 13 8 2 9 8 9 9 0 9 1 9 8 8 8 9 0 8 2 9 2 1 9 9 0 1 9 9 9 15 1 9 9 0 1 9 7 9 1 8 2
28 7 13 9 9 8 0 7 15 13 9 1 10 9 7 13 8 8 8 1 9 9 1 9 9 1 9 15 2
41 7 13 9 9 7 9 8 1 9 9 0 8 8 8 9 9 0 0 1 9 1 9 9 9 0 1 9 15 7 1 1 15 9 0 2 7 9 9 0 0 2
39 7 13 9 1 9 0 1 9 9 0 1 9 8 1 9 1 9 0 1 9 2 7 13 9 0 1 9 9 9 1 9 0 7 0 1 9 9 0 2
7 9 9 9 1 8 9 0
3 8 12 9
23 14 13 9 0 8 8 1 9 8 1 9 9 0 1 9 9 0 1 9 9 12 9 2
19 13 9 9 1 9 8 8 9 1 9 8 8 1 12 12 9 8 8 2
20 1 9 0 13 9 9 9 9 1 9 1 9 1 1 9 7 9 7 9 2
28 13 8 8 1 9 15 13 9 15 1 9 8 1 9 8 2 7 13 9 7 9 9 1 9 7 9 9 2
25 7 1 9 1 9 9 15 14 13 1 15 9 9 2 7 7 9 15 14 13 15 1 9 9 2
8 9 9 0 0 8 8 9 9
3 8 12 9
34 13 9 1 9 0 9 9 9 1 9 0 0 1 9 9 9 9 0 1 9 0 15 13 9 7 13 9 0 1 9 9 0 9 2
31 13 9 9 9 1 9 13 1 9 9 0 0 7 13 2 9 2 0 0 9 9 9 0 8 8 9 9 0 1 9 2
16 13 8 1 9 8 8 0 1 9 8 8 8 1 8 9 2
40 13 8 0 1 9 9 0 14 13 1 9 0 0 7 9 0 0 1 9 12 1 9 9 0 1 9 15 0 8 8 8 1 8 9 9 8 9 1 8 2
15 7 1 9 0 13 9 0 1 9 9 9 1 9 9 2
14 7 13 1 9 0 8 8 8 8 1 9 15 9 2
26 7 13 1 15 8 8 1 9 15 1 9 8 8 7 15 13 1 9 3 1 9 8 8 1 9 2
70 7 13 9 9 0 1 9 0 9 9 9 2 1 8 9 8 9 0 1 9 0 1 9 8 0 8 8 12 8 8 9 9 9 0 1 9 9 0 1 9 0 2 2 7 13 9 0 2 7 9 13 1 9 9 9 9 1 9 0 15 13 8 8 8 8 1 9 0 2 2
11 9 13 9 9 0 1 7 15 9 1 0
3 9 12 9
47 13 9 9 9 1 11 8 9 9 9 9 1 9 13 1 9 9 1 8 9 15 7 9 9 0 0 1 9 9 0 1 9 12 1 9 15 1 9 9 1 9 9 13 9 1 0 2
58 7 13 1 9 7 9 13 7 9 13 1 9 0 1 9 9 1 9 12 9 9 12 0 1 7 9 1 10 9 13 9 0 1 9 1 9 0 0 7 9 0 1 9 9 9 7 9 9 1 0 0 1 9 15 1 9 0 2
21 7 13 9 7 9 13 1 9 0 0 1 9 9 0 0 1 9 1 9 12 2
30 7 13 9 0 1 9 15 7 15 13 15 9 1 9 13 0 1 9 9 3 1 9 15 1 9 9 0 1 9 2
34 7 13 7 9 10 9 0 13 7 9 13 9 1 9 0 1 9 0 1 9 9 0 1 9 7 9 7 9 1 9 7 9 0 2
16 9 9 0 13 9 9 0 1 9 1 8 9 12 7 12 9
58 9 9 0 13 9 9 0 1 9 1 8 9 12 7 12 9 8 12 9 2 8 2 13 9 9 0 8 8 8 8 9 7 9 0 14 13 1 8 9 12 7 12 9 1 9 15 13 1 9 1 9 0 1 9 9 1 9 2
39 13 9 1 9 9 9 0 1 9 9 9 9 0 13 1 9 8 0 2 7 14 13 9 9 9 0 9 9 0 9 9 1 9 8 0 1 9 8 2
40 7 13 2 7 15 13 1 9 1 9 0 2 7 13 7 15 14 13 1 12 7 12 9 2 2 7 13 7 9 0 0 13 1 9 0 15 13 9 0 2
30 7 13 1 7 9 9 1 9 1 9 9 1 9 9 9 1 10 9 14 13 0 9 9 15 14 13 15 1 9 2
78 7 13 9 9 0 8 8 7 15 14 13 9 9 0 1 9 7 7 2 9 13 3 2 1 9 9 0 2 7 7 9 9 9 0 13 0 2 2 1 9 15 13 9 9 0 8 8 8 7 9 15 8 0 1 9 15 1 7 15 13 9 9 0 1 0 9 0 1 9 9 9 9 15 14 13 1 9 2
52 7 13 9 9 0 8 8 1 9 0 1 9 9 9 1 9 1 8 7 15 1 9 9 9 0 1 8 2 14 15 1 9 1 9 7 13 1 9 15 7 9 15 2 9 7 9 2 14 13 9 2 2
35 1 9 0 13 9 9 0 7 9 9 9 9 9 0 1 9 15 0 8 8 7 9 8 1 9 9 1 9 14 13 1 9 9 8 2
27 13 8 7 15 13 1 9 1 9 0 15 13 2 7 8 1 15 9 0 1 9 1 7 13 9 2 2
7 9 9 0 8 12 1 9
3 8 12 9
25 13 12 0 1 9 9 0 13 7 1 8 1 9 8 8 8 8 8 1 9 0 1 8 9 2
39 7 13 9 9 8 8 8 7 9 13 9 0 8 9 13 13 1 9 1 9 8 7 7 15 13 9 7 13 1 9 7 13 12 1 9 1 9 9 2
21 7 13 9 1 9 0 9 15 7 9 0 8 8 1 0 13 1 7 15 0 2
25 7 14 13 9 8 8 9 1 0 15 1 9 7 13 9 0 7 13 1 9 9 0 1 9 2
10 14 13 8 9 1 8 8 1 9 2
12 9 9 0 2 9 8 1 8 2 9 0 2
3 9 12 9
23 13 9 9 0 9 8 9 9 9 0 8 8 1 8 9 1 7 15 2 9 0 2 2
55 7 13 8 1 9 0 13 15 3 9 9 2 7 9 8 1 8 13 1 9 9 15 9 0 7 13 9 0 8 8 0 9 14 13 9 9 0 7 7 9 13 8 8 1 9 0 8 8 13 1 9 8 8 2 2
39 7 13 8 2 7 9 8 0 1 9 9 0 14 13 1 15 2 1 1 9 0 2 9 1 9 9 8 1 9 8 8 9 15 13 9 9 9 2 2
29 7 13 8 1 2 7 9 9 13 1 9 9 7 13 1 9 9 9 0 7 7 13 1 9 9 0 0 2 2
52 7 1 9 0 13 8 7 9 9 0 0 1 9 8 8 15 13 9 0 13 1 15 1 9 15 1 15 9 9 15 1 9 0 7 0 7 7 13 1 9 9 1 9 9 0 1 9 9 0 0 0 2
33 7 13 8 1 9 9 0 7 0 1 9 1 0 9 0 8 8 9 0 1 7 13 8 8 1 9 15 7 1 9 15 0 2
49 7 13 8 2 7 9 9 0 13 9 10 9 1 0 9 0 2 7 0 9 7 3 9 0 1 9 9 13 9 9 9 15 7 1 15 7 15 8 1 9 9 0 0 1 0 9 0 2 2
12 8 13 1 12 9 1 9 0 1 9 12 0
42 8 13 1 12 9 1 9 0 1 9 12 0 8 12 9 2 8 2 13 8 9 1 12 9 1 9 0 1 9 0 13 12 12 9 1 9 12 0 1 9 0 2
28 13 9 9 0 9 7 15 1 9 0 13 8 1 12 9 0 1 9 0 1 12 12 9 1 9 9 15 2
36 7 14 13 9 9 0 9 1 9 7 9 0 0 9 2 1 9 7 9 9 7 9 0 15 12 9 3 1 9 0 0 13 12 12 9 2
34 7 13 9 0 1 12 12 8 8 2 1 12 12 9 2 1 9 9 0 1 9 9 1 9 12 0 1 9 13 12 1 12 0 2
10 9 9 9 0 13 1 9 9 8 8
3 8 12 9
34 13 9 9 9 9 0 14 12 0 1 9 8 1 8 8 9 9 1 9 9 9 0 1 9 9 9 0 1 9 9 1 9 0 2
54 7 13 9 9 9 7 9 9 9 9 9 0 8 8 7 9 13 9 15 1 9 0 1 9 0 8 8 1 9 9 9 9 1 9 15 1 9 9 0 1 9 1 9 9 15 1 9 1 9 8 1 9 0 2
101 7 13 8 7 15 2 1 9 1 7 9 0 13 8 8 0 14 7 3 9 0 2 8 8 8 9 9 9 9 1 9 1 9 9 7 9 0 0 2 7 9 15 8 8 1 9 0 2 8 8 9 0 2 7 9 10 1 9 2 8 8 1 9 1 8 9 0 1 9 0 2 8 8 8 8 0 2 7 15 8 8 9 8 8 1 9 0 1 9 15 1 9 9 2 8 8 1 9 0 2 2
42 7 1 9 1 9 7 9 9 9 1 9 0 1 9 0 8 8 2 13 8 1 9 13 8 8 9 0 2 8 8 0 1 9 9 2 8 8 8 1 10 9 2
23 7 1 9 8 9 0 8 13 8 9 0 8 8 1 8 8 1 9 8 0 1 9 2
36 7 13 7 15 2 1 0 7 15 8 8 9 7 9 2 7 9 8 8 2 14 13 0 1 15 7 15 13 8 9 1 8 7 8 2 2
25 7 13 8 0 1 9 9 2 7 13 1 2 8 8 9 9 1 15 13 1 15 1 9 2 2
9 13 9 0 1 9 9 0 1 9
3 8 12 9
26 13 9 9 0 1 9 9 8 0 1 9 9 0 1 9 1 9 9 0 1 9 8 8 1 9 2
41 13 9 9 1 8 8 8 9 9 0 1 9 0 13 15 1 9 9 15 8 1 9 9 15 7 7 9 8 8 1 9 1 9 9 0 0 1 9 1 9 2
17 13 9 8 8 0 7 9 1 9 7 13 9 13 0 1 9 2
30 13 9 8 8 8 1 9 8 13 1 15 7 9 9 9 8 1 9 13 7 13 15 0 1 9 2 9 0 2 2
26 13 9 8 8 9 0 1 9 9 9 1 9 9 1 9 15 7 13 9 9 0 1 8 8 0 2
48 1 9 0 2 13 9 8 0 9 7 9 9 1 8 1 9 13 7 13 9 0 1 9 8 8 7 13 1 9 0 7 13 8 8 9 8 8 1 9 1 9 1 9 0 1 0 9 2
35 7 1 9 1 9 13 8 2 8 2 8 2 8 9 9 8 7 15 7 13 8 1 9 8 13 1 9 7 13 9 1 9 1 9 2
27 13 9 14 13 9 8 1 9 1 9 9 0 8 8 1 9 0 7 13 9 1 9 7 13 1 9 2
7 8 13 8 1 9 9 0
3 8 12 9
27 13 8 8 8 9 9 0 8 7 2 9 0 2 8 1 9 9 9 1 8 8 1 8 7 9 8 2
57 7 13 8 8 8 1 9 9 8 0 1 9 9 3 1 7 15 1 9 1 8 9 0 1 9 15 0 8 8 8 8 1 9 1 9 1 9 15 13 8 8 1 15 0 7 9 0 8 2 1 9 0 1 8 8 2 2
60 7 13 8 0 1 9 2 15 13 1 15 1 7 9 14 13 1 9 9 1 9 9 1 9 2 1 9 8 1 9 9 0 7 15 9 0 1 9 1 9 9 2 9 0 1 9 2 1 9 7 9 2 9 0 1 9 2 1 9 2
29 7 1 9 9 8 8 1 8 13 8 1 9 15 7 13 9 2 1 9 0 2 1 9 15 1 9 3 9 2
29 13 8 14 13 1 9 7 9 15 13 8 8 8 1 9 8 8 8 8 9 0 1 9 1 9 9 1 9 2
26 7 13 8 9 1 9 7 15 2 1 0 9 7 15 1 9 9 0 13 7 13 3 9 0 2 2
31 7 13 8 7 8 1 9 15 13 1 9 15 3 15 13 1 15 7 9 13 9 1 9 1 8 9 13 1 9 0 2
15 7 13 8 7 8 13 9 8 15 13 1 8 2 8 2
12 8 2 8 9 0 0 1 9 1 9 8 2
27 7 13 8 7 9 8 2 1 9 15 9 1 9 0 1 9 8 1 9 15 1 9 9 9 8 2 2
10 8 2 9 1 9 9 2 9 9 2
3 8 12 9
37 1 9 9 1 9 1 9 9 9 0 1 9 13 9 0 8 8 2 8 9 7 8 9 0 1 9 9 0 0 15 15 14 2 9 9 2 2
125 13 8 1 9 0 0 1 8 8 9 9 0 8 1 9 15 0 1 8 8 8 8 7 2 2 9 0 2 8 8 13 1 15 9 9 0 2 2 7 13 7 2 9 1 9 9 8 7 1 15 8 8 8 8 8 9 9 2 2 7 13 8 8 8 9 0 1 9 15 13 9 7 15 13 15 9 8 8 9 0 8 8 9 2 7 13 8 2 15 15 14 9 9 8 8 7 8 1 15 2 2 7 13 8 14 13 9 9 1 9 7 9 9 9 0 7 13 10 9 8 8 1 9 9 2
12 9 0 2 9 13 1 9 7 13 15 8 8
3 9 12 9
29 13 9 9 9 1 9 0 9 7 13 9 9 0 8 8 8 1 9 0 1 9 13 1 7 15 8 8 8 2
50 7 13 9 0 1 9 9 8 1 9 9 9 0 0 8 8 15 13 9 0 0 1 9 12 9 1 9 7 8 8 1 9 9 12 7 15 13 1 9 9 9 9 1 9 0 7 0 9 12 2
51 7 13 9 7 10 9 1 15 8 0 1 9 15 13 1 9 0 8 8 13 1 15 9 8 8 8 9 1 8 7 9 1 10 9 7 13 9 8 8 1 9 9 1 9 1 9 9 0 1 0 2
35 7 13 9 9 1 7 15 13 0 8 8 8 8 7 13 9 1 9 9 7 9 9 1 10 13 9 9 7 13 8 7 9 1 9 2
54 7 13 8 14 13 1 9 15 10 1 9 1 9 9 0 1 9 9 0 13 1 15 1 7 15 14 13 1 9 0 8 8 9 9 9 0 1 8 7 9 1 9 7 9 9 0 7 10 0 1 9 1 9 2
67 7 13 9 0 10 9 1 9 0 13 15 9 9 1 9 7 13 1 9 15 9 0 1 9 9 0 0 1 9 9 0 1 13 1 7 15 14 13 1 0 9 9 9 0 15 13 1 9 9 1 15 8 8 0 1 15 1 15 9 9 0 0 8 8 9 0 2
49 7 13 8 1 9 1 9 0 1 7 9 9 13 9 1 9 0 1 9 0 0 7 15 14 13 0 7 9 0 9 9 0 1 9 9 1 9 7 9 9 0 1 15 1 15 9 0 0 2
82 7 1 7 9 14 13 1 9 9 0 1 15 1 15 9 9 9 7 10 9 14 13 9 0 1 9 9 1 9 7 15 13 9 9 7 9 1 9 0 9 12 7 1 9 9 12 7 13 9 0 1 9 1 15 1 9 9 12 7 13 10 9 1 0 1 9 9 9 9 0 0 1 9 7 9 9 1 9 9 0 8 2
64 7 1 9 9 0 13 0 1 9 0 15 13 15 9 0 8 8 9 0 1 9 7 3 13 1 9 8 1 9 1 9 0 8 8 13 9 1 8 7 13 15 1 9 10 9 15 14 13 1 15 9 0 9 1 9 9 7 14 13 1 15 8 9 2
77 7 13 9 9 9 0 0 1 9 15 0 2 1 9 2 7 13 9 12 9 7 13 9 0 1 10 9 9 15 13 1 9 9 9 1 9 9 7 9 0 13 9 9 0 1 9 7 13 0 1 9 15 9 9 0 1 9 9 0 9 9 0 1 9 7 13 9 0 7 13 15 1 9 9 1 0 2
93 7 14 13 0 9 9 8 1 9 9 1 9 15 0 7 13 9 0 1 9 15 1 8 9 8 8 8 8 13 9 0 7 0 13 1 15 13 1 15 9 7 15 15 13 1 7 15 9 0 0 1 9 9 9 7 7 9 13 0 1 9 7 9 0 15 8 13 8 8 1 9 15 1 9 8 8 9 8 1 9 9 0 8 8 9 1 9 0 14 13 1 9 2
25 7 13 9 3 1 9 0 1 9 9 9 0 1 9 9 0 0 7 13 9 9 15 1 9 2
71 7 1 9 10 13 8 1 9 15 1 9 9 1 0 7 14 13 8 8 8 1 9 9 0 1 0 1 9 15 0 15 13 15 9 1 9 0 0 7 14 13 1 15 13 0 1 9 9 7 13 9 1 9 8 8 0 1 0 0 1 9 15 1 9 9 0 8 8 1 0 2
61 9 7 10 9 0 14 13 1 15 1 9 9 9 1 9 15 14 13 1 9 9 1 9 15 9 9 1 9 1 9 0 1 9 7 1 15 7 7 9 13 1 10 9 1 7 15 9 1 9 0 15 13 1 9 15 0 7 0 1 9 2
68 7 9 15 13 9 15 15 14 14 13 8 0 1 9 9 1 9 0 9 7 7 8 14 13 9 8 8 9 1 9 13 1 2 7 1 15 7 13 8 0 2 1 9 1 9 9 1 9 8 8 9 8 0 8 9 9 8 15 13 8 8 0 9 8 0 1 0 2
93 7 1 9 8 8 9 1 7 9 0 13 9 9 1 1 15 8 7 15 13 0 1 9 15 13 1 15 7 13 1 9 8 0 1 15 7 15 15 13 15 8 8 13 1 9 15 0 9 7 2 9 9 9 13 0 1 0 2 7 15 13 8 8 1 13 1 15 9 8 2 9 2 8 13 9 0 1 10 13 7 9 0 14 13 8 9 15 14 13 8 8 1 2
12 9 1 9 0 2 9 13 1 9 7 9 0
3 9 12 9
36 13 8 8 9 9 9 7 9 1 9 0 1 9 9 0 7 9 14 13 9 1 9 0 7 0 9 1 9 7 9 0 15 13 1 15 2
47 7 13 9 9 1 9 9 9 9 1 8 9 15 7 9 9 0 0 0 13 1 9 9 0 1 9 9 9 1 9 0 9 1 9 0 15 13 1 15 9 1 9 9 1 9 9 2
23 7 13 7 9 0 13 1 9 9 9 0 1 9 0 7 13 9 1 9 1 9 9 2
31 7 13 7 9 13 9 9 1 12 1 9 9 7 9 9 9 0 1 9 12 1 12 7 13 1 9 0 1 9 12 2
40 7 13 1 9 9 9 15 13 9 7 9 0 1 9 0 15 14 13 1 9 2 9 1 7 9 9 0 1 9 0 1 9 9 13 12 1 12 9 12 2
50 7 13 9 9 8 8 9 9 0 0 14 13 1 9 15 9 9 1 9 9 9 9 0 0 0 0 1 9 7 13 1 9 1 9 9 9 0 0 7 13 1 9 9 0 1 9 1 9 0 2
24 13 7 9 13 1 9 9 0 0 0 0 1 9 0 7 0 1 9 9 0 1 9 12 2
8 9 0 8 8 9 1 9 0
3 9 12 9
35 13 9 9 7 9 9 0 1 9 0 8 9 9 3 9 9 7 9 1 9 8 8 9 1 9 9 1 9 0 1 9 0 1 9 2
37 13 8 1 9 0 13 1 15 9 8 1 9 15 8 8 9 9 0 7 0 7 9 1 9 9 0 9 1 15 13 9 9 0 2 8 2 2
65 7 1 9 15 1 9 1 10 7 13 3 9 8 8 9 1 9 0 2 13 9 7 15 1 15 8 14 13 0 9 0 8 8 13 8 8 9 2 0 1 2 7 3 9 0 13 1 9 9 13 0 13 8 8 9 9 1 9 0 8 1 9 15 2 2
28 7 13 2 8 1 9 8 8 8 1 9 1 15 13 15 8 1 9 0 15 14 13 9 1 9 0 2 2
10 12 9 0 13 9 1 9 8 0 8
3 8 12 9
52 13 12 9 0 15 9 9 7 9 7 9 9 9 9 0 1 9 9 0 1 9 9 0 8 1 9 9 8 8 9 0 1 9 9 9 9 0 1 9 9 15 1 10 9 1 9 0 1 9 7 8 2
49 13 9 10 9 9 1 9 8 9 11 8 8 8 9 9 8 9 9 0 7 13 9 9 7 9 15 1 9 15 0 1 9 13 9 1 9 9 9 0 1 9 15 13 9 15 9 1 9 2
23 7 13 9 0 13 1 9 9 7 15 2 13 9 9 9 1 9 9 0 1 9 2 2
65 7 13 9 7 2 9 12 13 8 8 0 1 9 0 1 9 0 0 1 9 8 13 1 9 9 0 1 9 9 0 8 8 8 8 8 8 8 9 8 1 9 0 8 8 0 1 15 1 15 1 9 9 9 9 9 9 0 8 8 1 9 9 0 2 2
63 7 13 0 1 9 15 1 7 2 8 8 8 8 7 13 1 9 0 8 1 9 9 1 1 9 8 9 0 8 8 9 1 1 13 7 13 8 8 1 9 9 0 1 9 8 1 9 9 1 9 9 15 13 9 0 1 9 1 9 9 0 2 2
15 9 13 1 9 9 0 9 0 1 9 9 9 1 9 0
62 9 13 1 9 9 0 9 0 1 9 9 9 1 9 0 9 12 9 2 8 2 13 9 9 3 9 9 1 9 7 13 0 9 0 13 1 9 9 0 1 9 9 1 9 7 9 9 13 1 9 9 9 0 1 9 9 7 9 0 1 9 2
80 7 13 9 9 0 2 8 2 7 9 0 0 13 1 9 0 15 13 9 1 9 9 0 8 8 8 7 9 0 7 9 13 8 1 9 15 9 9 0 1 9 9 0 1 9 9 0 9 0 13 1 9 1 9 9 1 9 7 9 9 13 1 8 9 9 0 8 8 9 8 8 8 0 7 9 1 8 10 9 2
46 7 13 9 13 1 9 7 9 0 13 1 9 15 0 8 8 9 8 8 8 8 8 8 13 1 10 9 0 9 7 9 0 13 1 7 13 9 9 1 10 9 1 9 9 0 2
23 7 13 9 1 9 9 9 1 9 7 9 1 9 1 9 1 9 9 8 8 9 0 2
11 9 0 13 9 1 9 15 9 1 9 15
3 9 12 9
102 13 9 9 9 9 0 1 9 9 1 9 1 7 13 1 9 0 1 9 0 13 12 9 2 7 13 9 9 0 2 8 2 7 9 9 8 7 9 9 14 13 9 8 8 0 1 14 12 1 9 9 0 7 15 1 9 0 0 7 13 1 9 1 9 0 0 1 9 9 7 9 8 2 13 7 9 9 2 12 9 2 14 13 1 9 1 9 7 13 9 1 9 9 9 9 7 9 15 0 9 0 2
38 7 13 9 9 8 14 13 1 9 1 9 7 9 7 14 13 1 9 7 13 1 9 0 1 7 13 1 9 0 1 9 9 0 1 9 8 8 2
30 0 1 9 7 9 13 1 9 9 0 1 9 9 0 1 9 7 14 13 9 1 15 13 9 9 1 9 9 0 2
7 9 9 0 1 8 7 8
3 8 12 9
29 13 9 0 9 7 8 13 8 8 9 0 1 8 8 13 8 8 1 9 15 3 8 8 9 8 1 8 8 2
28 7 13 15 9 9 15 13 1 9 1 9 0 1 9 9 9 8 8 7 9 0 1 9 9 15 8 8 2
20 7 13 9 0 15 9 8 1 9 9 8 1 9 1 9 8 1 9 8 2
23 7 14 13 8 1 9 8 8 8 7 13 15 9 1 9 0 9 0 8 8 8 8 2
32 13 8 9 0 1 9 8 1 9 0 12 9 1 9 2 7 13 1 9 15 1 9 1 9 9 0 1 8 1 9 0 2
8 9 0 8 9 9 1 9 8
3 8 12 9
39 13 9 9 1 9 1 9 8 0 1 9 1 9 9 1 9 8 1 8 9 9 1 9 8 13 1 7 15 1 9 8 9 1 15 13 9 0 9 2
32 7 13 9 7 9 15 9 1 9 9 0 1 9 7 15 13 3 9 7 7 9 0 1 9 9 8 8 8 8 13 9 2
23 7 9 1 15 13 9 7 7 9 0 13 1 9 9 0 1 9 9 9 1 9 9 2
23 7 14 13 9 7 9 7 9 8 8 9 1 9 1 9 9 9 7 9 9 8 9 2
19 7 14 13 9 8 8 8 9 12 9 0 7 9 9 0 1 12 9 2
27 7 13 8 8 9 1 9 9 8 7 9 8 7 9 9 8 1 9 8 1 9 9 0 1 10 9 2
38 7 14 13 9 0 7 15 1 9 8 1 9 0 1 12 1 12 9 1 9 0 13 0 1 12 12 0 9 15 1 9 9 0 7 0 7 0 2
7 8 13 8 0 1 9 9
4 8 8 12 9
28 13 9 9 0 8 8 9 8 9 9 0 1 9 9 0 8 8 8 1 9 9 9 1 15 13 9 0 2
25 13 9 1 9 1 9 8 1 9 0 7 9 15 14 13 9 0 0 8 8 9 0 1 9 2
28 7 13 9 9 9 1 8 1 8 1 8 0 8 8 9 0 0 1 8 8 9 9 9 1 15 13 9 2
32 7 13 8 7 9 0 13 1 9 15 7 13 15 9 9 15 13 1 9 0 1 9 8 9 0 1 9 9 0 8 8 2
48 7 13 8 14 13 9 0 9 1 8 7 13 7 9 0 14 13 9 9 15 1 9 9 0 1 9 7 9 8 8 8 1 9 9 1 9 1 9 0 1 9 8 8 7 13 9 0 2
26 7 13 8 8 7 9 14 13 0 9 13 1 8 9 0 7 9 9 8 8 0 1 9 7 9 2
27 7 13 8 7 15 13 9 0 1 8 1 9 9 1 9 1 9 15 0 1 9 15 0 9 12 9 2
24 7 13 9 0 0 14 13 9 15 7 13 9 0 1 9 9 0 1 9 0 1 9 12 2
41 7 14 13 9 8 8 9 9 8 8 0 9 9 1 9 15 1 7 9 9 0 14 13 1 9 9 7 12 9 9 1 15 13 1 9 1 9 8 8 0 2
34 7 13 7 9 13 7 8 9 9 7 13 9 0 1 9 1 9 9 0 1 9 8 8 7 9 9 8 8 9 1 9 9 0 2
10 9 1 9 9 1 9 9 1 9 8
3 8 12 9
34 13 7 9 13 9 15 1 9 1 8 1 9 9 1 9 0 1 9 9 0 1 9 8 1 9 9 1 9 8 7 13 9 0 2
27 7 13 1 9 9 9 15 7 9 13 8 8 9 1 9 15 13 9 9 1 9 1 15 1 9 0 2
32 7 13 8 7 9 0 14 13 13 1 9 1 9 8 9 7 7 9 13 1 15 8 9 1 9 15 1 9 1 9 9 2
23 7 13 8 8 9 9 1 9 9 8 9 7 7 15 13 7 9 9 8 14 13 1 2
13 9 0 2 9 0 1 9 1 9 1 9 9 9
64 9 0 2 9 0 1 9 1 9 1 9 9 9 9 12 9 2 8 2 13 9 9 9 0 1 9 0 1 9 7 9 9 9 0 8 8 1 12 9 0 1 15 13 12 1 9 9 1 9 9 0 9 0 8 8 9 8 1 8 8 8 9 0 2
54 7 1 9 15 13 0 7 14 9 0 13 8 8 1 9 1 9 9 9 7 9 9 9 0 0 1 9 9 0 0 7 3 9 9 9 8 8 1 9 0 1 9 7 9 0 1 15 1 9 8 8 9 0 2
39 7 13 9 1 9 15 13 9 1 9 0 9 1 9 9 7 9 7 9 9 8 8 9 9 8 8 8 8 9 7 9 0 8 7 9 9 8 9 2
77 7 1 9 7 12 9 8 8 0 7 0 13 9 15 12 9 13 9 9 15 1 9 8 8 9 0 13 8 1 9 1 9 9 8 9 1 9 7 13 8 8 9 13 15 7 14 13 9 1 9 15 1 9 0 1 15 1 9 0 0 7 1 9 0 8 8 8 15 13 15 8 1 9 0 1 9 2
46 7 14 13 10 9 1 8 9 1 10 1 15 8 8 13 8 8 9 0 7 14 13 13 9 7 9 1 9 1 7 8 8 8 9 9 8 8 13 1 9 9 7 1 9 0 2
33 7 13 9 3 7 15 1 9 9 13 1 9 9 1 9 7 9 9 7 9 9 13 8 1 9 7 9 1 9 15 1 9 2
29 8 9 1 15 7 14 13 9 8 8 9 9 0 9 1 8 7 15 13 9 0 1 9 0 7 0 15 0 2
88 7 1 9 0 1 9 8 7 1 9 13 1 9 7 9 0 12 8 13 8 8 9 0 2 7 13 8 8 1 9 1 7 15 0 9 7 9 8 9 0 13 1 9 13 1 9 9 1 15 8 1 9 8 8 8 8 8 13 1 15 8 0 8 2 7 14 13 9 15 13 1 10 9 7 15 7 13 0 1 15 1 8 0 7 1 9 8 2
44 9 7 9 10 9 13 1 9 9 9 9 8 8 1 15 15 13 9 9 1 15 13 9 0 9 1 9 0 7 13 15 1 9 15 7 15 14 13 9 15 1 9 15 2
29 7 1 9 13 9 0 7 13 9 0 9 0 1 9 8 0 8 1 9 9 15 9 7 9 13 8 8 8 2
32 8 10 9 1 8 9 15 14 13 7 13 9 1 8 1 9 9 9 0 1 9 7 15 1 9 13 8 1 10 0 0 2
49 7 1 1 9 0 9 8 9 3 9 1 9 8 15 13 9 8 1 9 0 0 7 13 9 1 9 9 0 7 12 9 2 7 14 13 9 7 13 9 1 10 9 1 7 8 9 9 9 2
54 7 1 15 13 8 1 9 9 15 13 1 15 8 7 9 0 1 9 9 0 9 15 13 1 9 9 7 9 1 9 7 1 15 9 15 13 1 12 9 0 1 9 8 9 9 7 13 1 12 9 7 12 9 2
51 8 0 8 8 9 8 7 14 13 9 7 9 8 1 9 9 7 14 13 8 7 9 13 9 15 0 7 14 13 9 0 8 9 13 9 7 7 15 1 9 9 15 13 9 1 9 15 13 9 9 2
14 9 9 0 13 1 9 2 9 2 1 8 7 9 9
3 8 12 9
36 13 9 9 0 8 8 8 1 0 9 0 1 15 8 8 8 9 9 2 7 13 1 9 2 9 2 7 9 9 0 0 1 9 0 0 2
16 13 8 1 9 8 0 1 9 1 9 1 9 13 9 0 2
18 7 13 8 9 9 1 9 15 7 8 14 13 9 3 1 9 15 2
26 7 13 8 1 9 9 9 0 1 9 9 0 8 8 9 1 9 9 9 1 9 0 1 9 0 2
35 7 13 8 2 2 7 9 8 1 9 1 9 9 0 2 8 8 8 1 7 8 14 13 9 1 9 0 2 0 1 9 1 9 2 2
32 13 7 9 0 13 0 9 2 9 2 2 7 13 3 1 15 1 8 9 9 0 1 9 1 9 9 9 1 9 9 0 2
29 7 13 9 9 0 8 7 9 15 13 9 9 1 9 1 9 1 9 0 2 7 13 9 9 0 1 15 2 2
39 7 13 8 7 9 9 9 8 8 2 13 1 9 8 8 2 2 9 9 15 2 8 8 8 8 8 8 0 2 8 8 8 9 7 8 1 15 2 2
23 7 13 8 9 9 0 1 2 9 9 8 0 2 15 14 13 1 15 1 9 9 15 2
28 7 13 8 7 9 0 1 9 9 8 0 13 7 8 2 8 7 2 8 15 0 9 1 9 8 8 2 2
45 13 9 9 8 1 9 13 1 15 9 0 7 9 13 1 15 9 9 1 9 0 1 9 9 12 1 9 9 8 1 8 2 8 9 0 1 9 15 13 1 15 9 0 3 2
33 7 14 13 9 9 7 0 9 9 9 1 9 1 9 1 9 9 0 2 1 7 13 9 9 9 9 9 0 1 9 9 9 2
9 9 0 0 13 0 9 1 9 8
3 8 12 9
43 13 8 8 8 2 9 9 9 0 0 7 9 9 9 8 1 9 9 1 9 9 15 7 9 15 1 9 0 1 9 0 15 13 1 9 8 9 0 0 2 8 2 2
38 13 8 2 7 15 3 9 9 0 1 9 0 1 9 0 0 7 9 9 9 2 1 9 1 9 1 8 8 8 9 9 0 0 7 9 9 0 2
28 7 1 9 1 9 9 15 13 15 8 13 8 9 9 2 13 8 9 9 2 7 13 1 9 1 8 8 2
29 7 13 8 1 9 8 8 8 8 8 0 1 9 8 2 15 13 9 9 1 9 9 1 9 1 15 8 8 2
37 13 7 15 1 9 9 9 8 1 8 2 13 9 0 0 12 1 9 0 1 9 0 1 9 7 9 0 1 9 9 1 9 1 9 8 8 2
24 7 13 8 9 8 3 1 7 8 8 8 7 7 13 1 9 1 9 1 8 9 9 15 2
6 9 9 9 0 1 8
3 8 12 9
27 13 9 9 9 0 1 8 9 13 9 8 8 8 8 1 9 8 9 9 9 9 9 8 8 1 15 2
35 13 9 0 2 1 1 9 0 2 7 8 8 8 1 9 15 13 8 8 12 9 9 0 0 2 8 8 1 9 0 1 9 9 9 2
29 13 9 9 2 15 13 9 1 12 9 2 1 8 8 1 12 12 9 8 8 2 8 8 8 9 8 1 8 2
11 13 9 8 1 9 8 8 1 9 12 2
20 12 0 13 1 8 9 1 15 8 8 14 13 12 1 15 9 0 9 1 15
70 12 0 13 1 9 9 1 15 9 1 8 14 13 12 1 15 9 0 9 1 15 8 12 9 2 8 2 13 9 9 0 9 7 12 9 0 13 1 9 9 0 1 8 1 0 1 9 0 13 13 1 9 15 12 1 9 0 0 1 8 2 9 1 15 13 15 9 9 8 2
41 7 13 9 7 15 1 9 14 13 9 1 9 1 8 8 9 0 2 7 13 9 7 13 1 9 0 1 9 1 9 0 8 8 8 0 1 9 0 1 8 2
20 13 9 2 15 13 1 9 9 8 8 7 8 8 2 1 8 8 1 8 2
57 7 13 9 7 9 0 13 3 9 7 9 0 13 1 9 9 0 8 9 0 0 2 8 2 2 7 13 7 14 12 9 0 15 13 1 15 9 9 0 1 9 1 9 0 2 1 15 13 7 14 12 9 0 14 13 8 2
10 9 9 9 7 8 13 9 0 1 8
3 8 12 9
23 13 9 9 0 8 8 8 7 9 15 0 8 8 9 1 8 8 9 13 1 9 0 2
50 7 13 8 8 1 9 9 15 13 1 15 9 1 9 0 8 8 8 14 12 1 9 9 15 13 1 15 8 1 8 0 1 9 0 0 0 1 7 9 9 9 9 9 9 0 1 9 1 9 2
45 7 13 8 9 15 0 1 9 9 8 1 9 9 0 1 9 15 14 13 15 9 0 7 9 0 1 9 9 0 2 7 13 7 9 0 13 7 13 9 0 1 10 9 0 2
23 7 13 8 7 8 0 1 9 9 1 9 1 8 9 9 0 8 8 9 1 9 0 2
63 7 1 9 15 13 8 7 9 0 13 9 0 2 7 13 9 1 0 1 9 9 1 8 1 10 9 2 7 13 1 9 0 1 9 1 9 0 9 1 9 1 9 1 9 0 1 10 9 2 1 9 1 9 1 9 0 1 9 9 1 10 9 2
23 7 13 9 9 9 1 9 1 9 8 2 7 9 9 1 8 9 0 0 2 8 2 2
10 8 9 13 9 1 9 0 8 1 8
3 8 12 9
23 13 8 9 0 1 9 9 1 9 15 1 9 9 9 0 15 13 1 9 15 1 8 2
30 7 13 9 1 9 9 8 8 1 9 0 7 9 13 8 8 9 1 9 1 9 8 0 1 9 0 1 9 0 2
37 7 14 13 8 0 1 9 7 1 8 8 0 13 8 8 1 9 1 9 9 15 1 9 9 2 7 13 1 8 8 8 8 9 9 1 8 2
31 7 13 8 7 8 13 12 9 13 8 8 13 9 8 8 8 8 8 8 9 8 8 8 1 1 12 9 1 14 8 2
51 7 13 8 7 8 8 1 7 13 15 1 12 1 12 12 1 9 0 2 13 7 15 13 1 9 9 15 2 7 13 8 9 8 8 8 8 8 8 1 9 15 1 8 0 1 9 8 9 1 9 2
31 7 13 8 8 9 9 9 1 9 2 8 8 8 1 9 1 15 8 8 1 10 9 15 14 13 9 1 9 0 2 2
54 7 13 2 7 0 1 15 13 8 9 2 8 8 7 13 8 7 15 13 9 1 9 0 2 7 14 13 9 1 15 2 8 8 1 1 9 15 8 8 1 9 1 8 0 1 9 10 13 1 15 9 0 2 2
6 0 9 1 8 9 0
3 8 12 9
74 8 8 13 0 9 1 8 9 0 2 2 2 8 8 2 2 2 2 2 13 9 8 1 9 15 0 1 9 15 13 1 15 9 9 0 0 1 9 7 13 1 9 8 8 9 1 8 3 1 9 9 0 0 1 9 8 8 9 8 1 9 1 9 1 0 1 9 15 8 8 1 9 15 2
58 2 2 1 9 9 1 9 9 1 9 9 0 2 14 13 9 9 1 8 13 1 9 9 2 7 9 9 9 2 7 9 9 1 0 9 2 7 9 15 1 9 9 8 1 15 1 9 9 0 2 7 9 9 1 9 0 0 2
58 2 2 8 8 2 2 2 13 9 9 14 13 15 9 0 7 8 7 8 9 9 1 9 0 1 9 9 0 0 1 9 2 9 9 0 1 9 1 9 9 0 7 8 1 9 9 0 8 8 8 0 1 9 14 13 1 9 2
63 2 2 13 3 9 9 0 1 9 9 1 9 15 8 8 9 0 15 13 1 9 9 1 9 13 9 12 9 0 2 8 1 10 9 8 8 9 0 9 1 9 14 13 1 9 15 9 9 9 1 9 1 9 0 1 9 15 1 9 1 9 0 2
8 9 13 9 0 1 9 1 9
3 9 12 9
36 13 9 9 9 9 9 0 9 0 9 9 9 9 9 9 0 9 1 9 1 9 7 13 15 1 9 1 9 1 9 9 15 1 9 15 2
37 7 13 7 15 14 13 3 9 1 9 9 15 14 13 9 0 1 9 1 9 9 15 1 9 15 2 7 9 9 0 1 9 15 13 15 9 2
22 7 13 9 1 12 1 9 9 1 7 9 0 14 13 9 9 1 9 7 1 0 2
18 7 13 1 7 9 14 13 9 0 7 13 9 0 9 1 10 9 2
76 7 13 0 2 7 9 0 13 9 0 7 13 7 1 9 15 9 9 1 9 9 1 9 9 1 1 9 9 1 9 0 2 7 14 13 9 15 14 13 1 15 9 0 9 10 9 2 2 7 13 9 1 9 0 0 1 7 9 13 1 9 0 1 9 2 0 7 9 0 13 9 9 9 0 0 2
18 7 13 7 9 13 9 9 9 1 9 2 7 13 9 1 10 9 2
31 7 13 1 7 9 0 14 13 1 9 0 1 7 13 9 15 2 7 13 9 1 9 9 1 9 9 0 1 9 15 2
69 7 13 9 1 9 0 2 7 9 9 13 9 9 1 9 7 13 1 9 9 9 7 9 1 10 1 15 1 9 9 9 9 2 2 7 13 7 2 9 1 9 13 9 0 1 9 2 7 13 1 15 15 7 15 13 1 15 7 13 7 13 7 13 1 9 9 0 2 2
7 9 9 9 0 8 1 9
3 9 12 9
24 13 9 0 0 0 8 8 9 8 8 1 9 0 2 13 8 9 0 0 8 8 8 9 2
37 7 1 9 15 1 8 1 9 15 13 8 2 7 8 9 9 0 1 9 0 1 9 2 14 13 9 1 9 7 13 9 1 9 9 1 9 2
22 7 13 9 7 15 13 1 7 13 9 0 1 9 0 1 9 9 7 9 1 9 2
32 13 7 9 2 15 13 1 9 1 9 1 0 1 12 9 2 13 9 15 13 1 9 9 0 1 9 9 0 9 12 9 2
34 13 9 0 1 9 0 8 8 8 0 1 9 0 8 9 9 1 9 9 1 9 2 7 13 9 1 9 1 8 8 8 8 8 2
28 13 9 1 7 9 9 9 9 0 2 7 13 9 9 1 15 12 1 12 1 9 9 9 0 12 12 9 2
10 9 0 13 9 8 1 9 2 9 2
3 8 12 9
37 13 9 0 8 8 9 9 2 9 2 15 13 1 15 9 9 0 8 8 8 1 9 15 13 9 0 1 9 8 1 9 9 0 1 9 0 2
43 7 13 8 15 13 1 9 9 9 1 9 1 9 1 0 9 0 1 15 7 3 2 9 15 9 2 1 9 2 7 7 0 9 0 13 7 2 13 1 10 9 2 2
36 7 1 9 13 1 15 2 13 8 2 7 8 0 0 8 8 9 1 8 2 13 1 9 0 9 1 9 9 2 7 9 9 0 9 9 2
38 7 13 8 2 7 9 9 9 9 12 7 12 13 9 2 9 9 8 0 2 8 8 7 13 1 9 15 2 7 13 9 1 9 9 1 15 2 2
31 7 13 2 7 9 9 10 9 13 7 9 0 14 13 7 14 13 15 7 13 9 8 8 9 1 9 7 9 8 8 2
10 9 9 13 8 8 9 9 0 1 9
4 9 0 12 9
22 13 9 9 0 9 0 9 8 8 9 9 0 1 9 0 1 9 9 0 1 9 2
31 13 9 9 8 1 9 1 9 0 15 13 9 9 1 9 1 8 7 8 2 8 9 9 15 13 15 9 0 1 9 2
37 7 1 9 1 9 2 13 9 9 9 8 8 0 9 1 9 7 9 0 7 0 1 9 0 2 13 7 13 9 0 8 8 8 8 1 9 2
23 7 13 7 9 13 9 1 8 0 9 2 7 7 9 14 13 9 1 9 10 9 0 2
29 7 13 9 9 1 7 13 9 0 0 8 9 8 13 1 12 9 2 7 14 13 1 15 9 9 9 9 0 2
47 7 1 9 1 8 9 3 9 2 13 9 0 1 9 0 8 8 7 9 0 2 1 15 9 0 13 15 1 9 9 0 2 7 9 9 8 9 2 7 9 1 9 9 0 0 2 2
18 14 7 9 0 13 9 0 3 9 0 0 1 9 8 9 9 0 2
17 7 13 9 7 9 14 13 9 0 1 9 9 15 13 12 9 9
8 8 13 9 9 8 0 9 0
3 8 12 9
24 13 9 0 9 7 9 15 13 15 9 8 0 0 1 9 9 0 1 8 8 13 9 0 2
66 7 13 9 9 0 1 9 8 8 8 8 8 2 7 13 9 8 0 8 1 9 1 9 9 0 2 7 14 8 13 9 0 7 9 14 13 9 1 15 2 2 13 15 1 9 0 1 9 15 1 9 9 1 9 9 1 9 0 2 0 0 9 0 1 9 2
38 7 13 9 9 2 1 0 7 13 9 0 15 15 9 8 0 2 2 1 9 0 13 9 9 8 8 8 7 9 0 13 1 10 9 1 9 0 2
63 7 13 8 1 9 1 9 9 1 9 0 1 9 8 8 8 9 3 2 7 9 13 0 1 9 15 1 8 8 2 2 7 1 9 9 2 13 9 9 0 8 9 8 8 7 9 0 0 14 13 9 0 1 9 9 2 7 9 9 1 8 8 2
29 7 13 8 2 13 9 13 9 0 0 9 15 2 7 4 0 9 0 2 7 13 7 9 9 0 13 7 13 2
87 13 7 15 1 9 3 2 13 9 9 8 8 1 9 9 8 8 2 1 15 1 15 8 1 9 0 2 7 9 1 13 8 1 9 8 8 8 9 0 2 7 9 8 1 9 2 7 9 8 8 8 2 8 2 8 2 1 9 2 1 9 9 9 15 13 15 9 1 12 9 7 13 9 9 1 15 7 13 14 13 9 9 9 8 8 9 2
18 13 9 14 13 9 13 8 9 9 7 8 1 9 9 8 9 3 2
15 0 9 1 9 9 9 9 1 9 2 9 0 7 0 2
61 8 9 1 9 9 8 9 1 9 2 9 0 7 0 2 2 13 9 9 8 9 0 1 9 9 1 9 9 7 9 15 1 0 8 8 9 9 9 1 9 9 12 2 7 7 15 13 9 10 9 1 12 1 12 0 1 1 12 1 12 2
59 2 13 9 9 1 9 8 1 9 9 0 9 1 9 1 9 12 9 2 7 13 1 12 12 9 1 9 9 0 0 8 0 1 9 15 13 15 9 0 2 7 14 13 8 8 9 8 1 9 1 9 8 9 1 9 9 0 0 2
41 2 13 9 9 8 0 9 0 1 9 8 0 1 9 8 0 2 7 9 9 8 2 7 9 1 9 0 7 8 1 8 9 9 9 8 8 8 0 8 8 2
33 2 13 9 9 9 0 7 8 2 1 9 9 2 1 9 0 8 8 12 9 2 7 13 10 9 0 7 13 9 9 9 15 2
37 2 8 9 9 9 9 1 9 9 0 0 15 13 8 8 1 9 0 8 8 0 1 9 2 8 8 8 1 9 15 2 7 9 9 1 15 2
13 9 9 8 2 9 9 1 9 14 13 9 1 9
4 8 8 12 9
50 13 9 9 8 8 8 8 8 8 9 7 8 14 13 9 9 1 9 1 7 9 2 7 0 9 1 9 15 14 8 9 1 9 15 13 15 9 0 1 9 2 9 1 15 13 15 9 9 8 2
59 7 13 9 9 9 1 9 9 2 7 0 9 15 7 15 14 13 1 9 9 1 9 9 13 1 15 7 13 9 1 9 1 9 0 2 2 13 15 9 1 9 8 3 9 9 15 9 9 9 1 9 9 0 1 9 9 1 9 2
31 7 13 7 8 13 3 1 9 7 13 0 9 9 13 1 9 0 9 9 0 1 9 1 9 15 0 7 9 15 0 2
45 7 13 9 9 8 8 8 9 1 10 2 9 9 1 9 8 8 8 13 15 9 0 1 9 2 8 8 9 0 1 9 8 9 0 0 2 8 8 9 0 1 9 8 8 2
37 7 13 1 7 8 13 0 9 15 13 1 9 0 1 12 9 1 9 9 1 9 2 7 13 1 7 9 13 1 8 7 9 1 9 0 0 2
45 7 13 1 9 9 0 7 0 15 8 7 8 9 9 9 1 9 0 1 9 9 0 0 2 7 9 15 13 9 10 9 15 9 9 15 13 1 9 1 1 1 9 10 9 2
56 7 13 9 9 8 8 8 7 9 9 0 8 8 8 8 13 9 1 9 1 9 9 12 1 8 9 0 2 7 13 7 9 8 14 13 15 1 9 13 3 1 9 8 7 7 13 1 9 9 0 1 9 0 1 9 2
11 9 9 12 9 1 8 9 8 8 1 9
3 8 12 9
37 13 7 13 1 12 9 14 13 9 15 7 13 12 0 1 9 0 1 9 0 1 9 9 13 13 1 9 8 2 9 1 15 13 15 9 0 2
30 13 9 0 2 7 15 1 9 8 12 13 9 1 9 9 8 8 8 1 9 8 1 9 8 9 0 9 8 0 2
34 7 13 7 9 9 13 1 9 7 13 9 0 1 9 1 9 12 8 9 2 12 9 2 9 1 9 9 1 8 8 9 3 9 2
23 7 13 8 0 1 9 8 7 9 9 13 1 1 15 9 9 1 9 0 8 8 8 2
21 7 1 9 9 1 1 12 9 2 13 8 9 1 9 1 8 8 8 1 15 2
24 7 13 9 9 0 8 8 7 9 13 9 3 2 7 7 15 13 7 15 14 13 9 9 2
16 7 13 9 8 8 8 0 7 1 12 9 14 13 1 9 2
10 8 13 1 9 15 0 1 9 1 9
3 8 12 9
27 13 9 0 8 8 9 1 9 9 15 0 1 9 15 13 15 9 0 1 9 7 9 9 1 8 0 2
36 7 1 9 15 1 9 9 0 1 8 2 13 8 7 9 1 8 7 9 0 2 9 8 8 2 2 7 7 15 1 0 9 9 1 9 2
34 7 13 7 8 0 1 9 1 9 0 0 7 0 1 9 0 2 13 9 9 8 9 2 7 14 13 9 15 1 9 1 9 0 2
33 7 13 7 8 14 13 1 9 15 0 2 8 9 15 8 8 8 13 1 7 15 14 13 1 9 0 1 9 0 13 1 8 2
13 7 13 0 7 9 0 0 14 13 9 9 0 2
26 7 13 8 1 9 9 9 1 8 2 0 7 9 1 8 7 9 0 9 8 8 1 9 1 8 2
11 9 9 0 13 1 9 9 1 9 1 9
3 8 12 9
27 13 9 9 0 1 9 9 0 12 2 12 1 9 1 9 0 15 13 9 9 9 1 9 8 8 12 2
27 13 9 9 9 9 9 8 8 8 1 8 8 7 8 8 8 1 8 2 7 13 9 9 9 9 3 2
80 7 13 8 1 9 15 13 9 3 9 2 7 15 9 0 13 1 9 10 1 12 9 2 2 7 13 2 7 8 0 1 9 13 7 13 3 9 0 8 8 8 3 2 2 7 13 9 0 9 9 9 2 15 13 1 9 9 7 9 0 1 15 2 1 9 1 9 0 3 7 14 13 1 9 1 9 7 9 8 2
44 7 13 9 9 9 1 9 8 8 12 1 9 9 9 9 1 9 1 9 0 1 9 9 9 1 9 9 0 2 7 13 8 7 8 2 8 8 8 8 2 7 9 0 2
11 9 0 13 8 8 9 9 0 1 9 0
3 8 12 9
27 13 9 8 8 9 7 9 0 14 13 8 8 9 9 0 1 9 0 1 9 9 9 7 9 1 9 2
39 7 13 9 1 9 0 8 8 8 9 15 7 8 14 13 9 0 1 9 0 8 8 8 8 9 9 0 1 12 9 1 9 9 8 8 1 8 9 2
45 7 13 9 7 8 14 13 3 7 15 14 13 9 9 8 8 8 8 9 0 8 8 1 9 0 0 0 9 15 1 9 9 0 1 9 1 9 9 0 8 8 9 1 9 2
17 7 13 9 7 9 14 13 1 9 0 1 9 1 9 9 0 2
34 7 13 9 7 8 14 13 1 9 9 0 7 9 15 13 1 9 0 1 9 9 8 8 7 9 9 9 0 7 9 9 9 0 2
29 7 1 9 13 9 0 9 9 0 1 8 7 9 2 7 1 0 7 13 1 9 9 1 9 1 9 9 0 2
90 7 13 9 7 9 14 13 1 9 1 9 2 7 15 13 3 1 9 0 15 13 9 9 15 7 9 2 13 7 15 9 0 7 13 9 0 1 0 1 9 2 2 7 13 9 1 8 8 1 9 8 1 9 9 0 9 15 7 9 9 0 1 9 14 13 0 2 7 15 14 13 0 1 9 9 7 9 1 9 9 2 7 3 9 9 0 1 9 2 2
14 8 13 7 15 14 13 8 8 8 9 9 0 1 9
53 8 13 7 15 14 13 9 1 9 9 9 0 1 9 8 12 9 2 8 2 13 9 9 0 8 8 9 1 7 15 14 13 9 1 9 9 9 0 7 0 1 9 2 7 7 15 1 9 14 13 1 9 2
42 7 1 9 0 8 8 1 9 8 8 9 9 0 1 9 2 13 8 7 9 9 15 13 15 9 0 1 9 9 0 1 9 9 0 2 14 13 9 9 9 2 2
30 7 13 2 7 9 15 13 7 15 13 9 15 14 13 15 10 9 2 7 13 9 15 2 14 15 9 9 0 2 2
33 7 13 1 7 9 0 2 0 1 9 1 0 9 1 9 13 0 7 0 1 9 1 9 15 13 15 8 9 0 13 8 2 2
20 7 13 8 7 15 14 13 9 1 9 15 14 13 15 9 0 0 1 9 2
29 7 13 2 7 9 10 7 13 9 8 8 13 9 7 9 7 12 2 2 2 15 9 14 13 15 1 9 2 2
5 0 0 13 1 9
3 9 12 9
30 13 1 9 9 9 9 9 0 0 0 1 9 0 9 7 1 9 15 12 9 7 0 7 0 15 1 9 9 15 2
34 7 13 9 0 0 0 1 9 0 0 1 9 1 9 10 9 1 10 13 9 15 9 0 7 9 0 0 1 15 13 9 9 0 2
53 7 13 9 7 9 9 7 0 0 1 9 9 0 0 9 1 9 9 0 9 9 11 11 7 9 9 9 11 9 9 9 9 9 9 9 9 7 9 9 0 7 9 9 11 9 9 9 0 1 9 9 9 2
40 7 1 9 0 1 9 2 13 9 15 1 9 9 0 7 9 9 9 1 9 0 7 9 9 9 7 9 9 9 0 1 9 1 9 2 9 1 9 15 2
44 13 7 9 0 0 7 9 0 0 13 14 13 9 0 0 1 9 2 9 2 1 9 7 0 1 9 2 8 8 2 15 13 1 12 9 9 9 1 9 7 9 9 0 2
51 7 13 9 9 7 9 0 0 15 13 0 1 15 1 9 9 7 9 1 9 0 1 9 7 9 0 7 15 13 0 1 9 9 0 0 1 9 9 0 15 13 0 1 9 1 9 14 12 9 0 2
11 12 2 12 2 12 2 12 2 12 2 12
8 9 0 1 8 8 8 9 9
3 8 12 9
34 13 1 3 9 8 8 9 9 0 0 1 9 9 8 1 9 9 1 9 0 13 1 9 9 9 0 1 9 7 9 8 8 0 2
40 8 8 1 9 15 3 15 13 12 9 1 9 9 8 8 2 7 9 9 0 8 2 8 2 8 2 8 8 8 1 9 9 2 7 13 1 15 9 0 2
28 13 9 9 1 9 8 8 8 9 8 8 15 13 1 9 0 2 1 13 9 9 9 1 9 9 12 9 2
54 13 8 7 9 12 8 1 9 9 1 9 0 2 7 14 13 9 2 15 13 9 0 1 9 7 9 9 1 8 9 9 0 0 8 8 2 1 9 15 10 2 7 13 1 9 0 0 1 9 0 1 9 0 2
8 9 0 1 9 0 9 7 9
3 8 12 9
29 13 9 9 0 8 8 8 9 1 9 8 9 8 1 9 15 0 8 8 13 1 15 9 9 9 1 9 9 2
46 7 13 8 9 9 1 9 9 1 9 10 1 9 8 8 8 7 13 7 9 13 7 8 9 1 9 1 9 1 8 9 0 2 7 13 7 9 14 13 9 0 8 1 9 0 2
56 7 13 8 7 9 1 9 10 1 9 13 9 0 9 9 1 7 1 10 9 13 7 13 1 9 9 0 1 9 0 7 9 1 9 7 9 1 9 7 1 3 7 7 15 13 9 1 10 9 9 1 9 9 9 0 2
41 7 13 7 3 9 0 1 9 7 9 1 10 9 7 7 9 14 13 1 9 0 1 10 1 15 9 7 14 13 1 9 0 1 9 9 1 9 10 1 9 2
59 7 1 9 15 13 8 8 7 9 0 1 9 13 1 9 7 7 15 13 1 9 9 0 7 13 9 0 1 9 9 7 9 1 9 1 15 13 7 13 1 15 15 1 9 9 9 7 9 9 9 15 7 9 9 7 9 1 9 2
55 7 13 9 1 9 15 7 9 15 1 9 7 15 14 13 1 1 9 9 9 0 0 2 8 2 0 7 9 0 14 13 1 9 9 0 1 9 15 1 9 8 7 7 9 0 14 13 9 0 1 9 9 1 8 2
10 9 1 9 9 0 13 9 8 0 0
3 8 12 9
24 13 9 1 9 9 0 9 8 1 0 9 8 8 8 0 8 8 1 9 8 1 9 8 2
40 13 7 9 15 13 9 0 1 9 0 1 9 8 1 9 9 14 13 9 9 9 0 1 9 9 9 9 9 9 0 0 0 2 8 2 1 9 0 0 2
24 7 1 9 9 0 1 9 9 9 1 9 0 2 13 8 1 9 12 9 8 7 12 9 2
33 7 13 8 8 9 9 9 9 9 15 13 9 9 8 7 9 15 1 9 13 1 9 15 13 1 9 12 9 1 9 9 8 2
30 7 13 9 9 9 1 12 9 7 13 9 15 1 0 1 9 7 13 9 9 12 9 1 15 13 1 7 15 8 2
28 7 13 9 0 7 15 1 9 9 15 13 12 9 2 13 1 9 1 9 1 9 15 7 9 1 9 9 2
33 7 13 8 15 13 13 1 9 0 7 15 13 1 9 9 0 1 9 2 2 7 13 2 14 15 9 0 15 13 9 13 2 2
38 7 13 9 0 8 1 7 9 9 13 9 8 9 0 1 9 9 1 0 2 7 13 2 7 1 15 8 0 1 12 12 9 1 9 1 9 2 2
9 9 9 9 9 8 14 13 12 9
3 8 12 9
32 13 8 8 8 9 9 1 9 8 0 3 9 7 9 9 9 0 15 13 0 2 14 13 12 12 15 13 1 15 1 9 2
38 7 13 7 15 0 8 3 8 8 2 8 8 8 1 7 3 8 0 1 9 14 12 8 13 1 15 2 7 8 8 8 1 9 1 9 1 10 2
37 13 8 14 13 1 9 9 9 7 15 13 8 12 9 1 7 13 15 9 9 9 8 2 12 15 13 8 9 1 8 1 9 8 0 8 9 2
20 7 13 8 7 9 0 1 9 13 9 1 9 12 9 1 9 8 2 8 2
32 7 13 9 9 0 8 1 9 0 9 7 12 9 3 13 1 9 1 8 0 2 1 1 15 12 1 9 9 7 12 0 2
57 7 13 9 9 9 0 8 8 1 7 8 13 1 12 9 13 7 15 13 8 8 1 9 9 0 9 15 13 1 9 8 9 9 1 9 9 0 1 9 9 7 13 9 1 9 1 9 12 9 1 9 0 9 1 9 8 2
23 7 13 9 1 8 8 0 1 9 2 7 7 15 14 13 9 0 1 10 9 1 9 2
25 7 14 13 9 8 8 8 0 1 1 1 9 15 1 7 9 9 1 9 14 8 1 12 9 2
13 9 1 8 13 9 9 9 8 1 9 1 9 15
3 8 12 9
32 13 9 9 9 9 1 8 3 9 7 9 12 1 9 0 1 9 9 0 0 2 8 2 14 13 9 1 15 13 1 9 2
55 7 13 9 1 9 9 7 15 1 0 1 9 7 7 13 9 9 10 9 1 9 9 8 1 0 7 7 15 14 13 9 12 1 10 9 7 15 9 7 12 9 1 9 1 9 15 1 9 0 1 9 15 1 8 2
22 7 1 9 0 12 9 1 9 8 1 9 7 7 9 8 7 9 13 9 1 9 2
50 7 14 13 1 9 3 9 0 13 1 8 0 8 8 8 7 7 9 14 13 9 15 1 7 15 0 1 9 9 2 7 14 13 9 10 9 1 9 0 1 9 9 1 9 0 1 15 13 9 2
14 9 8 2 9 9 13 1 9 8 8 8 8 9 9
41 9 8 2 9 9 13 1 9 8 8 8 8 9 9 8 8 12 9 2 8 2 13 9 1 9 7 13 8 9 1 9 0 7 15 9 9 9 10 1 9 2
15 7 14 13 9 9 9 9 0 1 9 0 0 1 9 2
21 7 13 9 0 1 7 9 9 9 0 1 9 10 1 9 13 12 12 9 0 2
23 7 3 7 13 8 1 9 1 10 9 7 9 2 7 14 9 9 14 13 9 1 0 2
32 7 13 9 0 1 7 9 0 0 14 13 1 8 9 9 1 9 8 8 2 7 15 13 1 9 9 1 9 1 9 0 2
39 7 13 9 9 0 1 9 8 0 1 9 8 8 1 9 7 9 9 2 7 13 9 1 7 10 9 14 13 9 0 1 9 0 1 9 9 8 9 2
33 7 13 8 8 9 0 1 9 8 1 9 0 7 15 2 3 7 13 1 9 0 7 14 9 9 8 0 15 9 9 9 2 2
50 14 7 9 9 0 13 9 9 9 1 9 0 1 9 10 1 9 2 7 14 13 9 9 9 1 9 0 9 9 7 9 7 9 7 9 0 7 9 7 9 7 9 9 9 1 9 9 1 9 2
25 7 13 1 9 9 1 9 0 1 9 10 9 8 8 1 9 0 13 9 9 0 1 9 0 2
3 2 13 2
20 9 0 2 9 0 13 1 9 8 8 8 8 8 9 2 9 0 7 0 2
60 9 0 2 9 9 13 1 9 8 8 8 8 8 9 2 9 0 7 0 2 7 13 8 8 8 0 1 9 8 9 7 9 8 2 8 13 10 9 1 9 9 13 9 15 1 12 12 9 2 12 12 9 0 2 13 1 15 9 0 2
28 7 13 9 9 1 7 9 8 9 9 9 14 13 1 1 12 12 9 1 15 12 12 1 9 9 1 0 2
24 7 13 9 7 9 0 14 13 1 9 1 0 9 15 12 12 9 1 9 9 8 1 9 2
23 7 13 8 7 8 13 7 13 1 9 1 9 13 1 12 7 12 1 12 1 10 9 2
34 7 13 2 14 13 8 8 8 9 1 0 9 8 8 8 0 1 7 8 2 7 14 13 9 1 9 1 9 0 1 10 9 2 2
19 7 14 13 8 9 9 1 9 9 9 1 1 12 9 1 1 9 0 2
47 7 13 1 9 1 8 7 9 0 2 7 8 13 1 0 9 1 9 9 0 8 8 15 9 9 8 8 9 9 3 2 8 1 9 13 8 7 14 13 8 8 9 8 0 8 2 2
31 14 7 9 9 0 13 7 9 9 0 15 14 13 1 15 9 14 13 8 1 0 1 15 13 15 9 9 7 9 0 2
48 7 13 9 0 8 8 9 2 8 8 0 1 9 7 7 1 9 0 7 8 8 9 0 9 1 0 2 7 14 13 8 8 1 9 9 0 7 3 9 0 8 8 8 1 9 0 2 2
5 8 13 1 12 9
3 8 12 9
27 13 9 9 0 7 8 13 9 1 12 9 13 14 13 1 9 0 0 7 1 9 15 9 1 9 0 2
49 7 13 9 1 9 1 9 9 0 9 15 7 15 13 9 9 1 9 13 1 9 0 7 7 15 13 9 15 1 15 1 9 8 1 9 8 0 8 9 1 9 15 1 9 8 1 8 8 2
28 7 1 9 13 8 8 9 9 0 1 2 9 0 1 9 15 1 9 0 7 9 0 1 9 9 0 2 2
29 7 13 9 7 12 7 12 9 14 13 1 12 9 7 13 9 15 9 15 1 9 0 1 9 9 9 9 0 2
35 7 14 13 1 15 7 1 9 15 9 7 9 7 15 9 15 13 9 1 9 7 13 9 1 9 9 0 0 7 9 0 0 1 9 2
37 7 13 9 0 1 15 1 7 9 0 13 1 9 15 1 9 9 1 9 0 1 9 1 9 1 9 0 7 7 15 13 9 15 1 9 0 2
31 7 13 7 15 13 1 15 9 7 9 7 15 9 1 9 0 1 9 15 7 13 9 15 9 9 1 9 1 10 9 2
10 9 13 8 8 9 1 9 9 1 9
3 9 12 9
76 13 9 8 9 8 8 9 8 8 8 8 9 1 9 1 9 9 0 1 9 1 9 0 1 9 0 1 9 1 9 9 9 8 13 3 0 2 13 8 1 9 0 13 1 15 9 9 8 8 7 9 9 0 7 9 0 8 8 1 9 9 0 2 8 2 1 8 9 0 1 9 9 8 3 9 2
43 7 13 7 9 13 8 8 9 13 1 9 2 8 8 2 8 8 8 8 9 1 9 9 0 7 9 9 0 1 9 1 15 9 1 7 10 9 14 13 1 9 0 2
33 7 13 8 7 9 1 9 9 1 9 1 9 0 2 15 15 14 9 1 10 13 15 9 0 1 9 0 1 8 8 8 2 2
54 7 13 8 1 9 9 7 1 9 9 0 7 0 7 0 7 9 15 0 7 15 13 1 9 9 7 9 7 7 15 14 13 13 9 0 1 9 2 7 3 9 13 0 1 9 1 9 12 7 9 12 9 2 2
27 7 13 7 9 0 9 14 13 1 9 1 9 8 0 0 1 9 10 13 8 8 9 9 1 9 9 2
49 7 13 9 9 0 14 13 1 9 15 9 15 13 1 9 8 0 1 9 8 15 13 8 8 9 9 1 9 9 0 7 13 8 10 9 1 9 9 1 9 9 0 7 9 9 0 1 9 2
28 7 13 7 8 13 14 13 1 9 0 1 9 15 1 12 12 9 8 8 1 15 8 8 9 8 9 0 2
7 9 9 9 0 13 1 9
3 9 12 9
31 13 9 9 9 0 9 8 8 8 7 9 9 0 0 1 9 8 0 0 8 8 1 3 9 1 9 1 9 13 9 2
38 7 13 9 9 0 2 8 2 7 9 9 0 1 9 13 1 9 9 1 9 9 9 0 13 1 9 9 0 8 8 8 9 1 9 9 8 8 2
32 7 1 0 7 13 8 8 15 13 1 9 0 1 9 9 9 1 9 1 0 0 9 1 8 8 8 8 9 0 1 9 2
45 13 7 8 13 9 9 1 9 9 9 1 9 9 7 13 9 0 8 8 9 15 1 9 15 1 0 1 9 0 1 9 1 9 8 1 9 9 0 1 9 7 9 9 9 2
37 7 13 1 9 8 8 9 9 9 1 9 9 0 8 8 8 7 9 8 0 1 9 0 8 8 8 8 8 8 7 9 1 9 1 9 0 2
11 9 9 1 8 8 8 1 9 8 1 9
3 9 12 9
46 13 9 9 0 8 8 8 8 9 8 9 0 1 9 15 9 8 8 1 9 9 1 9 1 9 9 9 8 8 1 9 9 9 0 8 8 1 9 1 8 9 8 8 8 0 2
69 7 13 9 9 9 0 0 7 8 13 8 9 9 15 13 15 8 1 9 9 9 8 8 2 8 8 2 1 8 1 9 0 1 9 7 13 9 0 1 9 15 0 1 9 9 2 9 0 15 13 15 9 0 8 8 9 1 9 8 8 9 0 0 9 12 1 9 8 2
38 7 13 8 1 9 1 9 9 9 0 9 8 9 1 8 8 1 9 15 1 9 0 7 9 0 13 9 1 9 9 0 8 9 1 8 9 9 2
19 7 13 8 9 9 0 0 1 9 9 0 1 9 8 8 9 9 0 2
37 7 13 8 1 9 0 0 1 9 9 0 8 8 1 8 8 1 8 1 9 0 7 2 1 9 0 9 9 1 9 7 9 8 8 0 2 2
