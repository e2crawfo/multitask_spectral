27251 17
2 9 0
10 9 9 13 3 0 7 0 9 9 2
15 3 0 9 16 3 2 16 9 13 15 3 3 9 9 2
6 3 0 9 3 13 2
12 16 13 2 0 11 13 9 2 15 13 3 2
9 16 11 9 13 3 3 2 7 2
2 9 0
8 9 9 13 15 3 0 9 2
8 13 15 9 7 0 9 9 2
12 3 15 13 15 9 13 15 9 16 11 9 2
1 9
13 11 9 13 3 3 0 2 16 9 13 15 13 2
12 9 15 13 9 3 7 13 13 9 9 1 2
4 9 13 0 2
21 15 13 9 9 9 15 9 9 15 2 13 13 15 9 7 9 1 13 15 9 2
1 11
7 0 9 13 3 0 9 2
18 16 9 13 3 3 13 3 9 7 9 2 13 3 0 9 0 13 2
12 9 11 11 4 9 13 3 9 2 3 9 2
27 3 3 9 9 13 13 3 9 2 3 3 9 4 13 9 3 2 7 3 4 13 9 2 15 9 13 2
5 9 13 3 0 2
13 0 2 16 9 4 13 0 0 7 3 13 9 2
15 3 11 11 13 9 0 9 7 11 11 0 9 13 9 2
25 9 13 3 15 2 15 9 13 3 2 7 15 13 15 2 16 9 11 4 13 13 9 3 9 2
19 3 3 9 13 0 9 2 7 9 13 3 15 9 9 3 12 9 9 2
17 9 3 3 11 11 13 15 0 9 2 15 13 13 15 9 9 2
6 0 13 3 9 9 2
13 9 0 9 4 3 13 13 15 9 0 9 9 2
12 3 0 9 13 9 9 13 3 9 13 9 2
19 3 16 9 9 13 13 9 13 0 9 2 9 4 13 15 0 0 9 2
16 9 15 13 13 9 3 9 9 2 15 13 13 3 0 9 2
14 8 8 4 13 8 2 13 0 9 13 15 16 0 2
1 9
9 3 4 13 13 9 1 9 9 2
8 3 15 13 0 16 0 9 2
4 0 15 13 2
13 13 9 9 2 15 13 9 9 15 11 9 9 2
7 13 9 3 7 13 9 2
20 15 13 3 0 7 15 4 3 13 9 9 2 15 4 13 9 13 15 9 2
32 3 9 4 13 9 9 7 13 2 16 15 4 13 9 2 7 15 13 15 9 12 9 9 2 3 11 4 13 15 0 9 2
11 15 13 13 2 4 13 13 15 3 3 2
14 13 9 9 7 15 13 3 3 2 16 9 13 13 2
4 3 3 13 2
18 13 2 13 9 3 3 15 0 9 2 3 16 9 13 0 9 9 2
20 9 2 3 3 3 7 3 3 3 13 2 3 9 13 9 4 13 0 13 2
10 13 9 3 13 15 9 7 0 9 2
9 16 9 13 9 3 0 9 15 2
16 3 2 3 15 9 2 16 13 9 3 2 13 3 13 15 2
4 15 15 13 2
6 15 15 3 3 13 2
31 13 3 3 13 15 2 4 0 9 13 0 9 2 15 13 15 9 9 7 13 15 0 9 2 15 0 9 13 3 13 2
3 0 9 2
41 13 15 13 2 13 13 13 9 2 15 13 13 7 13 9 2 13 15 1 2 16 9 13 9 9 3 3 2 16 9 13 13 0 9 3 16 9 13 9 0 2
5 0 9 15 13 2
11 13 3 9 9 7 3 13 15 2 3 2
9 3 9 9 9 13 9 0 9 2
8 3 3 15 13 9 9 1 2
8 9 13 9 7 13 16 3 2
4 15 13 13 2
2 0 9
6 13 0 9 11 9 2
16 0 2 16 9 13 13 9 13 2 7 3 9 13 3 0 2
4 3 13 9 2
13 3 0 2 7 15 9 9 13 3 12 9 0 2
12 3 15 13 3 0 2 7 3 9 13 13 2
5 11 4 13 3 2
4 9 13 3 2
7 9 13 3 3 0 9 2
1 3
5 3 13 3 9 2
24 9 13 3 9 9 7 16 15 4 13 3 2 4 3 4 13 3 3 7 13 7 13 11 2
4 13 3 3 2
6 9 13 3 0 13 2
19 9 13 0 7 9 2 13 9 12 9 2 13 9 9 7 13 9 9 2
12 13 3 13 9 0 2 7 9 13 3 0 2
7 13 3 7 13 9 9 2
5 13 9 0 9 2
4 13 13 11 2
4 9 13 12 2
8 3 13 9 7 13 9 9 2
16 13 12 9 7 13 9 9 9 9 13 0 9 9 9 9 2
13 13 13 9 9 7 13 0 9 9 13 9 9 2
6 13 13 9 9 3 2
9 15 13 9 9 7 13 3 9 2
6 9 13 3 9 1 2
1 9
9 13 9 1 9 7 9 13 9 2
15 15 13 15 2 3 15 9 1 9 13 13 9 1 9 2
5 13 9 13 9 2
12 9 2 0 7 0 2 15 3 13 2 13 2
14 15 13 13 9 0 9 2 15 1 9 13 13 3 2
11 3 9 13 2 16 9 13 15 3 3 2
4 12 9 1 2
12 15 1 16 9 3 13 9 13 3 0 15 2
5 15 9 9 1 2
11 3 3 13 9 3 16 15 15 13 13 2
26 13 2 16 16 15 13 4 13 9 3 3 9 12 9 9 2 13 15 13 2 13 15 13 15 1 2
7 9 9 2 3 7 3 2
16 15 2 15 0 9 4 13 13 15 2 16 9 13 0 9 2
4 13 15 0 2
10 3 9 9 13 2 3 15 9 13 2
18 3 3 15 4 13 9 3 0 9 2 15 9 15 13 4 3 13 2
1 9
3 13 9 2
26 2 13 2 16 9 13 9 13 9 3 3 9 3 9 9 1 2 16 15 13 13 13 0 9 1 2
26 13 0 7 13 3 9 5 2 16 4 13 15 9 2 15 13 9 9 13 13 3 15 9 1 2 2
5 15 15 13 3 2
1 9
6 15 9 13 13 9 2
10 9 9 13 9 7 13 9 15 1 2
12 0 13 15 0 9 7 3 13 0 9 3 2
11 13 2 13 15 4 13 3 0 9 9 2
15 0 9 3 4 13 3 3 9 2 13 9 4 3 13 2
5 7 9 7 9 2
17 13 16 12 9 13 9 13 3 15 2 16 9 4 13 3 3 2
19 3 13 0 9 3 13 7 9 13 13 9 2 15 0 9 13 13 15 2
6 3 9 13 3 0 2
14 13 13 0 9 0 9 3 2 16 9 3 13 3 2
12 13 9 9 2 15 9 4 13 3 9 9 2
12 3 13 2 3 13 13 9 9 0 9 9 2
9 3 3 13 3 0 13 0 9 2
9 7 3 3 3 3 13 13 0 2
19 9 13 9 7 9 2 15 3 3 9 4 13 15 3 9 2 9 9 2
17 16 15 13 2 13 13 2 13 13 2 4 13 2 15 15 13 2
14 7 3 4 3 13 9 9 2 7 13 9 0 9 2
9 9 9 13 3 7 9 9 9 2
10 9 13 3 16 3 13 7 13 13 2
19 12 9 4 13 0 0 9 9 7 12 9 9 2 7 3 13 4 13 2
16 3 4 13 13 9 13 0 9 9 7 13 3 15 0 9 2
7 7 16 3 13 3 0 2
12 3 13 9 3 2 13 9 7 13 15 0 2
14 3 0 0 9 1 13 9 1 0 9 9 15 9 2
18 9 13 9 9 0 9 2 15 13 0 9 7 9 13 0 0 9 2
16 4 3 13 9 2 7 15 13 13 3 0 2 13 0 3 2
16 15 13 13 3 3 3 13 7 9 13 3 13 3 13 9 2
8 3 13 3 11 11 0 9 2
8 7 3 13 3 3 3 9 2
4 7 0 9 2
7 3 4 13 13 9 9 2
14 3 0 9 1 9 13 13 9 11 7 3 3 11 2
2 0 2
9 9 9 9 4 13 13 9 9 2
10 13 2 16 9 11 4 13 15 9 2
3 9 1 0
5 9 15 9 1 2
15 1 0 9 2 15 9 13 9 9 9 2 15 9 13 2
9 2 9 2 15 15 3 13 9 2
6 13 9 3 13 9 2
12 16 13 2 16 3 15 9 2 15 9 13 2
7 2 13 3 3 9 9 2
7 13 0 9 3 0 2 2
3 9 1 0
7 1 9 0 9 13 3 2
9 2 9 2 15 13 15 3 9 2
18 2 6 2 13 7 13 9 2 3 9 13 3 0 13 9 9 1 2
10 13 3 15 9 13 9 9 9 9 2
3 9 13 2
7 9 4 3 13 15 13 2
5 15 13 3 2 0
8 2 9 2 13 15 13 9 2
5 13 13 9 9 2
5 9 11 7 13 9
7 0 9 2 9 7 9 2
15 3 3 2 15 9 13 0 2 16 9 13 3 0 9 2
13 3 13 3 4 13 2 16 4 13 15 13 9 2
18 15 13 9 15 2 16 0 0 7 0 9 1 15 4 13 9 9 2
16 15 3 4 13 9 9 2 7 3 15 13 3 0 13 2 5
11 13 3 0 9 2 15 13 0 0 9 2
13 13 15 11 9 15 9 2 15 1 0 15 13 2
17 9 13 15 15 9 3 2 16 0 0 9 13 0 13 3 2 5
7 15 9 13 3 3 0 2
20 4 3 13 9 0 9 2 15 3 13 9 1 2 13 7 9 13 3 0 2
17 15 13 3 0 9 0 9 2 16 15 13 3 0 7 3 0 2
15 16 15 9 13 0 7 0 2 13 9 13 9 13 9 2
13 13 9 15 9 2 15 4 13 9 3 12 9 2
16 15 9 15 13 2 16 0 9 13 3 0 13 0 0 9 2
23 9 15 9 13 11 11 13 9 3 0 9 2 9 13 9 13 3 9 0 9 13 9 2
13 9 4 13 3 7 15 4 13 11 11 9 2 5
14 13 3 9 9 11 11 0 9 2 9 8 8 2 2
15 4 3 13 3 11 9 2 3 3 15 13 9 9 13 2
16 0 9 13 15 9 1 7 13 13 2 13 15 15 9 2 5
16 0 13 9 13 15 3 0 2 7 0 9 9 15 13 13 2
13 15 1 15 9 13 0 9 7 9 1 3 3 2
27 9 13 0 9 15 2 13 15 13 0 9 2 7 9 13 0 13 3 7 15 4 0 9 13 3 9 2
7 3 2 13 13 15 2 5
20 13 3 3 3 2 3 3 2 9 2 16 4 3 4 13 15 9 1 9 2
13 9 2 15 13 3 9 13 13 3 15 0 9 2
10 13 0 9 3 9 13 7 9 13 2
19 0 9 13 3 0 7 16 9 15 9 13 13 3 3 2 13 9 9 2
7 13 9 7 13 3 13 2
6 0 9 9 13 2 5
13 13 3 15 9 2 15 9 1 13 13 9 1 2
11 0 1 9 13 0 9 7 9 7 9 2
9 3 13 3 9 13 13 9 9 2
8 3 15 0 9 13 9 1 2
14 7 3 13 3 15 3 0 9 2 3 0 9 9 2
7 7 3 9 2 6 2 5
11 13 3 9 2 16 9 13 13 15 9 2
16 0 9 13 9 1 3 0 9 9 11 11 11 11 11 11 2
13 13 3 3 9 7 15 13 3 15 0 9 2 5
14 9 13 3 2 15 0 9 13 9 7 9 13 0 2
7 9 9 9 4 13 3 2
14 13 3 15 9 2 16 9 9 7 15 9 13 3 2
7 3 15 13 9 9 9 2
12 9 13 3 3 9 1 2 3 13 13 3 2
12 9 9 7 9 13 3 3 15 0 9 1 2
11 13 9 13 9 2 4 13 9 9 2 5
6 3 15 3 13 3 2
12 13 15 3 3 0 16 9 2 3 9 13 2
6 9 9 7 0 9 2
4 11 5 9 9
7 3 4 13 15 9 3 2
6 9 15 13 3 13 2
11 13 15 9 2 16 0 9 13 3 9 2
7 6 2 15 15 13 13 2
5 13 3 0 2 5
15 15 9 13 3 13 2 15 9 4 3 13 3 9 9 2
10 15 13 15 2 16 13 9 11 9 2
17 11 4 3 13 8 8 0 9 2 3 4 15 9 13 9 13 2
6 15 13 3 12 9 2
15 9 13 3 9 11 2 15 13 3 3 13 13 3 9 2
7 6 2 3 0 9 2 5
14 13 3 2 16 9 13 3 3 0 9 7 3 0 2
19 16 9 13 9 7 9 13 13 9 2 13 11 1 9 7 13 9 15 2
17 15 9 13 13 9 9 9 7 13 9 2 7 3 15 13 13 2
15 7 15 3 13 2 16 0 12 9 9 9 4 13 15 2
8 13 3 11 0 9 9 9 2
8 3 0 9 13 9 9 3 2
9 9 13 9 3 13 15 0 9 2
4 13 9 2 5
11 1 0 9 9 11 13 15 9 9 1 2
10 13 0 9 9 7 4 15 3 13 2
14 3 13 3 11 11 9 2 13 3 13 15 9 2 5
13 3 13 13 15 9 9 2 7 3 15 13 15 2
10 3 3 0 15 9 13 3 3 13 2
10 9 9 13 0 9 13 3 0 9 2
13 13 15 9 3 2 7 13 13 15 3 3 9 2
2 6 2
12 9 9 7 9 7 9 1 13 9 13 9 2
12 3 13 0 9 2 15 1 13 3 0 9 2
15 4 13 11 3 0 3 0 9 7 15 13 3 0 9 2
8 0 13 6 13 3 3 2 5
15 9 13 3 3 3 0 3 13 3 4 13 15 1 9 2
13 3 9 13 3 13 3 0 2 0 9 13 3 2
16 11 13 3 3 0 9 2 16 0 0 9 9 13 3 9 2
16 6 2 0 9 13 12 9 2 15 13 13 13 9 13 9 2
5 3 2 11 2 5
13 13 3 15 0 9 1 3 0 9 7 0 9 2
16 15 9 9 13 15 0 9 0 2 7 15 13 3 13 9 2
7 13 4 13 0 9 9 2
10 3 13 0 9 2 13 15 9 2 5
10 3 9 4 13 0 9 3 0 9 2
11 7 3 0 9 2 7 15 15 15 9 2
10 9 13 0 9 2 13 9 3 3 2
10 7 3 0 0 2 7 0 9 2 5
22 9 13 3 0 9 7 13 11 0 9 2 11 5 9 2 11 2 11 7 15 2 2
9 11 13 11 7 13 3 0 9 2
4 7 3 13 2
12 3 13 15 9 2 16 15 9 13 3 0 2
5 15 0 4 13 2
11 13 3 9 13 15 15 9 2 11 2 5
9 0 9 13 11 13 2 9 2 2
14 9 13 3 15 0 9 2 15 13 9 9 0 9 2
13 13 13 9 9 0 9 7 3 9 13 9 9 2
25 11 13 13 15 9 1 2 16 9 13 0 2 7 15 13 13 2 7 13 11 9 13 0 9 2
7 9 2 13 15 13 9 2
14 11 3 13 9 13 15 9 15 2 3 3 9 13 2
6 3 9 13 15 9 2
9 3 7 13 3 11 15 0 9 2
15 3 3 3 0 15 3 13 9 16 15 3 13 9 2 5
13 9 13 13 0 9 2 16 9 13 0 9 15 2
6 7 6 13 7 13 2
14 11 13 0 9 7 11 13 13 3 16 13 0 2 5
9 0 9 9 2 16 3 0 13 2
19 8 8 13 3 9 13 9 9 15 9 2 16 4 13 13 15 3 9 2
10 3 13 3 9 7 9 9 7 9 2
16 13 13 0 9 3 0 9 7 4 3 3 15 9 13 2 5
15 15 9 1 13 3 3 9 2 16 15 13 3 3 9 2
2 6 2
26 13 2 13 13 15 0 16 15 2 16 15 13 15 2 16 3 4 13 2 13 13 9 9 1 2 5
9 15 13 3 3 15 9 15 9 2
28 15 13 3 0 2 16 0 9 9 13 3 15 0 9 1 7 16 9 13 15 2 13 13 3 0 9 13 2
13 13 9 13 9 2 3 15 9 13 3 3 9 2
15 15 9 9 13 3 13 9 9 2 16 13 3 13 3 2
26 9 13 3 3 9 2 9 2 9 7 9 2 7 3 3 13 13 13 9 3 13 2 16 3 13 2
8 15 13 13 9 3 3 3 2
8 15 13 2 16 13 12 9 2
2 3 2
13 9 9 13 3 0 2 16 13 13 9 0 9 2
16 15 0 9 1 13 13 2 15 9 13 3 0 0 9 9 2
14 9 15 0 7 0 9 2 3 13 3 0 9 3 2
1 9
12 9 7 3 0 9 0 9 4 13 0 9 2
10 15 13 13 13 3 16 13 7 13 2
22 3 15 13 3 0 2 16 9 13 0 2 7 3 15 4 13 0 9 7 9 3 2
19 0 9 2 16 13 12 9 2 9 2 9 9 9 2 0 9 13 13 2
17 3 4 3 13 15 1 9 2 12 9 7 3 3 15 0 9 2
9 4 13 15 9 3 0 9 9 2
23 15 13 0 9 2 16 1 0 9 2 13 3 4 13 3 9 7 13 0 0 9 2 5
4 13 13 0 2
10 9 13 3 9 2 9 7 3 15 2
5 0 13 11 9 2
13 3 13 3 0 9 13 2 13 13 11 3 15 2
22 9 13 3 12 9 2 12 9 7 12 9 2 15 15 13 3 3 0 0 7 11 2
16 13 13 9 9 3 2 7 13 3 13 3 15 3 13 9 2
12 9 13 0 2 7 13 3 13 15 3 3 2
10 13 9 3 9 9 12 9 9 9 2
5 13 9 3 2 5
12 9 13 3 11 7 9 15 13 0 7 0 2
11 15 13 9 7 15 9 13 3 13 0 2
8 13 15 3 0 9 15 9 2
12 9 13 3 3 2 16 15 13 3 9 13 2
8 15 13 0 0 7 15 0 2
13 13 9 2 3 3 0 9 13 9 3 3 9 2
14 9 3 2 16 15 9 13 13 9 13 3 15 9 2
18 13 3 0 3 9 2 16 7 11 7 11 13 15 1 9 0 9 2
8 15 15 13 2 9 2 2 5
11 13 13 0 9 2 7 13 0 9 9 2
6 7 13 9 9 9 2
13 16 3 13 2 16 13 3 2 7 13 3 9 2
7 3 2 13 15 13 3 2
7 13 3 12 9 9 1 2
5 9 13 0 9 2
13 11 13 3 9 2 16 13 3 9 9 0 9 2
13 9 13 15 2 16 4 13 9 9 3 3 9 2
6 9 15 3 15 9 2
12 0 15 9 13 13 2 7 3 0 3 2 5
11 15 9 13 0 9 7 9 3 0 9 2
9 9 7 9 0 9 13 15 9 2
20 9 9 13 3 0 2 16 15 13 0 9 1 16 16 15 13 0 9 9 2
3 13 3 2
17 15 1 2 16 13 11 9 2 15 9 15 13 9 4 13 9 2
14 3 13 0 9 2 16 15 9 4 13 15 0 9 2
16 13 3 3 15 2 16 9 4 13 9 7 3 15 4 13 2
12 9 1 4 3 13 3 9 7 15 9 11 2
11 13 9 3 3 2 16 13 13 9 2 5
3 0 9 5
16 4 13 15 15 2 16 3 13 9 13 0 9 3 0 9 2
6 7 3 4 13 2 5
15 4 13 12 0 9 9 7 15 9 5 9 13 9 9 2
19 15 0 9 2 15 3 15 9 1 13 4 13 13 13 2 13 13 3 2
5 3 3 13 9 2
19 0 9 4 13 15 9 2 16 15 9 13 9 1 13 3 9 0 9 2
28 9 7 9 3 3 13 9 2 9 9 2 9 9 7 9 9 13 15 9 7 9 15 2 16 9 13 13 2
12 3 3 13 7 15 13 3 0 7 0 13 2
21 3 0 9 9 2 0 7 0 2 13 9 9 3 2 16 13 9 0 9 9 2
9 9 3 0 9 13 9 7 9 2
10 9 13 13 3 2 13 15 13 3 2
17 9 2 15 13 3 13 7 15 13 3 13 13 9 1 0 9 2
16 15 13 15 13 9 0 9 2 15 13 0 13 7 0 13 2
12 9 9 9 7 9 13 0 7 13 9 9 2
21 9 2 9 9 7 0 9 9 1 13 15 9 13 0 9 7 13 15 9 9 2
8 0 9 13 9 0 3 9 2
19 13 3 0 13 12 9 3 13 3 13 9 3 7 13 9 9 0 9 2
16 9 2 15 9 13 9 2 3 16 5 2 13 15 3 2 2
18 3 4 9 1 13 2 2 15 9 13 9 13 9 9 5 2 2 5
3 13 9 2
3 13 3 2
16 16 13 4 13 9 7 3 13 15 0 9 2 13 13 15 2
4 0 9 13 2
18 3 9 15 1 13 3 0 9 15 9 2 15 9 4 3 13 2 5
4 0 9 2 5
3 9 9 2
19 9 13 2 9 13 3 0 9 7 9 13 3 0 16 15 9 4 13 2
11 3 16 13 13 0 9 2 13 13 9 2
16 9 2 9 7 9 13 13 16 0 9 2 15 13 9 9 2
18 15 9 13 4 13 15 9 7 9 0 9 3 2 16 13 0 9 2
9 9 13 9 0 9 13 9 9 2
10 9 13 3 13 7 0 9 13 13 2
12 9 13 4 13 2 16 13 3 7 13 3 2
12 3 4 0 9 13 9 7 13 0 9 2 5
9 15 9 13 0 7 3 0 9 2
9 3 9 13 3 0 16 0 9 2
6 3 13 0 9 13 2
7 13 9 13 9 9 15 2
12 3 3 9 7 9 9 9 4 13 3 3 2
14 13 15 2 16 13 13 3 15 0 9 9 9 13 2
26 9 13 0 9 2 9 13 13 7 13 9 2 9 13 3 0 9 2 9 13 3 9 3 7 3 2
20 7 9 9 9 13 9 2 16 0 9 13 13 1 9 0 2 9 13 9 2
16 2 3 3 2 9 13 3 9 2 15 9 15 7 3 13 2
21 13 7 13 15 9 15 2 3 15 13 9 2 9 7 9 13 15 15 9 13 2
16 13 9 2 15 13 0 9 2 7 13 2 13 4 13 9 2
7 15 13 0 9 0 9 2
14 9 13 15 2 16 15 4 3 13 9 7 13 13 2
3 13 0 2
3 13 9 2
3 13 3 2
3 13 3 2
5 13 7 13 3 2
5 13 7 13 3 2
17 16 13 15 2 9 7 13 3 15 12 2 4 13 15 3 13 2
8 15 16 13 9 9 3 3 2
8 9 9 13 13 15 0 2 5
8 9 7 9 13 9 15 2 5
6 0 9 12 2 2 2
16 9 4 13 2 9 13 3 3 7 0 2 0 9 3 2 5
8 3 13 3 2 3 13 9 2
8 0 13 3 15 9 2 3 2
6 15 15 4 3 13 2
14 4 13 2 13 2 3 3 13 7 13 15 9 2 5
7 9 4 13 15 0 9 2
22 11 4 13 0 9 7 9 2 11 13 15 2 15 0 9 13 4 3 13 13 2 5
10 9 13 2 9 9 13 3 0 9 2
14 3 9 13 9 9 2 15 1 15 15 9 13 9 2
8 9 9 13 3 7 13 9 2
8 13 0 13 3 9 1 2 5
10 9 13 9 13 9 2 9 7 9 2
6 15 12 9 13 9 2
19 13 9 13 0 9 2 15 13 4 13 9 2 9 7 9 9 15 9 2
9 0 9 9 13 13 3 15 9 2
5 15 13 3 3 2
19 13 15 15 3 2 3 3 0 15 13 9 2 9 9 7 9 9 13 2
11 3 13 15 9 2 9 2 9 7 9 2
9 13 0 9 2 15 13 9 9 2
8 13 2 16 15 13 9 13 2
7 13 9 2 9 7 9 2
7 15 13 9 9 15 9 2
6 13 9 13 9 9 2
10 15 13 9 2 15 1 15 4 13 2
6 0 0 9 15 2 5
3 9 1 5
6 0 2 9 13 2 5
3 3 9 2
20 9 4 15 9 13 3 2 9 4 13 3 3 7 9 13 9 0 9 2 5
13 3 3 2 15 4 13 0 9 2 15 13 9 2
4 3 9 9 2
10 9 13 9 13 13 9 7 3 3 2
13 3 13 0 9 13 9 2 13 9 7 13 9 2
3 13 3 2
3 13 3 2
9 15 13 15 2 16 13 13 15 2
9 4 3 13 0 9 13 9 1 2
15 3 13 3 13 9 9 2 7 0 2 0 9 9 2 5
12 9 13 12 0 9 2 15 9 7 15 9 2
16 0 13 3 0 9 7 9 3 7 15 1 13 13 0 9 2
17 7 9 13 13 0 3 9 1 2 16 15 13 13 15 9 2 5
13 15 13 0 9 13 9 9 3 3 9 13 3 2
20 13 3 13 15 2 15 9 13 9 3 3 2 16 15 13 13 3 3 9 2
10 15 13 3 9 2 15 13 3 3 2
13 15 9 13 9 9 0 9 2 16 15 13 13 2
9 9 4 3 13 3 0 9 2 5
12 15 9 4 13 9 9 9 0 9 0 9 2
21 3 2 13 15 9 9 9 3 0 3 7 3 0 9 13 13 15 9 3 3 2
9 3 13 3 9 13 3 7 9 2
15 0 9 13 2 13 9 1 7 13 3 1 0 9 9 2
6 0 9 15 15 2 5
2 0 9
18 16 15 13 9 9 1 3 9 2 13 9 9 3 3 3 13 9 2
23 6 2 9 13 13 2 16 16 3 13 9 15 9 13 0 9 13 2 3 9 15 13 2
10 4 3 13 0 9 2 3 3 2 5
23 9 15 9 13 9 13 0 9 15 2 16 9 7 15 9 4 13 13 3 13 7 13 2
7 15 9 13 15 3 9 2
26 9 9 4 13 7 13 9 13 9 7 9 7 0 2 7 9 13 15 15 0 2 15 4 15 13 2
16 3 3 13 3 15 2 15 13 13 13 3 15 2 7 15 2
5 9 13 16 9 2
9 15 3 13 2 15 13 9 3 2
4 9 13 9 2
15 15 15 13 13 13 0 9 2 4 13 0 13 3 9 2
9 9 0 9 13 13 15 0 9 2
9 9 13 15 2 3 13 15 15 2
6 13 13 13 3 15 2
14 16 9 4 13 7 9 13 2 13 9 13 0 9 2
13 0 9 13 13 0 9 15 9 2 7 15 9 2
13 15 15 13 0 9 2 13 0 7 13 3 0 2
12 9 1 13 0 9 13 9 9 3 0 9 2
10 9 9 13 13 13 3 0 9 2 5
22 15 1 2 7 3 1 15 2 4 13 9 0 2 0 7 0 9 13 0 13 9 2
9 0 2 0 13 9 13 3 0 2
18 15 9 4 13 9 2 7 16 15 9 13 2 13 15 0 13 3 2
6 9 13 0 3 9 2
14 16 15 13 0 9 2 13 9 9 3 3 0 9 2
11 3 3 13 3 3 2 16 15 13 0 2
11 9 7 15 9 9 9 7 9 13 0 2
7 3 0 9 4 13 9 2
15 9 9 1 2 9 2 9 7 0 9 13 3 9 9 2
12 15 9 9 13 9 2 0 9 7 9 2 5
12 3 0 0 2 7 3 15 15 15 9 13 2
10 9 2 15 13 9 2 13 0 9 2
10 9 13 0 9 2 7 15 13 15 2
26 16 13 13 0 9 12 9 2 15 13 9 13 2 13 15 9 2 3 13 9 7 3 13 9 2 5
5 11 9 13 3 2
3 9 2 5
11 3 13 15 9 9 9 13 9 12 9 2
7 13 15 3 7 13 9 2
10 3 13 9 3 0 9 7 13 9 2
8 13 9 9 7 13 15 3 2
19 9 13 9 9 9 2 9 13 9 2 7 13 0 9 9 7 9 9 2
11 9 13 0 2 16 9 13 13 9 9 2
7 9 1 3 0 9 2 5
5 0 9 15 2 5
1 9
6 11 13 9 9 2 5
13 15 13 15 15 9 9 2 15 15 13 13 13 2
13 3 15 9 13 0 9 2 3 0 9 13 9 2
11 9 7 0 11 13 9 2 15 13 2 5
11 9 4 0 9 13 7 9 9 13 9 2
14 15 9 9 13 3 2 16 0 9 13 9 0 9 2
15 16 15 7 9 13 9 9 2 13 9 13 9 9 1 2
11 3 2 15 15 0 16 12 9 9 2 5
10 9 9 13 13 3 15 0 16 3 2
11 3 3 15 13 9 0 9 9 7 9 2
9 15 1 13 13 3 9 13 9 2
8 9 13 3 13 0 7 0 2
15 3 13 3 13 9 15 9 2 15 9 0 9 15 13 2
9 15 1 2 13 13 9 15 9 2
13 15 1 13 0 9 2 16 15 3 13 13 2 5
4 9 0 9 5
7 0 9 3 13 0 2 5
10 15 13 3 3 2 13 13 3 9 2
10 16 13 0 2 9 13 15 0 9 2
15 16 4 15 1 13 9 2 13 13 9 0 9 3 9 2
9 9 13 3 0 9 16 9 2 5
10 13 9 3 15 9 2 15 9 13 2
18 16 13 3 9 3 0 9 9 7 3 3 9 2 13 0 9 9 2
17 4 3 13 15 0 9 9 7 9 2 3 3 9 4 13 9 2
7 15 15 13 15 9 9 2
18 16 13 9 0 16 15 13 7 13 15 2 13 13 15 15 0 9 2
15 15 2 15 3 13 3 3 13 9 2 13 3 3 3 2
5 13 3 9 0 2
10 4 13 15 2 15 9 1 13 2 5
4 15 0 9 2
15 4 15 13 3 9 13 15 2 3 15 4 13 9 2 2
9 2 15 15 13 13 9 9 2 2
6 2 13 13 9 2 2
13 2 4 15 13 15 9 13 7 15 15 13 2 2
9 15 13 9 15 13 9 0 9 2
12 16 4 13 9 2 3 4 13 0 0 9 2
39 9 2 3 9 2 13 11 2 13 9 0 9 2 2 9 13 3 0 11 11 11 9 15 2 15 9 13 13 9 9 16 9 13 9 2 3 3 9 2
12 9 7 9 4 13 9 9 13 3 9 9 2
16 15 13 15 9 13 9 7 12 0 9 9 2 15 13 9 2
10 15 15 9 7 9 13 9 0 9 2
22 2 16 9 13 9 13 3 9 9 2 15 4 13 15 2 16 13 13 9 0 9 2
9 0 9 13 3 9 3 0 9 2
22 0 9 13 3 9 3 0 7 0 9 2 2 13 3 11 11 9 11 7 11 9 2
10 0 9 13 7 9 7 9 3 0 2
7 3 3 13 15 0 9 2
21 3 13 7 4 13 2 16 0 9 7 9 13 0 2 15 13 9 7 13 0 2
26 2 9 9 13 9 13 15 2 16 9 13 15 13 2 13 13 13 15 9 13 2 7 13 3 0 2
11 9 13 16 9 13 9 2 7 0 9 2
12 16 9 13 9 13 15 2 15 13 0 3 2
28 16 9 9 13 0 9 0 9 7 15 2 13 9 4 13 15 0 2 7 9 13 9 1 2 9 13 3 2
15 16 9 13 3 0 9 13 9 0 2 15 4 13 9 2
22 9 13 3 13 2 13 13 9 3 3 2 15 13 3 13 2 13 3 3 13 9 2
31 13 3 0 2 16 9 13 13 13 9 2 7 3 15 0 9 2 3 3 9 13 9 9 13 9 13 9 15 9 2 2
10 3 13 11 11 9 11 7 11 9 2
8 13 9 13 15 9 0 9 2
13 13 9 13 9 2 16 15 13 0 9 13 9 2
7 13 9 13 9 9 15 2
21 3 13 9 9 9 2 16 2 13 15 9 2 13 15 2 13 15 0 9 2 2
15 9 9 13 3 15 9 2 3 15 13 3 3 0 9 2
3 3 15 2
32 13 15 15 2 15 13 15 15 13 7 13 13 15 2 16 13 13 0 2 15 13 15 0 2 13 13 13 15 3 7 3 2
27 13 15 1 9 13 2 0 9 3 13 2 7 0 9 9 13 2 16 13 13 13 15 15 9 7 9 2
21 15 4 3 3 13 2 16 9 2 15 9 7 9 13 0 13 2 3 9 1 2
25 3 3 15 9 13 13 2 15 13 0 2 13 15 13 15 13 2 13 13 9 2 0 13 2 2
32 3 3 15 9 13 2 3 2 15 13 16 9 2 13 13 15 9 7 15 15 9 2 15 13 3 0 2 13 3 13 2 2
8 3 13 13 9 3 3 0 2
11 9 13 3 2 15 1 9 13 0 9 2
18 9 13 3 3 15 2 15 13 13 13 3 2 16 9 13 9 0 2
10 3 13 13 15 15 9 2 15 13 2
12 3 13 13 9 9 9 2 16 13 13 9 2
13 3 13 0 7 13 2 16 15 13 3 3 3 2
15 15 15 9 7 0 0 9 13 3 0 7 3 0 9 2
8 9 1 9 13 3 9 9 2
3 3 13 2
3 15 13 2
18 13 9 2 16 15 13 2 0 2 2 0 2 0 2 0 2 0 2
12 7 3 2 16 13 13 3 9 7 9 1 2
14 9 4 13 9 13 0 9 2 13 11 11 15 9 2
14 15 13 2 2 9 13 15 0 7 0 9 9 9 2
14 9 13 9 9 13 0 9 2 2 13 13 15 0 2
17 16 15 13 2 0 13 3 2 15 13 13 7 13 15 3 2 2
10 9 13 13 2 16 15 4 13 0 2
11 15 4 3 13 3 9 2 3 7 3 2
6 13 13 0 7 0 2
14 15 9 4 13 3 3 2 13 15 13 13 0 9 2
10 9 4 13 9 2 9 7 9 2 2
7 15 3 0 9 3 13 2
23 15 4 3 13 12 7 12 9 2 7 9 13 3 15 9 2 16 9 9 13 3 9 2
33 16 9 13 13 0 2 0 2 0 2 3 0 16 9 2 3 2 15 13 13 15 7 13 15 2 16 13 13 3 0 16 9 2
39 16 9 13 13 13 9 9 7 13 15 2 16 15 13 3 0 2 0 7 0 16 9 2 3 9 9 13 7 15 9 13 13 2 7 15 9 4 13 2
19 0 9 13 13 3 13 15 3 2 13 13 9 2 13 3 13 15 13 2
40 13 0 13 13 2 16 9 9 2 16 13 3 13 2 13 13 3 0 2 13 13 13 9 2 13 13 13 9 2 9 13 13 15 3 2 13 9 7 9 2
11 11 11 13 3 2 2 3 9 13 9 2
20 15 4 3 13 0 9 2 7 0 9 13 9 13 9 2 9 7 9 9 2
6 0 9 4 13 3 2
11 3 9 9 13 9 7 15 9 13 9 2
9 15 13 3 9 7 9 9 2 2
15 4 13 9 15 2 13 4 3 13 0 2 0 7 0 2
15 3 13 2 7 9 4 3 3 13 0 9 3 15 9 2
29 16 13 13 7 13 9 3 2 16 15 13 9 9 2 3 4 13 3 3 2 16 13 13 13 9 3 0 9 2
10 3 15 4 3 13 13 3 0 3 2
11 9 7 15 13 9 13 15 9 0 9 2
18 16 9 2 9 7 0 9 13 15 15 9 2 13 15 15 15 9 2
16 4 13 15 2 13 9 13 0 2 16 9 9 13 13 0 2
3 9 13 9
13 11 13 3 3 3 9 3 3 13 9 7 9 2
26 3 13 11 7 11 2 15 1 9 13 9 3 11 11 11 9 7 15 9 9 13 13 11 11 11 2
40 3 9 9 2 15 3 13 3 12 9 9 2 1 13 0 13 3 0 9 2 7 13 3 3 0 9 2 13 9 2 15 15 13 13 9 2 15 9 13 2
6 9 13 3 11 11 2
17 9 13 0 15 2 16 9 4 13 13 15 9 2 8 8 2 2
13 15 1 9 9 13 13 0 9 2 8 8 2 2
38 4 15 9 3 3 13 2 16 11 11 13 13 15 0 0 9 7 15 13 9 15 15 0 3 3 13 2 3 11 11 2 7 9 0 9 13 9 2
13 9 11 13 0 9 13 3 0 9 11 11 1 2
10 15 13 3 15 13 0 9 13 9 2
14 9 4 3 13 9 9 0 9 13 2 9 7 13 2
4 15 13 13 5
6 11 11 9 13 12 2
3 0 9 2
6 9 13 3 7 3 2
10 13 15 9 9 9 3 15 9 1 2
16 9 13 3 2 7 16 15 15 9 13 2 15 4 13 9 2
11 9 13 13 15 3 15 2 16 9 13 2
13 9 13 9 13 0 2 13 13 15 3 0 9 2
10 11 13 13 3 3 3 16 15 9 2
10 3 9 13 9 9 7 9 13 9 2
19 3 3 4 13 9 12 9 9 13 9 7 15 0 0 9 2 11 2 2
7 9 13 13 3 13 9 2
16 9 3 13 2 7 1 4 3 13 9 2 16 9 13 3 2
19 7 16 15 11 7 9 13 13 15 11 15 13 2 13 9 3 13 3 2
6 3 13 13 9 13 2
23 11 13 11 15 9 9 2 3 13 15 8 0 9 0 2 13 3 9 9 7 9 2 2
12 9 13 11 2 7 15 9 9 7 15 0 2
9 9 13 9 2 13 9 3 3 2
20 13 3 13 11 2 16 13 13 9 3 3 3 16 13 9 9 7 15 9 2
30 15 9 4 4 13 11 3 0 9 2 7 16 15 4 13 11 7 11 2 7 11 2 2 3 15 4 4 13 3 2
18 9 9 9 4 13 13 15 9 2 13 9 2 8 2 2 16 13 2
4 3 9 9 5
8 9 9 2 9 2 9 2 9
17 4 15 9 13 3 0 12 9 2 3 15 9 13 9 13 3 2
13 13 9 2 15 13 0 9 7 9 13 9 9 2
16 13 3 13 9 9 1 2 3 3 9 9 13 3 0 9 2
23 9 13 3 12 9 2 8 2 8 2 8 2 0 8 2 9 2 9 7 0 8 9 2
35 9 9 13 2 9 2 2 9 15 4 13 2 8 15 13 7 15 12 15 9 3 13 9 9 9 9 12 2 7 13 3 13 9 12 2
9 8 7 9 13 3 15 9 1 2
20 15 9 9 1 4 3 13 0 9 2 16 15 4 3 13 3 12 9 1 2
15 3 12 9 13 15 9 2 7 15 13 13 9 9 9 2
11 3 0 13 13 9 12 9 12 9 9 2
10 9 13 13 9 9 12 9 9 9 2
17 15 9 9 13 3 3 0 9 1 2 13 15 4 9 3 13 2
49 9 13 9 13 3 9 9 1 2 13 3 16 11 13 9 2 15 13 9 7 13 9 9 9 2 3 9 13 9 2 2 16 15 9 13 13 9 13 9 2 9 13 9 13 3 9 13 2 2
15 15 9 15 3 2 16 9 4 13 9 7 9 13 9 2
14 9 4 13 12 9 2 15 13 15 9 0 13 9 2
6 0 9 13 0 9 2
4 13 3 3 2
12 15 9 13 12 9 2 7 13 15 3 12 2
5 3 15 13 0 2
6 13 9 13 9 8 2
36 3 13 13 4 13 9 9 15 9 2 7 16 13 9 15 9 7 13 9 15 9 3 7 3 3 0 9 2 13 15 15 13 3 9 13 2
13 0 9 9 13 2 7 13 15 9 4 9 13 2
14 9 13 15 9 12 0 9 2 15 15 13 0 9 2
14 9 15 9 4 13 9 15 2 3 9 13 12 9 2
28 9 12 9 13 7 8 8 2 9 2 7 8 8 2 9 2 0 2 15 15 4 13 0 9 15 12 9 2
10 16 15 13 13 9 2 9 13 13 2
9 15 3 13 7 13 13 13 9 2
9 15 13 9 3 3 3 12 9 2
8 0 9 13 9 15 9 15 2
10 12 0 9 13 9 2 0 9 13 2
6 9 4 13 3 9 2
22 0 9 13 15 0 9 8 8 9 2 16 15 9 15 9 9 4 13 8 8 9 2
9 13 9 3 13 2 16 9 13 2
19 9 4 13 0 9 3 0 9 3 13 2 9 2 3 4 13 2 11 2
25 3 15 4 3 3 13 2 16 13 9 13 3 3 2 16 13 3 12 9 15 7 13 9 9 2
11 9 13 3 3 2 7 3 3 13 9 2
18 15 9 9 9 13 11 2 7 15 13 13 9 9 13 9 9 9 2
15 13 3 9 15 2 15 4 13 13 9 13 3 0 9 2
6 11 11 13 3 3 9
11 11 11 9 0 4 3 13 0 9 1 2
27 16 9 9 3 13 2 13 0 9 9 7 3 13 9 13 3 2 9 13 9 2 2 7 3 13 13 2
17 11 13 3 9 9 7 9 13 9 7 13 9 3 0 9 1 2
7 0 3 3 16 13 3 2
16 3 11 9 9 13 13 9 2 9 9 13 4 13 9 2 2
24 9 13 9 13 9 8 2 5 8 2 5 8 2 5 8 2 15 1 11 11 13 13 3 2
10 16 3 9 13 13 2 9 13 3 2
27 16 15 9 13 9 2 13 0 9 7 15 13 2 13 3 3 15 9 1 7 3 9 2 9 13 2 2
12 13 9 7 13 9 13 0 11 11 9 1 2
5 11 2 9 7 9
20 15 9 4 13 9 3 0 9 9 16 15 9 2 7 9 13 3 3 9 2
21 13 3 11 2 3 13 11 11 2 15 13 0 9 9 2 8 8 8 8 2 2
29 11 13 3 0 1 9 2 16 15 13 0 2 0 7 3 13 9 2 15 4 13 3 15 0 9 9 9 1 2
13 11 13 0 9 2 7 9 4 13 3 15 0 2
8 3 11 13 3 12 0 9 2
15 9 4 13 3 15 13 2 16 11 4 13 0 9 9 2
17 13 3 0 9 3 15 9 3 13 11 11 2 9 9 7 9 2
6 15 13 9 12 9 2
38 9 13 11 11 2 13 11 9 2 2 15 4 15 3 13 3 3 0 9 2 13 9 2 7 9 13 3 7 3 3 13 15 9 2 7 0 9 2
13 13 0 9 2 2 11 11 2 11 11 11 2 9
17 11 11 13 3 15 0 9 2 3 9 9 13 9 13 3 9 2
19 11 4 13 0 2 9 2 2 8 2 15 15 13 13 3 8 7 9 2
14 7 15 0 2 15 13 13 15 0 9 2 0 3 2
26 16 13 9 11 9 7 9 2 13 13 15 9 11 2 11 11 11 11 11 11 11 2 11 11 11 11
30 9 13 3 3 13 9 7 11 9 2 9 13 11 0 9 2 2 15 1 13 3 13 3 9 7 15 0 13 9 2
15 15 1 0 13 13 3 8 9 7 15 15 9 13 9 2
11 15 13 3 0 9 9 2 3 13 13 2
16 0 15 3 13 16 15 9 0 9 7 3 3 13 15 0 2
5 11 13 0 9 9
11 11 13 3 13 9 11 8 7 8 9 2
4 9 13 0 2
12 0 9 13 13 9 3 16 3 0 12 9 2
20 9 0 9 1 9 0 9 12 7 15 3 13 4 13 15 9 3 12 9 2
15 9 0 9 12 1 13 15 9 13 9 12 9 13 9 2
11 9 13 12 9 9 9 0 12 9 1 2
9 15 13 3 12 9 7 12 9 2
15 9 9 4 3 13 15 0 9 1 9 7 13 11 9 2
19 13 3 13 2 3 15 13 13 12 7 12 9 9 0 0 2 0 9 2
13 3 15 4 13 0 2 2 15 3 3 2 9 2
11 3 3 9 3 3 13 0 13 15 9 2
16 13 2 16 15 9 13 3 3 3 3 16 15 3 4 13 2
17 9 7 9 9 9 13 3 7 15 9 15 13 15 9 3 9 2
12 3 15 13 3 9 3 13 2 7 13 13 2
4 13 3 3 2
5 9 7 9 9 9
14 16 15 11 3 13 2 13 15 9 3 3 3 3 2
15 13 3 3 9 1 15 9 7 13 3 3 2 15 13 2
15 0 9 13 9 9 2 7 16 9 13 2 13 3 3 5
8 9 9 13 3 12 9 9 2
18 15 9 9 13 13 15 0 9 2 7 0 7 0 2 2 9 9 2
13 8 13 9 15 0 9 9 2 15 13 0 9 2
17 7 3 0 9 13 2 3 0 9 15 9 13 2 15 15 13 2
8 9 9 13 3 9 13 9 2
14 16 11 13 0 9 2 15 13 13 9 15 9 11 2
12 11 13 3 13 15 9 9 2 11 3 13 2
11 15 13 3 9 2 15 1 4 13 11 2
15 11 13 11 2 13 0 13 9 9 7 13 0 9 8 2
6 9 13 3 7 3 2
11 11 1 15 13 13 2 11 1 13 3 2
21 11 13 13 9 9 12 9 2 3 15 9 9 13 12 12 9 9 13 13 13 2
10 9 2 9 2 9 2 9 2 9 2
4 0 9 9 2
16 15 9 9 13 9 9 2 15 13 11 9 2 15 11 9 2
20 15 11 2 11 9 13 9 2 16 9 9 13 9 7 15 13 9 3 3 2
9 9 9 13 9 9 13 4 13 2
17 9 13 9 13 3 9 2 16 11 8 13 15 9 13 15 1 2
10 3 13 15 2 7 13 3 16 13 2
11 3 2 9 4 3 15 13 2 13 13 2
8 15 15 4 15 13 15 13 5
4 0 9 7 9
18 3 15 13 15 1 13 0 9 2 3 13 3 16 3 9 15 13 2
1 9
15 9 4 13 3 3 2 7 3 2 2 9 13 15 13 2
24 11 8 8 8 2 0 8 13 13 9 7 15 13 11 11 11 2 3 15 8 4 3 13 2
19 11 13 12 9 12 9 2 1 9 2 7 15 13 3 3 12 9 1 2
5 6 3 13 9 2
10 9 1 13 3 0 9 16 3 13 5
16 2 3 3 9 13 15 1 16 9 13 9 7 3 13 8 2
3 9 9 9
11 13 15 3 3 12 3 0 9 9 9 2
7 13 3 13 9 9 9 2
13 9 9 13 3 9 2 15 15 13 7 13 11 2
19 9 4 13 13 9 11 11 9 2 15 9 13 15 16 9 7 11 12 2
7 3 9 13 3 4 13 2
19 9 4 13 12 9 2 15 13 0 9 2 3 2 7 2 3 2 9 2
9 9 13 3 3 3 7 9 9 2
5 9 13 0 9 2
6 6 2 13 11 13 2
9 9 9 13 0 9 2 11 9 2
11 9 13 12 9 1 9 9 3 15 13 2
27 9 13 0 2 7 15 4 13 3 15 9 2 16 11 2 11 9 13 12 9 7 9 9 9 9 12 2
9 9 4 13 9 9 9 7 9 2
25 13 9 7 15 9 2 7 16 13 13 15 9 7 15 9 9 2 13 15 3 0 13 9 13 2
22 3 13 9 12 9 2 15 13 15 13 2 15 4 3 13 3 15 3 2 16 13 2
19 9 4 3 13 11 11 9 11 12 2 7 9 13 15 3 15 9 9 2
16 13 13 3 15 9 9 9 9 2 7 13 9 12 0 9 2
13 0 9 2 15 9 9 9 2 4 13 9 9 2
21 9 13 13 15 9 7 16 15 13 13 2 4 15 13 3 3 0 9 2 9 2
25 15 2 15 9 4 13 2 13 15 3 13 9 13 7 15 15 13 7 13 13 15 3 15 13 2
14 13 3 4 9 2 16 4 13 2 13 13 13 9 2
7 3 15 13 3 15 9 5
4 15 9 2 2
14 6 2 4 4 13 3 0 9 0 9 11 2 2 2
3 6 13 2
5 11 13 0 9 2
19 3 13 15 0 9 9 9 11 2 3 0 9 16 4 3 13 13 9 2
10 9 0 9 13 9 1 13 3 11 5
23 8 8 8 2 16 13 3 13 15 12 9 9 3 15 4 3 13 9 7 13 3 9 2
9 8 8 2 9 13 15 3 9 2
7 9 13 11 7 13 9 5
7 13 6 0 9 13 0 2
22 9 13 9 2 16 13 9 9 9 1 2 16 15 13 3 13 3 0 13 9 9 2
7 7 13 3 13 9 9 2
6 7 13 9 9 13 2
29 13 15 13 9 3 0 2 0 7 3 3 9 13 0 16 13 0 9 15 2 16 15 3 13 7 3 13 15 2
12 13 3 4 3 13 2 7 15 13 3 9 2
5 6 13 3 3 5
9 3 9 9 13 3 3 0 9 5
14 9 9 13 15 15 9 9 0 11 2 9 2 9 2
6 7 11 13 12 9 2
24 11 7 11 1 13 9 7 9 9 2 13 0 7 0 9 2 9 2 7 11 9 13 9 2
11 13 3 0 9 7 13 3 0 13 15 2
8 9 2 7 15 13 3 9 5
8 0 9 13 3 13 9 9 2
13 13 3 13 3 7 15 3 13 3 0 7 0 2
13 13 3 9 9 7 3 13 11 11 13 9 9 2
15 13 3 3 3 0 9 2 16 13 9 13 9 13 0 2
12 16 0 9 4 13 12 9 2 13 9 9 2
7 3 4 3 13 9 9 2
15 9 0 9 13 13 13 9 2 15 3 0 9 1 13 2
28 0 0 9 9 13 0 2 3 13 2 13 13 11 9 7 13 9 13 9 2 16 9 1 13 13 15 9 2
6 13 3 11 1 11 2
24 3 0 9 2 9 3 13 7 13 2 15 13 3 0 7 3 3 2 13 0 7 13 3 2
5 3 0 2 2 5
13 13 3 3 0 2 16 13 3 13 11 15 9 2
18 9 13 3 0 9 11 7 11 9 2 7 3 13 12 9 9 3 2
15 0 0 13 13 9 9 9 9 2 15 13 3 9 9 5
28 3 3 13 9 13 3 0 9 7 15 13 0 9 13 2 16 15 9 13 9 15 9 16 9 9 13 11 2
6 0 9 13 3 3 2
30 11 13 15 9 2 13 13 3 15 9 2 13 15 9 13 7 3 15 11 11 0 9 13 13 2 9 13 0 9 2
23 9 13 3 9 13 7 13 13 7 3 13 15 2 16 3 13 3 13 0 9 2 6 5
19 11 9 13 3 0 2 7 3 3 13 0 9 7 0 9 2 15 13 2
12 13 2 16 9 13 3 13 2 15 9 13 2
14 15 4 4 13 9 13 15 0 9 7 9 2 2 5
14 6 3 3 13 15 9 2 7 9 13 3 3 9 2
14 15 9 4 13 3 13 2 15 15 13 16 13 3 2
5 8 8 8 8 2
3 9 9 2
11 2 9 4 13 3 0 0 3 3 9 5
8 2 13 3 9 3 7 0 9
13 2 9 9 13 1 9 3 0 7 3 3 0 2
12 2 15 2 11 9 7 11 13 2 2 2 2
4 6 3 0 5
14 2 2 7 3 15 13 4 3 13 13 15 11 9 2
13 2 13 3 3 0 13 13 0 0 9 7 0 2
9 2 13 9 0 9 2 9 5 2
11 2 9 5 11 5 11 13 3 3 0 2
3 7 9 2
7 2 9 13 3 0 9 2
13 3 3 2 16 9 13 15 0 0 9 0 15 2
8 3 0 2 15 13 13 13 2
7 13 3 2 13 0 6 2
18 2 16 9 9 13 9 13 3 3 3 9 13 13 13 7 3 2 5
3 0 11 2
6 2 13 0 13 3 5
6 3 9 13 3 9 2
9 7 13 3 3 11 12 9 1 2
7 13 3 15 15 9 2 5
1 11
6 3 9 3 3 9 5
17 13 0 9 11 7 11 1 0 2 9 2 9 3 11 11 1 2
18 13 4 3 3 13 11 7 11 2 7 9 9 9 1 13 3 0 2
8 13 3 13 15 9 7 9 2
13 6 2 13 4 4 13 0 9 7 9 15 9 2
38 11 13 3 0 9 15 13 0 0 12 9 0 2 7 9 13 3 9 7 11 11 2 15 13 11 7 15 9 0 9 9 7 9 7 9 1 9 2
15 9 13 0 7 3 9 7 11 9 2 11 13 2 2 2
16 13 3 0 13 2 3 13 3 9 13 9 7 9 3 3 2
10 7 9 2 3 3 9 2 3 13 2
12 11 13 3 0 0 9 13 9 3 0 9 2
6 9 2 9 2 9 2
24 13 3 0 13 2 3 0 9 9 2 15 4 13 15 12 9 7 12 9 2 4 3 13 2
21 12 9 1 13 15 9 11 7 11 9 9 9 2 3 13 13 3 0 8 8 2
14 3 15 9 13 13 15 7 3 13 13 3 3 3 2
12 7 3 3 16 11 9 2 13 3 13 9 5
22 9 13 13 0 9 7 9 7 13 15 9 9 2 13 3 3 0 9 15 9 9 2
20 13 9 3 11 9 13 9 7 9 2 7 13 3 3 0 9 3 0 9 2
16 3 0 13 3 15 2 16 9 1 13 11 13 11 7 11 2
24 11 13 9 2 3 12 9 9 2 7 13 0 13 15 9 9 11 2 9 2 11 9 3 2
7 9 1 13 0 0 9 2
15 3 15 9 13 0 2 16 13 4 12 9 13 3 9 5
16 7 0 9 9 13 15 9 3 3 0 2 9 7 3 9 2
9 6 2 13 13 9 15 11 9 2
8 13 3 0 9 2 0 9 2
16 13 9 9 2 16 15 13 3 3 9 2 15 13 0 9 2
10 13 3 9 13 13 2 15 3 13 2
12 3 15 13 3 0 3 3 11 7 11 9 5
15 13 3 9 13 7 13 9 7 9 2 7 9 3 9 2
13 9 4 3 13 3 2 13 4 13 15 0 9 2
17 3 13 12 3 0 9 2 13 3 3 2 16 4 13 0 9 2
2 0 2
19 13 3 3 0 9 15 2 3 13 2 7 9 13 13 3 0 9 0 2
19 13 15 9 11 9 2 9 7 9 2 9 2 3 13 3 3 15 9 2
21 3 15 13 15 2 13 4 13 15 9 0 9 9 0 9 2 7 13 3 9 2
7 11 7 11 9 13 0 2
7 15 9 9 13 3 9 2
4 3 9 11 2
14 11 9 13 0 2 16 13 3 9 7 15 1 9 2
17 13 9 2 15 13 15 15 9 2 7 3 13 3 15 1 3 2
13 9 13 3 0 2 0 12 9 0 9 3 9 2
20 3 13 3 13 3 9 2 7 9 2 1 2 7 13 15 0 9 3 3 5
22 9 13 9 7 13 3 12 9 3 0 9 2 9 9 1 9 9 13 9 2 6 2
13 15 13 15 9 2 16 11 3 13 3 3 3 2
1 0
6 0 9 13 3 9 2
20 3 3 13 13 9 3 2 3 3 13 3 0 13 15 2 16 13 3 9 2
21 4 3 4 13 2 16 3 13 15 0 9 13 3 3 2 7 9 3 15 1 2
9 7 9 9 9 2 7 13 9 5
25 16 13 2 16 15 9 3 13 3 2 6 2 7 13 2 3 13 2 16 4 3 3 13 9 5
12 0 8 9 4 13 3 15 9 9 9 1 2
10 15 13 3 9 2 13 0 15 9 2
10 0 2 0 0 9 13 3 15 9 2
15 0 0 9 13 3 0 2 0 2 9 2 13 3 0 2
5 9 3 12 9 2
4 9 8 8 2
5 6 13 15 11 2
14 7 0 2 0 9 13 13 2 3 15 15 13 9 2
26 11 13 0 2 16 15 9 1 9 9 13 15 2 16 13 0 9 7 13 0 9 2 16 9 13 2
8 7 15 4 13 3 15 9 2
32 11 9 4 13 2 16 15 3 9 7 9 13 11 13 3 3 0 0 2 13 3 13 15 9 2 13 15 13 3 3 3 2
30 15 13 3 3 3 9 1 2 13 16 15 0 9 13 9 16 13 2 3 2 9 7 15 13 13 13 15 9 2 2
3 6 3 5
14 15 9 9 0 9 9 2 4 13 3 0 2 3 2
19 13 0 8 8 15 15 9 2 9 2 2 0 7 0 2 7 3 0 5
11 6 6 2 7 3 0 9 13 9 9 2
5 13 9 15 0 2
2 11 12
6 3 4 15 9 13 2
16 12 9 9 13 3 3 2 0 9 9 1 7 3 9 13 2
32 3 3 9 0 11 11 13 0 2 3 9 2 9 13 3 9 7 13 2 7 15 9 9 13 3 3 3 0 9 13 9 2
25 9 11 11 13 0 9 2 15 1 15 9 2 15 9 13 3 3 15 9 2 13 7 9 13 2
23 9 9 11 2 9 7 3 15 1 2 16 9 13 13 15 3 2 16 9 13 3 3 2
20 9 9 13 3 9 13 9 2 7 9 4 13 9 9 2 15 13 3 3 2
19 13 3 0 7 0 9 2 3 9 13 3 3 9 15 3 13 7 13 5
11 9 3 13 13 2 16 4 13 15 0 5
18 9 13 0 9 11 9 2 15 13 0 11 11 9 9 7 3 13 2
10 13 1 9 9 2 15 13 3 9 2
11 9 13 3 13 9 7 13 0 9 9 2
8 13 3 0 11 7 15 9 5
12 15 11 13 12 9 11 11 9 11 8 9 2
18 11 13 3 3 15 9 16 15 2 0 9 2 15 13 9 2 9 2
13 9 13 3 16 15 2 3 16 3 13 0 9 5
20 0 9 13 9 13 0 9 9 0 9 2 7 13 13 9 13 7 13 15 2
16 0 9 13 15 3 2 16 12 9 9 7 9 13 13 3 2
14 11 7 11 13 13 15 7 11 0 9 7 15 9 2
4 8 8 8 2
9 13 11 1 3 0 9 9 1 2
11 15 9 15 2 16 9 2 6 2 13 2
15 9 9 13 3 13 9 9 15 9 2 15 13 9 13 2
1 8
9 6 2 3 13 13 9 3 0 2
14 3 3 13 11 2 13 4 13 3 12 9 15 9 2
14 9 2 12 9 13 15 9 2 7 3 13 13 3 2
9 13 3 9 13 9 7 13 9 5
12 3 0 13 15 2 16 13 7 13 0 9 2
10 13 13 9 2 7 3 5 6 6 2
3 13 9 2
11 13 15 2 16 13 0 9 4 3 13 2
9 7 15 9 9 13 15 9 3 2
7 0 9 2 15 13 0 9
46 3 13 3 3 0 9 1 2 2 0 9 11 2 0 9 2 13 2 2 0 11 9 2 9 2 2 0 9 2 9 11 2 0 2 0 9 2 8 2 8 2 8 2 2 13 2
17 0 9 13 3 3 2 3 3 15 15 9 9 13 9 2 0 2
13 3 13 9 9 2 13 9 9 3 13 9 1 2
16 13 3 3 15 9 2 16 3 15 11 13 3 0 16 11 2
5 6 2 15 9 2
4 7 15 9 2
19 3 15 7 9 13 15 9 2 16 15 13 0 2 13 5 0 2 9 2
6 3 4 13 13 9 2
7 0 9 7 9 15 9 2
5 9 2 9 7 9
4 3 13 13 2
6 11 9 4 13 9 2
16 15 9 13 12 9 9 2 3 3 0 13 13 2 7 0 2
13 9 13 9 9 13 3 2 16 4 3 13 9 2
19 15 4 3 3 13 9 1 9 2 7 15 13 13 15 13 0 0 9 2
15 9 13 9 2 9 2 9 2 9 2 9 7 3 9 2
6 9 9 15 0 9 2
6 2 7 9 13 0 2
9 13 9 9 9 7 13 9 15 2
2 0 13
3 9 1 9
11 3 3 15 13 0 9 11 13 9 9 2
8 3 13 15 0 9 2 0 2
14 0 13 2 9 13 13 3 3 3 0 3 13 2 2
9 9 13 9 2 13 0 0 13 2
1 6
4 13 9 7 9
24 9 13 9 9 2 9 2 0 13 2 9 9 7 9 2 13 13 3 9 13 9 2 2 2
10 13 0 2 7 13 0 7 0 0 2
6 9 13 3 3 9 9
21 9 13 9 9 9 1 7 3 13 9 2 15 15 13 13 2 7 13 15 9 2
1 9
7 3 0 9 2 9 0 2
6 9 13 12 9 9 2
6 9 9 13 3 11 2
13 9 13 9 7 0 9 7 15 9 9 7 9 2
14 9 13 12 0 9 13 7 13 15 3 9 13 0 2
4 9 13 9 1
11 9 9 2 13 2 9 13 1 13 9 2
20 9 13 9 2 9 2 9 2 13 9 2 9 2 13 9 2 9 2 9 2
22 13 9 9 2 13 9 7 13 2 13 13 9 7 15 9 7 13 9 3 3 13 2
11 13 3 3 9 7 9 9 7 13 9 2
7 13 3 2 13 9 13 2
2 13 2
10 15 9 4 13 3 0 0 1 9 2
17 9 13 3 0 9 7 15 13 3 3 9 2 3 9 13 0 2
4 9 7 0 9
6 15 3 3 13 3 0
36 9 0 9 2 9 2 9 9 2 0 9 2 15 9 13 9 0 9 2 2 13 9 3 2 0 9 2 13 9 2 2 9 7 3 9 2
9 13 13 0 7 6 9 16 13 0
17 0 13 3 15 15 0 9 15 13 13 9 9 9 9 1 11 2
18 15 9 13 9 2 9 2 0 9 2 0 9 2 9 7 0 9 2
6 9 13 15 0 9 2
3 0 0 9
10 9 13 3 3 13 9 2 3 3 2
19 7 15 9 3 13 3 0 9 9 2 3 13 3 3 9 13 0 9 2
10 9 13 9 2 9 7 13 9 1 2
9 15 13 3 12 0 9 3 2 2
18 13 9 0 9 1 9 2 16 13 9 13 7 13 0 2 9 2 2
37 13 9 9 9 9 2 12 9 13 3 7 3 13 3 0 9 2 5 13 9 7 9 9 7 13 15 9 13 9 7 13 15 3 9 13 2 2
15 3 9 13 12 9 9 2 9 2 9 9 7 9 9 2
30 13 9 9 9 1 0 9 2 3 3 13 9 9 13 9 2 16 15 13 13 3 0 2 16 9 4 13 15 3 2
22 9 13 13 9 7 13 16 3 4 13 9 9 3 3 9 2 7 3 15 9 13 2
9 3 3 9 9 1 7 0 13 2
12 9 7 9 1 13 3 3 9 13 0 9 2
15 9 13 15 9 3 9 13 2 16 13 15 3 3 13 2
2 0 9
9 3 0 7 0 9 15 9 13 2
2 9 9
8 0 9 13 3 9 1 2 2
10 3 0 9 9 2 13 0 9 2 2
1 9
19 12 0 9 13 15 9 2 9 13 13 3 12 9 3 16 4 13 9 2
13 13 9 3 3 9 3 7 3 12 0 0 9 2
12 13 9 3 9 3 5 3 9 13 3 0 2
14 9 13 3 12 9 13 9 2 3 9 7 9 13 2
8 9 13 15 9 3 12 9 2
9 9 13 12 9 9 13 9 9 2
12 3 12 9 9 7 7 3 13 9 12 9 2
45 12 9 13 9 9 9 2 0 9 12 0 9 9 13 5 3 9 2 0 13 12 9 13 5 12 9 8 8 7 0 13 9 1 12 9 9 0 9 0 9 5 9 12 9 2
20 3 9 13 13 9 2 7 15 9 13 3 3 0 2 16 13 15 3 9 2
12 9 13 13 7 13 9 7 15 9 3 13 2
12 15 13 13 15 9 2 16 15 13 3 9 2
11 13 9 13 0 9 1 9 1 9 13 2
17 9 13 12 9 0 9 5 12 9 0 9 5 12 9 8 8 2
16 9 9 7 3 12 9 9 9 2 13 9 2 9 7 9 2
1 9
22 15 9 13 11 9 3 9 9 2 2 7 15 9 1 13 9 7 0 9 9 9 2
17 15 9 7 9 13 9 13 4 3 13 2 3 3 3 13 2 2
10 15 1 13 15 9 3 7 9 13 2
15 9 13 13 3 9 2 3 0 13 4 13 3 9 9 2
80 9 15 13 13 15 9 2 11 9 9 2 7 9 2 11 9 12 0 2 9 7 13 15 9 0 9 7 13 15 3 15 9 3 9 7 9 2 9 2 0 9 2 7 9 7 9 2 2 9 2 9 7 9 2 9 2 13 9 7 3 9 7 9 13 0 13 3 9 12 9 7 9 3 0 0 9 0 9 1 2
6 13 13 0 9 2 2
6 9 4 13 0 9 1
5 9 2 9 9 2
5 3 13 0 9 2
9 2 7 3 15 15 9 13 2 2
2 9 9
15 13 9 9 2 13 13 0 9 2 7 13 15 13 9 2
11 13 9 7 9 9 1 7 13 9 9 2
10 13 9 12 2 12 9 3 12 9 2
3 13 3 2
12 9 3 13 0 9 7 9 3 3 0 9 2
1 9
13 0 9 2 9 9 13 13 3 3 2 15 12 2
4 9 13 3 2
8 13 9 7 0 9 3 9 2
9 13 9 9 3 2 0 9 13 2
12 13 0 9 3 7 13 15 9 9 3 13 2
6 13 3 9 13 9 2
6 13 9 9 9 1 2
7 13 12 9 3 12 9 2
12 13 13 3 3 2 16 9 13 13 3 2 2
13 7 16 13 0 9 2 16 15 2 13 3 3 3
2 0 9
8 0 9 13 0 9 13 9 2
4 9 2 9 2
2 9 2
22 12 9 0 9 5 12 9 9 5 12 9 9 5 12 9 9 5 3 12 9 0 9
14 5 13 9 9 2 13 9 2 9 7 13 0 9 2
22 13 9 7 0 9 9 2 9 1 2 1 9 2 13 9 9 3 9 1 9 9 2
2 9 2
19 12 9 13 9 5 12 9 9 5 9 2 9 2 9 2 13 9 7 9
2 9 2
56 12 9 9 9 2 9 2 9 2 9 2 9 2 13 9 2 9 12 9 2 12 0 9 0 9 2 12 0 0 9 2 12 9 9 13 2 9 12 9 0 9 2 9 12 0 9 3 13 2 0 9 13 2 9 7 9
20 5 13 9 0 7 13 9 0 2 13 9 3 9 7 13 9 3 13 9 2
4 13 9 3 2
16 13 9 3 9 2 3 9 2 15 9 7 3 0 3 9 2
9 13 9 3 12 0 9 12 9 2
14 15 9 13 15 3 0 7 9 13 3 7 13 0 0
7 15 9 13 9 9 3 3
3 9 0 9
11 9 13 0 9 13 3 3 3 13 2 2
13 13 15 15 9 0 9 9 7 13 15 0 9 2
5 13 9 9 9 2
15 9 13 13 3 0 0 2 16 9 13 13 13 9 9 2
9 13 9 13 3 1 0 9 9 2
7 13 3 0 3 9 1 2
7 9 13 0 12 9 9 2
2 6 2
3 9 13 9
16 0 9 2 9 13 15 3 3 3 9 2 16 9 13 3 0
12 13 9 9 7 3 15 15 9 1 0 9 2
10 13 9 0 9 9 7 9 13 9 2
11 13 9 9 2 0 9 7 13 15 9 2
9 9 7 9 9 1 2 13 13 2
14 13 12 0 9 0 7 3 3 0 3 12 9 2 2
17 15 13 15 9 12 0 9 7 3 13 12 0 9 12 9 9 2
5 2 9 9 9 2
4 9 0 9 2
6 9 9 13 0 9 2
19 3 3 4 13 2 16 13 3 0 9 2 2 16 3 2 9 2 13 2
28 0 9 2 13 0 7 13 3 13 3 0 2 9 3 9 2 13 9 2 9 3 2 15 0 5 9 3 2
18 15 12 9 2 13 2 13 9 13 13 9 1 11 9 11 11 9 2
2 0 9
11 15 13 0 2 13 3 3 0 3 13 2
7 9 13 3 9 7 9 2
6 0 9 13 9 9 2
10 15 13 9 9 9 1 13 9 9 2
11 13 9 1 3 15 15 9 7 0 9 2
3 13 9 2
5 9 13 12 9 2
5 9 0 12 9 2
2 9 2
22 16 9 1 13 9 7 9 13 3 0 7 16 13 9 2 13 3 13 9 3 2 2
4 13 3 1 9
10 0 9 4 13 15 9 16 9 2 2
8 9 13 0 9 15 9 1 2
2 0 9
5 0 9 13 2 2
13 9 13 3 13 2 2 7 0 9 15 3 9 13
7 13 9 5 9 0 9 2
11 13 9 2 13 9 7 9 7 13 13 2
11 13 9 7 9 7 13 15 9 1 13 2
9 13 9 0 7 13 9 3 13 2
6 13 9 9 7 9 2
11 9 13 12 9 9 3 3 3 0 9 2
5 7 13 0 9 2
2 15 3
6 15 0 9 13 2 2
19 3 12 9 4 15 15 9 13 2 13 3 3 4 15 9 0 13 2 2
13 9 0 9 13 9 9 2 16 4 0 9 13 9
14 15 9 13 13 15 2 16 15 9 1 13 9 2 2
18 2 7 9 9 9 13 9 13 9 2 13 9 4 3 3 13 2 2
11 13 15 9 13 2 16 15 13 9 2 2
2 15 9
20 9 9 15 9 13 0 0 7 15 15 9 3 9 13 9 13 3 9 9 2
12 16 9 13 0 9 1 3 13 15 9 9 2
16 15 2 15 9 13 3 13 9 9 9 9 13 0 12 9 2
2 9 2
9 3 3 13 15 15 9 15 0 2
4 15 13 13 2
14 3 15 3 0 9 13 2 16 15 9 3 13 9 2
7 13 3 13 15 3 3 2
25 0 7 0 9 2 15 13 9 3 13 9 2 1 12 5 15 9 13 9 13 13 15 9 9 2
12 13 9 13 15 15 9 2 7 0 9 9 2
24 16 0 9 4 13 15 3 2 13 9 1 15 2 13 9 15 9 2 9 2 9 7 9 2
8 13 9 2 15 15 15 13 2
19 13 9 3 15 9 9 2 16 9 0 9 13 9 15 15 9 9 9 2
11 9 2 13 2 16 13 9 2 13 3 2
4 3 7 15 2
28 3 3 9 2 3 15 4 13 15 3 9 2 2 15 13 3 9 9 13 9 2 13 9 2 9 2 9 2
44 3 2 9 13 2 16 9 13 13 9 9 2 2 13 9 9 13 9 13 13 9 3 2 15 13 3 3 15 1 9 2 2 15 13 9 9 13 2 3 15 13 9 2 2
19 13 9 3 3 0 15 2 7 13 15 3 13 13 9 1 0 9 9 2
15 15 16 9 13 9 9 3 2 16 13 13 3 0 9 2
19 0 13 2 16 15 13 13 9 13 9 1 15 2 15 9 15 3 13 2
16 0 9 13 15 9 7 13 15 3 16 2 13 0 9 2 2
12 6 13 3 2 9 2 7 15 13 13 9 2
21 3 9 13 3 13 15 9 9 2 15 9 13 13 3 1 0 7 3 13 9 2
9 15 9 4 13 0 9 3 9 2
17 15 9 0 9 2 13 0 9 2 16 0 9 13 3 9 9 2
10 13 9 13 11 9 2 9 13 9 2
34 13 0 9 7 13 3 13 15 9 9 2 15 9 13 0 2 9 3 7 3 0 13 15 13 9 2 9 2 15 13 0 0 9 2
15 13 3 12 13 9 13 9 2 16 9 13 3 0 9 2
15 13 2 13 9 3 13 3 2 3 16 13 13 9 9 2
29 13 9 7 13 15 0 2 3 9 2 3 9 2 13 3 2 3 13 3 13 9 9 16 9 4 13 15 0 2
8 2 6 15 9 2 2 13 2
5 2 0 9 2 2
13 13 13 7 13 9 2 3 9 13 9 3 3 2
12 2 12 9 13 13 13 12 9 2 2 13 2
15 0 9 9 13 3 0 9 2 11 2 15 9 2 1 2
3 13 9 2
7 11 2 13 3 13 13 2
12 9 2 15 3 13 13 2 3 16 15 13 2
8 7 13 15 13 15 9 13 2
8 0 9 13 9 13 9 9 2
6 13 0 7 0 9 2
5 9 13 0 9 2
3 2 6 2
33 3 0 0 9 2 15 4 3 13 13 15 9 2 3 13 15 15 9 9 9 3 16 0 9 13 9 4 13 15 15 0 9 2
24 3 15 4 13 13 11 9 2 13 1 16 13 4 13 0 3 7 3 15 13 9 9 3 2
17 9 3 13 9 9 13 9 1 7 13 2 16 13 3 3 0 2
12 7 13 15 13 3 15 9 13 9 13 9 2
2 3 2
19 15 13 13 13 7 13 9 3 9 13 2 3 0 9 13 3 3 2 2
18 7 9 8 2 9 13 7 9 0 15 9 2 7 9 0 15 9 2
12 9 13 13 9 9 2 15 13 13 0 9 2
15 16 9 13 9 9 2 9 7 9 2 13 9 0 9 2
13 7 3 0 9 2 3 15 15 9 3 3 13 2
7 16 9 13 13 13 9 2
6 9 7 9 15 13 2
22 7 16 9 13 9 15 9 13 9 9 9 7 13 9 13 9 9 2 13 9 9 2
20 13 9 13 9 13 0 9 2 13 15 9 1 3 9 1 2 9 3 13 2
12 9 2 16 15 13 15 2 3 13 3 9 2
12 9 2 13 2 16 3 15 13 12 0 9 2
7 9 2 13 3 3 9 2
11 9 2 6 3 15 3 9 3 3 13 2
8 9 2 6 2 13 3 3 2
5 9 2 3 3 2
7 9 7 9 2 12 9 2
15 16 13 13 9 2 13 15 3 12 9 9 2 12 9 2
12 13 13 9 3 2 7 7 13 15 9 9 2
36 16 9 13 2 13 9 2 3 9 2 15 13 3 9 7 13 0 9 2 2 9 2 9 2 9 7 13 9 0 9 2 13 9 13 9 2
14 13 12 9 9 3 12 9 2 13 3 4 9 13 2
20 16 9 13 9 2 13 9 13 3 12 9 9 9 2 12 9 2 1 9 2
27 15 1 13 9 7 13 9 9 0 9 7 13 9 12 9 9 2 13 13 7 13 9 3 3 13 9 2
9 13 3 15 9 7 13 3 9 2
4 13 3 3 2
5 13 13 9 1 2
9 15 0 9 13 9 9 13 9 2
5 13 0 2 13 0
5 13 0 9 9 2
8 16 15 13 0 2 13 0 2
8 16 15 13 9 2 13 9 2
16 13 15 0 9 2 16 15 15 13 2 16 13 13 9 2 2
24 7 15 13 15 15 9 2 16 3 2 7 3 3 3 2 4 13 9 2 13 13 15 13 2
9 3 3 13 2 16 3 3 3 2
11 4 3 3 13 2 16 3 0 9 13 2
5 3 9 13 0 2
12 15 3 13 15 0 9 7 13 3 0 9 2
11 15 13 0 13 2 13 2 13 7 13 2
15 2 6 2 15 9 2 6 2 13 15 3 2 0 9 2
13 9 13 2 6 2 3 3 7 3 13 9 9 2
11 9 2 6 2 9 13 7 9 15 13 2
3 6 2 2
22 7 9 13 9 2 16 15 13 3 2 3 3 3 2 16 13 15 9 13 0 9 2
12 7 9 13 13 13 2 16 15 13 3 9 2
5 3 16 9 13 2
19 0 13 9 2 16 9 4 13 9 9 13 9 2 16 15 13 13 9 2
3 15 13 2
10 7 3 6 13 2 13 15 3 0 2
13 13 15 9 1 9 2 4 15 3 13 15 0 2
7 9 13 2 16 3 3 2
3 13 9 2
16 0 9 1 15 13 2 16 2 13 0 16 13 0 9 2 2
24 9 13 9 13 3 13 7 3 9 13 9 0 9 2 16 13 3 0 9 9 7 3 9 2
14 9 13 3 13 15 9 15 1 2 13 15 15 0 2
12 9 2 3 15 13 2 13 13 0 1 0 2
16 3 9 13 2 16 9 13 3 3 0 2 16 15 13 9 2
11 15 13 2 15 9 13 7 15 9 13 2
16 15 13 0 9 2 15 13 2 13 3 13 0 9 9 13 2
6 3 13 13 9 9 2
6 15 9 13 4 13 2
6 13 3 13 15 9 2
16 15 13 2 16 9 13 3 0 9 7 13 3 9 1 9 2
8 9 2 15 13 3 11 9 2
4 9 2 3 2
6 9 2 9 2 3 2
4 9 2 3 2
8 9 2 6 2 9 13 9 2
6 9 2 2 0 9 2
27 4 3 13 3 9 2 0 9 9 2 7 3 9 2 15 13 0 2 7 3 3 3 3 13 2 9 2
9 3 3 15 13 13 0 9 13 2
8 15 9 13 3 12 5 9 2
19 9 13 3 13 0 13 2 16 13 4 13 12 9 9 7 9 3 3 2
27 9 4 13 0 9 3 3 9 9 2 7 9 4 13 3 12 9 9 2 16 15 13 3 16 12 9 2
11 15 13 0 2 15 13 3 12 9 9 2
7 7 9 2 15 13 0 2
4 15 13 13 2
17 15 13 2 16 9 9 1 13 0 7 16 9 13 15 16 9 2
11 7 15 2 15 13 0 3 0 11 3 2
26 3 13 3 0 9 2 7 3 0 9 13 15 2 16 13 13 9 15 9 2 15 13 15 9 9 2
20 13 3 3 11 2 15 9 13 13 3 9 7 15 9 9 0 13 0 0 2
7 3 15 13 13 0 9 2
20 13 13 9 13 9 2 13 9 13 9 7 13 9 2 15 3 3 13 9 2
6 13 15 15 9 13 2
19 15 2 16 15 9 13 13 9 0 2 13 13 2 16 15 13 15 9 2
17 15 9 13 13 9 15 9 2 16 15 13 9 7 13 0 15 2
7 13 0 9 2 12 9 2
8 3 2 9 1 9 7 13 9
14 3 13 9 9 9 13 9 2 13 9 1 12 9 2
6 3 4 13 3 9 2
8 13 9 3 16 13 9 9 2
11 6 2 13 13 9 3 3 9 1 9 2
18 16 13 3 13 2 3 13 9 2 15 9 13 2 13 3 15 9 2
6 13 9 12 9 9 2
9 13 9 2 9 2 9 7 9 2
14 13 9 2 13 9 7 9 7 13 9 2 13 9 2
15 13 9 15 9 7 13 3 15 9 1 2 13 9 1 2
18 13 9 2 9 2 13 15 1 9 9 2 2 13 9 7 9 9 2
4 13 9 1 2
2 9 9
6 15 13 0 9 9 2
17 7 15 13 13 0 7 0 2 9 2 9 7 9 13 15 13 2
15 7 3 9 9 2 9 2 9 7 9 2 15 15 13 2
12 9 13 11 13 9 13 0 9 7 15 9 2
13 9 13 0 7 13 9 0 9 9 1 13 9 2
19 9 13 9 13 13 16 13 9 12 9 0 9 2 9 7 0 0 9 2
14 13 9 3 0 9 2 15 0 9 13 3 9 1 2
14 9 3 13 2 16 9 13 9 2 7 15 13 3 2
8 3 9 9 13 3 9 13 2
6 9 2 15 15 13 2
4 9 2 15 2
4 9 2 6 2
8 6 2 3 0 13 15 9 2
21 9 2 13 15 15 9 13 2 7 15 3 15 9 4 13 3 9 3 12 9 2
12 9 13 9 9 7 13 9 13 11 9 9 2
13 9 2 13 3 15 9 13 16 15 13 15 9 2
4 3 2 6 2
6 13 15 13 2 13 2
4 9 13 0 2
12 15 13 3 0 13 2 3 15 0 9 13 2
7 15 15 13 7 15 13 2
11 13 13 13 15 9 9 7 9 3 3 2
39 9 13 0 9 2 13 13 13 13 2 13 0 9 9 7 9 2 9 7 9 2 13 15 9 16 3 2 4 15 13 9 7 13 2 3 15 13 9 2
10 9 13 13 3 9 7 9 15 9 2
9 9 1 13 9 13 9 3 9 2
16 0 0 9 13 9 9 1 2 7 3 3 3 16 3 13 2
25 9 13 13 15 2 16 9 13 7 9 1 13 13 2 16 0 9 4 2 3 4 2 13 3 2
18 16 16 9 0 9 13 9 9 2 3 3 13 0 0 13 9 0 2
15 9 13 9 3 0 2 16 0 2 15 9 4 13 3 2
8 9 13 13 3 3 9 9 2
13 9 13 3 0 7 9 13 2 3 16 9 3 2
15 0 13 13 15 3 3 3 9 2 15 1 13 4 13 2
5 13 1 0 9 2
5 9 2 12 9 2
8 13 0 9 9 7 13 0 2
19 13 7 13 9 7 9 2 9 4 13 0 2 9 7 9 4 13 2 2
14 13 9 7 9 7 13 9 2 13 9 0 9 2 2
7 13 9 9 7 13 9 2
11 13 9 9 2 13 3 7 13 9 3 2
20 16 9 9 13 3 13 9 2 13 3 9 7 9 2 9 2 9 7 9 2
14 13 13 9 1 12 9 7 3 2 16 9 13 0 2
7 13 9 7 0 9 1 2
1 9
6 9 13 13 9 9 2
28 0 9 2 0 9 2 0 9 7 3 13 9 13 3 0 9 16 0 13 9 2 0 9 7 3 13 9 2
8 3 0 13 9 13 0 9 2
9 7 0 2 15 13 15 0 9 2
5 6 9 2 13 2
9 9 13 3 0 9 0 9 9 2
12 15 13 2 15 15 13 3 2 16 13 9 2
12 0 7 3 0 9 7 0 2 9 13 9 2
30 15 9 13 2 16 15 9 16 9 4 13 2 13 3 13 2 16 2 15 15 15 13 2 16 0 3 13 2 2 2
15 9 13 0 7 13 2 16 2 3 0 9 7 9 2 2
13 3 13 9 7 13 2 16 15 0 9 15 13 2
11 15 9 13 2 16 2 15 13 15 2 2
10 0 9 4 3 13 9 7 9 9 2
8 9 2 9 2 12 2 12 2
13 13 3 3 9 2 15 9 13 15 9 9 13 2
7 15 9 2 16 15 13 2
17 9 9 9 13 0 0 9 9 0 1 9 2 3 3 0 9 2
13 2 13 2 15 15 15 9 0 9 4 13 2 2
33 7 15 9 2 16 9 13 13 9 0 9 7 9 1 9 2 9 7 0 9 2 13 9 9 2 16 15 15 4 13 9 9 2
14 9 13 13 9 2 16 9 13 9 13 9 1 9 2
25 0 9 13 3 3 3 2 16 2 13 9 13 3 0 9 3 2 7 13 13 9 0 9 3 2
18 13 15 3 3 11 0 9 2 3 12 9 1 2 16 9 3 13 2
22 7 15 9 13 3 9 2 9 13 3 7 13 15 3 2 16 13 15 0 7 0 2
18 15 13 3 0 9 13 9 0 9 3 2 13 13 15 9 9 13 2
13 16 9 13 13 15 0 2 3 15 13 0 9 2
4 8 8 8 2
24 13 15 9 15 9 13 2 15 16 15 9 9 2 15 4 9 9 7 9 13 15 9 13 2
13 0 9 16 13 9 11 2 13 9 13 9 9 2
12 4 13 3 0 9 16 13 0 9 13 9 2
10 9 13 13 9 9 16 9 13 3 2
11 13 13 9 9 2 6 3 0 9 2 2
13 9 13 13 9 9 3 16 13 3 0 1 9 2
18 0 2 16 9 13 15 2 0 9 2 15 9 16 9 9 13 15 2
5 13 15 9 9 2
5 9 2 12 9 2
4 13 9 0 2
5 13 9 0 9 2
10 13 9 9 2 13 9 3 7 13 2
9 13 9 7 13 15 2 13 9 2
15 13 9 2 9 7 9 9 2 13 3 0 9 7 9 2
15 13 3 16 9 13 3 0 7 13 15 3 13 9 9 2
13 13 9 9 7 13 15 9 9 2 13 13 2 2
22 16 9 13 0 2 13 9 9 2 13 9 9 7 9 2 13 13 3 15 1 2 2
14 13 9 7 13 9 7 13 3 9 2 13 13 2 2
7 13 0 9 7 9 1 2
9 3 13 0 9 9 13 0 9 2
13 0 9 13 15 9 3 0 2 13 9 13 3 2
13 15 13 3 9 9 9 13 7 13 11 13 9 2
17 9 4 3 13 9 15 15 7 12 9 2 13 9 13 3 9 2
7 0 9 9 13 0 9 2
5 11 9 2 12 2
16 0 9 2 0 7 0 9 13 3 13 9 3 3 15 9 2
22 3 11 9 13 3 9 2 9 2 9 7 9 9 9 9 13 2 3 13 3 11 2
12 9 9 13 13 2 7 15 4 13 3 9 2
9 9 4 13 7 15 4 13 3 2
11 15 4 13 9 9 3 9 13 9 9 2
19 15 4 13 0 3 7 3 2 9 9 13 2 7 9 13 9 7 9 2
8 15 9 9 13 3 3 9 2
21 9 13 9 2 15 13 4 13 9 3 2 15 13 13 9 13 13 9 0 9 2
7 3 13 9 4 13 9 2
9 0 9 4 3 13 0 3 9 2
14 9 3 13 9 3 3 3 3 7 13 15 3 3 2
14 0 9 9 9 13 3 2 9 13 7 9 9 13 2
19 3 9 13 0 9 15 1 2 16 9 9 13 13 9 2 3 13 11 2
14 15 9 4 13 3 2 16 0 9 9 13 0 9 2
17 15 15 13 3 9 3 15 9 2 16 9 13 9 3 13 15 2
15 0 7 0 9 4 3 3 13 3 3 9 7 9 1 2
20 13 2 16 9 9 7 9 11 0 9 13 9 7 13 0 9 0 9 1 2
26 0 9 2 9 13 11 9 9 13 9 2 7 9 9 9 13 9 13 3 0 7 13 9 9 9 2
37 13 2 16 4 9 13 15 0 0 9 13 9 2 15 13 15 13 9 0 9 15 1 2 16 13 9 2 9 7 9 9 9 3 0 9 9 2
19 0 9 2 0 9 9 2 0 9 2 15 9 9 9 4 13 3 3 2
15 9 7 9 13 0 9 15 9 2 15 9 13 0 9 2
23 3 3 3 3 9 4 13 9 2 7 15 4 13 15 1 9 2 16 13 2 15 13 2
15 15 9 9 13 9 13 3 0 9 15 9 9 13 9 2
14 13 3 0 2 16 0 9 2 3 9 2 13 3 2
25 15 13 15 2 16 3 0 9 3 9 13 9 13 4 13 15 15 9 1 2 16 9 13 13 2
30 3 13 15 9 2 16 13 3 0 2 16 4 13 13 9 3 0 9 2 7 0 9 2 15 13 9 3 9 9 2
39 15 13 2 16 16 3 15 9 13 2 16 9 13 11 2 15 13 9 2 9 13 2 9 4 13 2 16 13 4 3 13 15 9 2 3 9 13 0 2
30 3 4 3 13 13 2 3 9 9 13 7 13 9 3 7 13 7 13 9 3 3 16 13 9 2 15 4 13 9 2
36 9 4 13 15 2 12 9 3 1 2 15 15 4 3 9 13 9 13 3 3 2 3 9 15 2 13 0 9 13 3 0 9 9 7 13 2
23 15 13 9 9 15 9 2 16 13 3 0 13 15 3 9 2 15 13 13 9 13 9 2
23 15 13 3 13 2 3 9 13 2 13 15 0 9 7 13 15 3 3 0 9 15 9 2
13 15 1 9 13 13 9 2 15 13 0 9 9 2
11 13 3 13 12 9 9 9 3 9 1 2
11 15 1 9 7 9 13 9 9 11 9 2
7 13 13 9 2 15 13 2
25 13 13 7 9 11 7 9 15 0 7 0 9 2 15 15 13 7 15 7 15 9 1 15 9 2
21 13 9 2 15 1 9 4 13 3 16 0 9 2 15 9 13 3 3 0 9 2
26 9 13 0 3 13 9 0 9 2 16 0 9 13 3 15 9 13 0 9 2 15 15 9 13 9 2
14 9 13 3 13 0 9 2 7 9 13 0 9 9 2
10 13 9 9 13 3 9 11 9 9 2
21 15 9 2 16 15 13 0 2 13 3 9 2 15 1 9 13 13 13 15 9 2
21 15 13 3 0 13 2 16 15 4 13 3 9 7 16 15 4 15 1 13 9 2
11 13 13 9 2 16 15 13 3 9 9 2
30 15 13 13 3 0 7 0 9 2 16 15 4 13 3 3 2 7 15 7 15 9 13 9 0 2 16 9 4 13 2
9 16 12 9 13 9 2 13 0 2
36 2 0 9 2 0 9 9 2 0 9 2 16 15 9 3 3 13 2 15 9 9 13 9 9 9 9 1 15 2 15 11 9 9 15 13 2
23 0 9 4 13 11 9 12 9 12 12 9 2 12 9 0 9 13 12 12 9 0 9 2
11 15 9 9 13 15 9 7 15 13 9 2
11 3 15 9 13 0 7 3 13 0 9 2
23 9 12 15 0 0 9 13 12 9 11 9 2 7 0 9 0 16 15 15 9 0 9 2
15 13 3 9 13 2 13 0 9 3 4 13 0 0 9 2
14 0 9 13 3 9 9 1 13 9 13 9 0 9 2
20 15 9 13 9 9 9 7 13 0 3 0 9 2 3 9 7 9 7 9 2
33 16 13 3 3 9 13 9 9 2 15 9 9 9 2 9 7 0 9 9 13 3 3 13 9 9 9 7 3 9 7 9 9 2
10 15 9 9 9 7 9 13 0 9 2
44 13 3 2 12 9 12 9 1 2 9 9 9 12 9 15 4 13 0 9 13 15 9 0 9 2 16 15 12 9 4 3 3 13 2 7 13 15 3 11 9 9 0 9 2
28 0 9 2 13 13 9 11 2 15 4 3 13 3 9 7 13 15 9 2 15 15 9 4 3 7 3 13 2
26 13 3 13 15 9 15 0 9 2 15 15 4 13 9 9 7 3 13 15 9 2 15 13 9 0 2
17 13 3 13 9 2 16 15 4 3 13 0 7 0 9 13 9 2
12 9 4 13 0 9 2 3 16 9 4 13 2
15 13 3 0 13 11 9 9 2 16 0 9 9 13 15 2
7 9 13 0 9 11 9 2
14 9 13 0 9 0 9 9 2 15 9 13 0 9 2
17 13 9 0 15 2 16 0 9 7 9 9 13 9 13 12 9 2
21 9 2 3 9 13 0 3 2 0 9 13 13 7 0 9 13 0 9 9 9 2
25 9 13 2 16 0 9 2 0 0 9 13 9 7 0 9 13 0 2 0 7 0 9 9 0 2
20 9 9 2 9 13 0 9 7 9 3 3 13 13 0 9 2 9 7 9 2
15 15 13 2 16 3 0 0 9 9 9 4 13 3 9 2
3 13 9 2
5 9 9 13 9 2
36 16 13 2 9 13 3 0 9 9 2 7 4 13 13 2 16 4 3 13 0 3 13 9 9 2 15 4 13 9 13 9 9 7 9 1 2
19 9 4 13 13 3 0 9 7 9 13 9 7 13 9 9 7 9 9 2
14 13 3 2 16 15 13 9 0 9 2 3 16 9 2
21 9 4 13 3 7 9 9 2 15 3 13 0 2 13 0 9 2 3 11 9 2
21 15 13 3 13 9 13 9 7 9 4 13 3 2 3 2 16 4 0 13 9 2
23 2 0 9 2 13 2 13 3 13 3 9 9 9 7 9 9 7 11 13 11 9 9 2
23 9 13 9 7 0 11 9 9 2 15 15 13 3 4 13 2 15 13 9 11 11 9 2
33 0 9 9 2 15 15 13 0 9 7 3 7 0 9 9 2 13 0 9 9 9 9 1 2 15 13 3 3 7 12 9 13 2
17 13 9 13 3 9 9 13 9 7 3 11 9 9 13 0 9 2
21 13 0 0 2 16 9 9 9 9 13 2 7 9 13 15 13 2 16 3 13 2
14 15 13 4 13 9 3 2 16 9 13 0 9 9 2
18 15 1 2 16 9 9 13 2 15 9 2 3 9 2 13 3 9 2
25 15 9 7 9 13 9 7 13 9 0 2 0 7 0 9 0 9 2 15 9 13 3 3 9 2
10 13 3 9 0 9 7 13 15 3 2
16 13 3 11 9 13 15 9 2 15 13 13 9 7 9 3 2
17 13 2 16 13 9 7 15 9 9 3 16 9 9 13 13 9 2
15 13 2 16 9 13 13 3 7 16 9 9 13 9 15 2
23 13 3 7 13 3 9 13 7 13 15 13 9 7 15 9 2 9 9 7 0 9 9 2
30 15 13 9 3 9 3 15 2 15 9 0 13 13 2 13 9 9 3 13 2 7 15 2 15 13 15 3 9 9 2
10 15 13 9 7 0 7 0 9 9 2
27 13 15 9 2 9 7 9 2 13 3 9 13 9 0 9 9 2 15 13 0 9 2 3 3 11 9 2
20 15 9 13 13 9 9 9 2 15 13 2 7 13 3 2 0 9 11 11 2
20 9 4 13 15 9 9 3 2 16 15 13 3 15 9 2 15 13 13 9 2
8 15 1 13 11 11 0 9 2
14 0 9 2 3 13 2 16 9 13 3 0 7 0 2
7 9 9 13 13 0 9 2
23 4 3 13 9 2 15 1 9 13 9 9 2 16 9 1 2 15 9 4 13 13 15 2
45 15 1 15 11 9 13 9 4 13 3 2 3 13 7 0 13 15 3 13 2 3 16 15 9 9 3 13 2 7 15 2 15 13 13 11 9 2 4 13 15 15 0 9 9 2
7 9 9 9 13 13 3 2
10 15 13 0 9 13 9 4 3 13 2
13 3 13 9 13 2 16 13 9 13 13 15 9 2
6 0 9 2 13 9 2
22 13 0 2 16 15 11 9 13 1 0 9 11 1 13 9 2 9 2 9 7 9 2
7 3 9 11 1 13 0 2
23 11 13 13 3 9 2 15 13 9 2 7 15 4 13 2 15 9 13 0 9 9 11 2
9 15 9 13 13 13 9 3 3 2
17 3 11 7 11 0 9 13 3 9 2 13 13 15 3 11 9 2
16 11 9 0 9 13 3 13 0 2 15 11 9 4 3 13 2
16 11 13 9 13 9 3 11 3 15 9 7 3 3 11 9 2
19 0 9 2 3 9 9 13 9 9 1 4 3 13 9 2 15 9 13 2
10 9 4 13 2 3 16 4 13 3 2
16 13 3 3 15 9 9 7 13 9 11 9 9 13 9 3 2
6 15 15 13 4 13 2
9 3 0 9 13 3 3 0 9 2
24 13 7 13 3 2 15 13 0 9 2 15 13 3 9 2 9 0 9 11 0 7 0 9 2
8 11 9 13 15 9 0 9 2
12 15 9 2 15 3 13 7 15 13 2 13 2
8 9 9 13 3 3 3 3 2
23 13 3 2 16 9 13 3 0 9 7 16 15 13 4 13 2 16 9 13 13 0 9 2
31 9 13 3 13 3 15 0 9 2 7 15 13 3 15 15 9 0 9 2 0 9 9 2 7 15 13 3 9 0 9 2
12 9 13 3 15 0 9 2 7 15 9 13 2
12 15 11 9 9 13 3 3 3 15 15 9 2
19 15 13 3 2 7 13 15 0 9 4 2 7 15 4 3 13 0 9 2
13 15 13 13 3 3 15 2 7 15 13 15 9 2
13 15 13 15 9 15 2 15 13 3 0 9 9 2
33 0 9 9 2 9 11 11 11 7 15 2 15 4 3 13 0 9 9 12 1 2 4 13 3 15 9 2 7 13 13 15 9 2
29 3 11 13 3 15 13 9 9 9 11 11 11 9 13 2 16 16 15 13 9 9 9 2 11 9 13 13 15 2
14 1 9 9 15 13 0 9 15 2 13 15 9 13 2
12 0 9 11 9 7 15 9 11 13 13 0 2
28 15 13 3 9 9 2 9 1 2 7 15 13 15 3 2 16 15 2 15 13 13 9 2 13 3 13 13 2
68 0 2 15 9 9 13 2 0 9 3 13 2 3 15 9 2 15 15 13 2 7 13 13 2 3 13 0 2 16 15 9 9 2 11 9 9 13 2 13 9 11 1 3 0 7 9 13 9 2 15 13 9 13 9 2 9 3 13 3 3 3 7 9 13 0 9 9 2
34 13 9 9 2 13 15 15 9 3 9 2 16 11 9 13 13 3 0 9 13 9 13 9 7 9 1 7 13 15 9 11 9 1 2
33 13 2 16 15 13 3 0 9 2 9 15 13 3 0 9 2 7 3 15 13 15 15 7 0 9 2 15 13 0 9 13 9 2
19 11 11 0 9 15 13 13 9 2 7 13 3 3 15 9 7 13 15 2
5 15 9 13 9 2
45 0 9 2 15 3 13 2 13 3 0 9 9 9 2 9 9 7 15 4 3 13 0 7 0 9 0 9 1 2 15 13 3 12 9 2 15 13 0 0 9 7 9 13 9 2
22 15 4 13 2 16 9 13 2 7 15 4 3 13 9 7 9 7 13 3 0 9 2
29 13 3 13 12 9 13 9 2 15 9 11 13 3 2 13 3 9 2 15 13 11 15 9 9 2 15 13 9 2
31 15 9 9 4 13 9 0 9 2 7 3 3 4 13 0 9 0 9 15 9 2 16 13 3 0 7 0 9 9 3 2
11 15 4 13 2 16 0 9 13 15 9 2
21 0 9 7 9 9 2 0 9 9 2 9 9 13 9 3 9 13 11 9 9 2
10 4 13 2 16 0 9 13 11 9 2
20 9 9 9 13 3 7 9 13 0 9 11 9 7 9 13 13 15 9 3 2
9 9 13 9 7 11 0 9 9 2
14 15 4 13 2 16 0 9 13 0 9 13 11 13 2
16 15 13 2 16 9 2 15 11 4 13 2 13 9 3 3 2
21 13 13 3 13 2 16 15 13 3 0 9 2 15 11 9 4 13 11 15 9 2
9 15 1 13 3 15 0 9 9 2
7 0 9 15 9 4 13 2
24 11 9 13 4 13 2 15 4 13 11 9 7 15 9 2 13 9 7 13 3 9 9 9 2
26 11 13 0 9 13 9 3 3 2 16 11 9 13 15 9 9 15 7 16 3 9 13 11 9 13 2
23 15 9 4 13 2 13 0 9 4 3 3 13 13 9 2 15 13 11 0 7 0 9 2
30 15 13 3 0 9 2 16 7 0 9 7 9 0 9 13 9 13 13 15 0 0 2 16 9 3 13 11 9 13 2
20 15 13 15 2 16 9 7 9 13 13 13 11 9 9 13 9 11 9 1 2
22 3 13 0 2 7 13 15 2 16 0 0 9 9 11 9 13 3 13 0 9 1 2
22 2 9 2 0 9 2 0 9 9 9 13 3 11 7 11 9 2 15 13 3 3 2
9 13 11 15 9 11 9 0 9 2
17 15 4 13 13 9 3 9 2 7 13 0 9 7 9 0 9 2
19 9 15 4 3 13 2 16 15 4 13 3 3 13 15 2 15 3 13 2
8 3 15 13 9 13 3 9 2
11 13 15 9 13 3 9 7 9 13 9 2
12 13 15 2 16 9 13 3 13 9 15 9 2
11 0 9 9 2 15 4 13 9 15 9 2
28 13 9 3 12 9 7 11 7 11 9 7 0 9 11 7 15 13 9 2 15 4 3 13 9 9 7 9 2
9 9 9 13 2 16 3 13 9 2
22 0 0 9 11 7 11 1 13 13 0 3 15 7 11 2 7 15 13 3 0 9 2
12 0 9 2 15 13 9 13 9 11 15 9 2
30 3 15 4 15 9 13 2 16 15 13 0 9 0 9 2 16 15 0 9 13 2 3 16 15 0 9 9 9 9 2
17 11 9 13 0 11 11 7 9 12 11 9 1 0 9 15 9 2
22 9 13 3 13 15 9 9 2 15 13 3 15 11 9 9 2 15 13 0 16 15 2
37 16 13 2 16 9 9 13 15 9 2 16 9 13 2 16 13 2 16 11 9 13 15 9 2 13 2 16 9 13 11 9 9 11 9 9 9 2
14 15 9 9 0 9 11 9 1 13 9 0 9 9 2
11 15 13 0 0 9 2 0 9 9 9 2
9 15 13 9 9 3 0 0 9 2
9 13 2 16 15 4 13 15 9 2
21 3 15 9 0 9 11 9 2 11 9 9 9 7 9 13 9 13 3 0 9 2
26 0 9 2 0 9 9 2 3 13 13 9 9 2 15 15 4 15 9 1 13 15 3 0 9 9 2
14 13 3 13 9 11 9 2 15 15 4 15 9 13 2
12 9 13 0 2 16 11 9 4 13 0 9 2
15 13 3 2 16 11 4 13 9 3 3 9 7 9 9 2
30 3 13 3 9 2 15 15 9 2 15 13 2 16 15 4 13 9 2 3 3 13 0 7 0 9 3 13 9 9 2
13 15 4 3 13 9 2 7 3 15 15 9 13 2
38 15 4 13 15 9 2 13 9 9 2 15 1 15 9 0 9 13 15 11 9 12 9 3 16 15 15 2 15 3 13 15 2 16 15 13 15 9 2
23 13 2 16 15 4 13 2 16 9 13 3 3 0 9 2 15 13 9 2 9 7 9 2
31 13 9 15 9 2 16 9 0 9 13 3 9 9 2 15 9 13 0 9 2 7 16 9 9 13 0 9 15 9 9 2
14 9 13 0 9 13 13 15 9 13 9 7 13 15 2
13 0 9 9 2 3 3 13 15 9 9 13 9 2
19 15 15 13 3 9 0 9 7 3 3 9 13 15 9 2 9 7 3 2
17 15 13 15 2 16 9 13 3 3 15 2 16 9 13 3 3 2
24 13 15 9 3 9 2 15 13 9 13 9 9 9 15 9 9 2 15 15 13 13 9 13 2
32 15 9 13 9 2 15 15 15 4 13 9 1 2 7 13 15 9 3 15 2 16 9 11 13 0 15 2 15 15 4 13 2
13 15 9 13 3 3 15 9 2 15 13 15 9 2
43 0 4 13 9 12 2 15 13 0 9 13 9 9 0 3 2 7 9 12 7 12 2 15 13 9 0 9 0 9 2 15 4 13 0 9 3 16 9 13 9 7 9 2
26 3 4 13 15 15 9 2 15 2 13 9 2 9 13 0 9 0 9 7 13 9 7 9 0 9 2
17 13 13 3 3 7 11 7 0 9 2 9 7 9 15 13 9 2
39 15 9 9 13 3 13 15 9 9 7 3 9 2 15 4 13 11 9 9 9 7 2 16 3 13 2 7 9 3 9 13 9 9 9 7 9 9 9 2
6 9 9 13 9 9 2
20 3 3 13 0 2 13 4 13 9 12 7 12 2 15 13 9 0 9 9 2
13 3 3 13 13 3 15 9 2 15 11 13 3 2
6 3 9 9 0 9 2
23 13 2 16 15 13 9 2 15 13 3 9 7 15 15 3 9 2 7 9 9 4 13 2
16 15 9 4 13 13 9 2 15 13 9 9 9 13 9 9 2
12 9 11 2 9 13 2 16 9 13 9 3 2
18 3 3 3 13 9 13 9 13 9 9 13 9 13 3 9 9 2 2
29 13 15 2 16 9 13 9 2 15 4 13 3 15 9 2 7 9 13 3 4 13 2 16 9 13 15 0 9 2
18 15 4 13 9 2 16 4 13 2 16 3 13 2 0 9 7 9 2
23 9 11 2 15 9 15 4 13 2 16 9 12 13 0 16 15 9 2 13 4 15 13 2
11 13 3 0 13 9 1 15 13 13 9 2
31 15 9 9 12 3 13 3 2 16 15 13 15 0 9 2 15 13 9 3 13 9 1 2 4 13 15 9 13 9 9 2
11 13 15 2 16 13 15 13 9 3 3 2
28 9 12 9 15 4 13 15 2 16 9 13 3 0 2 9 2 9 15 13 9 2 7 9 9 13 3 0 2
7 0 9 11 4 13 9 2
17 15 0 9 4 13 9 2 16 15 13 0 2 7 9 7 9 2
22 9 9 13 15 9 13 9 2 15 1 9 13 13 9 7 13 9 3 16 13 3 2
11 15 13 13 9 9 13 3 15 0 9 2
34 15 13 3 13 2 16 0 9 4 13 15 9 13 9 2 9 7 9 7 16 15 9 13 0 2 16 15 9 13 9 4 13 9 2
27 15 9 2 15 9 9 13 15 9 3 3 3 2 16 9 9 13 13 3 9 13 9 2 13 4 13 2
52 3 3 7 0 9 7 11 9 9 9 9 4 13 9 2 16 15 9 9 13 13 15 9 16 11 9 9 2 13 9 0 9 2 16 16 15 9 4 13 2 15 4 13 9 7 9 3 15 9 9 13 2
23 11 9 9 1 13 9 13 0 9 13 9 0 9 15 9 9 1 2 15 4 3 13 2
17 3 13 3 3 2 4 3 13 15 9 2 16 9 13 0 9 2
13 15 9 9 13 0 9 4 13 9 7 15 9 2
32 15 9 13 9 2 15 4 13 0 9 15 9 2 16 9 9 13 0 3 0 9 9 2 15 13 0 9 7 9 13 9 2
6 13 3 15 9 9 2
21 15 9 4 3 13 15 9 9 9 2 15 9 13 9 9 13 0 9 9 9 2
20 0 9 2 0 9 9 2 3 13 3 13 2 16 0 9 13 0 9 9 2
13 9 4 13 3 9 13 13 0 9 11 9 1 2
26 13 13 15 3 3 2 16 9 13 13 2 16 9 9 2 15 13 3 2 13 0 13 3 13 9 2
19 13 3 2 16 11 9 13 9 3 2 16 9 13 3 7 13 9 13 2
30 15 9 13 3 3 13 15 13 15 9 9 7 13 9 11 7 0 9 1 13 9 7 15 2 0 9 9 2 9 2
19 9 13 0 9 2 15 9 13 9 13 9 0 7 9 9 9 3 9 2
23 0 9 13 9 13 15 0 9 9 12 2 7 15 9 0 11 13 3 12 12 9 3 2
27 9 13 9 13 9 9 7 13 11 0 9 12 1 9 9 9 2 9 7 9 0 9 2 9 7 9 2
24 13 0 9 2 16 15 9 4 13 12 9 9 2 15 13 9 9 13 13 13 9 9 1 2
24 16 15 9 9 13 12 12 9 2 15 9 13 3 12 12 9 9 7 9 13 9 3 11 2
14 9 9 1 9 9 4 13 9 13 9 3 12 9 2
12 0 9 9 2 13 3 3 0 9 9 9 2
24 9 11 7 11 1 13 12 2 16 9 13 11 12 9 9 9 7 9 13 13 9 9 1 2
16 3 16 9 0 9 9 2 13 3 9 2 15 9 4 13 2
25 13 3 15 9 2 16 9 13 3 2 16 9 13 13 2 15 12 9 9 13 7 0 9 13 2
11 13 3 0 15 2 16 15 9 13 13 2
13 11 13 15 2 13 0 9 13 9 11 0 9 2
17 13 3 0 9 2 15 13 9 2 15 1 15 9 4 13 9 2
4 15 13 3 2
7 9 13 3 9 13 9 2
10 9 9 13 0 9 2 15 9 13 2
22 3 13 3 9 11 11 7 9 11 9 7 13 15 15 2 16 15 9 9 13 9 2
6 0 9 9 4 13 2
3 13 9 2
8 9 11 13 9 0 9 13 2
12 11 9 4 13 0 9 13 0 7 0 11 2
10 3 15 12 9 9 9 13 0 11 2
17 11 13 0 15 9 1 2 15 9 13 0 9 3 13 9 1 2
22 11 13 0 9 13 9 1 2 7 9 13 13 0 2 9 3 3 13 7 0 9 2
13 3 15 4 13 0 9 2 16 15 9 13 13 2
42 15 9 4 13 0 9 2 9 7 9 0 9 7 9 9 9 9 9 2 15 13 15 13 9 7 9 2 7 0 2 8 8 8 8 2 0 9 0 0 9 9 2
19 9 9 4 13 1 0 9 9 2 16 15 13 9 13 3 0 7 0 2
40 13 3 2 16 9 13 9 13 3 15 9 3 12 9 9 2 16 15 9 4 13 2 16 15 12 0 9 4 13 9 2 15 13 3 0 9 11 9 9 2
18 2 9 2 0 9 2 13 3 13 15 2 16 13 9 12 0 9 2
9 13 13 9 3 9 2 9 2 2
5 3 0 9 13 2
16 2 9 2 2 13 2 16 11 0 9 4 13 3 9 2 2
6 2 0 9 13 2 2
11 0 9 9 2 13 13 9 13 9 11 2
15 3 15 4 13 2 16 15 13 9 13 3 13 3 9 2
22 13 9 11 2 16 13 15 0 9 4 3 13 0 9 9 1 2 4 4 13 9 2
20 15 13 3 15 2 16 9 2 3 11 13 9 2 3 12 9 13 15 9 2
20 13 9 1 2 15 11 11 9 13 13 15 9 2 15 15 9 9 4 13 2
32 13 0 9 2 16 11 11 9 13 0 9 0 9 7 13 3 0 2 16 9 9 1 13 11 9 9 13 7 13 0 9 2
24 13 15 13 7 13 13 9 9 2 16 15 4 13 2 16 11 13 13 3 0 9 15 9 2
49 0 9 2 15 15 13 11 0 9 9 13 9 1 2 16 13 3 3 2 16 15 9 13 2 16 15 9 2 15 13 15 9 2 4 13 15 9 3 0 9 2 15 4 13 12 9 0 9 2
33 9 13 0 9 13 3 15 2 16 3 15 0 9 9 13 13 2 7 16 13 2 16 15 13 2 9 2 9 2 13 3 0 2
27 13 15 9 2 16 15 4 13 15 9 3 0 9 2 13 3 3 0 9 2 15 4 13 3 0 9 2
29 0 9 2 0 9 2 13 3 9 11 11 9 2 15 13 0 9 7 15 13 15 9 0 9 7 9 13 9 2
34 13 3 2 13 9 4 13 3 9 7 0 9 9 2 7 16 15 13 9 13 0 9 13 9 2 15 9 15 0 0 9 4 13 2
20 11 11 9 13 0 15 13 9 9 7 3 3 2 16 15 9 13 13 9 2
5 15 13 9 9 2
9 3 13 9 0 9 13 0 9 2
5 3 15 4 13 2
17 0 9 0 9 4 3 13 15 9 13 12 9 15 9 13 0 2
7 13 4 13 0 9 9 2
14 15 13 0 9 0 13 12 9 2 15 13 9 9 2
19 3 13 3 3 9 13 15 3 9 13 9 13 0 9 7 15 0 9 2
3 0 9 2
15 13 3 13 9 9 9 9 2 15 15 3 0 9 13 2
17 13 13 2 16 15 9 13 0 9 2 15 13 3 3 4 13 2
7 0 9 9 4 3 13 2
10 3 15 9 9 13 3 3 13 0 2
23 15 1 3 13 9 9 0 9 13 0 2 16 13 13 9 9 2 7 13 15 0 9 2
25 11 9 0 9 13 1 9 2 7 3 0 9 9 13 9 7 0 9 9 9 2 15 3 13 2
11 13 2 16 9 13 9 4 13 9 0 2
11 9 4 13 9 13 9 9 12 9 9 2
12 9 4 9 9 13 13 15 3 9 12 9 2
16 15 13 15 9 9 11 11 9 9 11 0 9 12 13 9 2
13 15 13 15 2 16 15 9 13 9 9 4 13 2
25 4 3 9 1 13 2 16 13 13 3 9 15 0 9 3 0 9 9 4 13 0 9 0 9 2
20 13 3 13 2 16 9 13 0 15 2 16 9 7 9 4 13 0 9 9 2
16 9 9 13 3 0 9 1 0 9 2 7 9 7 9 9 2
15 0 9 2 9 13 9 0 9 12 13 3 3 12 9 2
12 12 9 3 9 13 9 13 9 9 11 9 2
8 13 3 12 9 9 15 9 2
18 2 13 9 0 9 9 2 16 15 13 15 9 1 13 9 9 9 2
34 11 2 15 4 13 0 2 13 3 9 9 2 15 4 13 15 9 0 9 2 9 2 15 15 13 9 0 9 7 15 15 13 9 2
16 0 9 15 9 13 9 2 15 13 3 0 13 0 0 9 2
18 9 12 13 9 9 13 9 13 9 9 9 9 13 15 9 9 1 2
26 13 13 3 3 15 2 16 9 9 13 9 11 13 9 9 13 0 9 2 16 9 9 13 9 1 2
9 13 3 13 9 13 15 9 2 2
10 13 15 0 9 13 3 15 0 9 2
17 4 0 9 9 13 13 9 15 9 7 13 3 9 9 1 9 2
6 15 13 3 15 9 2
12 3 15 2 16 9 9 13 16 9 0 9 2
8 15 13 13 3 15 9 9 2
8 15 13 3 13 15 9 9 2
28 9 9 12 7 9 12 0 9 13 2 16 9 13 0 9 9 2 16 15 13 3 2 16 15 13 16 3 2
13 12 9 12 9 13 9 3 13 13 9 13 9 2
23 15 9 13 3 3 0 9 9 9 12 2 7 3 2 9 12 2 9 13 13 0 9 2
12 0 13 3 2 16 9 3 13 13 9 1 2
27 15 3 0 9 2 15 13 9 9 2 4 13 13 11 9 2 15 13 9 7 9 2 9 7 9 9 2
33 15 13 3 3 2 13 11 9 2 15 15 9 13 3 2 13 9 0 9 2 7 3 15 9 13 0 9 2 15 13 11 9 2
29 15 15 9 13 9 13 3 0 9 2 7 3 9 2 15 15 4 13 15 9 2 4 15 1 13 3 3 0 2
10 0 9 4 13 3 3 15 9 9 2
8 15 3 12 9 13 3 0 2
22 12 9 13 9 9 15 0 0 15 2 13 15 9 13 0 9 2 4 13 0 0 2
33 15 3 0 2 15 9 1 13 0 9 13 9 1 13 2 13 9 1 2 15 2 16 2 9 13 13 9 2 9 7 9 2 2
18 15 13 3 1 9 0 9 1 2 3 15 9 13 3 12 9 9 2
8 15 9 0 9 13 3 9 2
45 3 2 9 12 13 9 1 9 7 15 9 13 0 9 2 16 15 9 13 9 1 9 15 2 16 15 13 0 9 7 15 2 16 3 3 16 9 13 2 15 9 13 0 9 2
18 15 13 3 9 0 9 2 3 9 9 2 13 15 9 13 15 0 2
12 15 9 9 13 15 15 2 16 13 15 9 2
19 15 13 2 16 15 9 9 9 1 9 0 9 13 2 13 0 9 0 2
6 9 13 2 13 13 2
19 0 9 13 2 3 0 9 13 9 9 2 16 9 13 4 13 0 9 2
43 13 0 2 16 0 9 3 13 0 7 15 9 7 16 9 2 15 4 13 3 15 9 2 15 9 4 13 2 13 0 15 13 0 9 2 16 13 3 13 0 9 9 2
6 9 4 13 0 9 2
7 3 13 3 13 3 0 2
10 13 3 13 9 7 9 0 9 11 2
10 13 15 13 0 9 15 9 9 9 2
35 13 15 2 16 9 9 4 13 9 9 2 16 11 13 13 3 2 15 4 13 7 13 2 16 9 13 7 9 11 9 2 12 2 13 2
25 9 12 9 12 9 13 2 16 9 9 1 15 13 4 3 13 1 9 9 13 9 12 7 12 2
17 16 9 13 13 3 0 13 2 9 13 11 9 13 9 11 9 2
21 2 0 9 2 0 9 2 3 13 13 9 9 12 9 2 15 0 13 0 9 2
16 13 13 2 15 3 0 9 9 13 2 13 15 4 13 9 2
13 15 4 9 13 0 7 3 0 13 3 0 9 2
6 0 9 13 11 9 2
32 3 16 13 15 3 2 13 13 2 3 9 4 13 3 13 12 0 9 9 9 15 2 11 9 2 11 9 7 0 11 9 2
32 0 9 15 9 13 9 13 3 3 15 2 7 3 13 13 0 2 15 13 15 0 9 2 7 3 3 2 3 15 9 13 2
14 13 0 2 16 9 9 4 13 15 15 15 12 9 2
16 13 13 12 9 11 9 7 15 2 3 4 13 11 9 3 2
27 3 16 11 0 9 13 2 3 15 9 2 16 13 11 9 2 13 3 3 9 7 9 2 15 4 13 2
45 9 15 13 3 3 0 9 11 0 9 2 15 13 3 15 2 3 9 13 2 7 11 13 0 9 9 2 7 15 2 3 9 13 2 7 9 9 2 7 15 2 3 9 13 2
10 3 13 13 9 7 9 9 0 9 2
28 0 9 13 3 0 9 2 3 9 2 13 15 9 2 16 3 9 13 7 9 7 9 13 4 13 3 0 2
18 15 13 4 9 13 3 13 9 9 13 15 2 3 4 13 9 9 2
13 0 15 9 9 9 11 9 13 3 0 0 9 2
22 15 13 3 13 15 2 7 3 13 15 2 16 15 4 3 13 9 7 0 9 1 2
10 15 4 13 9 7 13 0 9 1 2
10 13 13 2 15 9 4 13 15 9 2
13 15 13 12 9 7 9 13 9 9 2 15 13 2
37 16 3 13 0 2 16 12 9 13 0 9 9 11 9 1 13 9 2 3 13 0 2 16 13 13 9 13 9 9 11 9 1 9 0 9 1 2
15 13 3 13 0 9 2 13 3 13 2 3 15 13 9 2
18 9 13 3 0 9 9 9 2 15 13 15 0 0 2 16 13 9 2
24 13 0 2 16 13 15 2 3 15 3 13 9 4 13 3 3 9 7 3 9 4 13 9 2
15 0 9 13 3 9 2 0 2 9 2 2 15 13 3 2
6 15 13 9 11 9 2
17 0 9 9 2 3 13 9 9 7 3 15 9 7 0 9 9 2
12 13 13 2 4 9 13 15 11 9 13 9 2
12 16 13 2 11 0 9 9 4 13 9 9 2
25 13 0 13 2 15 4 13 2 16 11 9 13 4 3 13 11 9 2 3 16 15 15 9 13 2
51 9 2 13 15 3 0 7 0 2 13 3 3 0 9 7 15 9 9 2 15 13 13 15 0 9 1 2 15 0 9 7 0 9 13 13 9 2 16 15 13 3 15 9 0 9 7 9 9 9 1 2
12 9 13 13 9 9 7 0 7 0 9 1 2
2 0 2
31 2 2 9 2 11 9 13 9 13 3 9 2 15 13 15 9 2 7 13 9 2 15 13 2 16 13 15 9 0 9 2
11 13 0 2 16 9 9 4 13 0 9 2
37 16 9 13 2 16 2 0 7 9 2 0 9 7 9 3 13 2 13 3 13 3 11 9 9 9 2 2 4 3 13 2 13 11 13 3 9 2
31 9 13 3 2 11 11 2 9 9 9 13 4 13 15 15 9 2 15 13 13 0 9 13 9 0 9 9 9 13 9 2
37 13 0 9 13 9 0 9 9 9 2 15 15 9 13 13 7 13 9 7 9 9 13 9 7 0 9 0 9 13 7 9 13 9 13 9 9 2
18 15 9 4 13 9 13 0 9 13 7 13 9 3 7 13 13 9 2
31 0 9 2 9 9 9 13 3 0 2 16 9 9 1 9 12 15 4 13 12 9 2 16 16 9 12 15 13 3 12 2
35 15 9 13 3 9 9 0 9 2 7 7 9 13 9 2 16 9 4 13 11 9 1 9 0 9 2 3 9 9 12 7 12 9 1 2
49 3 13 11 9 9 13 3 15 9 2 16 9 13 13 3 15 9 2 13 9 3 9 7 9 2 7 13 3 0 0 9 2 15 13 15 9 2 15 13 13 9 9 3 3 3 7 3 3 2
17 3 15 9 2 15 13 13 9 9 2 13 3 3 0 13 15 2
6 15 13 15 0 9 2
8 0 1 13 15 12 0 9 2
21 3 15 13 15 2 16 9 4 13 13 3 9 2 15 9 13 3 0 0 9 2
13 13 2 16 15 13 3 2 16 9 9 13 9 2
20 9 15 13 13 3 3 2 16 9 4 13 0 9 7 16 9 13 13 9 2
20 7 9 9 11 13 9 9 2 15 4 4 13 2 16 3 3 4 13 9 2
13 0 9 13 9 2 9 9 13 4 15 9 13 2
21 15 13 3 9 12 13 0 9 9 13 9 2 15 9 9 3 13 9 9 1 2
32 16 13 9 0 9 2 7 9 2 15 13 2 13 2 3 2 15 13 9 13 9 3 12 9 13 2 16 12 9 15 13 2
40 7 3 0 9 13 9 2 15 9 13 4 13 3 7 15 4 13 3 3 2 16 9 13 9 9 4 13 13 9 13 9 9 9 2 15 4 3 4 13 2
13 3 13 3 11 0 9 9 13 9 9 12 9 2
21 13 3 2 16 9 13 4 13 3 2 16 15 13 9 15 9 3 0 9 1 2
14 3 9 13 0 9 2 3 9 0 9 2 0 9 2
20 3 13 9 9 2 16 13 13 13 9 2 7 3 3 13 9 15 3 9 2
15 3 13 3 11 9 9 2 7 11 4 3 13 15 3 2
26 0 9 2 0 9 9 11 2 0 9 9 11 2 11 9 13 9 2 7 15 13 0 15 9 9 2
12 15 9 4 3 12 9 9 13 13 3 11 2
31 15 15 2 15 3 13 15 9 2 13 3 0 13 2 15 9 15 13 2 16 3 13 9 1 13 9 4 13 1 9 2
15 15 13 13 3 9 13 2 16 9 13 15 9 9 1 2
14 9 13 9 13 9 3 3 0 9 16 0 9 9 2
14 0 9 13 3 4 13 0 9 16 9 7 3 9 2
10 15 4 13 9 2 16 11 13 9 2
17 16 9 9 11 13 2 11 13 0 9 9 9 7 3 9 9 2
26 11 9 4 13 0 2 0 9 15 4 13 2 16 9 3 3 13 7 3 16 0 9 15 9 13 2
17 15 4 4 13 15 2 16 9 13 2 16 3 12 9 9 13 2
13 13 0 9 9 11 13 9 2 15 13 3 0 2
22 11 0 9 12 9 4 3 3 3 13 2 16 13 15 9 2 13 3 0 9 9 2
21 13 0 9 2 16 13 9 0 9 2 16 9 7 9 7 9 7 0 9 9 2
9 9 15 4 13 9 13 0 9 2
12 3 11 1 13 9 9 9 13 15 9 9 2
19 9 13 3 3 0 9 9 2 3 9 13 9 2 13 15 9 13 9 2
5 3 9 13 13 2
20 11 9 9 9 1 13 3 9 9 2 3 13 9 11 9 7 3 15 15 2
11 13 3 2 16 13 0 9 0 9 9 2
23 9 4 13 3 2 3 7 3 2 7 11 9 4 13 9 13 9 9 2 15 3 13 2
13 2 13 11 9 9 0 9 12 13 9 3 13 2
19 0 9 7 9 2 3 3 9 13 13 9 0 9 13 9 0 9 9 2
21 0 15 9 13 13 15 9 2 7 15 9 3 0 13 15 13 15 0 0 9 2
23 13 3 15 9 0 2 15 4 13 1 0 9 7 15 4 3 13 15 9 0 9 9 2
11 13 9 2 15 13 11 9 11 9 9 2
20 13 13 15 15 0 9 9 2 3 9 13 0 9 13 3 7 0 7 0 2
15 3 4 3 13 12 9 2 16 0 9 13 3 0 9 2
22 13 3 13 12 0 7 0 0 9 2 11 9 11 7 11 2 7 15 9 7 9 2
13 3 15 13 9 13 3 9 3 13 0 9 1 2
32 3 13 9 11 9 11 11 11 2 0 9 9 1 2 15 13 3 9 12 2 16 11 13 13 3 2 16 15 13 13 3 2
12 15 2 11 11 7 11 11 13 9 3 3 2
19 16 11 4 13 3 3 2 4 13 12 9 7 0 9 0 7 0 9 2
24 13 13 1 3 9 3 11 11 2 11 11 2 11 11 2 11 11 11 7 11 11 11 9 2
16 3 15 4 13 0 9 9 13 11 11 9 3 12 9 9 2
42 15 4 13 0 9 2 7 4 13 13 0 9 15 9 2 3 3 15 1 2 16 4 13 3 0 9 7 0 9 13 9 2 15 13 11 9 7 15 9 0 9 2
10 15 3 9 0 9 13 13 12 9 2
33 15 13 15 0 9 15 0 9 2 15 4 3 15 9 13 2 0 9 2 0 0 11 11 9 2 15 13 13 3 9 3 3 2
11 13 0 9 9 2 15 13 15 0 9 2
15 9 2 9 7 9 13 3 0 9 16 3 15 9 1 2
6 9 9 4 13 3 2
13 9 7 9 0 9 13 0 16 3 15 9 1 2
7 3 15 4 13 9 3 2
15 13 1 9 2 15 0 9 13 7 9 2 3 0 9 2
17 16 15 13 9 13 11 0 3 13 9 9 2 15 13 0 9 2
18 13 4 13 9 15 2 16 13 9 11 9 15 15 13 9 3 3 2
10 13 3 9 15 2 15 13 15 9 2
7 15 4 13 15 3 9 2
8 0 7 0 9 4 13 9 2
8 13 9 7 11 9 0 9 2
23 3 9 9 2 3 3 3 9 2 15 13 9 2 13 4 13 15 2 16 13 13 9 2
15 3 0 9 13 3 9 2 7 15 9 4 13 0 9 2
20 0 9 13 15 0 2 16 13 11 9 15 16 3 0 9 7 0 9 9 2
27 0 11 13 15 0 9 2 3 15 2 15 13 3 3 13 9 2 7 15 13 13 1 9 0 11 1 2
6 9 4 13 0 15 2
17 15 4 13 15 0 9 11 9 9 3 2 16 15 13 0 9 2
12 15 13 13 3 9 2 7 3 15 9 0 2
25 0 0 9 7 15 15 9 2 0 11 11 2 13 15 3 2 2 11 13 15 0 9 9 2 2
27 15 13 3 15 2 13 15 4 13 3 0 9 7 9 2 7 9 2 15 13 15 7 15 15 9 9 2
79 11 13 13 3 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 7 3 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 7 11 2
13 0 11 4 13 3 3 15 0 7 0 9 9 2
20 11 9 13 13 13 0 2 0 9 9 2 2 15 11 9 11 11 3 13 2
17 16 13 0 9 13 1 11 9 9 1 2 15 13 16 13 9 2
8 13 2 16 9 13 15 0 2
22 15 9 13 0 2 7 15 0 9 0 9 13 9 2 15 3 0 11 4 15 13 2
20 9 4 13 15 2 16 9 9 13 3 7 3 13 3 16 9 9 9 9 2
13 13 0 0 9 2 2 8 8 8 8 8 2 2
5 15 9 13 9 2
9 0 9 7 9 2 9 13 0 2
8 15 4 13 15 9 13 9 2
8 13 15 9 9 7 15 9 2
7 15 4 13 15 9 3 2
9 15 13 0 2 7 3 0 9 2
10 15 9 13 0 12 7 9 9 13 2
5 15 13 9 15 2
19 15 9 13 15 7 15 15 2 15 13 0 9 13 0 9 2 11 9 2
4 7 3 9 2
3 2 9 2
25 0 9 2 13 3 3 3 13 0 9 9 1 9 11 11 9 7 3 13 13 9 11 11 9 2
33 0 9 2 15 15 15 9 4 13 2 7 9 11 11 13 15 0 9 2 15 4 13 3 9 2 13 12 9 2 15 13 9 2
10 3 2 9 13 9 11 9 9 9 2
14 0 9 2 15 9 13 2 13 9 9 0 9 9 2
47 0 2 7 15 13 0 9 3 2 15 13 3 9 2 15 13 7 0 9 7 9 1 7 3 3 3 15 11 9 9 2 15 9 13 11 2 7 3 15 9 2 15 0 9 13 3 2
32 15 13 15 2 16 15 4 13 15 9 3 3 9 2 15 4 13 7 11 9 1 9 1 7 3 11 9 7 0 9 1 2
38 9 11 11 13 15 2 16 9 13 13 15 0 9 2 15 13 13 15 0 9 2 7 15 13 3 0 9 7 15 13 11 9 0 9 7 0 9 2
7 15 1 15 13 15 9 2
10 15 9 13 15 2 16 15 13 9 2
26 15 13 13 9 2 15 13 13 9 2 15 13 15 16 9 0 9 7 0 9 2 15 3 4 13 2
18 15 13 13 3 15 9 2 15 0 0 7 0 9 1 13 9 13 2
7 15 13 13 0 9 0 2
58 15 13 13 2 15 13 15 1 2 15 13 9 0 9 1 2 7 0 9 1 2 15 13 2 16 15 13 0 9 7 16 11 7 11 3 13 3 7 11 3 13 9 2 15 15 9 4 3 13 7 3 15 13 9 1 11 9 2
7 15 13 3 15 9 1 2
12 15 13 2 16 0 7 0 9 9 3 13 2
7 15 13 13 3 9 15 2
9 15 13 13 9 0 9 7 9 2
10 4 13 15 2 16 4 13 9 9 2
5 3 13 13 15 2
9 13 11 9 9 2 15 13 0 2
5 15 13 13 9 2
9 15 13 15 1 13 11 13 9 2
9 13 2 16 15 4 13 13 9 2
11 3 9 13 15 2 15 13 15 9 9 2
15 13 0 7 0 9 2 9 2 15 13 13 11 9 9 2
12 13 3 0 9 2 15 11 11 11 9 13 2
4 15 13 0 2
6 15 13 13 15 3 2
14 15 13 3 13 15 9 2 13 3 9 9 9 11 2
10 15 13 3 15 2 15 15 3 13 2
18 15 13 13 15 15 2 15 4 13 2 15 13 0 9 2 0 9 2
5 15 15 13 15 2
27 13 3 0 2 16 13 3 3 0 9 2 15 13 3 3 3 16 3 15 9 2 15 4 13 15 1 2
4 0 9 9 2
12 3 13 9 9 9 12 9 2 15 13 9 2
13 9 7 9 1 13 9 2 15 9 13 13 3 2
15 15 4 3 9 13 2 16 9 7 9 9 13 13 15 2
21 13 2 16 9 13 3 9 2 7 15 9 13 3 9 2 7 15 9 13 15 2
26 9 13 0 2 16 16 3 13 0 9 2 15 2 15 4 3 13 0 9 2 13 3 1 13 9 2
6 9 4 13 9 9 2
38 15 9 13 2 16 9 13 9 3 3 2 7 3 13 3 0 15 2 16 3 9 9 2 15 13 3 13 15 0 9 2 9 9 13 3 3 3 2
19 15 9 13 15 9 1 2 7 15 13 15 2 16 15 13 13 15 9 2
15 13 15 9 2 16 13 0 13 15 3 2 16 4 13 2
33 3 9 9 4 13 3 2 16 15 13 3 9 9 9 2 16 9 13 0 9 13 9 7 9 2 9 13 9 3 15 9 9 2
30 15 13 13 9 13 0 9 2 7 15 13 2 16 15 9 2 15 15 13 13 2 13 3 13 9 13 3 9 9 2
25 0 9 2 0 9 9 2 13 9 9 11 11 1 13 15 9 13 9 2 15 13 3 15 9 2
21 15 9 13 9 9 9 7 9 0 3 13 15 3 0 9 2 0 7 3 0 2
33 15 9 9 13 16 3 15 2 16 0 9 13 0 2 9 13 0 9 9 2 15 3 13 0 9 2 15 13 0 9 15 9 2
25 15 2 16 13 9 3 9 2 15 13 9 2 16 13 9 3 9 2 4 9 1 13 15 9 2
12 0 0 9 4 15 9 13 3 0 0 9 2
17 15 13 3 13 3 3 9 2 16 13 3 0 9 13 9 9 2
18 13 0 2 16 9 13 9 13 9 7 9 2 15 3 3 13 9 2
26 3 4 3 13 2 16 0 9 4 13 15 1 2 16 13 3 13 15 0 7 0 9 13 9 9 2
11 0 9 0 9 1 15 9 13 4 13 2
30 15 9 2 15 13 3 9 0 0 9 9 13 3 3 3 3 13 7 13 0 9 9 13 3 0 9 13 9 9 2
20 15 13 3 15 9 2 7 13 0 13 3 7 13 15 3 7 13 9 9 2
61 15 9 0 4 13 15 2 16 3 2 16 0 9 13 2 13 0 0 0 9 2 15 9 0 9 13 1 13 9 2 15 0 0 9 7 9 13 0 13 2 3 13 2 0 7 13 9 13 0 9 0 9 0 9 7 9 0 9 9 9 2
17 13 13 0 9 9 9 13 9 13 0 9 2 15 15 13 15 2
12 3 13 9 13 13 13 3 9 7 0 9 2
18 2 11 2 0 9 9 2 15 13 0 9 2 15 13 15 9 9 2
17 0 9 9 9 13 7 13 9 9 13 13 3 9 13 0 9 2
14 15 13 4 13 15 9 9 2 16 9 13 4 13 2
16 3 3 3 9 9 13 9 13 4 13 2 7 15 13 13 2
13 9 2 15 13 15 9 9 9 9 2 13 0 2
18 0 9 13 15 13 15 9 9 7 13 2 16 9 9 9 13 3 2
31 0 9 2 15 9 13 3 3 0 9 13 9 0 9 1 15 2 16 9 13 3 0 0 13 2 16 15 13 9 9 2
11 3 13 13 9 1 2 7 15 13 9 2
80 0 9 13 3 0 9 2 16 13 11 11 9 0 0 9 2 9 9 1 2 7 13 11 9 13 0 0 9 13 2 15 13 3 0 0 2 16 15 13 9 11 11 11 11 9 13 9 2 7 3 13 2 16 9 13 15 13 9 2 15 9 4 13 13 3 2 13 3 11 9 7 11 11 13 11 11 7 11 9 2
17 0 9 2 13 3 13 13 13 0 9 2 15 3 13 9 9 2
41 2 9 2 16 9 0 9 0 9 9 13 9 7 9 2 13 0 2 16 11 9 13 15 0 0 9 9 13 0 9 2 16 15 9 9 9 13 0 9 15 2
18 3 11 9 4 3 13 9 13 9 9 12 9 13 9 13 0 9 2
40 13 3 0 13 3 15 2 16 15 9 0 9 4 13 0 9 13 9 7 9 7 0 9 2 9 11 7 11 7 11 9 2 9 9 0 7 0 9 9 2
13 3 9 13 15 2 13 9 9 13 3 15 9 2
63 3 13 0 2 16 9 13 0 9 7 3 9 0 9 3 0 9 9 2 0 9 3 0 9 7 9 0 9 2 0 9 7 9 9 2 9 9 7 0 7 0 9 9 7 9 9 9 9 13 9 2 15 13 3 0 9 9 9 0 9 9 13 2
11 2 9 2 0 9 2 4 13 13 9 2
5 15 9 13 3 2
5 15 13 3 3 2
12 15 13 3 2 7 13 2 16 13 15 9 2
32 0 9 2 15 9 13 0 9 7 15 9 13 15 0 9 2 9 2 3 3 16 15 4 13 2 13 3 9 15 9 9 2
18 0 9 9 3 9 13 0 7 3 15 9 2 16 15 4 13 9 2
15 15 9 13 13 9 15 9 2 15 13 0 9 9 1 2
23 13 13 3 15 9 2 16 13 0 9 0 9 11 2 15 9 9 11 9 13 15 0 2
9 15 9 1 9 9 13 9 0 2
14 3 9 11 13 9 3 0 9 2 15 13 9 1 2
9 11 9 13 3 3 3 0 9 2
53 16 13 15 0 9 3 9 7 13 9 2 13 9 13 9 13 15 2 15 13 3 4 13 2 16 3 13 3 9 0 9 13 9 0 2 9 2 15 0 9 2 13 3 15 2 3 13 7 13 2 13 13 2
34 15 9 1 0 9 3 13 9 13 0 9 13 9 9 2 0 9 9 1 2 15 13 9 2 15 13 9 13 0 9 7 1 9 2
31 15 13 13 13 15 9 2 16 13 9 3 15 9 2 15 9 13 13 13 9 3 15 9 2 16 13 13 9 13 9 2
8 3 15 4 13 3 15 9 2
8 15 4 13 0 9 13 9 2
26 15 4 13 9 2 15 13 9 2 9 2 9 2 7 15 9 15 9 9 2 15 13 7 13 0 2
25 3 3 7 3 2 3 7 3 2 15 4 13 9 2 15 13 15 2 9 2 15 13 9 9 2
15 0 9 2 13 3 0 13 2 16 9 13 3 0 9 2
18 15 13 3 0 9 2 9 0 9 2 3 9 2 15 13 3 0 2
11 11 13 9 4 13 0 9 1 13 9 2
8 11 13 3 9 3 12 9 2
5 15 13 4 13 2
6 13 13 13 15 13 2
35 11 11 2 15 13 9 11 11 13 0 9 9 9 9 2 13 11 9 2 15 1 11 13 3 9 12 12 2 12 12 9 3 9 1 2
9 9 11 11 4 3 3 13 9 2
26 15 13 2 13 4 13 2 16 15 13 9 3 9 7 13 0 9 13 15 2 15 11 13 9 1 2
26 9 11 11 11 2 0 9 0 9 9 11 2 13 11 11 9 7 13 9 13 9 7 11 9 9 2
21 3 15 9 15 9 1 9 12 1 9 13 9 9 9 11 13 3 3 9 9 2
16 15 9 13 9 13 0 9 13 3 13 9 7 3 9 9 2
27 13 13 2 16 12 9 9 13 9 11 11 11 7 13 15 13 9 7 13 0 9 11 3 13 0 9 2
11 9 13 13 3 3 3 11 7 3 9 2
19 16 15 13 13 0 9 11 11 3 0 9 2 15 13 2 15 3 13 2
6 13 15 13 13 15 2
7 9 13 0 9 0 9 2
24 9 13 9 0 9 7 13 15 9 2 3 3 9 9 7 11 11 9 13 9 13 13 9 2
5 0 9 4 13 2
6 13 13 13 15 13 2
29 15 13 13 3 2 7 11 9 9 2 15 13 9 11 11 2 13 3 2 15 4 13 0 9 3 13 0 9 2
13 15 4 13 3 9 2 15 13 1 0 11 9 2
6 15 13 3 4 13 2
12 15 9 13 0 9 2 16 11 11 9 13 2
14 13 4 13 15 2 7 15 4 13 15 0 9 9 2
5 15 13 0 9 2
24 15 13 15 3 0 2 16 16 9 13 9 13 4 13 9 9 2 9 4 13 3 0 9 2
11 13 2 13 0 9 3 13 9 15 9 2
24 3 3 15 0 9 13 9 2 11 11 2 13 2 13 15 13 13 9 9 13 3 12 9 2
18 11 9 9 1 9 4 13 13 9 9 2 16 9 13 3 12 9 2
27 9 9 13 9 3 13 2 16 2 9 2 9 2 9 12 13 13 9 9 13 7 13 9 9 1 2 2
12 4 9 13 2 3 15 13 15 9 9 9 2
6 0 9 2 9 9 2
5 15 13 0 9 2
10 0 9 2 13 13 9 13 0 9 2
9 4 13 9 15 9 9 13 9 2
16 13 15 2 16 15 4 13 2 16 15 13 15 9 13 9 2
6 13 9 11 3 3 2
9 9 13 15 7 0 9 11 9 2
11 11 13 9 7 9 13 9 0 9 1 2
19 13 2 16 16 4 13 9 11 9 9 9 2 15 4 13 3 9 9 2
28 3 3 16 13 13 9 9 9 9 1 2 15 13 3 9 9 2 16 13 3 9 2 16 0 9 13 9 2
20 3 3 15 4 9 13 2 16 13 9 15 0 9 9 7 9 13 9 9 2
6 15 13 0 9 9 2
31 15 9 9 13 13 2 0 9 2 9 2 3 16 15 4 2 13 13 9 12 9 13 9 9 2 2 16 9 4 13 2
31 3 0 0 9 13 9 2 13 2 9 13 15 2 16 11 1 13 9 2 15 1 4 13 3 0 13 9 9 7 9 2
25 11 9 7 11 9 9 13 9 3 16 0 9 7 0 9 7 3 15 9 9 9 7 9 9 2
22 0 9 9 13 15 9 0 7 0 9 2 7 3 4 13 13 11 9 13 9 1 2
5 11 9 2 12 2
12 0 9 2 9 13 9 13 9 3 9 9 2
10 9 0 9 13 4 15 9 13 3 2
16 12 9 13 2 16 0 9 13 13 2 13 7 13 3 3 2
23 9 4 13 2 16 15 9 2 15 0 7 0 9 9 3 13 2 13 3 13 13 0 2
16 3 0 9 13 3 0 9 2 9 13 3 2 16 9 13 2
17 0 9 13 13 0 2 16 3 9 7 9 9 13 9 13 9 2
19 3 9 0 9 2 15 13 13 9 9 9 0 9 2 13 3 0 9 2
7 15 4 3 13 9 9 2
14 15 9 13 15 13 15 2 16 9 9 13 0 9 2
15 13 15 9 2 16 3 13 9 13 15 0 7 0 9 2
7 9 11 9 15 13 3 2
8 0 13 2 13 15 9 9 2
36 0 9 2 3 13 2 16 13 9 1 2 7 13 0 13 9 1 2 13 9 9 11 13 15 13 15 2 16 9 13 3 0 9 9 9 2
9 0 9 2 9 13 9 9 9 2
5 9 13 9 9 2
4 15 13 9 2
10 9 12 13 13 9 13 3 13 9 2
10 13 3 3 0 2 16 9 12 13 2
29 0 9 2 11 9 12 9 0 9 13 9 13 9 13 9 2 15 13 4 13 9 9 7 4 13 15 3 3 2
15 4 13 2 16 0 9 13 3 0 9 9 13 9 9 2
30 16 0 9 4 13 2 9 13 9 9 2 15 4 0 9 13 9 13 9 13 9 2 16 9 4 13 3 0 9 2
6 9 13 13 9 9 2
7 15 13 13 2 9 2 2
17 3 11 9 7 9 9 11 13 13 9 2 13 9 13 15 9 2
25 16 9 9 13 4 3 13 9 9 2 13 3 0 13 9 9 9 7 15 1 3 11 0 9 2
28 11 13 3 0 9 12 9 12 9 13 9 2 7 9 2 4 13 0 9 0 9 13 9 9 9 9 2 2
12 11 0 9 9 13 3 9 13 9 0 9 2
7 0 9 9 13 3 13 2
9 9 13 3 0 0 9 9 1 2
10 9 13 9 13 11 9 9 9 12 2
17 12 0 9 9 9 4 13 12 9 9 1 13 15 13 9 3 2
33 15 9 9 13 9 2 9 7 15 9 3 13 9 2 15 4 3 13 9 9 9 9 0 9 7 15 4 13 9 0 9 9 2
20 15 9 9 9 13 2 16 16 15 9 13 13 9 2 9 13 13 15 9 2
10 3 3 13 0 13 15 0 0 9 2
14 15 13 13 9 2 16 9 9 7 9 13 0 0 2
18 15 1 13 9 13 2 16 13 9 13 12 9 9 13 9 15 9 2
22 13 3 3 0 13 2 13 9 11 9 7 9 13 9 9 7 3 0 9 0 9 2
24 9 12 13 0 9 13 9 13 3 15 9 2 15 4 9 9 9 9 13 0 7 0 0 2
13 9 3 9 13 9 9 0 9 13 4 3 13 2
10 15 9 9 13 0 7 0 9 9 2
35 3 3 2 16 0 9 9 4 13 9 2 4 13 9 15 2 3 3 9 4 13 0 0 9 7 15 9 2 15 4 13 9 0 9 2
22 16 9 13 0 9 13 9 9 1 15 9 9 2 0 9 4 13 3 9 12 13 2
25 15 0 9 13 9 9 7 13 9 7 3 13 9 9 9 15 1 2 16 15 4 13 0 9 2
11 16 0 9 9 13 2 15 9 13 0 2
29 13 9 7 9 13 9 13 15 0 9 2 15 13 9 9 2 9 2 9 9 2 9 9 7 9 9 0 9 2
18 13 9 1 15 9 13 3 2 16 9 13 0 9 9 7 9 1 2
25 15 9 4 13 3 15 9 1 2 15 13 11 12 9 9 13 9 7 0 9 0 9 13 9 2
20 13 9 4 13 2 16 9 9 4 13 7 9 13 2 16 9 4 13 9 2
21 4 13 2 16 13 9 9 9 9 13 0 0 9 9 2 15 9 4 3 13 2
16 13 3 0 9 15 2 16 9 13 13 3 1 0 0 9 2
12 13 3 9 2 15 13 0 7 0 9 9 2
15 15 9 9 13 13 9 9 0 0 9 7 0 0 9 2
41 13 9 9 2 15 13 13 15 12 9 0 9 2 13 3 0 2 9 9 7 0 2 0 9 9 0 9 2 7 3 0 9 7 0 2 0 9 9 0 9 2
25 15 13 13 9 2 16 9 13 3 0 9 2 7 15 12 9 13 9 2 15 9 13 0 9 2
15 3 13 13 15 9 2 16 9 13 0 0 7 0 9 2
16 9 4 3 3 13 0 0 2 0 7 0 9 0 9 1 2
21 15 12 9 4 13 0 9 0 9 2 9 7 0 9 9 2 9 7 9 1 2
11 13 13 13 0 11 0 9 0 9 9 2
7 9 4 13 9 0 9 2
7 15 1 0 9 13 9 2
20 9 4 13 9 13 2 16 9 13 11 9 9 13 9 13 0 7 0 9 2
26 9 4 13 2 16 9 13 9 13 13 3 3 7 16 9 13 3 9 13 3 0 9 7 9 9 2
5 9 13 15 9 2
16 0 9 0 9 9 13 0 9 9 2 15 13 3 9 9 2
8 11 9 13 13 3 15 9 2
21 15 13 3 3 13 9 9 9 9 9 7 3 13 9 2 15 13 9 0 9 2
14 3 9 2 0 9 2 9 11 2 13 3 13 15 2
12 9 7 9 13 3 0 2 15 4 13 3 2
21 7 3 2 13 0 9 2 13 9 13 13 3 3 0 2 3 15 13 0 9 2
10 0 9 13 9 7 9 0 9 9 2
25 16 13 9 0 12 9 0 9 2 13 3 13 13 2 16 0 9 13 3 3 3 9 7 9 2
32 7 15 13 2 13 13 15 15 9 2 7 15 2 15 13 9 15 9 7 15 3 13 9 3 3 2 0 0 9 9 9 2
13 15 13 3 9 9 2 15 13 13 15 0 9 2
4 9 13 0 2
8 9 11 1 13 9 9 1 2
27 13 13 13 3 9 7 13 3 15 9 2 0 9 9 13 9 13 9 9 12 9 9 7 13 15 9 2
11 0 9 9 11 11 13 3 9 7 13 2
25 15 9 15 4 13 3 13 9 2 16 4 13 9 9 9 3 2 15 13 4 13 15 0 9 2
8 15 1 4 13 9 9 0 2
2 9 2
34 2 2 9 2 0 9 2 0 9 9 2 13 9 13 9 1 2 16 13 9 15 15 13 9 15 0 1 2 15 13 13 9 13 2
35 13 3 13 15 2 13 11 9 4 13 9 0 3 2 16 15 0 0 9 13 9 2 16 3 4 13 2 13 13 9 13 3 15 9 2
18 0 9 2 13 13 9 2 16 3 3 13 2 16 9 13 0 0 2
13 9 9 11 15 13 13 2 16 12 5 13 13 2
31 9 11 3 13 2 16 13 13 9 13 13 15 2 16 12 9 9 13 9 9 2 7 3 3 13 15 9 15 9 1 2
13 13 15 9 2 16 13 0 13 15 9 3 3 2
39 9 13 9 13 9 9 13 3 13 2 16 9 13 3 0 2 3 15 4 3 13 3 9 15 2 16 13 3 15 2 15 3 13 15 9 2 3 9 2
18 9 11 13 11 13 9 2 7 3 11 13 13 15 9 2 13 9 2
36 7 4 3 13 2 16 15 9 13 12 12 9 9 2 12 12 9 0 9 7 12 12 9 9 2 7 15 13 0 9 11 9 13 0 9 2
6 15 13 3 0 13 2
25 3 3 2 16 15 9 4 13 13 9 7 9 2 13 4 13 2 16 9 0 13 9 9 3 2
6 15 4 13 15 9 2
39 15 4 13 15 2 16 13 0 9 3 3 16 0 9 2 15 13 13 3 2 7 9 2 7 13 3 9 9 13 9 7 13 15 9 7 3 0 9 2
6 9 9 4 13 3 2
45 15 9 0 9 13 9 2 3 11 2 13 9 7 11 13 13 15 2 15 13 4 13 15 2 16 13 0 2 13 3 2 12 9 0 9 0 9 15 1 2 16 13 0 9 2
6 15 13 4 3 13 2
17 13 3 9 13 15 9 1 2 3 16 9 3 13 13 15 9 2
8 7 3 15 13 13 0 9 2
4 9 13 9 2
10 16 9 11 13 2 12 5 13 13 2
20 15 4 13 9 3 0 2 7 9 4 13 9 7 9 13 15 9 13 9 2
37 0 9 2 13 13 13 9 0 9 7 13 2 16 9 9 13 9 7 9 0 0 9 2 3 9 9 2 0 9 2 0 9 7 9 9 9 2
37 13 3 13 2 16 11 9 15 9 13 3 7 15 13 3 9 12 2 16 11 9 9 13 9 9 13 9 15 9 13 3 9 9 13 15 9 2
59 9 0 13 1 15 2 16 15 13 3 0 9 2 7 12 12 9 9 13 9 9 13 15 2 16 13 0 13 9 3 12 12 9 9 15 11 9 9 7 3 13 9 12 12 9 9 11 9 9 2 15 13 13 9 9 9 15 9 2
51 0 9 13 15 2 16 11 9 2 0 9 12 13 9 12 2 13 0 15 9 2 3 9 13 9 9 13 9 2 7 3 11 9 13 13 9 9 9 9 2 7 13 0 9 3 13 15 9 9 3 2
7 15 13 13 9 0 9 2
25 11 9 13 0 13 9 9 9 2 15 13 9 3 7 13 9 3 0 7 9 9 7 15 1 2
25 2 0 9 2 0 9 9 2 0 9 7 9 11 2 15 13 3 3 15 9 9 9 13 9 2
6 15 15 3 13 9 2
11 13 0 2 16 9 13 9 3 9 9 2
31 9 9 3 7 3 3 13 0 9 9 2 16 15 13 0 9 9 9 7 3 9 13 9 2 7 15 13 3 3 9 2
6 9 13 3 3 9 2
6 3 11 15 13 9 2
13 3 3 11 9 9 9 3 7 3 13 9 9 2
10 13 13 15 9 13 2 7 13 9 2
28 9 13 12 9 2 7 16 13 9 7 16 13 3 2 16 9 13 3 2 0 7 0 9 13 13 9 0 2
23 0 9 2 7 3 0 9 2 9 4 13 9 9 2 7 3 15 15 0 9 4 13 2
27 16 13 9 9 9 7 15 9 13 3 9 9 7 9 2 13 9 13 3 2 3 15 4 13 9 9 2
22 15 1 13 9 11 9 3 0 2 16 15 13 0 0 9 2 15 15 9 13 9 2
10 13 0 2 16 11 3 13 15 9 2
13 13 2 16 15 12 13 13 9 13 3 0 9 2
43 13 15 2 16 15 13 3 15 0 2 7 11 9 7 3 9 13 3 13 0 9 2 15 13 0 9 2 13 15 15 9 2 15 13 11 15 9 2 13 3 13 11 2
12 15 1 13 9 0 0 2 16 13 0 9 2
30 3 15 13 4 13 3 3 9 15 2 15 9 13 15 9 2 16 2 9 3 2 9 13 13 9 3 15 9 9 2
26 15 4 13 15 15 11 0 9 9 2 15 2 0 7 0 2 9 13 3 3 0 7 0 9 9 2
29 15 13 0 9 2 7 0 9 0 7 0 9 1 13 15 2 16 0 9 13 9 9 0 7 0 9 13 13 2
18 9 13 15 2 4 13 9 3 2 16 3 0 9 13 7 0 13 2
32 0 9 15 2 16 13 15 9 3 13 2 16 9 7 9 9 4 13 15 2 16 9 13 3 3 0 13 0 9 0 9 2
11 9 7 9 1 4 3 3 13 0 9 2
28 15 1 13 0 2 16 13 3 9 13 9 2 13 15 3 7 13 3 2 15 13 0 9 2 7 13 9 2
9 15 1 13 3 3 9 11 9 2
6 9 4 3 13 0 2
15 13 13 3 13 9 7 9 2 7 15 4 13 9 9 2
22 4 3 13 13 9 9 2 15 13 3 3 9 13 9 7 15 9 4 13 9 9 2
13 9 4 13 1 9 2 7 15 4 13 0 9 2
36 9 2 3 16 11 9 2 9 2 7 11 9 9 9 2 13 0 2 16 9 13 3 2 16 13 15 3 7 16 9 13 9 0 9 9 2
17 0 9 2 13 9 9 11 2 15 13 13 15 9 3 7 3 2
23 9 15 9 13 0 9 2 13 2 16 11 9 13 0 9 2 15 9 4 13 3 13 2
35 13 2 16 9 7 9 13 2 16 9 4 13 3 3 7 16 15 9 4 15 9 13 13 3 9 9 2 16 15 13 13 9 15 9 2
23 15 9 13 13 9 3 9 2 15 13 15 9 2 7 13 13 0 9 13 15 0 9 2
13 9 13 4 13 3 15 9 2 15 9 16 15 2
8 9 13 3 3 15 9 0 2
8 15 13 4 15 9 13 9 2
9 15 13 0 0 9 13 15 15 2
28 13 13 2 3 9 9 4 3 13 9 2 7 15 4 13 13 9 9 7 15 4 13 15 9 9 13 9 2
10 15 4 13 15 9 7 13 15 9 2
11 13 11 9 0 9 12 13 9 3 13 2
21 13 2 16 15 15 4 13 0 9 2 7 13 15 0 9 15 9 9 0 9 2
14 0 9 2 13 3 9 2 15 13 15 13 9 9 2
26 3 13 9 1 15 4 3 13 13 15 9 9 9 2 15 13 9 2 3 0 9 9 13 13 11 2
17 4 15 13 13 3 2 7 9 9 9 9 4 13 13 15 3 2
16 3 4 13 15 9 7 9 15 9 2 15 13 13 13 3 2
3 9 1 2
27 2 2 9 2 0 9 2 11 7 11 13 12 9 0 9 9 2 15 13 9 9 15 9 13 12 9 2
10 15 9 0 9 13 0 11 11 9 2
10 0 9 4 13 0 0 9 11 1 2
11 9 0 9 13 9 15 0 9 13 3 2
10 15 13 0 9 2 15 13 3 0 2
16 0 9 13 9 0 9 2 16 9 7 9 13 3 0 9 2
8 9 13 13 9 2 9 13 2
31 3 3 9 9 13 9 12 13 9 2 7 3 2 9 13 9 1 2 4 3 13 0 0 9 2 13 0 7 3 0 2
16 13 2 16 9 13 9 9 3 3 2 3 3 9 0 9 2
15 9 9 2 15 3 0 9 4 13 2 13 13 3 0 2
12 0 9 9 9 12 13 0 7 3 0 9 2
17 13 0 2 16 0 9 0 9 13 9 7 9 7 13 3 9 2
10 3 15 13 0 9 15 3 13 9 2
10 3 9 1 13 2 9 13 13 0 2
21 15 9 1 11 4 13 0 9 13 9 13 9 2 15 1 9 13 4 13 3 2
17 3 11 9 9 13 3 0 9 13 3 0 1 9 13 0 9 2
17 0 9 9 9 9 13 13 15 9 2 7 9 15 13 9 9 2
26 0 9 9 2 13 9 3 3 2 16 0 9 13 0 9 0 9 2 15 9 15 9 13 3 13 2
12 16 11 13 9 13 9 2 11 4 13 0 2
10 13 0 0 2 16 15 13 0 9 2
16 13 9 9 7 15 9 9 7 13 2 16 9 13 3 9 2
17 13 13 3 9 11 11 15 9 7 9 13 9 2 15 3 13 2
38 0 9 2 0 9 2 0 9 9 2 9 2 9 7 3 13 9 13 15 3 13 0 0 2 0 9 0 7 0 9 2 15 9 4 13 9 9 2
29 9 9 13 3 3 15 2 0 3 3 0 2 16 3 0 9 3 9 7 3 13 9 9 7 9 13 9 9 2
13 13 13 3 2 15 13 7 13 7 3 13 9 2
24 13 9 13 9 2 3 13 15 9 2 15 4 3 13 9 2 15 13 0 16 3 13 9 2
24 3 3 13 9 13 9 2 15 13 7 15 13 1 9 7 9 9 7 9 9 9 13 9 2
35 16 13 3 3 9 2 4 13 2 16 15 13 15 9 7 3 13 9 13 0 9 2 15 13 7 0 7 0 9 7 15 1 0 9 2
7 15 9 13 3 0 13 2
27 15 1 9 13 0 13 9 13 3 2 16 15 13 9 7 15 9 9 9 0 9 7 13 15 3 9 2
20 9 4 13 2 16 15 0 9 13 0 9 2 15 13 3 3 13 0 9 2
67 0 9 9 13 9 9 13 0 0 7 9 2 3 0 9 2 15 13 0 7 9 0 9 7 15 13 3 0 9 15 9 9 13 9 9 2 15 9 13 0 2 16 13 15 13 0 9 9 7 9 13 9 2 15 13 3 0 0 9 9 7 9 9 0 9 1 2
20 3 9 9 13 13 15 9 9 2 9 7 9 13 9 7 9 9 13 9 2
21 9 13 9 9 3 2 16 3 13 12 9 1 4 13 3 12 0 9 13 9 2
11 15 13 15 0 9 2 15 13 9 13 2
35 15 1 11 9 2 15 13 13 9 3 13 9 2 13 0 9 7 9 0 9 7 9 1 2 15 13 2 16 0 9 13 9 15 9 2
36 15 9 0 9 9 4 13 9 13 9 2 15 13 9 0 9 13 15 16 0 9 13 9 9 2 0 9 9 13 12 0 9 9 13 9 2
20 11 9 13 15 9 2 16 15 16 0 9 13 9 9 13 0 12 9 9 2
20 15 15 9 13 9 2 15 13 3 0 2 7 15 9 3 3 3 13 15 2
19 11 9 13 3 15 9 2 16 15 0 9 9 13 0 9 7 13 9 2
31 9 2 15 13 15 9 9 9 2 15 9 4 13 2 4 13 3 3 13 9 2 15 13 3 9 0 0 9 7 9 2
18 15 9 9 13 2 16 0 9 4 13 0 2 0 9 13 7 13 2
26 3 13 13 7 13 15 2 3 0 9 4 9 13 13 0 15 16 0 9 2 15 13 9 4 13 2
20 16 9 13 12 0 0 7 0 9 13 9 2 13 9 13 9 7 13 15 2
36 13 3 0 13 15 13 9 15 1 2 16 15 13 13 9 15 16 0 9 2 16 4 13 2 16 0 7 0 9 2 15 3 13 9 9 2
17 0 9 2 11 7 11 0 9 9 13 3 11 9 9 13 9 2
31 13 13 3 3 9 11 9 2 16 9 13 11 7 11 9 0 9 7 13 13 3 9 0 9 13 0 9 11 9 9 2
12 15 13 0 3 11 7 3 15 9 7 9 2
7 9 13 11 9 11 9 2
40 9 13 15 9 2 13 15 4 13 15 3 2 16 3 0 9 13 13 0 9 2 15 13 15 2 16 15 9 13 3 7 1 9 7 9 11 13 9 9 2
34 3 13 0 9 2 15 15 9 13 13 9 15 15 3 3 13 0 9 1 7 15 15 13 13 3 13 3 2 16 13 9 13 9 2
32 0 9 0 11 9 13 3 15 9 2 3 16 15 13 13 3 13 15 1 2 13 0 9 7 9 13 3 3 15 0 9 2
14 0 9 3 13 2 7 15 0 9 13 3 13 13 2
22 15 4 13 15 9 2 16 13 13 0 9 15 2 16 11 9 13 3 3 0 9 2
3 15 13 2
7 13 11 13 9 3 13 2
9 9 7 9 9 9 4 3 13 2
16 11 13 4 3 13 3 3 0 9 9 9 13 9 3 1 2
21 15 0 13 3 2 3 9 11 9 1 2 13 0 9 7 9 1 11 9 9 2
10 15 13 15 9 7 11 7 0 9 2
12 0 9 4 3 13 3 3 13 0 9 9 2
44 2 0 9 2 0 9 9 2 0 9 2 13 9 13 9 0 9 9 13 0 9 2 7 13 15 3 15 9 2 3 15 15 2 15 9 7 9 4 13 9 11 11 9 2
16 9 13 0 13 9 13 9 2 7 15 4 13 3 15 9 2
40 0 9 9 2 13 13 15 2 15 15 9 4 3 13 2 13 3 2 16 15 15 9 3 13 9 3 0 9 2 16 11 4 13 3 13 9 3 9 9 2
34 16 13 9 0 9 9 2 13 3 2 16 3 4 13 11 2 11 2 11 7 11 2 15 13 3 13 9 2 16 3 4 3 13 2
14 15 1 11 2 0 11 7 11 9 13 9 1 0 2
25 9 13 3 9 9 2 7 3 3 3 9 2 16 9 2 0 9 2 9 9 13 9 9 9 2
18 3 3 11 7 11 0 0 0 9 13 9 9 13 3 9 9 9 2
26 15 9 13 3 15 9 2 16 11 4 13 13 0 9 3 0 13 9 13 9 9 9 13 15 9 2
20 9 13 4 13 9 0 9 9 9 9 0 9 13 11 9 9 9 13 9 2
20 15 1 9 4 13 12 11 9 9 2 11 2 11 2 11 2 11 7 11 2
7 15 9 13 4 13 9 2
19 4 13 2 16 9 9 13 9 9 2 7 3 9 4 13 7 13 9 2
20 9 13 3 9 13 9 2 16 4 13 15 9 13 0 7 0 11 9 9 2
32 9 13 0 7 0 9 13 9 2 15 13 9 9 7 15 13 9 7 0 9 11 7 15 13 9 13 9 2 9 7 11 2
19 2 2 9 2 13 15 9 1 2 15 13 11 9 9 11 9 9 13 2
22 9 13 9 0 9 2 16 15 13 9 13 9 2 15 13 9 11 0 9 11 9 2
36 15 13 3 0 9 2 3 15 2 15 13 2 16 4 13 2 0 9 9 2 13 9 2 15 1 13 9 2 0 0 9 9 7 9 9 2
34 7 9 2 15 13 0 9 13 9 7 9 9 9 9 13 3 16 2 0 9 2 9 2 9 13 2 16 9 13 3 12 9 2 2
36 0 13 3 9 2 15 13 2 16 1 0 9 9 13 0 9 13 9 2 7 15 9 13 13 15 9 2 15 13 13 11 9 2 13 9 2
12 15 9 13 2 15 3 9 4 15 9 13 2
15 9 13 3 13 11 9 2 15 13 3 13 3 0 0 2
10 3 9 11 9 13 3 0 9 9 2
26 15 13 11 9 1 13 0 9 2 15 9 4 13 9 2 7 15 13 13 9 7 0 9 9 9 2
7 13 4 13 0 0 9 2
15 0 9 2 9 9 7 9 13 9 9 4 13 3 0 2
25 13 13 3 3 0 9 2 3 2 3 13 9 9 4 13 3 9 7 9 9 4 13 9 9 2
12 3 13 0 0 7 0 13 13 0 9 9 2
9 15 13 15 7 9 11 9 9 2
13 3 2 0 3 2 9 13 3 15 15 13 9 2
11 3 13 3 9 13 9 3 3 9 9 2
25 15 13 13 9 2 15 13 9 9 0 2 0 9 2 7 15 13 9 2 15 13 9 0 9 2
15 15 15 4 13 7 3 13 3 2 16 13 9 3 9 2
14 4 13 15 3 9 2 7 15 9 4 13 9 11 2
9 15 1 13 0 13 9 3 9 2
1 9
29 3 15 13 13 9 9 15 9 7 13 0 13 4 13 15 2 16 0 9 9 9 13 3 13 9 9 15 9 2
43 3 3 15 13 2 16 9 9 13 15 9 2 16 15 13 9 12 9 9 2 7 16 9 13 3 0 9 2 13 13 9 9 13 3 3 0 7 9 1 13 9 13 2
7 13 13 9 9 0 9 2
53 4 15 7 15 11 9 13 9 13 9 9 0 15 2 16 16 15 13 15 13 0 9 2 9 13 13 9 11 7 3 11 9 9 13 9 13 16 15 9 13 1 9 7 9 2 7 9 1 3 13 11 9 2
4 9 13 15 13
12 13 0 9 1 9 2 9 13 3 0 13 2
14 9 13 0 7 0 9 2 13 9 3 13 0 9 2
13 9 13 15 2 15 3 13 15 15 9 15 13 2
18 15 13 9 13 9 9 9 13 2 13 9 7 9 13 9 3 15 2
14 9 13 7 13 9 7 9 13 9 0 9 0 9 2
24 15 13 3 9 2 9 13 4 3 3 13 2 9 13 4 3 3 13 13 0 9 13 9 2
28 13 15 4 13 15 7 13 15 15 13 2 15 13 3 9 13 15 15 2 13 9 2 9 0 7 0 9 2
31 13 15 3 13 3 16 13 3 3 2 16 15 13 3 9 15 13 9 2 9 15 4 3 13 15 9 7 13 15 3 2
13 3 15 4 13 9 2 3 15 13 3 3 13 2
15 3 15 3 13 2 13 9 2 16 3 3 15 15 13 2
9 15 15 3 13 2 9 13 9 2
14 13 13 3 3 13 13 2 13 13 3 3 9 13 2
31 3 13 2 16 15 3 13 3 2 16 15 3 13 9 15 9 2 15 13 15 3 0 9 7 13 15 15 0 9 3 2
19 15 13 3 9 13 2 13 15 15 3 4 4 13 2 13 3 15 15 2
19 13 15 13 13 2 13 7 13 9 2 15 3 16 15 9 4 15 13 2
7 13 3 4 13 15 9 2
8 13 15 3 9 2 0 0 2
11 13 3 13 15 3 2 13 13 3 13 2
13 7 13 3 13 15 13 2 13 15 13 15 9 2
13 3 9 13 13 15 2 13 3 15 3 0 9 2
14 15 13 3 0 9 2 15 13 3 3 13 13 3 2
19 7 3 15 13 2 13 2 13 15 2 3 15 2 13 9 3 9 9 2
12 15 4 13 0 15 2 15 3 0 3 13 2
17 13 15 3 9 2 3 9 13 9 2 3 4 15 9 13 9 2
15 13 13 13 9 13 3 2 13 3 3 9 7 13 9 2
30 9 9 13 13 2 16 3 16 15 4 13 3 15 9 13 2 15 9 13 13 15 0 9 3 15 2 15 3 13 2
18 13 9 2 7 13 3 13 9 2 15 4 3 13 2 9 4 13 2
23 4 13 2 16 15 4 13 0 9 13 9 2 3 15 13 2 13 13 0 16 9 3 2
14 7 3 15 13 3 15 2 13 16 13 3 9 13 2
6 13 13 15 3 13 2
10 16 4 13 2 15 4 13 3 3 2
19 7 13 3 3 0 13 2 13 4 3 13 15 2 13 4 15 16 13 2
18 9 13 13 9 3 2 9 13 12 9 9 13 9 13 3 15 0 2
9 3 15 13 3 0 2 0 9 2
19 9 9 13 0 0 2 9 13 13 9 2 3 13 0 2 3 0 0 2
6 3 16 15 13 13 2
7 3 15 4 13 2 9 2
7 0 2 0 9 13 9 2
18 13 13 9 15 1 2 13 13 7 13 9 2 7 13 3 3 9 2
5 9 13 7 13 2
15 15 13 0 9 2 9 15 1 7 9 13 3 0 9 2
8 13 13 2 15 13 3 0 2
11 3 15 13 2 13 9 7 9 15 9 2
8 13 13 2 15 15 9 13 2
9 2 15 13 2 16 15 13 3 2
15 3 13 9 2 13 3 9 2 13 15 3 3 13 9 2
24 0 9 2 3 15 13 3 2 15 13 15 3 16 9 2 3 15 3 13 2 13 15 13 2
9 13 3 13 3 2 13 15 3 2
2 9 9
14 0 2 0 9 13 0 9 13 9 3 15 9 1 2
15 9 15 13 0 0 2 0 9 2 15 9 13 0 3 2
21 9 13 0 9 1 1 9 2 15 13 3 9 2 15 3 0 9 13 2 0 2
19 15 2 15 13 9 7 9 9 2 9 13 7 9 13 13 9 9 1 2
15 9 13 13 9 2 9 13 9 7 15 13 9 3 13 2
21 9 13 0 0 9 3 2 9 3 13 9 3 3 9 3 13 7 13 15 9 2
19 9 13 9 1 2 13 9 9 7 13 9 2 13 3 3 7 13 9 2
16 15 13 0 9 13 9 9 9 2 16 15 9 13 9 9 2
13 9 13 9 2 13 9 2 7 13 9 0 9 2
16 3 0 13 9 2 9 3 13 3 7 3 0 0 9 3 2
25 9 13 0 9 0 9 2 7 3 15 13 13 9 7 9 2 15 4 3 13 9 9 1 9 2
22 15 13 2 13 3 2 3 13 15 3 4 13 2 7 15 3 13 9 2 0 9 2
12 9 13 9 2 11 7 11 2 13 9 13 2
18 11 13 13 9 2 7 13 9 9 2 15 13 9 7 13 9 3 2
19 9 1 15 9 13 2 9 13 2 13 9 2 3 9 15 13 3 13 2
10 13 3 9 2 15 13 3 13 15 2
21 9 13 9 2 15 13 0 0 9 2 15 13 9 15 15 13 3 3 13 13 2
14 11 7 11 13 3 3 2 9 2 15 13 9 9 2
14 9 13 3 0 2 16 0 9 13 15 15 13 15 2
14 15 13 0 9 2 15 9 7 15 9 13 15 9 2
17 15 4 13 15 2 16 9 13 13 2 16 15 9 4 3 13 2
20 15 13 0 9 2 15 4 13 7 15 3 0 9 13 13 15 2 16 13 2
12 3 0 9 13 0 9 2 3 0 0 9 2
8 13 3 0 13 15 13 15 2
16 9 13 9 2 16 9 13 3 3 0 2 16 15 13 9 2
19 15 13 13 15 13 13 2 15 4 3 13 15 3 7 13 2 13 9 2
13 9 2 15 9 9 13 2 11 7 11 13 13 2
11 15 13 0 9 2 0 9 7 13 15 2
11 11 13 9 13 9 9 7 13 15 9 2
16 15 9 11 13 9 2 15 9 13 13 3 16 9 4 13 2
26 9 7 9 1 13 9 2 15 9 13 4 13 2 15 9 13 4 13 2 16 15 4 13 9 1 2
14 3 15 15 15 4 13 2 3 3 15 15 3 13 2
10 9 9 13 13 7 13 9 3 3 2
10 3 15 13 16 15 13 3 4 13 2
11 11 7 11 13 0 9 7 13 9 1 2
19 9 13 3 3 2 9 13 3 3 2 15 13 13 16 15 4 3 13 2
16 11 7 11 9 13 13 3 9 2 7 9 9 13 3 9 2
7 15 13 3 3 13 3 2
16 9 13 13 3 3 0 13 2 3 9 13 15 13 0 9 2
6 3 15 13 13 3 2
16 11 7 11 9 13 13 0 15 13 2 3 3 15 13 13 2
26 0 7 0 13 9 13 2 16 15 9 4 13 13 3 3 2 16 0 9 2 15 13 13 3 3 2
10 0 7 0 13 9 2 13 15 9 2
1 9
26 0 9 9 13 9 9 13 12 9 9 7 9 0 11 2 13 9 2 15 2 15 15 13 9 13 2
23 13 3 3 0 2 16 9 4 13 9 3 2 13 9 9 9 13 2 16 3 15 13 2
20 9 9 13 9 9 1 0 9 7 9 2 9 13 0 13 9 7 15 9 2
11 3 15 9 13 2 15 15 4 13 15 2
11 9 13 9 2 9 0 9 13 3 9 2
14 15 13 9 2 13 15 13 15 16 4 13 9 9 2
18 7 15 13 3 15 9 2 15 15 13 13 13 2 13 13 13 13 2
8 9 13 9 2 16 13 0 2
15 9 13 9 3 2 16 13 0 13 2 4 15 13 15 2
12 15 13 4 13 15 9 2 15 13 15 9 2
25 9 13 0 9 13 15 1 7 9 13 3 0 2 16 15 13 9 0 9 9 3 16 13 15 2
7 15 9 15 4 13 3 2
20 13 9 2 13 9 0 9 3 13 0 9 2 9 9 13 2 9 9 9 2
22 9 15 13 2 16 4 13 9 9 2 7 9 13 3 0 7 0 2 13 15 13 2
17 15 9 13 7 13 3 0 2 16 9 9 9 13 15 9 3 2
21 13 15 4 13 15 9 9 15 2 15 15 13 13 1 9 2 7 15 13 3 2
20 9 13 13 3 16 15 3 13 7 3 9 9 13 9 13 13 15 13 9 2
11 9 13 9 9 2 13 9 9 1 9 2
12 15 9 15 4 13 13 1 9 7 13 9 2
7 15 13 8 7 9 9 2
1 9
7 3 13 9 1 9 9 2
13 3 13 0 9 9 13 9 1 7 13 0 9 2
11 15 13 13 2 0 9 2 15 13 9 2
20 13 15 9 13 1 15 2 13 15 9 9 2 9 9 2 13 9 9 1 2
6 13 15 13 3 15 2
6 13 15 13 3 15 2
11 15 13 0 9 2 0 9 13 13 9 2
10 15 13 9 9 7 13 3 9 9 2
9 15 9 13 16 9 9 13 9 2
14 7 15 13 3 2 3 3 15 9 1 7 15 1 2
12 13 3 9 2 9 7 9 1 2 3 15 2
15 15 13 13 15 9 2 13 16 13 9 1 9 9 9 2
12 3 13 9 13 3 3 3 2 13 15 9 2
4 15 13 15 2
9 13 15 9 9 1 13 9 1 2
11 15 13 2 13 15 9 7 13 9 9 2
11 9 13 0 9 15 7 15 13 3 9 2
18 9 13 9 13 9 1 7 9 13 9 9 13 3 3 9 9 0 2
2 0 9
13 13 3 0 9 11 9 9 0 9 0 9 0 2
11 4 13 9 13 9 2 9 7 0 9 2
14 15 13 9 16 12 9 0 9 2 9 9 9 13 2
13 9 13 15 11 9 9 2 9 0 2 3 0 2
4 3 13 3 2
7 3 13 13 9 13 9 2
10 9 13 9 2 13 15 9 13 9 2
12 9 13 0 1 9 7 0 9 9 9 1 2
6 0 9 13 13 9 2
11 9 13 9 7 9 9 3 0 9 1 2
16 9 13 0 1 7 9 9 13 9 13 0 2 15 15 13 2
1 9
8 13 3 9 0 9 9 13 2
13 9 4 13 9 2 9 9 7 9 13 9 9 2
9 15 13 0 7 0 16 9 9 2
14 15 9 13 9 3 3 2 16 15 13 3 9 1 2
18 9 13 9 3 3 7 13 9 3 0 2 16 4 4 13 9 13 2
10 15 13 4 3 13 2 3 13 9 2
9 13 13 2 13 4 15 3 13 2
9 15 9 13 13 3 16 3 13 2
13 9 2 9 9 13 0 9 13 0 9 13 9 2
28 15 13 2 3 3 15 13 2 15 9 16 3 13 11 9 9 9 1 7 3 13 3 3 16 9 9 15 2
14 9 13 15 3 3 3 7 13 9 9 13 9 9 2
11 15 13 3 3 0 0 2 3 15 9 2
22 15 9 13 3 9 0 0 2 13 9 2 13 9 2 7 3 0 9 9 9 0 2
12 9 9 13 7 3 3 13 13 0 16 9 2
20 13 9 2 13 15 9 3 0 16 9 2 13 3 4 13 2 16 15 13 2
17 7 0 9 13 13 2 9 13 9 9 2 16 9 3 13 13 2
8 9 9 13 9 13 9 3 2
19 13 13 13 15 9 2 16 9 13 3 15 3 0 2 15 13 15 0 2
14 13 9 9 13 9 1 2 13 4 4 13 9 3 2
26 7 15 13 4 4 13 2 16 15 13 3 13 9 15 2 13 3 9 1 9 7 13 15 3 13 2
10 13 9 9 7 13 9 13 9 9 2
10 9 3 4 13 13 9 9 16 9 2
20 13 9 0 9 2 9 7 9 2 13 9 9 7 12 9 1 13 9 9 2
7 15 9 13 13 2 13 2
9 9 13 0 0 0 9 9 1 2
8 0 9 2 15 9 13 0 2
16 3 0 13 15 9 1 9 7 3 3 13 2 3 4 13 2
1 9
9 13 9 2 13 9 7 12 9 2
8 4 13 2 16 9 1 9 2
8 3 2 0 9 2 15 3 2
6 15 9 13 9 3 2
4 9 13 9 2
9 3 2 13 9 2 13 9 9 2
9 13 3 2 11 2 11 2 11 2
15 13 9 7 9 2 13 9 7 13 16 9 13 3 9 2
18 13 9 3 0 9 1 0 9 1 7 13 9 2 15 13 3 9 2
9 13 9 1 13 9 7 13 9 2
17 16 13 3 2 13 3 3 2 9 1 13 15 9 7 9 9 2
1 9
13 15 4 3 13 9 2 16 9 13 9 1 9 2
10 4 13 3 9 9 9 2 13 13 2
14 13 15 15 9 2 16 9 13 9 1 0 9 3 2
10 15 9 9 13 9 3 16 9 9 2
1 9
17 13 9 9 13 0 9 7 13 13 13 9 13 9 7 9 9 2
7 15 15 4 13 2 13 2
5 15 13 9 9 2
20 13 3 0 9 9 9 9 9 1 13 2 9 13 1 9 13 9 13 9 2
14 11 13 3 13 15 2 13 9 9 9 7 13 3 2
10 15 13 13 15 0 2 9 13 15 2
6 15 13 15 9 9 2
19 16 4 13 13 13 15 15 9 1 2 15 15 9 13 2 4 13 13 2
12 15 13 13 15 9 2 15 13 0 15 9 2
12 3 2 15 9 13 3 1 11 7 15 9 2
13 15 4 13 9 9 7 15 13 15 1 16 9 2
17 13 15 2 16 13 11 2 13 3 2 16 13 15 1 15 1 2
17 3 3 4 4 13 12 9 1 2 16 15 4 13 9 0 9 2
17 4 13 15 3 2 13 3 3 16 15 15 2 13 4 13 15 2
7 11 13 7 13 3 9 2
15 2 13 15 3 13 2 7 2 2 2 15 13 3 3 2
8 13 15 3 16 13 15 9 2
13 13 15 4 13 2 3 4 2 16 15 13 13 2
12 11 13 9 9 2 13 9 7 13 15 3 2
9 15 13 4 13 2 13 15 13 2
11 13 9 7 13 9 3 3 2 13 13 2
4 9 0 16 9
5 9 13 13 13 2
8 9 1 13 9 13 0 9 2
4 15 13 3 2
12 13 15 2 13 15 9 2 13 9 9 1 2
12 13 13 13 9 9 9 3 0 9 13 15 2
9 13 3 3 2 16 9 13 0 2
8 13 13 9 1 2 13 15 2
7 13 3 2 13 13 13 2
8 13 9 9 1 12 0 9 2
9 9 0 9 13 15 1 3 13 2
11 15 13 4 13 2 15 13 4 13 9 2
10 9 13 9 2 0 9 7 0 9 2
18 3 13 15 2 13 3 0 0 9 2 15 2 15 1 15 13 13 2
1 11
5 9 13 9 1 2
18 15 13 13 3 9 2 13 15 9 0 9 7 12 7 12 9 9 2
14 9 15 13 12 9 9 9 2 15 9 7 9 9 2
10 9 13 15 9 9 2 9 15 9 2
25 3 15 13 9 2 7 13 9 7 9 2 15 2 15 15 4 9 1 13 2 2 15 13 0 2
20 9 13 13 9 13 9 2 15 13 3 13 2 3 15 4 3 13 3 0 2
6 9 13 3 13 9 2
15 3 2 15 1 15 13 9 2 13 15 9 7 9 1 2
21 16 15 3 13 9 2 9 13 3 3 9 9 9 2 7 15 9 13 3 9 2
14 15 9 13 9 15 15 9 2 15 15 4 9 13 2
13 9 13 7 13 3 0 2 3 9 13 15 13 2
7 3 9 13 9 9 9 2
19 3 9 13 0 2 3 0 2 16 9 4 13 15 0 9 3 3 9 2
8 9 13 13 1 9 0 9 2
15 13 3 0 2 9 13 3 3 2 16 9 9 13 0 2
6 9 13 9 7 13 2
12 3 15 13 13 2 16 15 9 13 15 9 2
11 3 15 13 2 16 13 15 9 15 1 2
12 3 16 13 2 13 3 13 3 2 9 13 2
6 3 15 4 13 13 2
10 9 13 13 15 15 2 13 13 9 2
14 9 4 13 15 3 2 3 15 4 13 7 13 3 2
9 3 3 3 2 16 15 13 0 2
1 11
14 11 13 9 2 13 9 9 7 13 0 2 0 9 2
10 9 13 9 2 7 3 15 13 13 2
6 13 0 2 13 0 2
6 9 2 15 3 13 2
15 0 9 13 13 13 2 13 11 13 13 15 12 9 1 2
17 3 9 9 13 13 9 0 9 2 15 13 15 3 13 9 9 2
13 13 15 15 13 13 9 2 7 9 13 3 13 2
12 11 13 3 13 15 13 9 2 9 7 9 2
11 15 13 0 9 16 11 13 15 9 1 2
16 15 13 9 0 9 2 9 9 9 1 2 13 9 0 9 2
9 15 2 15 11 4 9 9 13 2
13 9 13 11 3 2 13 3 9 1 7 13 13 2
13 3 13 11 9 2 15 13 9 2 15 13 15 2
12 7 11 4 13 13 2 13 9 13 13 15 2
8 3 3 11 9 13 3 3 2
12 3 15 13 2 3 9 7 11 13 3 3 2
11 9 4 13 3 13 15 7 13 15 0 2
12 3 9 4 13 2 13 11 3 3 13 9 2
18 15 13 0 9 2 15 11 13 9 13 15 3 3 11 9 9 9 2
15 15 13 13 15 3 2 3 13 9 2 15 15 3 13 2
23 11 13 13 9 0 9 15 2 16 12 9 1 11 9 9 13 9 2 11 13 15 3 2
12 13 15 13 2 13 13 9 1 2 13 15 2
1 9
10 15 13 9 0 9 7 13 0 9 2
14 9 2 3 15 3 13 9 9 9 13 0 16 13 2
7 13 15 3 3 13 0 2
35 1 3 3 0 9 2 16 15 9 9 13 15 9 9 2 3 15 2 15 15 4 13 9 3 9 2 7 13 15 3 9 0 9 9 2
9 3 15 13 0 2 3 13 9 2
12 15 13 15 15 9 2 15 15 4 4 13 2
16 9 4 4 13 9 12 7 13 11 0 9 0 9 13 9 2
21 7 9 13 2 3 13 2 9 2 13 3 13 3 13 12 0 9 1 9 9 2
15 9 9 13 3 13 15 9 2 9 9 7 9 0 9 2
15 13 3 13 2 15 13 0 9 2 3 15 13 9 13 2
7 9 9 13 13 15 3 2
20 15 1 15 13 9 15 9 9 9 2 13 9 9 7 13 13 9 9 1 2
5 13 2 13 15 2
4 9 12 2 12
7 9 13 0 9 2 5 2
7 9 9 13 13 3 0 2
17 3 13 13 9 7 3 9 2 7 3 2 15 13 3 15 9 2
2 3 2
6 11 13 15 7 13 2
10 16 9 13 13 2 13 13 13 3 2
10 9 13 13 13 9 2 4 13 3 2
8 4 13 9 9 13 0 9 2
5 4 13 0 9 2
12 4 13 0 9 3 15 13 3 3 1 9 2
15 4 13 13 9 3 3 16 3 2 12 2 12 2 12 2
25 16 3 13 9 2 15 4 13 3 7 3 3 3 2 16 15 13 7 13 9 9 2 7 13 2
19 9 9 13 12 9 7 9 12 9 2 15 15 11 4 3 3 15 13 2
11 9 4 13 0 2 7 15 13 3 0 2
22 3 15 13 3 7 3 7 12 9 15 2 11 13 3 7 13 3 2 13 0 9 2
10 9 13 0 2 9 1 4 13 9 2
6 13 3 12 2 3 2
11 9 13 0 2 7 13 2 9 2 9 2
8 0 9 15 9 2 3 3 2
13 15 9 15 13 2 9 2 15 4 3 13 3 2
8 9 9 13 9 2 3 0 2
22 9 9 13 12 9 2 9 0 9 2 12 9 0 9 9 2 12 9 13 9 9 2
5 4 13 15 13 2
8 9 9 4 13 3 0 9 2
12 11 13 3 13 13 3 15 0 9 15 13 2
11 9 15 13 3 2 16 3 15 3 13 2
3 13 9 2
13 15 15 3 4 9 13 2 3 2 0 0 9 2
6 13 3 2 13 3 2
6 13 15 3 0 9 2
7 9 4 13 9 7 9 2
2 15 2
16 0 9 15 13 3 15 9 7 13 2 16 9 4 13 9 2
15 15 9 11 13 9 3 9 9 7 13 3 9 15 9 2
12 9 9 7 9 13 9 13 13 2 3 9 2
24 3 9 9 1 7 0 9 13 4 13 9 7 9 7 9 7 9 7 0 0 9 13 9 2
13 3 2 0 9 13 3 0 2 13 13 3 9 2
6 13 3 0 15 13 2
20 3 0 9 9 1 2 7 15 13 3 2 9 13 3 9 0 0 9 3 2
11 11 13 9 9 2 3 2 13 13 15 2
12 0 13 2 16 13 9 2 13 9 13 3 2
10 9 13 3 2 9 2 9 9 9 2
8 13 13 9 3 13 3 3 2
8 0 13 13 9 3 9 9 2
7 16 3 15 3 15 3 2
7 9 9 9 11 13 13 2
3 13 15 2
9 3 2 3 2 13 3 3 3 2
4 13 15 15 2
2 13 2
14 15 9 15 3 13 9 7 13 3 7 15 4 13 2
11 11 13 2 16 3 13 3 2 7 3 2
14 9 9 13 9 7 13 9 7 13 9 2 13 13 2
5 9 4 13 13 2
11 11 13 13 3 15 0 3 13 2 0 2
9 4 15 13 3 3 3 3 3 2
5 3 3 3 13 2
5 9 9 4 13 2
11 11 13 7 13 9 2 9 3 2 3 2
8 13 3 16 15 15 9 13 2
6 9 13 13 9 13 2
9 15 13 9 9 2 13 0 9 2
4 9 9 13 2
13 11 13 9 9 3 7 3 7 3 3 16 0 2
7 9 9 1 2 15 9 2
10 0 9 2 9 13 2 9 3 3 2
3 15 9 2
7 15 15 3 13 1 15 2
6 3 9 4 13 9 2
7 13 9 2 3 13 9 2
10 3 13 13 9 2 13 15 3 13 2
6 9 9 13 0 13 2
17 16 11 13 0 2 15 13 2 16 3 13 3 15 2 13 3 2
7 15 13 0 9 16 13 3
4 9 12 2 12
10 9 9 1 13 9 9 2 7 9 2
2 0 2
12 0 9 13 3 9 2 0 9 4 13 3 2
13 0 9 13 7 13 2 7 13 2 13 9 13 2
5 3 9 13 3 2
4 9 13 9 2
9 0 9 13 3 2 3 2 9 2
6 9 1 9 13 3 2
4 9 13 0 2
6 9 0 13 9 9 2
12 3 2 4 15 13 2 16 15 13 15 9 2
13 15 9 13 3 9 9 2 9 0 9 9 1 2
5 15 13 0 9 2
13 15 13 9 9 3 16 15 13 3 2 13 3 2
8 15 13 13 9 3 3 9 2
10 15 9 0 9 13 4 13 3 3 2
11 16 13 15 3 15 9 3 13 9 9 2
10 9 13 3 15 9 9 0 9 9 2
16 15 13 0 9 2 13 9 9 9 3 7 0 9 0 9 2
9 9 4 13 9 7 9 13 0 2
14 15 13 0 9 9 7 9 2 15 0 7 9 13 2
14 13 0 9 15 3 13 2 7 13 3 9 0 9 2
6 3 9 1 13 0 2
8 9 0 9 13 15 3 13 2
11 3 15 13 11 2 3 11 2 3 11 2
13 9 0 9 13 3 13 9 2 13 3 13 13 2
5 9 15 13 3 2
12 15 13 1 0 9 9 9 1 7 13 9 2
4 9 13 9 2
6 9 13 9 9 1 2
6 9 13 13 0 9 2
5 4 13 7 13 2
12 9 9 13 3 7 0 2 9 0 1 9 2
10 9 9 13 2 13 0 2 13 9 2
12 9 9 3 13 9 2 13 15 15 13 13 2
17 9 9 13 2 16 15 13 3 2 3 2 16 9 13 3 13 2
7 9 9 13 3 4 13 2
8 9 13 0 9 2 0 9 2
14 9 9 13 3 13 0 9 2 15 15 13 2 0 2
9 9 9 13 15 0 7 9 13 2
11 9 9 13 3 4 13 3 15 9 1 2
16 15 13 3 3 7 3 3 2 13 2 13 2 13 0 9 2
7 13 3 3 13 13 0 2
7 9 13 3 9 3 3 2
13 9 1 0 9 4 13 3 9 2 16 3 13 2
8 9 15 15 3 13 9 1 2
15 3 15 15 9 7 9 9 13 3 3 0 13 9 9 2
12 15 13 3 9 3 2 13 2 13 15 9 2
15 13 3 3 13 15 16 13 2 3 3 16 15 9 13 2
8 9 9 13 3 3 2 9 2
9 9 13 9 2 13 2 13 9 2
6 9 13 0 3 0 2
13 9 13 7 13 2 16 3 2 15 13 4 13 2
8 3 2 13 4 2 9 13 2
5 3 3 13 15 2
15 9 9 13 2 16 9 13 3 13 2 13 7 13 9 2
11 15 13 9 3 3 7 3 3 13 15 2
4 9 13 13 2
6 3 9 13 3 0 2
14 15 9 13 0 16 0 9 2 13 3 0 13 0 2
14 15 9 13 0 9 2 9 13 2 13 3 13 15 2
9 15 13 9 13 2 13 3 9 2
4 2 15 9 2
6 4 13 15 3 2 2
11 9 13 15 9 2 15 13 3 0 9 2
10 9 13 9 2 3 9 7 3 9 2
8 9 3 13 3 16 9 13 2
14 2 11 2 2 15 13 2 3 2 7 15 3 3 2
8 7 3 15 13 0 9 3 2
10 15 13 13 15 3 9 13 3 9 2
11 15 13 13 3 0 9 13 15 9 9 2
12 15 13 0 7 0 7 0 2 0 7 0 2
17 15 13 9 7 13 3 3 3 2 13 9 13 13 15 3 13 2
6 9 13 3 15 15 13
4 9 12 2 12
14 11 13 15 9 9 3 2 7 11 13 13 15 3 2
10 11 13 3 3 13 13 2 13 3 2
9 15 13 3 9 3 3 3 3 2
12 15 13 13 9 9 9 2 13 9 3 9 2
4 11 13 13 2
19 11 13 13 9 2 13 13 9 2 13 3 3 11 9 1 7 13 9 2
5 3 15 13 0 2
9 9 13 0 9 7 13 3 9 2
8 15 13 3 3 9 2 3 2
18 7 3 15 13 3 0 0 3 3 15 9 2 15 9 2 15 9 2
17 11 13 9 3 11 1 7 15 1 2 13 3 15 9 1 9 2
8 0 9 13 3 13 1 9 2
12 9 13 3 9 7 9 9 2 7 9 13 2
7 13 3 0 13 9 1 2
4 9 15 13 2
13 15 9 13 9 7 9 2 12 9 11 13 9 2
8 15 9 0 9 13 13 9 2
25 11 13 9 2 15 4 13 2 0 9 7 0 9 2 9 0 9 2 7 9 2 9 2 9 2
13 11 13 3 15 15 13 15 3 2 13 2 13 2
7 11 13 9 9 0 9 2
11 13 3 9 2 9 2 16 15 13 3 2
11 9 9 13 9 2 13 9 9 7 9 2
5 3 13 0 9 2
6 9 13 3 9 3 2
13 3 11 13 2 7 13 9 0 9 9 9 13 2
10 9 13 13 9 7 13 1 0 9 2
12 9 13 9 12 7 12 2 0 7 9 3 2
16 11 7 11 0 9 9 13 3 3 9 2 3 13 13 13 2
16 0 9 9 4 13 0 9 9 9 2 13 9 2 3 12 2
9 13 2 16 9 4 13 3 9 2
10 13 0 2 13 3 3 0 13 4 2
5 3 4 2 16 2
18 9 11 13 11 2 16 4 13 0 9 2 3 0 9 2 7 9 2
10 2 11 2 9 2 13 3 9 2 2
3 2 0 2
7 13 15 13 3 9 2 2
8 13 0 9 2 13 0 9 2
5 16 13 3 3 2
6 11 13 13 9 0 2
13 9 13 3 9 2 16 3 3 4 3 13 15 2
15 11 9 13 3 3 2 0 9 2 7 3 1 0 9 2
12 0 13 3 15 2 15 4 13 13 15 13 2
16 15 9 4 13 9 3 12 9 2 3 15 3 3 3 13 2
6 9 13 15 0 9 2
13 11 13 0 9 2 15 15 13 3 13 9 1 2
11 9 9 13 3 15 2 7 9 13 15 2
7 0 9 4 13 9 9 2
13 9 3 13 0 2 16 9 13 7 9 13 15 2
16 3 15 13 9 1 7 9 9 7 3 9 2 13 9 0 2
6 0 9 13 0 9 2
10 9 13 15 9 2 15 13 0 13 2
12 3 13 3 15 2 16 3 13 3 13 3 2
5 2 15 3 13 2
20 15 15 9 13 2 13 15 15 15 13 2 2 11 13 11 9 2 13 9 2
6 3 15 13 3 9 2
8 15 9 9 13 3 3 3 2
15 11 13 4 3 13 15 2 16 9 13 9 2 13 9 2
17 16 3 13 13 2 4 3 13 2 7 0 9 4 13 3 3 2
6 9 9 13 0 0 2
12 11 13 9 2 3 13 4 13 15 15 13 2
12 11 13 3 12 9 3 13 3 3 15 3 2
8 3 4 3 13 15 15 13 2
12 9 13 3 9 2 13 3 16 13 3 3 2
10 9 9 13 13 3 3 3 16 4 2
10 15 13 15 9 2 13 13 9 9 2
8 9 13 0 9 2 9 11 2
14 11 13 9 1 9 2 13 2 13 3 3 15 3 2
9 11 13 9 2 13 3 2 13 2
17 11 13 13 3 3 7 0 9 13 3 9 2 3 9 7 9 2
10 13 3 0 9 2 3 9 9 9 2
6 3 15 4 3 13 2
3 13 4 2
3 4 15 2
1 9
21 13 0 9 9 13 1 9 9 2 13 15 13 9 7 16 4 15 13 9 2 5
6 9 2 0 2 0 2
4 9 15 1 2
10 3 15 13 9 2 13 9 7 9 2
8 13 7 13 13 0 9 13 2
3 9 13 2
8 9 9 13 3 7 3 13 2
5 15 9 13 15 2
6 13 16 15 13 9 2
12 12 2 12 2 12 2 9 13 4 13 0 2
13 9 13 9 0 2 16 9 13 13 9 0 9 2
9 13 9 9 7 13 13 3 9 2
14 9 13 7 9 13 15 9 2 16 13 9 9 3 2
7 13 9 9 7 13 9 2
9 15 13 3 0 9 7 9 9 2
5 9 13 13 9 2
14 3 13 9 7 13 9 0 7 3 0 9 9 9 2
4 15 13 0 2
11 13 0 9 9 9 7 13 15 9 9 2
13 9 13 1 9 7 3 13 2 3 3 0 9 2
3 9 13 2
3 13 9 2
7 0 0 9 13 9 1 2
9 13 9 7 9 9 7 9 1 2
6 9 13 7 13 0 2
2 13 2
8 2 3 2 2 9 13 9 2
8 9 13 2 7 13 13 9 2
7 9 13 9 9 9 9 2
6 9 13 0 0 9 2
9 9 9 9 13 15 13 7 13 2
8 15 13 2 7 3 13 15 2
5 13 9 0 9 2
5 15 13 3 9 2
2 0 2
7 15 13 15 0 0 9 2
8 7 3 15 13 3 13 0 2
5 9 13 15 13 2
6 13 15 0 9 9 2
6 15 13 0 7 0 2
11 4 13 9 7 13 9 3 0 9 9 2
6 15 13 9 13 3 2
8 15 13 15 9 2 15 13 2
4 13 15 9 2
7 3 3 4 13 3 13 2
6 4 13 3 0 9 2
11 13 4 13 9 0 9 7 9 13 9 2
4 13 9 3 2
5 15 13 15 9 2
19 4 13 9 9 3 9 0 2 0 9 13 9 7 15 13 13 13 15 2
10 9 3 13 7 13 0 9 7 9 2
9 9 13 9 1 7 13 15 13 2
4 15 13 9 2
6 13 0 2 0 9 2
10 9 13 0 7 0 2 7 13 13 2
10 16 13 3 9 4 13 9 0 9 2
9 13 13 15 2 7 15 13 0 2
2 13 2
6 3 15 4 3 13 2
4 3 13 13 2
4 13 13 13 2
9 13 13 9 7 9 9 9 1 2
8 7 3 13 3 13 13 15 2
7 13 3 13 9 7 9 2
5 13 3 13 15 2
5 3 15 13 3 2
10 4 13 9 2 15 1 16 9 13 2
8 13 3 3 13 13 15 9 2
9 7 3 2 9 13 7 15 13 2
8 9 13 13 7 13 9 13 2
4 13 9 13 2
12 13 3 3 3 16 15 2 16 13 3 3 2
10 13 3 3 7 3 2 7 13 3 2
4 13 13 15 2
2 3 3
8 13 9 7 15 13 12 15 2
12 11 2 11 2 11 2 11 2 11 2 11 2
2 15 2
11 9 4 3 13 7 15 13 0 9 3 2
20 13 15 9 2 16 15 13 15 9 2 15 13 9 2 13 9 2 13 9 2
7 13 9 9 7 9 13 2
11 9 13 9 2 7 3 15 4 13 0 2
8 9 13 13 2 13 3 3 2
10 15 13 9 2 9 3 2 15 9 2
12 0 9 3 2 3 12 7 12 9 7 9 2
7 0 9 9 2 9 1 2
5 9 2 3 9 2
7 9 2 9 2 9 9 2
16 9 13 9 7 9 2 15 13 9 2 0 2 0 2 0 2
18 13 15 9 9 2 13 13 15 9 2 13 15 9 2 9 7 15 2
5 15 13 3 0 2
12 15 4 13 15 3 7 15 3 13 15 3 2
8 9 13 2 13 9 7 9 2
11 3 13 11 9 15 2 15 13 15 13 2
3 13 3 2
38 13 9 9 1 2 4 13 9 1 2 7 15 13 9 2 13 15 13 9 2 15 13 15 3 3 7 9 13 3 2 16 15 13 15 3 16 9 2
3 9 13 2
6 9 2 9 2 9 2
11 13 2 16 9 13 13 2 13 13 9 2
7 9 1 9 2 9 9 2
5 9 9 13 3 2
5 3 13 2 3 2
9 13 9 1 7 13 9 13 9 1
1 3
2 0 9
10 13 15 11 7 13 15 13 0 9 2
16 3 15 9 13 2 13 3 0 9 4 13 13 7 13 13 2
35 0 9 9 13 2 13 15 3 7 13 3 7 3 16 13 15 2 13 3 3 2 16 3 2 3 15 13 3 7 3 2 13 13 3 2
7 0 9 9 13 13 9 2
11 13 2 16 13 3 2 7 13 3 9 2
4 7 9 13 2
18 9 13 15 2 16 16 13 15 2 3 9 13 13 9 2 16 13 2
15 2 15 4 13 15 9 7 13 9 15 13 13 9 9 2
12 3 16 15 13 13 9 2 9 13 3 3 2
3 2 6 2
5 6 3 13 3 2
9 2 15 13 3 11 7 13 9 2
8 15 13 15 3 3 0 9 2
6 2 6 2 0 9 2
11 7 9 2 15 13 13 3 13 9 9 2
7 3 2 9 13 0 9 2
51 15 1 13 9 7 9 3 9 2 13 9 1 0 9 7 13 15 1 0 2 15 9 13 9 7 13 15 13 9 3 2 13 15 0 9 7 13 15 9 2 13 9 13 0 9 7 13 9 13 0 2
44 16 9 13 9 2 9 13 0 7 16 15 15 13 1 13 3 0 0 13 13 15 3 9 7 15 13 13 3 0 3 13 13 9 2 3 0 0 15 15 9 13 9 9 2
18 13 4 13 13 2 13 13 15 2 15 13 9 3 3 9 7 9 2
15 7 3 3 3 0 3 3 3 13 2 16 9 4 13 2
9 16 3 12 15 13 9 4 13 2
16 16 9 4 13 9 2 16 13 0 9 1 3 9 0 9 2
10 7 3 15 0 9 3 13 15 9 2
20 13 9 2 15 15 13 15 9 9 7 13 2 3 15 4 13 0 9 13 2
12 13 15 9 9 2 16 15 13 15 13 9 2
9 13 4 13 2 13 15 3 13 2
5 16 15 13 9 2
5 16 9 13 3 2
12 13 15 13 15 16 9 2 15 15 3 13 2
18 9 2 15 15 13 9 9 7 9 2 13 15 4 4 13 2 2 2
26 7 15 13 7 13 0 9 2 3 3 2 13 13 0 9 13 13 15 9 2 7 13 9 9 13 2
5 7 13 15 9 2
12 13 15 9 13 9 0 9 2 13 0 9 2
20 7 15 13 3 7 3 3 0 7 0 9 2 15 9 13 0 7 0 9 2
6 13 4 13 13 9 2
9 13 4 13 13 16 13 15 0 2
28 13 4 13 13 0 2 16 13 15 13 3 13 0 9 7 13 15 0 9 2 16 0 9 1 0 3 13 2
2 9 9
14 13 9 9 3 0 13 13 13 15 0 7 15 0 2
33 3 15 13 2 16 13 15 2 15 13 4 13 9 9 9 13 9 0 9 2 3 3 13 9 2 16 13 4 13 0 9 15 2
14 16 15 13 13 9 0 13 9 2 15 15 3 13 2
5 13 0 0 9 2
13 13 15 13 13 15 2 7 13 15 13 0 9 2
4 13 15 13 2
13 9 13 15 9 9 0 9 7 0 0 0 9 2
9 13 13 12 9 0 2 0 9 2
20 15 13 3 0 2 16 4 13 9 9 13 9 9 7 13 9 9 3 9 2
4 9 3 13 2
6 13 13 9 13 9 2
14 3 9 13 7 13 2 7 13 15 2 13 9 9 2
12 11 13 0 16 13 9 7 13 9 3 0 2
11 0 3 7 13 3 9 13 9 13 0 2
21 15 1 15 13 4 13 9 9 0 0 2 3 9 13 9 7 13 0 9 9 2
7 13 3 9 9 7 9 2
11 13 3 9 13 0 9 9 1 9 9 2
6 13 15 15 3 13 2
33 7 4 3 13 9 2 16 15 0 9 2 3 13 9 13 9 7 13 9 9 1 2 13 15 9 2 9 7 9 1 13 9 2
2 0 2
7 13 3 13 3 3 3 2
30 3 3 15 9 2 16 13 13 15 0 9 2 15 3 13 13 2 16 13 13 13 9 13 3 0 2 0 7 0 2
33 2 16 16 15 13 9 0 9 1 0 2 15 13 13 3 0 9 7 0 0 9 2 16 9 13 9 13 4 13 9 15 2 2
5 9 3 3 15 9
9 4 13 0 2 13 16 0 9 2
10 3 3 13 3 0 9 9 7 9 2
4 3 15 13 2
37 13 13 13 12 9 9 2 12 9 9 2 12 9 9 7 12 9 15 9 7 9 2 15 4 13 13 15 9 2 15 13 13 3 3 12 9 2
6 3 15 13 15 9 2
14 9 13 13 3 12 9 9 13 7 15 13 3 9 2
6 3 15 13 3 13 2
5 13 15 3 9 2
16 0 9 13 9 9 13 9 7 13 9 7 9 3 13 9 2
16 0 9 13 3 0 9 2 7 9 13 4 13 13 9 1 2
9 15 1 15 13 2 13 9 9 2
27 2 16 15 13 13 0 9 9 2 3 15 13 13 9 9 2 16 13 3 9 7 13 9 0 9 2 2
8 12 9 9 13 3 3 0 2
23 4 3 13 9 2 7 3 3 15 13 15 9 9 1 7 13 2 16 13 15 3 3 2
12 9 15 13 13 2 16 0 13 9 7 9 2
12 7 6 15 9 1 4 13 9 0 9 9 2
16 13 3 0 2 16 13 2 7 15 9 1 9 13 3 9 2
11 15 9 4 3 13 2 7 13 15 9 2
13 13 3 13 9 15 1 2 7 9 13 3 0 2
24 13 3 9 7 13 9 3 2 16 0 9 13 15 9 7 13 3 13 0 9 3 15 1 2
22 3 3 13 3 13 9 2 16 9 13 0 2 9 13 0 2 13 15 13 3 0 2
15 3 13 13 9 7 13 9 2 15 13 3 13 15 0 2
16 3 9 3 3 2 15 9 9 2 9 9 7 9 3 9 2
38 4 3 13 0 2 16 4 13 0 9 9 1 7 4 4 3 13 9 7 13 11 2 9 2 3 2 7 9 2 13 9 9 1 7 13 3 9 2
29 3 4 4 13 16 13 9 13 2 13 9 3 7 13 3 9 2 15 13 4 4 3 13 0 9 7 0 9 2
5 7 13 3 13 2
40 9 13 3 15 9 2 13 3 0 9 13 0 9 2 13 3 13 9 2 13 9 9 9 9 1 13 3 9 7 9 7 13 9 13 13 3 9 9 1 2
42 7 13 15 9 3 3 2 3 12 9 0 9 2 3 16 9 9 7 9 13 9 2 15 13 13 15 9 0 3 15 2 15 1 4 3 13 13 15 9 2 13 2
1 9
11 15 0 9 13 9 2 9 7 9 0 2
22 15 4 13 12 3 13 9 9 2 7 9 13 3 0 9 7 4 3 13 13 9 2
4 13 15 9 2
5 15 13 3 0 2
9 13 2 13 9 3 13 15 9 2
13 13 3 9 13 0 9 2 15 3 9 13 13 2
27 15 0 9 0 9 13 2 16 15 3 4 13 1 9 2 16 13 13 0 9 2 16 15 15 9 2 2
16 3 0 9 13 3 9 3 0 2 7 9 13 3 0 9 2
27 15 13 0 13 0 7 0 7 15 13 0 13 15 0 9 2 16 0 13 3 2 16 4 3 13 13 2
22 13 3 15 9 2 13 3 9 0 7 13 9 7 13 0 0 9 1 0 0 9 2
26 2 4 3 4 13 3 2 7 9 4 13 9 13 9 7 4 13 0 13 3 15 0 9 9 2 2
40 4 13 2 16 9 13 13 3 13 9 0 9 7 13 0 9 9 2 7 16 13 0 7 0 2 4 4 3 3 3 13 9 0 2 9 2 7 13 3 2
3 7 9 2
8 9 13 0 16 9 7 9 2
3 3 9 2
32 0 9 9 2 3 9 2 4 13 2 16 15 13 7 15 13 3 2 7 9 1 9 13 7 13 13 0 9 15 0 9 2
4 13 15 3 2
10 3 3 0 15 4 13 0 11 9 2
41 0 0 0 0 11 11 11 12 0 9 13 15 9 9 2 15 15 13 13 9 13 7 15 9 15 13 13 0 2 7 15 9 15 13 15 13 15 0 7 0 2
27 16 3 13 7 13 9 4 13 13 15 9 7 9 2 7 15 2 3 0 7 0 2 13 13 15 3 2
25 13 13 13 15 9 1 13 2 13 3 13 1 9 9 13 9 9 7 13 9 9 9 7 9 2
32 3 11 13 0 9 7 3 11 4 4 13 15 13 15 9 2 7 15 4 3 3 13 0 2 13 3 13 3 13 15 15 2
40 3 13 3 13 2 16 15 13 2 9 2 9 13 15 13 0 0 9 2 7 3 15 4 13 13 2 16 15 11 13 9 13 15 7 13 15 13 0 9 2
29 3 3 2 13 3 2 15 13 9 15 11 13 9 2 16 13 12 9 3 3 16 15 2 13 9 7 9 9 2
5 7 9 13 3 2
14 15 13 13 9 2 16 13 15 9 7 15 0 9 2
8 15 13 3 13 11 13 9 2
5 9 13 15 13 2
5 3 3 13 3 2
14 15 4 13 0 9 9 9 2 0 9 13 13 9 2
8 13 13 0 9 0 9 0 9
10 13 9 2 15 13 3 4 13 9 2
20 16 15 13 13 9 2 0 9 7 0 0 9 2 15 3 4 13 15 9 2
33 0 2 16 12 9 1 13 0 0 2 9 9 13 9 9 2 9 2 7 3 13 3 12 9 13 9 15 2 13 15 13 9 2
25 13 15 9 2 16 9 13 13 15 13 9 2 16 3 15 9 13 13 2 16 9 13 0 9 2
14 3 2 7 15 9 2 16 9 13 3 16 9 9 2
7 13 15 3 3 15 13 2
4 13 0 9 2
8 3 15 0 9 9 1 3 2
22 0 0 9 2 15 13 4 15 9 13 2 9 3 13 3 15 0 0 9 9 1 2
5 7 15 13 9 2
6 13 15 0 9 9 2
10 15 13 9 2 9 2 9 7 9 2
27 16 13 9 9 9 13 0 9 2 0 9 7 9 13 9 2 9 13 3 0 0 9 7 0 0 9 2
16 3 0 16 9 9 7 9 3 2 3 0 16 9 0 9 2
6 13 9 0 9 9 2
3 7 9 2
7 7 15 0 13 13 9 2
4 0 13 9 2
17 13 15 3 13 0 0 9 2 15 9 4 13 9 9 7 9 2
9 7 13 15 13 9 13 0 9 2
5 13 9 13 3 2
30 3 3 13 13 0 12 7 12 9 2 3 12 13 0 9 2 3 13 3 3 3 2 7 3 13 3 3 9 2 2
9 7 13 3 13 3 9 7 9 2
4 9 13 13 2
5 9 9 7 0 9
12 9 9 9 1 13 9 3 0 9 9 13 2
29 15 13 9 3 9 7 13 2 3 9 7 9 13 3 3 13 15 2 13 4 4 13 13 0 9 0 9 9 2
6 15 3 13 15 9 2
16 13 9 13 13 7 13 9 15 3 9 3 0 7 0 9 2
24 3 9 13 15 9 7 0 9 2 7 3 13 9 7 15 2 15 4 15 9 13 15 9 2
15 0 9 13 3 13 2 0 3 2 3 3 15 15 13 2
14 12 9 9 1 3 13 0 9 15 1 11 0 9 2
19 15 13 13 3 9 9 1 2 15 0 13 2 7 13 0 0 9 9 2
17 15 9 13 3 0 2 3 12 9 0 2 0 13 9 0 9 2
11 9 15 13 0 9 9 9 13 12 9 2
27 3 15 13 0 7 3 9 13 15 0 9 9 9 9 2 13 3 3 9 1 7 13 9 9 3 13 2
6 3 9 1 9 13 2
32 9 13 13 0 9 9 2 7 9 2 16 3 0 2 13 3 3 0 9 13 0 9 2 0 16 0 9 0 7 0 9 2
56 3 9 13 3 9 9 13 0 9 0 9 9 1 0 9 9 2 0 9 9 1 0 9 9 2 13 0 9 0 9 7 13 3 9 2 7 13 9 3 2 16 13 9 3 13 15 9 2 16 9 15 9 4 13 13 2
17 9 13 3 0 2 16 3 13 9 15 13 7 9 7 9 1 2
24 15 13 0 0 9 0 9 2 13 0 0 9 9 7 4 13 9 3 2 16 4 13 0 2
11 9 13 3 9 2 16 3 15 13 9 2
15 9 13 3 13 9 0 9 9 13 2 13 0 9 9 2
12 16 13 2 13 15 15 2 13 15 13 9 2
19 16 9 13 0 2 9 7 9 13 9 9 2 15 13 3 3 9 13 2
23 9 3 2 13 0 9 13 3 9 13 2 7 9 16 3 9 13 1 9 9 1 3 2
14 3 3 13 0 9 4 13 2 15 13 15 9 3 2
7 9 13 9 7 13 9 2
17 9 9 13 2 13 9 13 1 9 2 7 13 9 3 0 13 2
12 13 9 0 9 13 7 9 7 7 9 1 2
43 15 13 3 0 13 15 2 3 9 13 13 9 9 2 7 15 2 3 9 13 15 9 9 13 13 9 2 7 3 13 9 9 9 13 9 3 3 3 2 7 3 3 2
6 9 13 9 9 9 2
16 0 13 2 3 9 13 13 13 7 16 3 13 15 2 13 2
17 8 8 2 8 8 4 9 9 13 0 9 7 9 15 13 9 2
3 13 13 2
3 13 0 2
12 13 3 9 13 13 9 2 16 13 3 9 2
23 15 0 9 4 9 9 13 9 2 15 12 0 9 13 7 9 7 0 9 0 9 9 2
17 9 13 3 9 1 2 13 1 9 7 13 0 9 9 13 0 2
11 9 15 13 13 15 9 13 9 13 15 2
19 15 13 3 9 13 2 0 9 13 3 12 0 9 2 7 9 13 0 2
39 9 13 15 9 9 15 3 3 3 2 3 9 13 0 2 3 13 9 7 9 15 13 3 2 7 3 9 9 13 9 3 16 15 13 9 13 15 0 2
17 9 9 13 0 9 2 13 15 9 7 0 13 13 9 3 9 2
11 3 13 9 9 0 9 12 9 9 1 2
19 3 16 9 13 9 3 9 9 2 13 9 1 9 2 9 7 3 9 2
9 3 3 9 9 13 9 13 9 2
15 2 3 0 2 2 15 13 2 2 3 0 0 9 2 2
20 9 13 13 15 9 2 7 15 13 13 2 16 9 9 13 9 9 0 9 2
10 15 0 9 9 13 15 3 0 9 2
12 3 9 1 2 7 3 9 1 13 0 9 2
17 15 13 13 9 15 2 13 0 9 2 13 3 3 7 13 3 2
15 9 13 9 7 3 9 13 0 9 9 2 15 13 9 2
9 9 1 13 9 2 0 0 9 2
23 0 9 13 2 13 7 3 13 9 2 13 13 9 2 7 13 7 13 12 9 9 9 2
17 9 13 0 0 9 2 3 13 9 7 9 2 15 3 13 3 2
13 9 13 9 7 13 13 9 2 13 15 3 13 2
17 9 13 3 9 9 2 15 13 7 13 13 9 3 2 3 9 2
15 15 9 13 9 13 3 0 2 0 9 13 13 3 3 2
17 0 9 13 9 9 2 15 13 13 3 2 13 13 13 3 13 2
8 9 1 0 9 13 13 9 2
16 2 3 15 15 13 2 2 13 9 3 7 13 9 1 9 2
13 3 9 13 9 2 3 3 2 7 15 13 15 2
13 13 3 1 9 9 13 3 0 9 7 0 9 2
11 0 9 4 13 15 3 9 7 3 9 2
26 9 13 3 0 9 9 13 15 9 15 4 13 13 3 9 2 3 3 4 13 9 7 9 9 1 2
14 3 3 9 4 13 9 9 2 15 15 3 13 9 2
22 15 13 16 9 13 15 2 13 9 3 7 16 13 0 9 13 9 3 3 13 13 2
15 16 0 9 4 13 9 9 2 4 15 13 3 15 9 2
23 15 13 3 13 9 2 16 13 2 13 9 13 13 9 9 2 3 1 13 2 13 9 2
31 9 4 13 15 9 2 16 13 9 7 9 9 13 15 9 3 15 2 16 15 13 15 15 2 7 9 2 9 7 9 2
28 3 9 3 13 9 2 3 9 9 3 13 9 13 9 1 9 2 13 13 15 3 13 9 7 9 13 9 2
19 9 13 3 3 9 9 13 9 9 0 9 2 15 13 15 9 9 9 2
25 0 9 13 13 9 3 3 2 7 9 13 15 9 2 13 3 9 9 3 9 7 13 9 3 2
31 0 9 9 9 13 3 0 9 9 9 2 3 0 9 2 0 9 9 7 0 9 2 13 9 7 9 3 7 13 3 2
8 9 13 9 9 3 13 9 2
9 9 13 9 13 15 7 13 3 2
11 9 9 3 13 9 2 3 3 9 9 2
10 15 3 0 4 13 0 9 0 9 2
18 0 9 13 9 7 13 9 4 13 3 13 9 2 13 7 13 9 2
1 9
11 12 9 9 2 15 13 9 1 3 9 2
19 0 9 4 13 9 3 9 1 2 13 2 13 2 13 7 3 13 9 2
10 13 9 15 9 2 13 12 0 9 2
4 15 7 9 2
5 9 7 9 9 2
6 13 9 13 0 9 2
13 15 4 13 9 3 3 2 16 13 9 3 9 2
20 3 13 15 13 15 0 2 9 9 13 13 3 2 16 13 13 3 9 9 2
11 9 7 9 13 9 2 15 4 9 13 2
4 15 13 9 2
15 15 0 9 7 9 13 9 0 9 9 1 7 13 0 2
5 15 13 13 3 2
19 13 9 2 9 9 2 9 9 9 0 9 13 9 13 9 13 3 9 2
9 15 9 9 13 9 15 1 13 2
15 16 15 13 0 9 2 9 7 9 13 15 9 3 3 2
4 13 9 9 2
8 2 13 9 2 2 15 13 2
10 16 13 9 13 2 13 15 0 9 2
17 4 13 9 13 3 15 2 7 13 9 7 9 7 13 9 1 2
4 15 13 9 2
7 3 13 9 2 13 9 2
4 15 13 9 2
7 9 13 3 13 15 13 2
4 13 9 9 2
6 9 9 13 3 3 2
5 13 3 15 9 2
19 15 13 12 2 13 3 13 9 2 13 9 9 7 13 3 9 13 9 2
9 13 2 13 9 13 2 13 3 2
12 13 13 9 2 13 13 13 2 13 3 9 2
5 13 9 9 3 2
8 9 13 2 15 13 9 9 2
9 9 13 2 15 13 3 9 13 2
15 15 4 13 15 0 9 1 13 2 15 15 3 3 13 2
6 4 13 3 0 9 2
39 15 13 9 2 0 9 2 9 2 9 2 3 2 2 9 9 2 0 9 9 2 9 2 9 2 9 2 0 9 2 9 2 0 9 2 9 7 9 2
52 15 13 13 9 2 9 2 3 2 2 9 13 9 2 9 2 9 2 0 9 2 9 2 13 13 2 2 0 9 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 9 0 9 2 9 7 9 2
9 15 13 13 15 2 9 13 0 2
6 13 9 7 9 9 2
8 9 13 9 9 2 3 3 2
10 15 13 0 9 2 15 13 13 9 2
9 4 13 3 2 7 9 13 9 2
11 15 13 3 2 9 13 0 2 7 0 2
12 9 13 9 9 2 15 13 7 9 13 9 2
12 13 2 2 4 15 9 9 13 9 9 2 2
18 3 15 13 3 3 2 2 9 7 9 2 4 3 13 13 9 2 2
9 9 13 7 13 3 9 13 9 2
5 13 9 1 3 2
7 13 15 2 13 9 3 2
3 13 13 2
9 13 3 2 7 13 13 13 3 2
7 13 13 13 3 9 9 2
25 13 2 16 15 15 13 9 7 15 13 11 11 2 16 13 2 13 15 9 15 13 0 13 0 2
12 9 13 7 13 9 2 15 13 3 13 9 2
5 15 13 15 9 2
11 9 13 13 9 2 15 9 1 13 3 2
9 15 9 9 13 9 7 9 9 2
8 9 9 13 9 7 9 9 2
8 9 13 9 7 13 9 9 2
4 9 13 9 2
18 9 13 3 9 7 9 9 2 7 3 9 1 2 15 13 9 9 2
12 15 13 9 9 2 13 9 2 7 13 3 2
5 9 13 3 13 2
13 9 12 0 13 9 2 12 12 9 13 9 1 2
4 7 0 9 2
6 0 9 2 9 9 2
7 9 2 15 9 9 9 2
61 0 9 2 0 9 2 0 9 2 7 15 0 7 0 2 2 0 9 9 9 2 0 9 2 0 9 2 0 9 2 9 2 9 3 1 9 2 9 2 9 2 9 9 2 9 0 9 0 12 9 3 2 9 9 2 0 9 7 0 9 2
8 13 9 13 15 15 7 9 2
13 0 9 4 13 9 7 13 2 16 3 13 15 2
4 9 13 13 2
14 15 13 9 2 9 13 12 9 2 9 13 15 9 2
5 0 13 9 9 2
3 13 3 2
20 13 0 3 2 13 9 2 13 9 7 13 12 9 3 3 2 16 9 13 2
1 11
7 11 13 3 12 12 9 2
13 9 13 12 9 2 15 15 13 11 1 16 9 2
18 9 0 9 4 13 9 9 2 7 3 9 13 16 15 3 0 9 2
28 16 15 9 13 0 13 9 15 0 9 2 15 15 9 3 13 13 15 9 7 4 3 9 1 3 13 9 2
6 11 13 3 3 0 2
16 15 13 15 9 3 3 13 2 9 1 4 3 13 9 13 2
24 7 16 9 13 9 13 3 2 16 9 13 2 13 9 0 9 13 9 7 9 9 13 9 2
19 4 13 2 16 0 12 9 9 11 13 0 7 0 9 16 9 12 13 2
2 0 2
11 4 3 13 2 16 9 13 9 12 12 2
12 15 13 3 15 2 16 15 13 3 9 13 2
26 9 2 15 13 3 13 2 13 9 0 2 7 9 13 0 0 7 0 9 3 13 2 13 0 9 2
11 13 2 9 13 9 9 2 13 16 13 2
6 9 13 9 13 12 2
7 0 9 13 15 3 12 2
18 13 11 2 13 3 3 9 12 9 2 13 2 16 12 9 1 13 2
5 4 13 3 9 2
10 16 13 9 2 13 12 2 9 12 2
7 11 9 0 9 13 12 2
13 13 3 0 9 15 2 15 7 3 15 13 13 2
16 13 3 11 3 9 2 9 2 13 9 7 3 0 9 9 2
14 0 9 3 2 13 15 4 13 0 9 3 9 9 2
10 9 13 13 7 3 9 13 9 0 2
11 15 13 0 9 13 2 3 3 0 9 2
9 0 15 13 3 13 2 0 3 2
13 0 13 9 3 0 9 2 3 13 13 3 13 2
5 13 9 16 13 2
5 3 3 4 13 2
13 9 13 9 2 13 15 13 9 13 9 0 9 2
4 13 9 1 2
8 16 9 15 1 13 2 13 2
6 13 9 12 12 9 2
11 3 13 1 9 9 2 3 13 9 11 2
8 13 0 9 2 13 3 12 2
15 15 4 13 9 2 15 13 9 2 3 9 2 3 9 2
17 13 9 2 13 15 13 15 9 13 3 3 3 2 3 3 13 2
7 13 9 13 3 16 0 2
6 15 9 4 13 13 2
5 0 9 13 13 2
4 9 9 13 2
6 12 9 13 1 9 2
11 0 9 13 3 9 7 13 9 9 1 2
8 15 9 9 4 13 13 11 2
4 16 15 13 2
6 15 4 13 9 9 2
3 15 3 2
9 15 9 13 13 1 3 15 9 2
8 13 15 11 3 3 0 9 2
4 9 13 9 2
26 15 1 2 16 13 0 9 2 13 9 7 9 7 15 3 2 15 13 9 9 9 2 2 13 13 2
8 13 0 9 2 15 9 13 2
3 3 11 2
3 3 11 2
8 13 3 0 9 3 7 13 2
11 9 4 13 2 13 9 13 3 15 9 2
18 13 13 13 11 13 11 2 16 15 13 3 0 2 16 15 13 13 2
12 13 13 9 2 16 15 13 13 3 3 3 2
5 15 13 12 13 2
10 9 9 4 13 9 2 13 13 9 2
7 9 9 13 16 15 13 2
12 15 15 13 0 9 2 15 13 3 0 9 2
4 9 13 3 2
10 9 13 16 15 2 0 9 0 11 2
12 7 16 15 15 11 15 13 2 13 9 9 2
16 13 13 2 2 3 0 2 7 2 13 4 3 15 13 2 2
19 13 13 2 2 3 3 3 0 2 2 16 3 15 13 9 13 9 9 2
28 16 13 2 3 3 13 9 2 7 13 0 9 7 0 9 0 9 7 13 9 13 2 16 15 13 3 0 2
18 7 13 0 15 2 13 0 0 9 13 15 0 0 9 0 0 9 2
15 16 15 7 15 0 9 3 13 7 13 15 9 16 15 2
16 15 3 13 7 13 2 16 0 9 4 13 3 9 15 9 2
1 9
13 9 13 13 9 7 13 0 0 9 3 12 9 2
13 9 13 13 9 7 13 15 3 1 9 7 9 2
10 9 1 13 0 0 9 15 13 9 2
18 9 13 3 9 2 7 15 3 13 13 15 0 9 2 15 0 9 2
4 13 15 15 2
14 2 13 4 13 3 2 2 9 13 13 15 9 9 2
13 2 3 4 13 15 3 15 3 13 9 1 2 2
15 2 13 3 3 3 2 2 13 9 13 15 9 3 9 2
19 2 13 13 0 9 2 2 13 9 0 0 9 2 16 13 0 9 9 2
6 13 0 9 11 9 2
7 9 0 9 13 0 9 2
13 9 9 13 9 2 7 9 13 9 15 9 1 2
13 3 2 9 9 1 2 9 13 9 7 9 13 2
20 13 9 7 13 11 0 9 1 2 15 9 13 9 13 9 2 2 9 2 2
13 15 1 4 13 13 9 2 15 1 13 0 9 2
14 9 15 9 13 9 9 2 15 15 0 9 13 9 2
18 9 2 15 4 13 15 3 2 13 0 9 2 13 9 7 13 3 2
18 13 3 9 15 1 2 7 13 0 2 16 9 0 9 13 9 9 2
12 13 3 9 13 9 2 13 9 7 13 3 2
5 13 9 13 9 2
13 15 13 13 9 15 2 15 15 4 3 4 13 2
7 4 15 13 1 15 9 2
10 4 13 9 7 13 15 13 15 3 2
3 13 9 2
6 9 9 13 0 9 2
7 15 13 0 7 0 9 2
13 0 9 13 3 3 15 2 15 4 13 11 13 2
5 13 9 13 15 2
9 15 4 13 9 9 9 7 9 2
7 2 11 2 2 9 13 2
2 13 2
8 2 11 2 2 9 13 15 2
12 2 3 9 2 3 13 4 13 3 3 2 2
14 2 3 2 13 3 2 0 15 13 3 9 13 2 2
3 11 13 2
16 2 3 2 13 3 0 9 1 2 3 13 15 3 9 2 2
13 13 9 1 9 2 15 4 13 0 9 9 9 2
6 3 11 13 15 9 2
9 2 3 9 1 13 9 7 9 2
7 9 13 15 9 1 2 2
9 11 13 9 9 13 15 13 9 2
15 9 2 15 13 13 3 2 7 15 4 13 3 0 9 2
6 13 13 9 9 9 2
19 13 2 3 0 9 13 3 2 3 13 12 9 1 9 0 7 0 9 2
5 13 9 0 9 2
11 9 13 0 9 2 15 11 13 0 9 2
5 15 13 15 15 2
6 2 13 15 3 2 2
15 11 13 9 13 9 2 7 9 9 13 0 2 0 9 2
15 2 15 9 4 13 7 13 9 13 9 2 2 15 13 2
4 13 0 9 2
12 15 13 0 2 13 15 9 9 7 15 9 2
4 9 13 0 2
9 15 9 13 0 2 0 7 0 2
14 9 13 0 2 9 9 2 7 15 13 0 0 9 2
10 9 4 3 13 12 7 9 9 9 2
6 9 13 0 0 9 2
11 9 13 0 9 13 9 9 9 7 9 2
10 9 13 0 0 2 13 9 9 9 2
6 9 13 9 3 3 2
11 9 13 9 2 12 9 2 9 7 9 2
10 13 9 9 2 15 13 0 7 0 2
6 15 13 13 3 9 2
18 2 9 7 9 13 9 2 2 11 13 2 2 7 9 13 9 2 2
4 11 13 15 2
12 13 9 3 9 7 13 9 9 13 9 9 2
6 3 2 0 0 9 2
7 9 4 13 0 7 0 2
17 13 9 2 7 13 11 13 9 9 9 2 3 15 13 3 3 2
13 13 3 13 9 13 9 2 7 13 9 13 9 2
9 13 3 0 2 13 13 3 9 2
4 9 13 15 2
10 13 3 9 1 2 7 13 9 9 2
12 9 13 0 9 2 7 13 0 9 13 9 2
5 13 13 9 13 2
3 9 13 9
11 2 6 2 6 15 3 3 13 9 2 2
7 9 9 4 13 13 11 2
17 15 0 9 4 13 9 3 9 2 7 3 15 13 13 3 9 2
5 9 9 1 13 2
9 13 15 15 9 3 9 7 9 2
27 13 15 0 9 9 9 2 7 13 15 0 9 7 0 9 2 7 13 15 3 0 9 1 0 0 9 2
6 11 9 13 9 1 2
5 9 13 13 9 2
15 0 9 13 3 0 0 9 2 15 13 9 3 0 9 2
4 9 13 9 2
12 9 13 7 15 9 13 13 3 0 0 9 2
9 2 9 7 9 2 2 9 13 2
5 2 13 0 9 2
6 13 3 15 9 2 2
7 3 3 9 13 11 9 2
25 15 13 1 9 13 9 2 3 11 9 13 7 9 13 2 13 13 7 9 7 3 3 13 9 2
5 2 13 3 2 2
8 9 9 13 13 9 13 9 2
7 2 0 9 9 13 2 2
5 2 13 9 2 2
18 12 9 3 15 9 4 13 9 0 9 9 9 1 2 9 13 9 2
13 2 0 3 13 9 3 13 2 2 13 11 11 2
13 2 6 2 3 13 0 2 2 13 11 9 11 2
16 2 9 3 3 2 13 15 13 13 2 7 9 9 3 2 2
13 2 3 11 3 13 2 16 15 13 0 9 2 2
4 2 11 11 2
14 13 15 13 15 0 13 11 2 2 2 11 13 13 2
6 2 15 9 0 9 2
7 15 15 3 13 9 13 2
12 3 11 13 3 9 2 13 15 13 9 2 2
6 15 9 13 0 9 2
9 2 11 13 13 2 2 9 13 2
7 2 7 15 13 13 2 2
10 3 11 13 13 9 13 13 9 9 2
14 15 9 9 13 3 9 9 11 13 9 3 1 9 2
18 3 13 9 13 9 13 9 2 16 9 9 3 13 13 3 0 9 2
11 9 3 13 9 7 13 9 1 0 9 2
7 9 13 9 9 3 3 2
15 11 9 13 13 9 1 2 13 3 9 0 9 3 9 2
20 3 13 9 9 1 13 9 2 9 2 11 2 9 2 11 7 9 0 9 2
5 2 3 15 13 2
4 3 15 13 2
8 11 4 13 9 13 9 2 2
3 9 13 2
8 2 15 15 15 4 13 2 2
15 2 11 9 15 13 2 7 15 1 0 9 4 13 9 2
11 13 7 13 2 7 15 13 3 3 2 2
8 2 11 2 15 13 9 2 2
5 9 13 7 13 2
13 9 15 1 13 13 2 7 3 15 13 9 9 2
4 11 13 13 2
10 2 13 11 3 2 15 13 13 2 2
11 2 13 13 9 13 9 2 2 11 13 2
7 2 3 3 15 13 2 2
8 3 9 2 9 7 9 13 2
13 9 4 13 9 1 7 9 1 13 9 0 9 2
3 13 0 2
10 9 1 13 3 0 9 7 0 9 2
16 9 13 3 3 13 9 3 13 2 16 0 0 9 13 9 2
13 3 2 0 0 9 1 2 9 13 3 13 9 2
11 2 4 4 3 13 3 2 2 11 13 2
6 15 13 11 1 9 2
8 11 13 3 13 0 0 9 2
5 15 15 3 13 2
5 15 0 13 9 2
9 9 1 0 9 13 9 13 3 2
9 2 6 2 2 11 13 3 13 2
9 2 15 4 13 3 9 3 2 2
9 0 13 9 13 9 9 9 12 2
19 9 1 0 9 13 0 9 0 9 2 15 9 9 1 13 3 12 9 2
10 9 9 15 9 13 9 12 12 9 2
14 0 9 1 9 13 13 11 9 2 13 0 9 9 2
14 0 9 9 13 9 3 9 2 3 9 9 0 9 2
6 7 13 15 11 9 2
1 9
11 13 9 9 0 9 2 1 9 7 9 2
20 4 13 3 3 9 9 2 7 0 13 16 15 9 9 13 3 0 9 13 2
3 7 9 2
10 15 13 9 13 2 16 15 13 15 2
15 13 3 3 3 16 3 13 0 9 13 9 3 0 0 2
12 13 13 9 7 15 4 13 9 7 15 1 2
6 13 9 3 0 9 2
5 4 3 13 3 2
6 15 15 9 4 13 2
15 15 13 9 2 13 0 0 2 7 0 2 0 7 0 2
5 3 0 7 0 2
9 13 9 1 7 13 3 1 9 2
12 9 13 9 3 13 13 0 9 7 13 9 2
10 15 13 2 3 3 4 13 0 9 2
12 9 13 13 7 15 4 13 9 9 13 9 2
2 3 2
16 13 13 3 7 13 0 9 3 2 13 3 13 9 3 3 2
2 9 2
12 15 13 9 13 15 0 2 0 7 0 9 2
26 13 0 16 15 13 15 0 2 15 0 9 2 16 9 13 16 15 3 0 9 13 15 9 0 9 2
15 13 13 15 15 15 13 2 7 15 13 13 0 9 9 2
16 0 9 9 9 13 3 2 9 1 2 1 9 7 9 9 2
25 13 3 13 15 2 16 9 1 13 9 13 13 13 2 13 3 3 16 13 9 3 13 15 1 2
12 7 13 3 2 15 6 13 15 9 7 9 2
6 13 0 3 2 3 2
14 1 9 7 9 2 1 9 7 9 2 9 7 9 2
8 3 9 13 7 13 3 0 2
4 13 9 13 2
4 13 13 9 2
5 0 2 0 9 2
12 15 0 13 16 3 2 0 9 2 0 9 2
5 3 15 4 13 2
5 13 3 15 13 2
10 0 2 0 9 13 9 13 9 9 2
5 13 3 15 0 2
2 13 2
12 9 2 9 2 15 13 3 15 9 13 9 2
12 9 13 13 3 2 3 2 1 9 7 9 2
2 13 2
18 13 9 2 13 0 16 9 4 13 15 9 2 7 3 15 13 9 2
5 7 13 15 9 2
6 4 3 13 16 13 2
4 9 13 13 2
4 15 13 0 2
17 16 15 13 13 9 2 13 3 2 13 3 9 13 16 9 13 2
9 4 13 3 2 7 13 1 9 2
9 9 13 0 2 7 15 13 15 2
6 13 15 3 7 3 2
4 9 7 9 2
2 9 2
7 0 9 9 7 0 9 2
10 13 3 9 7 13 9 15 9 9 2
4 13 13 9 2
16 1 9 2 9 7 9 2 1 9 2 9 2 9 7 9 2
9 9 2 9 2 9 2 7 15 2
3 13 13 2
4 6 6 6 2
12 13 9 16 9 9 2 13 9 7 13 0 2
10 3 4 13 0 2 16 13 15 13 2
15 13 9 3 9 7 13 0 2 0 9 13 9 1 9 2
19 13 16 9 13 9 13 0 9 2 15 15 13 16 13 15 3 1 9 2
3 13 9 2
13 13 16 0 9 13 15 9 2 13 3 13 9 2
13 15 16 15 13 13 3 9 15 15 13 3 13 2
5 15 15 9 13 2
2 11 2
6 0 9 13 9 3 2
7 13 0 13 9 7 9 2
19 13 9 16 9 3 13 3 3 9 16 9 13 3 3 9 16 11 9 2
8 9 1 0 9 7 0 0 2
3 9 13 2
6 15 13 9 0 9 2
12 13 9 3 13 0 9 15 13 13 9 13 2
7 13 3 16 4 13 15 2
2 11 12
25 9 13 3 7 15 13 9 15 13 9 3 2 13 9 3 9 1 7 13 3 9 13 0 9 2
6 6 15 9 15 13 2
17 15 9 13 9 0 2 3 9 15 13 9 9 2 3 9 9 2
11 11 3 15 3 13 9 3 13 15 0 2
5 6 3 13 9 2
21 9 13 3 7 9 13 13 1 9 9 9 15 3 13 7 11 2 11 7 11 2
34 7 3 3 16 13 9 13 9 15 13 9 9 2 13 9 9 7 13 15 9 13 11 12 9 15 13 3 0 12 9 7 3 3 2
12 15 3 3 2 16 15 13 8 9 9 13 2
18 3 15 13 3 0 9 9 2 13 9 0 13 0 9 9 9 1 2
3 6 6 2
8 9 13 1 9 12 9 9 2
2 0 2
13 15 13 9 1 7 0 9 7 9 9 13 9 2
17 15 13 9 9 7 13 9 2 13 0 9 9 7 13 0 1 2
16 16 3 13 3 15 9 2 13 3 3 13 3 2 15 13 2
9 13 9 9 7 13 3 9 1 2
19 9 13 15 13 0 9 9 3 13 9 7 13 13 15 3 0 9 13 2
6 9 13 9 0 9 2
7 13 15 3 0 15 13 2
10 3 3 13 15 3 0 15 13 15 2
7 9 3 13 13 0 9 2
11 9 3 7 0 9 3 2 13 0 9 2
3 6 6 2
5 3 15 15 13 2
16 13 15 13 9 13 9 7 13 9 3 13 15 0 0 9 2
3 15 6 2
8 9 9 1 13 13 0 9 2
19 0 9 2 13 15 0 9 7 0 9 2 0 15 13 9 0 9 13 2
19 15 3 13 9 7 9 13 9 3 0 7 0 0 9 9 13 1 9 2
3 0 6 2
9 9 13 15 9 2 13 7 13 2
11 15 13 3 9 2 16 3 13 9 3 2
10 9 2 9 13 0 9 0 0 9 2
19 16 13 15 3 13 15 2 13 15 13 15 15 13 15 3 3 3 13 2
14 15 4 13 0 0 9 11 2 11 2 11 7 11 2
10 15 13 13 16 9 13 13 15 9 2
17 9 15 13 3 2 9 2 2 7 13 13 15 0 9 9 0 2
16 15 13 13 3 3 13 3 9 2 15 13 6 6 13 9 2
18 9 15 2 16 15 9 9 3 13 12 9 9 9 13 3 0 0 2
4 13 9 9 2
10 13 15 15 2 15 13 13 9 9 2
1 9
21 9 13 9 2 15 13 9 13 3 9 0 9 15 13 9 1 9 9 0 9 2
11 9 13 9 2 7 6 6 15 13 0 2
7 9 0 9 13 9 9 2
9 0 9 13 3 3 0 9 9 2
5 0 0 11 11 2
5 0 9 9 9 2
8 9 13 3 3 9 7 9 2
10 15 9 9 13 0 2 0 7 0 2
9 9 13 0 7 13 9 13 9 2
9 13 9 9 7 13 9 15 9 2
15 13 11 9 7 11 11 11 2 11 13 13 9 9 9 2
9 13 9 3 7 13 13 9 9 2
6 13 9 13 9 1 2
8 13 9 0 7 13 3 3 2
17 1 9 9 9 13 9 9 1 7 13 9 0 9 9 1 9 2
4 11 11 13 9
14 4 13 9 16 9 13 13 7 13 3 0 15 9 2
6 3 13 0 9 9 2
6 3 13 3 9 9 2
12 3 9 13 3 4 13 7 9 13 9 9 2
16 13 13 9 9 1 7 13 9 9 0 13 15 9 9 9 2
23 9 13 3 7 9 1 13 0 9 2 15 13 0 9 9 3 3 3 12 9 1 9 2
15 15 0 9 13 1 9 7 13 9 9 1 0 9 13 2
4 11 11 13 2
9 9 7 15 9 13 13 13 3 2
21 9 9 4 13 0 9 0 7 3 13 0 7 0 2 3 0 9 1 3 13 2
3 2 9 2
9 13 15 3 3 9 3 9 2 2
12 13 9 9 9 2 15 13 9 13 13 9 2
7 2 13 13 0 9 2 2
12 9 13 13 7 13 13 13 15 3 9 1 2
16 2 3 6 15 13 3 0 15 2 13 3 15 1 13 2 2
14 9 9 13 3 13 2 7 13 13 15 13 0 9 2
9 13 9 3 9 7 13 9 13 2
11 9 13 13 11 11 11 2 15 3 9 2
7 9 13 3 0 9 9 2
19 0 9 13 9 9 2 13 0 9 9 7 15 9 13 9 13 13 9 2
22 3 9 1 15 4 13 9 3 3 9 16 9 13 9 9 7 15 13 3 3 13 2
17 13 13 15 3 13 9 2 7 13 4 9 9 13 0 15 9 2
8 13 4 2 7 13 15 13 2
5 3 13 0 9 2
3 9 3 3
16 15 9 9 9 7 9 1 13 3 15 9 2 15 3 0 2
6 13 15 9 7 9 2
2 9 2
5 3 15 13 3 2
5 3 15 13 9 2
13 3 2 13 15 3 13 2 13 3 7 13 9 2
3 15 9 2
2 15 2
11 15 13 9 7 15 9 13 0 9 9 2
15 16 9 13 9 15 13 2 6 2 15 4 13 13 2 2
13 16 9 13 9 2 15 13 2 13 0 9 2 2
11 16 9 13 3 2 13 2 3 6 2 2
17 3 16 13 9 13 9 13 9 2 16 13 3 15 9 13 13 2
34 9 15 13 0 13 9 2 9 0 7 3 13 9 2 15 0 7 9 4 3 13 13 9 7 13 3 13 9 2 13 13 15 9 2
3 9 13 9
7 2 13 2 15 4 13 2
4 15 13 13 2
5 2 15 13 13 2
4 2 15 9 2
3 2 9 2
5 15 9 15 13 2
8 2 15 13 3 13 15 3 2
12 2 15 4 13 12 9 3 7 13 12 9 2
3 3 6 2
6 15 13 13 15 3 2
5 13 3 13 3 2
5 13 15 15 15 2
8 6 6 9 15 13 15 15 2
7 2 13 15 13 15 15 2
5 15 13 3 13 2
11 15 4 13 15 13 3 3 13 15 9 2
3 2 9 2
4 13 13 9 2
8 6 4 15 13 13 15 9 2
6 3 6 15 1 9 2
3 3 9 2
5 3 15 12 9 2
20 2 16 15 13 3 3 13 13 3 3 3 3 13 9 1 7 13 9 1 2
1 9
4 2 9 1 2
4 2 3 11 2
4 2 9 1 2
3 2 6 2
3 9 13 2
2 3 2
7 2 3 6 15 13 15 2
3 13 3 2
9 15 13 15 9 7 15 13 15 2
6 13 3 15 15 13 2
2 13 3
14 15 13 3 4 9 13 3 0 3 16 15 3 13 2
11 9 9 9 13 15 0 9 9 2 3 2
12 9 3 13 9 9 2 9 7 9 9 9 2
7 15 13 9 7 13 13 2
3 3 6 2
3 13 9 2
15 13 15 3 0 9 2 13 15 9 1 9 2 3 3 2
19 13 3 13 9 0 2 7 3 13 0 9 0 9 2 16 13 15 13 2
6 15 15 3 13 9 2
7 13 16 9 13 9 9 2
19 9 13 3 0 2 13 16 4 13 15 9 2 7 3 15 0 13 9 2
10 3 16 13 2 3 13 13 15 9 2
7 13 3 3 3 15 9 2
13 9 13 7 0 9 13 9 1 1 0 9 13 2
10 3 15 15 13 3 0 9 0 13 2
8 3 13 13 3 3 3 9 2
10 3 15 9 2 9 13 13 3 0 2
10 15 13 3 16 12 0 9 12 9 2
12 16 13 9 2 9 13 13 9 16 13 9 2
7 9 3 9 13 3 0 2
17 13 0 9 0 2 7 0 0 9 2 3 16 9 4 9 13 2
3 13 13 2
11 3 13 9 13 2 9 13 3 9 13 2
14 13 15 0 9 2 7 0 9 0 2 3 0 9 2
1 9
4 15 13 9 2
12 13 13 15 0 9 2 7 4 13 9 13 2
8 15 13 9 13 12 9 9 2
10 3 3 15 4 13 9 2 15 13 2
14 13 7 9 7 3 9 9 13 2 15 13 3 13 2
12 15 13 15 13 15 9 2 3 15 13 13 2
5 15 9 15 9 2
10 7 15 15 13 0 2 15 13 9 2
13 15 13 3 9 3 3 15 9 13 13 3 13 2
7 3 15 13 15 9 9 2
17 7 15 13 0 9 7 9 9 2 15 15 9 4 13 13 15 2
14 9 13 3 9 13 9 9 2 13 7 13 15 1 2
13 9 13 15 2 7 13 3 9 13 0 9 9 2
10 12 15 9 2 15 13 0 9 9 2
4 2 9 3 2
5 9 3 9 1 2
7 3 13 13 3 13 9 2
9 15 13 15 9 16 15 13 9 2
12 3 15 3 13 13 3 9 12 15 9 1 2
14 6 6 2 15 13 3 3 0 9 12 15 9 1 2
18 15 13 13 13 15 9 2 15 15 4 13 7 4 15 13 0 9 2
10 15 13 9 2 13 9 7 13 13 2
10 3 15 13 3 0 9 2 0 9 2
6 2 15 13 9 3 2
22 3 3 2 13 15 3 13 15 9 2 7 9 13 0 0 7 15 13 0 9 9 2
18 9 15 4 13 9 2 13 15 9 2 15 1 0 0 9 3 13 2
12 3 0 9 9 2 7 15 9 13 3 3 2
20 15 4 3 15 9 13 13 3 0 9 0 3 13 9 3 3 15 7 15 2
11 16 13 16 15 13 15 4 3 13 15 2
21 16 13 13 0 4 3 13 15 0 2 7 6 6 2 15 3 15 13 13 0 2
13 3 0 9 1 15 13 16 3 15 13 15 0 2
15 2 9 9 7 9 9 9 2 16 9 13 13 9 3 2
11 15 13 13 0 13 15 0 7 0 9 2
9 9 13 3 0 7 0 16 3 2
13 16 12 9 13 3 2 13 16 15 15 13 3 2
21 9 13 3 9 3 2 7 16 12 9 9 13 9 9 9 1 15 13 13 15 2
6 15 13 7 0 9 2
7 2 15 13 3 9 9 2
25 9 1 13 15 9 16 9 2 16 13 13 9 13 9 7 9 13 2 13 3 4 13 0 9 2
21 7 3 16 15 4 13 15 13 13 2 9 9 0 7 0 13 13 9 15 9 2
6 0 15 13 13 9 2
17 15 13 3 16 15 13 3 13 9 13 9 9 7 0 9 9 2
9 2 15 13 13 3 15 9 3 2
10 15 13 13 2 13 15 13 3 2 2
8 9 13 13 15 9 0 9 2
7 3 13 9 9 2 9 2
25 15 13 0 9 7 3 9 13 15 0 7 3 9 13 9 7 9 9 3 15 13 3 13 0 2
7 9 9 7 9 9 1 2
14 13 15 0 2 13 9 7 3 3 13 15 9 15 2
8 15 13 2 3 9 13 9 2
10 9 13 7 15 13 13 12 9 13 2
5 13 9 13 9 2
2 0 9
10 13 9 9 13 9 13 9 0 9 2
8 15 9 13 13 3 3 9 2
16 4 1 9 13 3 16 13 9 9 2 7 4 13 0 9 2
11 0 13 3 0 2 3 0 13 0 0 2
8 6 13 3 9 3 1 9 2
15 15 13 13 13 13 9 7 15 4 13 0 15 13 9 2
15 13 9 13 9 16 13 9 9 9 2 3 0 9 13 2
15 13 15 3 7 13 15 9 13 3 9 9 13 9 1 2
8 13 3 13 3 15 13 9 2
23 3 13 12 9 9 2 15 0 9 9 13 3 3 2 7 15 0 9 9 13 3 0 2
12 13 13 9 16 4 13 9 9 1 3 3 2
22 15 9 2 15 3 4 13 13 13 9 15 2 13 0 9 13 15 3 16 4 4 2
20 13 0 0 0 9 9 2 16 13 3 13 9 15 1 15 9 13 3 9 2
9 13 0 9 7 13 9 2 9 2
19 15 3 3 9 4 15 13 2 9 2 2 0 9 13 3 15 13 9 2
6 13 13 9 15 3 2
20 3 0 9 13 9 4 3 13 9 2 7 9 4 15 9 13 9 15 9 2
18 13 13 15 2 16 3 9 4 13 3 2 16 9 13 13 3 0 2
17 6 2 13 13 9 9 2 7 13 16 15 13 3 0 0 9 2
18 3 16 13 13 0 9 3 2 13 13 15 9 13 13 15 9 3 2
21 13 3 13 16 3 6 15 3 13 2 7 13 9 2 9 9 2 13 15 15 2
11 13 3 9 3 7 13 15 13 9 3 2
8 13 13 13 9 3 13 9 2
27 3 2 13 3 0 9 9 2 13 16 9 2 0 0 2 13 3 3 9 2 13 15 13 0 9 9 2
15 13 16 9 4 13 15 3 16 13 13 15 0 9 9 2
12 13 16 15 15 3 2 13 2 7 13 9 2
6 13 4 3 13 3 2
17 13 9 15 13 0 9 9 2 7 13 9 15 9 13 0 9 2
23 13 9 3 2 7 13 3 9 2 9 13 3 13 9 2 7 15 13 9 7 15 13 2
10 13 9 2 13 13 0 9 15 9 2
5 13 3 13 9 2
15 13 13 9 13 3 15 9 3 15 9 15 4 9 13 2
21 13 3 12 9 2 13 9 15 13 0 0 2 13 16 15 13 3 9 0 9 2
11 15 9 13 13 3 9 2 13 3 9 2
12 9 9 13 9 9 2 7 9 13 9 9 2
10 13 9 9 13 15 9 3 3 3 2
7 9 13 13 13 3 9 2
12 13 9 1 7 13 13 13 9 13 9 15 2
17 13 3 3 15 4 13 2 7 13 15 9 2 13 3 13 9 2
6 6 3 13 2 13 2
11 13 3 0 9 2 7 13 9 9 3 2
14 9 13 13 16 13 15 3 9 2 13 16 9 9 2
17 3 13 13 9 15 13 9 2 7 13 3 3 2 9 7 3 2
6 7 13 3 0 9 2
15 13 15 9 3 2 7 13 3 15 13 0 9 2 13 2
15 13 15 3 2 7 13 16 13 13 3 9 2 3 9 2
18 9 13 0 9 3 2 7 9 15 13 2 13 13 0 9 15 9 2
4 13 3 3 2
9 0 2 9 4 13 3 15 13 2
8 13 13 7 13 15 13 3 2
8 16 13 9 3 4 15 13 2
9 9 13 3 2 0 13 13 9 2
5 3 13 7 13 2
3 7 13 2
10 13 13 3 13 2 7 3 9 13 2
10 13 3 9 2 7 3 13 0 9 2
5 9 9 7 9 2
15 9 13 3 9 7 15 9 0 9 15 9 13 9 13 2
4 13 3 9 2
10 3 3 13 9 2 15 3 0 9 2
8 13 3 9 2 13 3 9 2
3 9 13 2
9 15 13 9 15 13 15 4 13 2
24 13 7 13 9 2 7 15 13 15 13 0 9 15 3 13 11 2 7 0 15 13 13 11 2
7 13 15 16 13 3 3 2
12 13 13 9 15 9 2 16 3 15 4 13 2
14 9 13 3 0 9 2 3 15 4 15 13 15 3 2
10 0 9 15 13 2 13 0 0 9 2
7 15 13 3 9 2 3 2
10 13 9 7 15 13 3 13 15 13 2
22 15 13 13 3 4 13 2 7 9 15 9 13 9 13 15 2 15 13 13 15 9 2
6 13 3 13 15 9 2
11 13 9 2 13 3 9 7 13 9 3 2
13 3 13 9 15 13 0 9 2 13 9 3 3 2
1 9
17 15 9 4 3 13 0 11 9 2 3 16 3 13 13 3 9 2
23 15 9 4 3 13 3 15 16 3 15 9 13 3 3 2 7 9 1 15 4 13 9 2
24 6 3 13 15 9 2 15 15 11 3 13 7 13 13 13 2 7 15 9 13 3 15 9 2
22 6 13 15 4 15 16 13 15 9 2 16 13 9 4 9 13 2 7 9 13 13 2
25 9 4 3 13 0 13 9 1 3 2 15 13 13 3 13 3 7 15 4 13 13 15 3 3 2
47 3 15 4 13 9 2 15 13 16 16 15 9 13 2 3 3 13 15 2 7 9 13 16 15 13 15 9 9 3 2 15 4 13 7 0 9 13 13 15 13 2 16 3 4 13 9 2
30 7 15 1 13 9 3 13 2 3 15 0 9 2 13 15 3 0 16 15 2 7 0 16 9 2 3 15 13 9 2
14 16 3 16 9 13 9 2 3 9 13 3 13 9 2
22 3 2 15 13 0 9 3 3 2 16 13 13 13 3 13 16 9 13 9 7 9 2
30 6 15 11 2 15 13 15 0 9 0 9 7 15 13 0 9 15 9 9 2 3 3 15 9 16 12 15 12 9 2
19 15 13 15 2 16 3 15 11 4 3 3 13 3 2 15 15 13 9 2
5 3 15 15 9 2
36 9 15 13 9 15 2 16 9 13 15 9 2 3 15 13 13 11 3 9 9 2 7 3 15 16 15 9 2 15 11 13 2 1 13 15 9
31 3 15 13 3 13 11 1 2 7 15 13 13 15 9 2 7 13 3 3 3 15 9 15 15 4 4 3 13 9 1 2
23 3 15 13 9 15 9 9 13 9 9 2 15 13 16 9 9 15 13 3 13 9 3 2
20 15 9 13 3 3 0 2 9 9 2 4 4 15 9 9 13 0 9 1 2
12 6 13 15 15 2 13 9 7 13 13 9 2
16 15 9 9 13 3 0 2 7 15 0 9 13 3 3 3 2
16 7 15 0 9 13 15 9 9 2 15 13 13 3 9 9 2
7 7 9 2 15 9 13 2
19 3 15 13 3 0 2 9 9 3 9 2 7 11 13 13 9 9 3 2
24 15 13 3 13 9 0 16 4 4 3 3 13 11 3 2 13 15 4 13 15 3 3 3 2
24 15 9 9 13 13 3 15 9 2 7 15 4 3 3 13 13 2 16 13 3 4 9 13 2
23 3 15 13 16 11 13 15 9 9 1 2 7 13 2 16 3 9 15 13 13 9 9 2
8 15 15 9 4 13 15 3 2
13 3 2 15 13 15 1 16 9 9 9 13 9 2
14 9 2 9 1 2 0 9 9 13 13 15 9 9 2
33 7 16 15 13 3 9 9 9 13 15 15 9 9 2 3 13 16 11 3 9 13 0 9 2 3 15 13 9 3 7 13 3 2
24 3 16 15 9 9 2 3 9 9 4 3 13 15 9 3 2 13 11 13 7 3 9 1 2
18 15 13 13 3 3 15 9 2 7 3 4 13 2 11 13 15 9 2
7 13 15 9 7 13 9 2
14 0 9 2 9 13 7 12 9 13 2 7 15 13 9
23 15 13 9 2 15 13 13 16 15 13 3 13 3 2 9 15 13 4 15 9 3 13 2
37 13 9 13 3 9 2 13 15 16 13 11 15 9 3 13 2 7 15 0 13 3 15 1 7 13 13 16 15 15 15 9 13 3 3 15 9 2
28 13 3 15 2 7 13 16 13 15 13 16 15 13 0 9 9 2 7 16 3 16 13 2 3 3 9 13 2
13 13 16 3 3 2 15 9 13 3 0 9 11 2
28 11 13 15 0 9 2 9 1 2 7 15 4 3 13 15 3 9 9 2 3 3 9 13 16 15 13 0 2
11 15 13 12 9 3 15 13 13 9 13 2
17 3 15 13 9 13 15 15 15 13 7 15 9 15 15 9 13 2
15 3 9 13 16 13 16 15 9 4 13 3 15 9 9 2
17 15 13 16 13 3 9 2 7 13 15 9 15 13 15 9 13 2
14 3 11 13 15 3 2 3 2 3 13 9 15 9 2
33 15 9 4 13 15 9 3 3 2 13 3 13 3 3 9 13 2 7 16 3 13 13 15 2 9 13 3 9 9 9 9 9 2
14 9 13 3 3 2 16 13 9 13 3 3 9 9 2
7 3 13 4 3 9 13 2
18 13 9 3 2 7 9 13 3 3 13 15 9 13 11 3 15 9 2
45 15 13 12 9 2 4 4 13 9 9 9 2 3 4 13 11 3 9 7 3 3 9 13 2 7 3 4 13 0 9 2 16 9 9 4 13 15 15 9 7 15 3 3 9 2
30 13 13 3 13 11 9 1 2 3 15 9 4 13 9 3 3 2 16 13 9 13 15 9 16 4 13 12 13 9 2
21 3 15 13 9 3 13 3 2 15 13 9 15 16 9 1 9 13 13 3 3 2
19 3 13 2 11 7 15 2 9 13 3 3 0 9 1 2 9 3 3 2
15 13 13 9 15 2 9 15 9 0 9 4 13 3 0 2
22 3 16 9 3 13 15 1 2 13 3 9 13 2 16 15 1 9 13 3 0 9 2
20 15 9 3 0 9 13 2 16 13 9 9 13 9 7 13 13 15 3 3 2
13 9 4 3 13 9 13 2 13 3 3 9 1 2
23 13 3 15 9 2 3 16 3 13 13 9 0 9 2 15 9 0 9 15 3 3 13 2
17 13 9 2 16 13 15 13 15 9 13 2 16 13 13 3 9 2
15 9 13 13 0 0 9 15 13 9 9 3 3 9 1 2
14 15 13 9 9 3 13 2 7 13 13 13 9 3 2
19 15 13 11 1 9 2 7 9 13 0 2 15 0 9 15 3 13 3 2
6 13 9 2 13 11 2
18 13 9 1 13 0 9 2 7 9 0 9 13 15 13 0 0 9 2
11 4 13 9 9 3 2 7 13 13 9 2
5 13 15 13 9 2
24 16 13 12 9 2 13 13 11 9 13 0 9 3 2 7 9 3 13 3 15 0 9 11 2
22 13 3 0 9 9 2 7 13 13 9 2 3 9 2 16 11 13 13 15 9 1 2
24 16 11 7 3 13 9 9 2 9 7 3 9 13 2 13 13 3 9 3 3 15 13 9 2
25 9 13 13 9 9 13 2 7 3 3 15 9 11 9 13 2 13 13 15 12 3 13 9 13 2
17 16 9 13 2 13 13 3 7 13 13 13 0 9 1 9 1 2
14 9 13 3 3 12 9 2 7 13 9 3 7 3 2
9 3 13 13 9 13 9 0 9 2
9 9 7 9 9 13 9 3 9 2
19 9 3 13 9 9 2 15 13 3 3 7 9 9 9 2 13 11 9 2
21 9 13 13 3 15 2 13 3 9 15 2 16 11 13 13 9 3 13 9 1 2
15 9 4 13 9 3 3 16 13 13 11 3 3 16 15 2
1 9
4 13 3 9 2
4 13 13 3 2
8 15 9 13 3 3 13 15 2
15 15 13 13 13 15 3 2 13 4 13 0 9 0 9 2
15 9 13 3 0 2 3 15 9 13 9 2 9 15 9 2
9 16 13 2 3 13 9 9 9 2
11 3 2 16 13 2 3 13 15 15 13 2
13 13 0 13 15 15 4 13 2 16 15 13 9 2
19 16 4 3 13 9 9 2 13 4 13 9 3 2 3 9 4 13 3 2
3 7 9 2
10 13 3 13 3 4 13 3 9 9 2
34 13 0 9 13 9 3 0 2 13 9 2 13 15 13 3 3 9 2 7 16 13 0 9 2 3 15 13 4 13 2 13 13 13 2
14 3 2 3 16 3 13 2 13 3 13 3 15 13 2
15 13 3 0 2 16 9 4 13 0 15 7 13 13 0 2
11 15 13 15 2 3 13 13 3 15 13 2
7 13 15 3 0 9 13 2
29 15 9 2 15 9 13 11 2 4 13 15 9 9 9 2 9 15 13 15 9 15 9 2 3 13 13 9 15 2
15 6 2 13 13 3 3 2 7 9 13 13 3 13 9 2
13 7 3 11 13 9 2 3 13 15 9 0 9 2
6 3 2 13 3 9 2
9 15 9 13 15 9 13 9 0 2
11 7 3 2 13 13 15 9 9 3 13 2
7 7 3 2 13 3 9 2
1 9
21 0 1 4 13 13 9 2 13 9 0 9 7 13 9 2 16 9 13 13 9 2
16 15 13 9 2 15 9 7 0 9 2 15 15 13 3 9 2
24 13 15 13 9 0 7 0 9 2 15 13 13 3 0 9 1 7 13 9 7 9 1 9 2
18 13 15 9 2 13 15 9 2 4 13 0 9 2 15 13 7 13 2
13 13 9 0 9 9 3 13 9 7 15 13 9 2
5 13 13 13 0 2
10 13 3 9 9 9 7 13 15 3 2
11 9 13 3 13 2 7 15 15 13 9 2
11 13 3 13 9 2 3 13 3 13 3 2
15 3 9 13 13 2 7 13 3 3 0 7 0 9 13 2
6 3 3 15 9 13 2
6 7 15 13 0 13 2
19 13 15 4 3 13 3 9 15 9 2 0 16 3 13 15 3 9 13 2
10 16 3 13 3 2 13 3 9 9 2
12 13 2 16 4 13 9 3 2 16 9 13 2
6 9 15 13 2 3 2
8 13 0 9 9 13 2 13 2
5 15 13 12 9 2
18 15 0 7 0 2 7 9 13 13 3 13 15 15 9 2 15 13 2
6 9 13 3 13 9 2
5 3 13 13 9 2
18 13 3 2 15 9 3 2 7 3 3 2 16 15 13 3 0 9 2
10 13 9 9 9 7 13 9 13 9 2
15 15 13 2 16 13 9 2 7 15 9 13 3 13 15 2
6 13 13 3 2 13 2
5 13 13 9 9 2
5 9 13 9 9 2
9 3 15 13 13 13 9 13 9 2
9 15 13 9 7 13 15 9 15 2
10 9 13 9 2 7 15 13 9 15 2
2 15 2
19 15 13 15 3 2 7 9 4 13 3 0 9 0 2 16 9 13 9 2
11 9 13 9 9 13 2 16 9 13 9 2
8 15 15 13 13 9 16 15 2
8 15 15 3 13 12 0 9 2
11 13 9 2 9 9 13 2 7 9 13 2
17 15 13 1 9 9 7 13 3 13 9 7 13 9 13 9 1 2
5 15 13 3 0 2
5 3 13 9 9 2
10 15 13 9 7 15 13 9 15 9 2
12 13 13 2 13 15 0 9 7 13 15 9 2
5 9 13 9 9 2
11 4 13 15 0 2 13 9 3 13 3 2
7 13 9 9 7 13 9 2
9 15 13 15 13 7 13 3 9 2
6 13 1 9 7 9 2
8 13 1 7 1 9 7 9 2
9 3 15 13 15 3 7 13 3 2
5 3 13 13 9 2
3 15 13 2
4 15 15 9 2
14 13 0 9 9 0 0 9 2 15 13 0 0 9 2
18 15 9 13 3 0 9 7 15 0 9 13 0 9 9 9 3 9 2
17 15 15 13 0 9 2 7 9 9 9 13 3 15 9 9 9 2
24 3 9 13 0 9 2 15 15 13 15 9 9 7 3 13 3 15 2 15 13 3 0 9 2
14 15 0 9 13 9 7 13 9 9 9 7 15 9 2
27 13 15 15 9 2 13 3 9 9 13 7 13 9 3 13 0 9 0 9 2 15 15 9 4 3 13 2
23 3 9 9 2 15 3 13 0 9 2 13 15 9 1 7 13 3 3 0 3 0 9 2
16 3 15 13 9 9 0 9 13 0 9 7 13 15 3 9 2
13 15 9 2 15 9 3 2 13 3 3 13 9 2
19 7 3 15 13 13 9 7 3 2 16 15 13 9 2 15 9 13 9 2
16 9 13 3 2 15 13 3 13 9 7 15 9 13 9 9 2
16 0 15 13 2 16 16 13 15 9 2 3 13 3 15 0 2
16 3 3 4 13 3 2 16 15 13 15 9 7 9 13 3 2
47 15 15 9 2 0 7 0 9 2 13 3 2 16 3 13 15 2 15 9 4 13 7 15 4 13 9 2 7 13 9 2 16 3 15 13 13 13 9 2 7 15 13 3 9 0 9 2
4 3 13 13 2
17 9 3 0 7 12 9 13 9 3 7 13 13 2 3 9 13 2
16 15 13 9 0 9 7 13 0 9 0 9 13 3 0 9 2
17 15 13 9 9 7 13 3 0 9 2 15 15 13 0 7 0 2
5 15 13 0 9 2
22 16 15 9 13 13 9 2 15 9 13 13 15 15 9 2 3 9 13 3 13 9 2
15 16 15 3 13 0 9 2 15 13 15 0 9 9 9 2
40 9 9 2 15 4 13 13 0 9 2 13 2 16 16 9 13 0 7 0 13 13 9 2 3 9 13 4 13 15 3 0 2 7 16 13 13 13 9 0 2
15 15 13 3 9 15 0 9 2 15 4 13 13 15 9 2
33 15 13 3 2 16 0 9 13 9 13 15 3 0 2 7 13 2 16 16 9 3 13 9 13 9 2 15 13 0 9 3 0 2
18 9 9 13 3 3 9 9 2 16 15 13 13 15 9 13 9 9 2
15 15 13 9 0 9 13 2 15 13 3 2 9 7 9 2
31 15 9 13 2 16 13 0 13 0 9 0 9 7 13 3 0 9 9 15 9 2 15 13 0 9 7 15 1 0 9 2
17 15 9 3 13 13 0 9 0 9 7 13 0 9 9 13 1 2
11 3 15 9 13 9 9 0 9 13 13 2
11 4 15 3 3 13 13 15 3 0 9 2
20 7 13 15 9 15 9 15 9 7 13 3 3 15 13 7 3 3 15 13 2
33 9 2 15 13 0 9 2 13 15 13 15 9 7 3 15 9 13 15 9 9 0 9 13 2 3 0 9 7 0 9 15 13 2
13 7 13 15 13 9 3 2 13 3 0 0 0 2
26 15 9 13 13 15 2 16 15 9 4 13 15 9 1 2 7 15 13 0 9 9 0 2 15 9 2
12 3 13 13 9 2 15 13 0 9 9 9 2
21 9 13 13 15 2 15 13 9 9 7 13 2 7 9 9 13 9 0 0 0 2
5 9 13 0 9 2
13 9 13 9 7 9 2 16 15 3 13 9 3 2
7 15 9 13 3 3 9 2
27 15 13 0 0 7 0 9 2 13 0 9 9 9 9 2 0 9 9 0 9 1 7 9 9 9 9 2
21 13 9 3 13 2 13 9 3 13 2 1 3 9 2 7 15 13 3 0 9 2
6 9 13 9 0 9 2
16 15 9 9 9 13 7 15 13 0 9 13 0 9 0 9 2
5 15 13 0 9 2
28 9 2 15 3 13 9 13 9 2 13 15 0 9 13 2 16 13 9 13 9 3 3 2 7 13 0 9 2
21 15 13 9 0 9 0 9 2 7 3 15 13 2 16 9 0 9 13 3 13 2
19 15 0 9 2 9 3 0 9 9 2 13 9 2 16 9 15 13 9 2
14 15 9 13 9 13 3 7 13 9 13 1 9 9 2
9 3 13 3 13 0 7 0 9 2
14 9 2 15 3 4 3 13 9 2 13 7 13 9 2
10 9 4 13 7 15 9 13 9 9 2
10 3 15 4 13 9 9 7 13 9 2
11 9 13 9 9 7 15 9 13 3 3 2
11 3 3 15 2 15 9 13 3 9 13 2
20 15 9 13 9 0 9 0 9 2 16 0 9 13 9 9 4 3 13 0 2
42 9 9 2 15 3 13 9 3 2 16 15 15 0 9 13 2 13 16 9 13 13 15 3 9 2 7 3 9 2 16 9 13 9 2 15 3 13 9 0 9 3 2
5 7 3 3 13 2
7 15 9 13 9 13 9 2
20 15 13 9 9 3 7 13 3 9 9 2 15 9 3 13 9 0 0 9 2
14 9 13 15 9 3 9 7 13 0 15 9 13 9 2
19 9 13 2 7 13 9 9 7 0 9 2 15 13 3 13 9 9 13 2
4 9 13 0 2
19 15 13 3 9 2 13 9 15 9 15 15 9 7 13 15 13 3 9 2
1 9
4 2 13 15 2
3 2 6 2
6 2 15 13 0 9 2
4 2 0 0 2
9 2 6 13 15 3 3 9 13 2
7 2 13 4 3 13 15 2
5 2 13 4 13 2
4 13 9 3 2
10 2 15 13 9 2 13 13 15 15 2
5 2 13 4 13 2
6 9 13 9 7 15 2
5 2 15 15 13 2
4 13 3 15 2
6 2 6 16 3 3 2
6 15 9 4 9 13 2
10 2 0 9 2 13 13 13 15 13 2
12 2 15 13 15 11 2 13 16 15 13 13 2
8 2 15 13 15 9 7 15 2
9 2 15 13 3 13 2 13 3 2
6 2 13 3 13 15 2
5 15 13 15 9 2
8 2 3 15 13 15 9 3 2
8 2 15 4 3 13 15 15 2
14 2 16 15 13 15 0 7 15 13 3 15 12 9 2
9 2 7 15 13 15 3 0 0 2
12 2 16 3 2 13 15 13 15 9 3 9 2
9 2 15 4 13 15 0 0 9 2
7 2 3 3 9 2 3 2
6 2 3 0 2 13 2
3 9 3 2
7 2 11 13 13 15 9 2
3 13 9 2
3 11 0 9
6 0 9 13 0 0 2
13 11 11 9 11 13 0 9 13 11 13 0 9 2
19 11 13 3 2 15 9 11 4 13 9 7 3 15 13 3 13 9 9 2
10 11 13 9 3 2 11 13 15 9 2
13 11 13 9 9 9 2 13 9 7 13 3 11 2
14 11 13 11 0 9 2 3 15 4 4 13 13 3 2
15 3 15 4 13 9 0 9 1 2 3 9 9 7 9 2
9 15 13 3 13 13 3 9 3 2
10 7 0 13 9 13 9 2 3 0 2
16 9 13 13 13 9 11 13 9 2 13 15 13 13 9 3 2
13 11 13 9 9 7 9 2 15 13 15 9 9 2
20 9 15 13 3 13 13 2 15 4 13 15 3 16 15 0 9 13 9 9 2
7 9 15 15 1 13 13 2
18 15 13 13 9 9 2 7 9 9 13 3 9 13 3 9 7 9 2
6 11 13 9 1 11 2
10 9 13 15 9 2 7 11 13 13 2
5 15 13 0 9 2
9 9 15 13 0 9 13 15 13 2
13 15 9 13 15 0 0 2 3 3 11 0 9 2
20 9 1 13 11 3 0 11 15 4 3 3 13 13 2 3 0 15 3 13 2
7 11 13 3 12 9 11 2
11 11 13 0 2 4 13 3 11 0 9 2
28 15 13 3 1 11 2 9 7 9 9 13 11 13 13 3 3 2 16 15 13 3 9 13 15 9 11 9 2
17 11 4 15 1 13 13 15 0 9 9 13 11 0 9 0 9 2
18 9 13 9 12 13 3 12 9 3 7 13 2 15 13 11 11 2 2
22 16 11 4 13 3 9 7 9 9 1 2 15 4 4 13 9 3 7 13 15 3 2
13 3 15 13 15 3 16 15 13 9 13 15 9 2
10 9 13 0 9 13 15 9 13 9 2
11 0 13 0 9 7 0 13 9 0 9 2
12 0 9 13 3 9 2 7 3 12 13 9 2
25 9 2 15 13 13 9 7 15 13 3 9 9 13 13 9 3 13 15 3 13 3 0 9 3 2
20 9 1 13 9 4 3 13 15 0 7 9 1 9 13 9 7 9 13 9 2
8 11 13 9 7 13 9 3 2
8 2 15 15 13 2 11 13 2
10 2 13 15 13 0 2 0 9 13 2
6 2 13 9 7 9 2
9 11 13 9 7 13 15 0 9 2
9 2 13 15 7 13 2 11 13 2
14 2 15 13 12 9 7 15 13 12 2 0 9 13 2
16 2 3 13 2 12 15 13 7 13 3 9 0 9 15 9 2
11 11 13 15 9 9 13 13 2 15 13 2
5 0 9 13 13 2
11 15 13 1 11 9 3 7 13 0 9 2
4 11 13 9 2
11 9 13 0 9 9 7 13 9 13 9 2
14 9 13 9 13 9 7 13 9 9 9 13 13 9 2
12 0 9 13 9 2 7 13 9 13 13 9 2
11 0 9 13 9 1 7 13 11 13 9 2
8 11 13 3 9 7 13 9 2
17 15 13 9 12 9 13 3 15 16 15 2 16 9 13 15 3 2
13 11 13 15 15 2 13 4 3 13 9 9 9 2
21 15 3 11 9 4 3 13 15 11 13 9 2 15 4 13 15 13 15 9 9 2
11 0 9 13 9 13 7 13 3 9 9 2
9 2 13 9 3 2 9 13 3 2
5 2 15 13 13 2
17 0 9 13 11 13 15 1 7 13 15 9 9 3 3 16 13 2
7 11 13 9 13 3 13 2
14 9 2 9 7 9 9 13 9 13 9 9 13 15 2
11 15 13 13 9 13 7 15 13 15 3 2
19 9 13 9 3 11 9 7 13 15 0 2 16 13 13 13 9 13 9 2
14 16 11 9 13 3 11 2 11 13 3 15 0 13 2
15 15 13 15 9 1 13 11 7 15 13 15 0 9 1 2
16 13 3 3 0 13 13 9 3 7 0 9 9 13 15 9 2
19 0 9 11 11 0 9 13 9 9 9 12 13 11 0 9 13 0 9 2
15 15 9 13 3 0 9 7 15 0 9 13 13 11 9 2
13 9 13 9 7 9 12 9 13 3 11 11 11 2
7 15 13 3 11 0 9 2
4 9 7 9 9
13 15 9 3 0 9 9 1 0 11 11 9 13 2
13 9 13 0 7 0 7 13 3 13 9 9 1 2
9 11 13 9 9 7 13 9 11 2
6 11 13 7 13 9 2
12 15 13 9 7 13 13 9 13 9 9 11 2
15 11 13 11 13 1 9 7 13 3 9 3 16 13 9 2
9 11 13 9 16 11 13 9 1 2
7 2 9 9 2 11 13 2
5 2 15 9 13 2
7 2 9 3 2 11 13 2
8 2 9 13 9 16 3 13 2
7 13 3 0 9 16 9 2
8 2 13 9 3 2 11 13 2
23 2 9 4 13 9 0 3 15 1 16 11 11 13 9 9 9 11 7 13 12 9 9 2
9 2 13 13 2 9 13 3 9 2
6 15 15 3 9 13 2
5 2 13 11 9 2
9 9 13 2 16 3 4 13 9 2
7 13 2 16 3 13 3 2
8 2 15 4 13 2 11 13 2
10 2 15 4 13 2 16 9 13 13 2
12 13 3 3 0 9 2 16 13 3 9 9 2
7 9 13 9 9 13 9 2
11 2 13 9 2 16 9 11 13 0 9 2
12 13 3 3 9 9 13 4 13 3 3 3 2
10 2 9 1 13 3 13 2 11 13 2
14 2 9 13 3 2 3 9 9 8 13 3 13 9 2
6 13 15 13 3 13 2
7 9 4 13 7 13 15 2
10 2 0 9 13 9 3 2 11 13 2
6 2 3 11 3 13 2
10 11 13 9 7 9 3 4 13 9 2
4 2 13 9 2
7 15 13 11 2 0 9 2
13 3 16 11 13 13 2 9 13 0 7 0 9 2
6 2 9 2 11 13 2
5 2 3 13 3 2
9 11 13 9 2 15 13 0 9 2
7 2 3 3 2 11 13 2
11 2 13 15 15 0 9 13 2 11 13 2
12 2 13 15 15 9 13 13 2 13 13 15 2
15 11 7 11 13 9 7 15 1 13 9 2 15 11 13 2
7 2 3 3 2 11 13 2
6 2 13 3 3 3 2
6 11 13 3 0 9 2
7 9 9 4 13 0 0 2
11 11 13 9 2 16 9 4 13 3 3 2
10 9 1 13 12 9 2 15 13 3 2
10 2 13 3 13 9 2 0 9 13 2
16 2 13 13 2 13 2 16 9 4 13 9 1 2 11 13 2
10 2 9 13 13 2 15 13 9 1 2
10 2 15 15 13 7 3 13 3 9 2
9 2 15 13 11 2 0 9 13 2
6 2 15 9 13 11 2
7 13 13 15 13 3 9 2
8 13 13 2 13 15 13 9 2
11 2 15 3 9 13 7 3 2 11 13 2
14 2 15 9 13 13 16 9 9 2 9 7 9 9 2
11 2 15 3 13 2 13 9 2 11 13 2
15 2 15 13 13 2 13 9 9 9 7 13 9 9 9 2
8 7 13 9 9 13 15 9 2
13 2 13 3 13 2 16 13 3 3 2 11 13 2
6 2 15 15 15 13 2
6 11 7 11 13 3 2
5 9 9 13 9 2
9 11 7 11 13 15 9 7 13 2
8 11 4 13 9 7 9 9 2
8 11 13 9 1 7 13 9 2
10 15 13 9 7 13 15 9 0 9 2
6 3 15 13 9 9 2
1 9
12 13 3 3 0 9 2 13 15 9 3 13 2
16 9 13 0 16 15 9 13 9 1 2 15 1 13 3 9 2
10 15 9 15 13 9 7 9 1 9 2
16 15 13 15 3 13 9 2 15 13 15 13 3 9 3 3 2
6 9 1 15 13 9 2
11 13 0 9 0 0 7 13 15 1 9 2
13 9 15 13 0 2 9 16 13 0 9 0 9 2
19 13 2 16 16 9 13 9 2 13 15 15 9 7 15 13 0 9 15 2
11 3 15 13 15 9 9 7 9 9 3 2
9 9 13 0 7 0 9 0 9 2
19 9 2 9 7 15 9 13 0 9 3 0 2 9 1 15 3 13 13 2
7 15 13 15 16 13 13 2
15 9 3 2 3 15 9 1 16 13 3 13 9 9 0 2
17 13 3 13 9 2 3 0 15 4 13 2 13 3 13 9 3 2
13 15 9 2 15 4 3 13 0 2 13 15 0 2
12 15 13 15 9 2 13 3 16 9 13 9 2
6 3 9 1 15 13 2
12 9 13 3 3 9 2 3 0 7 9 13 2
10 3 13 0 2 0 7 13 9 9 2
8 13 15 3 3 3 13 9 2
5 13 15 13 9 2
2 9 9
5 13 3 0 9 2
13 15 13 3 3 9 9 2 3 15 13 15 9 2
12 16 13 15 1 2 15 13 9 9 3 15 2
19 3 13 3 13 1 0 9 2 1 0 9 2 15 3 9 0 9 13 2
14 13 13 3 3 2 7 13 2 16 15 13 3 0 2
25 16 15 13 2 13 13 9 2 7 16 15 13 13 15 2 13 13 3 13 13 15 3 16 3 2
21 15 13 3 3 13 15 9 9 2 13 3 2 7 15 13 13 3 15 0 9 2
11 13 13 3 13 9 2 13 13 3 15 2
3 13 15 1
18 13 4 13 3 2 13 2 13 3 3 16 13 2 3 3 16 13 2
15 13 13 16 15 13 15 9 2 3 2 13 15 3 13 2
12 15 13 13 3 2 13 2 13 2 3 3 2
5 9 3 15 9 2
11 2 3 2 3 2 13 15 13 15 13 2
6 2 7 15 13 9 2
7 2 15 13 13 3 9 2
14 13 3 15 0 9 1 2 15 15 4 3 13 9 2
24 13 9 2 13 9 3 2 13 9 3 7 13 15 9 2 15 9 13 13 12 9 9 1 2
13 13 15 3 9 0 9 2 13 3 13 3 9 2
7 3 13 3 13 9 9 2
5 2 15 13 11 2
4 11 13 9 2
31 11 13 15 2 15 13 3 9 9 2 15 2 15 13 3 9 9 7 15 15 13 3 2 13 2 16 15 15 13 2 2
18 16 13 2 16 9 13 0 2 15 13 7 9 7 9 2 9 1 2
18 11 13 9 2 15 13 15 3 0 2 15 3 13 13 3 13 9 2
24 2 13 16 9 2 2 9 13 2 13 13 13 15 7 11 1 2 2 15 16 13 9 2 2
11 13 0 2 16 11 4 13 13 15 3 2
16 3 13 15 9 16 9 2 3 16 13 11 1 9 1 9 2
25 13 9 0 9 2 9 13 0 7 15 15 13 0 0 9 7 9 2 15 13 0 13 9 9 2
13 13 3 3 13 0 9 2 9 13 3 0 9 2
14 9 13 3 15 13 0 9 16 11 13 7 15 13 2
14 9 13 2 13 9 2 7 13 13 9 11 0 1 2
12 4 3 13 15 15 2 13 15 3 11 1 2
15 3 13 15 4 13 2 16 13 9 15 9 9 13 3 2
14 13 15 3 2 3 0 7 0 9 13 3 9 9 2
7 2 6 15 13 15 9 2
11 2 15 13 2 3 15 13 15 9 9 2
11 2 6 15 13 15 15 2 13 15 0 2
5 2 3 15 2 2
22 3 15 13 2 3 3 16 9 4 13 3 7 9 9 13 16 15 4 13 0 9 2
15 3 15 13 2 13 9 7 13 9 2 13 13 15 15 2
9 15 13 9 13 9 2 15 13 2
8 13 2 13 3 3 16 13 2
12 13 3 3 2 13 4 3 3 13 3 9 2
21 16 13 3 13 2 13 9 2 13 9 3 7 13 2 16 15 13 3 0 9 2
18 3 13 0 9 2 15 13 11 2 7 9 1 13 15 13 15 0 2
12 2 13 15 15 2 2 11 13 7 13 9 2
25 13 15 9 7 13 2 3 11 13 9 2 13 15 13 9 2 13 15 9 3 7 13 9 3 2
9 15 13 9 7 13 15 3 9 2
17 0 9 15 13 3 13 2 16 11 13 9 7 0 9 9 9 2
16 13 11 13 3 13 9 2 7 13 3 15 13 9 9 1 2
16 15 13 3 7 13 3 11 13 13 2 15 13 7 13 15 2
6 15 13 9 0 9 2
11 13 15 9 2 13 15 3 7 13 3 2
26 9 9 13 15 9 2 15 15 13 9 2 15 9 2 15 13 2 2 0 9 2 9 7 9 2 2
4 13 3 13 9
26 13 3 9 12 7 12 2 16 13 15 0 9 2 7 3 15 2 15 13 9 3 9 9 13 9 2
21 15 13 15 2 15 13 9 13 12 0 9 2 13 9 9 16 15 3 13 9 2
16 3 13 15 1 2 13 2 15 13 2 7 15 13 11 11 2
22 13 15 13 3 9 2 0 9 15 15 9 7 15 13 3 0 9 2 13 15 3 2
24 13 7 13 15 9 15 1 7 15 13 7 13 9 9 16 9 3 13 7 15 13 3 13 2
34 13 15 9 7 13 9 0 9 2 13 2 16 3 13 15 9 2 7 3 13 15 9 16 9 15 13 15 15 7 13 9 9 9 2
17 15 13 3 9 1 2 16 13 15 15 3 13 2 13 3 9 2
13 3 13 15 9 3 2 7 3 0 9 13 13 2
24 13 3 3 13 2 13 3 9 2 16 15 13 0 2 15 9 15 4 4 13 15 9 11 2
28 15 0 9 2 3 9 12 7 12 2 15 13 15 9 7 13 2 13 15 3 9 7 13 3 15 13 15 2
29 15 3 3 13 2 6 2 16 13 9 7 3 13 9 2 16 13 13 15 13 0 2 13 2 3 15 9 13 2
18 13 4 13 9 2 7 13 15 3 9 2 7 15 13 13 15 9 2
15 2 15 16 13 3 9 2 2 13 15 15 1 3 13 2
2 3 2
12 3 3 15 2 16 15 9 13 0 1 15 2
12 3 13 15 2 13 9 9 7 3 15 13 2
19 3 3 3 13 15 2 7 3 9 9 13 3 2 0 9 15 0 1 2
24 13 0 9 2 0 9 2 9 7 9 1 2 11 9 9 7 9 9 2 9 7 12 9 2
35 15 9 9 2 9 0 9 13 9 15 9 2 15 4 13 9 15 2 13 13 9 7 9 3 2 7 9 9 4 13 15 9 9 9 2
9 13 16 13 15 3 4 13 13 2
18 7 3 13 9 12 7 12 2 13 9 13 7 13 15 9 9 1 2
16 13 0 2 9 13 9 2 7 1 9 9 13 15 1 9 2
8 2 6 2 15 13 2 13 3
8 15 13 15 9 3 2 13 3
8 2 6 2 11 11 2 3 2
19 2 6 3 2 0 9 2 13 3 2 13 16 13 0 9 2 13 13 2
19 3 3 2 7 13 3 13 15 7 9 1 2 15 13 13 3 2 13 3
13 2 6 6 2 15 13 3 7 13 13 9 3 2
12 2 7 13 11 7 11 1 2 15 13 11 2
9 4 13 0 3 2 13 3 3 2
27 9 13 2 9 13 3 15 13 3 11 1 2 13 16 9 13 3 2 7 13 11 11 11 11 11 13 2
2 9 9
13 13 9 3 0 9 7 9 13 9 3 13 9 2
12 3 9 13 15 9 2 3 13 15 13 3 2
32 9 0 9 13 3 9 2 13 15 13 15 4 13 2 16 15 9 9 4 9 1 13 12 9 3 2 2 13 15 3 2 2
15 3 13 9 9 1 2 16 9 13 9 0 9 9 9 2
20 9 13 13 9 9 2 13 9 9 2 2 7 13 9 9 16 13 9 9 2
9 3 9 13 2 13 3 3 9 2
30 15 9 2 15 13 9 9 2 13 9 9 7 13 9 9 9 9 2 9 2 15 1 0 9 13 7 9 9 13 2
13 13 9 9 9 1 2 16 9 15 1 13 9 2
22 9 13 13 15 9 13 15 2 7 3 9 13 13 9 9 0 9 9 9 15 9 2
9 3 9 4 13 2 4 3 13 2
19 13 9 15 9 2 13 9 1 15 1 13 9 1 13 2 13 9 13 2
20 13 15 9 13 2 9 2 16 15 4 2 3 4 15 3 13 9 0 9 2
30 0 9 9 13 9 9 13 2 3 16 15 4 3 9 13 2 7 13 3 9 3 13 9 2 13 15 15 4 13 2
26 15 9 9 13 0 2 7 15 0 9 4 3 13 0 7 0 9 2 15 9 9 4 13 15 3 2
20 3 9 13 9 9 9 2 15 9 13 9 3 3 2 2 13 15 3 2 2
16 13 9 13 3 9 2 16 9 13 3 13 9 3 9 1 2
6 13 15 3 15 13 2
24 13 15 9 3 13 9 13 9 9 9 13 15 9 7 9 2 4 9 13 15 9 15 9 2
19 9 13 9 9 2 13 2 13 9 15 2 2 7 13 15 3 9 9 2
32 3 9 13 9 9 2 9 2 15 13 9 9 2 13 3 9 7 13 3 13 9 2 9 2 15 9 4 13 12 9 3 2
2 9 9
21 13 9 7 9 2 13 3 16 13 9 13 9 13 9 7 9 13 9 15 0 2
17 13 9 9 0 9 2 7 13 13 15 3 4 13 15 13 15 2
30 9 13 9 1 7 13 9 13 9 1 16 13 0 11 9 1 0 9 9 2 3 15 13 9 7 13 9 3 9 2
22 13 11 9 7 13 11 9 1 2 9 9 13 7 9 3 13 2 13 15 3 2 2
16 13 9 9 9 16 13 9 9 9 2 13 13 15 15 15 2
16 9 9 13 9 9 9 7 13 2 2 15 3 4 13 2 2
31 13 7 13 9 9 9 13 9 9 0 9 1 2 9 2 15 3 13 9 9 2 7 9 2 15 13 3 13 3 2 2
10 13 9 9 2 9 7 13 9 1 2
12 13 9 2 7 13 2 3 9 13 0 9 2
33 3 13 15 9 15 13 2 13 15 0 0 9 2 7 13 13 13 9 2 15 3 13 15 13 2 3 3 13 13 15 3 2 2
2 7 2
21 13 3 3 13 9 15 13 15 15 9 2 13 9 7 9 2 3 15 9 1 2
22 15 13 13 15 2 15 9 13 0 0 16 15 3 13 2 7 15 13 15 3 3 2
23 3 3 13 9 1 7 13 9 15 13 3 9 2 0 15 13 15 0 9 3 15 9 2
19 15 13 15 9 16 13 13 13 9 9 2 13 3 3 13 15 4 13 2
11 9 9 13 9 2 9 13 2 3 15 2
21 13 9 3 9 13 2 4 9 9 7 9 9 13 2 13 9 9 9 3 13 2
32 16 0 11 13 0 2 0 9 13 9 2 13 2 0 9 2 13 9 13 9 9 1 2 13 15 9 15 9 3 13 2 2
19 3 13 9 9 13 9 2 3 15 13 9 2 3 15 13 3 9 9 2
4 3 9 13 2
6 2 3 9 13 2 2
7 2 6 2 3 12 2 2
5 2 15 13 2 2
8 2 6 2 15 13 9 9 2
7 7 15 13 13 15 2 2
3 2 6 2
7 6 3 15 3 13 2 2
4 2 15 3 2
5 15 13 9 9 2
6 7 3 15 13 3 2
6 13 3 15 9 2 2
10 2 7 13 15 3 13 15 3 2 2
4 2 13 15 2
3 13 3 2
23 0 9 3 9 9 13 16 3 2 7 9 3 1 9 13 16 15 13 3 3 1 12 2
15 16 15 13 9 9 2 3 15 13 3 3 3 1 12 2
13 15 13 15 9 13 2 7 15 13 3 15 3 2
3 3 2 2
8 2 16 13 15 13 3 3 2
6 15 9 3 13 2 2
4 2 3 3 2
5 15 13 3 12 2
17 16 15 13 13 9 13 2 3 15 13 3 3 3 16 15 13 2
11 13 15 15 13 2 3 13 15 15 2 2
3 2 6 2
21 7 16 9 13 3 3 9 2 7 15 13 9 16 15 13 15 3 16 15 13 2
8 13 3 9 7 15 13 3 2
5 15 15 13 2 2
6 2 4 13 3 9 2
6 15 13 3 3 2 2
6 7 16 13 9 2 2
9 2 15 13 0 9 16 15 2 2
13 2 3 2 15 13 0 9 7 15 13 0 9 2
12 15 13 0 9 16 15 13 3 0 9 2 2
8 2 15 9 13 6 3 0 2
3 13 13 2
22 3 15 13 3 0 9 2 7 16 15 13 0 9 16 15 2 3 15 15 15 13 2
21 15 3 13 13 15 9 2 7 16 15 4 15 13 2 3 15 13 12 9 2 2
6 2 15 13 13 2 2
4 2 13 3 2
7 13 3 3 15 9 13 2
6 7 13 15 4 13 2
11 15 9 9 13 6 0 9 2 7 9 2
13 4 13 3 13 15 3 16 4 13 15 13 9 2
7 6 15 13 3 0 9 2
8 15 13 15 3 16 15 13 2
8 7 15 13 3 15 15 13 2
5 13 15 4 13 2
10 6 2 15 3 13 16 9 13 0 2
5 15 13 15 3 2
14 15 4 3 3 13 13 15 15 9 2 13 3 9 2
12 16 9 13 13 15 2 3 15 13 3 9 2
7 13 15 13 15 9 2 2
3 2 6 2
12 7 15 15 9 4 13 3 3 12 3 2 2
7 2 6 2 13 15 2 2
12 2 3 15 3 13 15 15 9 16 13 15 2
9 16 15 3 13 3 15 3 2 2
8 2 6 15 15 9 3 13 2
4 9 13 0 2
9 4 13 16 15 13 16 9 13 2
12 4 13 0 13 13 15 15 13 13 9 2 2
3 2 6 2
6 7 13 3 13 2 2
6 2 7 13 15 13 2
4 15 13 3 2
5 15 13 9 2 2
2 0 9
3 15 13 2
14 15 9 3 2 9 13 9 9 2 13 3 13 9 2
13 15 9 3 2 9 13 9 3 13 0 9 9 2
11 15 9 13 3 9 3 13 9 13 9 2
13 3 15 13 13 15 3 2 7 3 9 15 13 2
13 0 9 13 9 7 15 13 0 9 13 9 1 2
13 0 9 13 9 15 13 7 13 3 9 9 9 2
3 13 9 2
13 15 13 13 3 2 7 3 0 9 13 0 9 2
10 15 13 0 9 0 7 13 9 9 2
13 15 13 3 13 2 16 9 0 9 1 13 0 2
12 9 1 2 3 3 2 13 3 3 9 3 2
6 9 13 15 3 9 2
4 15 13 9 2
9 13 0 9 7 13 13 0 9 2
4 0 9 13 2
11 9 13 9 2 13 3 0 13 9 9 2
10 15 13 15 9 1 2 13 3 3 2
7 13 9 0 0 9 1 2
12 9 9 13 9 2 7 3 13 3 0 9 2
5 15 9 13 3 2
5 9 13 3 13 2
11 9 13 9 13 9 1 7 13 15 1 2
4 15 15 13 2
3 13 3 9
7 11 9 4 13 3 9 2
27 15 4 3 13 9 2 13 3 9 1 9 2 7 3 13 0 9 3 3 9 2 16 15 4 3 13 2
15 15 13 3 13 9 13 15 2 7 3 13 9 0 9 2
7 0 9 13 13 0 13 2
16 3 11 0 9 4 13 15 3 3 2 16 9 9 13 0 2
21 9 9 4 9 9 13 2 7 3 15 15 2 13 11 9 13 15 9 9 9 2
9 15 4 13 9 3 9 1 12 2
11 9 4 13 12 2 7 9 4 13 12 2
8 13 3 9 2 16 9 13 2
12 0 9 13 9 2 7 9 4 13 11 9 2
16 3 9 9 4 13 2 16 15 4 4 13 3 3 12 9 2
13 9 4 9 9 13 15 9 2 7 13 15 9 2
20 3 15 13 3 9 0 9 2 15 1 13 7 9 2 9 2 9 7 9 2
8 9 13 15 2 9 13 9 2
11 15 1 13 3 3 15 13 0 9 1 2
12 15 0 9 13 9 2 15 13 3 9 9 2
24 9 13 3 15 12 9 9 13 2 13 15 3 13 9 9 1 2 3 15 13 13 9 3 2
13 15 13 3 15 0 9 3 2 15 13 15 9 2
25 15 13 9 2 9 9 7 0 9 13 15 9 9 1 2 16 13 15 9 13 3 3 9 13 2
4 13 3 13 2
14 3 16 11 13 13 9 2 15 1 13 9 3 0 2
15 15 9 13 0 13 2 16 9 13 3 13 0 9 1 2
25 3 9 13 0 0 2 0 9 13 9 2 9 2 7 9 15 9 3 12 9 3 16 9 13 2
12 9 13 9 13 9 7 9 15 9 16 9 2
16 11 13 9 2 7 13 15 3 3 13 0 9 9 0 9 2
16 3 3 9 13 15 9 0 9 2 0 9 15 3 9 13 2
25 11 13 13 13 15 9 9 15 9 13 2 7 13 4 13 3 2 16 9 13 3 3 0 0 2
27 9 13 9 9 2 13 15 9 9 16 13 2 13 11 9 7 13 13 9 3 3 2 16 9 9 13 2
10 11 13 9 13 9 9 13 15 13 2
26 15 0 9 1 9 9 13 13 0 9 2 15 3 13 15 13 9 9 2 0 13 4 13 13 9 2
15 3 9 13 13 9 2 13 3 13 13 15 16 0 9 2
15 15 13 9 9 7 13 3 9 9 2 13 3 1 9 2
19 9 13 15 15 9 13 11 13 3 9 13 9 2 7 3 13 13 9 2
11 3 3 3 16 9 4 13 2 15 13 2
8 3 9 7 3 3 9 9 2
20 11 9 13 3 0 9 2 7 13 13 13 13 9 9 7 13 3 0 9 2
21 15 9 9 2 15 13 0 9 9 1 2 11 13 9 15 3 3 13 1 9 2
8 15 13 3 9 9 3 9 2
10 3 9 13 7 9 13 15 13 9 2
15 16 15 13 2 3 13 9 4 13 2 13 9 0 9 2
16 9 1 9 13 9 13 0 9 2 15 13 3 9 9 9 2
14 3 3 13 0 6 2 15 4 13 9 15 13 9 2
22 9 13 0 9 13 9 9 0 9 3 3 13 9 2 13 0 9 15 13 0 9 2
8 9 13 3 9 7 13 3 2
19 11 13 13 3 3 2 16 13 3 13 9 9 7 13 3 13 13 9 2
14 13 9 13 9 9 2 15 13 7 13 13 15 13 2
11 11 9 13 4 13 15 15 4 3 13 2
12 9 4 13 3 0 2 7 3 13 9 9 2
2 3 2
8 15 13 1 9 3 0 9 2
16 15 0 9 9 2 13 15 13 9 9 7 13 15 3 9 2
9 9 2 6 2 3 15 13 9 2
13 3 15 9 13 9 13 0 7 13 0 9 9 2
11 3 0 2 16 11 13 9 3 13 3 2
13 3 15 13 13 2 13 9 2 9 7 9 3 2
11 0 9 3 9 3 2 7 9 3 13 2
7 15 13 3 13 0 9 2
7 15 13 15 3 0 9 2
10 3 13 3 0 2 0 9 13 9 2
4 9 7 9 2
6 15 13 3 0 9 2
5 15 3 3 0 2
9 15 15 13 9 9 2 3 11 2
13 15 3 13 15 15 13 3 15 15 16 0 0 2
21 2 7 15 9 13 9 15 13 13 3 2 2 13 0 7 0 9 15 9 1 2
8 2 15 13 3 3 15 9 2
16 13 0 7 13 15 3 13 13 9 9 1 2 2 9 13 2
7 11 13 13 13 3 15 2
6 3 9 13 3 3 2
6 2 15 13 0 9 2
12 7 13 13 3 7 3 2 16 9 13 3 2
6 3 3 13 3 2 2
19 3 16 11 13 2 15 13 9 13 0 9 2 15 3 13 15 0 9 2
20 15 13 15 9 13 9 12 9 15 13 0 9 13 9 2 7 3 15 13 2
5 13 15 15 13 2
8 7 15 13 15 3 13 9 2
15 11 13 9 9 11 11 9 9 9 13 11 0 9 9 2
15 9 13 13 9 3 2 16 9 4 9 13 7 13 9 2
3 15 4 13
22 16 3 9 7 15 4 13 16 7 15 9 3 16 9 9 3 13 15 15 9 9 2
4 11 13 11 2
8 3 15 13 3 13 3 9 2
5 0 9 15 13 2
10 3 0 9 13 3 13 13 13 9 2
16 3 3 15 3 13 3 3 2 16 15 4 3 9 13 3 2
6 15 13 13 16 15 13
10 11 13 0 9 7 11 9 0 9 2
6 9 13 3 3 13 2
3 13 15 2
6 3 0 13 0 9 2
7 15 13 15 9 13 9 2
13 11 11 13 9 13 13 2 16 9 4 13 3 2
4 13 15 13 2
9 11 13 3 15 9 2 11 12 2
7 9 13 7 9 13 3 2
2 13 13
5 15 13 3 9 2
3 3 13 2
15 0 9 13 0 2 0 9 2 15 9 13 3 12 9 2
2 0 9
12 9 13 9 9 9 7 3 13 15 0 9 2
3 13 13 3
11 3 15 4 13 3 3 3 12 9 9 2
7 9 4 9 13 13 3 2
7 15 0 13 16 13 9 2
7 3 4 3 13 15 9 2
9 3 9 7 9 9 13 13 15 2
3 3 7 3
9 9 9 13 13 12 9 9 13 2
17 11 13 16 9 2 15 13 13 13 12 9 2 13 13 13 9 2
6 13 13 3 9 11 2
10 9 4 13 9 2 9 13 3 3 2
9 15 15 15 13 2 16 13 9 2
5 3 0 13 9 2
11 9 13 13 0 2 16 13 13 3 9 2
7 13 3 2 16 13 9 2
8 3 0 9 13 3 3 3 2
3 9 13 2
15 15 9 1 9 9 9 13 13 11 7 11 11 9 11 2
6 9 0 9 13 9 2
6 9 9 4 3 13 2
11 11 13 9 3 7 13 15 3 3 3 2
13 9 11 11 7 11 11 13 9 3 11 11 1 2
7 16 13 15 3 9 13 2
13 16 15 4 15 9 13 2 15 9 4 13 13 2
10 11 9 11 11 13 9 9 0 9 2
5 0 11 3 13 9
4 13 9 9 2
10 1 9 9 13 9 2 13 15 0 9
10 9 13 0 2 0 7 9 0 0 2
5 9 13 3 0 2
11 9 13 15 9 2 7 9 4 13 9 2
4 15 13 15 13
8 11 13 9 7 9 13 9 2
8 9 13 9 13 0 0 9 2
2 13 3
2 9 13
9 9 13 11 13 3 12 12 9 2
6 6 6 13 15 3 2
4 15 13 9 2
2 0 9
11 15 13 11 9 7 9 0 12 9 9 2
10 11 13 12 9 9 0 9 9 9 2
8 15 13 0 2 16 9 13 2
7 9 15 9 7 9 15 2
11 15 13 0 7 9 7 0 9 1 0 2
19 15 7 9 13 15 9 1 3 3 3 9 2 13 9 9 11 2 12 2
23 7 16 12 9 13 3 3 13 9 2 15 15 7 15 15 9 2 3 15 13 15 9 2
7 15 9 13 13 13 9 2
17 11 11 13 15 9 9 2 16 15 9 4 13 3 15 13 9 2
12 9 1 11 4 13 3 0 9 7 9 13 2
5 9 13 3 0 2
12 11 4 13 3 13 7 13 7 0 7 15 2
10 9 4 13 15 9 9 3 12 9 2
6 15 13 13 3 0 2
8 3 11 0 2 0 2 9 2
13 9 9 13 9 9 7 13 9 2 15 13 3 2
42 13 15 13 13 15 16 15 13 12 9 9 16 15 13 15 0 9 13 13 16 15 2 3 15 13 15 7 6 7 3 13 3 11 2 7 15 11 7 11 13 16 2
5 15 13 15 0 2
8 15 13 15 13 13 15 9 2
5 15 15 11 13 2
5 13 13 12 3 2
14 9 2 15 15 4 4 9 13 2 13 13 13 9 2
13 13 0 9 0 9 13 2 7 3 15 15 13 2
11 3 4 13 3 0 9 16 2 16 16 2
5 0 9 3 13 2
17 11 11 9 1 13 3 9 15 2 15 13 11 9 7 15 9 2
9 4 13 12 9 13 9 9 13 2
8 13 11 15 15 4 13 15 2
10 9 13 9 13 15 3 3 15 9 2
7 15 13 3 0 16 13 2
10 15 13 3 2 16 4 13 15 0 2
6 13 9 3 12 9 2
7 11 13 9 0 11 9 2
9 11 11 13 9 9 9 0 0 2
18 15 13 11 9 3 9 2 16 13 2 3 9 13 13 3 9 1 2
4 9 15 9 2
8 11 13 15 9 12 11 9 2
11 9 13 2 16 13 15 13 3 12 9 2
2 9 9
11 9 1 13 3 4 13 0 9 7 9 2
12 15 13 0 9 2 13 15 13 3 12 9 2
7 15 13 0 16 15 13 2
14 15 1 13 13 15 9 2 16 9 13 15 0 9 2
11 9 13 2 3 12 0 9 13 13 9 2
9 9 9 13 11 11 7 11 11 2
2 13 13
4 9 13 0 2
3 13 3 2
10 15 13 9 2 15 13 9 7 9 2
4 15 13 13 2
5 15 13 13 15 9
8 3 9 13 7 13 0 9 2
9 3 3 13 16 11 4 13 9 2
5 13 9 9 9 2
10 13 0 2 0 9 0 9 9 1 2
9 9 13 9 9 13 15 3 9 2
6 3 15 9 4 13 2
19 11 13 9 11 2 7 13 3 3 13 11 2 7 9 4 13 0 9 2
18 9 9 7 3 3 13 9 1 11 13 3 9 7 9 7 3 9 2
6 9 11 4 13 9 2
2 3 13
24 15 9 9 9 9 3 3 7 11 13 4 3 13 3 15 13 3 7 13 16 13 15 13 2
10 11 9 9 9 13 11 11 9 11 2
5 9 13 9 1 2
13 0 9 13 15 2 13 13 0 9 0 7 0 2
5 9 13 9 13 2
17 9 9 13 9 13 9 9 3 1 9 7 15 13 12 9 9 2
11 13 9 13 12 9 2 15 13 3 12 2
13 9 13 9 9 13 9 1 3 13 3 9 9 2
6 9 3 13 13 9 2
9 9 3 13 13 11 7 11 3 2
5 2 13 15 9 2
8 13 9 3 3 4 4 13 2
10 0 0 9 9 1 13 12 9 1 2
16 11 9 13 0 9 2 15 3 13 0 9 2 15 9 13 2
4 15 15 13 2
6 11 13 0 0 9 2
16 9 9 13 3 9 2 15 13 11 11 9 11 11 9 9 2
9 9 1 13 0 9 0 9 1 2
7 0 9 11 13 9 11 2
28 13 9 3 15 9 13 9 0 9 2 16 13 9 13 3 3 9 9 7 15 2 16 15 9 11 13 9 2
4 13 3 3 2
17 15 15 13 2 16 9 13 3 0 13 13 3 0 2 0 9 2
13 3 15 13 13 9 2 15 13 9 15 13 9 2
8 4 13 0 9 7 0 9 2
6 11 9 13 9 11 2
8 3 13 9 13 2 13 9 2
18 0 2 2 0 2 0 2 0 2 7 0 9 13 9 9 3 13 2
2 9 9
6 15 9 15 9 13 2
11 6 3 0 9 3 15 13 12 0 0 9
20 13 3 0 2 16 9 3 13 0 9 15 2 15 15 9 3 13 13 9 2
10 15 13 2 16 15 13 11 0 9 2
6 9 15 9 2 13 2
8 9 13 15 0 9 7 0 9
4 15 13 3 2
8 9 15 4 13 13 2 3 2
4 9 0 0 9
6 9 13 0 0 9 2
3 9 13 0
11 9 13 0 3 13 7 13 15 3 15 2
7 15 9 13 9 9 9 2
12 9 13 3 3 2 15 9 13 9 7 9 2
5 15 9 13 9 2
7 15 13 3 11 9 15 2
6 9 13 13 11 9 2
6 15 13 9 9 12 2
12 11 11 11 13 0 9 0 3 3 9 9 2
9 9 9 13 3 3 0 13 9 2
7 13 3 9 9 15 3 2
4 13 13 3 2
13 9 9 13 12 1 13 13 9 2 9 7 9 2
8 13 13 2 15 15 4 13 2
6 9 13 9 3 3 2
7 11 9 13 12 12 9 2
10 11 4 13 9 7 15 3 9 3 2
10 16 15 13 13 2 15 15 3 13 2
4 15 13 4 13
5 13 3 9 15 13
7 9 13 9 12 9 3 2
14 15 13 13 2 7 3 2 15 13 2 16 15 13 2
4 13 15 13 9
4 11 3 11 9
4 15 9 13 15
4 15 13 9 2
5 9 13 3 9 2
10 13 15 13 9 7 13 9 9 9 2
6 11 13 3 9 9 2
9 9 13 9 13 9 11 11 11 2
15 13 15 4 15 15 13 2 4 15 15 13 2 0 9 2
9 11 9 13 9 11 0 9 9 2
4 9 13 3 2
6 11 13 3 13 3 2
17 4 13 9 13 9 3 13 2 16 3 4 13 9 2 13 2 2
12 9 4 13 9 2 16 9 9 4 13 3 2
4 13 15 9 2
11 9 9 13 9 2 15 13 13 0 9 2
3 13 3 9
5 13 3 3 9 2
10 15 9 9 3 15 13 15 3 9 2
2 15 9
15 3 9 4 13 9 13 9 12 9 0 9 0 9 1 2
6 15 13 13 15 3 2
4 0 0 9 2
8 4 15 9 1 13 15 9 2
3 13 3 2
3 13 9 1
9 13 9 2 9 7 9 0 9 2
14 7 15 13 15 7 15 15 13 15 0 13 9 9 2
3 3 13 2
9 0 9 13 3 13 15 9 13 2
3 13 12 3
15 7 3 9 13 9 2 16 13 3 11 2 3 3 11 2
15 3 3 9 13 13 9 16 3 3 13 9 13 0 9 2
9 3 9 13 9 3 0 12 9 2
4 13 15 3 2
9 3 3 3 15 1 2 11 13 2
2 13 13
8 9 13 13 15 15 15 15 2
20 15 13 9 15 0 9 2 15 4 13 2 16 15 9 9 0 9 13 0 2
8 9 13 3 0 0 13 9 2
11 3 13 0 9 13 2 9 13 9 0 2
4 3 9 13 2
5 11 13 12 9 2
11 13 15 2 16 9 4 13 3 3 3 2
4 15 13 3 2
7 13 15 3 13 3 15 2
2 15 9
8 15 13 3 3 7 13 9 2
3 12 9 13
10 7 15 13 3 0 16 15 13 9 2
15 15 13 3 0 16 15 13 3 13 2 3 13 3 13 2
13 11 9 13 3 3 0 9 16 3 11 9 9 2
12 7 13 13 13 9 3 2 16 15 13 15 2
7 9 13 13 13 9 3 2
22 3 15 13 9 13 13 0 0 9 2 16 0 9 9 7 9 9 4 13 0 9 2
3 13 0 2
6 15 15 4 13 3 2
4 9 7 0 9
12 13 15 3 3 4 13 15 9 16 15 13 2
11 3 4 13 9 0 9 2 15 9 1 2
9 9 9 13 3 15 16 9 9 2
4 11 13 13 2
5 13 9 7 13 15
11 9 13 15 2 13 9 11 7 15 9 2
6 9 4 13 1 9 2
15 16 0 9 9 13 13 2 15 13 15 3 9 9 9 2
3 9 7 9
13 9 13 3 2 15 13 15 9 2 16 11 13 2
8 13 0 2 16 13 3 9 2
8 11 13 11 0 7 0 9 2
5 9 4 13 0 2
14 11 11 1 11 4 4 3 13 13 9 3 0 9 2
4 9 13 11 2
8 3 3 3 6 3 3 13 2
17 15 9 13 9 9 2 15 15 4 13 9 1 3 0 2 9 2
11 0 9 13 13 9 3 0 9 16 0 2
5 3 15 13 13 2
6 11 4 13 13 9 2
7 0 9 1 9 9 13 2
4 15 15 13 2
2 15 9
10 11 13 9 1 3 15 9 0 9 2
11 3 13 9 7 9 13 3 0 9 9 2
3 9 13 9
8 13 3 3 2 16 3 13 2
4 15 13 9 2
12 15 9 16 13 15 13 9 2 13 9 3 2
9 16 3 13 13 2 4 13 9 2
13 4 13 15 15 9 2 11 13 13 16 9 4 2
4 16 13 9 2
2 9 9
4 9 13 15 1
3 15 9 9
8 15 13 9 2 9 7 9 2
16 16 13 3 13 0 13 2 3 9 1 4 13 9 7 9 2
7 9 11 9 12 13 9 12
8 13 11 3 7 3 2 15 13
5 7 15 1 9 2
7 13 13 15 13 9 1 2
39 15 13 11 9 2 7 13 16 15 13 1 9 7 15 13 15 9 7 15 13 9 7 3 15 2 13 9 9 3 15 9 2 7 13 9 3 13 15 9
8 15 9 13 4 3 13 13 9
8 9 13 11 9 7 0 9 2
5 13 3 16 9 2
2 9 0
14 11 13 9 13 9 2 7 3 9 4 13 9 1 2
12 11 9 9 13 13 15 3 0 13 0 9 2
12 9 13 3 4 13 9 0 0 9 11 9 9
9 15 13 3 9 2 13 9 3 2
8 11 9 13 0 9 9 9 2
8 13 9 16 3 16 13 9 2
5 15 15 15 13 2
19 9 13 3 0 9 2 12 9 9 13 13 13 2 3 9 13 13 9 2
10 11 13 0 7 0 9 3 3 9 2
6 13 3 16 0 9 2
8 9 15 13 0 11 9 13 2
4 9 13 0 9
6 9 13 3 9 9 2
7 13 15 3 13 9 16 9
8 9 11 13 11 9 1 9 2
14 15 13 13 3 2 16 9 7 9 9 13 3 9 2
7 11 9 13 0 9 9 2
4 11 15 13 2
5 3 15 13 9 2
8 9 13 2 16 13 15 0 2
5 9 15 4 13 2
6 9 9 16 13 13 2
6 13 13 9 0 9 2
8 15 9 13 3 13 1 15 2
5 15 13 0 9 2
5 13 3 15 3 2
9 13 3 9 2 13 3 3 9 2
8 9 13 3 0 16 0 9 2
3 13 9 9
7 13 3 13 3 15 9 2
7 15 13 3 13 0 9 2
10 3 9 0 9 9 9 13 13 15 2
4 13 13 0 2
12 13 3 0 9 9 2 16 13 0 9 13 2
7 15 9 15 9 4 13 2
6 13 2 16 6 9 2
7 13 0 16 13 13 9 2
10 15 3 13 2 16 0 9 4 13 2
2 13 13
2 9 1
8 12 9 13 9 13 9 1 2
13 9 13 7 3 11 9 3 3 13 7 3 3 2
10 9 13 4 13 9 2 7 3 9 2
9 9 13 13 3 15 9 13 9 2
7 0 9 13 3 13 3 2
9 11 9 11 11 4 13 12 9 2
6 4 13 3 12 9 2
2 3 11
2 13 9
2 6 6
16 9 11 13 0 0 9 2 11 9 2 7 15 13 15 9 2
15 15 15 13 2 16 15 9 13 13 9 7 13 3 3 2
8 15 13 9 11 9 0 9 2
8 15 15 3 13 15 0 9 2
3 9 7 9
6 12 9 13 9 15 9
10 9 13 9 9 13 12 12 12 9 2
10 13 4 15 13 13 13 2 4 13 2
7 16 9 13 13 3 3 2
7 3 9 13 0 9 9 2
3 13 3 2
11 9 13 3 11 3 0 9 13 11 11 2
7 4 11 13 9 7 9 2
10 3 2 13 13 9 1 9 2 15 2
3 15 13 3
2 0 9
13 15 2 13 9 0 7 0 9 2 13 13 15 2
8 13 16 13 9 15 13 3 2
15 2 4 13 0 0 9 2 16 9 4 13 3 0 2 2
10 4 15 15 0 13 2 9 11 13 2
2 13 3
3 15 13 15
3 13 4 13
7 13 13 9 7 9 7 9
12 3 15 3 13 16 9 13 7 13 0 9 2
12 9 13 3 4 13 9 2 9 9 13 9 2
7 11 9 4 13 0 9 2
2 3 3
3 9 4 13
6 15 13 9 3 13 9
10 2 15 4 3 13 9 2 13 15 2
12 15 15 13 9 3 13 13 9 0 0 9 2
16 16 15 13 2 13 13 9 2 7 15 9 15 13 13 13 2
5 15 13 3 9 2
5 11 13 3 0 2
10 0 9 13 0 9 0 7 0 9 2
13 13 15 4 13 13 9 9 3 7 13 15 9 2
6 9 13 15 9 3 2
13 11 13 0 9 16 11 7 11 7 0 16 11 2
5 9 9 0 0 9
7 9 9 4 3 13 9 2
2 13 0
10 7 15 9 13 3 13 13 9 9 2
5 15 13 3 9 2
10 15 13 9 15 3 16 4 13 15 2
5 9 13 9 13 2
4 13 9 9 2
6 0 9 13 9 11 2
8 13 3 13 16 15 13 3 3
10 9 9 7 9 13 9 15 9 9 2
2 15 2
3 13 9 9
5 15 13 0 0 9
10 9 4 13 2 7 15 13 13 0 2
12 0 7 0 9 0 9 4 13 12 12 9 2
9 9 4 9 13 3 9 13 9 2
9 4 15 3 13 2 13 15 13 2
3 15 13 0
9 9 13 13 9 2 7 9 3 2
3 15 13 15
8 0 9 9 13 0 9 9 2
9 11 13 11 12 9 0 12 9 2
6 11 13 9 3 0 2
3 3 1 9
3 9 4 13
5 13 15 3 9 2
7 3 15 9 13 4 13 2
18 7 3 13 3 2 13 16 9 13 3 13 7 13 9 2 3 9 2
8 13 2 16 15 13 3 9 2
14 3 9 13 9 13 9 7 11 13 2 7 3 3 9
6 13 9 9 7 13 2
8 9 13 9 15 4 13 3 2
5 3 3 13 9 2
7 9 13 0 9 11 11 2
3 0 13 2
4 13 15 9 2
15 9 15 13 9 11 2 9 9 2 7 15 15 13 0 2
5 15 13 3 9 2
8 3 0 13 9 13 3 9 2
2 9 13
12 9 11 11 9 11 9 4 13 11 9 9 2
12 9 9 1 4 13 12 16 13 3 12 12 9
8 15 15 4 13 3 13 15 2
9 15 13 13 0 9 13 15 0 2
11 13 15 13 0 16 0 9 13 15 9 2
11 15 9 13 9 2 15 13 3 0 9 2
6 15 13 3 1 15 2
7 15 15 3 4 13 9 2
13 0 9 13 13 3 0 9 2 13 0 7 0 2
6 3 15 13 0 0 2
5 15 13 13 9 13
2 0 9
11 11 13 3 0 2 12 9 13 9 9 2
5 3 11 13 3 2
7 11 11 2 13 15 3 9
11 3 9 13 0 9 2 16 13 3 9 2
4 13 13 0 2
9 2 3 3 2 15 13 3 3 2
3 9 7 9
4 16 15 9 2
2 0 0
9 0 9 15 3 13 2 11 13 2
15 9 13 9 13 3 2 16 15 9 13 3 3 9 1 2
6 9 13 9 7 9 9
13 15 15 13 9 9 2 7 15 13 3 3 9 2
2 0 9
5 2 9 13 9 2
9 9 13 9 2 15 13 3 3 2
12 9 9 13 4 13 15 13 3 0 9 9 2
14 9 13 2 16 11 13 15 9 9 7 13 15 9 2
9 2 13 9 2 2 13 9 3 2
12 15 4 3 13 2 16 13 3 13 11 1 2
4 11 13 9 2
14 11 13 13 11 2 7 9 13 9 1 13 9 1 2
8 7 9 1 15 3 4 13 2
19 3 4 13 9 13 2 16 11 11 13 13 2 7 16 11 11 13 9 2
4 9 1 9 2
4 15 13 0 2
3 9 3 2
12 15 1 11 4 13 9 9 9 7 9 9 2
8 9 12 9 9 13 15 9 2
8 3 3 12 12 9 13 13 2
4 13 0 9 2
27 15 13 12 9 9 15 15 13 9 2 9 2 9 7 9 2 15 15 13 2 13 7 13 9 1 9 2
7 15 13 9 7 13 9 2
10 15 9 13 0 2 0 9 13 9 2
7 9 13 13 7 9 13 2
5 0 9 13 0 2
3 9 13 9
9 11 9 9 4 13 9 9 3 2
2 13 13
3 15 9 2
2 0 9
15 12 15 9 15 11 11 3 15 4 13 3 13 15 9 2
9 16 13 13 2 3 15 13 9 2
2 0 9
10 9 9 13 15 9 0 16 13 9 2
3 9 13 11
6 0 3 13 15 9 2
6 9 0 9 13 9 2
2 9 13
10 15 9 13 3 0 0 7 3 9 2
11 9 9 13 16 15 3 4 13 15 3 2
6 11 13 11 0 9 2
29 7 0 15 9 3 15 16 16 13 3 0 9 7 13 3 13 9 3 13 15 13 3 15 16 15 15 9 13 2
4 7 6 13 2
3 13 13 9
6 9 13 3 7 3 2
2 6 2
7 15 13 9 9 1 9 2
14 9 9 13 3 0 2 16 13 9 4 13 9 13 2
7 9 13 13 0 7 0 2
8 9 13 9 9 7 9 9 2
12 9 1 4 13 3 0 9 9 2 7 9 2
12 11 13 11 2 16 3 13 13 9 1 9 2
4 0 9 9 2
12 11 11 13 15 3 16 15 13 15 7 15 2
8 16 9 13 9 2 13 9 2
11 9 13 13 9 3 3 2 16 4 13 2
7 15 13 3 3 3 11 2
4 3 3 11 2
4 3 15 9 2
8 2 6 2 13 15 0 9 2
8 9 9 13 11 13 9 11 2
5 12 9 9 13 2
2 9 2
7 9 15 13 0 9 1 2
9 15 15 13 3 9 1 3 9 2
4 15 15 13 2
12 0 9 9 9 13 2 16 15 13 9 13 2
12 13 15 4 13 13 15 15 1 16 11 13 9
5 15 13 0 13 15
3 3 3 16
7 9 4 13 9 11 1 2
8 11 13 9 3 7 9 9 2
3 3 13 3
6 15 9 15 4 13 2
6 4 13 0 9 9 2
6 12 9 9 13 9 2
13 9 13 9 9 2 3 9 9 7 0 9 9 2
10 13 3 0 2 7 13 13 3 13 2
3 3 9 1
10 15 4 13 15 9 3 15 3 13 2
5 15 13 13 9 2
6 3 3 13 13 9 2
8 15 15 4 13 3 0 9 2
13 13 0 2 16 13 9 2 9 9 7 15 9 2
4 13 12 9 2
9 15 13 9 2 1 11 13 9 2
16 3 15 13 0 9 9 2 3 15 4 13 9 7 13 9 2
16 9 13 3 9 9 2 13 3 15 0 12 12 9 9 13 2
4 15 13 0 2
3 13 15 13
14 3 15 2 12 3 3 3 3 3 7 2 3 3 0
16 0 9 9 9 2 15 13 9 15 9 2 13 9 0 9 2
10 15 13 15 13 13 9 9 9 9 2
14 15 13 2 16 9 4 13 0 9 7 15 4 13 2
22 15 9 13 9 1 13 7 15 13 9 13 2 15 1 15 13 13 9 13 9 3 2
12 0 2 0 2 16 13 13 0 9 13 11 2
8 16 9 13 2 4 13 9 2
4 13 3 3 2
16 9 2 9 7 9 13 13 3 2 16 15 0 9 13 9 2
7 15 4 13 9 9 1 2
17 11 11 13 15 9 15 3 0 9 0 9 2 3 13 3 9 2
9 11 13 9 2 7 9 13 9 2
11 9 13 3 3 3 15 1 2 11 13 2
5 2 13 13 3 2
10 13 2 16 13 9 13 13 11 9 2
7 11 13 0 9 13 9 2
9 0 9 13 9 7 11 13 9 2
3 13 3 2
16 16 9 13 9 2 13 4 13 15 2 16 13 15 9 13 2
4 15 4 13 2
15 11 13 11 9 3 13 9 0 16 0 11 9 13 9 2
5 3 0 15 15 13
4 11 13 13 2
7 15 9 13 3 0 9 2
3 13 9 1
13 0 9 13 12 0 11 11 9 11 7 11 9 2
11 15 13 3 3 9 0 16 15 9 3 2
17 7 15 13 16 15 15 3 13 0 9 7 0 7 9 13 3 2
2 13 13
13 9 13 2 16 11 13 4 3 0 9 13 3 2
3 13 3 3
14 3 11 13 15 9 2 16 9 13 0 9 9 13 2
5 15 13 9 3 9
12 15 11 13 3 3 11 9 16 13 13 9 2
13 15 13 9 7 9 2 15 3 13 9 7 9 2
7 15 13 12 7 12 1 2
4 9 13 0 2
9 7 9 13 3 9 3 0 9 2
3 9 13 13
7 13 12 9 9 7 9 2
19 9 2 15 13 13 15 9 13 3 2 13 15 9 3 13 3 13 9 2
4 0 13 13 2
4 13 3 0 2
14 15 15 13 2 16 15 13 9 2 15 9 15 13 2
11 15 13 0 9 3 0 7 3 0 9 2
10 3 9 13 3 16 13 9 15 1 2
8 9 13 13 9 0 0 9 2
4 9 15 13 0
15 11 9 13 11 9 2 0 2 0 2 0 2 0 9 2
6 0 9 15 13 9 2
7 13 15 15 13 7 13 2
13 9 9 7 9 9 9 13 7 9 7 9 9 2
3 13 9 2
19 15 13 15 9 11 0 9 2 15 13 13 9 15 3 16 11 9 9 2
6 7 15 13 0 13 2
10 16 9 13 3 2 9 13 3 13 2
10 15 9 11 9 9 13 3 12 9 2
8 9 7 9 13 9 1 9 2
5 11 13 3 9 2
6 3 3 13 7 13 2
7 15 13 9 3 3 9 2
14 15 13 2 16 9 13 2 9 13 1 2 9 13 2
5 9 13 15 13 9
9 9 9 3 13 9 11 11 9 2
6 15 13 0 9 0 2
6 3 11 9 13 0 2
11 9 2 15 13 2 16 15 13 3 13 2
7 15 13 12 0 9 9 2
18 11 9 13 2 16 9 4 13 3 12 9 9 2 15 13 3 0 2
11 15 4 13 15 9 2 15 9 13 13 2
11 11 13 13 15 3 9 11 5 11 1 2
7 9 9 15 13 0 9 2
8 11 13 9 3 3 3 15 9
4 9 13 0 2
3 11 13 2
16 13 13 9 9 7 9 1 3 3 13 9 13 13 9 9 2
5 9 13 3 0 2
2 9 9
8 0 11 9 4 13 9 12 2
17 11 4 13 11 9 0 9 1 13 9 4 13 12 9 9 9 2
3 9 15 13
4 9 9 13 9
9 11 13 13 9 7 9 3 9 2
13 0 9 9 13 9 9 9 3 9 11 11 9 2
4 13 16 4 13
7 9 9 13 3 0 9 2
8 9 9 13 3 12 12 9 2
17 9 13 0 3 2 3 9 13 3 9 3 9 3 13 9 9 2
14 15 15 3 9 9 9 2 15 3 13 0 0 9 2
5 15 4 3 3 13
7 3 15 4 13 11 13 2
9 13 3 2 9 3 13 11 1 2
14 15 9 13 3 9 11 9 2 15 4 13 9 11 2
13 13 13 2 16 3 13 4 13 3 9 9 9 2
10 3 13 9 2 16 4 9 13 3 2
7 0 9 15 4 13 6 2
13 15 9 4 13 3 2 16 3 9 13 13 9 2
5 15 13 9 9 2
10 13 15 13 9 9 15 15 0 9 2
16 3 13 9 13 15 2 15 3 15 9 4 13 3 0 9 2
3 15 11 2
4 9 4 13 2
11 11 9 13 0 2 7 9 4 13 3 2
16 13 13 15 2 9 7 9 2 15 13 9 9 9 2 16 2
3 0 9 2
2 13 3
6 13 2 16 13 3 2
4 9 13 0 2
6 13 9 9 9 1 2
13 15 13 13 2 11 13 2 16 9 13 13 9 2
4 13 15 11 2
11 9 13 3 3 3 9 1 15 2 16 2
21 4 9 13 2 16 15 13 9 9 2 7 13 4 13 2 16 15 13 9 9 2
8 3 13 15 13 9 9 11 2
5 15 13 13 13 13
8 15 13 13 15 13 0 9 2
9 4 13 0 2 16 9 13 9 2
9 15 13 12 9 9 3 13 3 2
4 13 0 9 2
4 11 13 11 9
4 9 11 9 13
13 7 15 13 13 9 2 7 0 9 2 15 9 2
13 12 9 13 9 9 13 0 9 9 9 7 9 2
3 15 13 9
9 15 13 2 16 15 13 9 0 2
10 15 13 9 2 16 15 13 13 9 2
6 11 11 13 3 9 2
2 0 9
2 0 9
5 9 13 11 9 2
13 4 3 0 9 3 13 2 15 13 4 3 13 2
12 11 1 9 4 13 15 9 9 15 13 9 2
3 9 11 9
14 0 9 13 9 15 2 16 9 13 7 13 15 9 2
5 13 9 0 9 2
21 15 3 4 13 3 15 9 2 7 15 0 9 13 3 11 2 3 2 3 3 2
12 11 9 13 3 0 13 9 16 9 3 9 2
13 4 9 13 9 9 9 2 7 16 2 3 3 2
24 9 9 13 3 0 0 9 2 15 13 15 9 0 9 2 15 9 9 13 13 3 13 9 2
6 9 4 9 13 9 2
2 0 9
19 9 13 3 3 3 3 16 9 9 2 7 15 13 7 13 3 3 9 2
2 9 0
14 9 9 4 9 1 13 11 9 12 9 11 9 1 2
2 0 9
6 2 15 13 9 13 2
6 0 9 15 3 13 2
4 15 15 13 2
6 9 13 9 9 3 2
11 13 11 7 11 13 11 13 11 11 9 2
14 15 13 0 9 7 13 3 13 2 16 15 13 13 2
10 13 2 16 3 13 9 1 15 9 2
11 0 9 13 13 13 2 16 9 13 13 2
12 11 9 9 11 11 1 9 13 13 13 13 2
20 7 16 15 15 13 3 15 2 9 11 3 15 13 3 0 13 15 13 15 2
7 11 4 13 15 0 9 2
10 13 0 0 9 2 16 9 4 13 2
11 15 9 15 13 0 9 9 9 1 11 2
4 15 4 13 2
14 11 2 15 13 3 15 9 15 13 3 3 9 13 2
9 11 13 4 13 11 9 13 9 2
5 11 2 11 13 9
14 15 13 3 0 9 2 16 9 3 13 2 9 13 2
12 11 4 3 13 9 7 13 3 9 9 13 2
5 13 9 0 9 2
6 16 13 3 13 3 2
11 13 15 0 9 16 15 4 13 9 9 2
21 7 15 13 3 3 9 0 8 8 9 15 16 3 13 16 13 3 0 13 9 2
8 3 9 4 9 13 1 9 2
2 3 16
15 3 13 15 16 15 15 9 13 13 15 0 16 0 9 2
6 3 9 13 9 0 2
3 15 9 0
15 15 2 16 9 13 2 13 15 2 16 4 13 3 0 2
5 16 13 11 13 2
3 9 13 0
5 13 3 0 11 2
4 15 15 13 2
2 13 13
8 15 12 9 11 13 11 9 2
8 3 3 9 3 13 11 9 2
4 12 13 9 2
4 3 13 3 2
4 9 9 11 1
14 13 13 7 3 11 9 0 9 2 15 9 13 3 2
15 9 7 9 13 13 9 2 3 13 9 13 13 15 0 2
11 0 9 13 0 2 15 3 0 13 0 2
4 3 13 0 9
2 11 11
9 13 13 2 16 13 9 13 0 2
3 0 0 9
3 13 15 15
11 4 15 13 2 3 4 13 15 0 9 2
4 13 15 3 2
7 0 9 13 3 0 11 2
5 9 13 9 13 9
14 9 7 9 15 13 2 11 4 3 13 0 9 9 2
12 11 4 3 12 9 13 13 3 0 16 3 2
5 9 13 13 13 2
6 15 13 13 9 1 2
5 15 15 15 13 2
11 15 2 15 13 13 13 15 3 2 13 2
8 13 9 9 9 7 13 9 2
19 15 9 11 13 13 9 9 9 3 9 2 16 9 9 4 4 13 3 2
12 3 0 3 15 13 2 9 4 13 13 9 2
5 9 13 7 0 2
5 0 9 13 0 2
12 15 9 15 13 9 2 16 9 13 9 9 2
7 9 13 9 9 13 9 2
7 13 15 13 15 1 13 2
12 3 15 13 2 16 13 15 3 9 4 13 2
6 15 4 13 13 9 2
14 9 13 9 2 16 9 13 9 9 11 0 11 9 2
5 9 13 9 1 2
4 9 13 9 2
5 11 11 13 9 2
9 3 13 15 2 15 3 13 9 2
7 7 3 13 9 3 9 2
4 0 9 7 9
7 15 9 13 12 0 9 2
12 13 16 9 7 9 13 0 7 13 0 9 2
2 13 3
5 3 13 0 0 2
3 4 13 2
10 3 11 15 9 13 9 9 9 13 2
8 13 3 15 9 13 15 9 2
11 2 9 13 3 13 3 2 16 3 13 2
15 3 3 11 7 11 13 9 2 3 15 3 13 0 9 2
14 15 15 13 2 9 9 9 1 9 2 9 7 0 2
11 9 1 13 13 9 2 15 4 9 13 2
4 15 13 9 2
3 3 15 1
3 15 13 0
9 13 9 15 0 9 15 0 9 2
3 9 13 0
9 15 13 9 1 2 13 7 13 2
4 9 13 0 2
5 4 13 3 9 2
4 13 3 9 2
5 9 13 9 9 13
15 9 3 13 15 13 9 9 2 3 3 3 3 13 13 2
10 11 0 9 13 9 2 9 7 9 2
16 16 13 16 9 13 13 2 9 13 16 4 3 13 3 9 2
10 9 4 13 9 1 3 9 9 0 2
8 0 9 13 3 0 0 9 2
11 16 15 13 9 13 3 15 13 16 13 15
2 11 9
19 9 9 1 13 9 9 1 2 7 15 13 15 2 16 13 15 3 9 2
3 13 13 2
10 9 13 12 9 7 13 9 12 9 2
9 15 4 13 0 9 15 4 13 3
8 15 3 4 13 9 15 13 2
8 13 3 0 2 13 0 0 2
8 11 11 13 3 9 13 3 3
15 9 13 3 9 9 9 2 7 3 13 9 3 0 9 2
5 3 9 13 3 3
4 15 4 13 2
22 9 15 13 9 3 3 2 13 9 9 7 13 2 16 13 9 2 13 3 3 3 2
12 15 13 6 13 15 7 13 15 3 9 1 2
4 0 9 1 13
5 9 13 3 3 2
5 3 13 13 9 2
12 3 15 4 3 13 9 2 7 13 13 15 2
5 15 13 9 13 2
18 3 9 3 15 9 13 9 13 9 2 16 4 13 3 3 15 0 2
8 9 9 13 9 0 0 9 2
8 13 15 9 9 9 7 9 2
7 15 9 13 11 0 9 2
12 15 13 3 3 2 16 9 13 9 13 9 2
3 13 13 2
24 15 9 4 13 2 16 3 0 9 13 0 13 9 3 7 9 3 2 16 3 9 13 4 2
12 9 13 9 11 9 2 9 2 13 3 9 2
9 3 11 7 15 12 9 13 9 2
9 9 13 0 2 7 9 9 0 2
4 9 13 0 2
7 11 13 0 0 16 9 2
4 0 13 11 2
18 15 4 13 0 9 7 0 9 2 9 3 7 3 3 3 7 3 9
15 4 15 13 3 9 3 12 9 2 13 3 15 9 1 9
3 13 9 12
9 0 11 11 9 9 13 9 11 9
5 15 13 15 1 2
6 13 9 7 13 13 2
6 13 9 9 7 9 2
5 3 3 0 13 2
18 9 4 13 13 3 2 16 13 15 13 9 13 0 9 0 9 1 2
12 6 6 2 15 13 16 9 13 3 9 13 2
5 15 13 11 9 2
3 15 0 9
4 15 9 13 15
3 15 9 2
14 13 0 9 13 2 15 11 7 11 13 13 13 9 2
5 4 13 13 9 2
6 9 13 0 9 13 2
2 15 9
6 2 9 13 3 13 2
13 15 13 3 9 2 16 13 9 0 9 13 11 2
10 15 9 13 11 13 9 9 9 9 2
13 15 13 15 3 15 15 9 1 2 7 13 11 2
4 13 9 0 9
10 15 15 13 0 9 7 9 4 13 3
7 15 9 13 3 7 3 0
5 3 13 3 9 2
4 9 13 0 9
5 15 9 9 13 9
7 0 9 13 3 15 1 2
12 9 4 4 9 13 3 2 16 15 13 9 2
7 11 11 13 9 9 9 2
19 13 15 16 15 13 9 7 9 7 9 7 9 7 9 7 9 7 9 2
11 3 13 9 2 7 15 0 13 0 9 2
4 3 4 13 9
8 9 13 3 0 16 3 3 2
3 6 15 9
13 13 3 9 9 7 15 9 7 3 9 13 3 2
2 3 3
13 11 13 9 12 13 3 15 2 3 9 13 9 2
5 9 13 9 9 2
9 0 15 9 4 4 13 9 9 2
8 9 1 11 4 13 0 9 2
4 15 13 3 2
4 9 13 3 2
5 13 15 1 9 2
6 15 13 0 9 9 2
6 13 3 13 15 9 2
6 13 9 9 3 9 2
2 15 9
5 15 13 9 9 2
11 13 13 2 16 11 13 9 0 9 1 2
25 9 13 9 3 3 2 3 9 13 13 7 3 15 1 13 2 13 7 13 9 9 7 9 9 2
5 9 13 9 9 2
8 9 9 15 9 13 3 0 2
14 9 13 9 3 15 2 15 9 2 7 3 0 9 2
9 2 9 2 1 9 2 13 2 2
8 15 13 9 13 13 3 9 2
2 0 9
10 13 15 3 2 16 3 13 9 9 2
8 15 4 13 3 3 3 12 9
15 11 13 0 9 2 11 9 9 2 15 0 9 9 13 2
4 9 13 0 2
11 11 13 9 0 9 2 0 13 0 9 2
17 7 15 2 15 9 9 3 13 2 13 9 7 15 13 9 9 2
2 6 2
15 11 9 13 0 2 16 3 11 9 4 13 9 15 0 2
15 9 9 13 15 2 13 9 13 9 9 13 7 13 9 2
6 9 13 13 13 9 2
4 15 13 13 3
3 13 9 2
10 9 13 3 9 7 15 13 9 0 9
7 4 0 7 3 13 0 9
5 9 13 0 9 2
24 9 2 15 9 0 9 3 9 0 9 2 3 9 13 9 3 13 3 3 7 13 9 9 2
13 9 9 13 15 2 16 9 4 13 0 9 1 2
5 0 9 13 9 2
6 15 13 13 15 13 2
13 3 13 3 3 3 3 0 2 0 7 0 9 2
8 9 13 4 13 3 12 9 2
9 15 3 13 13 3 0 9 9 2
4 13 13 9 3
21 11 9 9 13 3 1 9 0 2 16 15 9 4 13 15 9 11 11 9 9 2
7 9 1 4 13 2 16 2
4 9 13 9 2
7 15 13 11 9 11 9 2
6 0 9 13 0 11 2
4 9 1 13 2
7 9 9 4 3 13 3 2
7 9 13 13 3 12 9 2
5 12 9 1 13 11
10 11 9 13 11 0 9 9 3 9 2
11 16 13 3 2 16 13 13 12 9 0 2
6 15 13 13 15 0 2
17 15 13 15 3 9 9 15 15 13 16 15 13 11 3 3 9 2
5 13 15 3 15 2
5 13 0 13 0 2
11 11 11 11 9 13 0 9 3 9 12 2
9 15 0 9 15 4 3 9 13 2
7 13 15 3 15 3 13 2
8 15 13 3 0 0 9 1 2
3 13 11 9
5 13 9 0 9 2
10 11 11 12 0 9 4 3 13 9 2
3 11 0 9
11 0 12 9 9 13 4 13 3 13 9 2
6 9 13 9 13 3 2
10 0 9 11 13 9 9 11 9 1 2
29 15 4 13 2 3 3 0 2 0 9 3 3 13 2 15 9 7 2 0 2 3 15 9 15 4 13 7 2 0
9 0 9 13 13 13 0 9 9 2
8 11 9 9 9 9 13 9 2
3 13 11 2
18 9 13 9 2 15 3 15 13 13 13 2 7 15 15 13 4 13 2
4 15 16 13 15
7 9 9 13 3 3 0 2
15 15 13 0 2 7 3 9 13 9 2 15 0 9 13 2
16 4 15 2 13 4 2 11 11 13 13 7 0 9 0 13 2
22 6 3 2 6 4 3 13 3 15 9 3 7 9 3 13 3 16 15 0 15 13 2
8 9 11 11 13 9 11 9 2
4 9 13 15 9
6 15 13 3 9 1 15
12 11 13 9 9 2 13 11 7 13 0 9 2
9 9 13 3 16 4 13 9 0 2
24 15 4 13 9 13 7 13 15 2 15 15 0 9 13 0 2 7 9 7 9 7 0 15 2
5 11 13 9 9 2
8 15 15 13 9 2 13 0 2
10 0 9 13 11 11 9 13 9 9 2
2 0 9
12 13 9 9 13 9 3 2 16 15 13 13 2
7 15 13 13 0 0 9 2
10 3 13 12 0 9 2 15 13 9 2
13 7 11 4 3 15 9 13 3 12 9 0 9 2
7 11 13 9 1 11 11 2
5 2 13 15 3 2
16 9 7 0 9 13 9 3 9 9 2 0 9 9 7 9 2
12 11 9 13 13 9 2 3 15 9 13 9 2
8 11 13 9 1 3 13 9 2
9 9 1 9 13 9 1 4 13 2
4 3 15 13 9
5 15 3 9 13 2
14 15 15 0 11 13 9 9 1 7 13 3 15 9 2
4 13 3 3 13
13 9 9 13 9 2 16 15 15 13 2 13 3 2
11 15 13 2 7 15 15 2 9 0 9 2
7 9 13 3 15 9 9 2
7 13 2 16 15 13 11 2
7 3 15 13 2 13 9 9
19 0 9 9 13 15 9 3 12 9 9 2 7 15 9 13 3 3 9 2
4 9 1 13 9
18 9 13 0 2 9 0 7 0 2 9 0 2 1 7 1 12 9 2
8 15 9 13 13 9 7 9 2
10 15 13 0 13 2 7 13 13 15 2
19 0 9 0 7 0 9 9 4 11 9 13 9 3 0 2 0 7 0 2
13 15 4 13 15 15 2 15 4 13 7 15 13 2
10 11 13 3 9 0 7 9 7 9 2
10 11 12 9 9 12 0 9 13 9 2
4 15 13 9 11
7 15 7 15 13 3 9 2
5 9 13 3 9 2
6 15 6 15 9 13 2
7 15 15 13 9 15 9 2
3 13 4 13
8 15 3 13 3 15 2 16 2
7 15 13 0 9 2 13 2
11 0 9 13 9 13 13 13 13 15 3 2
9 9 13 3 13 9 2 13 9 2
13 11 9 7 9 9 0 9 9 13 3 13 9 2
7 13 9 9 3 13 9 2
6 11 13 3 0 9 2
6 3 15 13 3 9 2
10 11 9 9 13 0 9 0 12 9 2
11 6 6 2 3 15 3 13 2 9 13 2
6 9 13 15 13 3 2
9 6 2 15 13 3 15 3 0 2
10 9 7 9 0 9 13 9 0 9 2
4 15 13 3 9
6 9 13 15 13 9 2
10 9 13 15 9 7 9 7 0 9 2
7 13 9 13 7 9 13 2
6 13 2 16 15 13 2
2 9 9
5 9 13 4 13 9
14 0 7 9 9 13 15 9 3 9 13 7 9 9 2
4 9 13 0 9
5 9 9 4 13 2
6 11 9 9 9 13 2
6 3 11 13 13 9 2
3 0 9 2
9 15 13 13 9 2 4 13 9 2
6 11 13 11 7 9 2
17 3 13 3 2 7 13 15 3 3 0 16 13 9 0 9 9 2
2 6 6
3 9 13 2
4 13 15 3 2
4 9 13 9 2
6 7 15 13 13 15 2
11 3 15 13 0 2 15 13 4 3 13 2
5 9 13 9 9 2
7 12 0 9 13 3 9 2
13 9 13 13 11 15 3 0 9 2 7 13 0 2
8 11 9 13 3 7 13 3 2
7 0 13 9 2 9 9 2
6 13 12 9 9 9 2
9 0 9 12 9 9 13 3 9 2
17 4 15 11 13 16 15 13 3 16 15 13 9 9 16 4 13 15
13 9 4 13 3 1 2 1 9 15 13 13 15 2
8 15 13 16 15 13 15 9 2
10 3 13 9 13 13 9 9 9 1 2
4 9 13 15 9
6 11 11 13 1 9 2
8 15 9 4 12 9 13 11 2
3 13 3 2
17 9 4 13 3 2 16 16 13 9 2 13 0 9 15 9 9 2
4 9 13 1 9
3 9 3 2
8 15 4 13 9 13 15 9 2
7 0 9 4 13 3 9 2
5 13 9 13 0 2
4 9 13 13 9
6 13 9 13 3 3 2
12 3 9 13 9 4 13 0 7 0 9 15 2
18 16 13 13 7 13 0 9 13 4 13 9 11 7 13 13 13 9 2
3 15 13 15
7 13 15 13 13 3 9 2
9 11 9 11 4 9 13 13 9 2
6 15 9 13 11 9 2
6 13 3 16 13 3 2
13 11 0 11 11 11 13 9 7 3 3 13 13 2
10 13 9 0 9 2 16 13 15 3 2
15 15 9 9 9 4 13 2 13 15 0 9 16 9 9 2
17 0 9 4 13 15 2 13 9 7 0 9 0 0 9 9 9 2
6 0 9 9 13 11 2
7 9 15 13 9 9 13 9
14 13 15 3 9 7 2 9 7 9 16 15 13 3 2
13 0 9 13 2 16 13 13 0 2 3 3 0 2
12 9 13 9 3 13 3 13 9 13 9 3 2
4 13 9 1 9
10 3 11 13 2 16 15 9 13 3 2
9 16 15 13 3 13 9 13 3 2
10 3 15 3 9 4 9 13 9 3 2
9 11 4 9 13 16 9 13 9 2
11 15 9 16 9 13 2 15 13 15 9 2
4 0 9 0 9
5 2 13 3 15 2
5 13 13 3 0 2
2 13 13
4 9 13 16 13
6 15 13 13 0 9 2
8 0 12 0 9 9 13 11 2
4 9 13 3 2
7 9 4 13 15 9 9 2
8 3 0 9 9 4 13 9 2
3 2 3 2
3 3 3 2
4 0 7 0 9
7 0 9 11 13 13 9 2
2 13 2
2 13 9
7 15 9 9 9 4 13 2
20 11 11 2 9 7 11 9 11 13 3 9 9 1 7 15 9 11 9 13 3
4 13 15 11 2
5 15 13 9 15 2
7 15 9 9 13 9 9 2
4 12 9 0 9
9 13 13 0 9 13 9 2 13 2
6 13 3 9 9 9 2
5 3 3 0 9 2
16 9 9 7 9 9 9 13 3 3 2 16 11 13 3 0 2
5 9 13 9 1 2
11 15 9 4 13 3 9 9 2 9 13 2
5 13 9 13 15 2
5 3 3 3 13 2
8 13 12 13 3 0 0 9 2
7 9 4 13 3 12 9 2
8 15 4 3 13 3 9 1 2
5 9 13 13 9 15
7 15 13 13 15 9 3 2
8 3 0 15 13 2 11 9 2
7 7 13 13 15 9 9 2
4 2 15 9 2
4 13 3 11 2
12 3 4 13 3 15 9 2 7 13 13 13 2
11 9 11 9 13 0 2 7 9 13 0 2
14 16 0 9 9 9 13 11 13 2 3 3 9 4 13
7 9 13 3 3 11 9 2
20 9 9 2 7 9 15 15 9 4 3 16 4 0 15 9 9 2 3 9 2
17 9 9 9 9 13 15 2 16 11 9 13 9 11 11 9 9 2
15 16 0 9 13 3 2 0 9 9 13 3 13 9 0 2
9 3 15 13 15 15 15 15 0 13
5 15 4 15 9 13
12 7 3 13 3 9 3 3 15 13 4 13 2
12 11 13 2 13 9 7 13 9 9 9 2 2
12 16 12 0 9 9 13 2 9 13 15 0 2
9 11 13 9 13 3 15 0 9 2
7 0 4 13 0 9 9 2
8 15 13 13 7 13 9 9 2
11 9 3 13 0 9 2 16 13 3 13 2
5 16 13 13 3 2
5 13 15 13 9 2
12 4 13 9 9 7 3 4 9 13 3 9 2
11 9 13 11 9 0 9 9 9 11 9 2
3 0 9 9
7 3 9 13 9 13 3 2
4 13 16 13 2
3 13 13 2
7 9 13 3 2 3 3 3
14 9 7 9 13 9 1 3 15 2 15 13 13 9 2
4 15 13 16 9
21 13 9 2 3 9 13 0 13 15 9 2 16 15 3 13 15 9 16 4 13 2
10 13 9 13 9 16 9 4 13 9 2
5 9 13 13 0 2
2 0 9
11 9 9 11 11 13 11 13 0 9 11 2
11 9 4 13 9 3 11 7 11 1 11 2
4 9 13 9 2
10 9 13 9 2 15 4 13 7 13 2
4 9 13 3 2
18 7 15 13 3 2 16 9 13 15 2 15 13 9 1 0 9 9 2
3 13 3 2
9 11 13 9 13 9 3 7 3 2
2 9 9
4 13 0 9 2
4 12 9 13 3
11 3 0 9 13 11 7 11 9 11 1 2
7 0 9 13 3 9 9 2
2 13 13
19 16 15 3 13 13 3 9 7 13 3 3 2 15 13 9 9 13 15 2
2 15 3
6 3 15 3 9 13 2
11 7 9 9 7 9 9 13 15 12 9 2
5 13 12 0 9 2
8 7 3 4 13 13 0 9 2
12 15 9 13 12 9 3 16 15 0 9 13 2
11 2 9 2 2 15 13 9 9 9 9 2
14 9 4 13 3 0 3 2 15 9 13 0 13 3 2
8 15 13 13 3 3 9 9 2
6 13 13 13 0 9 9
21 9 13 4 13 3 9 3 2 15 4 13 0 9 3 7 13 15 9 0 9 2
16 9 9 13 3 9 2 16 9 4 13 12 9 9 0 13 2
16 13 3 2 16 3 9 9 13 3 0 0 9 13 0 9 2
3 13 3 2
11 4 9 13 9 2 16 15 13 0 9 2
9 15 13 3 0 3 15 9 9 2
5 9 13 3 9 2
10 15 13 2 16 9 13 3 3 9 2
9 9 4 13 3 0 9 13 9 2
7 15 9 9 13 9 9 2
10 9 13 3 0 7 13 15 1 3 2
7 9 13 9 3 9 12 2
12 9 4 13 2 16 9 13 9 3 0 13 2
4 13 3 9 2
2 13 13
2 15 9
8 9 13 9 0 9 9 9 2
4 15 13 0 9
9 12 9 13 16 4 13 9 9 2
3 9 9 11
4 9 13 9 9
4 9 13 11 2
7 9 9 7 0 9 7 9
4 11 13 11 2
5 13 3 0 9 2
14 0 9 4 13 9 3 9 2 16 3 13 3 9 2
5 15 13 0 3 2
17 16 9 13 3 9 2 13 9 9 13 3 3 16 0 15 9 2
18 0 9 9 13 15 3 0 2 16 0 9 13 3 4 13 15 3 2
10 11 13 13 0 9 1 9 9 9 2
6 9 9 2 12 9 12
9 0 15 9 9 13 3 13 9 2
7 13 2 16 15 13 9 2
7 12 0 9 13 9 1 2
9 9 13 11 9 13 15 9 0 2
8 13 9 2 16 13 3 9 2
7 0 9 13 9 7 9 2
11 11 3 13 11 13 3 15 9 11 9 2
5 7 9 15 13 2
17 13 11 11 7 13 16 11 13 9 7 4 13 3 0 9 3 2
7 11 13 3 9 9 12 2
11 15 13 9 9 13 7 3 4 3 13 2
8 15 9 16 13 15 13 9 2
7 15 13 9 3 9 13 2
6 9 13 11 4 13 2
3 15 13 2
16 9 13 13 3 9 3 0 9 2 7 7 13 0 9 1 2
4 0 9 11 11
5 9 13 3 3 9
7 15 0 9 13 3 0 2
5 13 16 13 13 9
8 9 13 9 13 9 0 9 2
2 0 9
3 0 3 2
10 3 13 13 15 3 0 7 0 9 2
7 15 13 9 0 9 9 2
5 9 13 12 12 2
16 9 13 9 2 13 0 2 9 13 13 9 1 7 13 3 2
5 15 4 13 3 2
11 0 9 9 13 12 9 2 16 15 13 2
14 15 4 13 2 7 9 9 13 4 13 3 0 9 2
7 4 9 13 9 7 9 2
9 9 13 3 9 7 15 9 0 9
9 4 9 4 3 3 13 15 9 2
5 15 1 13 0 13
3 9 9 9
3 3 3 2
12 15 9 13 3 9 15 9 2 11 11 11 9
12 11 1 13 9 13 9 1 9 13 13 0 2
3 9 13 2
11 9 11 7 11 11 13 0 13 0 3 2
8 13 15 0 13 2 7 0 2
13 9 4 13 3 3 0 9 2 7 3 3 0 0
5 11 13 3 3 2
7 13 13 0 9 13 9 2
6 9 9 13 13 9 2
8 7 13 9 11 0 9 13 2
10 15 9 1 9 13 0 9 13 9 2
8 9 7 13 9 1 7 1 2
2 3 15
5 15 13 11 1 2
8 15 13 9 15 13 15 3 2
5 16 3 13 15 2
14 9 9 13 3 9 15 13 9 2 7 15 13 3 2
19 15 13 9 13 0 9 9 2 15 13 3 13 3 0 16 3 9 9 2
7 9 13 9 12 9 9 2
8 13 16 13 4 3 13 15 2
14 15 13 13 9 2 3 9 9 9 13 3 9 9 2
13 11 11 13 15 9 16 9 2 3 1 0 9 2
8 15 9 13 9 13 0 9 2
19 13 9 11 13 9 3 15 9 16 11 2 13 0 7 13 0 0 9 2
5 15 13 9 3 2
5 3 3 3 3 2
4 13 9 3 2
19 3 15 13 2 16 15 13 13 2 7 13 15 2 3 15 4 9 13 2
12 9 13 9 0 9 7 13 15 13 9 9 2
6 11 13 16 13 0 2
3 0 0 9
12 9 9 0 9 13 3 3 3 12 9 1 2
13 11 2 11 7 11 13 3 2 7 9 3 0 2
5 15 13 13 15 2
8 13 11 11 13 13 2 16 2
2 9 1
2 15 9
12 15 9 9 13 11 2 11 15 4 13 9 2
7 13 13 13 1 9 9 2
6 9 9 13 9 9 1
5 9 13 3 0 2
20 15 2 3 9 13 7 9 13 2 9 13 3 0 2 9 2 2 9 9 2
10 9 13 3 3 2 7 13 9 0 2
3 13 9 2
10 15 13 15 7 15 13 0 13 9 9
3 2 13 2
4 15 13 0 9
15 3 15 9 13 16 9 2 13 9 9 13 0 9 9 2
6 3 13 3 9 3 9
23 7 16 9 4 13 3 9 2 4 15 13 9 2 16 9 9 13 4 13 13 7 13 2
16 15 4 3 3 13 11 9 2 3 3 0 9 15 4 13 2
14 0 7 0 9 2 9 1 2 13 15 11 0 9 2
6 15 13 3 0 9 2
2 0 9
7 11 7 11 9 13 0 2
8 9 9 13 9 13 12 9 2
4 3 13 0 9
6 15 3 11 13 3 2
9 9 13 3 16 9 13 9 9 2
7 11 11 11 13 1 9 2
6 3 13 9 15 9 2
3 13 13 2
4 3 13 9 2
6 0 13 2 0 13 2
7 3 1 15 13 13 13 2
4 13 3 3 2
15 9 13 0 9 2 16 13 12 9 2 16 13 15 3 2
3 13 9 2
5 13 9 7 9 2
7 11 13 3 13 9 9 2
7 13 13 15 0 9 2 2
6 9 13 9 13 9 2
30 13 3 6 15 13 9 9 9 7 6 15 3 15 13 3 12 7 3 13 2 15 9 16 13 3 4 13 3 3 2
9 9 4 13 9 16 9 13 9 2
9 0 9 4 13 9 13 13 9 2
13 9 13 0 7 0 9 9 2 9 7 3 13 9
9 9 9 9 4 13 9 9 8 2
37 15 13 9 7 9 2 15 4 13 15 7 15 13 9 1 15 2 13 15 9 2 9 2 9 2 9 2 9 2 9 2 9 7 0 9 9 2
5 9 9 13 3 0
22 11 4 4 13 9 1 11 9 2 7 13 15 4 13 16 13 13 3 4 13 3 2
12 11 9 9 4 13 2 16 15 13 0 9 2
7 13 15 15 16 13 9 2
13 9 0 9 3 15 13 9 9 2 0 9 13 2
6 15 13 3 13 9 2
6 15 13 3 12 9 9
10 16 9 13 2 15 4 13 9 1 2
3 13 11 5
9 9 13 0 9 13 9 3 3 2
5 9 13 9 0 2
2 3 9
20 11 7 11 0 9 13 0 9 15 2 3 12 9 13 9 4 13 15 9 2
5 9 13 9 13 2
10 13 13 13 15 0 16 3 3 13 2
2 13 13
6 13 9 0 9 1 2
8 13 13 2 15 13 0 9 2
5 1 9 13 3 2
2 0 9
19 13 4 3 3 13 0 2 3 15 4 13 12 9 16 13 9 0 9 2
11 9 13 3 12 12 7 9 12 12 9 2
6 9 9 4 13 3 2
6 15 13 13 9 9 2
8 9 1 13 13 0 7 0 2
6 12 9 4 13 9 2
4 13 15 3 2
19 11 1 9 13 9 15 2 16 9 13 13 0 2 3 16 9 13 9 2
11 9 13 9 12 9 9 12 9 9 11 2
2 15 9
6 2 13 3 0 9 2
6 13 3 7 13 13 2
7 15 13 13 9 9 13 2
3 9 13 2
3 9 13 2
5 11 13 3 9 2
9 9 13 3 9 7 9 13 9 2
16 0 9 9 11 11 13 11 9 0 9 7 9 11 9 11 2
8 9 9 13 3 3 0 9 2
4 15 13 9 1
8 13 3 13 3 9 9 0 9
13 3 11 13 9 9 9 9 2 3 9 9 13 2
20 15 3 0 15 4 13 3 2 3 9 2 9 2 9 2 9 7 0 9 2
6 9 1 13 3 9 2
11 15 13 11 3 7 13 13 15 9 9 2
11 13 2 3 9 13 9 2 3 9 13 2
2 15 9
9 9 9 4 13 13 12 9 9 2
4 9 13 9 15
14 15 13 13 9 7 15 13 3 0 9 9 15 9 2
5 9 15 1 4 2
16 11 11 9 4 13 3 9 16 9 4 4 13 3 15 1 2
10 3 16 15 13 9 2 13 4 13 2
8 9 13 15 12 3 0 9 2
12 0 9 9 3 13 7 9 13 0 9 3 2
4 13 15 15 2
5 15 13 9 13 2
11 4 3 13 2 16 13 3 13 15 13 2
8 11 4 13 3 15 9 9 2
18 9 7 9 9 11 11 13 12 7 13 12 9 1 9 7 0 9 2
14 9 9 13 9 2 15 9 13 3 13 13 15 9 2
8 13 15 13 2 15 15 13 2
3 9 13 9
6 6 13 3 4 13 2
9 13 15 15 2 16 13 9 9 0
8 9 13 13 9 9 4 13 2
4 15 3 13 2
4 15 11 13 2
7 9 13 9 7 9 13 2
2 0 9
17 9 13 0 2 15 9 13 13 2 13 3 3 2 7 3 3 2
12 11 13 11 9 3 3 9 11 13 0 9 2
2 11 9
7 9 2 0 9 2 9 2
4 15 13 3 9
7 9 1 9 13 9 13 2
5 15 13 9 9 2
33 2 13 13 9 2 13 13 9 2 9 4 13 0 9 7 11 11 4 13 15 3 3 2 16 13 4 3 13 2 2 11 13 2
3 15 9 9
10 9 13 13 9 0 9 2 13 11 2
15 11 13 15 3 9 9 2 16 13 15 3 0 13 13 2
9 3 3 15 13 3 0 9 13 2
7 11 7 11 13 9 12 9
12 9 15 13 15 9 2 3 15 3 9 13 2
19 9 13 9 2 15 13 15 2 16 15 9 9 9 4 13 7 9 13 2
2 13 9
5 13 3 13 13 2
12 3 13 9 13 0 7 0 2 7 13 0 2
17 11 13 13 9 2 7 3 0 2 16 15 4 13 0 9 13 2
6 9 13 3 0 9 2
6 3 13 13 0 9 2
2 13 13
10 9 13 9 2 13 9 3 3 3 2
6 13 13 9 4 13 2
6 15 13 13 15 0 2
16 9 9 13 3 0 2 16 15 13 2 16 15 3 4 13 2
10 9 1 13 9 7 13 15 13 9 2
7 13 3 15 13 3 3 2
18 9 1 9 9 4 4 13 9 9 0 9 2 16 9 9 13 9 2
14 9 11 11 1 0 9 9 13 0 13 1 0 9 2
3 13 3 2
15 9 13 13 9 15 2 16 15 3 3 13 9 7 9 2
6 9 13 15 9 9 2
14 11 7 11 13 3 2 7 3 3 13 3 3 13 2
2 13 9
4 15 13 13 3
15 9 13 15 9 2 9 0 9 7 13 15 12 9 9 2
2 13 13
11 3 15 13 3 0 7 15 13 3 15 9
8 15 13 3 13 13 11 3 2
11 15 4 9 13 15 2 7 13 13 9 2
8 13 15 0 15 0 9 9 2
2 9 9
6 15 4 13 13 9 2
8 0 9 9 11 11 11 13 9
6 3 13 9 1 9 2
3 13 13 9
17 7 16 15 13 9 2 15 13 0 0 9 0 9 13 3 9 2
7 15 13 9 13 15 9 2
2 0 9
13 13 7 13 0 9 0 9 9 12 9 9 2 2
4 7 15 13 13
11 13 0 16 11 9 13 9 3 0 9 2
11 13 3 11 11 2 15 13 9 3 9 2
6 15 13 9 3 9 2
3 13 4 13
8 15 13 9 13 0 0 9 2
16 13 11 7 9 11 7 3 13 3 0 2 16 3 13 13 2
19 9 2 15 13 13 9 9 2 13 15 12 9 13 15 9 9 0 9 2
22 16 11 12 13 11 11 2 11 9 7 3 15 9 13 15 7 0 9 13 9 9 2
7 13 3 4 13 15 9 2
8 0 9 9 13 9 3 3 2
10 15 13 2 9 2 0 7 0 9 2
6 13 9 9 9 1 2
6 9 13 9 15 9 2
8 15 9 13 13 9 12 9 2
10 9 13 3 9 7 9 7 9 9 2
9 7 15 13 9 2 13 3 9 2
7 15 13 3 13 9 3 2
18 0 9 7 9 13 0 9 2 15 13 0 7 3 3 0 16 0 2
2 9 4
5 15 13 3 3 2
5 9 13 9 9 2
6 9 13 9 0 9 2
13 11 13 3 0 2 16 11 13 13 9 3 3 2
5 12 2 7 0 9
3 0 12 9
18 3 9 9 13 2 13 3 3 9 2 7 15 9 15 13 13 9 2
4 0 15 13 2
15 11 9 11 13 9 9 9 11 11 7 9 11 11 9 2
4 11 13 9 2
12 15 13 15 11 15 2 16 13 15 15 13 2
2 0 2
7 9 13 0 12 12 9 2
9 3 9 13 9 9 3 0 0 2
7 7 15 9 13 9 3 2
8 4 13 0 13 0 9 9 2
5 9 13 0 9 2
21 15 13 13 11 2 16 3 15 15 9 13 2 13 7 13 2 16 13 9 3 2
17 9 13 9 9 2 9 13 13 0 0 9 7 3 0 9 13 2
6 7 3 13 3 13 2
16 11 13 13 0 13 9 2 15 3 15 13 13 9 11 9 2
8 13 13 9 9 15 13 3 2
6 13 2 16 15 13 2
16 9 13 9 2 15 13 9 2 16 0 9 13 9 7 9 2
15 3 3 9 9 13 3 0 9 16 15 2 15 11 13 3
8 9 13 0 9 2 13 13 2
12 15 9 2 9 7 9 15 0 0 9 13 2
15 13 13 9 2 16 13 3 9 13 7 13 0 9 9 2
4 13 0 16 13
2 13 13
12 11 9 13 9 13 9 0 9 7 9 9 2
5 15 13 9 9 2
4 6 3 0 2
9 9 9 9 13 0 3 12 9 2
13 0 9 9 13 9 13 0 12 9 11 11 9 2
7 9 2 3 3 0 3 9
5 9 1 15 13 2
10 15 13 15 11 2 13 4 0 13 2
10 13 2 11 2 4 13 12 3 9 2
8 9 9 13 9 3 9 12 2
8 11 13 15 9 9 0 9 2
16 3 9 0 9 9 4 3 13 11 11 11 9 13 9 12 2
9 13 0 2 16 15 13 0 9 2
8 13 4 13 2 16 13 9 2
10 9 13 0 9 3 7 3 15 1 2
11 15 13 15 9 2 15 1 15 13 9 2
5 0 0 13 13 2
10 9 13 2 16 9 4 3 3 13 2
11 11 1 4 3 13 2 13 9 7 9 2
12 0 9 9 13 9 9 13 7 15 1 9 2
7 13 0 2 16 13 15 9
7 15 13 15 9 3 13 9
10 9 9 13 9 12 7 13 3 9 2
4 15 9 13 2
18 16 13 15 9 2 3 11 11 2 15 3 4 13 9 3 9 13 2
9 15 15 13 13 3 0 7 0 2
4 15 9 9 2
6 4 9 13 3 3 2
14 16 15 13 2 16 15 13 3 2 15 13 3 3 2
20 0 9 3 13 9 15 2 16 15 13 13 9 0 2 13 7 13 0 9 2
6 9 13 12 3 12 2
18 9 13 9 0 9 2 0 15 13 3 4 15 9 13 2 11 13 2
11 15 13 2 16 0 9 13 3 15 9 2
6 15 13 13 9 13 2
9 13 9 3 4 0 9 9 13 2
10 11 9 13 9 13 9 7 13 9 2
7 9 9 13 9 0 9 2
15 11 13 9 7 13 0 2 3 16 11 13 3 0 9 2
3 9 9 2
3 13 13 2
4 9 13 13 2
6 3 15 13 11 11 2
16 9 13 3 2 3 3 16 9 13 13 2 9 15 1 13 2
4 9 7 15 0
9 11 4 13 0 9 3 9 1 2
5 9 13 0 9 2
6 15 13 0 9 13 2
9 9 13 13 3 9 16 13 9 2
13 9 13 3 9 1 9 0 7 0 9 9 1 2
12 9 2 3 0 9 4 13 9 13 0 9 2
8 3 15 9 13 13 9 9 2
5 0 9 13 9 2
6 0 9 13 9 9 2
3 11 9 9
12 9 13 11 11 13 2 16 15 13 9 3 2
10 11 11 13 2 16 9 13 9 9 2
11 9 9 15 13 3 7 13 0 9 9 2
9 11 9 13 3 3 0 16 13 2
6 13 3 12 9 15 9
6 3 15 13 2 9 2
12 15 13 9 13 0 9 9 13 7 9 13 2
5 15 3 4 13 2
17 3 0 15 13 0 13 9 9 9 2 7 15 4 13 0 9 2
12 11 13 9 3 7 13 0 9 9 9 3 9
19 9 13 0 9 15 2 16 7 0 7 0 7 0 9 13 9 13 9 2
2 0 9
4 13 3 9 2
4 9 13 9 2
5 15 13 9 9 2
15 15 3 4 13 9 2 3 2 9 7 9 13 13 2 2
8 9 2 9 7 9 4 13 2
23 15 3 13 11 13 15 9 2 16 12 9 4 13 0 9 9 2 15 4 13 15 0 2
8 9 13 13 2 15 9 13 2
11 3 13 2 16 9 3 3 13 13 0 2
3 9 13 13
19 0 9 4 13 3 3 12 12 9 2 15 3 12 13 13 0 9 9 2
3 9 11 9
2 15 9
12 13 15 13 9 15 2 13 9 9 7 9 2
5 15 13 9 3 2
20 3 13 9 9 3 13 3 15 9 13 15 7 15 9 9 3 3 11 9 2
18 9 4 13 3 0 2 16 9 4 13 7 13 9 9 13 9 1 2
3 3 7 3
2 0 9
5 0 9 13 3 2
2 13 13
4 9 13 3 2
12 13 9 3 3 13 15 13 3 9 1 9 2
4 9 13 9 2
11 11 13 13 13 2 15 9 9 4 13 2
8 9 13 3 9 11 11 9 2
15 15 13 3 0 9 7 15 9 4 13 9 9 1 9 2
14 0 9 9 13 9 2 7 13 15 9 9 13 9 2
10 9 3 13 13 9 13 0 9 9 2
13 9 12 13 11 12 9 2 0 9 9 13 12 2
2 9 9
2 9 9
2 3 2
46 3 15 13 3 0 16 3 11 13 3 3 3 15 13 11 9 15 13 3 0 9 15 13 3 13 3 13 13 15 13 3 13 16 2 11 3 13 3 13 3 9 7 15 13 15 9
5 9 13 9 13 2
6 13 15 13 15 9 2
13 13 9 2 16 13 0 0 9 13 3 15 1 2
3 13 15 2
8 3 13 9 13 2 3 9 2
12 9 9 13 2 16 9 9 13 9 9 9 2
2 0 9
6 7 13 15 13 9 2
4 3 9 0 2
4 3 15 13 2
21 16 11 13 9 13 3 13 13 2 9 9 13 0 9 0 11 11 2 9 2 2
12 9 13 3 0 9 2 16 15 13 15 0 2
11 11 4 13 12 9 3 16 13 11 13 11
8 3 15 11 9 15 13 13 2
11 9 9 4 13 3 0 7 0 16 9 2
6 13 15 11 15 9 2
2 3 3
9 15 13 9 3 9 0 9 1 2
7 13 13 16 13 9 13 3
16 15 13 13 11 1 15 9 16 15 13 2 13 15 3 3 2
14 9 13 15 0 9 7 15 3 15 16 0 0 9 2
9 13 3 9 15 0 0 9 11 2
12 3 15 13 13 13 2 16 9 13 15 13 2
9 9 1 11 13 2 16 9 13 2
8 9 13 9 9 11 11 11 2
7 11 4 13 7 13 9 2
16 3 13 0 9 7 9 2 3 0 16 15 4 4 15 13 2
11 9 9 4 13 12 12 7 9 12 12 2
2 11 9
12 0 9 13 0 9 2 9 7 9 7 9 2
12 13 4 13 0 9 2 16 9 13 15 9 2
3 13 9 2
11 0 9 13 11 9 9 13 9 9 9 2
17 13 9 9 13 12 9 2 15 13 7 9 13 13 12 12 9 2
8 12 9 1 9 3 13 12 2
2 9 9
11 13 4 3 13 9 16 15 13 3 15 9
3 0 9 9
66 9 9 2 13 12 9 9 12 2 9 0 9 2 11 2 7 0 9 13 9 9 2 11 2 9 13 9 9 7 13 9 13 15 9 9 13 9 9 9 1 13 9 9 7 9 12 9 0 7 0 9 2 13 9 12 12 2 2 11 9 0 9 2 2 12 2
49 11 9 9 2 15 13 9 11 9 9 2 13 9 9 9 13 9 13 13 9 7 9 9 12 9 9 12 13 9 9 12 2 12 2 2 7 3 15 12 9 12 7 12 9 2 7 13 0 2
17 2 12 2 9 9 12 2 12 2 13 7 13 0 9 13 9 2
50 9 9 13 13 9 13 9 2 15 9 4 13 13 9 9 7 13 9 13 9 4 13 13 9 13 13 9 9 12 7 0 0 9 9 2 0 9 2 11 2 7 0 9 13 9 9 2 11 2 2
25 2 12 2 11 13 12 9 9 12 13 9 2 16 9 13 11 9 13 9 9 11 11 11 11 2
10 9 4 9 13 13 9 9 12 1 2
22 9 4 3 13 9 0 9 2 15 13 9 9 13 9 12 12 13 12 9 0 9 2
27 2 12 2 13 9 13 9 12 12 9 0 2 7 15 4 15 1 13 7 9 12 9 0 4 13 3 2
15 16 9 4 13 13 9 2 9 4 13 12 9 9 9 2
24 2 12 2 11 13 12 9 9 12 13 9 2 16 9 12 9 0 13 12 9 13 9 13 2
15 9 4 13 11 9 9 13 9 1 13 9 15 0 9 2
14 9 13 9 12 9 0 13 12 9 13 9 13 9 2
8 9 13 9 4 15 1 13 2
18 2 12 2 15 9 12 13 2 11 7 11 13 9 4 3 13 9 2
21 15 9 4 13 13 9 9 2 7 15 4 13 9 9 12 2 12 2 9 0 2
11 15 9 4 15 1 13 9 12 9 0 2
11 2 12 2 9 12 4 15 1 13 3 2
18 2 12 2 15 9 13 9 13 9 7 9 9 13 0 9 9 0 2
5 4 13 15 9 2
2 12 9
39 0 13 11 13 9 9 12 12 9 12 9 0 9 13 9 9 9 12 7 0 0 9 9 2 0 9 2 11 2 7 0 9 13 9 9 2 11 2 2
41 0 13 11 13 2 9 12 12 9 12 9 0 9 13 9 9 9 13 9 12 7 0 0 9 9 2 0 9 2 11 2 7 0 9 13 9 9 2 11 2 2
2 12 9
5 13 9 12 3 2
10 12 2 13 9 0 15 9 9 0 2
10 12 2 13 9 0 15 9 9 0 2
2 12 9
14 9 4 13 3 13 9 13 9 2 9 7 0 9 2
2 12 9
7 15 9 4 13 15 9 2
7 13 11 12 9 9 12 2
6 9 1 11 11 9 9
27 2 8 2 2 11 9 9 2 11 12 12 12 0 9 9 9 2 11 9 2 11 9 7 9 7 9 9
3 0 9 9
7 9 0 9 9 9 11 9
1 9
3 0 9 12
6 0 13 0 9 9 12
6 0 1 0 11 9 12
3 0 9 12
2 11 12
2 0 9
14 0 9 7 0 9 9 9 13 3 9 13 11 9 2
11 9 9 4 4 13 9 7 9 13 9 2
14 9 13 3 0 9 3 0 2 7 3 15 0 9 2
25 9 9 4 13 9 7 9 13 9 1 9 2 7 9 13 13 2 16 9 13 3 4 13 13 2
18 16 9 9 2 9 7 0 9 13 15 2 9 13 13 0 0 9 2
9 15 9 13 9 15 1 13 9 2
17 11 13 7 13 0 9 9 9 4 13 9 3 0 9 0 9 2
13 9 12 9 7 9 9 13 13 9 13 0 9 2
16 9 12 13 9 13 9 7 13 9 13 3 9 9 7 9 2
14 9 13 9 2 9 7 9 13 9 9 13 0 9 2
23 0 9 9 7 9 9 13 13 9 9 2 11 11 11 11 11 11 11 2 13 9 12 2
21 9 12 9 12 13 9 13 11 9 13 9 13 3 0 9 7 9 13 11 9 2
21 11 9 1 0 9 13 9 4 13 9 11 0 9 2 15 13 0 9 7 9 2
22 9 7 9 9 13 0 9 12 0 9 2 15 13 0 9 9 9 13 0 11 9 2
14 11 9 9 13 13 0 9 13 9 1 9 12 9 2
15 9 13 0 9 0 9 0 9 13 9 9 13 11 9 2
13 0 9 13 2 16 9 13 9 4 13 0 9 2
8 9 13 3 0 11 9 9 2
13 9 3 7 3 13 9 9 13 3 11 9 9 2
19 9 13 7 13 9 9 2 15 13 9 2 9 7 9 7 9 0 9 2
14 9 13 3 9 9 2 16 9 9 4 13 3 9 2
17 0 9 7 9 13 13 9 9 13 13 9 2 15 13 9 9 2
14 9 3 13 9 13 9 2 9 7 9 0 9 9 2
8 11 9 13 0 9 9 9 2
41 9 13 9 2 9 9 7 0 9 15 2 9 2 9 13 9 2 15 13 9 7 9 0 9 2 16 4 13 9 2 0 9 7 15 0 9 13 13 0 9 2
28 13 11 0 9 9 12 7 11 9 0 9 9 12 13 0 9 2 15 13 9 15 9 7 15 13 9 9 2
6 9 13 0 0 9 2
7 11 13 9 9 0 9 2
37 0 9 9 9 13 9 2 11 2 4 13 0 9 13 0 9 9 7 13 9 7 9 2 9 7 9 7 15 9 0 9 9 7 0 9 9 2
15 9 4 13 3 9 2 7 13 13 9 13 4 13 9 2
14 9 4 13 9 12 9 1 0 9 9 0 9 3 2
11 15 9 13 0 9 9 9 13 0 9 2
28 9 9 13 11 9 9 2 7 3 13 9 2 15 4 13 9 9 9 13 0 9 2 15 13 9 9 9 2
17 9 9 2 15 13 11 9 9 12 2 13 3 13 9 0 9 2
7 3 11 9 13 15 9 2
15 15 9 13 9 0 9 9 9 13 9 13 0 11 9 2
20 9 9 13 9 0 9 2 15 0 9 13 3 2 7 0 15 13 11 9 2
17 9 13 9 11 3 13 9 7 13 0 9 7 0 7 11 9 2
7 9 13 13 0 0 9 2
16 3 13 0 9 2 15 13 11 9 13 7 0 9 0 9 2
5 0 13 0 9 9
10 0 9 13 9 7 11 7 9 9 2
18 13 9 2 15 13 9 9 2 13 9 9 2 9 7 13 11 9 2
24 9 13 13 0 13 9 4 13 9 2 7 9 4 13 13 9 7 9 0 9 7 9 3 2
11 9 13 3 0 7 11 9 9 0 9 2
15 15 9 4 13 9 9 7 13 3 9 9 7 9 9 2
19 0 2 9 13 0 0 9 2 15 9 7 9 7 9 9 4 13 2 2
6 0 9 2 11 9 2
12 13 13 9 9 13 0 9 13 9 13 9 9
9 13 0 9 2 15 0 9 13 3
19 13 9 3 9 2 9 7 0 9 9 3 9 9 2 16 15 13 3 9
7 13 13 9 9 7 9 9
7 13 0 9 0 9 9 9
10 13 9 7 0 9 9 9 2 9 3
11 13 9 9 1 3 13 9 0 9 9 2
25 13 9 0 9 2 3 9 7 0 9 2 15 9 13 0 9 9 9 7 9 7 0 7 0 9
18 13 9 7 9 2 15 13 0 9 13 9 9 9 9 7 9 9 2
9 0 2 9 13 11 9 9 9 2
6 0 9 2 11 9 2
13 13 9 9 9 7 15 13 0 9 9 13 9 2
18 3 13 13 2 16 9 13 0 7 0 9 7 13 15 7 13 15 2
10 13 0 9 9 9 13 9 0 0 9
12 13 13 0 9 2 15 13 0 9 11 9 2
21 0 2 9 13 0 9 9 2 15 13 0 9 9 13 3 7 3 13 9 9 2
6 0 9 2 11 9 2
8 13 0 9 2 15 13 9 9
9 13 9 9 13 9 9 7 9 2
16 13 9 7 9 9 9 13 9 2 16 4 13 9 9 7 9
16 13 3 13 9 1 0 9 2 15 13 9 9 2 9 7 9
14 13 9 2 9 9 7 9 9 9 2 15 13 3 9
24 13 9 9 13 9 9 9 9 9 3 3 13 2 16 9 9 13 9 13 13 15 13 13 9
13 13 9 13 9 13 9 7 0 9 7 15 9 2
12 13 9 9 1 3 13 9 7 15 9 9 2
10 13 9 2 15 0 9 13 9 9 9
9 13 9 13 9 2 15 13 9 9
14 13 9 9 7 3 13 0 9 9 9 13 9 9 2
23 0 2 9 13 13 1 9 13 9 9 2 9 7 9 2 9 4 13 9 13 15 9 2
6 0 9 2 11 9 2
15 13 9 9 9 3 13 1 9 9 9 7 9 7 9 9
27 13 0 9 9 9 7 15 9 2 16 15 13 9 0 9 9 2 9 2 9 2 0 9 2 9 7 9
14 13 0 9 2 15 13 9 0 9 7 0 9 13 9
21 13 9 9 13 9 13 7 9 2 9 2 9 2 0 7 0 13 9 7 15 9
13 13 9 9 9 7 9 2 9 7 9 7 9 2
11 12 0 9 9 11 13 0 9 9 2 0
38 11 9 9 9 0 9 11 9 7 9 9 9 0 9 9 2 9 7 9 9 11 13 0 9 9 2 12 2 12 2 12 2 2 9 2 0 9 2
16 11 9 2 15 2 13 9 9 0 9 2 12 2 12 2 2
17 2 13 9 0 9 13 9 9 9 11 9 7 9 2 12 2 2
10 2 13 9 9 13 9 2 12 2 2
10 2 13 9 9 9 12 9 12 9 2
7 2 13 9 9 12 9 2
15 2 13 9 9 2 9 7 9 9 0 9 2 12 2 2
6 0 13 0 9 3 2
10 0 13 9 13 9 9 9 7 9 2
6 13 9 12 2 12 2
6 13 3 13 0 9 2
6 13 3 13 0 9 2
13 9 12 9 9 2 12 12 2 2 9 2 9 2
21 11 9 9 9 12 13 9 9 9 4 13 9 12 2 11 9 9 3 9 9 2
36 11 9 7 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 9 9 9 13 9 9 2 9 2 9 12 9 2 11 9 0 9 2
58 11 9 7 11 9 9 2 15 13 9 11 9 9 7 3 15 12 9 12 9 2 13 9 9 9 2 12 2 2 13 9 9 7 9 9 2 12 2 2 4 13 9 9 2 13 9 12 9 13 9 2 12 2 2 7 13 0 2
19 2 12 2 13 0 13 9 0 9 2 16 9 13 9 13 9 0 9 2
31 2 12 2 11 13 9 12 9 9 12 0 9 15 0 9 13 9 9 2 15 13 0 0 9 9 0 9 13 9 9 2
18 15 9 13 9 12 13 11 9 7 15 3 13 9 9 2 12 2 2
14 2 12 2 11 9 13 3 3 11 9 9 0 9 2
14 2 12 2 11 9 13 0 9 9 9 7 9 9 2
17 2 12 2 9 4 13 11 9 7 13 9 13 15 9 13 15 2
40 2 12 2 13 3 13 9 9 9 9 12 9 9 12 13 9 9 2 9 2 9 12 2 12 2 15 9 11 9 0 7 13 3 9 0 9 13 0 9 2
33 2 12 2 15 9 7 11 9 13 9 7 15 9 9 2 13 15 4 13 3 2 16 15 9 0 9 13 15 9 15 9 9 2
31 2 12 2 0 9 13 3 13 0 7 0 9 2 15 1 11 9 1 13 0 13 0 7 0 9 7 0 7 0 9 2
18 2 12 2 9 3 13 0 13 9 9 0 9 9 15 9 9 9 2
19 2 12 2 0 7 0 9 9 9 7 9 9 13 0 13 0 9 9 2
43 2 12 2 9 9 9 13 4 4 13 3 11 9 12 9 12 9 2 13 15 13 2 16 9 13 13 9 9 7 15 9 13 9 7 15 9 9 7 0 9 7 9 2
48 2 12 2 9 9 2 9 7 9 7 9 13 9 13 0 9 9 2 15 13 15 9 9 9 13 9 2 13 0 7 0 9 7 9 7 9 2 7 15 9 9 4 13 2 3 13 9 2
23 2 12 2 9 9 9 13 13 0 13 0 9 9 0 9 2 7 0 13 9 9 0 2
19 2 12 2 9 9 7 15 13 0 9 0 9 13 0 13 3 9 1 2
18 2 12 2 11 9 12 9 13 9 13 2 16 9 9 13 3 0 2
29 15 9 13 13 3 13 9 9 9 9 9 12 9 9 12 13 9 9 2 9 2 9 12 12 9 2 12 2 2
21 2 12 2 15 9 4 13 9 9 13 9 2 16 15 4 13 13 9 1 9 2
21 2 12 2 15 9 13 9 13 3 13 3 9 7 11 9 9 9 0 9 9 2
35 2 12 2 15 9 16 11 9 3 9 13 3 15 9 15 9 9 2 15 9 2 9 2 9 12 13 13 2 9 9 13 13 15 9 2
5 4 13 15 9 2
2 12 9
9 13 9 2 9 2 9 12 3 2
33 12 2 13 9 9 3 2 2 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 7 15 9 9 13 9 9 9 2 2
7 12 2 13 12 9 3 2
3 2 12 9
20 15 9 13 3 11 9 13 9 7 15 9 9 13 9 7 13 0 0 9 2
11 15 3 13 15 9 9 9 0 9 2 2
7 12 2 13 12 9 3 2
3 2 12 9
5 0 15 9 13 2
14 9 2 2 9 9 2 9 2 15 13 3 13 9 2
26 9 2 2 9 9 9 2 9 9 2 15 13 9 2 9 2 9 12 9 0 9 13 3 13 9 2
21 9 2 2 9 13 9 2 9 7 9 2 15 13 9 3 13 9 1 13 9 2
27 9 2 2 9 2 2 13 15 4 3 13 2 11 9 12 9 12 9 13 9 0 7 13 7 0 9 2
12 9 2 2 0 9 2 0 9 13 0 9 2
47 9 2 2 11 9 2 15 0 9 13 9 9 11 12 9 9 12 13 9 2 7 11 9 2 0 16 15 13 13 11 12 9 9 12 2 7 11 12 9 9 12 13 11 9 13 9 2
21 9 2 2 11 9 2 11 12 9 9 12 13 15 0 9 13 9 9 13 9 2
21 0 15 9 13 9 2 15 13 13 12 9 2 13 15 16 11 9 13 9 2 2
7 12 2 13 12 9 3 2
3 2 12 9
19 0 9 7 15 9 13 9 9 9 9 13 15 0 9 13 11 9 9 2
56 0 9 2 9 2 9 12 12 9 13 9 13 2 15 9 16 15 13 9 13 9 2 13 2 16 9 9 9 4 13 0 9 1 2 15 13 13 2 16 15 9 13 9 13 0 15 2 15 15 13 13 15 9 3 2 2
6 12 2 13 9 3 2
4 2 12 9 9
63 9 2 15 9 9 9 4 13 11 9 12 9 12 9 3 2 3 16 9 4 3 13 15 9 9 2 15 13 9 9 9 2 4 13 9 2 15 13 9 0 9 9 7 9 13 9 2 15 13 0 9 9 7 9 2 15 4 13 3 9 9 0 2
8 9 4 13 9 9 13 2 2
6 12 2 13 12 9 2
7 12 2 13 12 9 3 2
3 2 12 9
43 0 9 9 9 4 13 7 3 12 9 13 15 2 16 9 13 0 9 9 4 13 2 13 9 2 15 13 0 9 0 0 9 7 15 13 9 15 2 15 15 4 13 2
23 0 9 0 9 4 13 3 12 0 9 13 9 9 9 1 2 13 3 13 12 9 9 2
48 0 9 9 13 13 9 9 2 7 15 4 13 9 9 9 9 9 13 0 9 2 7 15 4 13 3 3 11 9 12 9 13 9 7 16 9 2 15 9 13 2 13 13 9 13 9 2 2
7 12 2 13 12 9 3 2
3 2 12 9
48 0 15 9 9 13 9 9 4 13 2 16 9 13 15 9 2 9 7 11 9 13 9 3 13 2 9 0 9 7 15 9 13 9 13 9 3 13 9 9 13 9 7 9 13 9 0 9 2
12 15 9 9 9 9 9 4 13 9 13 9 2
20 0 9 7 9 13 4 13 9 9 2 13 15 9 9 7 11 9 9 9 2
23 0 3 12 9 13 9 1 15 9 9 4 13 9 13 7 13 9 9 15 9 3 9 2
19 2 0 9 13 9 9 9 9 9 7 9 9 2 16 0 9 13 13 2
35 2 0 9 13 9 9 9 9 9 9 2 9 7 9 9 7 9 2 16 0 9 0 9 4 13 9 9 7 9 4 13 15 1 9 2
13 2 0 9 13 9 9 9 9 9 13 9 9 2
36 0 16 9 9 9 13 15 9 2 12 7 12 9 13 9 3 13 9 4 13 15 2 15 13 15 9 2 13 9 9 9 3 13 0 9 2
25 16 9 0 9 9 13 15 9 2 12 7 12 9 13 3 9 2 9 7 15 1 13 9 2 2
7 12 2 13 12 9 3 2
3 2 12 9
26 9 13 3 12 9 13 15 2 16 9 2 9 2 9 12 2 12 2 13 13 2 9 15 9 9 2
26 9 13 3 9 13 11 9 9 13 9 13 9 0 9 7 0 9 2 11 2 9 13 9 1 2 2
6 12 2 13 9 3 2
10 2 9 9 9 9 9 7 15 9 9
17 15 9 13 9 9 9 7 11 9 13 9 9 9 9 13 9 2
5 9 9 7 9 9
11 9 9 7 9 9 9 13 4 3 13 2
20 3 12 0 9 0 2 0 9 0 9 2 9 9 9 9 13 4 13 9 2
21 15 9 0 9 9 9 4 13 9 1 13 2 13 15 4 13 3 7 3 3 2
1 9
27 16 9 13 7 13 2 9 9 4 13 9 0 0 9 9 12 9 13 15 2 16 9 13 9 4 13 2
16 9 15 9 4 13 3 12 0 9 2 0 9 0 9 2 2
4 9 9 13 9
27 9 13 9 9 13 9 2 3 16 15 4 13 15 9 13 9 9 9 7 16 0 9 13 13 0 13 2
17 9 9 13 9 9 9 13 12 0 9 2 0 9 0 9 2 2
17 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 9 9
46 11 9 9 2 15 13 9 11 9 9 7 3 15 12 9 2 13 9 9 13 9 2 12 2 13 9 11 9 9 2 12 2 2 13 9 9 7 9 9 2 12 2 2 7 13 2
43 16 2 12 2 4 13 15 13 0 9 13 9 9 4 13 9 0 2 0 2 3 7 3 13 2 0 9 9 13 9 13 9 9 9 7 9 7 15 9 13 9 9 2
67 2 12 2 0 9 9 13 9 9 9 12 9 9 12 13 9 9 12 2 12 2 13 13 0 9 13 9 2 15 13 13 0 3 2 16 0 9 13 2 0 9 13 9 13 0 9 15 1 2 13 9 0 7 0 9 2 13 15 13 0 9 15 9 13 9 9 2
17 2 12 2 13 3 13 0 0 7 9 7 9 13 9 13 9 2
49 2 12 2 9 12 13 9 4 15 1 13 2 16 13 3 15 2 16 9 0 9 0 9 7 9 13 15 9 16 0 9 2 7 16 13 9 9 7 9 13 9 1 13 15 9 13 9 9 2
35 2 12 2 9 3 0 9 9 0 9 9 13 9 2 15 4 13 3 3 9 2 16 9 13 15 9 0 9 9 13 9 7 9 9 2
43 2 12 2 9 9 12 9 9 12 13 9 9 2 9 2 9 12 2 12 2 13 9 15 9 9 2 3 15 9 2 15 13 0 9 9 2 13 13 9 9 7 9 2
15 2 12 2 0 13 9 9 9 13 3 9 0 9 9 2
9 2 12 2 9 0 9 4 13 2
13 2 12 2 9 9 4 13 9 3 0 9 9 2
20 2 12 2 13 3 13 13 9 15 9 9 7 15 9 0 7 0 9 2 7
18 2 12 2 9 12 2 12 2 13 9 4 13 0 9 12 9 3 2
7 9 4 13 13 15 9 2
5 4 13 15 9 2
2 12 9
3 9 7 9
27 0 15 9 4 13 9 9 2 15 13 9 13 2 0 9 13 9 9 13 9 9 7 15 9 13 9 2
13 0 15 9 13 9 9 3 1 0 9 13 9 2
19 9 2 9 13 9 9 2 15 0 9 7 9 13 0 0 9 13 9 2
26 9 2 9 2 9 7 0 9 7 9 13 9 2 3 1 0 9 7 3 9 13 9 13 9 9 2
27 15 9 13 9 13 15 9 9 1 0 9 13 9 9 2 15 9 7 0 0 9 13 13 0 9 0 2
21 15 9 13 4 9 9 13 3 12 9 13 0 9 0 13 9 9 3 12 9 2
2 12 9
1 9
4 15 9 13 2
16 2 2 9 9 2 15 9 9 2 15 13 9 13 9 9 2
32 2 2 9 9 2 9 9 2 15 15 9 13 9 7 15 13 3 9 7 9 9 9 7 9 7 9 9 13 9 9 9 2
22 2 2 9 13 9 9 2 3 7 3 9 13 9 9 2 9 2 9 2 9 2 2
33 2 2 9 13 9 9 2 9 13 0 9 9 2 9 2 7 9 9 9 2 7 9 2 0 9 2 7 9 2 0 9 2 2
12 2 2 9 2 3 7 3 9 13 0 9 2
25 2 2 9 2 0 9 9 2 15 4 3 7 3 13 15 16 0 9 9 2 3 9 2 9 2
16 2 2 9 2 9 13 9 9 2 15 4 13 9 9 13 2
32 2 2 9 2 9 13 9 9 2 15 13 13 9 7 15 4 13 3 2 16 9 15 9 7 0 9 15 9 9 13 9 2
11 2 2 9 2 9 9 7 15 13 9 2
15 2 2 9 2 9 13 9 2 15 4 13 0 7 9 2
11 9 2 15 4 13 9 2 13 15 9 2
21 2 2 13 2 9 0 9 13 9 9 9 9 1 15 2 13 0 9 9 9 2
45 16 9 13 0 9 9 9 7 9 2 0 9 2 7 9 2 0 9 2 2 15 9 9 2 9 7 9 2 7 9 7 9 4 13 0 9 2 9 9 13 9 9 9 3 2
13 2 2 9 2 9 9 0 9 13 9 0 9 2
20 16 9 13 9 13 9 7 0 7 9 2 9 9 13 9 7 9 9 9 2
26 2 2 0 0 9 2 9 9 0 9 13 1 13 7 0 9 2 7 9 9 2 7 9 0 9 2
16 2 2 11 2 9 9 2 15 13 9 13 9 9 9 9 2
2 12 9
1 9
8 0 9 13 0 9 13 9 2
6 9 2 9 13 9 2
6 9 2 9 13 9 2
6 9 2 9 13 9 2
18 0 15 9 13 0 9 2 15 9 7 15 9 13 9 9 13 9 2
15 0 9 9 13 9 13 9 13 13 9 9 0 9 9 2
14 0 9 9 9 7 9 9 13 12 9 13 9 13 2
2 12 9
2 9 9
26 9 9 7 9 4 13 3 2 16 9 13 0 9 13 9 13 9 2 15 13 9 9 9 0 9 2
8 9 13 12 9 13 9 13 2
2 12 9
3 9 9 11
27 0 9 4 13 11 3 12 9 13 7 9 9 13 9 13 7 3 13 9 9 13 9 2 9 7 9 2
17 9 13 13 15 0 9 13 9 2 15 4 3 13 3 0 9 2
22 0 3 12 9 13 9 7 13 0 9 13 9 9 13 9 13 12 9 13 9 13 2
11 0 9 13 12 9 13 15 0 9 9 2
8 0 9 13 9 12 0 9 2
43 0 9 4 12 9 9 12 13 7 12 9 3 13 9 0 9 13 9 9 13 5 9 12 2 12 2 12 7 12 9 7 5 9 12 7 12 9 13 9 9 13 9 2
4 13 9 13 2
10 2 0 9 9 2 9 9 0 9 2
8 2 0 9 9 2 0 9 2
36 0 3 12 9 13 9 9 13 12 9 13 9 13 3 16 0 9 13 0 0 9 7 0 7 0 9 9 9 9 13 12 7 12 9 3 2
2 12 9
2 9 9
24 9 9 13 0 9 9 13 9 2 3 13 13 9 9 7 9 2 13 12 9 13 9 13 2
2 12 9
1 9
14 0 3 0 9 9 9 9 9 13 11 9 13 9 2
11 13 9 13 11 3 9 13 9 0 9 2
33 9 9 9 13 7 13 9 9 9 9 13 9 9 2 9 2 9 12 12 9 12 9 3 2 12 2 2 11 9 0 9 2 11
2 13 9
3 9 9 2
18 9 2 15 13 9 2 9 2 9 12 12 9 12 9 9 9 13 9
23 2 8 2 2 11 9 9 2 11 12 12 12 0 0 9 11 9 9 9 2 9 13 2
2 0 9
31 15 0 9 9 13 13 15 0 9 13 9 11 9 9 2 11 2 11 11 11 2 9 7 15 0 9 7 9 13 9 2
24 11 13 9 12 9 7 9 2 16 4 13 2 16 9 7 9 15 9 13 9 9 4 13 2
33 15 9 13 13 9 7 9 0 9 0 2 0 7 0 9 13 7 13 3 9 3 13 13 9 7 13 9 7 0 9 13 9 2
19 15 9 11 13 9 13 0 9 7 9 2 15 9 11 9 13 7 13 2
27 16 9 9 13 9 12 2 13 9 13 0 9 7 13 15 0 9 9 9 15 2 3 9 13 0 13 2
4 0 0 0 9
25 11 9 13 3 9 12 0 9 7 9 13 9 2 3 0 13 13 9 9 9 0 11 3 3 2
6 9 13 9 9 12 2
23 11 9 12 13 9 9 9 9 13 2 13 0 9 9 2 9 7 9 13 9 9 2 2
8 15 3 11 13 9 9 12 2
15 9 1 13 2 16 9 9 13 0 9 9 13 0 9 2
20 11 9 12 13 9 13 11 9 7 13 4 2 13 9 13 0 9 9 2 2
32 3 9 2 15 13 12 2 13 9 9 9 13 11 9 2 16 2 11 9 7 9 9 13 9 4 13 9 15 9 0 9 2
22 0 0 13 13 0 9 9 2 9 7 9 15 0 9 9 7 13 15 9 3 2 2
3 0 0 9
23 9 7 11 9 7 9 13 3 9 7 9 0 9 2 15 11 0 9 4 13 9 13 2
15 9 13 3 9 12 13 9 7 13 11 9 12 13 9 2
29 3 2 16 15 0 9 13 9 13 0 9 3 9 2 9 13 13 0 13 3 2 16 15 13 3 13 3 13 2
27 3 0 9 13 7 13 9 2 15 4 13 3 9 2 13 3 0 11 9 7 9 2 7 9 7 9 2
26 0 9 7 9 0 7 0 9 7 9 7 0 11 13 4 13 3 0 2 0 7 0 9 7 9 2
12 11 7 9 9 0 9 13 3 3 3 9 2
16 3 11 7 9 4 3 3 13 3 9 9 7 9 13 9 2
19 15 9 9 13 0 9 2 15 9 15 9 13 7 15 13 0 0 9 2
17 0 13 3 0 2 13 9 7 9 13 0 2 0 7 0 9 2
24 3 13 9 9 9 9 7 0 9 13 9 9 13 15 9 2 7 0 9 9 13 3 3 2
5 0 11 9 9 9
21 15 9 13 11 9 7 15 9 2 9 7 9 2 15 9 13 0 0 9 13 2
4 12 9 7 9
18 15 9 11 13 9 13 12 0 9 2 11 2 8 8 8 2 9 2
14 9 13 9 9 2 16 15 13 9 7 9 7 9 2
16 0 0 9 13 4 3 13 9 2 3 15 13 11 9 9 2
9 15 15 13 13 11 9 9 12 2
32 0 9 13 9 9 7 9 2 9 7 9 9 7 15 9 13 9 2 9 7 9 9 13 9 2 7 9 0 9 0 9 2
14 9 13 3 3 2 3 3 2 16 9 9 13 3 2
13 9 12 13 0 9 9 9 7 9 13 9 9 2
2 12 9
8 9 7 9 13 0 9 3 2
34 15 0 9 2 15 13 9 9 9 7 15 9 2 13 13 9 9 7 9 0 2 0 9 13 9 7 9 13 9 9 13 9 1 2
27 9 9 13 9 12 9 1 12 12 9 2 7 9 12 9 9 13 12 12 2 15 13 9 13 9 12 2
18 3 13 9 12 0 9 7 13 9 13 9 9 9 7 9 9 1 2
6 12 9 7 9 0 9
30 11 0 9 1 15 9 9 13 13 9 2 9 7 9 3 9 0 2 0 7 0 9 9 7 9 0 9 7 9 2
23 15 13 9 13 13 3 7 13 13 3 13 13 9 7 13 3 7 13 13 13 0 9 2
15 11 13 12 15 13 9 2 3 9 7 9 7 3 9 2
30 15 13 9 9 2 9 2 9 7 9 13 9 9 7 13 0 9 0 9 13 9 9 7 0 9 9 0 9 1 2
10 9 9 13 0 9 11 9 7 9 2
8 11 9 13 9 13 0 9 2
30 13 15 9 0 9 0 9 13 9 2 9 7 9 2 11 9 0 9 9 12 3 15 9 4 15 9 9 13 3 2
1 9
15 0 9 9 13 9 3 13 3 13 0 9 11 9 9 2
20 9 12 13 9 13 9 7 9 2 16 9 13 0 9 13 9 9 3 9 2
7 15 13 3 9 7 9 2
16 9 4 3 13 3 0 2 3 15 9 9 13 3 9 9 2
30 0 9 4 9 12 9 1 13 9 3 12 12 9 2 7 3 4 13 0 9 13 9 7 0 9 0 9 7 9 2
13 9 13 9 9 13 3 13 13 0 9 9 9 2
35 13 0 2 16 9 4 3 13 3 9 2 16 11 9 4 13 0 9 0 7 0 9 7 0 9 9 2 9 13 9 7 9 3 9 2
3 9 7 9
12 11 4 13 0 15 9 7 9 7 13 9 2
54 9 4 13 9 12 9 9 9 0 9 2 9 11 0 9 9 9 12 13 9 9 9 7 9 7 13 9 13 9 2 9 9 9 9 12 13 9 2 15 13 9 9 9 9 7 15 9 13 9 2 7 15 9 2
26 13 9 9 12 0 9 13 3 3 0 9 9 9 9 9 3 13 0 9 9 7 0 9 9 9 2
42 16 13 3 3 0 13 11 9 9 9 9 2 4 13 2 16 0 9 4 13 0 9 2 15 13 9 9 9 3 13 0 7 0 9 2 15 9 4 13 9 9 2
3 9 7 9
10 0 9 0 9 4 13 9 9 13 2
18 0 9 15 4 13 13 0 9 13 0 9 7 13 9 9 9 9 2
13 0 9 4 13 9 9 9 0 7 0 0 9 2
13 9 4 13 13 3 15 11 9 13 9 7 9 2
21 15 13 3 4 13 9 9 2 15 13 3 2 16 11 4 13 9 7 13 9 2
21 11 9 9 9 13 15 9 0 2 16 3 15 15 9 4 2 3 2 9 13 2
12 15 1 9 9 9 13 3 4 13 13 9 2
21 9 9 13 3 15 2 16 9 4 13 9 3 0 2 3 15 0 9 13 9 2
15 15 9 13 3 15 9 13 11 9 7 13 15 9 0 2
2 12 9
16 9 12 9 13 3 0 9 2 15 0 11 4 13 9 13 2
12 12 0 9 13 0 9 9 7 9 0 9 2
28 3 0 9 0 9 7 9 7 15 9 13 9 7 9 7 0 9 13 0 9 2 3 9 9 13 3 0 2
23 3 9 4 13 0 9 7 15 3 13 3 2 15 13 7 9 7 9 9 0 9 9 2
27 9 9 2 13 12 9 9 12 2 9 7 9 7 9 9 9 3 13 9 9 12 7 12 9 2 12 2
157 11 9 9 2 15 13 9 11 9 9 2 13 9 9 9 9 3 12 9 9 12 13 9 9 12 2 2 2 0 16 15 13 3 13 9 9 12 2 2 2 7 3 15 12 9 9 2 13 9 9 7 9 9 9 3 12 9 9 12 13 9 9 12 2 2 2 0 16 15 13 3 13 9 9 12 2 7 3 15 12 9 9 7 13 2 16 0 7 0 9 9 9 9 12 9 0 7 9 12 9 0 4 13 3 2 16 0 9 9 7 0 9 7 9 9 13 9 13 11 11 9 9 9 15 16 11 11 9 7 9 15 16 11 11 9 2 7 15 9 13 9 13 9 2 9 7 9 13 9 7 9 13 0 9 9 0 2
5 4 13 15 9 2
2 12 9
5 13 9 12 3 2
133 0 13 9 0 13 0 9 12 9 9 9 9 12 9 3 0 13 9 9 13 9 3 0 13 9 2 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 11 11 12 11 11 11 11 11 11 11 11 11 12 11 11 11 11 12 2
136 0 13 9 0 13 0 9 12 9 9 9 9 12 9 3 0 13 9 9 13 9 3 0 13 9 2 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 12 11 11 11 11 12 11 11 11 11 11 11 11 11 11 12 11 11 11 11 12 2
2 12 9
5 13 9 12 3 2
42 13 9 0 13 0 9 12 9 9 9 9 12 9 3 0 13 9 9 13 9 3 0 13 9 2 11 11 11 11 12 11 11 12 11 11 11 11 12 11 11 12 2
2 12 9
14 9 4 13 15 9 9 13 9 3 12 9 9 12 2
7 15 4 13 15 9 3 2
2 12 9
7 15 9 4 13 15 9 2
7 13 11 12 9 9 12 2
5 9 1 11 11 9
27 9 9 2 13 12 9 9 12 2 9 12 9 15 11 9 9 9 2 15 0 9 9 9 13 2 12 2
238 11 9 9 2 15 13 9 11 9 9 2 13 9 9 7 9 9 13 9 9 7 9 7 0 9 9 0 9 12 9 9 12 13 9 9 12 2 2 2 0 16 15 13 3 13 9 2 9 2 9 12 2 2 2 7 3 15 12 9 12 9 7 12 9 12 9 2 13 9 0 9 13 2 0 9 3 13 0 9 9 12 9 9 12 13 9 9 12 2 2 2 0 16 15 13 3 13 9 2 9 2 9 12 2 7 3 15 12 9 2 7 13 2 16 9 11 9 2 15 0 9 9 9 13 2 13 3 9 9 12 2 2 2 0 16 15 13 3 13 9 12 2 2 2 9 12 12 9 7 9 13 9 9 2 9 7 0 9 9 0 9 13 9 12 9 9 12 13 9 9 12 2 2 12 9 12 9 3 13 0 9 4 13 2 16 15 9 9 9 4 13 0 9 2 15 9 4 13 2 16 12 0 9 13 9 12 12 9 9 2 15 1 15 4 13 13 0 9 9 2 9 13 15 1 3 13 2 7 15 9 13 9 13 0 9 9 0 2
5 4 13 15 9 2
2 12 9
8 13 9 12 9 15 9 9 2
2 12 9
7 15 9 4 13 15 9 2
7 13 11 12 9 9 12 2
5 9 1 11 11 9
33 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 12 9 12 9 9 9 7 13 9 9 13 9 9 12 9 2 12 2
46 11 9 9 2 15 13 9 11 9 9 7 3 15 12 9 2 13 9 9 9 2 12 2 2 13 9 11 9 9 2 12 2 2 13 9 9 7 9 9 2 12 2 2 7 13 2
122 16 2 12 2 9 9 12 9 13 9 13 9 12 9 12 9 3 9 2 15 3 13 9 9 9 12 7 9 12 7 12 9 0 9 2 12 2 9 2 16 9 12 9 12 9 13 13 0 9 9 13 3 0 9 9 2 15 9 13 3 12 9 7 15 15 9 13 15 9 9 15 2 16 15 13 0 9 3 15 9 13 3 13 9 9 2 7 15 9 13 15 9 9 15 2 13 15 13 0 9 13 3 15 16 15 9 2 7 15 15 12 9 4 13 15 9 9 7 9 9 1 2
78 2 12 2 9 4 9 9 12 1 3 13 12 9 9 12 9 2 9 2 9 12 9 12 9 12 9 9 9 9 2 12 2 7 9 2 9 2 9 12 9 12 9 12 9 9 9 9 2 12 2 7 12 9 9 12 9 2 9 2 9 12 9 12 9 12 9 9 9 9 2 12 2 2 3 2 9 2 2
38 2 12 2 9 13 12 9 9 12 0 9 2 9 9 7 0 9 2 2 15 13 0 0 9 9 12 9 12 7 12 9 9 0 9 7 13 9 2
42 2 12 2 9 2 11 9 2 9 7 9 2 9 9 7 0 9 0 9 1 13 9 13 2 16 9 9 9 0 9 9 13 3 3 2 15 13 3 13 9 9 2
48 2 12 2 0 9 4 13 0 9 9 7 0 9 9 2 13 15 9 4 13 9 3 9 13 3 3 0 9 7 9 13 9 2 9 15 9 0 9 13 3 9 9 3 0 16 0 9 2
57 2 12 2 15 1 2 16 3 13 9 13 9 9 13 9 9 7 13 9 7 9 2 15 9 13 13 13 2 9 13 3 15 9 2 15 13 9 2 0 9 13 9 13 3 3 0 0 0 9 2 15 9 7 9 13 3 2
105 2 12 2 13 9 13 3 0 9 13 0 9 9 2 15 9 13 7 9 9 7 9 7 15 13 0 7 9 9 7 9 2 15 9 1 13 3 3 0 9 2 15 4 13 0 16 12 9 1 2 0 9 7 9 13 9 7 9 7 13 13 9 7 9 9 7 9 13 9 2 0 9 0 9 4 3 3 13 9 12 9 12 9 9 3 9 0 9 9 2 15 4 13 9 9 13 9 9 7 13 0 9 3 0 2
62 2 12 2 0 9 9 13 9 13 3 3 2 16 13 9 2 15 12 9 12 7 12 9 13 2 13 9 13 3 9 0 9 0 9 2 13 9 0 9 2 15 13 9 9 0 9 3 13 9 0 9 9 2 4 13 9 0 9 9 0 9 2
101 2 12 2 9 4 3 3 13 9 13 9 13 3 13 9 13 2 0 7 3 13 9 2 15 4 13 0 0 9 2 0 9 13 9 9 0 9 4 13 9 2 3 9 2 15 13 15 9 2 15 0 9 13 9 13 9 0 0 9 1 13 2 9 9 4 13 9 0 9 9 2 0 0 9 0 0 9 2 3 9 7 0 9 7 0 0 0 0 9 9 2 4 13 9 9 1 0 9 9 1 2
138 2 12 2 9 13 4 15 9 9 12 13 9 9 13 3 13 9 2 15 13 0 0 9 2 13 9 12 9 12 9 9 9 7 12 9 9 9 9 4 3 3 13 3 2 16 15 13 15 12 9 12 9 9 13 9 2 15 9 13 3 12 9 0 9 1 9 7 9 0 9 13 9 7 15 13 9 2 15 1 9 4 13 2 13 7 13 0 9 7 9 2 2 0 9 2 2 3 13 9 2 9 7 9 7 0 9 13 9 7 15 9 2 0 13 9 0 0 0 9 7 0 7 0 9 9 7 15 9 7 0 9 7 15 9 0 0 9 2
123 2 12 2 13 9 13 9 9 9 12 12 9 3 9 13 0 9 9 13 9 2 16 15 9 7 0 9 9 13 15 0 9 12 9 12 9 13 9 1 0 9 2 9 0 9 7 9 9 0 9 9 13 0 13 2 16 16 0 9 13 9 3 12 9 9 7 15 9 2 15 13 15 0 9 9 2 0 9 0 9 4 13 9 9 9 13 9 2 15 9 13 0 9 9 2 3 3 13 3 13 9 9 12 12 9 2 16 4 13 9 2 15 9 0 9 4 13 9 9 13 9 2 7
116 2 12 2 0 9 13 9 9 13 9 0 9 9 0 9 2 9 4 13 9 2 15 13 0 9 4 13 15 9 0 9 1 2 9 4 13 3 0 9 9 9 2 9 13 13 9 2 16 0 9 0 9 13 3 13 9 2 3 9 4 13 3 12 9 0 9 2 15 13 9 9 0 9 15 9 13 2 15 9 2 15 13 9 13 9 0 9 13 9 9 2 13 9 9 12 9 9 3 2 9 13 0 9 1 1 0 9 9 7 9 9 3 1 9 9 2
5 4 13 15 9 2
2 12 9
6 13 9 9 12 3 2
7 12 2 13 12 9 3 2
7 9 2 13 12 9 3 2
30 2 0 9 4 2 15 3 13 9 9 12 9 2 9 12 9 12 9 3 9 13 2 16 12 9 12 9 13 13 2
39 9 2 0 9 0 9 1 9 7 9 0 9 13 12 7 0 9 0 9 9 2 15 13 9 2 15 3 9 4 13 2 13 7 13 0 9 7 9 2
53 9 2 0 9 9 2 15 9 13 3 12 9 7 15 13 9 9 2 3 9 2 9 2 9 7 9 2 9 7 9 7 0 9 2 15 9 7 9 1 4 13 9 7 0 9 9 7 9 13 9 2 2 2
20 9 2 13 12 9 9 9 9 2 15 9 2 15 9 4 13 2 7 2 2
7 9 2 13 12 9 3 2
14 2 0 15 12 7 12 9 13 13 3 13 9 2 2
5 12 2 13 9 3
4 2 12 9 9
67 3 12 9 13 9 4 13 15 9 2 15 9 15 9 1 4 13 0 0 9 7 13 9 9 0 9 2 9 4 13 9 2 16 15 9 13 2 7 13 9 2 15 13 12 9 0 9 13 3 13 0 9 7 13 9 15 9 2 9 4 13 3 12 9 2 2 2
9 12 2 13 12 9 12 9 3 2
13 2 0 9 13 9 9 7 0 9 13 0 9 2
18 9 2 12 9 13 9 9 1 9 9 9 0 9 7 1 9 9 2
20 9 2 12 9 9 13 9 9 1 9 9 9 0 9 7 1 9 9 2 2
16 12 2 13 12 9 9 3 2 3 0 15 9 13 12 9 2
78 2 0 16 9 7 13 9 2 15 4 13 12 9 13 9 13 0 9 9 12 9 12 9 13 9 1 0 9 2 15 13 15 9 9 7 15 9 2 15 13 15 0 9 9 2 15 9 0 9 4 0 9 7 9 7 0 0 9 7 9 9 2 15 13 9 13 15 0 9 2 13 0 9 9 13 9 2 2
2 12 9
18 15 9 13 3 0 9 15 1 2 16 15 4 13 11 9 0 9 2
14 15 9 13 15 9 13 2 7 15 13 0 15 9 2
7 13 11 12 9 9 12 2
8 9 1 11 11 9 2 12 2
3 9 9 2
34 9 9 12 9 4 13 3 2 16 15 13 9 11 9 12 9 0 11 9 9 9 9 2 3 3 9 13 9 9 12 9 12 9 2
24 9 9 2 13 12 9 9 12 2 11 9 13 9 9 2 0 9 2 9 7 9 2 12 2
58 11 9 9 2 15 13 9 11 9 9 2 13 9 11 9 9 13 9 9 9 13 9 13 9 7 3 9 9 12 9 9 12 13 9 9 2 9 2 9 12 2 12 2 7 3 15 12 9 2 13 9 9 9 2 7 13 0 2
23 2 12 2 11 13 9 13 2 16 9 13 9 13 0 9 7 13 9 13 9 0 9 2
43 2 12 2 9 2 9 2 9 12 13 2 16 9 13 9 9 9 15 9 13 9 13 9 2 0 9 2 9 7 9 0 16 15 13 15 9 7 15 13 0 0 9 2
24 2 12 2 9 9 9 9 13 0 9 9 7 3 9 13 9 9 7 9 11 13 9 9 2
21 16 0 9 13 13 2 9 4 9 9 9 13 0 9 15 3 9 13 9 9 2
23 2 12 2 11 13 9 13 2 16 9 13 9 9 7 9 9 9 9 13 9 13 9 2
20 2 12 2 9 9 12 9 13 0 9 11 9 7 13 9 9 1 0 9 2
16 2 12 2 9 9 11 4 13 9 9 9 13 0 9 9 2
15 15 9 4 13 9 9 13 9 13 0 9 7 9 9 2
30 2 12 2 11 13 3 13 2 16 15 13 9 13 9 9 9 2 9 2 9 2 9 7 9 13 0 7 0 9 2
4 4 13 0 2
2 12 9
33 9 2 9 2 9 12 12 9 3 11 9 13 9 13 9 2 0 9 2 9 7 9 13 15 9 9 2 15 13 0 9 9 2
2 12 9
18 9 13 9 9 13 9 13 9 7 0 9 9 2 15 9 13 3 2
2 12 9
18 15 9 13 3 0 9 15 1 2 16 15 4 13 11 9 0 9 2
7 13 11 12 9 9 12 2
7 9 1 11 11 11 11 9
22 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 9 9 0 9 0 9 9
46 11 9 9 2 15 13 9 11 9 9 7 3 15 12 9 2 13 9 9 9 2 12 2 2 13 9 11 9 9 2 12 2 2 13 9 9 7 9 9 2 12 2 2 7 13 2
29 16 12 2 9 12 9 9 3 9 13 9 2 15 13 13 0 9 7 15 3 9 0 9 13 9 12 9 3 2
33 12 2 0 9 9 3 3 2 16 9 0 9 15 9 0 9 9 9 13 2 4 13 0 9 9 0 9 7 0 9 0 9 2
45 12 2 13 9 13 9 9 7 3 9 0 9 9 13 13 13 0 9 7 13 0 9 2 15 4 13 9 9 2 3 7 15 4 13 15 0 7 0 9 9 0 9 9 9 2
13 12 2 0 9 13 13 13 9 2 3 13 9 2
28 12 2 15 9 13 13 9 9 2 15 4 15 9 13 3 9 9 13 9 9 2 13 13 9 15 9 9 2
33 12 2 9 13 0 9 0 9 9 7 0 9 9 7 15 9 2 15 9 15 9 7 9 13 0 7 0 9 0 9 9 9 2
16 12 2 9 7 9 4 13 3 7 3 9 9 0 9 9 2
74 12 2 9 2 15 9 9 0 9 13 9 2 4 13 15 0 7 0 9 9 0 9 9 3 3 9 2 16 13 9 2 16 9 13 9 7 9 13 2 13 7 13 7 16 9 7 15 9 13 9 13 13 2 15 4 13 9 7 13 15 9 9 2 15 15 4 13 7 4 13 15 9 9 2
26 12 2 13 9 0 9 9 4 13 0 9 9 2 15 1 9 4 13 7 9 4 13 15 9 2 3
19 12 2 9 13 13 15 12 9 13 9 1 15 9 15 9 9 13 9 2
5 4 13 15 9 2
2 12 9
4 15 9 13 2
34 0 2 9 2 0 9 0 9 0 9 9 2 15 13 9 7 15 9 7 13 9 1 2 7 15 4 13 9 12 9 9 3 15 2
30 9 2 13 3 7 15 9 0 9 9 0 9 13 2 13 7 13 15 9 9 2 15 9 9 7 15 9 9 1 2
12 9 2 13 0 9 9 2 15 9 13 2 3
17 9 2 13 0 9 9 13 9 7 9 9 2 9 7 9 9 2
37 0 2 13 9 2 9 2 15 9 0 9 13 0 9 9 13 9 13 13 15 0 7 0 2 15 9 13 9 9 9 7 9 0 9 9 9 2
2 12 9
24 15 9 13 13 13 3 2 16 15 13 9 9 2 3 3 9 2 9 0 16 15 9 13 2
19 15 9 4 3 13 9 7 9 13 9 9 13 9 0 9 13 15 9 2
2 12 9
11 0 16 9 13 7 13 13 9 15 9 2
27 9 2 15 3 9 2 13 15 0 9 7 13 2 2 15 13 9 13 9 2 4 13 9 3 9 2 3
22 9 2 9 13 3 9 0 9 7 15 15 0 9 13 9 2 15 15 13 9 13 2
30 0 0 9 4 13 3 3 9 7 15 9 13 9 13 9 9 7 9 9 7 9 2 15 9 4 13 7 4 13 2
9 9 3 13 9 4 13 3 9 2
2 12 9
52 0 16 9 13 2 7 16 12 9 15 13 2 0 9 4 9 2 13 15 0 7 0 9 3 2 16 9 0 9 9 9 13 9 3 2 7 9 2 13 3 9 9 2 15 15 9 4 13 7 4 13 2
14 0 9 13 12 9 9 9 1 13 9 3 15 9 2
2 12 9
48 0 16 9 13 2 16 9 4 13 9 2 15 13 0 9 9 2 15 9 9 4 13 0 9 2 7 13 9 13 15 0 7 0 9 0 9 9 0 9 13 2 15 15 13 9 9 1 2
10 0 9 13 9 13 9 12 9 9 2
26 0 9 4 13 0 9 13 9 9 11 9 0 9 2 7 15 13 15 3 15 9 2 15 15 13 2
45 0 9 4 12 9 13 9 9 7 2 13 9 9 2 15 15 4 13 7 4 13 12 9 3 9 2 7 2 13 13 9 15 2 13 4 13 9 2 15 13 9 12 9 9 2
27 0 9 4 9 13 9 0 9 13 9 2 16 9 13 9 13 2 3 13 9 7 13 9 4 13 0 2
14 15 9 13 15 9 13 2 7 15 13 0 15 9 2
7 13 11 12 9 9 12 2
5 9 1 11 11 9
28 9 9 12 2 13 12 9 9 12 2 9 9 12 2 12 7 12 9 11 9 9 9 2 11 9 0 9 2
143 11 9 9 2 15 13 9 11 9 9 2 13 9 9 9 9 12 9 9 12 13 9 9 12 2 12 2 2 0 16 15 13 3 13 9 9 12 2 12 2 2 7 3 15 12 9 2 13 9 9 3 13 9 7 15 9 13 9 9 9 12 9 9 12 13 9 9 12 2 12 2 2 0 16 15 13 3 13 9 9 12 2 12 2 2 7 3 15 12 9 2 13 9 9 9 9 0 9 3 13 9 2 3 13 9 7 9 2 12 9 9 12 13 9 9 12 2 12 2 2 0 16 15 13 3 13 9 9 12 2 12 2 2 7 3 15 12 9 2 7 13 0 2
55 2 12 2 9 7 0 9 9 2 9 7 9 3 13 2 9 9 13 0 9 2 15 13 9 0 9 13 0 0 0 9 9 13 15 3 2 16 9 13 3 0 7 3 0 3 9 7 9 9 9 13 13 9 9 2
26 0 9 9 9 9 13 15 2 3 3 9 13 9 13 9 7 0 9 2 13 13 9 9 0 9 2
20 9 13 9 9 13 0 9 9 2 15 9 4 13 3 16 0 9 4 13 2
20 2 12 2 9 9 9 13 3 3 2 7 15 13 0 9 7 9 9 9 2
63 9 9 13 9 9 2 16 9 0 9 13 13 9 7 15 9 13 13 9 9 7 16 0 9 13 13 7 16 9 13 9 9 13 4 13 0 9 7 16 0 9 9 9 13 4 13 0 9 7 9 4 13 9 9 9 9 3 13 9 7 15 9 2
27 2 12 2 11 9 15 9 13 9 13 13 0 9 9 9 12 12 9 3 2 16 9 9 9 13 9 2
8 9 13 9 9 9 9 9 2
34 2 12 2 9 0 7 0 9 15 9 9 13 11 9 9 4 13 9 13 9 7 9 1 13 3 9 9 9 13 9 2 12 2 2
14 4 13 2 13 15 9 13 9 9 13 9 0 9 2
35 2 12 2 9 0 9 15 9 15 0 9 9 2 15 4 13 9 2 4 13 13 9 13 9 7 9 1 13 3 9 9 9 13 9 2
19 9 13 2 16 15 9 13 9 9 13 7 15 0 9 13 13 0 9 2
25 2 12 2 9 9 4 13 15 9 13 9 9 9 9 9 7 15 15 9 13 9 4 13 9 2
11 2 12 2 9 13 9 9 4 13 9 2
18 3 4 13 9 9 7 9 2 15 13 13 9 9 13 9 9 9 2
16 2 12 2 9 12 2 12 7 12 9 4 15 1 13 3 2
18 2 12 2 15 9 13 9 13 9 7 9 9 13 0 9 9 0 2
5 4 13 15 9 2
2 12 9
17 13 9 12 9 0 13 9 9 0 9 2 2 5 9 9 5 2
2 12 9
17 13 9 12 9 0 13 9 9 0 9 2 2 5 9 9 5 2
2 12 9
7 13 9 12 9 0 3 2
15 2 13 9 12 9 0 15 9 9 13 11 9 9 2 2
2 12 9
16 9 4 13 7 13 15 9 9 13 9 3 12 9 9 12 2
7 15 4 13 15 13 9 2
10 15 4 13 15 9 12 9 9 12 2
20 15 9 13 9 4 13 15 9 7 15 4 13 0 9 2 16 15 3 13 2
9 9 4 13 15 2 3 9 13 2
2 12 9
18 15 9 13 3 0 9 15 1 2 16 15 4 13 11 9 0 9 2
2 12 9
7 15 9 4 13 15 9 2
7 13 11 12 9 9 12 2
6 9 1 11 11 9 9
31 9 9 12 2 13 12 9 9 12 2 11 9 9 9 7 0 9 13 9 7 9 9 11 13 9 12 9 9 7 15 9
48 11 9 9 2 15 13 9 12 9 9 12 13 9 0 9 12 11 9 9 9 7 0 9 13 9 7 9 9 7 3 15 12 9 3 11 9 13 9 12 9 12 9 1 2 7 13 0 2
26 2 12 2 9 13 12 9 9 12 11 9 9 9 7 0 9 13 9 7 9 9 11 13 9 12 2
14 2 12 2 9 12 9 13 7 9 13 3 9 12 2
34 2 12 2 15 0 9 13 4 13 13 12 9 9 12 1 2 3 9 12 9 13 9 13 2 7 15 9 4 13 3 13 9 1 2
5 0 9 13 0 2
15 2 12 2 9 12 9 4 3 3 13 7 9 4 13 2
4 4 13 0 2
2 12 9
5 13 9 12 3 2
20 9 2 13 12 9 12 9 13 9 9 2 12 9 2 9 2 12 9 2 2
22 9 2 13 12 9 0 9 9 2 12 9 9 12 2 9 2 12 9 9 12 2 2
6 9 2 13 12 9 2
10 9 2 13 9 15 9 9 13 9 2
2 12 9
9 15 9 13 3 12 9 9 12 2
2 12 9
7 9 13 11 9 0 9 2
7 13 11 12 9 9 12 2
5 9 1 9 11 11
23 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 15 16 11 9 9 13 9 9
89 11 9 9 2 15 13 9 11 9 9 7 3 15 12 9 2 13 9 9 0 9 9 13 9 7 9 12 9 1 13 9 2 15 13 9 9 13 9 2 7 3 15 9 9 2 15 13 9 13 15 0 9 2 16 0 9 7 15 9 13 9 4 13 3 15 9 13 9 2 13 9 9 9 2 12 2 2 13 9 11 9 9 2 12 2 2 7 13 2
33 16 2 12 2 9 2 9 2 9 12 2 12 2 9 13 9 0 9 2 15 13 9 7 9 15 16 11 9 9 13 9 9 2
65 2 12 2 15 0 9 13 9 13 13 0 9 3 7 3 0 9 3 2 15 13 9 7 9 13 9 2 3 2 9 2 2 0 9 2 9 0 9 9 13 9 2 9 12 9 2 7 9 0 2 0 7 0 9 9 7 9 13 9 2 9 7 9 2 2
62 2 12 2 9 12 0 9 4 13 0 2 9 0 9 9 13 9 2 7 15 1 9 9 4 13 15 0 9 9 2 13 9 9 7 9 13 0 9 0 9 13 0 13 0 9 9 15 9 2 15 1 9 9 7 9 13 0 9 13 0 9 2
30 2 12 2 9 13 9 7 9 9 9 15 9 13 13 3 0 2 16 9 13 9 15 2 3 15 0 9 13 15 2
94 2 12 2 0 9 9 7 9 9 7 9 13 9 12 0 9 9 2 3 2 9 12 9 2 2 13 0 7 0 9 2 15 13 3 9 9 2 9 9 7 15 0 9 13 9 2 3 13 9 9 7 9 2 0 9 9 9 2 9 9 7 9 2 9 9 7 9 7 9 13 9 9 2 9 9 1 7 0 9 0 7 0 9 9 9 9 4 3 3 13 0 9 0 2
108 2 12 2 13 0 13 0 7 0 9 9 9 2 3 0 9 4 15 9 13 0 9 2 15 4 13 9 0 9 9 2 13 0 13 9 2 15 13 0 9 4 13 0 7 15 4 13 9 7 4 13 3 13 9 7 0 9 7 9 0 9 2 3 13 0 13 9 0 9 3 9 2 4 3 13 9 9 7 9 9 7 9 2 0 9 9 13 3 3 13 9 2 15 13 9 2 0 9 7 15 9 7 15 9 13 9 9 2
48 2 12 2 9 9 15 16 9 13 0 13 9 2 15 1 9 13 0 9 2 15 13 9 2 13 2 7 13 0 0 9 4 13 2 4 13 15 2 16 9 4 13 15 3 15 0 9 2
34 2 12 2 4 13 9 7 13 15 0 9 2 15 4 13 15 9 2 15 13 2 16 0 9 13 9 13 13 9 0 9 0 9 2
67 2 12 2 9 7 9 0 0 9 9 4 13 9 7 15 9 3 13 9 7 13 0 9 9 9 7 9 13 9 2 16 9 9 4 13 2 3 13 0 2 16 9 4 13 13 0 9 2 16 0 9 4 13 0 9 2 16 9 13 0 9 2 9 7 9 1 2
60 2 12 2 13 0 2 16 13 0 7 0 9 9 2 15 4 13 2 4 9 13 9 13 7 13 15 13 0 9 2 16 13 13 2 16 9 9 13 9 13 9 13 9 9 7 9 2 13 9 13 9 15 9 9 7 3 0 9 9 2
56 2 12 2 4 13 9 2 9 9 2 7 13 15 2 16 9 9 13 9 4 13 15 9 1 2 7 4 13 9 2 9 2 2 3 13 3 13 15 2 16 9 4 13 9 0 9 9 1 2 7 13 0 9 9 9 2
51 2 12 2 13 3 13 2 15 4 13 9 13 9 2 7 15 9 9 2 15 9 9 13 9 9 2 7 13 3 0 9 13 9 2 9 7 9 13 9 2 4 3 13 9 9 7 9 9 13 9 2
97 2 12 2 13 3 13 2 15 9 9 4 13 9 13 9 2 7 4 13 15 0 9 13 15 0 9 7 13 9 2 3 13 0 13 3 9 13 13 9 7 9 7 3 9 15 2 3 9 4 13 2 13 9 7 13 9 0 9 2 16 15 4 13 9 2 4 3 13 9 2 15 3 9 4 13 15 9 13 9 9 7 13 9 15 2 9 9 9 4 3 13 9 9 7 9 1 2
69 2 12 2 4 13 9 2 15 3 0 9 4 13 9 2 7 4 3 13 15 2 16 15 13 4 13 9 2 16 9 9 4 13 3 16 12 9 7 3 16 12 9 2 0 9 13 3 3 13 2 16 9 4 15 9 13 0 9 9 3 12 9 7 3 12 7 12 9 2
68 2 12 2 13 3 13 9 7 9 13 9 9 15 1 2 16 13 9 0 7 0 9 2 4 3 13 9 9 7 9 9 7 13 15 2 16 0 9 4 13 9 13 9 1 7 16 9 13 3 9 9 2 9 13 4 13 2 16 13 9 7 15 9 13 13 0 9 2
93 2 12 2 13 3 13 15 16 2 13 0 9 7 13 2 9 4 3 13 12 9 7 3 12 9 13 15 9 2 9 7 9 4 13 2 16 9 13 9 7 9 0 2 7 15 9 4 13 2 16 9 4 13 9 2 13 3 13 9 9 7 15 2 16 9 9 4 13 9 0 2 16 0 0 9 13 0 13 9 2 7 13 3 13 9 9 9 2 16 9 13 9 2
53 2 12 2 13 3 13 0 9 0 9 2 16 15 13 0 2 7 13 9 2 15 9 4 13 3 2 16 13 15 2 16 13 0 9 13 9 2 3 13 3 13 9 0 9 2 16 9 13 7 16 15 13 2
89 2 12 2 13 3 13 15 2 16 9 9 13 12 9 13 2 3 16 9 13 2 16 15 4 13 2 16 9 4 13 13 9 0 9 2 13 3 3 13 0 9 9 7 9 15 9 2 13 13 9 9 0 2 3 4 13 15 2 16 16 9 9 13 9 9 2 9 13 13 13 9 7 9 0 9 2 16 15 9 13 15 9 9 2 15 9 9 13 2
39 2 12 2 13 3 13 3 15 2 16 9 7 9 4 13 3 2 16 9 13 9 0 9 9 13 7 16 9 13 13 15 9 9 2 15 9 9 13 2
66 2 12 2 9 12 9 13 13 9 9 9 2 16 0 11 9 13 9 9 7 4 13 11 9 13 2 16 0 9 4 15 1 13 7 11 9 9 9 13 13 3 13 0 9 9 0 9 2 3 9 7 0 9 13 0 9 9 9 2 15 0 9 13 9 9 2
19 2 12 2 4 13 9 13 9 2 16 9 0 9 13 15 9 3 0 2
27 2 12 2 13 3 13 15 2 16 9 9 13 9 4 13 9 3 2 16 15 9 1 4 3 13 9 2
33 2 12 2 9 0 9 9 13 3 2 16 9 13 9 7 13 9 9 9 7 9 9 13 9 9 7 15 9 3 13 9 9 2
31 2 12 2 13 3 13 15 2 16 9 0 7 13 9 4 13 0 9 2 9 13 9 9 2 7 15 9 13 9 9 2
23 2 12 2 13 3 13 9 9 7 9 13 13 9 9 9 13 3 0 9 13 9 9 2
21 2 12 2 9 9 13 9 13 0 0 13 9 2 16 9 7 9 9 13 0 2
42 2 12 2 13 3 13 15 2 16 16 9 13 13 9 0 9 2 4 9 13 15 9 7 16 15 9 4 13 0 9 3 0 16 15 13 2 16 9 4 13 9 2
13 2 12 2 0 9 9 4 13 9 9 9 9 2
37 2 12 2 13 0 2 16 9 13 9 13 3 0 9 7 9 7 16 9 13 2 9 9 9 13 2 0 9 13 2 16 9 13 9 13 9 2
40 2 12 2 13 0 13 9 2 15 4 13 9 9 9 9 9 2 3 13 9 9 9 2 7 13 9 2 15 13 9 13 9 4 13 2 7 13 9 9 2
50 2 12 2 9 15 16 11 9 9 13 9 9 12 9 9 12 13 9 2 9 2 9 12 2 12 2 9 13 9 2 9 2 9 12 7 13 9 0 0 9 9 15 16 11 9 9 13 9 9 2
20 2 12 2 9 2 9 2 9 12 9 13 0 9 13 3 2 16 15 13 2
12 2 12 2 15 1 0 9 4 13 12 9 2
36 2 12 2 9 2 9 7 9 1 0 9 4 15 1 13 7 13 2 13 3 13 0 9 7 9 2 9 2 9 12 1 3 13 9 9 2
5 4 13 15 9 2
2 12 9
1 9
17 0 9 4 13 9 13 9 2 16 9 9 0 9 9 13 9 2
22 0 9 13 9 13 2 16 15 9 9 13 0 16 0 9 13 0 9 0 9 9 2
6 0 9 13 3 9 2
31 15 4 3 13 9 13 9 2 3 16 9 3 3 13 15 1 2 0 9 13 13 9 7 9 13 13 0 9 15 9 2
50 0 15 9 9 2 0 9 2 4 13 13 9 2 15 13 0 2 3 3 15 9 0 16 9 13 9 2 7 0 9 13 2 15 9 2 15 2 16 15 13 13 15 9 0 2 13 9 0 9 2
2 12 9
2 9 9
2 9 9
15 0 9 13 3 9 0 9 0 9 13 7 13 13 9 2
19 16 9 13 13 7 13 0 9 9 2 9 13 15 9 7 9 9 9 2
37 0 9 2 15 1 13 13 9 7 9 2 0 9 13 4 13 0 9 13 7 15 4 13 9 9 3 2 16 13 2 16 0 9 13 13 9 2
27 0 9 9 13 3 9 9 13 0 9 9 2 16 9 9 13 3 12 9 9 9 13 9 9 9 9 2
17 0 9 9 4 3 13 3 3 2 16 13 9 13 0 9 13 2
60 0 16 0 9 13 13 0 9 7 9 13 0 7 0 9 13 0 9 9 13 4 13 0 9 2 0 9 9 13 9 9 9 13 0 9 9 2 9 7 15 9 7 9 2 7 0 9 13 0 9 13 9 9 13 2 16 9 13 0 2
72 0 16 0 9 13 9 9 7 0 9 9 2 15 13 0 16 9 2 0 7 0 2 9 13 9 2 9 7 15 9 2 9 4 9 1 13 13 0 9 13 7 15 4 13 9 13 9 13 3 2 16 13 9 13 13 9 13 0 9 7 9 2 15 13 4 13 15 9 0 9 13 2
24 16 9 2 15 13 9 9 0 2 13 9 9 13 9 2 4 15 13 13 9 0 9 13 2
52 13 9 13 3 9 7 3 12 9 2 7 9 0 9 13 9 13 9 0 15 9 13 2 16 13 2 16 9 13 9 13 13 0 9 0 7 16 9 0 9 13 9 9 13 3 12 9 9 9 13 9 2
38 0 9 13 3 9 9 13 9 9 9 15 9 2 16 15 9 4 13 0 9 3 13 9 3 7 15 13 0 0 9 0 9 9 7 9 13 9 2
18 9 0 9 13 9 13 9 2 16 13 2 16 0 9 4 3 13 2
12 16 0 9 13 13 2 13 3 9 13 9 2
28 9 13 3 15 0 9 1 2 15 13 0 7 0 9 2 13 0 9 3 4 13 9 15 9 13 9 9 2
58 16 9 15 9 13 0 9 9 13 0 2 0 9 13 9 9 7 9 0 9 0 9 7 15 9 13 13 9 1 2 9 0 9 13 3 13 9 3 13 9 9 9 2 7 0 9 9 15 13 12 9 0 9 13 13 0 9 2
23 9 9 13 9 13 9 7 9 0 9 3 2 7 15 13 13 0 9 9 13 0 9 2
29 0 9 13 9 9 9 9 13 2 9 0 13 9 13 9 3 2 16 15 13 1 9 7 12 9 13 9 9 2
32 0 9 2 9 7 15 9 7 9 1 13 9 4 13 0 9 2 15 13 13 13 9 7 9 0 9 9 7 9 0 9 2
94 16 0 9 13 3 4 13 2 15 4 13 13 0 9 2 9 2 15 9 9 13 9 7 9 9 13 0 9 13 9 0 9 9 7 9 9 9 9 2 0 9 7 9 13 7 13 0 9 15 0 9 9 9 7 9 0 9 9 9 9 2 15 3 15 0 9 15 9 2 16 3 13 9 9 13 13 9 2 15 15 9 7 9 3 13 15 0 9 13 9 9 9 9 2
87 0 15 16 9 3 13 9 7 3 0 9 2 15 13 9 9 2 9 2 9 12 2 12 2 2 3 13 9 9 13 0 9 2 15 13 9 2 13 9 7 0 9 9 7 0 0 9 15 9 2 3 9 2 13 9 9 7 2 16 15 13 13 0 2 15 3 0 9 2 3 13 0 9 3 9 13 7 13 9 2 15 4 13 13 0 9 2
20 0 0 9 2 15 13 9 2 13 0 9 13 9 15 9 13 13 0 9 2
18 3 9 13 9 7 13 13 15 9 9 13 0 9 2 15 13 9 2
24 9 9 13 13 9 9 1 13 0 9 2 15 13 9 2 7 15 13 12 9 9 13 9 2
2 9 9
17 0 9 13 3 13 7 13 9 9 2 15 4 13 9 9 9 2
70 0 16 9 13 13 7 16 13 15 2 16 9 13 13 0 2 16 9 7 9 7 0 9 1 13 9 7 9 2 9 4 13 15 9 9 2 15 13 9 13 0 3 0 9 2 7 16 9 13 13 0 9 7 15 13 13 0 9 2 15 15 13 13 2 15 3 15 0 9 2
26 0 9 13 9 9 7 9 0 0 9 2 3 9 7 9 2 7 9 9 9 0 9 9 9 9 2
27 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 9 9 9 9 2 9 2 9 12 13 9 9
40 11 9 9 2 15 13 9 11 9 9 2 13 9 9 0 9 12 9 9 12 13 9 9 2 9 2 9 12 7 3 15 12 9 12 9 2 7 13 0 2
24 2 12 2 9 9 2 9 2 9 12 4 13 9 2 15 13 9 0 9 13 9 9 11 2
31 2 12 2 9 9 2 9 2 9 12 12 9 3 9 4 9 2 9 2 9 12 12 9 13 9 13 13 9 9 9 2
19 15 9 4 13 9 3 9 2 9 2 9 12 12 7 12 9 13 9 2
16 9 13 15 9 9 2 15 9 13 9 9 0 7 15 0 2
23 2 12 2 3 13 9 9 0 9 0 9 13 2 16 9 9 4 13 12 9 13 9 2
13 2 12 2 15 9 13 9 13 9 9 9 0 2
5 4 13 15 9 2
2 12 9
31 9 2 9 2 9 12 13 9 9 12 7 12 9 9 12 0 9 13 9 9 9 9 9 13 12 9 12 9 9 1 2
2 12 9
9 15 9 13 3 12 9 9 12 2
14 15 9 13 15 9 0 2 7 15 13 0 15 9 2
7 13 11 12 9 9 12 2
7 9 1 11 11 11 9 9
38 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 9 9 9 9 0 9 13 9 9 2 9 2 9 12 9 0 9 2 11 9 0 9 2
65 11 9 9 2 15 13 9 11 9 9 2 13 9 9 9 9 9 9 0 9 12 9 9 12 13 9 9 2 9 2 9 12 2 12 2 2 0 16 15 13 3 13 9 9 2 9 2 9 12 2 12 2 2 7 3 15 12 7 12 9 2 7 13 9 2
29 12 2 9 2 9 2 9 12 3 9 9 4 13 3 15 3 13 9 2 15 13 9 9 13 9 13 13 9 2
30 12 2 9 9 4 13 3 2 16 9 4 13 15 9 13 9 0 9 9 9 0 9 9 7 15 9 9 0 9 2
39 12 2 0 9 13 9 9 13 4 13 15 9 2 15 9 4 13 2 0 9 15 13 9 13 9 2 9 2 7 9 9 9 0 9 9 2 9 2 2
18 12 2 9 9 9 9 3 9 9 4 3 13 9 2 9 7 9 2
23 9 7 9 13 3 3 0 9 13 9 2 7 15 1 9 13 3 13 3 9 7 9 2
24 12 2 0 9 2 9 13 9 7 9 13 13 9 9 9 4 13 3 9 2 9 7 9 2
20 12 2 11 11 9 7 11 11 9 4 13 9 2 9 2 9 12 9 0 2
53 12 2 4 13 0 9 1 15 9 9 2 16 9 4 13 15 9 9 9 9 13 9 0 9 9 9 13 9 2 15 4 13 9 9 12 2 12 2 2 0 16 15 13 3 13 9 12 2 12 2 2 3 2
12 12 2 15 9 13 9 13 0 9 9 0 2
5 4 13 15 9 2
2 12 9
14 13 9 2 9 2 9 12 9 0 15 9 9 3 2
2 12 9
18 15 9 13 3 0 9 15 1 2 16 15 4 13 11 9 0 9 2
12 15 13 0 9 15 1 2 16 15 4 13 2
14 15 9 13 15 9 13 2 7 15 13 0 15 9 2
7 13 11 12 9 9 12 2
6 9 1 11 11 9 9
31 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 13 0 9 9 9 12 9 9 12 7 12 9 9 12 0 9
42 11 9 9 2 15 13 9 11 9 9 2 13 9 9 0 9 12 9 9 12 13 9 9 2 9 2 9 12 7 3 15 12 9 12 9 0 9 2 7 13 0 2
72 2 12 2 9 2 9 2 9 12 12 9 12 9 13 2 16 15 9 12 9 12 9 13 9 13 7 0 9 9 9 13 13 9 12 9 12 9 9 7 9 9 13 9 2 13 9 9 9 13 9 7 9 12 13 3 0 9 2 11 2 2 3 16 15 13 9 2 4 13 13 9 2
46 2 12 2 9 9 2 9 2 9 12 9 13 0 9 0 9 13 9 9 9 9 9 12 9 9 12 13 9 9 2 9 2 9 12 13 2 16 0 9 13 0 9 13 9 9 2
27 2 12 2 9 2 9 2 9 12 12 9 13 2 16 0 9 9 4 13 3 15 9 12 9 13 9 2
13 2 12 2 15 9 13 9 13 9 9 9 0 2
5 4 13 15 9 2
2 12 9
28 9 2 9 2 9 12 12 9 13 0 9 9 13 12 12 9 12 9 9 12 7 12 9 9 12 0 9 2
2 12 9
9 15 9 13 3 12 9 9 12 2
14 15 9 13 15 9 0 2 7 15 13 0 15 9 2
7 13 11 12 9 9 12 2
7 9 1 11 11 11 9 9
23 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 9 9 2 11 9 0 9 2
53 11 9 9 2 15 13 9 11 9 9 2 13 9 9 9 12 9 9 12 13 9 9 12 2 12 2 2 0 16 15 13 3 13 9 2 9 2 9 12 2 12 2 2 7 3 15 12 9 2 7 13 0 2
20 2 12 2 9 12 12 9 9 9 3 11 3 9 9 13 9 9 13 9 2
17 9 4 13 12 9 2 16 15 0 9 12 9 9 0 9 13 2
26 2 12 2 15 9 9 13 11 9 13 9 9 9 4 13 2 16 9 12 12 9 9 13 9 13 2
22 11 9 4 3 13 7 13 0 9 9 9 0 9 0 9 12 9 9 9 9 3 2
24 2 12 2 9 9 13 9 4 13 0 9 11 9 9 7 0 9 9 15 9 9 13 9 2
17 2 12 2 15 9 13 9 13 9 7 9 9 13 9 9 0 2
5 4 13 15 9 2
2 12 9
19 13 15 9 9 13 11 7 15 9 9 13 9 9 9 0 9 13 9 2
2 12 9
17 15 9 13 3 15 9 13 9 2 15 15 13 11 9 0 9 2
14 15 9 13 15 9 13 2 7 15 13 0 15 9 2
7 13 11 12 9 9 12 2
6 9 1 11 11 9 9
15 12 9 0 9 13 9 7 0 9 7 9 13 9 9 9
17 11 9 9 9 0 9 13 9 7 0 9 7 9 13 9 9 9
39 11 9 2 15 2 13 9 9 12 9 2 2 13 9 0 9 12 13 9 9 0 9 13 9 7 0 9 7 9 13 9 9 2 0 13 9 9 3 2
23 2 5 2 9 11 2 11 7 11 13 7 11 9 2 11 2 0 9 13 9 2 12 9
23 2 5 2 9 11 2 11 7 11 7 11 7 11 2 3 13 11 2 13 9 2 12 9
12 2 5 2 9 11 7 11 0 9 2 12 9
12 2 5 2 9 11 7 11 0 9 2 12 9
12 2 5 2 9 11 7 11 0 9 2 12 9
10 2 5 2 9 11 13 9 2 12 9
30 2 5 2 11 7 11 2 11 7 11 7 11 7 11 0 9 13 7 9 11 2 11 7 11 13 9 2 2 12 9
20 2 5 2 9 11 7 11 2 11 7 11 7 11 7 11 0 9 2 12 9
10 2 5 2 9 11 13 9 2 12 9
13 2 5 2 9 11 9 13 9 13 9 2 12 9
20 2 5 2 9 9 7 11 9 9 2 3 13 11 2 13 9 2 2 12 9
11 2 5 2 9 9 13 9 2 2 12 9
15 2 5 2 9 11 9 3 13 11 13 9 2 2 12 9
11 2 5 2 9 11 13 9 2 2 12 9
11 2 5 2 9 11 13 9 2 2 12 9
11 2 5 2 9 11 13 9 2 2 12 9
12 2 5 2 9 11 9 13 9 2 2 12 9
13 2 5 2 9 11 9 9 13 9 2 2 12 9
11 2 5 2 9 9 13 9 2 2 12 9
11 2 5 2 9 11 13 9 2 2 12 9
12 2 5 2 9 11 9 13 9 2 2 12 9
20 2 5 2 9 11 9 7 11 0 9 9 2 11 2 13 9 2 2 12 9
20 2 5 2 9 11 9 7 11 0 9 9 2 11 2 13 9 2 2 12 9
12 2 5 2 9 11 9 13 9 2 2 12 9
13 2 5 2 9 11 7 11 13 9 2 2 12 9
11 2 5 2 9 11 13 9 2 2 12 9
13 2 5 2 9 11 0 9 13 9 2 2 12 9
13 2 5 2 9 11 7 11 0 9 2 2 12 9
13 2 5 2 9 11 7 11 0 9 2 2 12 9
13 2 5 2 9 11 7 11 0 9 2 2 12 9
16 2 5 2 9 11 7 0 11 9 11 0 9 2 2 12 9
13 2 5 2 9 11 7 11 0 9 2 2 12 9
13 2 5 2 9 11 7 11 0 9 2 2 12 9
13 2 5 2 9 11 7 11 0 9 2 2 12 9
14 2 11 2 9 9 7 11 0 0 9 2 2 12 9
11 2 11 2 9 0 9 2 2 12 9 2
12 2 8 2 2 11 9 9 2 11 12 12 12
2 0 9
2 9 9
26 9 9 11 9 7 15 9 7 11 9 0 9 13 9 12 9 9 13 9 13 9 9 2 9 13 2
1 9
13 0 9 13 11 9 7 11 9 13 9 9 9 2
30 0 11 7 0 11 9 9 13 3 3 0 2 16 9 7 9 13 3 2 15 1 9 9 9 4 13 13 15 9 2
17 15 9 9 13 9 4 13 9 13 9 0 9 9 7 9 9 2
12 0 11 7 11 9 13 3 12 9 9 12 2
32 12 9 4 3 13 2 9 2 9 2 9 7 9 2 9 2 9 7 9 2 9 7 9 2 9 7 9 7 9 7 9 2
9 3 4 13 9 7 9 13 9 2
40 0 9 7 9 13 3 7 0 0 9 9 2 15 13 11 9 7 15 11 9 13 9 9 7 3 11 9 2 9 9 7 11 9 9 1 13 0 9 1 2
34 0 15 1 9 13 11 7 11 1 13 9 13 9 3 2 16 9 13 7 15 13 9 7 9 1 13 3 0 9 7 9 13 9 2
12 0 9 9 13 11 9 15 9 16 9 9 2
27 16 13 9 2 15 13 11 9 13 9 0 7 0 9 2 9 9 13 9 9 2 15 13 3 9 9 2
12 3 9 13 9 9 3 9 9 7 9 9 2
12 0 9 9 7 9 7 9 13 9 13 9 2
11 9 9 7 9 4 13 3 11 9 1 2
1 9
2 9 9
22 9 9 11 9 7 15 9 7 11 9 0 9 13 9 12 9 9 13 9 13 9 9
29 11 9 9 2 15 13 9 11 9 9 7 3 15 12 9 12 9 0 9 2 13 9 9 9 2 7 13 0 2
29 2 12 2 11 9 7 15 9 7 11 9 0 9 13 9 12 9 9 12 2 7 15 13 3 12 9 9 12 2
18 2 12 2 9 12 9 1 9 4 13 9 9 13 9 7 9 9 2
4 4 13 0 2
2 12 9
33 11 9 7 15 9 7 11 9 0 9 13 9 13 9 13 9 9 2 15 13 0 9 12 9 9 2 13 9 13 9 9 9 2
2 12 9
21 9 13 11 9 7 15 9 7 11 9 9 9 2 7 15 9 13 15 9 3 2
20 11 9 9 13 9 9 11 9 7 15 9 1 7 13 9 9 9 13 9 2
22 9 2 15 13 11 9 13 9 0 7 0 9 2 11 9 13 9 9 13 9 9 2
6 11 9 0 9 13 2
10 9 13 9 9 7 15 13 15 1 2
14 13 11 2 2 2 9 2 2 2 9 2 2 2 2
3 9 1 9
1 9
5 9 2 12 2 2
11 11 7 11 9 9 9 7 9 13 9 9
25 11 7 11 9 2 15 13 9 11 9 7 15 9 7 11 9 0 9 13 9 2 7 13 0 2
28 0 9 9 2 9 7 9 9 13 0 7 0 0 9 9 2 15 13 11 9 7 15 11 9 13 9 9 2
24 0 9 9 2 9 7 9 13 9 13 15 9 1 9 0 9 7 15 13 3 9 13 9 2
24 0 9 13 0 9 2 15 13 0 0 9 9 2 9 2 9 9 2 0 9 7 9 9 2
19 0 11 7 0 11 9 9 9 13 3 0 2 16 9 7 9 13 3 2
11 0 4 13 9 0 9 9 7 9 9 2
28 11 9 13 9 9 9 7 9 11 9 9 1 9 2 15 13 9 2 16 0 11 9 4 13 0 7 0 2
19 0 9 4 3 13 13 9 9 9 0 0 9 9 9 9 7 9 1 2
14 0 9 12 9 1 4 13 9 9 13 9 7 9 2
4 4 13 0 2
2 15 9
20 11 9 7 11 9 9 13 9 7 9 13 9 7 13 15 9 2 15 13 9
23 0 9 7 9 13 9 9 13 9 4 3 13 9 0 9 9 11 7 11 0 0 9 2
14 9 13 15 0 9 9 9 9 9 7 13 9 9 2
10 15 9 13 3 9 2 15 15 13 2
2 13 2
2 9 1
2 9 12
1 9
9 11 7 11 9 9 12 9 7 9
4 0 9 7 9
13 9 13 11 9 7 15 9 7 11 9 9 9 2
7 15 9 13 15 9 3 2
2 0 9
13 9 13 9 9 2 15 15 13 9 15 9 1 2
5 9 13 13 9 2
7 15 4 3 13 9 9 2
2 0 9
8 9 13 9 9 3 13 9 2
23 9 13 3 0 0 9 13 3 9 7 9 13 9 2 15 13 11 7 11 9 13 9 2
12 15 13 3 9 9 2 9 7 9 13 9 2
11 13 9 13 9 0 9 9 13 9 3 2
19 9 13 3 13 9 13 9 2 13 15 3 13 9 7 13 9 15 9 2
24 0 9 9 7 9 2 3 9 7 9 9 2 9 9 2 9 13 9 15 13 7 15 9 2
22 0 9 9 7 9 13 0 0 9 9 7 9 7 9 11 13 9 13 0 9 9 2
8 0 9 0 9 0 9 9 2
30 9 13 13 0 2 7 9 4 3 11 7 11 0 9 9 9 13 15 15 9 13 9 2 3 0 9 2 3 9 2
11 3 0 9 4 13 9 15 3 9 9 2
14 15 9 9 4 13 15 2 0 7 15 3 13 9 2
2 0 9
14 11 9 9 7 11 9 9 9 13 3 9 0 9 2
7 15 9 13 9 13 9 2
2 0 9
14 9 13 3 2 16 9 15 13 2 7 3 3 9 2
15 9 4 13 3 15 9 9 2 15 0 9 13 15 9 2
14 15 9 9 13 9 9 3 9 13 9 12 9 13 2
12 9 9 13 9 3 13 9 7 3 13 9 2
8 0 9 13 9 3 9 13 2
21 11 9 9 2 9 2 9 12 2 13 12 9 9 12 2 9 13 9 2 12 2
73 11 9 9 2 15 13 9 11 9 9 13 9 12 9 9 12 13 9 9 2 9 2 9 12 2 12 2 7 3 15 12 9 12 9 7 12 9 12 9 2 13 9 11 9 13 9 12 9 9 12 13 9 9 2 9 2 9 12 2 12 2 7 3 15 12 9 12 9 2 7 13 0 2
41 2 12 2 9 13 9 12 9 9 12 13 11 9 9 2 9 2 9 12 2 12 2 2 12 2 4 3 13 9 2 9 2 9 12 2 12 2 2 12 2 2
22 16 0 9 13 3 0 0 9 2 13 0 2 16 0 9 13 3 12 9 15 9 2
17 2 12 2 11 9 2 11 2 13 9 13 9 9 4 13 9 2
21 15 9 9 13 13 11 9 2 11 2 0 9 9 9 12 9 13 9 13 9 2
28 15 9 13 13 9 7 9 2 15 13 9 2 0 9 9 9 2 7 3 9 3 13 9 13 9 13 3 2
41 2 12 2 11 13 9 11 9 9 2 3 2 9 2 2 9 3 7 11 9 7 11 9 9 2 3 2 9 2 2 1 3 3 16 15 13 3 11 9 9 2
17 15 9 4 13 9 7 15 9 9 12 9 12 9 13 9 9 2
28 2 12 2 9 12 9 13 2 16 11 13 0 9 9 0 9 7 0 0 9 7 3 0 9 11 9 13 2
20 9 12 9 13 2 16 0 9 13 2 3 3 16 0 2 12 9 13 9 2
51 2 12 2 0 9 4 13 0 13 0 9 9 11 9 9 13 9 9 0 9 13 9 2 15 15 13 0 9 13 9 9 7 0 9 7 0 9 3 7 15 13 15 9 2 16 11 9 9 13 13 2
10 15 9 4 3 13 9 9 13 9 2
15 9 9 9 4 15 9 13 2 16 9 13 15 9 1 2
13 9 11 4 13 0 15 9 13 9 0 9 9 2
39 2 12 2 9 2 9 2 9 12 12 9 13 2 16 11 4 13 0 9 9 9 9 1 2 7 13 11 9 13 15 9 9 3 7 3 9 13 9 2
28 15 9 12 9 12 9 13 2 16 11 4 13 9 9 2 15 3 4 13 9 13 9 7 13 0 9 9 2
43 2 12 2 11 13 9 2 9 2 9 12 12 9 13 9 7 13 9 9 9 9 2 13 9 15 2 3 9 15 9 13 3 7 13 9 2 7 13 0 9 0 9 2
34 9 2 9 2 9 12 12 9 11 13 9 13 9 9 9 13 9 7 9 13 15 9 9 7 9 2 15 9 13 13 13 9 9 2
22 13 0 2 16 9 9 13 9 9 9 13 9 13 3 11 9 0 9 9 0 9 2
35 2 12 2 9 2 9 2 9 12 12 9 13 2 16 9 4 13 9 9 0 9 7 13 11 1 0 9 13 9 12 9 13 9 9 2
39 2 12 2 16 13 13 2 16 11 9 12 9 1 13 9 13 13 15 9 13 13 15 9 9 0 9 2 9 12 9 13 7 9 13 7 15 0 9 2
51 9 2 9 2 9 12 13 2 16 9 12 9 7 9 12 9 13 3 15 2 16 9 0 9 4 13 7 13 0 9 15 0 13 9 11 9 13 9 9 7 13 9 13 9 3 0 13 9 13 9 2
19 2 12 2 9 4 13 3 15 9 0 9 11 9 7 9 9 9 9 2
10 9 4 3 4 13 9 7 13 9 2
22 9 9 7 9 13 9 13 13 9 9 13 3 0 9 7 13 3 3 13 0 9 2
24 2 12 2 9 13 9 7 9 13 0 9 13 3 13 2 16 15 9 9 9 9 4 13 2
17 15 9 13 9 7 9 13 9 13 9 13 9 13 9 0 9 2
9 15 9 4 13 15 9 9 0 2
10 15 9 13 13 9 13 9 9 1 2
36 2 12 2 11 0 9 4 13 9 2 9 2 9 12 2 12 2 3 13 9 9 2 15 13 9 7 9 0 9 7 15 13 9 9 9 2
31 3 9 13 3 9 9 9 13 0 9 13 9 9 2 15 13 9 9 0 9 2 7 9 2 9 2 15 9 3 13 2
13 16 13 9 15 9 9 2 9 9 9 13 0 2
39 2 12 2 13 0 13 0 9 2 16 13 0 9 9 3 7 3 9 2 3 7 9 9 9 2 9 7 9 1 2 16 15 9 13 0 9 9 9 2
10 15 13 9 2 15 3 13 3 3 2
15 2 12 2 13 3 13 0 9 7 15 9 9 7 9 2
31 13 9 9 13 9 13 15 9 2 15 13 9 2 15 9 9 9 7 9 9 2 9 7 15 0 9 2 3 9 9 2
24 2 12 2 13 0 13 9 9 2 9 13 2 3 13 7 0 9 9 13 15 13 9 9 2
7 3 9 9 4 13 9 2
21 2 12 2 9 13 0 9 2 9 2 13 7 13 9 2 9 13 9 2 9 2
15 15 9 13 9 13 9 13 9 7 13 15 0 9 1 2
9 0 9 4 3 13 9 9 9 2
17 2 12 2 9 9 4 13 9 9 2 15 13 0 9 13 9 2
5 4 13 15 9 2
2 12 9
1 9
34 15 9 9 2 9 2 2 2 9 13 9 2 7 2 15 9 13 2 13 15 9 16 15 4 13 9 2 9 2 9 12 12 9 2
2 12 9
3 0 9 9
12 0 0 9 9 13 9 13 9 9 13 9 2
48 9 1 9 13 9 13 9 2 3 16 15 4 13 9 9 2 7 15 15 9 13 9 2 15 13 3 9 7 15 0 9 15 16 9 7 13 9 7 13 9 0 9 2 3 0 9 2 2
32 0 0 9 4 13 0 9 9 9 2 16 13 9 1 13 9 9 13 3 12 9 15 9 13 9 15 9 9 13 13 9 2
22 0 9 13 15 9 9 3 3 2 16 15 4 13 13 7 13 9 15 9 9 1 2
2 12 9
4 9 13 9 9
34 0 11 13 7 13 9 0 13 12 9 0 9 13 9 3 9 13 9 9 13 9 0 9 11 9 9 13 9 9 7 9 13 9 2
12 9 13 9 9 9 7 9 13 11 9 9 2
28 0 11 7 0 9 13 9 13 9 9 7 15 9 0 9 0 9 2 3 3 11 1 7 0 9 9 9 2
10 0 9 13 9 9 4 13 3 9 2
37 16 12 9 0 9 0 13 13 9 13 3 0 2 11 13 13 9 9 2 15 13 4 3 13 9 15 9 16 15 4 0 9 13 0 9 9 2
2 12 9
3 9 13 9
36 0 9 13 9 0 9 9 7 9 0 9 9 13 3 9 9 9 7 9 9 2 9 7 9 9 13 9 9 15 9 9 2 15 9 13 2
8 15 9 13 9 13 3 9 2
10 0 13 9 4 13 15 9 9 0 2
22 0 13 9 13 15 9 9 0 13 9 9 2 9 2 0 9 7 9 13 9 3 2
20 0 0 9 13 7 13 0 9 9 13 15 9 2 15 0 9 9 4 13 2
34 0 9 13 2 16 15 9 13 13 9 7 16 15 9 4 3 13 3 12 9 0 9 9 2 9 2 0 9 7 9 13 9 9 2
17 0 9 12 9 12 9 13 9 9 13 13 9 9 13 9 3 2
23 2 15 9 2 15 13 0 9 2 13 0 9 2 0 16 15 4 13 15 9 9 0 2
24 2 15 0 9 2 15 13 13 9 2 13 0 9 2 0 16 15 4 13 15 9 9 0 2
14 0 9 4 13 13 13 9 7 13 15 1 9 3 2
26 0 0 9 4 13 9 9 9 9 9 13 9 9 13 9 2 15 3 13 12 9 12 9 13 9 2
29 0 0 9 4 13 9 9 9 9 7 9 9 7 13 15 9 3 13 3 13 9 9 2 13 16 0 9 13 2
29 2 9 13 0 9 0 9 9 2 3 13 0 9 15 2 3 0 9 15 3 13 0 9 4 13 0 9 13 2
22 2 16 4 13 0 9 2 0 9 13 9 13 9 13 9 15 9 2 15 9 13 2
59 0 16 9 13 9 7 9 7 15 9 2 15 4 13 9 13 9 9 2 9 13 2 15 1 16 9 0 9 9 4 13 0 2 7 3 16 9 7 9 4 13 3 2 0 0 9 13 9 2 15 3 15 9 13 9 13 9 13 2
2 12 9
13 13 9 9 9 2 9 2 9 12 2 12 2 3
49 0 15 9 13 15 9 3 13 9 9 9 9 9 12 9 9 12 13 11 9 9 2 9 2 9 12 2 12 2 2 12 2 3 2 0 16 15 13 13 9 2 9 2 9 12 2 12 2 2
14 15 9 13 15 9 3 13 2 13 15 9 9 9 2
38 0 9 0 9 4 9 2 9 2 9 12 2 12 2 12 9 13 9 3 13 9 9 7 9 15 3 13 9 15 9 12 9 7 9 0 13 9 2
14 0 11 9 9 13 9 7 9 13 15 9 9 0 2
16 15 9 9 13 9 2 9 2 9 12 2 12 2 9 1 2
2 9 9
2 9 12
20 0 9 11 9 13 9 2 3 0 9 9 13 3 13 9 13 9 7 9 2
2 9 9
19 9 13 9 2 16 0 9 9 13 0 9 1 11 9 9 9 0 9 2
11 9 13 3 3 2 16 9 13 13 9 2
16 9 9 13 3 13 7 13 3 3 0 9 13 0 13 13 2
17 15 9 13 9 0 9 2 15 4 13 3 0 9 3 7 9 2
7 9 13 3 0 9 9 2
14 9 9 9 9 9 13 3 0 2 3 9 13 0 2
15 9 13 12 0 9 2 7 9 13 3 13 15 9 9 2
19 11 9 9 13 9 13 2 9 11 1 13 11 9 13 9 0 9 9 2
38 15 9 13 3 0 9 13 9 9 7 15 9 7 9 1 13 0 9 15 15 15 0 9 9 13 3 7 9 1 7 9 7 15 9 9 3 13 2
2 0 9
14 13 9 9 3 15 2 15 9 13 3 15 9 0 2
7 15 13 3 11 9 13 2
19 13 15 9 9 9 1 2 11 9 11 13 0 9 9 2 2 13 2 2
2 9 3
3 13 9 12
14 3 3 0 9 1 0 9 3 11 7 9 9 9 2
22 0 9 13 9 3 0 9 13 9 9 7 15 9 13 13 3 11 9 9 9 9 2
15 9 7 9 4 13 3 7 9 0 9 4 3 3 13 2
17 9 13 3 3 12 2 7 3 9 9 13 3 9 13 2 8 2
4 9 3 8 2
9 8 8 8 8 8 8 2 8 2
24 9 13 3 0 7 0 9 3 13 2 7 9 9 9 11 5 11 13 13 0 13 15 9 2
12 3 11 9 4 13 13 9 13 9 0 9 2
11 6 2 15 13 15 13 2 8 2 8 2
14 3 13 0 9 0 9 9 9 7 0 9 9 9 2
13 9 1 3 9 4 13 11 7 11 13 9 9 2
15 9 13 7 13 2 7 0 9 13 0 9 7 0 9 2
15 9 13 3 9 2 9 7 3 3 12 9 1 13 9 2
18 9 4 4 13 3 2 7 3 3 9 0 9 13 3 9 13 9 2
21 15 13 11 9 13 0 9 0 9 2 7 2 0 9 15 3 13 2 0 9 2
6 13 15 13 2 8 2
7 6 11 13 9 2 8 2
24 9 7 9 1 0 9 13 11 9 2 15 11 9 4 3 13 13 9 1 9 0 9 9 2
25 9 9 9 9 4 13 2 7 3 15 13 4 4 13 13 11 11 9 13 7 9 9 13 9 2
10 0 9 13 9 13 9 3 9 2 8
6 2 9 0 2 8 2
14 9 13 13 11 11 2 7 9 13 3 1 9 13 2
23 9 2 9 2 4 13 1 3 0 11 11 11 2 7 9 3 13 13 15 13 15 9 2
29 13 3 3 2 16 11 9 4 3 13 13 9 3 7 3 7 0 9 9 2 7 13 4 3 13 13 0 9 2
19 13 3 13 2 13 9 13 2 16 9 9 9 13 9 13 9 0 9 2
17 7 3 2 15 9 7 15 9 2 0 9 7 9 3 0 9 2
2 6 2
4 9 2 11 9
4 9 13 9 13
6 11 9 9 0 9 2
13 9 13 9 2 13 9 9 7 13 9 9 3 2
4 7 15 9 2
22 9 1 1 11 13 12 11 9 2 15 13 3 9 13 2 7 3 0 3 1 11 2
17 9 4 13 15 9 2 16 12 0 9 9 4 13 11 1 9 2
15 3 3 11 0 9 13 9 9 4 13 3 3 11 9 2
13 11 11 7 11 11 13 15 3 11 11 9 9 2
13 13 9 9 2 9 7 9 7 13 9 1 13 2
26 9 7 9 1 13 3 9 7 13 2 15 3 13 11 0 9 2 7 3 0 9 4 11 9 13 2
3 9 13 0
13 3 9 13 2 16 15 3 0 9 13 13 9 2
18 11 13 9 12 9 2 7 3 9 9 13 9 9 13 12 12 9 2
26 11 9 13 9 9 0 12 2 7 9 13 0 9 2 7 9 12 9 13 9 13 0 12 0 9 2
12 9 9 9 13 12 2 11 2 11 7 11 2
9 3 15 11 3 13 0 9 13 2
22 11 7 11 13 2 16 11 9 13 3 12 9 2 9 9 2 9 7 9 7 9 2
18 15 9 13 9 9 3 0 9 9 2 7 9 9 13 3 3 0 2
12 11 9 13 3 7 15 13 9 7 0 9 2
17 0 9 15 0 9 13 9 13 3 11 2 11 2 11 7 11 2
7 9 9 4 13 9 9 2
28 2 16 13 0 9 1 2 13 0 13 9 1 13 9 9 2 2 11 9 13 7 15 1 9 13 11 13 2
4 15 15 13 2
8 9 11 9 15 9 13 3 2
15 9 1 9 13 0 9 13 9 13 0 9 9 1 13 2
18 2 16 15 13 9 2 13 0 0 9 9 2 2 11 13 11 13 2
11 15 13 13 3 0 9 9 2 3 9 2
10 9 13 3 2 7 9 7 9 9 2
10 11 13 13 3 0 9 9 9 9 2
25 9 9 13 9 9 13 3 9 2 9 9 2 9 9 2 9 2 9 7 3 0 9 9 1 2
12 7 11 7 11 13 3 3 11 9 13 9 2
29 3 15 1 2 16 9 13 3 3 9 2 13 3 13 9 2 15 13 13 2 2 2 7 9 9 3 3 13 2
8 3 9 13 3 11 9 13 2
11 2 9 13 13 3 3 2 2 11 13 2
22 0 9 13 11 9 9 2 7 9 9 13 9 9 3 7 3 2 7 15 13 9 2
18 9 11 13 11 7 11 1 0 9 9 9 7 3 9 13 15 3 2
16 0 13 9 13 13 2 7 3 15 15 4 13 0 13 9 2
10 11 9 13 0 9 7 15 3 13 2
7 3 13 3 3 3 13 2
24 2 0 9 13 3 13 9 16 15 0 9 2 15 15 13 15 9 13 13 2 2 11 13 2
23 9 9 9 13 0 9 13 11 1 3 9 7 9 0 9 2 7 3 9 7 9 13 2
23 9 13 15 9 2 7 15 1 13 13 9 13 15 0 9 2 3 9 2 9 7 9 2
12 9 13 9 2 7 0 9 9 13 4 13 2
6 8 8 8 2 8 8
17 11 9 11 11 13 9 9 1 13 13 9 9 9 15 9 3 2
20 16 0 9 9 13 0 9 9 9 2 13 3 15 9 3 1 13 0 9 2
21 15 1 9 0 9 9 13 0 9 2 9 0 9 9 7 0 9 9 13 9 2
23 3 9 13 9 13 13 3 0 9 2 7 13 0 9 1 13 9 13 15 3 0 9 2
30 0 7 0 0 9 13 9 15 4 3 13 15 9 3 2 3 16 9 13 3 9 2 3 15 9 2 3 15 3 2
21 0 0 9 9 13 2 7 15 13 3 0 9 2 3 9 7 9 1 13 9 2
6 9 1 13 3 9 2
12 13 9 2 16 3 11 4 9 13 9 11 2
4 9 13 0 2
13 2 9 13 3 0 9 2 15 4 13 3 9 2
10 11 0 13 0 13 2 2 11 13 2
17 2 16 3 11 13 0 9 2 15 13 13 15 0 9 9 2 2
3 3 9 1
17 16 3 13 4 13 9 9 9 2 13 11 0 9 13 0 9 2
7 15 4 13 9 13 9 2
21 9 1 3 12 9 13 0 9 3 13 9 0 9 2 7 11 9 9 13 0 2
23 2 15 9 13 15 1 2 3 9 13 15 15 2 13 9 13 9 1 9 7 9 2 2
22 16 9 13 0 2 13 15 13 15 9 1 2 15 1 9 13 12 3 9 0 9 2
31 16 15 13 3 2 3 13 9 3 0 9 2 7 16 15 1 13 4 13 13 9 0 9 2 4 9 13 9 3 3 2
16 16 13 13 3 13 0 9 2 3 9 9 7 9 13 9 2
8 11 13 0 9 13 0 3 2
10 2 9 9 13 0 9 13 0 9 2
12 11 13 3 9 1 7 9 13 3 9 9 2
15 15 1 15 0 9 13 3 9 7 0 9 3 9 2 2
8 11 9 13 3 13 9 9 2
31 16 11 4 13 3 3 11 11 11 11 11 11 13 9 11 0 9 0 9 9 2 13 3 9 3 4 13 0 9 9 2
6 3 15 0 9 13 2
20 2 3 4 3 13 0 9 2 16 9 13 3 2 2 11 13 12 9 9 2
23 2 3 3 4 3 13 9 15 0 9 2 15 13 15 9 13 3 2 2 13 11 3 2
9 2 3 15 15 9 4 13 2 2
4 11 11 13 9
2 0 9
13 9 12 9 11 13 15 9 13 9 1 0 0 2
21 11 7 11 9 13 3 9 3 0 9 7 13 3 9 0 9 11 11 9 12 2
9 0 9 13 16 9 13 9 9 2
16 0 7 0 9 11 11 13 9 9 12 16 9 9 13 3 2
33 9 15 9 2 15 4 13 11 12 7 13 9 12 2 7 13 13 16 12 13 0 9 0 9 2 11 11 7 11 11 2 9 2
26 1 9 13 3 3 9 11 11 2 11 2 11 11 2 0 9 9 2 11 12 2 9 7 11 11 2
5 0 9 7 15 9
10 0 9 4 13 9 9 3 0 13 2
9 0 9 4 3 3 13 9 1 2
17 9 13 3 13 13 3 2 3 13 13 3 9 7 3 13 9 2
7 15 9 13 0 9 9 2
6 3 9 13 13 9 2
19 9 3 0 9 13 15 2 16 9 13 15 9 13 2 9 13 3 0 2
26 3 3 9 9 2 7 6 15 15 2 3 15 0 9 13 3 9 2 16 13 13 3 9 3 0 2
18 0 9 13 3 11 2 9 7 11 11 2 15 3 13 0 0 9 2
21 0 9 11 11 7 11 11 13 0 9 2 15 9 0 9 2 13 0 9 2 2
21 16 9 13 9 3 0 2 4 9 13 3 0 16 0 11 13 9 9 0 9 2
2 9 9
16 0 9 9 13 9 13 9 13 9 7 13 3 13 9 9 2
21 16 13 4 13 9 2 4 13 0 9 9 16 11 3 13 2 13 13 9 3 2
11 9 13 3 15 9 9 7 15 13 13 2
13 9 1 0 9 13 11 9 1 13 11 11 9 2
10 9 13 11 9 9 7 13 3 9 2
23 11 9 13 3 9 2 16 9 13 3 15 9 16 9 0 9 9 9 1 13 9 9 2
32 11 11 9 13 3 0 2 7 11 11 2 11 11 7 11 11 7 11 11 1 4 13 13 11 11 2 15 13 3 9 11 2
20 13 11 9 15 3 2 13 15 11 7 11 9 0 9 9 2 3 15 9 2
2 9 9
25 9 13 13 3 13 7 16 9 13 3 0 7 9 0 2 13 9 13 13 11 9 13 7 13 2
17 9 9 13 3 11 11 13 9 12 3 2 9 9 13 12 9 2
19 11 9 9 13 15 9 11 11 2 15 13 0 9 7 9 3 15 9 2
13 9 13 0 13 7 15 13 13 15 0 0 9 2
15 3 13 15 9 9 13 11 9 2 15 13 13 0 9 2
25 15 3 13 9 9 9 7 13 3 2 0 9 0 9 2 9 9 9 2 9 9 13 9 9 2
2 9 9
13 0 0 9 4 3 13 9 9 11 9 11 11 2
10 9 13 15 9 1 0 11 9 9 2
5 9 13 15 9 2
19 15 0 9 3 3 3 0 9 13 0 9 2 15 4 13 9 9 9 2
4 3 0 0 2
14 9 9 13 13 13 2 16 13 9 13 13 13 9 2
5 9 13 3 11 2
3 0 9 2
10 9 7 9 9 9 13 3 13 9 2
29 15 13 4 13 9 9 13 0 9 2 7 13 13 13 9 16 15 13 3 0 13 9 7 0 9 7 3 0 2
23 9 13 3 13 0 9 1 2 7 9 13 0 13 0 7 0 9 13 9 3 13 9 2
3 12 9 12
9 13 9 13 3 9 11 9 1 2
13 9 13 13 0 16 13 9 9 7 13 12 9 2
17 9 13 0 9 9 13 13 9 2 3 0 9 4 13 9 9 2
14 9 9 15 9 4 13 9 2 15 3 13 13 13 2
15 9 13 0 0 9 2 15 1 13 3 13 15 9 13 2
15 13 9 1 9 12 9 9 9 2 12 9 2 9 0 2
35 9 13 9 9 9 13 2 15 13 15 9 3 3 16 13 13 9 2 3 13 9 12 0 2 9 9 7 0 9 9 0 9 9 2 2
6 9 13 13 3 3 2
14 13 15 9 9 7 13 3 3 13 15 9 0 9 2
9 0 12 9 13 3 3 9 13 2
6 9 13 3 3 12 2
9 0 9 13 9 13 12 9 1 2
21 3 12 9 9 13 15 9 9 1 2 13 9 1 7 13 3 0 12 9 9 2
15 0 13 9 0 9 2 7 9 13 3 0 9 15 9 2
24 0 13 9 2 0 9 13 3 2 15 12 9 9 9 13 4 13 15 15 13 4 13 9 2
2 9 2
4 0 9 13 2
15 11 9 13 9 13 9 7 13 0 9 1 13 9 13 2
17 15 0 9 13 9 9 9 9 7 13 9 16 13 13 0 9 2
14 15 13 9 15 0 9 2 9 13 9 13 0 9 2
9 9 9 13 3 15 13 0 9 2
10 13 9 9 9 7 13 3 13 9 2
4 13 13 9 2
2 15 9
22 11 9 9 9 7 9 13 13 3 0 9 13 9 9 9 7 15 1 9 13 9 2
9 9 9 9 9 13 13 15 9 2
19 9 13 3 12 9 13 3 3 2 16 9 4 13 7 9 9 13 0 2
20 15 9 9 13 12 9 2 15 12 13 16 15 13 9 2 7 12 13 9 2
6 15 12 13 15 9 2
15 12 9 13 13 9 2 7 15 9 16 15 13 3 3 2
39 9 13 3 9 2 15 4 13 9 9 9 7 3 9 0 2 9 13 9 0 9 13 13 9 2 7 9 9 1 13 0 2 16 15 13 9 3 3 2
6 15 13 0 9 9 2
58 9 9 13 2 12 9 2 0 9 2 9 2 12 5 2 2 0 9 2 8 8 2 2 0 9 9 2 9 11 2 12 5 2 2 9 2 11 9 2 12 5 2 2 9 2 15 11 13 9 7 15 15 13 2 16 3 13 2
16 9 11 0 2 13 2 13 3 9 2 13 13 13 9 1 2
22 9 2 9 13 2 2 15 4 3 13 13 13 15 2 13 0 9 9 7 9 9 2
4 9 13 9 2
9 9 9 7 11 9 11 12 2 12
18 9 0 2 9 2 13 3 9 9 9 2 15 0 9 13 9 11 2
15 11 0 9 9 13 15 9 13 3 12 9 7 9 9 2
8 9 9 13 3 12 9 9 2
16 15 9 9 13 11 0 9 3 9 13 0 2 7 15 0 2
9 9 9 9 13 13 3 9 9 2
10 9 13 9 9 7 13 9 9 9 2
4 9 13 3 2
9 11 13 9 9 13 13 0 9 2
6 11 13 0 3 9 2
8 11 13 9 13 9 0 9 2
3 13 9 2
10 9 13 9 13 3 9 2 11 11 2
11 13 3 9 2 15 9 13 9 9 9 2
7 13 0 9 9 13 9 2
13 3 9 4 13 9 2 15 3 13 0 9 1 2
8 3 13 9 0 9 2 9 2
22 9 3 3 13 9 7 0 9 0 9 13 9 9 13 0 16 15 0 9 4 13 2
19 9 3 13 13 9 9 9 9 13 9 11 2 15 13 13 15 9 9 2
22 9 13 9 9 13 7 3 9 11 13 13 9 1 9 2 15 13 3 9 9 9 2
5 9 13 9 0 2
6 9 13 0 9 9 2
12 9 13 3 9 16 15 9 13 3 13 3 2
7 15 13 3 9 13 9 2
13 3 13 9 1 13 9 9 8 8 7 11 9 2
20 9 9 4 3 13 9 13 9 16 0 13 3 9 13 9 3 0 9 13 2
12 9 13 0 9 3 4 3 3 13 1 9 2
4 9 7 9 13
7 9 13 9 7 9 9 2
6 0 9 13 9 9 2
10 15 0 9 13 3 0 11 9 9 2
7 9 13 3 13 13 9 2
12 3 0 9 13 9 1 7 13 13 9 9 2
8 0 9 4 13 9 15 9 2
14 9 9 13 0 16 11 4 13 9 9 15 9 13 2
6 0 9 2 6 6 2
5 0 9 13 9 2
25 9 13 13 9 9 13 9 2 9 13 9 2 15 3 12 9 1 13 9 2 15 4 13 9 2
12 9 13 9 1 0 9 13 9 7 0 9 2
12 9 13 9 13 7 3 13 9 13 9 9 2
7 11 7 11 9 13 9 2
7 4 13 9 9 2 6 2
11 9 0 9 9 13 9 0 13 9 11 2
10 9 4 13 0 9 7 9 13 0 2
10 0 9 9 7 3 9 1 13 9 2
6 0 9 9 13 9 2
7 3 13 12 9 15 9 2
8 9 13 7 13 3 9 9 2
10 0 9 4 13 9 15 9 13 13 2
6 3 9 13 13 9 2
11 9 9 13 0 9 9 9 13 9 1 2
12 0 9 4 13 2 15 13 12 9 3 2 2
11 11 4 3 13 15 9 1 9 0 9 2
7 0 9 13 3 0 15 2
12 9 15 12 9 13 0 9 9 13 9 1 2
23 9 13 13 1 9 11 9 13 9 7 13 15 9 7 3 13 9 7 13 15 9 9 2
9 9 4 13 9 13 9 1 9 2
20 9 1 15 9 13 9 12 9 2 7 9 1 9 9 13 12 9 1 9 2
8 11 13 9 3 13 11 9 2
10 9 13 13 13 12 1 12 9 1 2
16 0 9 13 3 0 0 9 1 0 9 7 11 9 13 9 2
9 11 13 15 9 9 7 3 13 2
2 9 9
10 13 9 13 9 2 15 13 9 9 2
10 9 13 13 2 7 9 9 13 9 2
16 9 9 11 9 13 0 2 11 9 13 0 3 3 9 12 2
10 9 9 13 3 2 9 9 13 13 2
16 9 13 3 0 9 2 16 0 9 4 13 3 16 0 9 2
9 9 9 4 13 15 13 3 9 2
11 11 13 3 3 9 9 7 13 9 3 2
12 9 1 13 16 11 4 13 15 0 11 9 2
3 9 15 2
5 9 13 9 9 2
9 15 9 9 1 13 9 3 11 2
5 9 13 3 12 2
3 9 11 9
1 9
10 11 9 13 11 9 9 0 9 9 2
6 9 13 12 9 3 2
9 9 13 9 7 13 9 9 9 2
10 3 9 9 13 9 2 9 7 9 2
15 13 9 13 15 9 15 9 3 16 0 9 13 13 3 2
11 9 11 9 9 13 3 12 0 9 9 2
20 9 9 13 3 9 16 9 4 13 3 9 9 7 9 13 3 9 3 9 2
16 9 13 3 1 0 15 9 9 13 13 12 9 13 9 3 2
7 0 9 13 9 9 1 2
20 3 9 0 9 7 0 9 9 2 9 13 0 9 9 13 3 12 11 9 2
21 9 13 3 3 2 7 9 9 2 12 12 1 2 13 3 11 9 0 9 12 2
9 0 9 9 13 0 7 3 13 2
10 1 13 15 9 3 12 9 3 9 2
4 9 13 11 2
14 0 9 11 9 13 3 3 9 7 9 13 0 9 2
11 0 9 9 9 13 2 7 9 13 13 2
24 9 9 7 9 3 13 15 9 13 11 9 9 0 9 13 9 2 15 13 3 13 0 9 2
12 0 9 13 3 9 9 7 9 9 13 9 2
19 9 13 9 13 3 0 2 0 9 13 9 9 7 0 9 13 3 9 2
5 0 13 11 9 2
5 9 13 9 12 2
7 0 9 13 3 9 1 2
14 9 13 9 13 0 9 3 3 7 9 13 3 15 2
10 9 13 7 3 13 0 7 0 9 2
14 9 0 9 13 13 7 9 13 3 13 0 9 9 2
6 9 13 3 12 9 2
8 15 13 3 9 9 0 9 2
12 9 13 3 3 7 9 13 3 0 0 9 2
3 9 13 0
6 3 11 13 9 1 2
17 9 13 15 9 9 2 16 9 9 9 13 4 13 0 9 9 2
7 0 9 3 13 0 9 2
14 9 4 3 13 7 9 7 9 7 9 13 15 13 2
14 9 13 13 0 9 2 3 9 13 12 11 9 0 2
11 9 9 13 7 0 9 13 13 3 0 2
5 9 13 9 12 2
7 11 11 13 3 0 9 2
24 3 9 1 13 0 2 16 9 9 13 0 3 3 7 9 13 3 3 9 9 11 9 9 2
15 3 13 11 9 15 9 2 7 9 13 3 0 9 1 2
8 9 11 12 9 2 11 12 2
9 9 0 9 9 13 9 0 9 2
6 3 13 0 9 9 2
16 11 13 3 12 9 9 3 3 9 4 13 15 9 0 9 2
5 9 13 3 0 2
9 3 0 9 13 12 9 9 9 2
11 9 9 13 0 9 15 9 3 3 13 2
15 9 0 9 15 9 2 13 2 9 13 3 3 15 3 2
7 9 13 3 12 9 9 2
11 9 9 9 13 9 1 3 0 9 9 2
10 13 12 9 9 2 16 9 13 9 2
16 16 9 13 13 9 15 9 2 3 9 9 13 4 3 13 2
10 9 13 3 0 7 9 4 13 9 2
11 15 9 11 13 0 7 13 9 9 12 2
1 9
13 11 9 7 9 9 13 9 2 15 13 0 9 2
7 11 9 13 3 9 9 2
6 9 13 1 12 9 2
13 9 13 12 12 9 7 9 13 3 3 9 1 2
10 9 13 9 7 12 9 12 12 1 2
18 9 11 9 13 9 9 3 0 9 2 13 0 9 11 7 13 11 2
6 9 13 3 9 11 2
13 11 13 9 3 0 0 9 7 9 13 3 3 2
13 3 11 13 9 7 13 9 2 15 3 13 11 2
14 9 9 9 13 3 0 2 7 9 13 0 9 9 2
10 11 13 3 3 13 9 12 9 9 2
7 11 13 3 9 9 3 2
14 16 9 13 9 3 2 9 13 3 9 3 9 0 2
15 3 11 9 13 13 9 7 9 13 13 9 9 9 1 2
12 9 13 3 11 2 7 0 9 13 3 9 2
4 0 9 9 12
16 11 9 0 9 9 9 2 11 2 13 9 12 0 9 9 2
23 11 13 3 11 11 13 9 2 15 9 13 13 0 9 9 7 13 3 9 9 15 9 2
9 15 9 11 13 0 9 9 9 2
14 9 13 9 3 12 0 9 7 0 9 9 9 9 2
27 9 9 13 9 3 11 9 11 2 11 2 11 7 9 7 9 11 9 2 11 11 7 11 11 11 9 2
13 9 9 9 13 13 12 9 7 12 12 9 9 2
2 9 9
10 9 9 13 11 11 11 11 11 11 2
12 9 9 13 11 9 0 9 2 3 9 9 2
18 9 13 9 0 9 15 2 15 15 11 3 13 7 15 15 13 3 2
20 9 13 3 11 1 13 9 9 15 9 7 9 2 7 3 15 0 9 13 2
12 11 11 1 9 13 11 11 9 0 11 11 2
12 11 11 13 7 13 0 9 1 11 9 9 2
29 9 13 3 9 7 9 9 2 15 9 9 7 0 9 4 13 2 7 3 3 13 15 13 9 7 9 7 9 2
19 3 0 13 3 11 11 11 11 0 9 11 12 2 15 13 3 11 9 2
12 3 9 13 9 11 7 9 15 9 13 9 2
4 9 7 13 9
11 9 13 9 0 9 9 13 11 9 9 2
9 11 13 0 9 7 9 13 9 2
12 11 11 11 13 0 9 0 7 0 9 9 2
18 3 9 13 3 3 0 9 9 2 13 0 7 0 9 13 3 3 2
19 3 9 13 15 2 13 0 9 9 9 1 13 0 9 0 3 9 9 2
9 9 1 9 13 11 9 11 11 2
24 11 9 13 2 3 9 9 2 9 0 9 15 2 3 0 9 7 11 13 0 9 13 9 2
17 9 13 0 9 2 9 7 9 9 2 15 13 9 1 13 3 2
9 3 13 3 3 11 9 15 9 2
9 11 9 13 3 3 0 9 9 2
3 9 0 9
14 0 9 1 0 13 3 9 13 9 7 9 9 9 2
15 9 13 9 12 9 9 0 2 3 3 9 9 13 2 9
13 9 9 13 3 11 9 9 7 0 0 9 11 2
18 3 3 0 9 9 13 0 2 3 3 9 9 1 13 9 9 13 2
14 9 13 3 11 9 9 2 15 11 9 4 11 13 2
18 13 3 15 2 15 15 9 13 3 0 9 13 2 13 9 0 9 2
2 13 15
9 0 9 2 15 13 13 3 0 2
21 4 13 9 13 15 0 9 2 9 9 3 7 3 13 13 0 9 9 13 15 2
14 7 3 13 15 0 9 2 15 9 13 3 0 9 2
10 9 13 4 3 13 3 0 7 0 2
9 7 3 15 9 4 13 13 15 2
28 9 3 4 13 9 2 3 0 4 13 3 9 9 7 15 0 9 2 15 0 9 4 13 15 0 9 9 2
15 0 9 13 0 9 3 0 9 3 9 9 9 9 9 2
9 9 13 3 9 3 3 0 9 2
5 6 3 15 9 2
18 15 15 1 4 13 7 1 15 2 15 15 0 13 3 9 9 3 2
4 6 6 13 2
24 15 4 9 1 13 9 0 9 9 15 9 0 9 9 2 13 15 3 9 9 7 0 9 2
16 9 1 15 11 9 13 9 1 3 15 0 7 0 0 9 2
20 15 11 4 13 9 13 13 11 9 1 9 3 15 9 7 13 11 0 9 2
11 9 4 13 13 0 12 9 15 3 13 2
10 13 2 16 15 9 13 15 0 9 2
15 3 9 4 13 0 2 15 13 3 0 9 9 9 9 2
6 3 13 0 9 9 2
23 4 9 9 13 15 9 9 13 11 9 9 7 9 9 2 9 7 9 9 9 9 13 2
15 13 13 2 16 9 13 0 9 3 15 1 7 15 0 2
19 9 9 13 0 13 15 13 15 2 7 4 13 0 15 0 9 9 9 2
19 11 13 9 9 3 0 9 2 15 0 9 9 13 9 9 9 13 9 2
10 9 13 3 9 9 13 0 11 9 2
8 9 13 9 9 11 9 9 2
12 9 11 4 13 9 9 11 11 0 9 9 2
25 9 9 13 3 3 9 9 13 9 9 7 9 9 9 9 9 9 2 9 2 9 7 11 9 2
9 9 13 9 11 13 9 9 9 2
15 0 9 13 3 9 7 9 2 15 11 13 3 12 9 2
27 3 13 11 4 15 9 13 9 2 16 0 11 11 13 9 0 0 9 13 7 0 9 13 9 13 9 2
20 3 9 9 15 9 13 3 15 15 9 13 9 3 13 9 9 11 11 9 2
36 9 13 13 3 12 0 0 2 16 9 4 15 9 13 2 16 9 9 9 11 9 13 3 13 3 9 9 9 9 13 3 0 9 9 9 2
12 3 3 11 13 3 9 15 0 9 0 9 2
17 9 4 13 15 3 3 3 9 7 3 9 13 13 9 9 1 2
16 13 15 13 9 2 16 13 9 0 0 9 7 15 9 9 2
28 13 13 2 13 9 2 7 3 1 15 2 13 9 9 7 13 13 3 0 13 9 9 9 3 13 3 9 2
12 15 13 9 2 7 13 13 13 3 0 9 2
17 11 13 13 15 1 7 3 3 9 0 9 9 9 7 9 13 2
6 13 9 7 13 9 2
6 3 3 9 7 9 2
9 13 15 7 3 2 16 13 15 2
2 9 9
6 13 9 15 0 9 2
7 13 0 9 9 9 9 2
19 4 3 13 9 9 3 2 16 13 13 13 9 7 13 9 1 13 9 2
28 3 13 13 15 9 9 0 9 1 9 2 7 9 0 9 7 9 0 9 13 15 13 9 1 3 12 9 2
26 9 13 3 0 13 3 9 9 13 15 2 13 13 3 13 9 2 4 3 13 9 13 0 9 15 2
37 9 0 9 13 0 9 11 9 9 2 7 9 13 15 9 13 12 9 9 13 0 9 7 15 13 9 1 2 15 1 13 9 3 9 0 9 2
5 2 13 13 2 2
18 0 9 9 9 13 15 9 13 9 2 9 9 9 7 15 0 9 2
38 3 9 1 13 13 15 2 16 9 13 15 7 9 3 13 9 2 9 7 9 2 7 3 13 13 15 9 2 15 13 15 13 2 3 0 4 13 2
29 11 11 13 0 9 7 9 2 15 13 9 3 0 9 9 16 15 2 7 15 3 13 9 13 9 11 9 9 2
30 11 13 2 16 0 9 13 0 9 9 13 0 9 2 0 9 7 9 2 7 3 13 3 3 3 13 9 7 9 2
13 3 16 13 9 3 3 2 16 15 13 3 13 2
16 16 13 9 3 9 7 15 9 2 7 13 9 3 9 1 2
22 11 1 13 9 3 2 16 0 9 13 7 0 9 13 13 9 3 9 0 9 9 2
30 9 9 9 2 11 11 11 2 12 2 11 13 9 7 13 15 0 9 2 13 9 2 3 13 9 2 9 7 9 2
27 15 1 16 13 15 0 9 3 13 9 9 2 13 15 13 9 2 13 0 9 9 7 13 13 0 9 2
6 11 13 13 9 3 2
18 9 9 4 13 9 0 0 7 0 2 7 9 13 0 9 9 9 2
24 9 2 15 9 9 3 13 9 2 4 13 9 13 9 0 9 2 3 9 0 7 0 9 2
23 9 13 15 9 2 3 9 13 0 9 9 2 15 13 7 9 9 2 3 9 7 9 2
8 0 9 4 13 3 3 9 2
15 9 4 3 13 0 9 9 2 15 0 9 13 13 9 2
35 3 13 7 3 13 9 4 3 13 9 2 13 9 3 16 3 13 7 13 9 13 9 2 7 3 9 9 13 9 9 0 13 3 0 2
19 9 13 9 9 0 9 2 7 0 13 15 2 16 13 15 2 15 13 2
25 3 9 9 9 13 9 2 16 15 13 3 0 7 13 3 9 2 0 9 15 13 9 7 9 2
56 15 9 9 3 9 9 13 3 9 11 11 9 9 11 11 11 11 2 12 2 2 2 13 15 13 15 2 16 15 13 3 3 9 2 13 3 9 2 15 9 13 9 7 13 9 7 9 3 2 7 3 9 13 2 2 2
33 3 9 13 3 3 9 9 13 0 9 2 15 9 13 13 9 2 7 1 13 13 0 7 0 9 7 9 0 7 0 9 1 2
23 0 9 9 2 16 0 7 3 0 13 2 13 9 9 0 9 9 0 7 3 0 9 2
15 15 3 13 4 2 13 4 13 13 15 15 13 0 9 2
35 16 0 3 13 13 1 9 9 2 13 3 9 1 7 13 9 0 9 11 2 4 13 0 9 7 13 0 9 2 9 13 3 8 8 2
7 9 9 4 15 9 13 2
19 13 3 2 3 3 13 13 0 2 0 9 1 13 2 15 15 13 9 2
17 9 13 0 2 16 9 13 0 7 0 9 2 15 9 13 9 2
19 16 13 13 2 15 9 13 9 7 13 2 13 2 16 0 9 15 13 2
10 15 13 13 9 2 15 13 15 9 2
36 16 3 13 0 13 2 13 9 9 7 9 2 7 13 15 9 7 9 2 13 13 15 9 3 2 16 13 15 13 9 2 9 9 7 9 2
11 15 9 13 9 2 9 13 9 0 9 2
5 13 13 13 3 2
8 3 2 13 15 3 9 9 2
27 13 15 3 3 9 2 3 9 9 2 15 1 16 13 13 3 13 9 2 9 7 11 11 9 0 9 2
21 9 13 3 0 9 9 2 16 15 15 13 13 13 9 13 4 9 3 13 15 2
19 16 3 13 9 9 3 9 1 2 13 0 2 16 9 9 9 13 0 2
17 3 7 13 15 9 9 9 2 13 15 0 9 3 3 13 9 2
5 9 13 0 9 2
25 9 13 9 0 9 16 3 15 13 9 13 2 15 13 3 13 3 15 13 2 7 3 15 13 2
14 7 16 9 13 9 9 2 9 9 9 13 0 13 2
6 0 9 2 0 9 2
10 9 9 0 9 13 0 2 3 0 2
14 13 0 13 9 2 13 0 9 2 13 9 1 9 2
34 16 15 13 9 9 9 2 9 13 3 13 2 16 9 3 13 9 2 16 9 2 9 9 7 9 9 1 9 13 9 13 9 0 2
25 9 13 3 15 16 0 9 2 15 13 0 9 2 0 9 7 9 2 15 13 3 0 0 13 2
24 15 13 2 16 9 13 3 16 13 9 15 15 13 9 13 2 13 3 4 13 15 9 9 2
18 9 9 9 4 3 13 9 0 9 2 7 15 4 3 13 3 13 2
21 9 2 16 9 9 13 0 13 9 0 9 7 13 9 9 9 2 13 0 9 2
10 9 9 9 3 13 12 9 0 9 2
5 0 9 3 13 2
22 9 13 0 2 16 0 12 9 9 13 13 2 13 13 9 9 2 9 7 9 9 2
7 3 2 9 13 0 9 2
38 4 3 13 9 2 13 3 13 13 9 0 0 2 7 13 13 0 9 13 9 2 15 9 13 13 0 9 7 9 2 7 15 13 13 3 0 9 2
18 9 13 3 9 2 13 15 3 9 2 16 9 0 9 13 13 9 2
15 13 13 2 3 3 15 13 9 9 13 3 9 7 9 2
12 13 15 2 16 9 13 13 0 2 13 0 2
17 13 9 13 15 15 9 2 15 9 13 3 0 2 13 9 3 2
14 13 2 16 0 9 4 13 0 16 0 7 0 9 2
14 15 3 13 13 13 0 9 2 0 9 7 0 9 2
15 7 0 9 9 9 9 2 3 3 3 4 15 9 13 2
7 15 13 3 13 9 13 2
11 0 2 0 9 1 9 13 3 3 0 2
6 9 3 13 13 9 2
13 9 9 13 9 4 3 3 13 13 0 9 9 2
5 3 3 13 9 2
15 0 9 3 13 9 1 3 3 3 13 9 16 0 9 2
12 9 13 9 13 9 9 2 16 9 13 9 2
12 3 3 16 9 13 9 2 9 9 13 3 2
11 3 9 13 9 2 7 0 9 15 13 2
11 0 3 9 9 4 3 13 3 0 9 2
14 0 9 2 9 7 9 9 4 13 9 2 3 9 2
18 15 13 9 7 9 13 9 7 9 0 9 2 13 3 13 9 9 2
10 9 9 3 13 9 7 13 0 9 2
13 3 9 7 9 13 9 4 3 13 9 3 9 2
16 2 13 13 2 13 0 9 2 13 9 9 15 13 3 0 2
15 3 4 3 13 3 13 13 9 15 2 16 9 13 0 2
6 3 3 11 9 9 2
4 12 9 9 2
7 9 13 9 3 0 9 2
8 12 9 13 3 12 9 9 2
12 9 11 9 13 13 9 9 3 3 12 9 2
11 9 13 2 7 15 9 9 13 9 9 2
8 3 0 2 15 13 13 9 2
19 9 13 13 3 3 0 2 7 15 13 9 0 3 3 3 9 9 1 2
23 9 13 3 15 2 13 15 13 13 3 0 0 9 15 2 15 15 12 9 9 9 13 2
11 15 13 2 3 9 0 9 4 9 13 2
11 7 3 3 3 0 9 15 4 9 13 2
20 9 0 9 7 9 9 4 13 3 0 2 7 9 9 4 13 3 0 9 2
4 13 3 9 2
16 0 15 9 9 0 9 9 2 12 9 9 2 12 9 9 2
5 9 2 12 9 2
12 0 0 9 13 9 2 12 9 9 7 9 2
6 9 2 3 12 9 2
30 0 9 13 9 2 9 13 9 9 2 3 3 12 9 2 7 9 9 13 12 9 0 9 2 15 13 9 7 9 2
17 15 9 4 13 15 9 9 0 9 2 15 15 9 13 7 13 2
6 9 2 3 12 9 2
29 13 3 0 9 9 2 3 3 9 13 3 3 0 2 7 15 9 15 12 0 9 13 13 9 3 0 9 13 2
14 15 9 1 9 1 13 3 3 15 9 9 13 9 2
10 0 9 0 9 13 3 13 3 0 2
21 3 9 9 13 9 13 3 0 9 9 7 9 13 15 2 13 9 9 7 9 2
21 3 3 0 7 0 9 4 13 9 0 2 7 9 1 15 13 9 13 15 9 2
9 9 9 13 3 13 9 0 9 2
28 15 15 9 13 13 9 3 9 2 15 15 9 0 9 13 9 13 3 0 9 2 7 13 9 15 9 9 2
22 13 13 13 9 2 15 13 9 15 2 13 13 9 13 7 13 16 9 13 13 3 2
39 9 13 9 4 13 3 0 2 13 3 3 13 15 2 16 9 9 1 4 3 13 3 2 13 3 3 13 16 9 15 9 3 3 15 3 3 13 2 2
19 13 3 9 9 2 16 0 9 13 9 13 9 2 7 3 9 13 9 2
13 9 13 0 9 2 7 9 9 13 9 7 9 2
19 0 0 15 9 13 15 2 13 3 4 3 3 13 3 9 12 9 13 2
14 9 13 13 9 2 15 9 7 0 9 13 3 13 2
6 9 13 9 13 9 2
14 7 3 3 9 13 9 15 11 13 2 13 9 13 2
13 0 9 9 9 13 3 7 2 7 3 9 13 2
31 3 0 9 9 13 9 4 13 15 2 16 9 13 15 7 9 0 7 3 0 9 1 15 9 2 15 13 9 3 13 2
9 15 3 13 0 0 9 15 9 2
21 13 3 9 9 9 13 9 11 11 2 15 13 15 9 0 9 13 12 9 1 2
36 9 11 0 9 13 13 0 2 7 3 15 13 2 16 13 15 9 3 0 9 2 16 9 13 9 13 9 9 2 16 4 13 13 9 9 2
4 13 15 9 2
6 9 13 3 9 9 2
52 3 3 3 16 13 0 9 2 15 9 9 13 13 9 2 7 15 3 3 13 9 9 2 2 13 3 9 2 7 3 0 9 1 13 0 7 3 0 9 15 2 3 3 7 0 9 9 12 9 1 13 2
2 9 9
16 9 13 3 9 9 7 9 1 13 0 3 13 2 11 2 2
10 0 0 9 13 3 0 9 0 9 2
18 13 3 9 2 16 9 13 13 9 9 7 11 9 13 3 13 9 2
3 13 9 2
5 15 15 3 13 2
15 9 13 13 13 3 0 9 7 15 2 0 2 4 13 2
15 11 9 4 13 2 11 13 3 15 15 7 11 13 9 2
4 15 3 9 2
9 3 13 15 9 1 15 9 1 2
23 9 13 0 9 11 2 11 11 11 11 11 11 11 11 2 13 13 3 15 13 13 2 2
12 11 13 0 2 3 7 3 0 0 9 9 2
11 9 13 12 0 9 2 15 13 0 9 2
10 11 0 0 9 13 13 9 1 11 2
14 3 4 9 9 13 12 12 9 7 15 11 13 9 2
13 9 9 13 13 0 9 12 9 3 13 0 9 2
5 9 13 9 9 2
8 15 13 3 9 9 11 11 2
9 7 13 13 0 13 9 9 11 2
15 3 11 11 11 11 9 2 15 13 12 9 13 1 11 2
10 15 15 13 0 16 13 9 0 9 2
12 2 13 0 2 7 13 15 13 3 0 2 2
3 13 3 2
18 9 13 3 12 5 7 15 13 9 2 9 9 7 12 9 15 9 2
5 9 13 3 3 2
14 13 4 15 3 2 15 13 9 7 9 13 9 9 2
10 9 13 1 11 2 9 13 3 9 2
24 13 2 16 13 9 9 1 13 3 0 12 9 3 3 2 16 15 13 3 9 2 13 9 2
15 9 11 9 13 9 9 2 7 0 9 13 9 13 12 2
9 3 13 13 3 3 9 13 13 2
9 11 2 11 2 11 7 3 11 2
15 13 3 3 9 11 9 2 5 2 7 13 13 0 9 2
6 11 13 9 0 9 2
9 4 15 3 13 9 13 13 9 2
4 0 9 9 2
5 7 13 3 9 2
9 13 13 2 3 9 13 11 9 2
16 11 13 9 2 15 13 13 9 0 2 16 15 4 13 9 2
14 15 13 9 9 9 2 7 13 0 9 9 13 9 2
12 9 13 13 9 9 13 9 13 9 9 9 2
7 0 9 13 3 0 9 2
16 3 9 13 0 9 1 2 7 13 15 3 13 9 7 9 2
17 9 9 1 11 4 13 9 2 15 4 13 9 9 1 13 9 2
13 3 3 9 13 3 3 2 3 12 9 13 15 2
17 7 3 16 9 9 13 0 0 9 2 13 11 13 9 9 9 2
15 11 9 13 9 2 15 13 13 9 9 7 15 9 13 2
9 3 3 2 13 9 13 9 1 2
19 16 9 13 13 0 3 2 13 9 13 13 13 15 9 7 0 9 1 2
9 11 9 4 13 9 3 13 11 2
15 3 9 13 13 2 13 9 3 9 7 13 15 3 11 2
2 9 9
4 9 13 0 2
6 3 13 2 15 13 2
12 3 13 13 9 9 2 12 9 2 3 3 2
5 9 13 12 9 2
12 9 4 13 15 9 2 15 13 15 0 9 2
14 9 13 13 15 9 0 9 2 7 15 13 9 1 2
9 15 13 3 13 13 0 9 9 2
17 3 15 13 13 13 15 2 7 3 9 13 13 3 0 7 0 2
24 15 4 13 3 15 2 16 15 15 13 13 9 2 3 15 9 13 13 15 9 16 0 9 2
14 13 3 12 0 9 2 15 9 13 16 9 13 9 2
10 9 13 2 16 13 13 3 0 9 2
8 3 9 3 13 1 0 9 2
20 13 0 13 0 9 2 13 13 9 0 9 7 13 2 16 9 13 0 9 2
11 9 13 3 0 9 2 15 3 13 13 2
17 0 9 13 3 3 0 0 9 7 9 2 15 13 3 0 9 2
9 2 6 2 3 15 13 0 2 2
14 15 1 13 9 0 9 2 9 13 9 3 0 9 2
20 13 3 13 2 16 13 13 0 0 2 13 2 9 2 9 2 9 9 13 2
18 13 15 3 0 2 16 4 0 9 13 15 9 2 13 13 3 0 2
22 9 3 9 9 13 13 9 13 9 9 9 2 16 9 13 13 13 15 13 9 1 2
14 9 9 7 9 13 15 9 13 2 7 15 13 9 2
5 3 3 13 9 2
23 15 4 13 9 9 2 3 9 13 3 0 9 13 9 2 7 3 9 13 0 9 9 2
7 3 13 9 0 9 9 2
11 9 13 3 3 9 7 9 9 13 9 2
12 9 13 3 0 2 0 7 3 9 13 9 2
17 15 13 9 15 9 2 16 3 13 13 9 9 15 9 13 9 2
21 3 13 15 3 0 9 2 16 15 13 13 15 9 7 13 13 0 16 15 9 2
17 9 13 9 2 15 9 9 13 9 4 13 9 2 7 3 15 2
8 9 9 9 9 13 0 0 2
11 9 1 15 13 2 0 9 13 2 9 2
20 15 9 13 9 7 9 0 9 2 7 9 13 3 13 0 13 13 0 9 2
10 15 9 3 13 3 12 5 0 9 2
13 9 13 9 2 15 12 9 13 13 12 15 13 2
13 3 9 13 9 2 15 4 13 2 9 3 2 2
13 13 0 13 15 9 3 15 9 7 9 1 9 2
10 13 3 13 2 15 9 13 12 9 2
5 13 3 13 13 2
13 0 9 9 13 3 12 2 12 2 12 7 12 2
8 11 13 0 9 7 11 9 2
31 9 9 13 9 2 15 13 3 9 9 13 9 2 2 9 11 11 2 13 0 9 2 7 2 11 11 2 13 0 9 2
15 9 13 3 3 0 9 2 15 13 9 3 9 13 9 2
8 0 9 9 13 9 4 13 2
11 9 13 12 9 2 16 9 13 9 9 2
6 11 13 9 1 9 2
11 11 2 15 3 13 0 9 2 13 9 2
2 9 9
14 2 9 13 2 16 3 15 13 13 15 13 11 11 2
4 3 11 13 2
9 9 13 7 13 2 2 0 2 2
13 2 9 13 9 2 15 1 9 13 0 13 0 2
14 11 13 15 3 9 2 2 13 15 13 15 9 2 2
11 3 13 9 13 7 13 2 2 13 2 2
18 3 11 13 13 2 16 0 3 13 9 4 13 11 9 9 9 3 2
12 15 13 0 9 7 9 9 7 0 9 9 2
12 2 9 13 7 13 3 2 2 15 13 9 2
7 6 15 13 15 9 2 2
15 2 15 9 13 2 16 9 4 15 13 9 2 9 2 2
5 9 13 15 9 2
15 3 11 13 2 2 7 15 4 13 9 13 9 11 2 2
8 0 9 13 2 7 11 13 2
6 11 11 11 11 11 12
7 15 9 11 13 9 11 2
10 13 9 13 9 2 0 9 7 9 2
20 0 9 13 9 9 0 9 2 12 9 13 9 11 9 7 13 9 0 9 2
15 9 0 9 7 0 9 13 9 15 11 2 15 13 9 2
11 9 13 9 12 2 15 13 9 9 9 2
19 0 9 13 3 3 9 2 7 13 13 15 2 15 9 13 13 3 9 2
12 3 9 0 9 13 15 11 9 0 9 9 2
9 9 9 13 9 2 7 15 13 2
17 11 9 13 0 9 3 0 9 9 2 15 13 0 9 13 9 2
9 9 13 9 13 0 9 7 9 2
8 15 1 11 13 0 9 9 2
15 9 9 13 15 0 9 0 9 2 13 11 9 13 13 2
16 9 13 12 9 4 13 9 9 2 13 3 0 9 13 9 2
19 11 9 4 3 13 15 9 9 9 0 2 15 15 13 0 9 11 11 2
13 15 13 9 9 7 9 3 3 12 9 13 9 2
14 9 1 9 13 9 2 15 9 9 13 9 9 9 2
7 3 9 9 13 9 9 2
18 11 0 9 13 9 9 9 7 13 9 13 15 2 13 13 0 9 2
17 13 9 0 2 8 8 8 8 8 2 9 7 9 9 0 9 2
13 0 9 13 9 2 3 13 0 9 0 9 13 2
18 9 9 13 9 2 0 9 2 9 2 9 2 9 7 11 9 9 2
14 15 9 13 0 9 9 2 7 9 4 13 3 9 2
16 3 9 13 11 13 9 9 2 7 4 13 13 3 9 9 2
6 0 9 13 0 9 2
19 15 9 9 9 4 13 9 9 7 9 9 2 13 15 13 9 3 9 2
10 9 3 13 9 9 9 2 3 3 2
16 9 13 13 3 7 0 2 15 13 9 15 0 9 9 13 2
16 15 9 9 1 4 13 9 9 13 9 2 15 9 3 13 2
16 11 9 13 0 9 7 13 3 3 2 9 13 13 9 3 2
16 9 13 9 13 2 16 9 9 13 3 3 16 11 13 3 2
25 9 13 0 9 13 3 0 0 9 13 2 16 15 9 9 13 13 9 3 3 2 3 1 9 2
23 9 2 15 9 9 13 9 9 2 9 9 2 13 2 16 9 9 13 3 9 7 9 2
11 9 13 3 12 12 9 7 15 13 9 2
14 9 9 13 3 13 9 2 15 13 9 9 15 13 2
13 0 9 13 11 1 9 13 16 13 11 13 9 2
14 9 13 9 13 9 7 13 9 9 9 0 9 9 2
14 0 9 13 13 11 9 9 2 15 13 0 9 9 2
9 9 9 9 9 1 13 0 9 2
7 9 13 13 3 0 9 2
10 9 1 3 12 9 3 13 9 9 2
14 0 9 9 13 9 9 9 13 9 9 7 9 13 2
20 9 13 9 9 13 13 9 9 1 2 16 3 15 13 13 9 9 1 9 2
15 9 13 13 3 9 0 9 2 16 15 9 13 9 9 2
7 9 13 13 0 9 1 2
12 9 9 13 13 9 9 7 15 13 9 9 2
17 9 13 13 9 2 7 13 13 9 9 9 2 3 1 9 9 2
18 9 9 13 3 0 2 3 3 0 2 16 9 13 15 3 0 9 2
18 9 13 9 9 3 2 13 0 9 1 13 9 2 7 13 9 3 2
12 0 9 13 3 9 7 13 9 0 9 13 2
7 9 9 1 9 13 3 2
14 9 13 2 9 13 2 9 13 0 7 9 13 13 2
15 9 1 9 3 13 9 13 3 7 13 9 0 0 9 2
13 9 13 3 9 2 16 11 11 13 13 9 9 2
8 9 13 9 13 9 15 3 2
31 0 9 13 3 15 9 2 15 13 0 9 9 2 12 0 9 7 9 1 11 11 11 13 9 13 11 1 9 0 9 2
16 9 13 2 16 9 13 9 13 0 7 13 9 7 11 9 2
21 0 9 13 9 13 11 11 13 0 9 2 15 3 13 11 9 7 11 0 9 2
17 9 13 0 2 16 9 13 3 7 9 13 11 9 4 13 9 2
12 3 11 9 13 9 13 2 3 0 0 9 2
21 15 9 1 9 13 0 9 7 13 1 9 13 2 9 13 0 9 11 2 9 2
16 9 1 11 9 9 13 9 9 13 13 9 13 0 9 9 2
10 9 13 3 13 3 15 0 9 9 2
7 9 4 13 11 9 1 2
10 9 9 13 9 7 11 9 9 9 2
2 9 9
6 9 2 0 2 9 9
13 11 9 0 9 13 3 9 8 2 2 9 2 2
15 9 13 0 9 2 15 9 13 3 0 9 7 13 9 2
21 15 9 9 13 3 0 9 2 3 9 9 0 9 2 0 9 9 7 3 3 2
26 9 13 2 3 9 13 3 0 9 7 13 15 9 2 0 13 9 13 7 3 15 13 13 7 13 2
7 9 13 9 13 3 9 2
11 9 4 3 13 15 9 7 9 9 9 2
8 15 9 13 9 13 9 11 2
20 9 13 3 13 9 0 9 15 9 2 16 3 0 0 9 13 9 4 13 2
21 9 13 3 15 9 2 15 13 3 15 9 9 2 15 13 13 3 9 9 1 2
21 9 7 9 4 3 13 9 9 9 2 15 4 3 13 0 9 9 9 7 9 2
14 0 9 4 13 0 0 13 9 2 15 13 1 9 2
7 15 9 13 13 0 9 2
24 3 11 9 9 13 0 2 3 13 9 2 9 2 15 13 0 2 0 7 0 9 7 9 2
17 3 3 13 9 2 0 9 2 15 13 3 0 9 2 9 9 2
18 15 12 1 13 0 9 2 9 9 2 15 13 9 7 9 0 9 2
12 1 15 0 13 9 15 13 4 3 3 13 2
9 9 13 1 9 2 15 0 9 2
21 3 9 13 13 9 2 16 9 13 0 9 7 9 2 3 13 3 3 0 9 2
18 9 9 9 9 13 9 13 9 9 1 13 0 9 13 9 9 9 2
13 13 3 13 9 2 13 9 9 13 0 9 9 2
10 9 7 9 13 3 13 0 0 9 2
17 9 13 13 3 0 2 3 15 4 13 2 16 9 13 9 13 2
21 9 13 3 0 2 7 15 4 13 3 0 9 2 15 13 13 0 15 13 13 2
12 3 9 4 3 13 0 9 2 3 11 9 2
16 11 9 13 0 9 2 15 13 0 11 9 2 3 9 9 2
7 9 3 13 13 0 9 2
25 0 13 9 9 2 15 1 13 13 0 9 2 15 13 0 9 2 15 9 9 13 9 0 9 2
7 15 1 9 13 3 13 2
8 13 3 13 9 9 2 9 2
14 9 13 0 9 2 15 15 13 9 7 15 15 13 2
13 9 13 3 9 9 2 13 9 9 4 9 13 2
12 3 9 13 3 9 2 9 15 0 9 13 2
4 9 9 7 9
14 9 7 9 4 13 3 2 16 13 9 7 13 9 2
20 16 13 11 9 2 9 2 13 4 13 9 13 3 2 6 2 13 3 15 2
20 13 3 4 13 15 9 2 16 9 2 9 2 9 2 9 2 13 13 9 2
5 3 15 3 13 2
17 3 15 9 13 2 0 7 13 4 13 0 13 9 2 9 9 2
12 13 3 2 15 3 13 9 1 2 15 9 2
7 9 15 9 13 3 0 2
18 9 13 3 13 9 13 9 2 3 15 1 4 3 13 7 9 13 2
24 16 9 13 3 3 2 9 2 9 2 9 7 9 13 15 0 9 2 4 9 13 15 9 2
13 16 9 13 13 13 9 0 2 15 13 9 9 2
7 3 9 13 13 9 9 2
18 16 9 13 13 3 3 2 15 13 9 3 3 7 13 9 9 9 2
23 13 9 7 9 13 9 13 3 13 9 2 13 15 0 2 16 3 0 2 9 9 9 2
14 9 13 0 0 9 2 3 9 0 9 15 9 9 2
27 15 13 3 9 7 3 9 9 2 15 13 9 9 9 2 9 7 9 9 0 9 9 2 7 3 9 2
8 15 9 9 13 3 9 1 2
33 3 11 11 11 0 9 4 13 9 15 2 3 0 9 9 13 0 9 2 15 9 9 3 13 0 9 7 13 0 9 1 0 2
7 13 9 9 7 9 9 2
13 9 13 9 0 9 2 7 15 13 9 15 1 2
11 16 9 13 13 9 9 2 13 0 9 2
22 9 13 9 9 2 15 15 9 13 13 15 2 16 15 3 13 0 7 0 9 1 2
4 3 9 13 2
23 3 11 9 0 9 0 13 9 2 15 9 9 13 9 13 3 9 7 3 3 9 9 2
9 3 15 4 13 3 9 2 9 2
20 9 9 13 9 9 2 9 13 3 9 9 13 9 2 15 15 9 13 15 2
10 16 9 4 13 9 2 15 13 9 2
18 15 0 4 3 13 2 9 4 13 0 2 15 4 13 0 9 15 2
47 15 4 13 3 7 3 2 9 13 4 13 3 9 2 7 0 9 4 3 13 9 2 15 13 15 0 9 9 13 2 15 13 9 7 9 13 0 9 2 15 9 13 9 4 13 0 2
20 16 9 4 13 9 9 2 4 0 9 3 13 15 9 2 3 0 0 9 2
19 0 9 9 13 3 13 0 9 9 3 2 9 2 9 7 9 2 1 2
10 9 13 3 13 3 0 13 9 9 2
11 7 15 15 9 13 16 9 0 9 9 2
3 9 9 2
20 0 9 9 7 9 13 13 9 15 2 7 9 13 3 9 15 12 9 1 2
8 15 4 13 9 0 0 9 2
11 16 9 13 13 13 2 0 9 4 13 2
22 0 9 13 0 9 13 3 13 2 7 9 15 13 9 0 9 7 9 9 7 9 2
7 9 3 13 13 0 9 2
14 15 13 9 2 0 9 7 9 2 15 1 13 9 2
25 15 9 2 9 2 3 0 9 7 9 9 13 9 4 13 15 9 2 15 13 9 0 13 9 2
16 9 13 13 3 9 2 9 2 15 9 13 15 9 13 3 2
6 9 13 2 15 13 2
1 9
3 0 9 9
12 9 9 13 9 9 9 13 13 2 15 13 2
5 13 3 13 3 2
17 3 13 9 7 9 2 3 9 4 3 13 9 7 13 9 9 2
13 9 13 3 15 0 2 16 9 13 13 9 13 2
25 15 9 3 9 13 15 2 16 0 9 13 13 13 3 0 13 9 2 7 15 4 13 13 9 2
9 13 9 13 2 9 13 13 0 2
8 3 4 15 9 13 0 9 2
16 7 3 15 9 9 13 0 3 13 2 7 9 0 9 13 2
11 3 15 9 13 0 9 7 9 13 13 2
5 9 9 7 13 2
15 9 1 13 3 0 9 2 16 13 13 9 9 0 9 2
18 9 7 9 13 3 2 13 3 0 9 9 9 2 3 0 9 13 2
14 9 4 13 2 16 9 13 9 13 13 1 15 9 2
10 9 13 9 9 13 0 9 13 9 2
14 9 9 13 2 16 9 13 11 2 7 3 3 13 2
9 9 1 9 13 0 9 0 9 2
31 9 1 13 3 0 9 2 9 13 15 9 2 16 0 8 2 7 15 9 2 16 9 1 13 9 7 3 13 0 9 2
7 7 3 2 11 15 3 2
15 3 7 3 13 3 3 9 7 12 7 15 3 13 9 2
11 9 13 13 2 15 9 13 3 3 13 2
10 15 9 9 3 9 13 13 1 9 2
21 9 13 11 9 7 9 1 13 15 9 3 0 0 0 9 9 9 2 3 9 2
6 7 15 9 3 13 2
5 7 3 13 3 2
10 0 0 9 13 11 7 11 9 13 2
13 3 16 11 0 11 11 9 9 13 13 1 15 2
9 3 13 15 0 2 3 13 9 2
26 3 3 9 13 3 0 2 16 3 0 9 13 2 0 2 3 13 9 2 16 15 13 3 0 9 2
30 13 15 2 16 3 9 11 7 11 2 11 2 13 0 0 9 9 2 0 9 2 2 7 15 9 13 15 13 0 2
16 3 15 9 9 13 15 9 9 3 0 2 15 13 13 9 2
9 3 9 13 3 9 9 9 1 2
15 9 3 13 9 1 13 9 2 7 0 9 13 3 0 2
21 9 9 13 3 3 0 13 9 0 9 13 9 7 4 13 0 9 9 3 9 2
8 9 13 3 0 16 13 13 2
16 3 9 9 15 9 13 13 0 2 13 9 7 9 13 9 2
6 9 13 9 7 9 2
11 9 9 13 2 3 2 12 5 9 1 2
11 3 0 9 13 2 13 9 9 3 0 2
12 3 15 3 2 16 13 15 0 9 9 1 2
22 9 13 3 13 7 3 3 13 9 9 9 0 9 9 2 9 13 13 3 3 0 2
24 9 15 9 4 13 9 7 9 2 13 13 13 9 15 9 9 9 2 7 3 13 9 3 2
17 9 13 3 9 13 3 12 0 9 3 2 3 9 13 9 3 2
9 9 4 3 13 3 0 9 9 2
8 3 4 13 9 15 3 9 2
12 9 13 3 0 9 2 16 13 15 9 1 2
12 13 2 16 9 13 3 0 9 15 0 9 2
15 16 9 4 13 9 0 9 2 15 13 3 13 0 9 2
8 13 3 9 3 0 0 9 2
18 7 3 15 2 15 13 3 13 2 15 13 9 2 4 13 0 9 2
4 9 13 2 9
6 9 13 9 0 9 2
32 15 13 2 13 2 13 2 13 2 13 2 13 2 13 2 13 2 13 7 13 2 4 15 9 9 13 9 9 13 9 9 2
20 15 9 0 9 13 11 0 9 7 13 2 15 9 7 0 9 13 9 13 2
10 9 13 12 0 9 0 9 9 13 2
9 15 9 13 9 13 13 7 13 2
15 9 9 13 3 7 3 7 3 0 9 13 15 9 9 2
16 3 0 9 0 9 13 11 9 2 15 9 13 13 15 9 2
12 15 9 9 13 7 0 2 0 7 3 0 2
2 11 9
3 9 2 11
8 9 2 11 11 2 9 12 2
11 0 9 1 13 3 0 9 9 13 9 2
10 0 9 13 0 9 13 0 0 9 2
16 3 13 0 9 13 9 7 9 13 11 13 9 9 9 9 2
8 11 9 9 13 4 16 13 2
18 9 13 9 3 3 2 9 7 9 1 9 13 3 9 7 0 9 2
12 9 13 0 0 7 9 3 1 0 9 9 2
10 3 9 13 0 9 13 0 9 9 2
9 9 9 13 9 9 9 9 0 2
11 9 13 0 2 0 0 7 0 9 13 2
13 3 9 13 3 2 13 0 9 9 13 3 0 2
20 9 1 13 9 13 9 9 2 13 9 9 7 13 0 9 9 9 15 9 2
9 9 13 0 0 7 3 0 9 2
14 9 9 13 3 9 2 15 3 4 3 13 9 1 2
12 9 13 0 7 9 15 9 1 13 9 1 2
12 9 13 3 9 0 9 9 7 15 0 9 2
12 15 9 13 9 9 2 3 9 13 0 13 2
7 9 9 13 3 1 0 2
14 15 1 9 13 9 1 0 13 13 0 9 0 9 2
9 13 2 9 2 9 2 9 2 9
9 13 2 9 9 7 9 13 9 9
3 9 2 12
16 9 2 2 3 13 12 9 2 16 15 9 13 0 9 2 2
1 0
3 9 2 9
11 9 2 0 13 9 2 0 0 9 9 2
18 11 11 1 13 9 13 9 0 9 1 0 9 9 0 0 7 0 2
8 9 9 13 3 11 9 0 2
18 3 9 13 13 13 13 7 9 9 13 9 2 3 0 9 13 13 2
4 13 2 0 9
4 13 2 0 9
3 9 2 9
5 9 2 13 15 0
1 0
5 9 2 9 9 12
11 9 2 11 11 2 9 0 7 0 9 2
9 9 9 12 13 9 13 9 9 2
20 15 0 9 13 13 0 9 9 2 7 9 1 9 13 13 0 3 0 9 2
8 9 9 13 9 13 0 9 2
16 9 9 13 0 7 3 9 9 1 15 13 9 0 0 9 2
16 9 13 2 7 15 4 13 3 9 2 15 9 13 13 0 2
11 9 13 0 0 7 9 9 13 0 9 2
18 9 9 0 9 13 3 13 0 2 16 0 9 9 13 1 9 9 2
6 3 0 9 13 13 2
8 9 9 13 3 9 0 9 2
13 9 9 13 0 0 2 7 9 7 9 13 13 2
22 0 9 13 3 9 9 2 15 13 15 15 9 13 9 3 13 9 9 0 9 13 2
9 9 13 3 0 13 3 0 9 2
12 9 13 9 2 0 9 7 3 0 9 9 2
15 9 13 9 9 3 9 2 16 9 9 15 4 13 13 2
16 9 13 9 7 9 7 9 2 3 9 9 13 0 7 0 2
15 9 13 3 15 9 11 9 1 2 15 13 0 9 9 2
14 9 13 3 9 7 15 0 9 9 13 13 15 9 2
7 13 2 9 2 9 7 9
8 13 2 3 0 9 7 0 9
3 9 2 12
6 9 2 2 9 2 2
1 0
5 9 2 9 9 12
9 9 2 11 11 9 2 9 9 2
8 9 1 13 9 4 9 13 2
11 9 13 9 9 9 7 3 13 0 0 2
16 9 13 9 9 13 9 7 13 0 2 16 3 13 13 9 2
9 3 9 13 0 9 9 0 9 2
5 0 9 13 3 9
12 9 9 9 9 13 0 7 9 13 9 0 2
4 13 3 3 2
9 13 2 3 3 9 9 13 9 2
3 9 9 2
3 9 13 2
9 15 9 4 13 0 9 9 3 2
14 9 4 13 0 2 16 9 9 4 13 3 3 0 2
27 3 9 0 9 1 13 0 0 2 9 11 9 13 9 13 2 16 9 9 9 4 13 9 9 3 3 2
17 9 9 13 9 4 13 9 0 12 9 3 16 0 9 0 9 2
14 9 3 0 9 7 9 11 4 13 9 3 12 9 2
5 9 13 2 3 9
20 9 9 1 0 9 7 9 9 13 9 0 9 9 9 13 12 9 0 9 2
6 9 9 13 12 9 2
10 9 9 4 13 3 0 9 15 0 2
6 15 9 13 3 9 2
16 15 9 9 9 9 13 3 3 2 11 9 9 11 11 13 2
22 2 9 9 4 13 3 2 7 16 9 3 13 2 13 9 2 13 9 3 0 9 2
26 0 9 2 13 3 2 13 2 16 12 9 0 9 11 13 4 13 3 3 12 12 9 9 9 9 2
14 0 9 13 0 9 0 9 3 12 12 9 0 9 2
22 9 12 9 9 9 9 11 13 3 12 9 0 16 0 9 0 9 2 3 12 9 2
26 2 16 13 2 16 9 9 1 13 3 9 2 15 9 13 13 2 3 9 13 13 9 2 11 13 2
10 9 9 4 13 13 0 9 9 11 2
10 9 0 9 9 9 13 12 9 9 2
9 3 12 9 9 9 13 12 9 2
7 3 9 9 13 15 0 2
19 0 9 9 13 0 9 0 9 12 9 9 0 9 7 12 9 9 9 2
5 13 9 9 9 2
11 9 9 0 9 9 13 12 9 9 9 2
12 9 9 3 13 11 0 9 9 9 0 9 2
22 9 11 11 13 2 16 9 13 3 3 9 15 2 3 15 13 3 9 9 9 9 2
10 3 2 13 0 9 9 0 9 0 2
13 3 3 13 9 12 9 9 13 3 12 12 9 2
23 11 13 2 16 9 9 13 3 0 2 7 7 9 9 7 9 9 13 3 3 16 3 2
11 0 9 9 13 9 12 9 9 12 9 2
8 9 13 2 15 9 9 13 2
13 3 4 13 9 2 9 7 9 7 9 9 13 2
7 9 9 4 13 13 9 2
12 15 4 13 0 9 9 0 9 13 9 9 2
16 11 9 13 0 9 2 16 13 9 13 9 9 9 0 9 2
11 15 3 4 13 9 3 0 11 9 9 2
21 2 9 13 3 2 13 15 0 9 13 9 2 13 13 0 11 9 2 11 13 2
4 9 9 0 9
10 9 4 13 0 9 1 0 9 9 2
13 9 13 3 15 9 2 7 11 2 11 7 11 2
11 9 13 3 13 0 9 12 9 13 9 2
14 0 9 9 13 2 16 9 9 13 15 15 16 0 2
11 11 9 13 9 13 9 9 9 0 9 2
13 9 13 2 16 11 9 11 13 13 9 9 12 2
10 9 4 13 9 9 13 9 9 12 2
7 9 9 13 0 12 9 2
9 3 12 9 9 13 3 9 9 2
28 2 9 0 9 13 15 3 3 13 9 1 0 2 16 9 9 13 15 16 3 0 9 13 2 11 13 9 2
8 3 0 13 9 11 7 11 2
11 9 9 13 9 12 7 0 3 9 12 2
14 11 7 11 9 13 9 12 1 9 9 4 13 11 2
20 3 15 9 13 13 3 0 2 9 9 13 9 13 9 0 9 3 9 12 2
3 9 9 13
16 9 11 1 9 0 9 13 9 2 9 2 7 0 0 9 2
25 2 9 13 9 15 2 16 9 9 13 7 3 7 0 9 2 9 11 11 9 11 11 13 9 2
17 11 9 9 13 3 0 16 9 2 9 4 13 3 3 12 9 2
25 11 1 2 0 0 3 13 9 13 3 13 0 9 3 9 0 9 2 15 13 9 9 13 2 2
12 2 11 4 13 15 15 16 3 0 0 9 2
9 9 9 4 13 7 0 9 13 2
14 15 13 0 0 9 2 11 9 11 11 13 9 11 2
5 9 9 2 13 2
7 11 9 13 9 1 9 2
20 9 9 13 9 2 16 9 3 0 0 9 13 9 9 0 3 3 12 9 2
16 0 9 9 9 13 12 9 2 16 9 4 13 12 9 9 2
10 9 13 0 0 9 12 9 12 9 2
17 9 13 2 13 2 2 11 11 11 9 11 11 13 11 9 9 2
11 9 13 3 9 9 13 9 0 9 11 2
3 9 13 9
14 11 9 9 13 9 9 9 2 13 9 9 9 13 2
10 9 11 11 13 15 9 2 9 2 2
7 9 13 9 7 13 9 2
22 11 13 9 1 9 13 0 9 4 13 9 9 2 15 9 0 9 13 9 9 3 2
10 2 3 13 2 0 9 9 3 13 2
18 15 13 13 13 0 13 9 9 2 0 11 11 9 11 11 13 11 2
8 2 9 4 3 13 0 9 2
11 3 15 13 3 9 2 7 3 0 0 2
17 13 0 2 16 9 13 13 9 2 13 3 0 9 9 11 11 2
9 0 9 9 13 15 13 3 9 2
20 15 11 9 0 9 13 0 9 2 7 9 7 9 12 9 13 13 3 9 2
7 15 9 4 3 13 9 2
17 9 9 9 13 2 16 11 13 0 9 3 16 9 4 13 9 2
7 11 13 9 9 2 13 2
17 11 9 0 9 13 11 2 15 0 9 3 12 9 13 0 9 2
12 0 11 0 11 11 9 13 9 3 11 9 2
11 9 13 3 11 13 9 9 2 9 13 2
9 2 9 4 9 9 13 9 1 2
35 13 9 3 11 0 0 9 7 11 0 0 9 2 15 4 13 0 9 7 13 0 9 2 16 15 13 13 0 9 13 0 9 7 13 2
18 2 3 0 3 15 13 2 9 9 13 2 16 9 13 9 0 3 2
25 13 3 3 0 7 9 9 2 16 11 13 9 7 13 9 12 12 9 2 7 3 0 2 9 2
6 11 2 0 0 7 0
4 9 13 9 2
16 13 3 0 2 7 3 11 9 2 9 11 11 13 11 11 2
16 11 9 11 13 9 3 3 9 7 9 2 16 9 13 13 2
12 11 11 7 11 9 13 3 13 0 9 9 2
12 11 3 13 2 13 11 9 13 0 9 3 2
19 2 15 4 3 11 13 0 0 9 7 13 0 9 2 16 15 13 9 2
18 3 13 9 3 15 3 2 16 11 13 13 2 11 13 11 11 11 2
16 11 1 11 4 13 9 3 3 2 16 15 9 13 11 13 2
10 9 11 13 3 9 0 15 9 9 2
8 2 0 11 13 3 0 9 2
16 15 9 13 13 9 2 16 11 7 11 9 9 13 0 9 2
14 15 13 0 0 7 0 9 2 11 13 11 11 9 2
15 9 13 13 11 9 0 13 11 13 9 7 9 11 9 2
14 0 13 2 16 11 7 11 9 13 0 9 9 9 2
20 2 2 0 0 2 9 4 13 3 0 9 0 9 2 16 15 13 9 9 2
14 7 9 2 9 9 7 0 9 2 11 13 11 11 2
2 9 13
8 9 13 3 11 9 9 9 2
14 11 9 9 13 3 2 15 15 9 13 2 0 9 2
7 3 15 9 13 9 0 2
10 9 11 13 13 3 13 15 9 3 2
11 11 9 9 11 13 9 3 12 9 9 2
7 11 9 13 0 12 9 2
11 9 11 9 13 9 2 7 15 9 13 2
11 11 1 15 9 9 9 9 13 3 0 2
8 11 9 9 13 9 12 9 2
10 15 9 13 11 9 2 7 3 3 2
6 9 13 9 1 11 2
11 11 11 11 9 13 12 9 3 9 13 2
11 9 9 13 3 2 7 9 13 12 9 2
16 11 11 11 4 13 9 13 9 9 12 9 2 9 11 13 2
15 9 13 3 3 9 11 0 9 7 9 11 7 11 9 2
12 9 13 9 9 0 9 2 12 12 9 9 2
7 9 4 13 9 12 9 2
7 0 9 2 9 4 13 9
11 3 0 9 7 15 9 4 13 9 9 2
19 0 9 9 4 13 2 16 9 4 13 2 13 9 11 11 9 7 9 2
8 9 13 2 7 0 9 13 2
11 9 9 1 9 9 4 13 12 12 9 2
15 9 7 9 9 11 11 13 0 9 2 9 4 13 9 2
15 11 1 0 9 13 9 9 3 0 7 15 13 3 3 2
7 2 15 13 3 15 9 2
9 9 13 12 2 16 9 13 0 2
10 11 1 9 13 3 0 0 9 1 2
21 2 13 2 16 9 13 3 0 2 13 13 0 13 9 9 3 3 16 13 3 2
22 2 9 13 3 3 2 7 15 13 9 15 9 2 16 15 4 3 13 9 13 9 2
3 9 4 13
9 11 11 1 9 13 9 7 9 2
13 2 16 9 13 3 3 2 15 13 13 3 13 2
8 9 9 13 3 3 3 9 2
11 16 9 13 2 15 13 3 13 13 3 2
11 11 13 2 16 9 9 9 1 13 0 2
13 15 1 0 13 13 9 3 16 9 13 13 0 2
7 2 9 9 13 0 13 2
4 9 13 13 9
8 9 7 9 13 13 0 9 2
10 11 11 13 9 0 9 7 9 9 2
13 2 9 9 9 13 9 9 13 15 9 3 9 2
18 9 9 13 0 2 7 11 13 2 16 3 13 9 4 13 3 13 2
15 2 9 9 13 0 9 2 3 0 9 13 3 16 9 2
13 2 3 13 0 9 2 7 9 13 0 9 3 2
8 15 13 13 3 3 13 9 2
9 11 13 2 16 9 13 13 9 2
26 2 0 9 13 4 3 13 15 2 3 3 9 13 2 7 15 4 3 13 15 2 3 0 15 13 2
15 2 9 13 9 9 9 2 7 15 13 4 13 3 13 2
5 11 13 9 13 3
4 11 9 11 11
11 11 9 0 9 13 0 9 0 9 0 2
11 9 1 9 13 3 12 9 12 12 9 2
8 9 7 9 9 13 3 9 2
9 9 13 15 1 13 0 9 9 2
14 0 9 9 7 9 13 9 12 9 0 12 12 9 2
7 9 9 9 13 12 9 2
9 9 9 15 1 13 3 12 9 2
5 9 13 15 3 2
7 3 11 9 13 12 9 2
7 9 13 3 7 12 9 2
10 9 9 13 12 12 9 12 12 9 2
8 9 13 12 9 9 7 9 2
15 11 0 9 9 1 9 13 12 9 0 9 12 12 9 2
14 2 9 13 0 7 9 9 0 1 9 13 9 12 2
6 9 13 9 0 9 2
13 0 0 13 9 9 9 2 9 11 11 13 9 2
12 11 13 2 16 0 9 9 13 0 9 0 2
3 11 13 11
9 11 13 12 12 9 9 11 12 2
12 11 13 9 2 15 13 3 0 9 11 9 2
6 11 4 13 9 9 2
9 11 13 3 3 9 11 9 9 2
12 11 11 13 11 11 9 13 3 0 11 9 2
35 0 11 11 9 7 9 1 9 4 15 9 13 16 11 9 2 9 13 11 2 0 9 13 15 7 3 9 9 13 0 9 4 13 11 2
9 9 13 0 7 12 12 9 0 2
13 11 0 9 13 11 11 11 4 13 9 9 1 2
22 2 11 13 3 0 13 9 3 2 16 9 4 13 0 13 3 15 2 15 11 13 2
20 16 15 9 13 15 9 2 15 4 13 9 9 2 11 9 11 11 13 11 2
9 11 11 11 13 9 3 9 9 2
26 2 0 2 15 4 13 13 0 9 9 2 13 13 0 9 3 7 13 11 9 9 2 9 13 9 2
8 11 4 13 11 9 9 12 2
9 15 13 9 12 9 7 9 9 2
7 11 1 13 3 13 11 2
15 11 13 9 3 9 11 9 9 2 9 7 9 13 9 2
9 15 4 3 3 13 11 9 9 2
7 11 2 9 13 13 0 9
9 9 9 4 0 9 13 9 9 2
18 9 13 9 13 9 9 9 2 15 13 13 1 9 2 13 11 9 2
20 9 9 9 9 1 4 13 9 2 15 4 13 3 9 15 13 9 0 9 2
16 12 9 7 0 9 9 9 4 13 3 3 2 12 9 9 2
10 2 0 9 13 3 12 9 1 9 2
21 9 13 9 2 13 15 4 13 3 3 2 9 11 9 9 11 11 13 11 9 2
5 3 13 15 3 9
7 9 9 13 7 9 13 2
13 9 13 9 13 9 2 7 9 13 9 9 9 2
7 15 13 0 13 9 9 2
14 11 13 12 0 9 2 15 9 13 15 3 3 9 2
22 9 7 9 9 9 13 15 9 13 0 9 2 9 9 7 9 13 9 9 0 9 2
9 15 9 9 9 4 13 0 0 2
10 9 0 9 9 9 9 13 0 9 2
10 3 9 13 9 9 13 9 0 0 2
24 9 13 0 13 2 7 15 9 9 4 13 9 9 2 13 11 9 7 9 9 9 11 11 2
18 15 7 15 9 9 13 11 12 9 2 15 13 13 15 3 3 9 2
7 0 13 3 2 13 7 13
11 13 0 9 13 9 9 7 15 9 9 2
13 16 9 13 2 9 7 9 13 13 3 3 13 2
4 9 9 13 2
3 9 13 2
8 2 15 13 3 13 0 9 2
19 0 9 4 3 3 13 2 16 9 9 7 9 13 3 2 11 11 13 2
13 3 11 9 9 11 11 13 9 9 9 0 9 2
18 2 9 9 4 15 9 13 13 9 9 3 2 16 0 9 9 13 2
14 11 13 2 16 9 4 13 2 16 0 9 13 0 2
14 3 13 0 9 9 2 3 9 2 0 9 7 9 2
15 2 3 0 9 0 4 13 13 7 13 9 9 3 3 2
12 9 4 13 3 3 3 9 7 15 9 9 2
15 9 13 3 3 2 16 9 13 3 9 9 2 15 13 2
11 9 13 9 13 0 13 3 9 1 9 2
10 3 9 9 7 3 9 9 13 3 2
5 0 13 3 12 9
6 9 13 13 11 12 2
6 0 9 13 3 15 2
5 9 13 9 9 2
12 9 9 13 15 9 3 3 12 12 9 9 2
7 13 9 13 3 9 9 2
10 9 9 13 9 3 3 12 12 9 2
12 0 9 13 15 2 16 0 9 9 13 0 2
18 9 12 0 9 9 2 9 2 13 12 7 9 3 3 12 12 9 2
22 9 13 3 0 0 9 7 9 7 9 2 13 0 9 9 7 9 9 3 13 9 2
27 11 11 11 1 0 13 9 13 2 16 13 9 13 13 3 3 0 9 2 0 9 0 7 3 13 9 2
11 9 0 9 13 3 12 2 3 12 9 2
8 9 3 13 9 3 0 9 2
8 3 9 9 13 9 9 0 2
7 0 13 12 9 2 13 15
15 13 4 13 0 9 3 3 13 9 7 13 12 9 9 2
27 2 3 13 2 16 13 9 13 13 15 12 0 9 7 13 3 15 15 2 11 9 7 9 11 11 13 2
17 9 4 3 13 3 9 15 2 16 9 13 9 9 2 15 13 2
9 11 1 0 9 13 13 0 9 2
26 15 4 13 3 12 0 7 12 0 9 9 7 9 13 2 3 9 13 9 3 7 3 9 13 13 2
11 2 3 3 4 13 3 9 9 7 9 2
13 3 9 1 4 3 13 7 13 9 2 11 13 2
10 16 9 13 3 2 13 9 13 9 2
20 9 13 13 9 2 9 7 9 13 9 3 2 3 9 7 9 3 15 1 2
4 9 13 0 2
10 9 0 9 13 9 4 13 3 3 2
14 9 4 13 0 9 3 2 16 9 13 12 9 3 2
16 9 13 3 9 0 9 13 9 2 16 9 13 13 13 9 2
6 0 13 2 4 13 9
10 0 9 9 4 0 9 13 0 9 2
6 9 13 7 9 13 2
12 11 11 1 9 13 3 3 0 9 9 9 2
13 9 4 13 9 7 15 9 13 9 7 9 9 2
7 9 13 3 9 13 11 2
19 11 13 9 13 9 4 0 9 13 3 3 3 9 2 13 9 11 11 2
16 9 13 15 1 2 16 9 13 3 9 13 9 9 13 9 2
12 2 9 9 9 13 0 2 16 9 13 0 2
16 3 9 9 13 0 2 7 0 9 9 13 0 2 11 13 2
6 0 13 15 9 3 3
17 9 9 13 7 9 13 3 12 7 15 9 2 9 13 9 9 2
14 15 9 3 9 7 9 13 3 13 9 2 3 9 2
7 3 3 9 9 13 3 2
17 11 11 11 13 2 16 9 13 13 13 2 13 9 9 15 3 2
5 9 3 13 9 2
17 9 13 9 7 9 9 13 9 2 7 15 4 13 15 3 13 2
16 2 15 13 3 13 9 0 9 1 9 13 9 2 11 13 2
4 9 2 13 9
7 9 9 13 13 0 9 2
7 0 9 13 9 13 9 2
11 9 13 0 0 9 9 13 9 13 9 2
12 3 0 13 13 3 3 13 9 2 3 9 2
11 0 9 13 13 9 9 0 2 9 13 2
9 9 13 0 9 3 12 9 9 2
17 9 13 3 9 9 2 15 13 12 9 0 9 2 13 11 9 2
11 0 9 13 3 3 9 2 9 7 9 2
13 11 9 9 11 11 13 9 0 9 0 9 9 2
16 2 0 0 9 9 13 9 3 3 13 0 7 9 9 9 2
22 3 13 9 2 3 9 7 9 2 4 13 13 0 9 2 15 13 3 13 0 9 2
12 9 9 13 15 9 9 9 2 9 13 11 2
3 9 0 9
20 11 11 13 2 16 9 13 13 3 3 0 15 2 3 0 9 9 13 9 2
16 9 13 0 9 3 2 7 9 0 9 9 3 13 3 0 2
16 3 15 2 3 9 4 13 2 4 13 13 9 9 13 9 2
15 9 7 3 0 9 9 13 13 9 2 15 13 9 9 2
9 2 9 13 9 9 13 0 9 2
10 9 13 9 9 1 4 13 15 9 2
16 4 3 13 2 16 12 9 3 3 13 13 0 2 11 13 2
3 0 9 0
12 9 11 11 13 2 16 0 9 13 0 9 2
9 2 9 4 13 1 3 0 9 2
23 9 13 3 0 9 2 16 13 0 3 13 2 15 9 13 15 0 9 0 9 15 9 2
20 2 16 9 13 0 9 0 9 2 15 4 13 0 9 7 9 9 13 0 2
18 9 9 9 13 9 0 9 2 15 4 13 13 9 3 2 15 13 2
6 9 13 2 13 9 9
10 11 9 11 13 9 9 9 0 9 2
8 9 4 13 12 12 9 9 2
35 11 0 9 9 4 13 11 9 9 7 9 9 12 9 2 9 11 11 7 9 11 11 12 12 9 9 9 0 9 9 2 9 13 9 2
7 9 13 13 9 13 9 2
16 9 9 13 13 15 0 9 2 15 13 9 13 0 9 9 2
14 0 9 9 13 9 9 0 0 9 2 3 13 9 2
18 9 9 0 9 2 3 13 9 2 9 7 9 13 4 13 3 3 2
18 2 9 9 0 9 13 3 9 9 7 0 9 13 9 1 7 13 2
17 15 13 15 9 9 2 7 3 2 3 0 0 2 11 13 9 2
11 11 7 11 13 13 9 13 9 0 9 2
16 2 13 0 13 9 0 9 2 16 15 1 9 13 9 13 2
19 13 2 16 0 9 13 0 9 2 15 4 13 0 0 9 2 11 13 2
9 9 13 9 9 0 9 9 9 2
8 0 9 13 0 9 13 9 2
11 9 13 2 16 9 13 9 9 13 9 2
16 15 2 15 13 3 0 9 2 3 13 0 9 9 9 13 2
6 15 13 3 0 9 2
7 15 7 13 13 12 9 9
9 11 9 13 9 9 0 9 9 2
8 9 13 13 0 12 9 9 2
11 13 2 15 9 7 9 12 9 9 13 2
18 11 13 15 15 15 9 2 15 13 15 0 7 12 9 9 0 9 2
23 9 9 4 13 3 9 2 16 9 4 13 11 9 9 2 16 9 13 13 9 9 9 2
7 9 11 13 11 0 9 2
18 3 12 15 0 9 2 11 5 11 7 11 11 2 13 11 9 9 2
15 9 13 3 3 2 16 11 9 7 9 13 9 9 9 2
6 3 0 9 9 13 2
18 11 13 3 9 2 16 11 9 13 12 9 9 2 16 9 9 13 2
15 9 3 13 0 2 15 13 15 2 16 9 9 9 13 2
12 9 9 4 13 0 9 1 13 9 0 9 2
10 0 9 13 9 7 9 15 0 9 2
7 16 9 13 2 9 13 2
11 12 9 9 9 13 0 7 15 9 0 2
3 12 9 9
17 11 7 11 5 11 12 9 9 13 11 1 12 15 9 7 9 2
10 11 5 11 9 13 3 15 9 0 2
19 11 5 11 13 2 16 15 13 9 3 2 16 13 13 3 3 13 9 2
18 11 9 13 11 1 11 2 3 9 13 3 0 3 1 11 7 11 2
12 11 9 13 3 3 0 11 2 11 7 11 2
11 9 3 13 11 2 11 2 11 7 11 2
5 0 9 13 15 9
4 2 11 11 11
3 2 11 11
4 2 11 5 11
2 2 11
8 11 13 11 9 9 0 9 2
7 9 1 11 9 13 0 2
12 11 4 13 0 9 3 11 5 11 7 11 2
4 11 9 13 2
17 11 11 11 13 9 2 16 11 1 11 12 9 9 4 13 13 2
24 0 9 11 4 13 11 15 2 16 15 13 3 13 9 9 9 2 16 9 13 13 0 3 2
9 11 9 9 13 12 9 9 9 2
19 9 9 1 13 11 11 11 1 3 11 2 15 9 9 9 13 12 9 2
17 11 9 9 13 13 0 11 9 2 13 11 7 11 15 0 9 2
5 12 9 3 12 9
11 9 12 9 9 0 9 13 3 0 9 2
22 11 5 11 4 13 15 9 3 12 9 7 11 2 11 2 11 11 7 11 5 11 2
10 0 9 9 13 3 11 11 11 11 2
12 9 3 13 12 9 9 0 9 0 9 1 2
11 3 9 9 0 9 13 9 13 3 12 2
14 12 9 9 12 9 0 11 13 11 7 11 11 11 2
8 9 4 13 9 7 9 9 2
17 11 1 15 12 9 13 13 9 13 9 2 16 11 9 9 13 2
6 11 9 2 13 13 9
17 9 11 11 13 9 9 2 15 1 15 4 13 9 13 11 9 2
23 9 11 11 2 9 2 13 9 9 2 15 1 15 4 13 0 9 13 11 9 11 9 2
9 2 13 4 13 16 3 13 9 2
5 15 13 0 9 2
11 15 13 15 13 0 9 2 15 13 9 2
11 11 13 9 0 9 2 15 13 11 9 2
8 11 13 3 9 9 0 9 2
16 11 13 3 9 9 2 15 1 11 13 9 13 3 0 9 2
6 2 15 13 13 9 2
17 16 9 13 13 2 11 13 13 9 1 2 7 15 13 0 9 2
20 9 11 11 4 13 9 9 11 2 16 11 4 13 9 13 11 9 0 9 2
7 11 2 9 13 13 9 9
7 9 13 3 9 9 13 2
16 9 13 3 9 9 9 2 7 9 13 0 9 2 13 11 2
7 9 13 3 9 9 13 2
12 9 9 4 13 9 13 9 9 2 13 11 2
12 9 13 3 13 9 2 7 9 13 0 9 2
10 9 13 9 4 13 0 9 0 0 2
9 3 9 11 13 0 9 9 9 2
14 9 13 9 9 4 3 13 2 7 9 13 13 9 2
9 0 9 9 13 13 9 0 9 2
10 9 13 2 16 9 13 13 9 9 2
17 3 15 9 13 9 9 2 15 9 9 4 13 3 3 9 13 2
4 9 13 11 11
9 9 9 11 3 13 9 0 13 2
14 11 15 1 4 13 3 9 9 1 2 13 9 9 2
7 9 11 13 12 12 9 2
15 11 13 9 13 12 12 2 15 13 9 12 9 0 9 2
10 11 13 9 13 9 7 3 9 9 2
14 15 3 9 13 9 12 12 9 13 1 9 13 9 2
7 9 13 12 9 0 9 2
18 9 9 13 9 3 12 9 2 15 13 12 9 9 0 9 9 1 2
10 3 15 0 15 9 13 9 0 9 2
6 9 13 9 7 9 2
20 9 13 3 9 9 9 9 2 15 13 12 12 11 13 0 9 9 13 9 2
6 9 2 11 9 13 9
13 9 13 2 7 11 9 0 9 9 13 9 9 2
19 9 11 11 11 13 9 3 12 9 9 13 2 13 11 0 9 13 9 2
16 9 13 9 13 0 0 2 16 11 13 13 13 9 3 3 2
10 11 11 11 9 9 9 13 3 13 2
19 9 13 9 3 12 9 13 3 11 9 13 9 0 7 0 9 0 9 2
12 11 0 9 15 1 3 13 9 2 9 13 2
16 3 12 9 13 13 3 9 9 9 7 0 9 9 13 9 2
10 9 13 12 0 0 0 9 9 9 2
13 12 9 13 9 13 3 12 9 0 12 9 13 2
10 3 12 9 13 9 3 12 9 9 2
7 12 9 13 9 13 9 2
6 9 0 9 13 9 2
12 12 9 13 2 16 9 13 0 9 13 9 2
18 3 12 9 13 9 0 9 11 7 12 9 9 9 13 3 3 11 2
17 16 11 9 4 13 3 2 3 12 9 9 9 13 0 9 9 2
22 9 9 13 2 16 11 9 4 13 9 9 1 2 16 9 13 3 3 16 1 9 2
9 11 9 4 13 9 3 3 11 2
4 9 13 11 9
14 9 11 9 1 9 13 9 3 9 0 9 0 9 2
5 3 9 13 9 2
16 9 13 3 0 9 9 3 7 13 9 7 9 13 0 9 2
13 11 9 1 9 13 9 12 9 0 12 12 9 2
8 0 9 13 12 9 12 9 2
10 9 13 9 0 12 9 12 12 9 2
13 9 13 9 3 13 12 9 7 13 12 12 9 2
16 11 11 11 11 9 9 13 12 9 7 11 11 9 12 9 2
23 2 9 13 9 13 0 9 9 9 0 9 7 9 9 13 9 2 9 11 11 13 9 2
13 2 9 13 3 9 2 3 13 9 13 0 9 2
6 11 13 9 9 3 2
9 9 9 9 7 9 13 9 12 2
10 9 9 13 11 9 9 9 9 9 2
6 11 13 2 3 13 11
5 11 13 9 11 2
17 11 9 13 13 0 9 7 9 9 9 2 13 11 9 0 9 2
12 11 13 9 12 11 9 2 15 13 12 9 2
16 11 9 9 1 9 13 13 3 3 2 13 9 13 9 9 2
13 2 11 9 13 4 13 9 7 9 9 9 11 2
14 7 0 9 2 7 0 9 2 9 11 11 13 9 2
15 9 3 12 9 0 9 13 0 9 7 9 9 13 0 2
13 0 9 13 0 13 12 9 7 9 13 12 9 2
13 2 0 9 9 9 4 3 13 11 3 3 0 2
22 15 9 4 13 9 9 7 9 9 9 7 9 1 13 9 13 9 9 2 11 13 2
11 11 13 2 16 3 9 9 13 3 9 2
6 11 9 1 2 9 2
26 11 9 11 11 11 11 4 13 9 2 16 9 9 9 13 3 0 9 7 13 9 1 12 9 9 2
14 3 11 2 11 7 11 9 12 9 9 13 9 9 2
27 11 1 11 9 0 9 9 4 3 13 9 9 2 16 9 13 13 9 13 9 9 9 7 13 9 9 2
14 0 9 11 13 9 2 16 11 13 2 9 9 2 2
15 15 9 9 11 13 2 16 9 9 13 9 3 13 9 2
21 9 11 9 0 9 9 4 13 12 9 7 9 11 9 0 9 9 13 12 9 2
20 9 13 9 2 15 1 11 13 13 9 7 13 9 13 15 9 3 12 9 2
11 11 0 9 9 4 13 12 9 12 9 2
9 11 13 9 2 2 15 13 9 2
11 11 9 11 11 13 9 13 9 9 9 2
10 9 9 1 11 4 13 0 9 9 2
18 11 9 11 11 13 9 13 9 9 13 9 2 11 11 11 9 13 2
15 9 9 13 13 2 16 11 11 13 9 13 9 9 9 2
10 9 13 2 16 15 9 13 3 9 2
23 2 15 13 0 0 2 0 7 0 9 11 0 2 0 7 0 9 2 9 13 9 13 2
9 11 9 11 11 4 13 9 0 2
16 9 13 0 9 0 9 2 15 9 9 13 15 9 7 9 2
11 0 9 4 13 9 2 15 13 3 9 2
9 3 11 4 13 9 11 13 9 2
19 2 11 4 13 0 9 7 9 9 2 15 4 13 11 9 2 9 13 2
10 3 15 9 13 4 13 9 11 1 2
22 2 13 3 3 2 16 15 9 13 15 9 2 11 11 11 13 11 11 9 11 13 2
12 9 9 9 1 9 4 13 11 0 9 9 2
6 11 13 7 3 13 9
8 11 9 4 3 13 0 9 2
8 3 3 11 9 4 13 0 2
6 11 13 3 3 3 2
7 11 0 9 13 9 3 2
7 11 9 13 9 0 9 2
22 3 9 9 13 3 9 9 2 15 3 13 0 0 9 9 9 13 9 3 9 3 2
11 11 9 9 11 4 9 12 13 12 9 2
7 13 9 13 12 9 9 2
13 9 4 13 12 12 9 2 15 11 12 12 9 2
11 11 1 9 13 11 2 11 9 7 11 2
17 9 11 5 11 13 13 11 0 9 9 12 9 9 11 9 11 2
6 0 9 9 13 11 2
12 0 9 11 13 2 16 11 13 0 11 9 2
9 9 1 0 9 11 13 11 1 2
9 11 9 4 13 12 9 12 9 2
13 9 11 13 2 16 15 4 13 9 9 11 9 2
18 11 3 13 12 11 7 15 0 9 11 11 9 11 2 11 7 11 2
15 9 9 11 13 9 12 12 0 9 11 7 11 11 9 2
7 11 9 4 13 12 9 2
21 9 11 11 13 13 11 11 9 9 2 0 2 2 16 15 3 13 2 13 2 2
10 11 11 9 9 4 9 13 12 9 2
9 9 11 11 9 13 12 9 9 2
14 9 11 11 13 3 11 9 9 0 12 9 12 9 2
10 9 11 13 13 9 7 13 9 9 2
7 9 9 13 9 9 1 2
6 9 13 3 9 9 2
7 9 9 13 12 9 9 2
6 12 0 13 13 13 9
14 9 9 9 13 13 13 3 2 16 0 9 13 0 2
11 11 11 11 0 9 4 13 11 0 9 2
17 0 9 4 13 11 1 15 9 15 2 15 4 13 13 9 9 2
12 15 3 4 13 9 7 13 3 9 7 9 2
19 11 13 3 3 0 9 0 9 2 15 1 9 7 9 13 3 12 9 2
8 13 7 9 1 7 15 1 2
6 13 9 7 13 15 2
6 13 7 0 7 0 2
13 15 0 9 13 3 3 9 7 0 15 13 9 2
7 9 9 13 0 9 9 2
10 16 9 13 2 15 13 3 4 13 2
24 15 9 0 9 13 3 0 9 2 15 13 13 3 3 2 16 9 13 0 13 0 9 9 2
19 15 9 15 4 13 9 2 16 9 9 13 13 2 7 15 13 9 1 2
2 9 9
8 9 9 4 13 0 0 9 2
11 9 1 13 3 9 2 16 9 13 9 2
12 11 7 11 0 9 4 13 9 0 0 9 2
15 15 9 13 3 9 2 16 9 13 3 15 9 13 9 2
8 3 9 13 13 7 13 9 2
8 9 9 13 13 3 16 9 2
9 3 0 9 13 13 15 9 0 2
19 0 9 13 3 3 9 11 11 9 2 15 15 13 9 9 13 9 9 2
9 11 1 9 13 9 3 3 9 2
17 11 9 1 13 9 2 16 9 9 9 13 3 0 16 9 9 2
9 9 13 4 3 13 3 9 9 2
19 13 0 13 0 9 2 16 15 9 13 2 16 15 9 9 13 13 13 2
10 9 9 0 9 13 3 9 16 9 2
14 15 13 2 16 15 9 1 13 9 1 12 9 9 2
12 3 4 13 2 16 2 9 9 13 9 2 2
3 9 9 1
13 3 3 13 13 2 3 12 9 9 13 0 9 2
8 9 9 15 9 13 3 3 2
12 3 15 9 13 13 7 13 9 9 7 15 2
11 15 9 9 9 3 9 4 13 13 13 2
12 15 9 9 13 13 0 2 13 9 9 2 2
8 0 11 13 15 9 3 9 2
12 9 4 13 0 9 2 15 9 13 13 13 2
10 4 13 3 3 9 2 9 7 9 2
9 3 15 4 13 9 1 3 9 2
10 11 4 13 11 0 9 13 9 9 2
20 9 4 13 15 9 13 9 0 9 2 16 3 9 4 13 3 9 16 9 2
16 9 9 11 2 9 13 9 2 9 13 15 9 3 0 9 2
4 9 13 13 11
11 11 9 11 13 13 9 15 9 0 9 2
18 9 4 13 12 12 9 9 9 2 15 13 9 9 13 9 0 9 2
14 11 9 13 13 13 9 9 13 13 11 7 0 9 2
23 9 4 13 12 12 9 2 3 12 12 9 2 9 9 2 15 13 9 13 0 9 9 2
9 11 13 9 9 3 11 0 9 2
14 9 12 13 9 9 13 9 13 11 9 13 3 11 2
30 9 13 3 12 0 9 9 2 7 13 3 3 9 3 2 11 0 9 2 7 2 9 11 2 2 11 11 11 13 2
15 9 13 11 7 11 12 0 9 4 13 3 0 7 0 2
8 9 13 13 3 11 13 9 2
13 7 11 7 11 13 9 9 7 13 13 9 3 2
3 11 13 9
11 9 11 0 9 13 0 9 0 9 3 2
6 9 13 7 9 13 2
6 0 9 9 13 3 2
15 2 11 9 11 9 1 13 9 9 4 0 9 13 9 2
15 4 3 13 3 15 3 0 9 2 9 11 11 13 9 2
16 11 9 9 4 13 2 15 11 1 13 3 11 13 9 9 2
8 3 15 9 4 9 13 3 2
7 3 3 9 4 13 9 2
11 9 11 13 9 12 9 0 12 12 9 2
10 9 13 12 12 9 7 12 9 9 2
10 0 9 9 13 3 0 2 12 9 2
11 9 1 9 13 12 12 9 12 12 9 2
5 9 13 3 9 2
10 9 11 13 9 9 13 12 12 9 2
7 9 13 12 12 9 9 2
8 0 9 13 12 9 12 9 2
8 11 4 13 0 9 9 3 2
15 9 13 9 13 3 15 9 0 9 7 9 1 9 13 2
6 11 2 11 13 16 9
21 11 9 11 11 13 11 9 9 2 15 13 13 9 1 7 13 9 9 15 9 2
17 11 9 11 11 13 11 9 2 9 2 2 13 11 11 11 11 2
22 2 11 13 13 0 9 2 15 13 9 15 13 9 2 11 13 0 9 13 9 3 2
6 2 11 13 9 9 2
13 11 1 9 13 11 9 3 2 13 0 9 2 2
17 11 13 2 16 16 9 9 13 0 9 2 11 3 13 9 9 2
9 11 9 13 15 9 9 9 9 2
20 3 9 12 11 13 9 12 9 9 2 7 15 9 9 13 13 12 9 9 2
8 11 13 9 3 12 9 9 2
17 16 9 9 13 3 2 11 9 13 11 11 9 1 9 9 9 2
8 9 2 11 13 11 7 11 9
16 9 11 4 13 9 11 7 9 11 9 9 2 11 9 13 2
8 9 13 9 7 9 9 9 2
24 11 4 13 0 0 9 9 9 2 9 7 9 9 2 7 11 1 9 13 4 13 12 9 2
18 11 13 3 13 9 9 2 7 9 7 9 1 11 13 9 13 15 2
7 11 13 3 3 3 9 2
22 11 9 1 15 4 13 0 9 9 3 12 9 9 2 7 0 9 13 15 0 9 2
8 9 9 13 0 9 11 9 2
7 11 1 11 13 9 9 2
15 11 4 13 9 9 2 7 3 9 7 9 13 9 9 2
10 11 1 3 9 13 4 13 12 9 2
9 11 13 4 3 13 9 9 13 2
11 11 13 2 16 15 13 13 9 1 9 2
25 11 9 13 11 11 13 11 9 2 16 11 13 13 9 3 9 2 15 15 9 13 13 15 9 2
13 11 13 3 13 13 11 13 9 7 11 13 9 2
3 9 13 9
11 9 11 1 9 13 9 13 3 15 3 2
17 11 4 13 9 0 9 2 7 15 9 9 9 9 13 12 9 2
10 9 0 9 9 13 12 9 0 9 2
16 11 13 9 9 12 9 2 7 15 11 13 0 9 12 9 2
11 9 13 9 12 9 0 12 12 13 9 2
9 9 13 3 0 11 7 11 9 2
8 3 13 0 9 12 12 9 2
21 9 2 11 2 11 7 11 2 13 12 12 7 0 7 0 11 3 12 12 9 2
12 11 4 13 0 9 0 9 1 9 0 9 2
10 9 4 13 0 2 13 15 13 9 2
16 15 9 0 9 0 9 9 13 12 9 0 9 12 12 9 2
27 11 9 13 15 2 16 9 13 0 0 9 3 11 2 11 2 11 2 11 2 11 11 2 11 7 11 2
14 11 13 0 9 3 11 2 15 15 9 13 12 9 2
3 11 11 9
9 9 9 11 1 13 9 11 9 2
16 9 9 13 11 9 13 12 9 7 9 13 3 12 12 9 2
10 9 9 11 13 11 1 9 0 9 2
13 11 9 4 13 11 7 11 1 9 0 0 9 2
17 11 9 4 13 0 13 9 2 11 2 11 2 11 7 11 2 2
10 9 1 11 4 13 0 3 9 9 2
8 11 1 11 4 13 11 1 2
13 9 0 9 9 13 0 9 12 9 12 12 9 2
26 2 11 9 13 2 16 15 0 9 9 4 13 3 3 3 0 9 3 11 2 11 9 11 11 13 2
13 2 11 13 3 0 9 13 9 9 7 13 9 2
4 11 9 9 0
13 11 13 11 1 3 2 7 9 13 13 9 0 2
24 15 9 16 11 7 0 9 9 4 13 3 3 0 2 4 11 9 13 9 9 13 0 9 2
17 0 9 0 9 13 12 12 9 2 12 9 3 16 0 9 9 2
10 0 9 9 9 9 13 0 9 0 2
9 11 4 13 3 9 11 7 9 2
19 9 11 2 15 13 7 11 7 11 9 9 2 13 11 13 9 12 9 2
13 15 9 11 9 11 13 12 9 0 9 12 9 2
19 9 11 11 11 2 11 2 9 13 11 12 9 0 9 0 9 12 9 2
17 11 0 9 13 3 0 11 13 2 15 11 13 9 12 9 9 2
7 11 2 9 13 13 9 9
13 9 13 0 7 9 13 9 2 11 13 9 13 2
13 9 13 3 0 13 9 7 9 2 16 9 13 2
15 9 13 9 2 15 13 0 3 2 16 9 13 0 9 2
19 11 9 13 9 9 9 13 3 2 16 9 0 9 13 3 12 12 9 2
21 3 12 12 9 9 9 13 9 12 9 13 9 3 7 12 9 4 3 13 15 2
20 12 12 2 12 12 9 9 12 9 13 9 3 7 12 9 4 3 13 15 2
9 9 9 13 2 7 3 9 13 2
24 16 0 9 13 3 12 12 9 2 3 12 9 13 9 3 7 3 12 9 4 3 13 15 2
16 9 1 9 13 0 3 13 9 13 9 9 2 16 9 13 2
20 3 3 9 3 12 12 9 9 13 9 13 2 16 9 9 13 9 9 9 2
22 9 13 13 0 13 2 16 12 12 9 9 9 13 3 0 2 16 9 13 9 0 2
8 9 13 9 13 3 12 9 2
6 9 9 13 12 9 2
6 9 2 11 7 11 9
18 12 11 7 11 0 9 13 13 13 9 7 9 9 1 2 11 13 2
15 11 7 11 0 9 13 9 12 9 2 16 11 13 9 2
16 9 13 13 12 11 13 9 9 2 16 9 4 13 11 9 2
17 9 13 13 13 9 2 16 11 9 9 13 0 13 9 0 9 2
11 0 9 13 9 13 12 9 9 11 11 2
15 16 9 13 13 9 2 15 9 13 13 13 2 11 13 2
3 9 13 9
6 9 9 4 13 9 2
8 9 1 9 13 13 9 13 2
7 0 9 1 9 9 13 2
9 15 9 13 9 13 3 3 3 2
18 9 9 2 11 2 7 11 9 9 2 11 2 0 9 4 13 9 2
12 11 7 11 13 9 11 11 9 3 0 9 2
8 9 13 13 9 13 9 1 2
11 9 13 9 9 2 9 7 9 0 9 2
11 9 9 13 9 13 3 13 9 9 13 2
13 9 1 9 13 0 9 12 1 12 9 0 9 2
13 9 13 3 12 9 9 9 13 9 1 13 9 2
13 0 9 9 9 13 0 9 1 12 9 0 9 2
11 3 0 9 13 9 9 13 13 13 9 2
8 9 13 3 0 9 12 1 2
15 11 9 11 11 13 11 2 16 9 13 0 7 0 9 2
19 2 9 13 3 13 3 0 2 7 3 3 9 15 13 2 11 13 11 2
11 2 9 13 0 0 7 15 9 3 0 2
21 15 9 13 2 16 0 9 13 0 16 9 9 2 11 9 11 11 13 9 11 2
7 11 2 9 9 4 13 9
17 9 13 9 13 9 0 9 2 15 4 13 9 9 2 13 11 2
8 11 1 9 13 3 0 9 2
12 3 0 9 13 12 9 3 9 16 0 9 2
6 9 13 3 3 9 2
10 2 3 9 0 9 13 15 9 0 2
17 15 9 13 3 15 9 0 2 9 7 9 9 9 11 11 13 2
19 0 9 9 1 9 7 9 9 9 13 3 0 11 2 11 7 11 1 2
9 9 13 3 0 9 7 0 9 2
7 3 3 9 11 7 11 2
8 11 9 13 3 16 15 9 2
25 2 3 11 4 13 3 0 9 2 7 13 9 9 3 2 9 9 7 9 11 9 11 11 13 2
3 9 13 9
9 0 9 9 13 0 9 9 13 2
6 3 9 13 3 3 2
9 15 9 9 4 13 12 12 9 2
10 9 13 12 9 0 9 0 9 13 2
7 9 13 12 12 0 9 2
10 9 0 13 0 9 13 12 9 3 2
8 9 13 0 9 12 13 9 2
10 9 13 12 9 3 16 0 9 9 2
20 13 9 4 13 12 12 0 9 2 15 13 12 9 3 0 9 0 9 13 2
8 9 13 3 9 9 13 9 2
6 9 13 9 9 3 13
14 16 9 7 9 13 9 2 9 13 15 15 9 3 2
8 3 3 13 9 13 15 3 2
7 9 13 3 11 9 9 2
11 9 13 0 9 9 2 15 13 9 9 2
11 9 9 9 13 3 16 15 15 9 9 2
8 3 12 9 9 13 15 9 2
13 9 7 9 1 13 9 13 3 9 3 16 9 2
13 11 13 13 3 9 9 0 9 2 9 9 13 2
18 16 12 12 9 7 9 13 9 0 9 2 3 9 9 13 15 9 2
5 9 9 13 13 2
8 9 12 9 13 9 0 9 2
6 3 11 9 13 3 2
7 11 7 11 9 13 3 2
14 9 12 9 13 13 15 2 16 9 9 13 9 9 2
8 0 9 9 0 13 12 9 2
10 9 9 3 0 13 9 9 0 9 2
6 3 13 12 9 9 2
10 9 13 0 12 9 7 9 12 9 2
5 11 0 9 13 11
7 9 11 9 13 3 9 2
11 9 13 11 11 2 15 13 3 9 9 2
9 9 1 11 9 9 13 13 0 2
12 9 11 13 7 13 11 11 13 15 12 9 2
12 9 13 12 12 9 2 15 11 12 12 9 2
13 11 1 0 9 13 11 2 11 2 11 7 11 2
7 9 11 13 13 9 11 2
4 9 13 13 2
14 9 13 2 16 9 13 9 9 11 2 11 7 11 2
5 9 13 12 9 2
10 9 11 9 13 12 9 13 11 9 2
10 3 11 11 9 13 0 12 9 9 2
13 9 11 11 13 11 11 9 9 12 9 12 9 2
12 9 13 3 13 11 13 9 11 11 0 9 2
9 9 13 9 9 13 9 11 9 2
6 9 9 13 12 9 2
7 11 7 11 13 3 9 2
14 11 13 2 16 9 0 9 9 13 0 9 9 1 2
9 9 9 13 12 9 9 9 13 2
11 9 11 13 9 0 9 7 0 9 9 2
7 9 9 9 13 12 9 2
7 9 11 13 3 9 9 2
8 9 1 0 9 13 13 0 2
5 9 13 12 9 2
4 9 9 13 3
7 9 13 11 9 9 12 2
11 9 13 9 7 9 9 9 3 0 3 2
11 3 9 9 13 13 3 2 0 9 13 2
16 9 11 13 9 13 12 9 2 15 13 3 12 9 15 9 2
8 9 4 13 12 9 9 13 2
13 9 1 9 13 13 9 3 12 12 9 0 9 2
8 9 13 3 12 9 9 13 2
8 3 13 9 9 7 9 9 2
22 2 9 4 13 7 13 13 0 0 9 9 9 2 11 9 13 9 11 11 13 9 2
14 9 9 13 0 9 2 16 0 9 9 13 12 9 2
6 11 9 2 3 12 9
11 11 7 11 0 9 4 13 15 9 9 2
11 12 9 9 1 4 13 3 12 12 9 2
10 11 7 11 0 9 13 9 9 9 2
8 0 15 13 13 0 11 11 2
22 11 11 11 7 11 13 9 12 12 9 2 15 13 12 9 0 16 0 9 9 1 2
7 11 11 13 3 3 9 2
17 15 13 12 12 9 2 15 13 12 9 0 16 0 9 0 9 2
7 0 9 13 12 1 9 2
10 0 9 13 9 11 9 13 11 11 2
13 15 13 9 13 11 9 12 9 3 12 12 9 2
15 11 0 9 13 12 12 9 2 15 13 9 9 12 9 2
7 3 9 11 13 15 9 2
17 3 11 2 11 7 11 11 9 13 11 7 11 1 12 12 9 2
18 16 3 13 12 9 13 11 11 9 2 9 9 9 13 3 12 12 2
16 9 13 0 9 9 2 3 3 13 9 9 13 0 12 12 2
9 3 0 13 13 11 11 0 9 2
21 9 9 13 9 1 11 13 9 13 9 9 2 16 9 9 13 12 9 0 9 2
9 11 13 15 9 11 1 11 9 2
6 11 9 2 11 13 11
13 11 7 11 9 13 3 13 9 13 9 9 9 2
19 11 9 13 2 16 9 11 11 11 11 13 9 13 9 7 13 11 9 2
11 11 13 9 1 9 9 2 9 11 13 2
14 11 13 3 9 9 9 11 11 7 9 9 11 11 2
8 9 4 3 13 9 0 9 2
13 11 13 9 9 12 13 15 0 9 7 9 1 2
23 2 15 2 16 11 4 13 9 2 13 16 9 13 0 2 9 9 11 11 13 9 11 2
2 9 13
29 9 0 11 9 13 9 4 13 13 12 9 7 15 9 2 15 13 3 3 16 11 2 11 7 11 4 13 9 2
16 0 9 9 13 9 9 9 2 11 12 9 7 11 12 9 2
23 9 11 11 13 13 3 12 9 13 9 7 9 15 2 16 11 13 13 9 9 0 9 2
16 11 9 11 11 13 9 11 9 7 9 9 9 9 11 11 2
18 11 13 2 16 9 13 2 15 9 2 2 15 12 9 9 13 3 2
10 11 3 13 9 2 0 7 0 2 2
7 11 2 9 9 13 13 9
12 11 1 15 9 4 13 2 7 9 13 9 2
5 9 13 3 0 2
8 11 13 9 13 9 0 9 2
19 0 9 4 13 9 9 2 3 0 9 9 13 13 3 9 13 9 1 2
21 9 13 3 9 12 9 9 2 16 11 9 7 9 9 0 9 13 13 3 9 2
12 9 13 9 3 3 9 9 2 9 7 9 2
3 0 9 9
12 0 9 13 0 9 7 9 3 12 9 9 2
12 11 9 9 11 13 0 9 7 9 9 9 2
19 9 7 9 13 3 12 12 9 9 13 9 2 9 9 13 9 11 11 2
21 9 13 2 16 15 4 13 9 3 9 2 16 9 4 13 0 9 9 0 9 2
12 3 9 13 2 13 9 13 9 3 9 11 2
12 11 4 13 0 9 2 15 13 3 9 9 2
7 3 15 13 2 9 9 9
10 11 9 4 13 9 9 0 0 9 2
6 9 9 13 3 13 2
7 9 13 9 9 3 9 2
17 9 9 13 11 0 9 9 13 0 0 9 9 0 9 11 9 2
14 9 13 3 9 12 3 13 0 9 2 11 2 9 2
22 11 7 11 4 9 9 1 9 13 0 9 9 9 15 9 16 0 9 11 0 9 2
8 9 13 9 13 9 13 9 2
18 3 9 4 3 13 9 9 2 16 9 9 11 13 9 9 13 13 2
8 9 9 13 15 11 9 9 2
10 9 13 9 13 9 15 13 9 9 2
6 2 9 13 11 9 2
16 11 13 9 13 9 3 0 9 11 2 0 0 9 13 9 2
15 11 0 9 13 2 16 9 1 11 9 4 3 13 9 2
21 0 9 9 9 2 15 13 13 9 2 7 9 9 13 0 9 1 9 0 9 2
16 2 4 13 11 9 9 9 2 11 9 11 11 13 11 1 2
28 9 1 3 11 9 11 11 2 15 4 3 13 9 11 9 2 13 2 16 2 9 0 9 4 3 13 2 2
8 2 9 13 13 1 0 9 2
13 0 9 7 0 9 4 13 9 9 13 0 9 2
21 15 13 15 2 16 9 13 0 9 7 9 2 7 9 7 9 13 15 9 0 2
29 11 11 9 9 9 11 11 13 3 2 16 9 13 0 0 9 2 9 9 2 7 9 0 9 7 3 9 9 2
14 11 9 9 13 13 9 2 15 9 4 13 11 9 2
11 2 15 13 3 0 9 11 0 9 1 2
21 3 13 0 0 9 16 11 2 3 3 9 2 11 9 9 9 9 11 11 13 2
15 11 1 9 9 4 13 3 2 7 9 9 9 3 13 2
13 3 13 9 9 9 9 9 9 4 13 13 3 2
30 2 3 3 4 13 9 2 16 9 9 4 13 0 9 9 9 2 15 9 7 9 9 4 13 3 3 2 11 13 2
6 2 0 13 13 9 2
14 11 11 13 3 0 2 16 9 13 9 13 3 9 2
18 16 9 13 13 7 13 3 2 15 13 13 13 9 2 16 9 13 2
16 2 13 3 13 13 3 15 2 15 0 12 9 9 4 13 2
21 15 9 13 0 9 2 15 13 0 3 13 3 0 9 7 9 9 2 11 13 2
6 9 4 13 3 9 2
13 11 9 13 0 9 0 9 2 15 13 9 9 2
9 2 9 9 13 13 3 16 13 2
19 3 4 13 0 9 3 7 13 2 16 1 0 0 9 0 9 13 0 2
14 0 9 13 3 3 0 9 2 16 9 4 13 9 2
6 2 9 13 0 9 2
11 9 15 13 9 9 9 9 2 11 13 2
7 2 11 13 11 13 9 2
16 0 9 0 0 9 11 11 1 9 9 9 13 4 13 3 2
14 15 1 9 9 0 9 4 13 0 9 1 0 9 2
16 2 0 9 9 13 13 9 2 15 1 9 13 13 9 9 2
14 15 13 13 12 0 9 2 12 9 7 12 0 9 2
23 9 13 13 3 0 2 16 0 9 9 13 13 0 7 13 9 9 7 9 2 15 13 2
20 11 9 1 11 9 0 9 13 13 7 9 13 3 9 13 7 9 13 9 2
14 11 9 13 0 9 0 2 16 15 13 9 0 9 2
17 11 13 3 3 13 11 11 11 9 11 0 0 9 2 11 13 2
22 11 9 11 11 13 11 9 13 2 16 15 13 9 13 9 2 15 13 3 9 9 2
11 2 13 15 3 0 13 2 16 13 3 2
7 15 13 0 0 9 9 2
10 9 11 9 9 13 13 15 0 9 2
11 2 15 9 4 13 13 3 3 12 9 2
7 15 13 3 3 0 9 2
4 9 1 15 9
23 11 13 11 9 7 9 9 13 9 2 15 0 9 4 13 11 9 9 11 11 11 9 2
33 11 0 9 9 0 9 2 9 9 2 9 7 9 11 9 9 2 13 2 0 9 7 9 9 7 9 13 1 9 12 0 9 2
10 9 13 13 0 9 0 9 7 9 2
8 9 9 13 9 3 16 3 2
17 9 13 15 0 9 2 15 9 7 9 13 13 9 9 7 9 2
12 9 13 2 15 13 0 9 9 7 9 9 2
9 3 9 13 9 7 9 9 9 2
10 3 9 0 9 7 9 9 13 9 2
13 0 13 9 0 9 0 9 2 9 7 0 9 2
9 0 9 13 9 9 1 9 3 2
27 9 13 2 0 0 7 0 9 9 2 9 2 9 7 0 9 13 9 13 7 3 15 13 9 7 9 2
8 12 9 13 3 3 9 9 2
25 9 13 3 15 2 3 13 0 9 7 9 9 2 15 13 3 0 9 2 9 2 9 7 9 2
11 9 13 0 9 7 9 9 9 0 9 2
10 11 9 9 9 13 9 13 9 9 2
26 2 3 0 0 9 9 13 0 9 9 2 15 15 3 13 9 2 13 3 13 0 9 13 11 11 2
22 9 7 9 13 3 3 0 2 16 9 7 9 13 9 2 15 13 13 7 9 1 2
11 0 9 0 9 13 13 9 9 7 9 2
15 0 11 13 3 13 2 16 3 0 9 13 9 13 9 2
7 13 9 13 3 0 9 2
14 0 9 13 3 3 3 3 9 9 7 9 9 9 2
26 2 15 1 16 11 9 0 9 13 9 7 0 9 9 2 13 9 7 9 13 11 15 9 1 9 2
19 9 12 11 9 11 13 9 0 9 4 13 9 11 4 3 13 9 9 2
15 15 1 11 9 9 13 13 9 13 11 11 7 11 11 2
3 9 13 9
10 9 9 13 13 9 0 9 9 9 2
13 9 13 9 9 9 2 15 4 13 0 9 9 2
14 15 1 9 9 13 9 7 13 13 0 9 9 9 2
22 2 15 13 15 15 9 9 9 2 3 4 13 3 0 9 2 13 9 13 11 11 2
14 9 13 9 9 9 13 0 9 9 2 3 0 9 2
6 3 9 13 9 9 2
17 2 9 9 13 9 13 13 9 15 2 16 9 4 13 0 9 2
16 15 13 15 2 16 9 13 13 9 7 13 9 2 11 13 2
7 11 11 13 9 9 9 2
5 15 9 15 13 2
15 2 9 9 13 9 13 0 9 9 9 7 15 9 9 2
18 16 15 13 2 15 4 13 9 15 9 2 13 0 9 2 11 13 2
6 15 15 9 3 13 2
14 9 9 9 9 4 13 3 0 9 9 3 0 9 2
23 2 11 11 2 15 13 9 2 13 9 2 15 13 13 9 9 7 9 13 3 9 9 2
15 9 4 13 3 0 3 13 0 2 16 9 13 3 0 2
8 11 7 12 9 9 13 9 13
11 9 13 9 9 0 9 11 9 13 9 2
8 9 9 11 9 13 9 9 2
18 11 9 13 0 2 7 9 13 0 13 2 16 0 9 13 3 13 2
17 2 13 3 11 9 7 9 13 3 11 11 2 13 9 11 11 2
29 9 0 9 13 9 2 16 9 13 11 9 13 11 7 12 9 9 2 15 13 0 7 0 9 9 9 7 9 2
14 11 7 12 9 9 13 0 9 11 9 9 13 9 2
17 2 9 13 13 9 2 15 9 9 3 13 2 13 9 11 11 2
10 11 7 12 9 9 13 9 9 1 2
13 11 11 13 9 2 16 9 9 13 11 0 9 2
14 2 3 9 13 13 13 9 2 13 0 9 13 13 2
8 11 11 9 13 9 9 9 2
11 2 13 9 13 0 9 2 11 13 9 2
13 2 9 13 3 13 13 2 13 9 3 0 9 2
14 16 9 13 3 9 7 9 2 13 15 9 3 0 2
15 11 13 2 16 11 4 13 0 9 2 16 13 9 9 2
9 2 13 15 13 9 2 11 13 2
6 15 13 3 2 9 2
11 15 1 9 9 13 13 3 3 0 13 2
4 9 13 9 2
6 12 9 13 9 9 2
26 11 13 2 16 11 2 11 7 11 13 15 11 0 9 13 15 9 3 16 9 13 7 9 13 11 2
12 11 13 2 16 11 7 12 9 9 13 0 2
15 2 9 13 15 2 3 9 4 11 13 15 12 9 2 2
6 11 11 13 9 9 2
5 2 9 13 15 2
19 11 13 13 9 2 11 11 7 11 11 2 15 15 13 9 2 9 9 2
9 13 9 1 11 9 2 11 13 2
3 9 9 9
18 11 9 13 9 11 9 13 9 9 7 9 9 3 3 12 12 9 2
8 9 11 11 13 11 11 9 2
15 9 11 11 13 11 11 9 9 9 9 7 0 9 9 2
17 9 13 11 9 9 11 11 13 11 11 13 0 9 9 9 9 2
29 9 9 13 9 13 9 9 11 11 7 11 11 9 11 9 13 9 2 16 15 9 13 9 2 9 13 9 13 2
11 0 9 4 13 9 13 15 9 13 9 2
10 11 11 4 13 0 9 9 9 9 2
19 15 13 13 7 13 9 2 15 13 2 16 13 9 9 9 13 0 9 2
11 3 3 15 9 4 13 0 9 9 9 2
23 11 4 13 9 1 9 2 7 3 11 7 11 9 4 3 12 9 13 3 0 16 11 2
7 3 9 13 3 12 9 2
12 11 9 9 13 3 3 9 9 0 9 9 2
17 9 13 3 12 9 2 15 12 13 9 2 12 9 7 12 9 2
12 9 13 11 9 9 11 11 9 11 11 13 2
15 0 9 13 2 12 12 9 9 13 12 7 0 9 12 2
25 0 9 13 9 11 11 2 9 11 11 7 9 9 11 11 7 9 9 11 11 7 9 11 11 2
12 3 0 9 9 4 15 9 13 9 9 9 2
10 9 13 9 7 9 12 12 9 9 2
8 9 9 13 12 11 9 9 2
26 9 9 13 0 3 7 3 13 9 7 9 11 1 2 15 1 15 9 13 3 9 9 3 3 0 2
20 9 9 0 9 13 9 11 11 2 15 13 9 3 9 11 11 1 9 12 2
12 11 11 13 11 9 9 9 13 15 9 9 2
14 9 13 9 11 11 9 9 2 0 9 7 13 9 2
27 2 15 0 9 2 3 9 11 11 2 4 13 3 0 9 7 13 9 13 3 3 9 9 2 13 11 2
6 11 9 13 0 9 11
17 2 0 9 4 13 3 2 2 11 11 13 9 9 9 13 9 2
19 9 13 9 0 9 13 9 13 11 13 9 7 9 13 9 13 9 9 2
18 9 13 9 11 11 2 11 2 11 2 13 11 9 13 0 11 9 2
15 2 9 13 13 3 0 9 2 15 7 13 7 13 13 2
15 3 13 9 2 15 13 9 2 16 15 9 13 15 9 2
13 11 11 2 9 0 2 1 11 13 13 3 9 2
23 2 11 11 13 7 3 0 2 16 15 4 13 2 7 3 0 2 16 15 13 4 13 2
14 9 13 3 9 2 15 11 9 7 15 9 4 13 2
7 2 15 4 13 1 9 2
9 0 9 4 13 3 2 11 13 2
17 9 11 11 11 9 13 13 0 9 2 11 2 9 11 9 9 2
9 2 9 13 9 13 2 11 13 2
17 11 13 11 9 9 3 9 15 2 3 11 9 3 13 9 9 2
23 15 13 3 2 16 11 9 7 15 11 9 13 9 13 3 9 13 11 9 9 13 9 2
10 9 11 11 13 9 3 11 0 9 2
14 2 13 9 2 16 0 9 13 7 13 15 13 9 2
9 9 7 9 9 13 13 9 9 2
12 9 11 11 13 2 16 9 4 13 0 9 2
11 9 13 11 9 9 9 7 9 9 9 2
13 2 9 4 13 2 15 4 13 9 3 0 9 2
6 9 13 13 0 9 2
12 9 13 3 1 11 9 0 9 7 0 9 2
10 11 13 9 3 9 11 9 9 9 2
8 2 9 4 9 13 3 3 2
6 3 0 9 13 3 2
3 9 0 9
14 11 9 13 3 12 9 0 9 7 9 9 13 9 2
12 11 9 13 9 9 9 13 3 12 12 9 2
12 9 9 9 9 13 3 12 9 7 12 9 2
6 9 12 13 11 9 2
20 9 11 11 13 9 0 7 0 9 7 9 9 11 13 9 13 12 12 9 2
36 9 11 11 9 11 11 11 11 11 11 11 2 11 11 11 13 12 12 9 7 9 11 11 11 13 11 11 11 11 11 2 9 12 12 9 2
39 0 0 9 13 9 2 9 11 11 13 9 2 15 9 13 11 11 11 11 11 11 11 11 2 11 11 11 11 11 11 11 11 2 2 12 12 9 2 2
51 15 13 9 13 11 9 9 9 9 2 12 12 9 2 2 9 11 11 9 7 9 13 9 11 9 2 12 12 9 2 7 9 9 11 11 9 9 7 15 9 9 13 9 13 9 2 12 12 9 2 2
11 11 9 9 9 11 11 13 11 9 9 2
15 2 3 0 9 11 9 9 9 13 9 9 9 11 9 2
20 12 13 9 13 3 3 9 0 9 2 0 9 7 0 9 9 2 11 13 2
25 11 9 13 3 3 13 9 2 15 9 13 13 0 9 7 13 9 0 9 0 9 7 9 9 2
13 9 9 9 9 13 13 9 9 7 0 9 9 2
24 11 9 9 4 13 0 9 2 9 0 9 4 13 3 3 12 9 2 9 2 9 7 9 2
14 2 9 4 3 13 0 9 7 9 9 13 0 9 2
17 13 0 9 13 9 13 9 9 3 2 11 9 9 11 11 13 2
7 2 9 13 9 0 9 2
12 11 9 13 0 9 9 7 9 9 15 9 2
8 9 13 0 9 9 9 9 2
16 9 13 3 9 9 7 13 9 4 13 12 9 7 9 1 2
18 2 15 9 13 9 11 9 1 7 15 9 13 3 0 2 11 13 2
13 15 0 9 13 11 9 13 11 9 9 11 11 2
7 2 13 13 9 9 9 2
10 9 13 11 9 9 9 2 11 13 2
9 9 13 0 9 0 13 9 1 2
9 12 9 13 3 12 9 9 0 2
21 9 13 11 9 9 2 15 9 13 13 0 9 2 9 7 9 2 9 3 9 2
4 9 13 9 9
11 0 9 9 12 13 9 9 7 9 9 2
8 0 9 9 13 0 9 12 2
7 15 9 9 13 9 9 2
18 9 13 0 2 16 11 9 4 13 9 9 7 15 13 3 13 9 2
19 11 9 9 9 4 13 3 9 9 13 9 2 13 9 13 9 11 11 2
14 2 9 9 4 13 3 2 16 15 13 3 9 9 2
12 9 13 13 9 9 9 0 9 2 11 13 2
15 9 9 13 9 3 9 9 9 2 9 9 7 9 9 2
5 11 2 9 7 9
21 11 9 9 9 13 9 9 9 2 15 13 12 9 0 9 7 13 11 11 9 2
17 9 11 11 4 13 9 11 11 9 7 9 9 9 7 11 9 2
16 9 13 15 13 11 9 13 9 11 9 9 0 7 0 9 2
18 11 9 1 9 9 13 0 9 2 16 9 9 0 9 9 13 0 2
23 3 2 9 13 11 2 13 0 2 16 11 13 3 3 11 7 15 11 9 13 0 9 2
20 9 11 13 11 1 13 9 9 3 13 9 7 3 3 0 7 0 9 1 2
14 9 4 13 9 9 7 9 2 7 13 3 0 9 2
26 9 9 11 4 13 9 12 13 9 7 13 13 9 9 9 9 9 7 15 13 9 13 9 9 9 2
15 9 9 13 0 9 9 13 9 7 15 9 9 7 9 2
16 9 13 9 15 0 9 2 15 9 9 9 9 13 0 9 2
8 3 13 0 12 9 11 9 2
7 3 13 15 9 9 9 2
11 3 9 12 9 13 9 3 3 12 9 2
26 9 2 9 7 9 2 13 11 1 3 11 13 0 9 2 15 0 9 13 9 9 2 9 7 9 2
10 9 9 13 0 9 11 11 13 9 2
23 15 13 9 13 3 9 2 15 13 0 2 13 0 9 9 7 13 15 0 0 9 9 2
13 9 13 9 9 11 11 9 9 9 7 11 9 2
12 9 13 9 0 9 7 9 7 9 9 9 2
18 11 13 9 9 9 2 9 2 9 7 15 2 0 2 13 9 9 2
7 9 13 9 3 0 9 2
9 11 13 0 9 9 7 13 9 2
10 3 9 9 13 3 3 9 9 9 2
17 12 9 1 13 9 11 4 3 13 9 9 9 15 0 9 13 2
8 0 9 13 9 12 9 7 9
13 9 13 9 9 9 2 15 13 3 0 9 9 2
8 9 13 9 7 9 11 11 2
11 2 9 13 0 9 2 7 9 13 0 2
24 0 9 9 7 9 1 4 13 3 0 0 9 2 0 9 2 9 9 11 11 13 9 13 2
9 2 15 9 4 13 13 15 3 2
17 9 13 13 2 3 9 13 9 1 7 0 15 13 15 9 9 2
20 0 9 9 13 9 7 9 9 13 9 15 2 3 9 9 7 9 13 9 2
11 11 11 13 2 16 9 13 13 3 9 2
9 9 9 13 9 11 11 7 9 2
13 11 4 13 9 11 9 7 13 9 12 0 9 2
29 2 15 4 13 9 0 9 7 13 9 15 2 15 0 0 9 4 13 2 13 9 9 9 7 11 13 9 11 2
11 2 11 4 13 9 3 15 11 9 9 2
27 15 4 13 3 11 0 0 0 9 2 11 9 13 11 11 9 16 15 13 15 2 15 13 3 13 9 2
17 9 0 9 13 11 13 2 16 9 13 13 3 3 9 7 9 2
16 11 11 13 3 0 9 0 9 7 9 9 0 9 0 9 2
30 2 15 9 3 13 2 16 13 0 9 15 0 7 9 2 16 9 7 0 9 4 13 3 3 7 3 1 0 9 2
14 12 9 13 9 11 11 2 15 9 13 11 11 9 2
17 2 11 9 13 2 3 9 9 13 13 13 0 0 9 13 9 2
18 9 13 13 13 3 9 9 1 2 13 9 9 9 13 9 11 11 2
9 2 11 4 3 13 13 9 9 2
5 11 9 12 0 9
9 11 9 9 13 0 9 0 9 2
17 11 9 9 7 9 9 9 13 12 9 2 15 13 12 0 9 2
19 11 9 9 13 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2
11 9 7 9 9 9 9 3 13 12 9 2
8 12 9 9 12 13 11 9 2
14 15 13 11 11 2 11 11 2 11 11 7 11 11 2
12 9 13 9 9 13 3 0 9 7 15 9 2
15 9 13 0 9 9 9 7 9 13 9 3 12 9 9 2
14 9 13 9 13 9 9 7 13 13 9 13 3 9 2
10 9 9 13 9 9 7 0 0 9 2
5 11 11 11 9 9
14 11 9 0 9 11 11 4 13 11 9 9 0 9 2
25 9 9 13 9 9 9 9 13 2 16 11 4 0 9 13 11 9 0 9 0 7 0 9 9 2
14 9 13 3 9 0 0 7 3 0 9 11 9 9 2
9 11 11 13 12 1 11 11 9 2
21 11 4 3 13 3 11 9 0 9 9 12 2 12 2 3 15 13 11 9 9 2
15 15 4 13 3 11 9 9 9 9 9 7 0 9 9 2
11 11 13 0 9 1 0 0 7 0 9 2
12 15 13 3 11 9 9 2 11 2 9 9 2
15 11 9 9 9 11 11 13 9 12 1 3 0 9 1 2
12 15 1 11 4 13 9 9 1 9 0 9 2
22 11 9 9 0 9 13 11 9 9 9 2 15 3 13 11 15 13 9 11 9 9 2
10 9 9 0 9 9 13 9 11 11 2
13 11 9 9 0 9 13 9 12 11 9 9 9 2
10 9 9 13 9 13 11 9 9 9 2
4 0 9 11 9
16 11 9 9 11 9 9 13 9 12 11 9 9 12 12 9 2
20 9 13 13 0 0 9 7 9 2 15 11 9 7 9 9 3 11 9 13 2
28 2 3 13 9 13 9 9 9 2 16 3 13 9 0 7 0 9 9 3 9 2 13 9 11 11 11 9 2
27 2 13 0 2 16 11 9 4 13 1 11 9 9 7 9 7 13 9 9 2 11 9 9 11 11 13 2
11 11 9 9 9 13 9 9 7 9 9 2
16 9 13 0 9 13 9 1 2 12 9 13 12 9 9 0 2
10 9 9 13 3 12 12 9 9 9 2
5 0 9 13 3 9
10 0 9 0 9 13 9 9 9 9 2
32 2 0 9 9 4 9 3 13 9 9 2 9 7 9 9 9 1 2 9 9 13 11 11 7 11 11 11 9 9 9 13 2
16 9 13 9 3 13 9 0 9 9 2 9 7 9 0 9 2
20 16 9 13 3 9 12 2 15 13 3 13 13 0 7 15 0 9 13 9 2
17 0 9 13 9 15 9 16 9 9 2 7 0 9 9 13 0 2
7 9 4 13 0 9 1 2
8 0 9 1 0 9 13 9 2
9 15 13 13 9 0 9 7 9 2
18 3 3 0 9 13 9 2 16 9 4 3 3 13 2 15 13 9 2
22 9 13 9 7 0 9 1 0 9 11 7 11 13 0 9 9 4 3 13 13 9 2
7 9 4 3 13 13 9 2
13 15 13 0 9 9 2 0 9 7 0 0 9 2
7 9 9 13 0 7 0 2
29 15 9 13 3 9 2 15 13 0 9 9 0 9 7 9 7 9 9 2 15 4 13 3 2 3 13 3 9 2
15 15 9 13 3 9 2 16 0 9 13 13 3 9 9 2
10 9 9 13 3 3 9 7 9 9 2
18 9 13 0 2 9 1 13 2 7 3 9 9 13 0 9 13 9 2
24 11 7 11 9 13 3 3 2 16 9 3 13 15 9 2 7 9 9 9 13 3 9 15 2
22 2 9 13 3 13 3 3 9 9 13 2 16 3 0 9 13 0 9 2 9 13 2
6 3 13 9 9 1 2
17 0 9 13 13 3 2 9 2 7 13 9 0 9 7 9 9 2
4 9 9 13 0
15 11 9 9 9 13 9 11 9 1 3 9 13 9 12 2
4 9 13 9 2
11 9 9 9 13 9 11 11 11 11 9 2
11 9 9 9 3 13 8 11 11 11 9 2
6 9 13 9 11 11 2
5 9 13 0 9 2
17 9 13 16 13 3 16 9 13 0 7 13 3 16 15 13 0 2
6 2 9 13 13 13 2
6 15 4 3 13 13 2
11 0 9 13 0 0 9 2 11 11 13 2
9 9 13 2 16 9 13 0 9 2
8 2 9 9 13 3 9 0 2
23 15 1 9 9 13 3 12 9 2 15 1 13 3 12 9 9 0 8 9 2 11 13 2
11 9 13 7 15 3 13 4 13 0 9 2
7 12 9 13 0 9 9 2
19 2 11 4 13 2 16 9 12 1 12 9 11 9 4 4 13 13 9 2
32 3 11 9 13 9 3 2 16 15 3 2 15 13 9 7 13 15 9 9 2 13 3 0 9 13 3 13 9 2 11 13 2
11 0 9 13 3 16 13 13 15 13 9 2
5 9 13 3 9 2
11 2 13 9 2 15 13 3 12 0 9 2
9 3 15 4 13 0 13 0 9 2
22 13 0 2 16 15 0 13 13 15 9 2 15 4 13 0 9 9 2 13 11 11 2
19 11 1 9 9 13 13 9 9 9 2 7 3 3 13 15 15 13 13 2
6 2 9 13 3 9 2
10 15 9 13 13 13 9 7 13 15 2
14 9 9 13 12 9 0 11 9 0 9 7 9 9 2
13 9 13 11 11 11 9 7 9 11 11 11 9 2
5 9 13 11 11 2
18 15 9 9 13 2 9 9 9 9 2 11 2 11 11 11 11 2 2
11 9 4 13 9 11 11 7 9 11 11 2
5 9 9 9 11 11
14 0 9 11 4 13 9 9 9 9 2 11 11 11 2
14 15 13 11 9 9 9 7 0 9 9 7 9 9 2
11 11 11 4 13 3 9 7 9 9 9 2
16 15 13 11 9 0 9 9 9 9 7 9 9 0 9 9 2
12 11 13 3 3 9 7 0 9 9 7 9 2
18 9 13 2 16 11 11 4 13 9 11 9 0 9 9 12 13 9 2
19 15 9 9 9 9 4 13 3 9 9 11 9 0 9 13 9 12 9 2
17 11 13 9 9 9 9 7 13 3 9 15 0 9 13 0 9 2
13 12 12 9 0 9 13 12 11 9 9 9 11 2
18 0 9 11 13 9 12 9 9 9 2 15 9 13 9 9 9 9 2
19 9 13 15 0 9 3 9 9 2 9 7 9 7 9 0 9 13 9 2
8 9 13 9 13 0 9 9 2
11 2 0 9 1 9 4 13 3 9 9 2
7 9 0 9 13 0 9 2
31 9 13 3 9 13 2 3 9 4 13 2 11 9 9 11 11 13 13 0 9 9 13 2 0 9 7 9 2 9 12 2
20 9 11 11 7 11 11 13 9 2 15 9 9 0 9 13 15 13 9 9 2
17 11 9 9 9 13 9 12 11 7 11 13 9 0 9 7 9 2
16 9 1 11 7 11 13 12 0 9 13 9 13 9 0 9 2
14 2 9 13 13 3 0 9 7 13 9 3 0 9 2
14 13 3 13 0 9 7 12 9 9 2 11 11 13 2
19 9 9 13 9 9 9 2 9 9 2 9 7 9 9 9 7 9 9 2
11 11 13 2 16 9 3 3 13 9 1 2
11 2 9 7 9 13 9 3 13 9 3 2
10 9 13 2 16 13 1 12 9 9 2
8 15 4 13 13 3 9 9 2
10 9 9 4 11 7 11 1 13 3 2
18 3 9 13 15 1 3 3 15 2 16 0 9 13 9 13 9 9 2
8 2 9 13 13 0 9 9 2
10 9 11 11 13 9 3 9 0 9 2
12 2 9 9 9 13 2 16 15 13 13 3 2
9 15 9 3 9 13 9 9 3 2
10 9 7 9 4 13 9 7 0 9 2
11 3 15 4 13 0 0 9 2 11 13 2
23 12 9 0 9 9 13 9 13 9 2 9 7 9 2 15 11 9 9 9 11 11 13 2
20 11 13 9 11 9 7 9 9 2 15 13 0 9 11 11 11 2 11 2 2
13 11 13 11 2 8 8 7 0 9 9 7 9 2
16 0 9 1 0 9 13 3 0 9 11 11 7 11 11 11 2
12 2 9 13 9 0 0 9 7 0 9 9 2
19 9 9 15 13 9 3 0 9 11 11 11 2 15 9 13 3 9 9 2
13 0 9 13 11 7 11 11 11 9 2 11 13 2
3 9 13 9
11 9 13 12 0 9 9 9 9 7 9 2
16 11 11 9 11 11 13 0 9 7 15 9 11 11 13 9 2
10 9 13 3 9 9 9 7 9 9 2
18 15 1 9 9 13 0 9 9 9 7 9 13 0 13 15 9 9 2
10 9 9 9 13 3 9 9 0 9 2
7 9 13 9 0 9 1 2
6 9 9 13 3 9 2
15 9 9 9 0 9 9 13 13 13 9 1 3 0 9 2
12 9 9 11 11 7 11 11 13 0 9 9 2
29 2 9 9 13 13 0 9 2 16 3 9 4 13 2 16 13 13 9 2 13 11 11 9 11 11 7 11 11 2
15 3 3 11 9 13 2 16 9 9 13 15 15 13 13 2
13 2 13 0 2 16 13 9 9 7 15 0 9 2
12 7 15 1 3 9 7 9 15 13 0 13 2
12 3 4 13 3 9 0 9 2 13 13 15 2
18 11 9 13 3 2 16 13 9 7 13 2 9 13 9 13 13 9 2
13 2 16 9 13 2 15 1 13 9 13 0 9 2
4 11 9 13 9
9 9 11 9 13 3 12 12 9 2
8 9 13 9 3 16 0 9 2
18 9 9 0 9 13 9 15 2 16 9 13 1 0 9 11 9 13 2
8 11 9 7 11 9 13 12 2
12 2 9 13 9 0 9 9 13 12 9 1 2
10 0 2 0 0 11 9 3 13 9 2
22 3 0 13 3 15 2 16 11 9 4 9 11 9 13 13 9 2 9 11 11 13 2
16 9 13 0 9 11 9 2 9 9 2 0 9 7 0 9 2
17 2 3 0 9 4 13 9 7 9 9 3 3 9 0 9 9 2
12 9 9 15 9 13 3 2 9 11 11 13 2
12 15 11 9 9 11 9 9 13 3 12 9 2
6 9 9 13 12 9 2
9 9 11 9 13 9 12 3 12 2
15 0 9 9 9 13 9 9 7 9 9 9 1 9 9 2
5 9 13 13 0 9
15 11 11 9 4 13 11 9 13 9 9 2 9 11 11 2
14 11 9 9 13 11 11 9 11 11 0 9 9 9 2
13 9 2 9 9 2 9 9 2 13 9 9 9 2
8 11 13 9 11 9 9 9 2
15 15 13 9 9 9 0 9 13 9 2 15 13 9 9 2
10 9 3 13 9 2 15 13 15 13 2
9 13 9 13 2 15 9 13 9 2
11 9 13 13 0 2 0 7 13 0 9 2
18 9 13 2 16 9 13 2 13 2 13 9 7 13 2 15 9 13 2
12 3 9 13 2 16 9 13 7 13 15 1 2
8 9 9 13 9 9 7 9 2
15 9 13 3 2 16 0 9 13 9 2 9 7 0 9 2
21 13 9 13 2 16 9 13 13 0 9 7 16 9 13 9 9 4 13 0 9 2
13 9 13 9 13 9 13 12 9 9 9 13 9 2
8 11 11 13 11 9 9 12 2
6 11 13 9 9 9 2
11 9 13 11 9 11 11 11 9 9 9 2
4 9 13 13 9
13 11 11 9 13 9 2 9 7 9 9 13 9 2
12 2 11 11 13 15 9 0 9 15 9 11 2
15 15 4 13 0 9 3 11 9 9 9 7 13 0 9 2
12 9 9 1 15 4 13 1 3 11 9 9 2
17 15 13 9 7 0 9 0 0 9 2 13 9 13 9 11 11 2
13 13 9 9 11 2 9 0 9 13 9 11 11 2
14 15 13 13 9 7 3 9 9 2 9 7 9 11 2
25 11 13 2 16 13 0 9 0 9 4 13 0 0 9 2 0 9 7 9 7 9 9 0 9 2
14 2 0 9 7 9 0 9 13 9 0 16 15 9 2
14 11 1 9 13 9 4 13 9 2 16 9 13 13 2
10 15 13 2 16 9 0 9 13 0 2
9 11 13 3 9 13 9 9 9 2
15 2 15 13 13 0 9 7 13 0 7 0 9 9 1 2
26 11 13 9 11 11 13 3 15 9 2 15 13 2 16 9 13 11 9 9 7 9 13 13 0 0 2
21 2 11 0 9 13 2 16 1 9 13 9 2 9 7 9 13 0 13 0 0 2
3 9 9 9
10 0 9 9 9 4 13 9 9 9 2
17 9 13 0 9 1 13 0 9 2 15 4 13 9 9 9 3 2
18 9 13 9 2 15 4 13 3 0 9 13 7 3 15 13 9 9 2
11 3 4 13 0 9 3 3 13 9 1 2
8 9 9 13 11 9 9 9 2
9 2 9 13 0 9 7 9 9 2
22 9 9 4 13 9 9 0 9 7 9 1 7 13 0 9 9 2 9 11 11 13 2
11 15 9 9 0 9 4 13 0 9 9 2
20 9 13 9 9 13 9 0 9 7 15 4 3 13 2 3 0 13 13 9 2
19 13 3 9 0 9 4 3 13 3 3 9 13 9 7 15 1 0 9 2
11 3 13 9 4 13 9 7 9 13 9 2
19 15 4 13 3 9 13 9 9 2 7 13 3 2 3 3 9 13 9 2
12 9 9 13 0 7 0 2 7 9 13 0 2
6 9 13 3 0 9 2
14 3 9 4 13 9 9 9 2 16 9 13 0 9 2
24 9 13 9 9 9 7 15 4 13 13 9 2 7 7 0 9 13 9 2 7 0 9 13 2
7 9 13 13 13 9 9 2
11 9 13 0 9 2 15 9 4 13 11 2
9 9 4 13 9 7 0 15 9 2
7 9 9 13 3 0 9 2
4 9 13 9 5
5 9 9 9 13 9
11 11 9 7 0 9 9 13 9 9 9 2
9 0 9 9 13 0 9 9 9 2
13 0 2 3 0 9 9 13 0 9 9 7 9 2
8 15 9 9 13 3 0 9 2
8 2 9 4 13 15 9 3 2
44 15 4 13 0 9 13 0 0 9 9 9 2 15 4 13 0 9 7 9 2 0 9 2 9 9 9 2 9 7 9 9 7 9 9 2 13 11 9 7 0 9 9 9 2
10 9 13 9 7 9 9 0 9 9 2
13 9 13 0 9 9 9 4 13 0 9 11 9 2
27 2 9 13 3 3 3 9 9 7 0 9 9 13 9 9 7 9 2 9 11 11 11 9 9 9 13 2
38 9 13 15 9 11 9 9 7 9 9 2 11 11 11 11 11 2 11 2 2 11 9 2 11 11 11 2 11 7 9 13 9 2 3 11 7 11 2
27 2 9 9 13 0 9 11 9 0 9 7 9 2 0 9 7 9 9 13 0 9 13 9 2 11 13 2
14 9 13 9 9 11 11 9 3 9 0 9 7 9 2
12 0 9 0 9 13 3 9 9 9 11 11 2
11 11 9 9 13 9 11 9 9 9 9 2
11 9 4 13 9 13 9 7 0 9 9 2
13 9 9 13 9 13 9 9 12 13 11 0 9 2
4 9 1 12 9
12 11 9 9 7 9 13 9 13 9 9 9 2
6 9 9 9 4 13 2
12 9 13 3 9 9 2 9 2 9 7 9 2
17 9 13 9 9 0 2 0 9 2 15 13 3 0 7 0 9 2
8 9 13 3 12 9 1 11 2
25 11 9 9 7 9 13 0 0 9 9 9 13 13 9 9 7 9 7 9 9 7 0 9 1 2
7 9 7 9 13 9 9 9
6 13 9 15 16 9 2
5 13 9 15 9 2
5 15 9 9 13 2
7 9 9 9 13 9 9 2
18 9 12 9 9 9 13 9 9 9 13 9 9 7 9 9 7 9 2
18 11 9 9 11 11 13 9 2 0 13 13 9 7 9 12 9 1 2
15 9 13 9 0 9 2 11 11 9 15 9 11 9 1 2
10 9 9 13 9 9 0 9 3 9 2
18 9 13 3 9 9 13 0 9 7 9 2 9 9 7 9 9 0 2
12 3 9 13 9 13 3 9 9 9 13 9 2
13 2 9 13 13 9 13 9 2 7 9 13 3 2
7 9 13 15 9 0 9 2
19 9 13 0 9 7 9 2 3 15 13 3 0 7 0 9 2 9 13 2
7 9 9 1 0 13 9 2
21 9 13 3 9 9 2 16 9 13 2 13 9 0 9 9 7 13 9 0 9 2
8 9 9 9 9 9 13 9 2
10 0 9 9 11 11 13 9 9 9 2
15 11 13 9 9 9 0 9 2 15 3 13 9 0 9 2
7 3 9 13 9 13 9 2
26 9 9 13 0 9 2 16 11 11 13 13 9 9 9 2 0 9 0 9 7 9 3 0 13 9 2
18 9 9 13 9 9 2 16 15 9 9 9 9 13 0 9 9 9 2
11 0 9 13 9 13 9 3 3 9 9 2
32 16 9 13 9 7 9 2 13 15 9 9 9 7 9 2 15 9 11 11 13 9 9 7 9 11 11 13 9 9 7 9 2
9 9 9 9 13 3 12 0 9 2
8 9 7 9 9 13 3 3 2
12 9 12 11 9 13 9 9 4 13 0 9 2
10 9 13 9 13 0 9 9 0 9 2
3 9 9 11
22 11 9 9 13 9 12 9 0 9 12 9 0 9 13 11 11 11 9 9 9 9 2
14 9 13 11 9 9 3 0 7 3 0 9 3 0 2
19 11 9 9 9 13 9 13 2 3 9 13 9 9 7 9 13 9 9 2
9 11 11 13 9 11 9 9 9 2
9 9 4 3 9 13 9 9 9 2
12 15 13 9 13 9 9 2 16 13 9 13 2
22 2 0 2 16 15 9 4 3 13 3 0 9 2 13 9 11 11 9 7 9 9 2
21 9 0 9 9 13 11 9 9 11 11 7 11 11 9 9 9 2 15 13 9 2
5 15 13 12 9 2
14 9 11 11 7 9 9 11 11 13 9 9 9 12 2
12 9 13 3 12 9 2 12 9 7 12 9 2
6 9 9 13 0 9 2
11 9 4 13 13 9 15 3 9 9 13 2
16 9 9 9 13 13 9 2 16 9 9 4 13 12 0 9 2
8 9 13 3 12 9 12 9 2
3 15 9 11
16 2 11 13 11 9 13 3 3 0 9 2 13 11 9 11 2
20 0 12 9 11 11 9 13 11 11 13 9 11 9 0 9 11 7 15 9 2
11 9 13 7 0 9 2 9 7 11 9 2
21 7 11 9 7 11 9 13 9 11 13 2 16 11 0 9 11 13 13 0 9 2
28 9 13 9 7 9 2 7 13 2 16 0 9 7 9 9 13 3 9 13 2 16 9 9 13 3 13 9 2
12 9 0 9 7 9 9 4 3 13 9 1 2
11 9 11 1 11 13 13 0 9 13 9 2
10 2 0 9 9 13 2 3 13 9 2
8 9 13 13 15 9 0 9 2
18 9 13 3 2 16 11 13 9 1 15 9 0 0 9 9 9 9 2
10 3 9 1 11 13 13 15 9 1 2
13 15 1 11 13 9 2 15 11 13 4 13 3 2
21 9 11 13 2 16 16 11 13 3 3 0 9 9 2 13 15 3 3 0 9 2
13 11 9 9 13 13 9 9 4 11 1 13 3 2
6 2 9 9 13 9 2
14 9 13 3 9 7 9 7 9 2 15 4 13 11 2
17 11 13 9 0 9 2 15 15 4 13 2 16 9 3 13 0 2
9 3 9 13 9 2 15 13 13 2
23 11 13 9 2 16 11 9 9 13 0 0 9 2 16 0 9 11 7 11 1 13 9 2
17 11 7 11 0 9 9 11 13 9 2 15 1 9 4 13 11 2
14 9 13 0 9 11 7 11 9 1 13 15 9 0 2
12 2 15 9 4 3 13 9 9 9 0 9 2
19 11 9 13 11 9 12 9 11 9 0 9 11 11 11 11 11 11 9 2
14 11 13 9 2 16 11 9 13 0 0 0 9 9 2
21 3 9 3 9 13 0 2 16 9 13 3 11 7 11 2 13 9 7 13 9 2
3 9 13 9
19 9 9 11 11 13 9 12 0 9 13 9 11 9 9 9 9 9 9 2
16 9 9 7 0 9 13 3 0 9 7 0 9 0 0 9 2
24 9 2 9 7 9 9 2 0 9 2 13 15 1 0 13 9 7 9 9 7 9 0 9 2
9 9 13 0 9 0 9 7 9 2
16 11 1 13 3 0 13 0 9 2 15 9 13 13 15 9 2
5 9 13 12 9 2
19 3 9 4 13 0 9 7 9 0 9 2 15 13 0 9 9 7 9 2
18 0 9 4 13 0 0 9 0 9 2 15 13 0 9 9 7 9 2
22 2 15 13 3 0 9 2 15 0 9 9 13 3 9 0 9 0 9 2 13 11 2
29 2 3 9 15 9 4 13 2 16 15 9 2 0 9 2 9 7 9 2 13 9 0 7 3 15 13 4 13 2
15 0 9 13 9 7 13 7 13 13 9 15 2 11 13 2
19 0 9 4 13 0 9 0 9 2 15 13 13 0 9 9 2 3 9 2
7 15 9 13 3 0 9 2
11 9 13 4 13 9 2 16 9 13 0 2
30 9 9 13 3 13 9 2 15 0 9 13 9 12 3 3 9 7 9 2 9 2 9 7 9 2 9 7 9 9 2
9 9 13 13 3 9 2 0 9 2
6 15 13 9 0 9 2
17 2 16 13 9 9 2 4 15 9 13 3 0 9 2 11 13 2
12 0 0 9 9 9 9 4 13 9 9 9 2
22 2 3 0 9 3 9 2 9 7 9 2 15 13 11 9 2 13 3 2 11 13 2
20 11 1 4 3 13 2 16 9 13 4 13 3 9 7 16 9 13 3 9 2
5 3 15 13 9 2
26 2 0 9 1 13 9 13 3 0 2 16 3 9 4 13 3 2 8 8 8 2 9 2 11 13 2
15 11 13 2 16 9 13 13 9 7 13 3 0 0 9 2
15 9 13 3 9 11 11 2 9 11 11 7 9 11 11 2
7 9 9 13 9 11 11 2
3 9 9 0
8 9 9 13 11 9 9 9 2
14 11 9 9 9 7 9 13 11 9 9 13 0 9 2
12 9 13 9 0 9 9 13 9 9 9 9 2
9 9 9 9 4 13 0 9 9 2
14 9 0 9 9 13 3 3 0 9 9 0 16 0 2
12 9 9 9 9 13 9 9 15 3 15 0 2
14 13 9 1 9 9 4 0 9 9 13 13 9 9 2
9 9 13 9 13 3 13 0 9 2
7 9 9 9 13 9 9 2
12 3 3 0 9 13 9 13 3 0 9 9 2
12 9 13 9 4 13 9 9 3 9 13 9 2
11 0 9 9 12 9 12 13 9 13 3 2
6 9 9 13 13 9 2
10 11 9 9 13 9 9 7 9 9 2
5 0 9 9 13 11
8 11 13 15 9 3 12 9 2
13 4 13 2 16 12 9 13 11 9 9 4 13 2
22 2 3 3 13 12 12 9 9 13 11 9 0 9 12 7 9 2 13 9 11 11 2
20 11 4 13 9 12 13 9 11 9 2 9 2 9 7 9 9 2 11 2 2
11 9 9 13 11 9 11 9 7 9 9 2
14 0 9 13 11 9 0 9 7 13 9 3 3 9 2
16 2 9 9 13 3 7 9 13 13 7 13 3 2 11 13 2
17 15 13 2 16 0 9 13 9 0 9 4 13 0 9 9 9 2
12 2 3 9 9 4 13 0 9 7 9 9 2
19 11 9 13 13 13 0 9 2 3 15 2 15 9 9 13 7 15 13 2
12 0 9 7 9 9 4 13 11 0 0 9 2
24 11 13 2 16 11 4 13 13 9 9 9 9 2 16 15 13 9 11 9 9 7 9 9 2
7 2 9 9 13 13 0 2
22 3 11 13 0 9 2 15 13 3 9 13 11 9 9 2 0 9 2 0 9 2 2
18 11 9 9 13 11 11 13 2 16 0 9 13 9 7 9 0 9 2
7 2 0 13 3 9 9 2
10 3 0 9 7 9 13 9 13 11 2
13 11 11 13 9 13 9 2 15 4 13 0 9 2
20 2 11 9 11 4 13 13 9 0 9 2 11 9 11 9 7 11 9 9 2
17 16 9 13 2 15 13 0 9 3 11 9 9 9 2 11 13 2
12 11 9 4 13 9 9 11 9 7 0 9 2
26 3 13 11 9 2 9 2 9 7 9 9 9 13 9 1 0 9 3 3 9 9 2 9 7 9 2
4 9 9 0 9
33 2 9 4 13 13 3 3 9 2 9 9 2 0 9 0 9 2 9 2 9 2 9 7 9 2 13 11 11 9 9 0 9 2
26 8 11 11 13 9 2 11 11 11 11 11 11 11 11 11 11 2 13 15 2 3 0 9 13 0 2
8 0 9 13 13 3 0 13 2
13 0 9 7 9 9 13 11 1 13 9 3 0 2
11 2 9 4 13 15 0 13 0 13 9 2
15 2 9 1 9 13 3 9 3 9 1 13 2 11 13 2
24 0 9 9 7 9 13 3 15 2 16 0 9 9 4 3 13 3 3 0 2 0 7 0 2
7 2 3 9 13 9 13 2
18 3 3 15 13 13 9 13 0 9 3 16 15 9 13 2 11 13 2
13 0 9 9 13 3 0 9 7 0 9 9 15 2
6 15 13 3 9 0 2
25 11 1 0 9 0 9 1 2 15 9 4 13 9 2 15 9 13 15 9 9 7 9 13 9 2
11 0 9 13 3 0 7 13 3 0 9 2
6 13 9 0 13 9 2
14 2 0 9 4 3 13 0 2 3 0 2 13 11 2
11 2 3 0 9 9 13 9 13 13 9 2
16 0 9 13 9 3 3 9 2 9 2 9 2 9 7 9 2
3 9 7 11
10 9 11 11 13 9 9 9 11 9 2
12 9 7 9 9 11 9 13 9 7 9 11 2
29 11 2 11 11 11 2 11 11 11 11 11 2 13 11 9 2 11 11 11 11 11 2 11 11 11 11 11 2 2
23 11 3 3 13 9 9 2 15 1 15 13 0 9 7 15 9 9 9 2 11 7 9 2
7 11 13 11 9 12 9 2
27 11 9 1 9 4 13 0 9 2 3 15 13 3 3 0 7 9 13 9 2 16 13 3 13 9 9 2
24 9 0 2 7 9 9 11 13 9 7 9 11 11 2 15 0 9 15 13 13 0 9 9 2
6 9 4 3 13 9 2
7 11 1 15 9 13 0 2
17 0 9 11 13 9 2 15 13 13 9 2 7 13 3 13 9 2
17 11 13 2 16 15 9 13 15 1 2 15 13 15 0 9 11 2
16 11 13 9 13 2 13 0 0 15 0 2 15 15 9 13 2
12 0 9 7 9 13 15 2 15 13 9 13 2
9 9 9 13 9 13 9 9 11 2
12 9 13 3 3 9 9 9 2 11 7 11 2
5 9 13 0 9 9
11 11 11 13 9 9 0 9 0 9 13 2
6 3 13 3 9 9 2
24 11 11 9 11 11 13 11 13 3 9 15 2 3 13 9 13 0 9 7 9 0 0 9 2
11 11 1 9 7 9 13 13 15 9 13 2
8 15 12 9 13 9 7 9 2
11 15 13 9 9 2 0 9 7 0 9 2
10 0 9 13 3 3 15 9 9 9 2
6 15 9 13 3 9 2
26 0 9 13 3 9 2 15 4 13 0 0 9 2 13 9 9 1 3 4 13 7 9 13 9 9 2
14 11 1 9 9 4 13 3 3 9 2 9 7 9 2
20 2 0 9 4 13 0 2 16 15 4 13 9 0 9 0 9 2 13 11 2
8 9 9 9 13 9 7 9 2
16 2 9 13 3 9 7 3 9 13 15 0 9 2 11 13 2
23 9 13 15 2 16 9 13 9 3 3 16 9 13 13 15 2 16 15 13 3 0 9 2
22 11 13 13 0 0 9 3 13 0 9 2 16 9 3 13 7 9 1 13 0 9 2
11 11 3 13 9 9 7 9 9 9 0 2
7 3 15 13 9 9 1 2
25 2 9 4 13 2 16 13 2 16 9 4 13 9 9 3 3 0 16 9 9 9 2 11 13 2
4 0 9 13 9
16 9 9 11 11 7 11 11 0 9 13 9 3 9 7 9 2
11 9 7 9 9 0 9 13 9 9 3 2
8 9 0 9 4 13 11 12 2
16 9 0 0 9 9 13 12 9 9 9 9 7 15 9 9 2
12 11 9 13 9 9 13 9 9 13 0 9 2
16 0 9 9 13 9 0 9 13 9 9 9 3 9 0 9 2
21 0 9 9 13 9 11 11 13 0 9 2 3 0 0 9 13 13 13 0 9 2
26 9 1 0 9 9 9 13 13 9 9 2 9 11 11 13 2 16 9 13 3 0 9 0 0 9 2
9 2 9 13 3 9 2 11 13 2
14 9 7 9 9 9 13 9 3 12 9 13 0 9 2
21 0 9 9 13 3 9 13 9 13 3 9 3 15 2 0 9 1 9 4 13 2
20 9 9 13 2 16 7 9 0 9 13 9 7 0 9 13 13 9 0 9 2
17 15 9 9 4 0 9 13 3 9 13 9 3 3 9 0 9 2
4 11 9 9 13
18 11 0 9 13 9 0 9 3 12 9 11 11 9 9 7 0 9 2
14 11 0 9 13 9 11 9 12 9 7 12 0 9 2
8 9 9 13 3 12 12 9 2
13 9 13 9 13 9 12 9 7 0 9 12 9 2
14 11 0 9 13 9 12 13 9 9 0 9 9 11 2
19 3 9 13 11 9 9 3 3 9 7 13 9 9 9 9 7 9 1 2
18 9 9 13 9 13 9 9 9 11 11 7 9 9 9 9 11 11 2
11 11 11 9 4 13 0 9 9 9 12 2
16 9 13 3 9 3 9 9 13 9 7 3 9 13 0 9 2
3 9 9 9
13 11 9 9 9 13 9 13 9 9 9 9 1 2
12 9 9 13 12 9 11 7 11 9 1 9 2
9 9 13 2 0 9 9 13 13 2
27 2 3 13 9 13 9 15 9 2 15 15 9 13 15 9 2 9 11 11 13 13 9 13 9 0 9 2
13 0 13 3 13 2 0 9 7 15 9 9 13 2
21 9 9 13 9 9 13 15 2 16 9 13 9 2 15 13 15 0 9 7 9 2
8 9 4 13 13 13 9 9 2
15 2 9 15 13 15 2 16 9 4 13 7 13 9 3 2
11 9 4 13 9 2 15 9 15 13 13 2
19 9 9 13 13 2 7 9 4 13 15 9 2 13 9 3 13 13 9 2
12 9 13 9 13 0 2 16 9 13 15 13 2
9 9 4 13 9 9 9 7 9 2
7 2 9 13 4 13 15 2
19 15 1 9 4 13 9 13 9 7 13 15 2 16 15 9 9 13 13 2
21 9 11 11 11 9 9 9 13 9 9 2 15 13 9 9 7 9 7 9 9 2
7 2 15 9 13 3 0 2
7 3 13 3 9 9 0 2
15 3 9 13 9 3 9 0 9 2 15 13 15 9 9 2
9 0 9 4 13 3 0 9 13 2
10 2 0 9 13 9 3 9 7 12 2
9 3 3 9 13 13 9 13 0 2
7 0 9 13 9 9 9 2
4 0 9 13 11
11 11 9 0 9 4 13 0 9 9 11 2
15 9 13 11 11 7 11 11 2 3 11 11 7 11 11 2
27 11 9 9 11 11 7 0 9 9 9 11 11 7 9 11 11 13 9 12 11 9 11 13 9 13 9 2
31 9 13 0 11 7 11 11 13 9 7 9 13 11 11 9 2 15 13 9 0 9 7 9 9 11 9 7 15 0 9 2
13 9 13 11 11 9 2 3 12 9 1 11 9 2
11 9 13 3 12 9 9 7 9 7 9 2
10 0 9 13 9 0 9 0 9 9 2
6 9 9 1 13 11 2
22 9 4 13 15 9 1 0 9 0 9 7 9 2 9 3 9 7 0 9 7 9 2
8 0 9 9 11 11 13 9 2
30 2 9 13 9 7 9 0 9 0 9 9 9 2 15 4 13 0 9 9 7 9 9 7 9 9 9 2 11 13 2
4 9 9 13 9
12 9 12 13 11 11 9 13 9 9 0 9 2
7 15 9 13 11 11 9 2
20 0 9 13 11 11 9 11 9 2 11 11 7 11 9 3 12 9 13 9 2
17 11 9 9 9 13 11 11 1 9 9 4 13 9 7 9 9 2
16 2 9 9 9 13 9 9 9 7 9 9 9 2 11 13 2
6 9 13 3 9 9 2
16 2 9 9 13 3 0 2 16 15 4 13 9 2 13 11 2
10 15 3 13 9 13 2 11 11 2 2
9 15 9 13 13 0 9 9 9 2
15 9 13 9 2 15 4 13 0 9 9 7 9 9 9 2
12 9 13 9 9 2 9 7 0 9 9 9 2
17 2 9 9 4 13 9 7 9 7 13 9 9 2 13 11 11 2
14 9 13 12 9 2 15 13 0 9 1 3 0 9 2
9 9 4 13 9 1 0 9 1 2
15 11 9 9 11 11 13 9 13 3 9 9 13 1 9 2
13 2 0 9 13 3 9 11 7 11 2 11 13 2
16 9 13 15 9 3 11 11 9 2 15 4 13 3 9 9 2
12 9 13 1 12 9 2 3 3 11 7 11 2
14 9 13 11 11 11 13 9 9 7 9 7 9 9 2
26 2 15 13 13 3 9 2 7 3 13 13 9 2 16 9 13 9 1 0 9 2 13 9 11 11 2
14 0 9 9 11 11 13 11 11 13 0 9 9 1 2
10 2 9 9 13 0 9 2 11 13 2
8 9 11 13 9 3 0 9 2
2 9 13
12 11 9 12 0 9 13 9 12 0 9 11 2
32 11 9 13 12 0 9 2 9 9 2 11 11 11 11 11 2 11 2 7 9 9 2 11 11 11 11 11 11 2 11 2 2
20 0 9 13 12 9 9 13 0 9 13 9 13 9 2 9 7 9 13 9 2
31 9 0 9 9 2 11 9 9 2 9 11 11 13 2 16 16 3 9 9 13 9 13 0 9 2 15 13 3 0 9 2
9 15 13 0 9 9 0 9 9 2
17 9 13 3 11 9 9 11 11 2 15 13 9 7 9 0 9 2
17 11 11 11 9 7 9 9 13 11 0 9 13 9 9 7 9 2
12 9 11 11 11 11 11 13 9 0 9 9 2
12 11 11 11 9 13 9 9 0 9 7 9 2
11 9 0 9 9 13 9 11 11 11 9 2
10 9 9 13 11 9 2 9 11 11 2
29 9 13 9 9 1 9 11 9 7 11 9 9 9 13 11 0 9 9 2 15 13 3 0 9 2 9 7 9 2
16 9 0 9 13 9 12 7 15 9 13 12 9 9 12 9 2
12 9 9 13 9 12 0 9 1 12 0 9 2
20 9 9 11 11 2 11 2 7 11 11 2 11 2 13 9 9 13 3 3 2
19 9 0 9 2 9 11 11 13 2 16 11 9 9 4 13 9 3 3 2
29 2 9 7 9 9 13 3 0 9 9 1 2 16 15 9 13 9 2 15 15 2 7 15 9 13 2 11 13 2
19 9 9 9 13 13 3 9 7 11 13 2 13 11 0 9 9 13 9 2
30 2 0 13 9 0 9 7 9 0 9 9 2 15 13 3 3 0 9 9 7 9 7 0 0 9 9 2 11 13 2
5 9 9 9 13 3
11 9 9 9 13 9 13 0 3 3 0 2
9 11 11 13 9 9 7 9 9 2
11 11 9 13 9 9 9 13 9 9 12 2
6 11 13 9 9 12 2
9 9 9 13 11 0 9 0 9 2
5 0 13 9 9 2
18 3 3 9 9 9 9 2 9 9 7 9 9 9 13 9 13 0 2
4 9 13 3 2
10 2 3 9 13 9 9 13 11 0 2
9 9 4 13 9 13 9 9 9 2
30 9 13 2 16 0 9 13 0 9 0 2 3 9 4 3 13 7 3 0 9 3 13 9 2 9 11 11 9 13 2
11 11 13 9 9 11 9 0 9 0 9 2
15 2 11 13 0 9 2 15 13 9 0 9 9 9 9 2
17 9 13 13 9 2 7 15 9 9 9 13 3 9 2 11 13 2
11 11 11 13 9 12 11 9 0 9 9 2
15 15 13 9 9 9 9 13 15 2 15 9 13 9 9 2
10 11 11 4 13 11 9 0 9 9 2
17 2 16 9 4 13 0 9 7 15 9 4 13 2 13 9 9 2
13 9 13 9 13 3 3 0 9 2 15 13 9 2
17 11 13 0 11 9 0 9 2 15 12 9 13 3 0 9 9 2
21 2 13 0 2 16 9 13 9 3 9 9 9 9 13 9 2 3 15 9 9 2
10 11 13 2 16 9 13 9 9 9 2
17 3 3 9 9 9 9 11 9 13 4 13 9 9 9 7 9 2
10 2 3 9 13 9 3 9 16 9 2
17 9 11 11 7 11 11 11 9 0 9 4 13 9 9 9 11 2
11 9 13 9 2 15 9 9 13 15 9 2
13 2 9 13 9 0 9 9 9 7 9 9 9 2
11 9 11 13 0 0 9 9 2 11 13 2
28 0 13 15 2 16 11 9 13 3 3 7 15 4 13 0 9 15 9 16 9 9 4 3 13 3 3 13 2
18 2 3 13 0 9 13 3 9 7 15 9 3 0 3 2 11 13 2
18 11 11 2 13 12 2 13 9 7 9 9 0 13 11 9 9 9 2
16 15 4 13 9 11 9 7 11 9 7 13 9 9 9 9 2
14 11 4 13 3 9 9 9 9 2 9 7 9 9 2
16 15 4 13 9 11 2 11 7 11 7 13 9 11 9 12 2
12 11 13 15 9 2 15 4 13 9 0 0 2
17 11 2 9 11 2 13 11 9 3 12 9 1 9 13 9 11 2
14 9 13 3 12 9 2 15 0 13 11 7 11 11 2
16 11 13 3 0 2 0 9 11 11 13 3 12 9 9 1 2
5 11 9 13 0 2
9 11 13 0 9 7 0 0 9 2
13 3 11 13 0 9 2 9 2 9 7 0 9 2
10 9 9 13 3 9 7 9 7 9 2
6 9 13 9 3 0 2
5 9 13 3 0 2
9 3 15 9 13 3 9 7 9 2
19 9 4 13 3 13 2 3 11 7 11 11 4 13 9 3 3 9 9 2
7 9 13 9 3 9 1 2
12 9 9 13 2 16 9 13 13 9 9 1 2
10 3 0 9 11 13 9 13 13 9 2
8 9 11 13 3 9 7 9 2
12 3 9 13 3 3 3 3 3 9 7 9 2
5 3 9 13 11 2
5 11 13 0 9 2
14 3 13 3 0 2 0 2 0 2 0 7 0 9 2
16 9 13 0 9 3 3 9 2 9 2 9 2 9 7 9 2
15 4 13 2 16 11 9 4 13 9 1 9 7 9 9 2
9 9 9 1 9 13 9 11 9 2
13 0 9 1 15 9 11 4 13 9 0 9 9 2
21 15 13 9 0 9 2 9 9 2 9 2 9 2 9 2 9 7 9 9 9 2
9 0 9 9 13 3 11 7 11 2
44 0 9 13 3 3 11 9 2 5 12 5 12 2 2 11 2 5 12 5 12 2 2 15 9 9 12 2 11 2 5 12 5 12 2 7 11 11 2 5 12 5 12 2 2
9 15 9 13 3 11 3 13 9 2
7 0 9 13 13 3 9 2
23 15 0 9 9 4 13 0 9 2 3 11 7 11 11 2 9 3 4 3 3 3 13 2
21 0 9 1 11 9 9 9 13 13 11 11 11 3 9 2 15 9 3 15 13 2
25 0 13 0 9 9 13 9 12 2 3 11 9 13 9 9 11 11 7 15 9 11 13 3 13 2
16 0 0 9 2 11 7 11 9 0 9 2 13 3 11 9 2
15 4 13 9 2 16 3 0 9 4 15 9 13 11 12 2
9 11 9 13 3 9 9 13 9 2
17 3 9 4 13 9 7 13 9 3 1 0 9 9 7 15 1 2
16 11 13 9 11 9 13 9 9 13 3 3 9 9 11 11 2
8 0 9 11 13 13 9 1 2
9 3 9 9 13 3 9 7 9 2
5 9 9 9 13 2
11 12 7 9 13 9 3 12 0 9 9 2
12 9 9 11 9 13 9 1 9 13 12 9 2
12 9 9 1 3 13 0 9 3 11 9 9 2
12 9 11 13 2 16 11 9 13 9 9 12 2
7 3 9 13 9 13 9 2
7 11 4 13 3 0 9 2
10 3 9 9 11 13 3 11 9 9 2
26 11 13 13 9 0 9 13 9 11 9 1 3 11 2 5 12 5 12 2 2 15 13 9 7 9 2
16 0 9 13 9 11 2 5 12 5 12 2 13 3 3 9 2
10 9 2 9 11 2 13 9 13 9 2
10 15 9 9 9 13 0 9 0 9 2
13 9 0 9 13 11 2 9 13 12 7 9 12 2
12 9 13 0 15 9 2 7 15 3 13 9 2
15 9 13 3 3 0 9 2 7 15 13 3 15 9 1 2
11 9 13 3 3 0 9 9 7 9 1 2
14 13 9 3 12 9 2 9 12 5 2 15 13 13 2
15 13 9 13 3 9 2 9 2 9 7 15 15 9 1 2
13 15 13 3 3 9 1 13 9 2 9 7 9 2
7 9 13 9 12 0 9 2
9 3 9 9 13 3 15 9 3 2
29 11 2 2 11 2 2 11 11 2 13 0 9 12 11 2 11 2 11 2 13 9 7 9 7 9 0 0 9 2
8 3 15 4 13 11 11 9 2
30 11 13 3 9 7 0 9 2 7 9 2 7 4 3 13 9 7 9 2 3 11 9 11 11 7 11 9 9 2 2
23 15 9 11 13 11 0 9 7 12 9 11 2 13 12 2 7 11 2 13 12 2 1 2
9 11 4 13 11 7 11 11 11 2
24 11 11 0 9 13 9 1 13 2 7 15 1 15 13 9 0 12 9 0 9 7 9 1 2
35 15 9 13 3 11 1 13 13 2 7 13 9 3 0 7 9 11 11 2 2 0 9 2 2 2 15 1 15 15 9 13 0 16 15 2
12 9 13 15 3 9 11 2 2 9 2 2 2
31 15 9 2 7 15 16 0 11 9 9 11 13 3 2 13 3 9 9 2 7 11 1 15 9 13 3 9 7 9 9 2
12 11 13 3 13 11 7 11 13 0 9 9 2
16 3 15 0 9 13 11 11 11 2 15 9 15 4 13 9 2
11 0 15 13 9 2 11 11 2 13 9 2
8 9 15 13 0 9 11 9 2
23 15 9 15 3 13 0 9 2 11 11 2 11 11 7 11 11 7 11 0 9 2 11 2
17 9 9 13 11 11 11 16 9 13 15 9 3 15 13 9 13 2
13 9 13 0 9 7 9 16 15 9 13 0 9 2
8 9 1 11 11 11 13 11 2
17 15 0 9 11 11 13 9 7 13 2 7 13 9 9 7 9 2
10 9 12 11 7 15 0 9 13 9 2
14 11 13 1 0 9 2 7 9 13 9 0 9 9 2
26 15 13 11 9 7 9 15 4 13 11 9 2 11 2 2 2 11 11 2 2 7 2 11 11 2 2
13 13 11 9 9 7 9 9 2 15 13 11 9 2
8 15 13 3 0 9 0 9 2
13 0 9 15 3 3 13 9 11 9 7 13 15 2
24 15 9 15 3 13 11 11 2 9 15 4 9 12 13 0 9 11 9 7 9 9 9 9 2
24 11 11 4 3 13 9 2 2 11 11 11 11 2 2 2 11 2 2 13 0 9 11 1 2
9 9 12 15 13 11 0 9 9 2
14 11 11 11 3 13 12 16 15 15 9 4 13 9 2
10 15 13 9 0 9 7 13 9 11 2
7 9 13 9 13 0 9 2
11 9 13 3 0 9 9 7 15 9 1 2
9 9 0 9 13 3 11 0 9 2
12 15 1 9 13 9 7 13 0 9 7 9 2
13 9 4 3 13 9 9 2 0 9 7 9 9 2
5 9 9 13 9 2
29 3 0 9 4 15 9 9 0 9 13 0 0 9 7 13 1 0 9 2 15 13 0 0 9 2 13 3 9 2
12 0 9 4 11 11 9 1 13 0 0 9 2
9 0 9 11 9 13 3 0 11 2
22 9 13 7 13 3 0 9 15 4 3 13 0 9 13 9 2 15 3 13 0 9 2
8 11 15 9 13 11 7 11 2
7 11 0 9 13 0 11 2
20 0 7 0 13 3 11 2 11 2 11 9 2 11 2 7 15 9 3 11 2
19 9 9 9 2 9 9 9 1 12 1 9 9 13 9 4 13 9 9 2
22 9 9 7 11 9 0 9 9 11 11 1 3 13 4 13 2 16 9 13 9 9 2
18 11 0 13 3 3 0 9 2 7 0 0 9 3 0 9 13 0 2
9 3 15 9 9 13 0 9 1 2
9 9 2 9 7 9 13 0 9 2
25 11 9 4 13 9 2 9 2 9 2 9 2 9 2 9 2 0 9 2 0 9 7 0 9 2
13 11 11 13 11 13 9 2 15 13 9 9 12 2
17 11 11 9 13 11 13 0 7 9 4 13 9 9 0 9 9 2
28 12 12 9 13 11 13 9 9 0 0 2 9 13 9 2 9 7 0 9 13 4 13 2 13 3 0 9 2
17 11 11 11 2 13 0 9 12 2 11 2 13 0 9 7 9 2
10 11 13 11 7 13 9 11 7 11 2
5 3 15 13 9 2
10 9 12 15 13 9 9 7 12 9 2
6 11 4 13 3 9 2
7 15 9 9 13 11 11 2
32 11 2 9 8 2 11 2 7 9 2 9 8 2 8 8 2 13 11 13 7 11 9 7 11 9 13 0 9 9 11 9 2
11 9 13 11 9 7 11 9 0 9 9 2
7 9 4 9 13 3 11 2
23 9 9 13 0 9 11 9 7 11 0 9 2 7 9 4 13 11 9 7 9 0 9 2
11 9 13 3 12 7 15 9 13 12 9 2
19 0 9 9 13 9 2 11 2 9 8 2 7 11 2 9 8 2 1 2
10 9 0 9 2 12 9 2 13 11 2
9 3 9 13 11 11 9 11 9 2
25 11 9 9 4 13 15 9 12 2 3 9 13 9 13 13 9 0 11 9 7 9 13 13 11 2
16 0 9 1 9 13 9 1 11 9 7 13 3 11 9 9 2
18 11 1 0 9 9 9 13 9 12 2 7 9 4 13 9 11 9 2
25 16 11 13 11 11 9 12 2 11 13 11 1 9 11 15 0 9 2 15 13 11 0 9 1 2
14 0 0 9 13 2 16 9 9 13 0 9 9 9 2
29 11 9 2 3 9 11 9 2 2 0 9 11 11 11 2 13 0 0 9 2 15 13 0 9 11 11 9 12 2
14 9 13 9 11 2 15 13 11 7 9 13 9 11 2
12 9 13 0 9 11 11 9 11 11 11 11 2
17 9 9 4 3 13 3 3 11 11 2 11 11 7 11 11 11 2
7 9 0 9 9 13 11 2
10 9 0 9 13 0 11 11 9 12 2
16 3 9 4 13 3 3 11 7 11 2 11 11 7 11 11 2
21 11 2 9 1 11 7 11 11 2 3 11 2 13 15 0 9 0 9 13 9 2
13 15 9 13 9 9 2 15 13 0 0 9 9 2
6 11 13 15 0 9 2
26 2 11 11 2 15 13 9 9 9 9 1 9 9 1 11 2 11 7 3 3 11 2 11 7 11 2
15 15 13 0 0 9 2 15 9 13 0 9 7 9 9 2
27 11 9 4 13 3 0 2 0 9 7 9 9 2 7 0 9 2 0 9 2 2 9 7 9 9 9 2
13 11 9 13 3 9 9 2 9 7 9 0 9 2
13 15 13 0 0 7 9 2 15 13 3 0 9 2
19 2 0 9 9 2 15 13 9 1 9 9 0 9 11 9 7 11 9 2
8 15 13 3 9 7 0 9 2
19 2 11 9 2 15 13 11 9 9 1 9 9 9 1 11 7 11 9 2
7 15 13 3 9 0 9 2
10 11 7 11 9 15 13 3 11 9 2
8 9 13 0 0 7 0 9 2
4 9 13 0 2
18 2 11 9 2 15 13 9 9 9 11 7 11 0 7 0 9 9 2
7 15 13 9 7 13 9 2
11 2 11 9 2 15 9 9 4 13 3 2
4 2 11 9 2
13 9 13 0 9 2 15 13 3 0 9 9 9 2
15 11 2 11 2 11 7 11 2 9 11 2 13 0 9 2
19 9 13 11 9 12 9 11 11 9 11 11 11 2 3 15 13 3 9 2
7 9 12 9 13 13 9 2
9 3 9 12 9 13 12 9 9 2
15 9 12 9 11 11 13 9 9 2 3 15 9 13 0 2
6 11 11 13 9 12 2
10 9 3 15 9 9 13 11 0 9 2
5 12 9 13 9 2
5 11 13 12 9 2
11 2 11 11 11 2 12 1 11 11 11 2
7 2 11 11 11 2 9 2
7 2 11 11 11 2 9 2
12 9 13 9 13 13 9 7 13 0 9 9 2
30 0 11 9 9 12 7 0 2 11 11 2 9 13 9 7 11 13 3 3 12 12 9 3 9 13 3 12 12 9 2
11 11 4 13 3 0 9 2 3 0 9 2
16 15 9 4 13 0 9 11 11 2 11 11 7 11 11 11 2
11 9 12 13 11 0 9 9 2 11 11 2
9 15 9 13 13 9 11 11 11 2
7 11 13 9 13 11 11 2
8 3 11 4 13 3 9 9 2
18 3 15 4 13 9 9 2 15 0 12 9 9 9 4 13 11 9 2
8 12 1 11 4 13 3 9 2
10 0 11 11 13 11 11 11 9 12 2
10 0 9 9 4 3 13 9 7 9 2
10 9 9 11 13 9 9 0 9 9 2
14 9 9 4 13 9 0 9 2 11 2 11 7 9 2
17 9 9 9 4 13 11 9 7 9 15 11 9 9 3 9 1 2
25 9 13 9 12 0 9 7 0 11 9 9 11 11 2 7 0 9 11 11 2 7 9 11 11 2
9 11 11 1 13 9 13 11 11 2
8 13 9 13 5 9 11 11 2
16 11 11 9 13 11 9 7 9 1 11 9 2 12 2 9 2
10 11 13 3 9 7 13 9 11 3 2
8 11 11 13 0 11 9 9 2
6 15 13 11 9 11 2
26 15 11 9 13 11 9 0 9 2 7 3 15 9 13 11 9 2 15 11 11 9 13 3 9 0 2
14 9 13 11 11 2 0 11 2 11 9 0 9 12 2
7 11 9 13 3 9 9 2
23 11 11 2 13 0 9 12 11 2 11 2 13 0 9 2 15 13 11 9 13 11 11 2
5 15 13 9 9 2
14 9 11 11 13 13 9 9 9 11 1 0 9 12 2
11 9 12 9 13 0 9 12 9 11 1 2
12 9 12 11 13 3 9 9 12 9 11 1 2
10 11 13 0 9 9 12 9 11 11 2
12 11 11 13 3 9 2 15 13 13 15 9 2
8 12 13 9 11 13 12 9 2
6 9 12 15 13 11 2
7 11 9 13 11 13 9 2
18 15 13 9 12 9 11 9 2 7 0 9 4 13 9 9 12 9 2
9 11 9 9 13 9 12 9 11 2
9 9 12 9 13 3 12 12 9 2
7 11 9 13 12 0 9 2
18 15 13 9 7 9 2 15 15 13 11 9 2 9 9 7 9 11 2
9 9 5 5 5 13 15 9 9 2
6 15 13 9 0 9 2
22 9 4 13 0 9 0 9 2 7 13 3 3 15 13 9 13 7 9 3 13 9 2
7 9 13 15 0 13 9 2
8 0 9 11 11 13 15 9 2
21 3 9 13 13 3 9 9 2 16 9 4 13 4 13 3 9 7 13 3 3 2
19 9 0 9 5 13 3 0 9 13 9 9 7 13 3 9 0 9 3 2
29 3 9 13 9 2 15 1 9 0 9 13 3 0 9 9 9 3 2 13 0 9 9 9 5 7 9 0 9 2
26 3 9 13 9 13 9 7 13 15 5 9 2 3 3 5 2 7 13 13 9 9 7 9 3 9 2
8 9 3 13 0 13 0 9 2
24 0 9 0 9 13 15 0 13 9 2 0 0 9 2 15 13 11 11 7 11 1 11 12 2
10 0 9 13 9 13 13 12 2 5 2
15 9 13 9 13 7 3 9 13 13 5 13 9 9 9 2
6 9 13 15 12 9 2
10 9 13 3 13 9 3 3 9 9 2
21 3 9 5 5 5 5 5 5 5 5 5 7 5 13 9 0 9 7 0 9 2
33 9 5 13 3 9 9 2 16 9 13 5 2 9 13 5 2 3 9 13 7 9 2 5 5 2 7 13 13 2 5 5 2 2
10 3 15 13 9 13 0 2 7 0 2
17 15 13 3 0 9 5 5 5 2 15 13 3 3 0 11 11 2
30 5 5 5 13 11 9 2 16 9 4 13 3 3 5 7 5 5 5 5 5 5 5 5 0 5 5 5 5 12 2
14 5 13 0 9 9 9 11 11 7 11 11 0 9 2
22 3 9 9 5 2 11 9 2 7 5 2 11 9 2 13 0 2 7 13 9 9 2
27 11 9 5 13 3 0 0 9 2 15 9 13 3 9 9 9 1 2 7 3 0 9 13 0 9 3 2
10 9 13 15 9 3 0 7 0 9 2
14 16 9 3 13 5 2 9 4 13 5 13 9 9 2
9 11 11 13 3 5 0 5 5 2
16 9 4 13 9 5 3 5 2 7 9 5 4 13 0 9 2
22 0 5 13 9 2 16 9 4 13 5 15 13 5 5 5 5 7 9 13 0 9 2
9 11 9 13 3 3 9 13 9 2
6 9 13 9 13 5 2
7 9 13 15 9 12 9 2
9 5 13 9 9 7 13 9 5 2
18 5 13 9 13 5 2 15 1 9 13 13 9 9 5 5 13 9 2
14 9 4 13 15 9 2 7 15 13 3 0 7 0 2
21 9 11 9 5 5 13 5 0 2 7 15 13 0 9 2 13 9 0 9 5 2
11 0 9 13 5 2 3 9 13 12 9 2
9 5 2 15 13 11 9 7 5 2
19 9 5 5 9 4 13 5 2 11 9 2 7 5 2 11 9 2 1 2
11 0 13 3 0 9 13 5 7 9 3 2
16 11 9 9 4 3 13 9 5 2 16 9 4 13 3 5 2
26 11 11 13 3 0 9 2 0 0 9 2 15 9 13 11 9 2 0 5 5 0 5 5 0 5 2
16 3 9 4 13 9 2 7 15 13 12 9 13 0 9 3 2
9 9 13 3 0 9 9 0 9 2
8 11 9 4 13 13 5 5 2
13 11 9 9 13 5 9 13 9 5 13 11 9 2
18 11 9 5 13 9 0 9 2 9 4 13 9 13 9 5 5 5 2
10 3 9 3 13 3 5 0 5 5 2
5 15 13 0 11 2
10 5 2 13 5 5 2 4 13 9 2
8 9 4 3 3 13 13 9 2
8 11 9 5 13 3 13 3 2
10 9 9 13 0 5 5 13 3 9 2
34 15 9 9 4 13 0 9 9 9 2 5 5 5 5 5 5 5 5 5 5 5 5 5 13 0 9 5 7 9 9 9 13 0 2
29 11 9 2 5 5 5 5 5 5 2 13 15 9 11 9 1 2 7 15 4 15 9 13 13 5 5 5 5 2
12 9 9 13 0 9 5 2 7 9 13 3 2
19 11 9 2 5 5 5 5 5 5 2 13 9 5 2 7 3 3 5 2
11 9 13 0 2 7 13 3 0 9 13 2
14 13 9 11 11 1 12 9 11 13 13 0 9 9 2
17 12 11 13 9 9 2 7 13 9 2 15 13 13 9 9 3 2
19 9 13 0 9 2 3 9 4 3 13 3 2 3 15 13 0 9 2 2
21 9 13 3 15 9 0 9 13 9 2 7 15 9 1 9 4 13 9 3 3 2
12 9 13 9 3 3 0 7 3 13 11 9 2
15 11 11 11 11 11 13 9 12 13 0 9 11 0 9 2
12 15 13 9 12 11 7 13 15 9 0 9 2
10 9 13 11 2 11 7 11 9 9 2
21 9 13 0 15 13 13 13 12 0 9 13 11 11 11 2 9 13 9 0 9 2
20 9 4 13 9 9 9 9 0 9 1 3 16 0 9 11 11 11 11 11 2
19 9 9 2 11 11 2 13 15 11 9 2 15 0 9 11 11 13 13 2
8 15 1 9 13 9 11 11 2
10 9 13 11 9 9 0 9 9 12 2
8 9 13 13 3 9 12 9 2
17 11 11 2 12 2 0 9 12 2 13 0 9 7 15 9 9 2
18 0 9 11 13 13 11 9 2 15 15 13 11 11 7 15 9 9 2
17 3 15 9 13 13 2 11 9 2 2 3 15 13 9 0 9 2
10 12 9 3 9 11 0 13 9 9 2
11 13 15 9 11 9 11 11 13 9 11 2
20 3 15 9 13 0 0 9 13 9 2 15 1 15 15 13 0 9 11 9 2
21 15 9 13 3 13 9 0 2 15 1 9 9 13 11 4 13 15 9 0 9 2
14 16 9 13 13 2 11 13 11 7 0 9 13 13 2
11 9 13 15 0 2 9 7 9 9 2 2
6 9 15 13 9 11 2
20 0 9 11 13 3 9 9 11 7 11 2 16 0 9 15 13 3 13 11 2
7 9 15 13 3 1 9 2
11 11 11 13 11 11 11 11 0 7 9 2
23 0 9 4 13 11 13 2 7 11 11 1 15 9 13 11 2 15 13 3 11 11 9 2
16 11 11 13 15 9 16 0 9 11 2 0 9 9 13 9 2
15 3 3 2 11 11 11 11 4 13 15 9 1 0 9 2
26 11 11 13 9 2 11 11 2 2 9 11 11 9 2 11 11 11 11 2 7 11 9 2 11 2 2
11 9 7 9 13 0 9 11 11 0 9 2
5 15 13 9 12 2
20 11 11 2 13 0 9 12 11 2 13 0 9 12 11 2 13 9 7 9 2
20 11 9 13 9 7 9 11 11 11 7 9 9 11 11 0 9 11 11 11 2
14 15 9 13 11 11 2 9 11 11 7 9 11 11 2
13 11 11 13 3 11 11 11 1 11 0 9 12 2
15 15 13 12 9 2 11 2 11 2 11 2 11 7 11 2
9 11 13 9 9 0 0 0 9 2
10 9 9 9 9 11 13 0 9 9 2
16 9 12 11 13 9 11 11 7 11 11 1 11 13 9 9 2
7 11 13 3 9 11 9 2
9 11 11 13 9 3 9 11 1 2
15 3 2 16 11 13 0 9 11 2 15 13 3 11 9 2
7 13 15 15 13 0 9 2
18 15 1 11 13 9 2 15 13 9 7 13 9 7 9 11 11 9 2
21 15 13 13 2 13 9 13 9 7 0 9 7 9 7 0 9 9 7 9 9 2
9 15 13 9 2 0 7 13 9 2
33 3 13 9 2 15 13 3 9 9 2 13 0 9 2 15 13 13 13 9 13 9 7 9 9 3 9 2 7 9 13 3 9 2
26 0 0 9 13 15 0 2 9 9 13 3 0 9 2 9 2 1 7 9 13 9 7 2 9 2 2
29 9 13 9 9 4 13 9 7 15 9 13 9 13 0 2 15 1 3 13 3 3 0 2 3 0 9 13 3 2
39 9 9 2 16 9 13 13 7 13 9 13 3 0 2 16 9 7 3 9 13 3 9 9 13 9 2 9 2 16 9 7 9 9 13 9 4 13 9 2
8 15 9 1 13 3 13 9 2
24 9 9 13 9 13 3 13 2 7 9 13 13 9 3 2 13 9 13 9 13 9 0 9 2
14 0 9 13 9 2 15 13 9 0 7 9 13 9 2
23 0 9 13 0 2 16 15 13 9 0 2 9 9 13 9 13 0 9 1 15 9 9 2
11 9 13 9 2 15 4 13 9 9 3 2
21 0 0 9 9 9 13 15 1 13 7 13 15 9 9 2 3 9 9 0 9 2
14 0 0 0 9 9 13 3 3 9 2 9 7 9 2
20 3 0 9 13 9 7 9 2 15 9 9 4 13 9 7 0 9 7 9 2
27 0 0 9 9 4 13 9 3 0 9 2 3 9 2 2 0 9 7 0 9 2 3 0 9 9 2 2
11 11 9 13 9 13 0 9 15 16 9 2
20 9 9 13 11 9 9 7 9 13 11 11 9 9 7 11 9 9 9 9 2
8 11 13 9 13 11 9 9 2
7 9 13 11 9 9 9 2
24 11 13 0 9 9 9 11 2 9 11 7 11 2 7 3 11 9 0 9 7 9 11 9 2
9 11 13 9 1 11 9 7 9 2
9 15 1 4 13 11 11 11 9 2
19 11 11 2 13 0 9 12 2 11 2 11 2 13 0 0 9 7 9 2
8 11 13 11 9 9 9 12 2
8 15 13 11 9 9 12 9 2
10 9 2 11 11 2 13 9 13 9 2
7 9 9 13 9 13 9 2
9 9 13 0 2 9 13 0 9 2
5 9 9 13 0 2
12 9 13 3 0 2 16 9 9 13 3 0 2
17 9 13 12 9 2 9 9 12 9 7 9 12 2 12 2 9 2
17 9 2 0 2 0 2 5 2 2 15 13 9 7 9 9 13 2
13 0 0 13 9 4 13 3 12 9 12 9 0 2
7 15 13 3 11 0 9 2
7 9 13 0 9 9 9 2
15 9 13 11 11 9 7 3 11 1 11 9 3 11 1 2
12 11 9 13 9 2 9 13 3 12 12 9 2
5 3 9 13 3 2
8 15 13 3 9 9 9 1 2
11 9 13 9 4 13 3 3 11 9 1 2
9 9 7 9 7 9 7 13 9 2
7 13 9 3 3 0 9 2
13 9 13 9 9 1 9 2 3 15 9 9 9 2
15 15 4 13 9 2 9 7 9 2 7 13 9 7 9 2
6 9 13 3 9 9 2
14 9 13 12 2 3 12 9 2 15 3 13 12 9 2
5 9 4 13 3 2
4 15 13 9 2
13 9 13 9 12 9 0 2 7 9 13 3 3 2
8 9 13 9 9 2 9 9 2
9 9 13 3 9 13 2 3 9 2
9 3 9 9 9 9 13 13 9 2
10 9 4 13 3 9 7 3 15 9 2
9 11 13 0 2 11 9 13 9 2
5 9 9 15 9 2
7 9 13 3 9 7 9 2
11 15 9 13 13 2 3 9 13 9 9 2
12 9 9 13 9 9 9 9 8 15 13 9 2
10 11 13 9 3 9 7 13 9 9 2
13 9 13 3 9 13 3 9 7 3 13 3 9 2
9 3 15 13 9 13 3 15 9 2
6 9 11 13 9 9 2
20 11 13 12 9 2 15 0 13 9 2 11 11 2 7 9 2 11 11 2 2
8 9 13 3 0 11 0 9 2
25 9 2 11 11 2 13 0 9 2 15 0 9 13 9 2 11 11 2 7 9 2 11 11 2 2
9 9 2 11 11 2 13 9 12 2
11 11 9 9 12 13 11 0 9 0 9 2
19 15 13 11 9 11 11 9 11 0 9 12 3 0 9 4 13 12 9 2
10 9 13 9 0 2 0 9 13 9 2
14 9 9 13 9 9 15 15 1 9 7 9 13 9 2
50 9 9 13 2 16 9 13 9 9 0 9 2 7 15 9 13 13 2 13 3 9 13 9 9 2 7 9 13 9 7 9 1 9 13 2 3 9 12 1 9 13 15 9 15 9 16 9 15 13 2
8 9 12 9 13 9 9 9 2
9 11 13 9 11 9 11 9 11 2
7 9 9 9 12 13 12 2
6 11 9 13 12 5 2
16 11 11 0 13 0 11 11 9 2 15 13 11 11 2 11 2
11 11 9 9 3 9 13 0 7 3 0 2
18 9 13 9 9 12 7 15 13 15 0 9 11 11 7 11 11 1 2
8 9 11 13 3 0 11 1 2
18 0 11 9 13 9 13 0 8 2 13 3 0 8 16 4 4 13 2
17 11 4 13 3 9 2 15 13 13 13 11 11 11 1 11 9 2
31 9 12 13 5 9 11 11 0 9 2 15 9 9 13 12 0 11 7 15 13 0 11 9 7 0 9 7 9 16 9 2
16 15 12 0 9 13 15 9 0 9 2 15 11 4 9 13 2
9 9 12 13 11 11 9 11 9 2
13 9 13 0 12 9 11 9 7 13 9 7 9 2
13 3 13 0 9 7 9 7 9 13 11 9 3 2
34 11 11 9 13 3 3 13 3 12 0 9 2 15 13 2 11 11 2 2 9 9 9 12 11 7 2 11 11 2 9 3 9 12 2
7 0 9 13 3 3 11 2
14 9 12 13 3 11 11 0 9 11 11 9 9 12 2
25 15 9 13 15 12 0 11 9 16 5 2 7 9 13 0 2 11 11 2 7 15 13 0 9 2
9 15 9 13 3 13 12 9 9 2
29 11 11 11 2 11 7 11 2 7 11 11 11 2 11 2 13 9 11 11 9 2 15 13 11 2 11 9 12 2
8 11 9 13 0 9 2 12 2
12 15 13 9 9 1 2 15 13 12 9 9 2
12 11 7 11 9 13 0 9 2 12 1 9 2
9 15 13 9 0 9 9 11 11 2
8 2 9 13 12 9 9 1 2
26 2 11 11 11 11 2 4 13 2 11 11 11 11 2 1 7 2 11 11 2 2 11 11 2 1 2
21 2 11 11 11 11 2 13 9 11 11 11 11 9 9 2 11 11 11 11 2 2
17 2 11 11 2 9 13 9 11 11 9 2 11 11 2 11 2 2
22 2 9 0 9 13 13 9 2 7 9 13 13 0 9 9 2 3 9 13 13 9 2
16 11 11 11 2 13 0 9 12 2 11 2 13 0 0 9 2
6 9 15 13 11 9 2
10 11 13 12 9 9 11 9 11 12 2
8 12 9 9 9 15 13 12 2
29 12 9 11 13 3 9 12 2 12 9 9 12 7 12 7 9 12 7 12 7 12 9 9 12 2 12 7 12 2
18 9 11 13 9 12 9 12 7 12 7 12 9 12 2 12 7 12 2
37 11 11 13 11 11 9 0 9 12 12 9 9 9 12 2 15 13 3 11 0 0 9 11 11 9 12 1 7 3 15 13 15 9 0 0 9 2
19 12 9 11 9 13 12 2 9 12 2 7 12 9 12 2 9 12 2 2
32 9 11 11 2 11 11 2 11 11 7 11 11 13 12 12 12 9 9 0 9 12 9 12 2 15 13 15 9 0 0 9 2
27 9 11 11 2 11 11 2 11 11 7 11 11 13 0 9 12 9 12 2 15 13 15 9 9 9 12 2
13 11 11 2 13 0 9 12 11 2 13 0 9 2
7 15 9 13 0 11 11 2
16 11 13 3 11 9 2 7 4 3 13 3 11 9 9 12 2
7 9 12 11 13 11 9 2
7 11 11 13 9 0 9 2
9 15 4 13 11 12 7 12 9 2
10 11 4 13 0 9 3 12 11 9 2
11 9 9 12 7 9 12 9 3 9 12 2
7 9 11 11 13 11 9 2
16 9 2 8 8 2 13 0 9 2 15 13 11 12 9 9 2
7 9 13 11 11 11 12 2
17 0 9 9 13 0 0 7 0 9 9 2 15 13 3 9 13 2
13 15 9 13 13 9 2 16 9 13 9 7 9 2
8 9 13 0 2 16 9 13 2
12 9 13 9 0 2 9 0 7 9 9 0 2
16 9 12 9 2 9 9 3 12 9 7 9 12 2 12 9 2
13 9 13 0 11 7 11 0 9 7 11 7 11 2
22 11 0 9 4 13 11 7 11 9 2 7 9 4 0 9 13 3 7 3 13 3 2
10 3 11 9 13 3 3 11 7 11 2
14 15 9 4 13 9 9 2 9 2 9 9 7 9 2
11 9 9 9 13 12 12 2 12 12 9 2
5 9 9 13 0 2
15 0 7 0 9 13 9 2 15 13 11 9 7 11 9 2
11 9 13 12 2 3 12 9 9 13 9 2
9 9 13 3 13 9 7 9 9 2
9 9 13 12 9 2 15 9 13 2
7 9 13 3 0 9 13 2
6 9 13 3 15 9 2
9 15 9 13 9 2 15 13 0 2
7 15 13 13 12 9 0 2
14 13 0 3 3 3 0 2 7 4 3 13 3 0 2
7 11 13 11 9 9 9 2
8 9 9 13 7 9 13 3 2
21 9 13 9 9 9 7 9 13 0 9 3 9 2 9 2 9 2 9 7 9 2
11 9 2 15 13 3 9 2 13 0 9 2
12 3 9 9 13 9 9 9 13 9 7 9 2
11 9 9 13 9 9 2 9 9 13 9 2
19 3 9 9 4 13 9 2 9 9 13 9 9 2 0 9 13 1 9 2
20 9 9 13 3 9 15 1 2 0 9 9 13 7 0 9 9 13 9 9 2
11 9 9 9 9 13 9 7 9 9 9 2
9 15 9 4 13 15 15 9 9 2
20 11 11 2 13 0 9 12 2 11 2 13 0 9 2 15 13 9 12 11 2
5 11 13 3 9 2
10 11 11 13 0 9 11 9 9 12 2
16 0 11 9 13 9 13 9 11 9 1 2 15 9 13 12 2
16 15 3 11 13 9 9 12 9 9 9 2 7 9 13 13 2
15 11 13 3 3 9 9 12 2 16 9 13 3 3 12 2
12 15 9 13 12 9 13 3 13 9 9 9 2
19 9 12 11 13 3 13 13 9 13 9 2 7 11 4 13 9 0 9 2
15 11 13 12 9 12 9 2 7 13 15 9 9 0 9 2
18 9 12 13 13 11 9 0 9 2 7 3 11 13 9 13 0 9 2
11 16 11 13 3 15 9 2 13 9 12 2
21 0 9 11 13 3 9 9 2 7 11 4 13 13 9 0 9 2 11 11 9 2
14 11 13 13 9 13 13 9 2 7 0 9 13 11 2
19 11 11 13 0 9 2 7 12 9 13 12 9 9 13 0 9 13 9 2
9 9 12 13 11 11 11 0 9 2
11 11 9 13 2 7 9 13 13 11 11 2
17 9 13 3 0 9 2 16 11 13 9 11 11 7 11 11 9 2
14 9 9 13 13 0 9 2 3 1 13 3 9 9 2
9 11 13 11 11 11 1 9 12 2
19 9 13 3 13 9 2 7 9 13 11 1 13 11 11 9 13 13 11 2
27 9 13 0 2 16 9 12 11 13 3 12 9 2 7 13 3 11 9 3 0 9 11 13 3 9 0 2
14 11 13 3 13 9 2 7 0 9 13 9 0 9 2
12 12 9 12 9 13 2 7 11 13 11 9 2
15 3 11 11 4 13 9 7 13 9 11 9 9 7 9 2
17 9 12 11 13 9 9 3 12 9 2 7 3 13 11 13 9 2
18 9 12 11 13 9 3 0 2 7 11 13 3 9 0 9 12 9 2
19 3 3 11 13 9 9 12 2 16 15 9 13 3 0 9 1 3 0 2
15 11 13 9 12 9 3 12 2 7 13 15 9 9 9 2
7 11 13 3 9 9 9 2
9 9 12 11 13 3 9 12 9 2
9 11 13 11 11 9 12 13 9 2
39 9 11 11 11 7 11 11 11 11 9 13 8 9 2 7 15 1 9 4 13 3 0 9 2 15 4 13 9 15 9 2 3 8 2 9 9 7 8 2
12 11 13 3 3 0 9 9 0 9 11 1 2
20 3 12 9 9 9 9 4 13 9 3 2 13 15 9 3 0 9 4 13 2
11 11 9 4 13 3 0 9 2 11 11 2
17 11 11 2 13 0 9 12 2 11 2 11 2 13 0 0 9 2
8 11 13 11 9 3 0 9 2
21 11 13 11 0 9 7 13 9 9 9 1 2 7 3 9 12 3 11 9 9 2
32 11 3 0 0 9 13 11 9 2 16 9 13 15 9 11 9 9 12 2 11 9 9 12 7 12 7 11 9 9 9 12 2
9 15 13 3 11 15 9 0 9 2
31 11 13 11 12 9 2 13 13 3 9 9 2 16 15 13 9 13 0 9 9 2 3 11 11 2 11 11 7 11 11 2
7 11 9 9 13 0 9 2
26 9 0 0 2 12 2 3 12 9 2 15 13 13 3 0 9 2 7 13 3 0 9 7 0 9 2
17 0 9 9 9 13 0 9 15 9 2 15 9 13 3 9 9 2
19 11 13 11 0 9 3 12 9 2 12 9 2 2 15 15 13 12 9 2
13 3 15 15 9 13 0 9 9 11 1 9 12 2
17 11 13 11 13 3 0 11 7 11 9 11 2 11 7 11 11 2
12 9 1 15 4 13 11 11 7 11 11 9 2
7 11 13 3 11 11 9 2
8 9 12 13 9 9 0 9 2
9 11 13 7 9 7 0 9 9 2
7 9 13 11 7 9 11 2
9 11 11 13 9 12 9 9 9 2
11 11 13 9 0 9 2 15 11 13 1 2
25 9 9 13 15 2 16 11 9 13 15 9 3 13 11 9 2 7 9 9 15 9 13 1 9 2
11 11 11 11 11 13 11 11 9 0 9 2
6 15 13 3 9 12 2
20 9 12 9 2 11 11 2 2 2 11 11 11 2 7 2 11 2 13 9 2
16 9 13 9 0 9 12 11 7 15 13 0 9 12 12 9 2
19 9 9 3 3 2 11 11 2 13 11 0 9 7 13 3 0 9 9 2
34 11 0 2 12 2 0 9 12 2 13 11 9 7 11 9 11 0 9 7 15 9 11 11 0 0 9 7 3 9 11 11 0 9 2
11 9 9 3 11 13 9 12 13 11 9 2
11 9 12 15 13 9 11 11 9 13 9 2
19 11 0 13 9 11 9 0 9 7 13 9 15 9 11 9 1 9 12 2
19 11 13 3 11 9 11 11 7 11 11 9 11 2 7 3 11 2 1 2
5 15 13 12 9 2
23 2 11 2 12 2 2 9 11 9 11 0 1 7 0 9 11 11 11 2 11 9 1 2
20 2 11 0 2 12 2 2 13 9 9 1 2 15 13 0 9 11 9 2 2
20 11 11 2 3 11 11 11 2 13 12 2 13 0 9 2 15 13 3 11 2
6 15 4 13 11 9 2
18 11 11 9 11 11 4 13 11 11 13 2 15 0 0 9 11 2 2
8 9 12 11 13 13 3 11 2
9 11 11 4 13 9 11 7 9 2
24 9 15 4 13 3 13 9 2 2 11 9 7 11 11 11 11 9 7 11 2 11 7 11 2
15 11 11 13 0 9 11 11 0 9 2 15 13 9 12 2
15 9 11 11 13 11 11 1 9 9 7 13 11 11 9 2
10 9 12 9 13 9 11 11 13 9 2
6 11 11 13 9 9 2
13 3 11 2 3 11 11 13 9 0 9 13 9 2
9 9 9 12 13 13 9 0 9 2
15 11 11 13 3 9 9 5 12 2 11 9 13 5 12 2
14 9 2 11 11 11 2 7 2 11 11 2 13 9 2
8 11 13 9 7 0 9 11 2
11 15 13 11 9 7 4 3 13 3 11 2
12 11 13 0 9 9 7 11 13 9 9 9 2
16 9 4 13 3 12 9 9 2 15 13 3 12 12 9 9 2
16 0 11 13 9 13 11 11 2 11 11 11 7 11 11 11 2
20 11 9 13 9 0 9 11 11 11 11 9 12 2 15 13 11 9 9 12 2
6 9 9 13 9 9 2
9 9 13 9 2 16 11 13 9 2
5 15 9 9 13 2
11 3 11 13 3 9 2 9 13 3 13 2
11 11 13 12 9 0 11 9 11 2 11 2
7 9 9 13 12 12 9 2
13 15 9 13 11 11 9 2 9 9 0 9 11 2
9 0 9 9 1 13 11 7 11 2
6 9 13 0 9 11 2
10 15 0 9 13 3 0 9 9 9 2
12 11 11 13 11 11 11 13 9 13 0 9 2
18 15 13 15 9 11 11 2 11 11 11 11 11 11 11 2 12 2 2
14 11 11 13 3 0 9 16 0 9 2 3 12 9 2
7 15 3 9 4 3 13 2
15 9 4 13 3 9 2 15 13 9 15 15 9 16 9 2
15 11 11 9 0 9 13 9 3 3 11 11 7 11 11 2
21 5 7 5 2 9 7 9 2 13 0 9 13 9 13 9 7 15 3 13 9 2
19 9 13 3 9 7 9 2 2 12 9 9 5 12 9 3 12 9 2 2
41 9 4 3 13 9 1 7 9 2 9 2 7 2 15 2 7 9 13 9 7 15 9 2 3 2 12 5 12 2 13 15 16 2 12 2 7 2 12 12 2 2
26 11 2 11 11 2 13 11 11 13 9 13 0 9 0 9 2 15 13 15 9 7 13 3 9 9 2
18 15 4 3 13 0 9 13 9 2 15 13 3 3 9 7 9 9 2
14 11 9 13 3 0 15 9 16 11 13 0 0 9 2
23 11 0 9 13 2 13 15 9 4 13 9 2 3 9 2 15 9 2 3 9 2 9 2
12 11 13 9 15 9 13 13 9 3 11 0 2
5 11 13 0 9 2
15 11 13 12 9 2 9 2 9 7 9 2 11 11 2 2
10 9 13 9 2 15 13 16 11 13 2
8 11 13 15 9 13 9 9 2
8 15 9 13 3 9 13 9 11
8 9 13 13 3 9 9 9 2
10 15 9 11 13 15 13 9 13 9 2
7 9 13 13 9 9 9 2
11 15 13 9 13 9 7 9 13 13 9 2
9 11 4 13 13 9 9 2 9 2
8 2 9 9 7 13 9 9 2
10 2 9 13 9 0 0 7 0 0 2
16 2 9 0 9 2 11 11 2 2 7 2 0 0 9 2 2
14 9 4 3 3 13 9 7 3 13 2 13 7 13 2
17 2 9 9 2 15 9 4 13 9 7 13 15 3 0 9 9 2
19 2 11 4 13 0 9 2 9 4 13 0 9 7 15 9 0 9 3 2
9 2 11 13 0 9 13 9 9 2
9 2 9 2 15 4 13 9 9 2
13 2 9 9 2 15 13 9 3 9 9 9 9 2
21 3 13 3 12 9 0 9 7 9 4 3 13 15 2 7 13 15 0 9 9 2
18 2 11 13 9 11 2 11 7 11 7 15 4 3 13 13 9 11 2
10 2 2 2 13 9 1 13 9 9 3
10 2 5 2 13 9 1 13 9 9 9
9 2 2 2 2 13 9 3 13 9
8 2 5 2 13 9 1 13 9
12 2 5 2 13 9 1 13 9 7 12 0 9
8 11 11 13 11 9 9 12 2
15 15 1 11 4 13 0 9 2 15 15 13 9 9 9 2
11 9 1 11 13 0 3 9 7 9 1 2
11 9 12 11 13 9 2 15 15 13 9 2
13 15 4 13 13 11 2 7 15 13 4 13 11 2
11 11 13 9 0 13 9 7 13 13 15 2
13 3 9 13 13 13 15 15 2 15 11 13 13 2
18 3 11 13 9 7 13 13 3 0 9 2 3 9 2 11 11 2 2
9 15 13 0 9 11 0 9 12 2
8 9 13 3 3 9 11 11 2
12 15 9 13 9 13 11 3 3 11 7 11 2
8 9 1 11 13 3 3 9 2
10 11 13 11 9 2 3 13 11 11 2
8 3 0 9 13 13 0 3 2
20 15 9 11 13 11 3 0 9 7 13 15 3 9 2 15 13 15 0 9 2
14 3 15 13 11 0 9 7 15 13 3 12 0 9 2
14 11 13 3 3 11 11 9 0 9 9 9 9 12 2
18 11 2 11 2 11 2 13 0 9 12 2 13 0 9 7 0 9 2
10 9 12 1 15 4 13 11 11 9 2
7 11 13 9 11 11 9 2
20 11 13 3 13 13 9 9 7 13 9 11 11 2 15 13 0 13 9 9 2
12 9 13 11 13 9 0 0 9 1 0 9 2
16 9 9 15 13 13 1 9 12 11 11 9 3 11 11 1 2
17 9 1 9 13 11 2 15 15 11 7 11 9 3 13 3 11 2
7 9 1 11 13 3 9 2
13 9 12 9 13 12 0 9 7 11 9 9 12 2
15 11 13 9 9 9 9 12 1 7 13 0 11 11 9 2
12 9 12 11 11 13 3 9 11 13 0 9 2
17 11 0 9 11 13 9 12 9 2 15 3 11 9 11 1 13 2
12 9 12 11 13 9 11 9 3 13 9 1 2
16 0 11 11 13 11 11 9 9 9 12 1 11 13 0 9 2
27 9 12 11 9 13 11 9 9 13 0 7 9 13 0 2 16 11 9 11 13 11 3 9 12 7 12 2
9 9 12 11 13 9 11 11 9 2
21 9 13 3 3 0 2 16 11 13 9 9 12 9 9 11 13 11 0 0 9 2
15 11 13 9 9 12 16 11 1 13 11 11 13 15 9 2
8 15 13 3 13 13 9 9 2
31 11 11 2 3 11 11 11 2 0 9 12 2 11 2 11 2 0 9 12 2 11 11 2 11 2 13 0 9 7 9 2
12 13 9 9 9 11 2 11 13 9 9 12 2
26 15 13 9 16 15 9 11 11 2 15 13 9 11 11 2 13 9 2 13 9 0 9 9 9 12 2
12 11 11 13 9 12 12 9 9 12 9 9 2
16 9 15 9 13 0 2 13 4 9 13 2 13 9 3 13 2
12 11 11 13 11 2 3 0 9 0 9 2 2
18 11 12 7 11 11 13 11 9 13 0 9 2 15 9 13 12 5 2
7 9 9 11 13 12 9 2
7 9 4 13 12 9 9 2
12 15 9 9 11 13 12 9 2 12 9 2 2
4 0 9 12 2
6 9 12 5 12 5 2
10 9 12 11 9 2 9 12 11 9 2
7 9 7 0 9 12 11 2
11 9 7 0 9 13 3 12 5 11 9 2
14 9 13 11 0 2 16 15 9 5 9 12 5 12 2
20 15 13 3 3 15 1 2 16 9 13 0 2 9 12 2 12 5 12 9 2
5 9 13 9 9 2
6 11 12 13 12 9 2
15 11 11 11 13 9 12 7 0 9 15 13 0 9 9 2
13 3 9 13 9 2 9 2 9 0 9 7 9 2
10 9 12 11 11 13 13 12 0 9 2
11 12 9 3 13 3 0 9 11 11 11 2
7 15 9 13 12 11 9 2
15 11 11 11 9 13 12 11 9 7 9 9 12 11 9 2
21 11 11 11 3 1 13 9 13 9 1 2 7 15 9 13 0 2 12 11 9 2
8 15 13 3 3 16 15 9 2
20 16 9 9 13 3 0 2 13 16 9 13 3 9 2 3 15 4 13 9 2
15 9 9 2 9 2 9 7 9 9 9 13 3 3 0 2
11 9 9 11 11 11 9 13 0 9 12 2
17 9 9 13 3 12 11 9 2 15 13 15 9 0 3 13 9 2
9 11 7 11 13 9 9 11 11 2
12 15 13 11 0 0 9 2 9 3 12 9 2
7 0 9 13 9 12 9 2
12 11 13 9 11 0 9 2 9 0 9 9 2
9 15 9 13 11 11 3 13 9 2
15 9 13 0 7 9 0 2 9 0 11 9 3 12 9 2
6 9 13 9 7 9 2
26 11 1 9 13 15 9 9 13 9 2 9 2 9 7 9 2 15 13 9 2 9 2 9 7 9 2
11 9 13 0 9 0 9 9 7 9 1 2
6 15 13 3 0 9 2
7 9 13 13 3 0 9 2
6 0 9 13 0 9 2
7 15 13 3 3 12 9 2
8 11 0 9 9 9 13 9 2
8 11 9 13 3 0 9 9 2
4 9 13 0 2
12 9 9 4 13 9 2 15 13 13 15 9 2
30 0 9 11 9 1 13 0 13 9 2 13 0 9 0 9 9 7 13 9 9 9 9 9 7 9 9 1 15 9 2
18 9 13 0 9 9 2 15 1 9 0 9 7 9 4 13 11 1 2
21 3 9 0 9 13 0 9 2 15 13 13 9 2 13 9 9 2 9 7 9 2
10 15 9 4 13 9 7 9 7 9 2
6 9 9 13 9 9 2
23 16 9 4 3 9 3 13 2 4 13 9 2 16 9 13 15 9 0 9 9 12 9 2
17 0 9 1 13 11 11 9 1 3 12 12 9 9 13 0 9 2
16 11 9 13 13 3 12 12 0 9 9 7 9 13 0 9 2
10 11 7 11 9 13 3 3 13 9 2
7 9 13 11 9 9 12 2
16 9 4 13 12 9 2 12 9 9 7 0 9 12 9 9 2
16 9 11 4 13 3 12 9 2 15 13 9 12 9 9 11 2
17 9 12 11 9 13 0 7 0 9 13 9 9 7 9 12 11 2
9 3 9 13 15 9 2 13 9 2
15 9 13 3 9 12 11 9 12 9 11 11 13 9 9 2
19 11 2 11 2 11 2 13 0 9 12 11 2 13 0 9 7 9 9 2
16 11 11 13 9 9 13 11 11 7 11 11 1 9 9 12 2
18 11 13 9 2 15 13 11 1 3 11 7 11 2 9 12 9 9 2
13 11 13 11 2 15 1 15 13 9 9 11 1 2
13 15 13 9 9 9 2 13 13 13 2 9 12 2
17 15 1 15 13 9 2 3 3 13 2 7 13 11 11 11 9 2
12 15 1 11 13 12 9 7 9 7 11 1 2
12 0 9 15 13 11 11 2 9 13 12 9 2
17 15 13 3 9 9 11 2 11 7 11 2 15 11 13 11 9 2
16 9 12 11 13 9 2 15 15 9 13 9 11 7 11 11 2
8 11 13 13 2 7 13 3 2
10 9 9 1 11 4 13 9 0 9 2
5 15 13 9 9 2
19 11 4 13 11 0 9 9 7 11 2 11 2 11 7 11 9 9 12 2
20 9 12 15 13 11 11 11 11 9 3 9 12 2 3 15 13 9 9 9 2
7 15 4 13 3 11 9 2
14 15 13 9 12 9 5 9 9 9 9 0 9 1 2
5 12 13 3 0 9
4 11 13 11 9
22 11 11 11 2 0 9 12 11 2 0 9 12 11 2 13 0 2 0 11 13 9 2
10 11 13 9 9 12 7 9 9 12 2
14 1 9 15 13 9 9 11 9 7 11 0 9 9 2
10 15 13 9 9 12 11 9 0 9 2
11 15 13 9 9 9 2 0 9 7 9 2
8 11 13 9 9 9 12 9 2
30 15 13 0 9 3 11 9 9 7 9 9 2 9 9 7 9 9 2 11 11 9 7 9 9 7 9 11 9 9 2
12 9 12 9 1 15 13 3 11 9 9 9 2
10 11 11 13 3 11 11 1 9 12 2
14 15 9 13 9 2 9 11 11 11 7 11 11 11 2
10 11 13 9 9 12 11 13 11 9 2
16 9 9 13 9 2 15 0 9 2 11 11 2 1 13 9 2
8 9 15 9 13 9 11 11 2
12 11 11 4 13 2 13 7 13 9 15 9 2
8 9 2 0 9 13 9 9 2
12 9 0 9 13 13 0 11 7 9 9 9 2
24 11 11 2 11 2 0 9 13 9 13 9 2 7 13 9 0 2 15 4 13 15 0 9 2
19 9 13 0 9 9 2 3 11 11 2 11 11 2 11 11 7 11 11 2
15 9 13 15 9 11 7 9 9 1 7 3 9 9 9 2
4 9 13 15 2
5 15 9 13 9 2
6 11 13 3 9 11 2
11 11 13 11 0 9 2 12 12 9 2 2
19 9 13 0 9 0 9 2 9 8 2 9 8 2 9 8 7 9 8 2
14 11 13 12 9 9 11 9 7 12 9 9 11 9 2
10 11 13 0 9 7 13 3 0 12 2
9 9 11 13 11 9 9 9 1 2
21 16 9 13 3 11 9 2 11 13 11 9 7 13 15 9 9 2 3 9 11 2
12 11 4 3 13 11 9 7 13 0 9 9 2
8 11 13 0 9 11 13 9 2
19 9 4 13 9 12 1 7 9 12 1 9 4 13 11 3 12 12 9 2
7 9 13 12 11 0 9 2
15 9 13 11 13 0 11 9 11 11 9 13 0 9 9 2
11 9 13 0 9 9 0 9 7 0 9 2
7 9 9 13 0 0 9 2
11 0 9 9 13 3 3 9 7 0 9 2
14 11 9 13 13 9 0 9 12 3 2 12 9 3 2
7 9 13 0 9 9 12 2
17 12 9 9 13 11 11 13 11 11 2 15 4 13 9 9 1 2
17 9 13 9 7 9 2 15 9 3 12 9 13 9 7 13 9 2
15 3 12 9 1 9 3 12 9 9 13 9 13 9 13 2
28 3 9 13 9 2 15 9 3 12 9 13 9 15 9 2 7 15 13 9 15 15 0 9 3 12 9 9 2
7 11 13 11 9 13 9 2
8 11 13 11 2 9 9 9 2
24 15 13 11 2 16 11 13 9 12 3 12 0 9 11 9 11 9 2 15 15 13 9 9 2
14 15 9 0 9 4 13 9 2 3 9 4 13 3 2
10 3 9 13 2 9 13 11 9 9 2
13 9 9 13 3 12 11 2 7 3 15 13 9 2
15 9 13 13 9 2 9 11 2 3 13 2 0 2 2 2
13 0 0 9 2 15 9 4 13 2 13 9 12 2
11 9 13 11 13 9 9 9 11 7 11 2
8 0 9 11 11 13 0 9 2
9 11 13 11 9 13 9 11 11 2
18 9 9 13 3 12 5 2 9 9 12 9 7 0 9 3 12 9 2
6 9 9 13 3 0 2
7 11 13 11 11 11 1 2
6 9 9 13 12 5 2
27 3 9 13 11 9 2 7 13 9 3 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 9 2
15 11 13 9 11 11 9 13 11 2 9 9 12 5 2 2
12 11 13 11 1 11 7 3 11 9 13 11 2
12 11 13 9 11 11 2 15 9 3 13 11 2
24 15 9 13 11 11 7 11 2 3 11 9 7 9 9 2 15 0 13 11 2 11 7 11 2
35 9 11 13 11 9 13 11 2 15 9 13 11 11 2 11 11 7 11 2 3 11 9 2 11 11 7 11 9 2 3 11 7 11 11 2
7 9 11 13 11 1 11 2
15 9 11 13 11 11 9 13 11 2 9 9 12 5 2 2
21 15 13 11 11 9 1 11 2 11 7 11 2 3 11 9 13 11 9 13 11 2
12 11 13 9 11 9 9 11 2 11 7 11 2
10 9 11 2 3 11 9 11 13 11 2
20 11 9 13 11 9 13 11 9 9 2 11 2 11 2 11 2 11 7 11 2
22 11 13 3 11 9 7 11 9 3 13 11 9 2 15 9 13 11 9 3 3 9 2
14 11 9 13 9 13 9 11 9 11 0 11 9 9 2
25 15 9 3 9 0 9 13 3 3 0 9 2 15 3 13 12 13 11 2 9 0 9 11 1 2
9 0 9 1 9 11 4 13 3 2
15 11 9 9 13 9 12 2 12 7 12 7 15 13 12 2
15 3 9 13 3 9 2 12 0 9 7 9 9 13 9 2
14 9 11 11 9 9 13 9 0 9 2 15 13 12 2
7 3 9 9 13 3 9 2
7 9 13 9 11 0 9 2
14 15 13 0 9 2 9 2 9 7 9 9 9 9 2
16 0 9 9 13 9 11 11 15 13 9 12 13 9 0 9 2
8 3 9 11 11 13 9 9 2
18 0 11 9 2 9 2 13 0 9 11 11 12 9 0 9 13 9 2
24 15 13 9 9 9 11 11 11 13 9 9 2 7 11 13 2 16 9 13 3 12 9 9 2
7 13 9 7 9 13 0 2
18 9 7 9 13 0 3 3 2 9 7 9 13 9 7 9 13 9 2
16 7 13 13 0 9 2 15 13 3 12 9 13 9 9 2 2
18 9 9 3 13 0 9 12 15 9 2 16 9 9 13 13 3 3 2
8 3 15 9 9 13 9 13 2
9 9 13 4 13 0 9 7 9 2
9 9 4 9 12 1 13 9 9 2
18 0 9 4 3 13 9 15 4 9 13 9 7 15 9 3 1 9 2
18 0 9 0 9 1 4 13 2 16 9 0 9 1 0 4 3 13 2
18 11 9 9 11 11 13 9 0 2 7 13 13 9 9 3 3 0 2
7 11 11 9 13 13 9 2
22 11 11 4 13 11 9 9 2 16 9 4 3 13 15 9 2 15 9 13 0 9 2
15 9 13 0 9 13 9 2 15 13 9 0 9 13 9 2
8 3 11 9 9 13 0 9 2
18 9 9 11 11 13 2 16 12 0 9 9 13 9 4 13 0 9 2
14 9 12 11 9 9 13 0 9 3 13 9 0 9 2
18 9 4 13 9 9 9 13 2 16 9 13 13 11 9 9 13 9 2
9 0 9 9 13 9 13 3 0 2
16 9 13 11 11 1 9 13 9 13 3 12 9 9 13 9 2
17 11 11 11 2 11 2 13 0 9 12 2 13 0 0 9 9 2
4 11 13 11 2
18 13 11 11 11 11 15 13 11 9 11 11 7 13 9 12 11 9 2
11 15 13 11 9 9 12 7 13 9 9 2
10 11 9 11 11 13 11 9 9 12 2
15 0 11 13 11 9 11 9 12 7 13 9 9 9 12 2
18 15 13 3 9 9 9 9 2 12 2 7 11 9 11 2 12 2 2
13 11 13 9 12 9 9 2 7 13 9 0 9 2
9 15 13 9 12 11 11 11 11 2
8 15 0 9 13 11 11 11 2
21 11 11 11 2 0 9 12 2 11 2 12 11 2 2 13 11 9 0 9 9 2
10 15 4 13 11 2 7 13 0 9 2
8 15 13 9 9 0 9 12 2
15 9 1 15 13 0 9 2 7 15 13 9 0 9 12 2
20 0 9 15 13 9 9 2 7 9 12 15 13 9 2 7 9 12 9 9 2
22 9 9 15 13 0 0 9 9 2 7 13 3 0 9 2 0 9 7 3 0 9 2
12 0 9 9 15 13 0 11 9 0 9 9 2
8 9 15 4 9 12 13 9 2
12 15 9 13 11 2 7 13 9 11 9 1 2
10 9 1 15 13 11 9 9 9 12 2
7 15 13 9 12 0 9 2
17 11 9 2 9 2 13 9 0 0 9 2 15 13 7 13 11 2
13 11 13 11 11 9 7 11 9 11 11 13 9 2
12 15 13 3 3 0 9 2 0 11 2 9 2
14 9 9 4 13 3 2 16 15 12 9 4 13 9 2
9 11 13 12 9 11 9 11 9 2
14 15 13 3 0 9 16 0 11 2 15 11 13 13 2
7 3 11 13 15 0 3 2
13 13 2 16 11 9 11 7 11 11 13 15 9 2
29 11 0 9 13 3 15 2 13 15 13 9 0 9 13 15 2 15 13 9 13 7 9 1 2 3 16 11 13 2
15 15 1 11 13 2 16 0 9 13 0 9 7 0 9 2
15 15 4 13 2 16 15 9 13 3 0 9 16 11 9 2
27 11 2 9 11 2 13 11 9 9 12 11 13 0 0 9 2 15 9 13 3 12 0 9 9 9 1 2
12 15 9 13 15 9 2 15 13 9 9 1 2
11 9 13 3 15 15 7 15 15 1 9 2
12 9 13 9 0 0 7 0 13 0 9 1 2
9 15 13 0 9 9 0 9 12 2
13 0 9 13 13 3 13 0 9 7 0 9 1 2
25 9 9 13 9 0 9 12 12 9 1 9 13 2 16 9 4 3 13 7 13 9 12 9 1 2
10 9 9 13 2 16 15 13 0 9 2
20 9 13 15 1 2 16 11 0 13 0 9 12 0 9 11 7 11 9 1 2
10 11 2 9 11 11 2 13 9 11 2
5 15 13 11 9 2
12 11 13 0 9 11 2 11 7 11 9 1 2
5 9 9 13 11 2
16 11 9 13 12 12 9 7 9 3 12 12 12 2 12 2 2
8 11 13 0 9 9 9 9 2
8 9 13 9 13 4 13 9 2
7 9 13 11 13 0 9 2
27 15 13 12 9 9 2 3 7 3 2 7 15 9 13 12 12 9 2 9 12 2 9 13 3 12 5 2
11 9 13 11 9 2 7 15 9 13 11 2
16 9 13 11 1 11 2 11 2 11 7 11 9 7 11 11 2
7 9 12 13 9 0 9 2
5 9 13 12 9 2
10 0 9 13 9 13 9 13 11 11 2
8 11 9 4 13 11 7 11 2
16 9 13 0 2 16 9 11 2 11 11 7 11 13 9 1 2
13 9 13 11 11 2 9 11 11 7 9 11 11 2
7 9 9 13 15 9 0 2
9 11 13 11 11 7 9 13 11 2
7 9 13 11 7 11 11 2
16 11 13 9 11 13 11 11 9 9 12 2 12 2 12 2 2
7 9 13 11 9 0 9 2
11 15 13 11 11 11 7 11 11 11 11 2
7 9 9 13 11 11 11 2
15 11 11 11 2 13 11 2 13 0 11 11 9 13 9 2
19 0 9 13 11 11 9 12 13 9 9 2 15 13 3 15 9 13 9 2
32 11 11 2 13 0 9 12 2 11 2 13 11 0 9 2 15 13 9 9 0 9 9 2 11 9 9 0 9 2 9 3 2
20 9 13 9 11 0 2 0 9 2 15 13 9 11 11 7 11 11 0 9 2
22 11 13 3 0 0 9 2 3 3 11 11 11 9 2 15 4 13 9 9 9 1 2
15 9 1 3 11 11 11 4 13 15 3 3 0 0 9 2
16 9 9 11 13 9 1 9 9 7 9 0 9 13 0 9 2
14 11 9 0 9 13 11 13 9 11 7 13 0 9 2
9 9 11 13 3 9 11 2 11 2
7 11 13 15 9 13 11 2
42 11 11 2 3 11 11 11 2 13 0 9 12 11 2 11 2 13 0 9 2 9 2 9 2 13 9 7 9 2 15 13 3 13 9 11 7 11 2 7 9 9 2
20 11 13 11 2 7 13 11 2 11 11 2 15 15 13 11 11 0 11 11 2
15 11 9 11 11 13 9 7 9 11 11 9 2 7 9 2
9 11 13 11 9 11 11 9 12 2
6 11 13 11 2 11 2
18 5 11 13 0 11 13 9 9 2 15 13 9 7 13 3 15 9 2
6 9 13 9 9 9 2
6 11 13 9 9 12 2
6 9 13 9 13 9 2
8 3 0 9 9 9 13 3 2
30 9 13 0 15 9 2 9 13 3 0 9 2 15 13 0 9 0 9 9 0 9 2 3 9 13 7 13 0 9 2
24 9 13 9 3 7 9 13 3 15 1 13 0 7 3 13 9 2 15 3 13 9 4 13 2
16 15 9 13 11 12 2 15 9 2 12 9 9 7 12 11 2
21 0 9 13 0 9 2 15 13 3 12 9 0 9 2 15 9 13 9 13 9 2
16 15 0 9 13 0 9 2 9 0 9 2 3 13 0 9 2
7 9 13 9 9 13 9 2
25 15 9 13 9 11 7 11 1 3 11 9 13 11 9 9 2 9 13 11 7 11 9 15 13 2
9 9 9 13 9 2 11 1 9 2
20 9 13 0 9 2 3 9 13 13 9 9 9 3 9 2 13 13 9 13 2
10 9 9 13 15 9 9 2 9 9 2
30 3 3 9 9 13 3 2 9 13 15 9 7 9 2 16 9 13 0 9 3 0 7 3 0 9 13 0 9 1 2
8 15 9 9 4 13 9 9 2
14 3 0 11 9 9 11 13 9 9 3 3 9 9 2
28 9 9 13 15 9 2 3 9 13 13 0 9 2 15 9 13 9 1 13 9 2 9 13 9 13 9 1 2
31 3 9 13 13 9 2 15 13 3 11 9 9 13 0 0 11 9 9 13 9 9 9 2 3 9 13 9 13 3 9 2
14 9 13 9 9 13 13 0 9 9 2 9 11 11 2
28 3 13 13 3 3 9 13 9 2 15 13 3 9 9 2 3 9 11 9 11 11 4 13 0 9 9 1 2
16 9 9 9 13 13 2 16 0 0 9 13 3 3 9 1 2
18 11 11 2 13 0 9 12 11 2 13 0 0 9 2 9 7 9 2
13 15 13 9 9 11 9 12 7 9 11 9 12 2
5 15 13 11 9 2
16 11 9 12 11 13 12 9 0 2 9 0 7 12 9 12 2
21 11 13 9 12 9 9 2 11 9 12 9 9 12 7 11 11 12 9 9 12 2
8 15 13 0 9 9 12 9 2
28 9 9 11 13 9 9 3 0 7 0 9 2 16 15 9 0 9 11 11 7 11 11 13 3 0 9 9 2
7 11 13 9 9 7 9 2
11 3 15 13 9 7 9 9 7 13 9 2
8 11 13 3 3 11 9 9 2
12 0 9 13 9 7 15 13 0 9 13 9 2
14 16 9 13 9 2 15 13 15 0 9 13 9 13 2
19 15 13 3 15 15 0 0 9 13 9 9 13 0 2 15 13 3 9 2
19 11 11 2 13 0 9 12 11 2 11 9 2 11 2 13 0 0 9 2
10 15 13 0 9 12 0 9 13 9 2
11 11 4 13 9 11 2 11 7 11 9 2
11 9 12 15 13 11 11 11 11 11 9 2
19 9 9 15 4 13 0 11 12 2 11 9 12 7 12 7 11 11 12 2
25 11 12 9 13 9 13 9 12 3 3 0 11 11 0 9 13 9 2 15 15 13 9 7 9 2
16 15 13 9 13 9 3 9 9 12 1 2 7 3 0 9 2
10 9 2 11 11 2 13 9 13 9 2
27 15 13 0 9 7 11 2 11 2 11 2 11 2 11 2 11 7 11 2 7 13 3 9 12 9 9 2
13 9 9 4 13 7 9 9 7 12 9 9 9 2
6 9 13 12 9 9 2
9 9 15 13 1 0 7 1 0 2
8 9 9 7 9 13 13 3 2
13 15 13 3 0 9 7 13 15 15 9 9 9 2
8 9 13 9 9 3 3 9 2
7 9 15 4 13 0 9 2
6 9 9 13 9 0 2
18 15 9 13 9 13 9 2 15 13 15 9 2 0 9 4 13 9 2
8 9 13 3 15 9 13 9 2
8 3 9 0 9 13 9 9 2
29 11 2 11 2 11 2 0 9 12 11 2 11 2 0 9 12 11 2 11 2 13 0 9 1 13 9 7 9 2
11 11 13 3 3 11 11 7 11 11 9 2
13 9 15 13 11 11 11 11 1 7 13 9 9 2
12 15 13 3 9 7 13 9 11 11 9 1 2
28 11 2 13 2 0 9 2 2 13 0 2 3 12 9 0 11 9 15 13 11 0 9 3 12 9 9 1 2
20 15 0 9 15 13 9 12 2 13 13 0 9 2 7 9 15 13 3 9 2
21 9 13 4 13 9 2 16 15 13 3 9 0 2 7 3 3 0 13 3 13 2
6 3 9 13 13 9 2
7 15 0 9 13 3 9 2
9 15 13 15 2 16 9 13 9 2
14 11 11 2 13 0 9 12 2 11 2 13 0 9 2
22 0 11 4 13 9 9 9 2 7 9 13 9 7 11 9 2 11 11 7 11 9 2
14 11 9 11 4 13 11 9 3 2 9 12 7 12 2
22 11 11 2 13 0 9 12 11 2 11 2 13 0 9 2 15 9 13 0 0 9 2
29 11 13 11 11 11 9 9 12 7 13 15 1 12 9 2 11 11 11 7 11 2 3 16 13 9 7 13 9 2
10 11 11 13 11 11 9 11 11 9 2
14 15 4 13 9 3 11 11 9 12 13 11 11 9 2
16 9 12 15 13 11 11 11 9 2 11 11 11 2 9 9 2
9 11 9 11 11 11 13 11 12 2
10 11 13 7 13 9 15 9 3 3 2
6 15 13 3 3 9 2
15 9 13 2 11 11 11 11 2 9 11 11 11 11 9 2
23 11 13 9 3 9 9 9 9 9 7 11 2 11 11 11 11 2 2 7 0 9 9 2
9 11 11 11 13 9 12 3 11 2
18 9 0 9 2 11 2 11 11 11 2 13 3 9 0 11 11 9 2
5 9 13 3 11 2
10 9 13 0 9 11 9 9 9 12 2
17 11 11 4 13 11 3 2 9 12 11 11 7 9 12 9 11 2
10 11 0 9 2 11 2 13 9 12 2
32 11 11 2 9 8 2 8 2 2 11 2 2 11 2 11 2 11 2 11 2 13 0 9 2 15 4 13 0 0 0 9 2
17 9 0 9 13 11 11 2 9 8 2 8 2 2 11 11 2 2
16 11 9 12 13 9 11 13 9 2 15 11 9 9 13 3 2
10 11 7 11 9 13 9 1 13 11 2
12 9 13 3 0 9 1 9 9 7 9 9 2
7 0 9 9 13 0 3 2
8 9 13 11 7 9 0 9 2
12 11 13 9 2 15 13 11 9 11 9 11 2
22 9 9 13 3 12 12 2 12 2 2 7 3 13 9 12 9 11 7 12 9 11 2
9 9 7 15 9 9 11 11 11 2
13 11 2 3 11 2 13 15 0 9 9 0 9 2
13 15 13 3 3 0 2 0 2 0 7 0 9 2
22 15 13 0 9 9 7 9 2 3 0 9 9 2 9 7 9 7 3 9 7 9 2
7 9 9 13 9 13 9 2
26 9 9 9 13 9 2 7 15 13 7 9 7 9 2 9 15 9 2 16 3 9 4 13 9 9 2
16 11 4 13 3 0 9 7 9 9 2 3 0 11 11 2 2
18 9 7 0 9 13 9 2 15 1 2 0 9 2 15 9 13 9 2
15 3 9 1 9 13 0 9 9 2 3 9 13 9 1 2
9 9 9 4 3 13 3 9 9 2
17 3 9 13 3 3 9 9 13 9 0 9 2 9 2 13 9 2
6 9 9 15 13 9 2
16 9 1 13 9 4 13 9 9 9 9 7 9 13 7 3 2
10 15 3 0 0 9 13 3 9 9 2
7 0 9 9 13 9 9 2
10 11 13 0 11 11 9 12 13 9 2
5 9 13 11 0 2
7 15 13 0 9 11 9 2
4 15 13 9 2
16 9 13 9 12 1 13 11 9 2 3 11 7 11 11 11 2
12 11 11 2 13 0 9 12 2 13 0 9 2
14 11 11 13 9 11 12 9 7 0 9 12 9 9 2
9 11 11 13 9 11 9 9 9 2
9 15 13 11 9 0 7 0 9 2
14 11 11 9 13 12 9 7 9 12 12 2 12 2 2
12 9 13 11 9 11 0 0 9 12 9 11 2
9 9 4 3 13 9 0 9 1 2
22 0 9 1 2 11 13 2 9 13 3 11 11 2 15 9 15 4 13 3 9 1 2
12 0 9 9 9 13 9 9 2 9 9 9 2
19 9 12 13 11 11 1 13 11 7 11 0 9 2 15 13 3 9 9 2
17 9 9 9 4 13 2 7 3 3 9 13 13 0 9 11 9 2
15 0 9 13 0 9 1 9 0 9 2 0 9 9 2 2
6 9 13 3 12 9 2
11 2 12 2 9 11 11 13 9 9 11 2
11 2 12 2 11 11 11 11 13 11 9 2
6 9 11 0 13 9 2
10 2 12 2 9 13 11 0 9 9 2
8 9 11 13 0 7 13 11 2
9 2 12 2 0 11 9 13 11 2
21 2 12 2 9 11 11 13 15 9 0 9 3 1 15 11 9 13 7 13 9 2
13 2 12 2 0 9 2 11 9 13 9 0 9 2
19 2 12 2 9 11 11 13 9 13 2 9 1 15 9 7 13 9 2 2
11 2 12 2 9 11 0 0 9 1 13 2
15 2 12 2 0 11 11 9 2 11 11 11 2 13 9 2
14 2 12 2 11 11 7 11 11 13 11 9 11 11 2
12 9 13 9 12 9 3 13 11 11 9 3 2
10 2 12 2 9 2 11 13 3 9 2
17 2 12 2 0 9 2 0 9 11 7 0 9 11 11 13 11 2
10 2 12 2 0 9 11 11 13 9 2
15 2 12 2 11 13 9 0 0 12 9 9 2 11 12 2
20 2 12 2 9 2 9 13 12 13 9 11 1 11 11 2 12 9 13 9 2
8 2 12 2 11 0 9 13 2
13 2 12 2 11 9 11 13 0 9 13 11 3 2
8 15 13 11 9 0 0 9 2
22 2 12 2 9 13 2 16 9 12 0 0 9 9 13 11 11 9 13 3 13 9 2
7 2 12 2 11 13 9 2
11 2 12 2 11 11 13 11 0 9 9 2
19 9 7 9 2 11 2 13 9 15 13 0 9 2 15 13 13 0 9 2
21 9 13 0 9 2 15 13 13 9 0 2 3 3 9 2 9 7 9 7 9 2
12 9 0 9 13 9 9 2 9 7 9 13 2
20 16 9 13 13 2 4 9 13 7 13 2 0 9 13 3 9 1 13 9 2
10 9 13 9 9 13 7 9 3 13 2
13 11 11 2 13 0 9 12 2 13 0 0 9 2
9 9 13 11 13 11 9 12 9 2
17 9 15 13 11 11 0 0 9 9 12 7 12 7 9 9 12 2
11 3 15 13 12 9 7 13 15 12 9 2
6 9 12 15 13 9 2
10 11 9 13 11 9 9 11 9 12 2
19 9 2 8 2 8 2 2 12 2 13 15 11 12 9 9 9 13 9 2
5 15 9 13 11 2
12 9 13 11 9 13 0 9 9 11 11 9 2
16 9 12 15 13 9 11 11 2 11 9 2 7 12 9 9 2
8 9 13 9 2 11 9 2 2
19 3 15 9 11 9 4 13 12 9 9 2 3 11 11 9 7 9 2 2
13 9 12 11 11 13 9 11 11 2 11 9 2 2
18 11 11 13 12 7 15 9 11 11 13 11 9 9 7 9 0 9 2
35 15 9 11 11 13 0 9 15 7 13 13 9 2 7 11 2 11 2 9 11 11 13 3 15 9 9 7 9 11 11 13 3 9 12 2
6 11 13 11 11 12 2
17 3 3 9 12 11 11 2 11 0 9 2 13 9 7 13 9 2
18 11 2 11 5 11 13 0 11 11 9 11 9 2 15 13 9 12 2
9 15 13 0 9 9 11 13 9 2
13 9 12 2 9 12 2 9 12 13 3 0 9 2
9 9 13 9 9 11 9 9 12 2
45 0 9 11 2 11 5 11 13 2 11 11 11 11 11 11 2 7 2 2 11 11 11 2 11 11 2 2 15 9 13 3 9 12 11 11 9 1 0 2 0 2 0 11 11 2
11 9 9 13 11 11 15 3 13 15 9 2
12 9 13 3 9 2 15 13 15 3 9 11 2
13 3 15 11 9 9 3 13 9 4 13 7 13 2
19 2 11 2 9 13 3 0 2 0 9 11 11 9 13 0 9 11 11 2
9 9 13 9 9 9 9 13 9 2
7 9 15 4 13 9 9 2
17 9 4 13 9 3 9 2 3 16 15 13 9 9 7 9 9 2
27 9 13 9 9 3 15 9 9 2 3 0 9 9 0 9 13 9 13 9 2 9 3 4 13 9 9 2
22 3 3 3 9 7 9 9 2 2 9 9 2 2 13 9 2 3 15 9 13 9 2
15 9 9 13 2 13 7 13 9 7 13 9 1 9 9 2
22 9 13 13 0 13 3 3 2 15 9 13 7 15 9 13 9 7 15 9 9 9 2
9 9 9 7 9 13 13 0 9 2
18 0 9 7 9 1 9 13 0 9 2 9 4 13 3 9 9 1 2
12 0 13 16 9 13 15 3 9 9 13 9 2
24 0 9 1 9 13 3 9 2 16 13 13 0 9 7 0 9 0 7 3 13 9 0 9 2
10 9 13 3 13 9 9 0 0 9 2
12 16 9 13 9 1 13 9 3 13 0 9 2
18 3 9 13 0 9 2 16 3 13 9 9 4 13 0 7 0 9 2
13 9 13 4 13 0 9 9 13 9 9 7 9 2
26 9 13 9 3 2 13 15 13 0 2 3 0 7 9 0 2 13 9 7 16 15 13 9 11 9 2
13 9 1 9 13 9 0 9 9 9 7 9 3 2
15 3 15 13 2 16 9 13 0 7 9 4 0 9 13 2
17 9 9 4 3 13 9 0 9 13 2 7 9 7 9 3 13 2
15 9 13 9 13 9 7 9 2 9 9 2 0 9 3 2
16 9 9 13 13 9 2 7 9 7 3 3 9 4 13 3 2
8 9 7 9 13 3 9 9 2
16 9 1 13 13 0 9 9 15 13 9 15 15 9 9 13 2
19 9 9 7 3 9 13 9 1 9 9 2 9 2 9 7 0 9 1 2
9 9 9 9 13 9 15 13 9 2
9 9 13 9 1 0 9 0 9 2
12 13 9 0 9 4 13 11 9 13 9 3 2
9 13 9 9 4 13 11 9 9 2
15 9 9 13 9 2 9 13 9 9 13 7 13 3 15 2
21 16 15 9 13 3 13 9 3 2 9 13 3 3 0 9 3 9 9 11 11 2
10 9 13 2 0 0 9 9 4 13 2
13 9 13 9 9 4 13 13 0 16 15 9 13 2
12 9 9 13 0 9 9 7 13 9 3 9 2
7 9 9 13 9 0 9 2
22 9 9 13 9 13 9 13 0 9 9 7 9 3 15 9 13 7 0 9 9 9 2
5 9 9 12 9 2
7 9 13 13 9 13 9 2
7 9 13 9 13 9 9 2
5 9 9 12 9 2
13 9 13 3 12 9 9 7 12 9 0 9 9 2
11 9 13 9 9 7 3 9 7 0 9 2
9 9 13 9 13 9 7 9 9 2
14 13 3 0 9 7 13 13 3 15 11 2 9 9 2
10 3 15 12 15 3 0 9 13 3 2
4 9 9 12 9
15 9 13 3 12 9 0 9 7 12 9 0 13 9 9 2
11 9 9 13 9 7 3 9 7 0 9 2
18 9 13 9 13 0 9 7 9 9 7 13 9 9 2 9 7 9 2
10 11 9 9 12 9 13 11 9 9 2
9 9 13 3 3 0 0 9 9 2
21 3 0 9 9 9 4 13 3 9 9 7 3 13 7 13 3 13 9 7 9 2
12 3 9 9 9 7 9 13 9 13 0 9 2
14 11 13 9 9 0 9 2 15 9 4 13 9 9 2
17 9 13 3 9 2 7 15 4 13 3 13 9 7 13 0 9 2
9 0 13 9 13 3 12 12 9 2
13 11 13 0 9 9 13 0 11 11 9 0 9 2
6 15 13 9 11 9 2
8 9 9 13 9 3 11 11 2
8 11 13 0 9 1 11 9 2
10 12 11 9 13 0 9 9 9 13 2
6 0 0 9 13 12 2
7 12 11 13 11 9 9 2
16 9 13 3 13 9 2 16 15 13 13 13 9 0 9 9 2
6 11 13 3 9 9 2
12 11 4 13 11 2 11 2 11 7 11 1 2
10 9 9 11 13 9 0 9 9 9 2
17 11 0 9 13 12 9 2 11 9 13 11 7 9 9 13 11 2
5 9 9 13 11 2
11 0 9 13 11 13 13 9 0 9 11 2
7 9 9 13 3 0 9 2
29 9 9 13 11 2 15 0 9 13 11 2 11 2 11 2 0 11 2 11 2 9 11 2 0 11 7 9 11 2
18 11 13 9 2 15 13 2 0 9 2 3 9 7 3 0 9 2 2
19 9 13 15 11 13 2 7 9 12 1 9 13 9 13 9 7 13 9 2
8 9 13 0 9 11 11 9 2
15 15 0 9 13 0 9 2 0 9 7 0 0 11 9 2
8 11 0 9 13 11 0 9 2
19 9 7 9 2 9 8 2 13 11 2 3 11 2 7 0 11 9 9 2
10 9 9 13 3 11 9 7 3 9 2
9 9 13 3 0 9 7 9 9 2
17 9 13 9 3 9 12 7 13 11 7 9 11 9 13 13 0 2
30 16 9 13 11 9 3 9 12 2 9 13 12 0 9 13 7 0 9 7 0 9 7 0 9 9 3 9 9 1 2
7 3 0 9 13 15 1 2
30 0 0 9 1 0 9 11 0 2 13 12 2 13 11 9 15 9 2 15 9 13 9 2 11 2 2 11 0 9 2
14 11 13 3 0 9 2 9 0 9 11 0 9 1 2
19 11 9 13 9 13 11 2 3 4 13 2 16 0 9 4 13 9 9 2
8 9 0 9 13 3 3 13 2
36 11 9 13 13 9 11 2 11 2 3 3 3 15 3 3 2 3 0 9 4 7 13 11 9 9 7 9 2 11 2 13 0 9 13 9 2
12 9 11 11 4 13 2 16 9 13 9 9 2
12 15 13 15 11 12 0 9 7 0 9 9 2
31 9 12 15 9 13 3 11 7 11 9 2 15 13 12 11 9 9 2 15 12 9 2 9 2 9 7 9 2 13 3 2
31 0 9 11 11 4 3 13 9 0 9 7 13 15 0 9 2 15 13 15 0 0 9 2 15 13 13 0 9 3 0 2
18 15 9 0 9 4 4 13 11 9 2 16 15 13 11 9 9 9 2
17 9 9 11 9 13 9 15 2 16 9 4 13 11 9 9 9 2
11 9 0 9 13 13 7 0 9 3 13 2
17 9 9 11 0 2 13 12 2 13 11 9 9 9 11 9 1 2
19 11 9 9 12 11 9 11 3 13 2 7 11 13 15 1 11 11 9 2
12 11 13 3 13 0 9 7 13 0 9 11 2
22 9 13 3 2 16 0 9 11 13 11 2 15 9 11 7 15 9 9 9 12 1 2
20 9 3 13 3 11 1 9 11 2 7 13 3 13 11 11 13 9 11 0 2
10 15 1 13 11 13 11 0 9 12 2
30 11 9 11 13 9 9 7 13 11 9 9 12 2 7 11 9 7 9 11 0 2 13 12 2 13 13 13 9 9 2
25 9 12 1 9 4 3 3 13 11 9 13 9 11 0 9 2 13 12 2 7 13 13 11 9 2
14 9 3 13 13 11 11 1 13 11 9 1 9 12 2
14 0 9 7 9 9 13 11 9 9 7 9 9 11 2
19 0 9 3 13 9 13 0 9 2 15 13 0 0 9 9 9 9 9 2
34 16 11 9 13 9 2 15 13 3 3 0 0 9 2 16 11 0 11 2 13 12 2 13 9 9 12 7 13 9 7 9 1 11 2
18 15 13 3 3 0 11 9 7 15 4 3 13 11 0 9 11 9 2
24 15 13 0 9 11 0 11 1 0 9 9 1 7 13 0 2 3 0 13 9 9 9 1 2
16 11 0 9 1 9 12 9 13 7 15 13 11 3 3 9 2
10 9 13 9 0 9 11 0 9 9 2
16 16 9 11 0 13 9 12 2 9 13 9 3 7 13 9 2
8 11 9 13 3 13 15 9 2
18 11 0 9 13 13 9 2 0 9 11 9 7 0 9 11 7 11 2
29 0 9 9 11 0 2 13 12 2 13 9 12 9 1 7 13 9 11 9 11 2 15 1 15 13 0 0 9 2
8 15 13 13 11 9 9 9 2
17 11 13 9 9 12 9 2 15 11 13 11 7 11 1 3 11 2
19 11 9 7 9 11 0 2 13 12 2 13 3 13 9 7 13 11 3 2
23 11 9 11 2 13 12 2 13 3 0 9 9 9 1 7 13 11 0 9 1 9 12 2
21 11 0 13 13 11 0 7 13 15 9 11 13 9 11 11 0 2 13 12 2 2
32 16 9 4 3 13 9 11 9 2 9 13 11 13 9 2 7 11 0 2 13 12 2 3 12 2 13 9 13 9 9 9 2
8 9 13 3 3 0 0 9 2
43 11 0 2 13 3 12 2 9 1 0 9 7 11 0 2 13 12 2 3 12 2 13 9 2 7 0 9 13 3 9 11 2 15 9 13 0 9 2 11 9 9 11 2
8 15 13 9 9 9 9 12 2
23 16 11 13 2 15 0 9 11 2 13 3 12 2 13 11 13 9 11 2 11 2 11 2
25 15 0 9 11 2 13 12 2 3 12 2 3 13 11 7 13 3 9 9 9 11 9 11 1 2
14 9 13 12 9 0 16 0 9 2 15 13 9 12 2
9 16 11 13 9 12 2 15 13 2
20 0 9 13 1 9 9 11 7 13 9 2 8 2 9 2 15 13 9 1 2
7 9 9 13 15 9 9 2
29 11 0 11 11 2 9 8 8 8 2 12 9 2 12 9 2 3 11 11 2 13 11 9 12 9 2 12 9 2
8 15 9 13 9 11 0 11 2
14 11 13 11 0 9 7 11 9 0 9 0 9 9 2
16 11 13 9 1 11 9 2 7 15 13 3 9 11 9 1 2
28 0 9 2 12 9 2 12 9 2 15 13 0 9 11 7 11 9 13 9 2 3 15 13 13 12 12 9 2
20 11 13 3 11 2 7 9 11 13 15 9 9 12 9 7 11 4 13 9 2
13 0 9 2 12 9 2 12 9 2 13 0 9 2
18 0 9 2 12 9 2 12 9 2 0 9 11 7 11 13 11 3 2
11 11 13 7 13 15 13 9 11 0 13 2
8 11 13 11 2 11 9 9 2
19 15 9 13 9 11 0 11 7 9 9 11 2 15 13 3 11 0 9 2
13 11 0 13 11 9 0 9 7 13 9 9 11 2
12 3 11 7 11 13 11 9 1 11 0 9 2
14 9 12 9 7 12 9 11 0 13 9 9 9 11 2
17 11 13 15 1 11 0 9 11 0 9 11 11 7 11 11 9 2
17 11 11 2 15 13 9 11 0 2 13 0 7 9 9 3 0 2
13 3 13 3 0 2 16 11 13 0 9 11 11 2
8 11 9 9 11 13 11 11 2
5 11 13 3 9 2
27 15 2 3 3 13 9 1 11 13 9 0 11 7 11 11 9 2 15 15 13 9 7 13 9 9 1 2
10 11 13 3 13 9 9 15 9 9 2
14 0 9 11 13 13 12 2 0 7 3 12 0 9 2
6 9 13 13 12 9 2
14 3 9 12 11 13 11 2 13 9 7 13 9 11 2
17 15 9 11 11 13 3 13 9 2 7 15 9 1 11 13 15 2
9 13 9 11 13 13 9 11 9 2
7 3 15 13 11 11 9 2
9 15 9 15 13 3 9 0 11 2
24 3 9 12 9 7 12 9 1 11 13 9 11 11 2 15 0 9 13 9 9 7 11 1 2
15 11 13 9 12 9 9 11 9 7 3 3 12 15 9 2
13 9 13 0 9 1 2 7 11 13 0 11 9 2
12 3 11 9 13 11 7 11 13 9 11 9 2
8 9 13 11 9 13 11 9 2
18 3 11 0 9 7 3 0 0 11 9 7 11 11 13 11 9 1 2
7 15 1 13 11 11 9 2
6 11 13 11 9 9 2
11 15 9 13 0 9 15 9 3 13 9 2
17 9 13 3 3 11 9 13 11 9 9 7 9 3 15 0 9 2
21 11 13 9 12 9 1 11 7 11 2 7 15 4 13 3 11 7 11 9 9 2
17 9 12 7 12 1 11 13 0 9 7 9 9 7 0 9 9 2
13 15 13 11 9 7 9 11 11 7 9 11 9 2
20 11 9 9 13 0 9 11 11 7 11 2 16 15 13 3 13 11 9 9 2
8 11 4 3 13 9 11 1 2
18 9 13 3 13 3 0 11 9 2 16 15 13 3 11 9 7 9 2
14 3 9 12 9 11 13 13 3 9 11 7 11 9 2
19 9 12 9 11 7 15 9 11 9 11 0 11 13 11 7 13 9 3 2
22 3 9 13 4 13 11 9 2 7 3 15 13 11 1 9 2 15 13 9 13 9 2
13 11 13 13 9 9 2 15 15 13 9 13 0 2
16 15 1 11 13 3 9 11 2 15 3 15 9 4 4 13 2
8 11 13 3 0 9 11 9 2
23 11 9 4 13 9 11 11 9 11 0 9 2 7 11 15 4 3 3 13 11 0 9 2
17 11 13 3 9 12 9 9 12 9 2 3 15 13 0 9 11 2
7 11 13 13 15 9 1 2
19 11 9 11 13 11 9 2 16 15 7 11 12 9 13 3 3 0 13 2
23 11 9 13 3 12 9 2 16 9 12 9 11 9 11 13 11 7 13 11 13 3 3 2
19 11 13 15 3 2 15 13 11 9 9 9 7 13 9 11 0 11 9 2
15 3 3 13 2 16 11 4 13 11 11 13 3 0 9 2
13 13 13 15 11 13 9 9 7 9 9 13 9 2
13 11 13 13 11 12 12 9 7 12 12 9 9 2
7 3 15 4 13 12 9 2
6 9 13 3 3 13 2
12 11 13 4 13 2 16 11 0 13 9 9 2
22 11 13 9 11 0 11 9 2 7 11 13 11 0 9 2 16 0 9 13 3 0 2
8 15 9 13 3 12 9 9 2
22 3 15 9 9 1 11 9 13 11 2 7 15 13 13 13 9 13 11 7 11 9 2
17 3 11 7 11 4 13 13 11 9 15 2 16 15 13 11 9 2
17 9 11 11 13 3 11 9 7 13 11 9 12 9 7 12 9 2
16 15 13 13 11 2 16 15 13 7 13 9 0 7 13 15 2
26 3 9 12 9 11 9 13 9 11 0 9 1 7 13 0 9 9 2 15 13 13 11 2 13 9 2
8 11 13 3 7 13 9 11 2
26 16 15 13 2 11 9 11 13 3 9 7 13 13 15 9 2 15 15 13 13 9 11 0 0 9 2
16 11 13 11 7 9 11 13 2 16 11 0 4 13 9 0 2
17 11 13 3 11 11 7 13 2 16 15 13 0 9 11 0 9 2
23 9 13 13 13 9 15 3 2 7 13 11 13 11 7 2 3 3 2 3 11 13 11 2
6 15 9 13 3 0 2
14 11 13 11 2 7 9 9 13 15 0 9 2 11 2
17 0 9 2 11 11 2 13 0 0 9 11 11 13 11 11 9 2
19 0 9 13 13 3 12 9 9 2 7 15 13 9 9 2 15 13 9 2
6 9 13 13 0 9 2
22 9 13 3 15 12 9 2 9 7 9 2 15 13 9 13 9 2 9 3 13 9 2
8 9 9 15 13 9 0 9 2
22 15 3 13 3 0 9 9 11 2 7 9 11 11 2 15 9 9 2 3 9 11 2
31 9 13 3 9 3 0 2 16 9 1 9 13 13 13 3 15 2 7 3 9 9 9 13 9 7 13 15 3 3 9 2
16 0 9 13 3 9 0 9 11 2 15 13 9 9 11 11 2
12 9 15 13 9 9 2 7 3 13 9 9 2
18 11 11 13 9 11 11 9 0 9 2 7 15 13 0 9 11 11 2
8 3 15 13 9 7 13 9 2
7 3 15 9 13 7 13 2
5 9 13 0 9 2
12 0 9 0 9 13 9 15 13 9 9 1 2
9 9 9 13 13 0 9 3 9 2
18 0 9 0 13 11 12 9 11 9 1 2 3 12 9 9 9 2 2
14 0 9 9 13 3 11 11 1 12 9 11 9 1 2
12 11 13 9 2 15 13 0 9 7 11 0 9
38 9 9 13 12 9 2 11 11 9 0 2 0 9 2 11 11 9 0 2 9 9 7 11 11 9 0 2 11 9 2 7 15 11 11 9 7 9 2
10 11 13 11 0 9 11 9 11 1 2
14 3 13 0 9 2 15 1 9 11 9 13 9 9 2
17 11 13 4 13 9 2 16 11 9 11 4 9 13 12 7 9 2
15 11 9 15 1 13 11 0 11 9 13 11 9 0 9 2
27 11 11 9 2 11 9 7 9 2 0 9 12 2 0 9 12 2 2 13 11 9 9 11 11 9 9 2
34 11 2 11 11 11 11 11 2 11 11 11 11 11 2 13 11 9 7 0 9 11 11 7 15 9 11 2 3 9 11 2 0 9 2
25 9 1 15 13 11 9 7 0 9 12 9 11 11 13 0 9 15 11 0 9 2 11 9 9 2
10 15 9 15 13 0 9 2 3 9 2
12 9 11 13 11 0 9 9 7 13 3 9 2
14 15 1 15 13 11 9 9 7 13 3 0 9 9 2
5 9 13 9 12 2
15 0 9 13 7 3 3 13 2 11 13 9 0 9 12 2
13 9 7 15 13 12 9 9 9 15 13 9 9 2
11 9 7 9 9 9 11 13 3 13 11 2
14 9 13 9 15 13 0 9 9 15 0 11 0 9 2
17 9 13 9 12 11 9 13 13 9 2 7 9 1 11 7 11 2
21 16 3 9 13 9 13 9 2 3 9 7 9 9 13 11 11 9 11 11 9 2
8 9 13 9 9 0 9 12 2
23 11 13 9 9 0 9 12 1 2 15 1 9 13 3 0 9 11 11 1 9 11 11 2
15 11 9 9 13 3 9 9 9 7 11 9 7 15 9 2
9 15 13 0 9 2 0 9 2 2
13 9 9 9 9 7 9 13 9 3 15 15 9 2
14 9 13 3 15 2 16 9 9 9 13 12 0 9 2
16 3 3 0 13 0 9 12 13 9 2 15 13 9 3 9 2
10 15 13 0 9 0 2 0 9 2 2
15 9 4 13 9 12 9 0 9 2 7 13 3 13 15 2
14 3 9 13 3 3 9 9 7 9 2 16 0 9 2
23 3 0 9 9 13 12 9 2 15 9 11 13 0 1 13 0 9 9 7 15 9 9 2
7 9 9 13 3 9 0 2
15 11 13 3 9 1 0 9 2 15 13 9 9 3 3 2
8 2 12 11 13 9 9 9 2
8 2 12 11 13 9 0 9 2
10 2 12 11 13 11 9 2 11 2 2
8 2 12 11 13 11 9 9 2
19 3 9 13 3 11 13 9 7 13 13 11 9 9 11 9 7 9 9 2
12 16 9 9 9 12 13 2 3 11 13 9 2
13 15 13 3 11 2 0 9 13 11 9 13 9 2
5 9 15 13 9 2
8 15 13 3 0 9 9 9 2
8 3 15 13 7 13 3 3 2
6 15 13 0 9 9 2
17 9 15 13 7 2 11 11 11 2 7 3 2 11 11 11 2 2
18 11 11 2 3 13 9 11 11 11 2 13 11 7 11 3 13 9 2
34 9 9 13 3 3 11 11 2 9 2 9 2 2 11 11 2 9 2 0 9 2 2 7 11 2 11 2 11 2 9 2 9 2 2
12 0 9 11 11 11 13 0 11 9 9 12 2
9 11 11 13 9 12 13 0 9 2
4 9 13 9 2
15 9 13 9 0 9 2 3 3 3 11 9 13 11 9 2
12 9 12 1 9 4 13 3 9 0 11 9 2
12 11 11 13 9 0 9 3 12 12 9 9 2
31 9 13 9 15 9 13 7 13 9 2 15 13 0 9 1 15 0 9 2 3 9 2 9 2 9 2 9 2 9 3 2
10 0 13 3 9 2 9 7 9 9 2
11 9 13 9 3 0 7 3 15 13 9 2
14 15 4 13 9 9 2 9 9 7 9 9 13 9 2
19 9 4 13 3 9 3 9 2 15 0 9 9 13 9 13 7 9 13 2
15 9 9 13 13 9 9 9 2 16 9 9 13 9 9 2
7 3 9 13 9 13 9 2
15 11 11 11 2 13 0 9 12 2 13 0 9 0 9 2
12 15 13 9 0 9 12 7 9 0 9 12 2
11 9 13 11 13 11 9 9 11 9 12 2
8 9 12 15 13 11 9 9 2
15 11 11 11 2 12 2 0 9 12 2 13 11 13 9 2
12 15 13 9 0 7 13 0 9 9 13 9 2
9 0 9 13 0 9 13 9 9 2
18 0 0 9 13 9 9 9 9 2 7 15 4 13 9 13 15 9 2
19 0 0 9 9 13 9 0 9 2 9 13 8 2 9 8 7 9 8 2
12 9 9 13 0 9 9 13 9 0 9 9 2
19 15 3 2 5 2 13 2 5 2 9 7 2 5 2 2 5 2 9 2
21 9 13 9 2 15 13 3 9 13 9 7 9 2 3 9 2 9 2 9 3 2
11 16 13 9 13 0 2 13 9 3 9 2
6 0 9 13 9 9 2
16 11 11 2 13 0 9 12 11 2 11 2 13 0 0 9 2
14 0 9 13 11 13 9 12 11 11 11 9 12 9 2
8 9 15 4 13 11 11 9 2
12 9 13 9 13 9 2 15 13 3 11 9 2
16 9 13 13 9 0 9 7 15 9 9 3 13 3 9 9 2
6 15 9 13 9 9 2
10 0 9 13 0 9 1 9 0 9 2
10 9 13 3 12 9 2 9 12 2 2
11 2 12 2 11 11 13 9 9 11 9 2
13 2 12 2 9 11 11 9 2 9 2 13 9 2
8 2 12 2 11 13 11 15 2
7 2 12 2 9 13 11 2
15 2 12 2 11 9 2 11 9 11 0 4 13 11 11 2
5 11 13 9 11 2
10 2 12 2 11 11 9 11 9 11 2
23 2 12 2 11 13 15 2 9 11 9 2 2 11 11 11 2 2 12 12 9 9 11 2
32 2 12 2 11 9 11 0 13 9 0 11 0 9 1 9 12 7 0 0 9 2 15 9 13 13 11 7 11 1 9 12 2
9 2 12 2 11 11 13 0 9 2
23 2 12 2 2 11 2 13 0 9 3 13 9 9 0 9 2 2 11 11 11 2 2 2
9 2 12 2 11 11 13 11 9 2
22 2 12 2 11 9 2 3 2 12 9 9 2 2 13 3 9 3 12 9 9 1 2
18 0 9 13 3 0 9 0 7 0 13 9 13 3 9 7 9 9 2
8 15 9 0 9 13 13 9 2
29 9 13 3 15 2 7 9 13 9 9 2 15 13 3 13 3 2 16 13 13 9 2 13 3 9 13 0 9 2
18 0 9 4 13 0 9 2 15 13 9 13 2 16 0 9 13 13 2
6 11 13 9 0 9 2
8 9 15 13 9 7 9 1 2
25 3 12 9 9 4 13 0 2 13 9 9 2 9 13 9 9 7 9 0 9 13 0 9 9 2
17 3 0 13 9 13 3 13 13 0 9 2 13 0 9 15 13 2
10 16 9 13 0 2 9 9 13 9 2
11 0 9 9 13 3 9 7 3 12 9 2
7 9 13 9 9 7 9 2
32 16 0 9 3 4 13 0 9 9 2 4 15 1 13 9 2 7 16 0 9 13 9 0 2 3 12 7 3 12 9 9 2
26 9 3 0 13 4 13 0 9 9 9 9 2 16 15 4 13 13 9 0 9 9 7 0 9 9 2
33 9 4 13 0 9 13 3 2 16 13 13 9 9 2 15 9 9 1 15 4 13 0 9 7 15 9 4 13 9 13 9 9 2
19 9 4 3 13 0 9 13 3 9 2 3 9 13 15 9 0 0 9 2
10 3 9 13 9 4 0 9 13 0 2
13 9 13 3 13 0 9 2 7 9 1 13 9 2
24 11 13 0 0 9 13 9 2 7 3 13 0 9 2 15 13 13 15 0 9 9 13 9 2
23 0 9 13 9 2 15 13 13 0 9 13 0 9 15 1 2 13 3 13 4 13 9 2
11 9 13 9 4 3 3 13 15 16 11 2
11 11 13 11 11 11 13 0 9 9 12 2
25 15 15 13 11 11 2 9 2 15 13 3 13 0 9 7 13 13 0 9 13 2 15 3 13 2
26 11 11 2 13 0 9 12 2 13 0 0 9 0 9 7 15 9 13 0 9 12 2 0 9 12 2
11 15 13 9 7 13 3 0 11 13 11 2
11 11 11 13 0 0 9 0 9 7 9 2
12 15 13 9 9 7 4 13 9 12 0 9 2
22 11 4 13 9 11 11 2 2 8 8 8 8 8 2 11 9 9 9 11 9 11 2
14 9 4 13 3 11 2 7 15 9 9 9 13 3 2
14 11 13 12 0 9 9 11 7 13 9 15 9 11 2
28 9 13 15 9 2 7 15 4 15 1 13 9 9 7 9 1 7 13 11 11 13 9 0 9 11 11 9 2
14 11 4 13 9 3 9 11 11 11 11 11 11 11 2
9 9 2 11 11 2 13 0 9 2
22 9 9 13 3 12 9 2 15 9 9 12 9 2 9 9 12 9 7 9 12 9 2
15 9 13 9 3 9 9 7 15 13 0 0 9 0 9 2
10 15 13 0 9 2 15 3 13 3 2
4 9 13 0 2
13 9 13 0 7 9 13 3 11 7 13 3 0 2
8 9 13 0 7 3 3 0 2
5 3 9 13 0 2
5 9 13 3 0 2
23 9 9 13 0 2 9 0 2 7 9 9 13 0 7 9 0 2 9 9 13 3 0 2
16 0 9 13 0 7 15 9 13 0 2 9 0 7 9 0 2
13 9 13 11 9 2 11 9 7 11 7 11 9 2
8 15 9 9 13 12 12 9 2
18 9 13 3 9 2 3 0 9 4 3 13 2 13 15 4 13 11 2
19 9 13 9 7 0 9 9 2 3 9 2 9 3 12 12 9 9 1 2
12 11 9 13 3 9 7 9 7 0 9 9 2
24 9 13 9 2 15 13 12 0 13 9 7 9 13 9 2 15 13 3 15 9 9 0 9 2
12 9 13 0 9 7 9 13 13 0 9 1 2
9 15 3 9 0 9 13 3 0 2
14 9 9 13 12 9 7 3 15 4 13 0 9 9 2
14 9 13 13 3 7 3 3 0 9 9 13 9 9 2
19 9 13 9 9 7 9 12 9 0 7 3 3 0 9 9 7 9 1 2
15 3 3 0 9 13 9 9 7 3 3 9 15 9 13 2
22 9 13 9 1 9 7 0 9 13 0 0 9 2 15 13 13 0 9 12 9 3 2
7 9 13 12 12 0 9 2
10 3 4 12 7 0 9 13 15 9 2
11 0 9 13 9 3 7 9 15 9 3 2
5 9 13 12 9 2
15 15 9 9 13 7 13 9 2 15 13 9 12 9 9 2
10 9 4 13 12 7 3 12 9 9 2
6 9 13 0 3 9 2
22 16 9 13 0 9 3 2 4 0 9 13 9 3 12 9 13 0 9 7 13 3 2
31 9 13 9 0 9 2 16 12 9 13 9 13 3 3 9 16 0 9 13 9 2 13 9 9 9 2 3 9 4 13 2
9 9 4 13 9 13 9 0 9 2
8 9 1 9 13 3 7 9 2
4 9 13 0 2
23 15 13 7 9 7 9 7 9 2 9 2 9 2 9 2 0 9 2 9 7 9 9 2
7 15 13 9 9 7 9 2
11 9 4 13 9 2 15 15 13 3 13 2
7 3 9 13 9 7 9 2
12 11 11 11 13 9 12 9 13 9 1 9 2
14 15 9 13 13 11 9 0 9 15 13 11 11 11 2
14 11 11 11 13 3 9 15 9 7 9 13 15 9 2
29 9 12 11 13 0 11 3 2 7 15 13 12 9 7 15 13 11 9 2 11 11 11 2 2 0 11 9 2 2
23 9 12 11 4 13 3 9 7 15 13 12 9 15 13 12 0 9 11 0 7 0 9 2
10 9 12 13 3 11 11 11 0 9 2
21 15 13 3 12 9 2 11 11 11 11 7 11 11 11 11 5 11 11 11 11 2
26 9 12 11 13 0 9 11 2 11 2 11 2 11 2 11 2 11 11 2 11 11 2 11 7 11 2
3 7 11 2
7 3 15 13 0 11 11 2
6 3 11 13 12 9 2
17 9 12 11 13 0 7 0 9 0 9 9 12 2 11 9 2 2
26 15 13 11 0 11 11 11 7 15 13 11 9 2 7 15 13 12 9 2 0 9 1 3 12 3 2
3 3 9 5
11 11 2 9 11 2 13 11 9 13 9 2
18 9 13 0 3 15 9 13 11 11 11 9 13 9 7 0 11 9 2
15 11 9 13 3 12 9 7 15 9 13 3 12 0 9 2
14 11 9 13 3 11 9 2 15 13 9 12 0 9 2
9 11 4 13 15 3 0 0 9 2
6 11 9 13 9 9 2
14 16 9 13 11 9 2 13 11 9 9 9 9 1 2
15 9 13 9 13 3 0 9 2 15 15 13 3 9 1 2
12 11 9 9 13 9 9 13 12 9 9 9 2
14 16 9 13 0 9 2 0 9 13 3 9 9 9 2
21 15 0 9 13 9 11 11 11 9 9 12 2 15 13 12 12 9 13 11 9 2
14 9 9 13 0 9 7 9 13 9 3 3 9 9 2
17 0 9 13 9 13 15 9 0 9 2 0 9 7 0 9 9 2
13 11 11 2 13 0 9 12 11 2 13 0 9 2
13 15 4 13 9 3 3 11 11 7 11 11 1 2
11 11 13 0 9 7 4 13 0 3 9 2
13 11 11 11 2 13 0 9 12 2 13 0 9 2
5 11 13 11 11 2
14 11 4 13 3 9 11 11 2 11 11 7 11 11 2
10 11 13 3 9 9 9 2 11 11 2
14 11 11 2 13 0 9 12 2 11 2 13 0 9 2
11 11 13 0 9 9 7 12 9 11 11 2
7 15 13 9 11 9 9 2
8 15 13 11 9 9 9 12 2
8 11 13 9 1 11 11 9 2
15 9 12 15 13 11 11 13 11 11 7 13 3 11 9 2
27 11 11 2 13 0 9 12 2 11 2 13 3 3 0 9 2 15 0 9 13 11 11 0 9 0 9 2
11 11 4 13 3 9 12 9 11 7 11 2
6 9 1 11 13 9 2
9 9 12 15 13 11 11 9 9 2
9 9 12 15 13 9 11 11 11 2
8 11 11 13 9 11 11 9 2
6 11 13 0 0 9 2
16 15 13 3 15 13 9 2 7 15 9 4 13 3 9 9 2
10 11 13 11 9 2 9 13 11 11 2
14 11 13 3 9 2 9 2 0 9 7 15 9 9 2
10 3 11 13 3 7 3 15 9 1 2
6 11 13 9 3 3 2
6 11 13 13 3 9 2
14 15 4 13 9 9 9 9 2 7 0 9 13 13 2
16 11 13 9 2 13 13 9 9 13 0 9 9 11 9 0 2
9 11 4 13 0 9 13 9 9 2
16 11 13 9 9 2 7 15 13 9 3 15 4 13 0 9 2
13 11 0 9 13 5 2 9 12 9 7 9 12 2
12 11 4 13 0 9 3 12 9 7 12 9 2
23 9 11 11 13 3 12 9 2 12 9 0 9 2 7 9 13 3 12 9 2 12 9 2
14 11 13 13 13 9 2 9 2 9 7 3 9 1 2
8 15 4 13 9 2 9 3 2
8 9 7 9 4 13 9 3 2
8 9 2 11 11 2 13 9 2
15 9 13 9 3 12 9 0 2 9 15 9 13 9 15 2
6 15 13 9 0 0 2
12 9 7 9 13 0 0 9 2 9 0 9 2
7 9 7 9 13 9 0 2
7 9 9 13 3 0 9 2
7 9 13 11 9 7 9 2
21 15 13 9 7 9 2 3 9 9 9 12 9 9 1 2 7 9 7 0 9 2
6 0 9 13 3 9 2
11 11 2 9 8 2 13 9 11 9 11 2
13 15 13 11 7 11 13 9 9 12 9 11 9 2
6 9 13 11 9 9 2
10 3 13 11 2 11 7 11 13 9 2
10 9 13 12 12 9 2 9 12 2 2
6 9 13 9 12 1 2
11 9 15 13 9 9 7 9 1 9 9 2
9 9 12 11 13 11 9 13 9 2
11 3 9 13 9 2 9 2 9 7 9 2
32 9 13 9 12 13 0 11 9 2 0 11 9 2 12 2 2 11 9 2 12 2 2 0 9 2 12 2 7 0 0 9 2
48 11 11 2 11 2 11 2 13 0 9 12 11 11 11 2 11 2 13 0 9 2 15 4 13 0 3 3 13 9 15 13 9 2 11 11 2 2 12 2 7 11 2 9 11 2 12 2 2
12 15 13 12 9 0 9 1 7 12 0 9 2
14 11 13 15 3 9 12 13 11 11 0 9 9 9 2
30 11 9 0 9 0 9 2 12 2 7 11 11 2 12 2 13 9 9 2 7 3 15 13 9 0 9 9 9 9 2
39 11 4 3 13 0 9 2 3 11 2 15 9 3 9 2 12 2 2 11 11 11 2 12 2 7 11 11 13 2 12 2 2 15 15 13 11 11 9 2
17 9 9 15 13 9 11 11 7 11 11 2 3 11 11 2 9 2
9 9 9 1 11 4 3 13 9 2
47 11 0 9 13 9 11 11 9 15 13 9 2 11 11 2 2 11 9 9 9 13 9 2 12 2 2 11 11 9 9 9 2 12 2 7 9 11 2 0 11 11 9 9 11 11 11 2
7 9 13 9 9 13 9 2
11 15 13 9 3 13 7 13 7 13 9 2
12 9 13 3 9 2 16 9 9 13 9 0 2
16 3 15 0 9 2 3 9 2 11 11 2 4 13 9 9 2
6 9 9 13 0 9 2
14 9 13 9 13 9 2 9 7 9 15 9 16 9 2
15 9 9 13 3 9 13 13 9 2 16 9 9 13 0 2
10 15 1 9 13 13 9 9 13 9 2
12 15 1 9 9 13 13 9 3 0 16 9 2
10 9 15 1 13 3 0 2 12 5 2
12 9 13 15 9 13 3 0 9 7 3 9 2
14 15 9 15 13 9 0 9 2 7 13 13 0 9 2
10 9 13 3 9 7 9 3 9 1 2
9 13 13 9 13 0 9 0 9 2
5 15 13 9 12 2
15 11 11 11 13 9 7 0 9 11 13 11 11 0 9 2
9 3 15 13 11 11 11 11 9 2
16 11 9 9 13 3 11 9 11 2 15 11 9 4 15 13 11
7 11 13 12 9 0 9 2
15 0 9 11 11 13 0 9 11 2 15 3 13 9 12 2
14 11 11 11 11 11 13 11 11 9 12 13 0 9 2
10 9 13 0 9 11 7 0 9 11 2
7 9 0 9 13 9 11 2
22 0 9 13 3 9 2 11 2 11 11 11 2 7 2 11 11 11 2 11 11 2 2
7 9 13 9 9 12 9 2
27 11 11 2 11 2 11 2 0 9 12 11 2 0 9 12 11 9 2 13 0 9 2 9 7 9 9 2
11 11 9 13 0 11 11 7 11 11 11 2
14 15 13 12 9 9 7 13 3 9 11 12 7 9 2
23 11 13 11 9 11 9 12 2 9 11 11 12 2 9 7 9 11 12 7 0 9 12 2
11 15 13 9 9 9 12 7 13 9 9 2
33 11 9 1 11 13 9 0 9 12 7 13 15 13 3 11 9 0 9 9 9 7 11 9 9 9 12 7 13 9 9 9 12 2
8 15 13 13 3 9 9 1 2
10 11 13 11 9 9 12 7 9 12 2
15 15 13 11 9 9 9 9 12 7 13 9 11 9 12 2
9 9 1 11 13 9 11 9 12 2
11 11 13 11 9 12 13 11 9 0 9 2
21 15 13 3 11 9 9 7 9 9 15 13 1 11 7 9 9 11 9 13 9 2
9 11 13 3 9 12 11 11 11 1
19 11 11 11 11 11 2 13 0 9 12 11 2 13 0 9 13 0 9 2
15 15 4 13 9 3 3 0 2 0 2 0 7 0 9 2
12 3 11 11 3 13 9 0 11 11 13 9 2
16 11 11 9 13 11 9 9 11 11 11 11 7 9 11 11 2
10 15 13 9 12 7 13 11 9 12 2
14 15 9 13 3 3 11 11 2 11 11 7 11 11 2
13 3 11 11 4 13 11 12 9 9 9 12 1 2
14 9 11 11 13 9 12 11 11 9 15 13 3 9 2
12 15 13 12 11 9 2 15 9 13 11 11 2
33 11 11 0 9 13 9 11 1 13 0 9 2 15 15 9 13 3 3 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2
13 11 11 13 3 12 11 9 7 12 9 9 12 2
13 0 9 13 9 11 11 9 9 11 2 12 2 2
27 3 11 11 4 13 3 3 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 7 11 11 9 2
7 11 11 4 13 3 3 2
14 9 13 9 11 11 1 2 12 2 15 13 12 9 2
9 9 11 11 1 15 4 13 12 2
17 11 11 11 2 13 0 9 12 2 11 2 11 2 13 0 9 2
10 15 13 3 0 9 7 3 0 9 2
17 11 9 4 13 3 3 11 11 2 11 2 11 11 7 11 11 2
11 11 11 11 9 13 11 15 9 0 9 2
21 11 11 9 4 13 3 11 9 9 2 15 13 3 9 12 9 11 11 7 11 2
11 11 13 9 0 11 9 9 11 13 9 2
26 3 11 13 9 11 9 2 7 15 13 3 15 11 7 13 0 9 2 15 1 15 9 13 0 9 2
17 11 13 9 11 0 9 2 9 11 9 7 9 7 9 11 9 2
13 0 9 11 13 13 7 9 13 0 11 9 9 2
17 1 11 9 9 2 9 12 2 11 13 11 9 2 9 11 9 2
9 9 11 9 13 0 11 9 9 2
20 9 11 13 13 2 7 9 12 9 1 15 4 3 13 7 9 13 3 11 2
22 9 9 13 3 9 12 7 9 13 13 9 2 7 12 4 9 3 13 7 9 13 2
14 3 9 13 15 3 9 2 7 9 13 13 0 9 2
14 11 12 7 11 12 13 0 11 9 12 11 13 9 2
10 11 12 13 0 9 12 9 12 9 2
6 9 9 13 12 9 2
8 11 9 15 13 0 9 12 2
8 3 9 13 11 9 9 1 2
15 12 9 9 9 13 7 9 9 13 9 9 13 9 9 2
19 11 12 13 9 5 0 2 5 0 2 9 12 9 9 11 12 9 9 2
12 9 1 11 12 9 13 9 7 13 11 9 2
17 9 13 12 9 0 12 5 7 12 9 9 2 12 9 2 9 2
9 9 13 9 9 9 13 9 9 2
20 0 9 9 13 11 12 13 0 15 9 9 13 9 2 9 9 12 13 0 2
13 11 9 2 9 8 8 8 2 13 11 0 9 2
6 15 13 1 11 9 2
7 11 9 13 11 0 9 2
8 11 13 3 15 0 9 11 2
14 11 11 2 5 12 2 12 2 13 11 11 9 9 2
19 9 9 11 11 11 1 13 11 9 11 2 15 9 13 12 15 13 9 2
20 12 11 11 13 9 11 11 9 9 13 15 1 9 2 15 13 9 0 9 2
11 15 13 9 7 13 0 9 11 0 9 2
9 15 4 13 9 9 7 11 9 2
15 11 9 13 13 9 12 2 7 11 11 13 13 15 9 2
12 11 11 13 9 9 1 7 13 3 9 9 2
12 12 15 13 11 7 13 3 0 9 15 9 2
11 9 12 11 11 11 13 9 11 11 9 2
10 15 9 13 13 0 9 9 9 1 2
11 11 11 13 15 9 0 11 9 11 11 2
12 12 11 11 13 11 9 13 3 13 13 9 2
14 0 9 9 3 13 7 11 11 13 13 15 0 9 2
12 15 13 9 9 0 1 15 13 3 13 15 2
8 13 11 9 15 13 12 9 2
18 0 9 11 11 13 13 9 3 16 11 11 11 4 13 9 0 9 2
22 12 13 0 9 9 7 9 1 11 11 2 9 13 11 11 15 13 11 11 9 9 2
18 16 11 11 13 13 9 3 0 15 13 9 11 11 9 7 13 11 2
12 15 13 9 13 12 7 15 13 0 9 12 2
18 11 11 2 13 0 9 12 2 11 2 11 2 11 2 13 0 9 2
13 15 13 3 9 11 9 2 15 15 13 9 11 2
22 15 4 13 3 9 11 11 2 11 11 2 9 9 2 9 11 2 11 7 11 11 2
7 15 4 13 3 9 11 2
13 11 13 0 9 2 15 13 9 11 9 12 9 2
14 9 0 9 13 9 11 11 2 11 11 7 11 11 2
7 9 13 13 9 7 9 2
10 9 9 13 0 9 9 9 13 9 2
12 9 13 9 2 11 9 2 15 13 9 12 2
7 11 13 9 12 13 9 2
14 0 9 9 9 13 11 11 13 0 9 11 11 12 2
19 9 12 9 9 13 11 11 11 2 15 3 13 15 9 12 9 11 11 2
15 3 3 0 9 13 9 12 0 2 7 9 9 13 11 2
11 9 9 9 13 2 7 3 0 9 9 2
16 11 11 13 9 9 0 9 12 7 13 9 15 9 9 1 2
14 9 2 11 11 2 13 11 7 3 11 13 0 9 2
5 15 13 9 9 2
10 11 11 13 9 2 15 13 9 12 2
11 15 13 9 2 15 13 9 7 0 9 2
13 15 13 11 0 9 7 11 11 11 9 15 9 2
15 0 9 11 13 3 13 9 11 11 11 2 15 13 11 2
20 11 0 0 7 0 9 13 0 7 0 16 0 2 15 13 11 9 11 11 2
9 11 13 11 11 9 11 2 11 2
23 11 11 11 13 11 9 11 2 11 9 12 2 7 9 12 9 1 3 15 4 13 11 2
29 11 9 15 15 0 9 2 11 11 2 11 11 2 11 11 7 11 11 2 13 15 16 15 13 12 1 12 9 2
18 15 13 0 2 3 12 9 2 16 0 9 3 11 11 7 11 11 2
15 0 9 11 13 3 0 9 12 7 13 9 12 11 9 2
8 11 13 13 15 9 9 11 2
33 9 13 9 0 16 9 2 15 13 0 16 0 9 7 0 16 0 9 7 9 3 11 11 2 11 11 2 11 11 7 11 11 2
15 9 13 13 0 12 9 0 0 7 0 12 9 0 0 2
12 9 13 13 0 12 9 0 0 8 8 9 2
19 11 2 9 11 2 7 11 2 3 11 2 11 2 13 12 9 11 9 2
5 9 13 11 9 2
6 15 13 3 12 9 2
5 9 13 9 9 2
14 0 9 11 4 13 0 9 9 9 0 0 9 11 2
12 9 11 4 13 15 2 16 9 13 3 9 2
13 9 4 3 13 11 1 2 7 4 13 3 3 2
7 3 11 13 3 9 11 2
17 0 9 9 9 13 0 0 9 11 2 15 11 7 11 13 9 2
11 11 13 9 11 9 2 11 11 2 11 2
13 11 9 13 12 12 2 7 15 13 3 0 9 2
24 11 13 3 9 9 9 11 11 2 15 4 13 11 15 9 2 9 7 9 3 15 9 9 2
15 9 2 9 8 8 2 13 9 13 9 0 9 13 9 2
19 9 13 0 0 9 15 9 13 9 9 7 0 9 15 1 13 9 9 2
6 9 13 9 3 3 2
8 9 13 9 0 9 9 13 2
18 9 13 9 13 9 2 15 4 13 9 7 15 13 9 9 9 5 2
8 9 13 9 3 13 9 9 2
12 9 0 9 9 13 9 2 15 13 0 9 2
6 9 9 13 9 9 2
6 9 4 3 13 9 2
11 9 13 9 2 7 15 13 3 9 3 2
10 9 9 13 9 4 13 13 13 9 2
9 9 9 13 15 9 1 13 9 2
18 9 9 13 9 9 2 3 9 13 13 9 3 2 7 9 13 9 2
16 9 4 13 9 3 15 2 7 9 13 9 4 13 0 3 2
12 16 9 13 2 15 9 13 7 9 13 9 2
15 9 4 13 7 9 3 7 15 15 9 13 9 13 9 2
23 11 11 11 2 0 9 11 11 11 11 2 13 0 9 2 15 13 11 9 2 11 11 2
12 9 13 0 9 11 9 9 2 15 9 0 2
37 9 0 9 4 13 12 9 2 9 13 0 8 8 9 11 2 0 0 8 8 9 0 9 2 0 8 8 9 9 7 0 0 8 8 9 11 2
26 9 9 13 0 0 8 8 9 11 2 0 9 11 11 7 0 9 11 2 15 9 9 13 13 3 2
12 9 9 13 9 9 13 8 8 8 9 11 2
17 9 13 3 3 9 13 9 9 2 7 15 13 3 13 13 3 2
13 9 13 9 2 15 13 0 9 7 9 9 9 2
13 9 13 0 9 11 11 11 13 9 11 11 11 2
16 9 13 9 9 9 13 9 2 15 9 13 9 0 11 11 2
10 9 13 9 0 9 7 9 12 12 2
9 9 13 9 0 9 9 11 9 2
7 9 13 3 3 12 12 2
16 9 9 13 0 11 11 2 15 13 9 1 3 3 11 9 2
17 9 9 13 0 8 8 9 11 2 15 13 9 0 9 7 9 2
11 9 13 9 9 2 15 9 15 9 13 2
12 11 11 11 12 13 3 0 3 11 9 9 2
5 9 13 3 12 2
19 9 13 9 11 2 15 1 13 11 7 11 1 13 0 8 8 9 11 2
12 9 3 0 9 13 0 2 0 9 13 11 2
19 9 13 0 11 7 0 11 2 15 9 13 9 11 11 11 11 11 9 2
19 15 9 1 11 11 11 9 13 13 9 3 0 9 2 13 9 0 9 2
16 11 2 9 11 7 11 2 13 11 9 9 7 9 0 9 2
7 9 1 11 13 11 9 2
9 11 13 13 9 0 9 0 9 2
9 9 1 11 13 9 9 1 11 2
12 9 13 12 9 9 11 2 15 13 0 9 2
23 9 9 13 3 9 1 9 2 15 13 11 13 13 9 0 0 9 2 15 13 15 9 2
10 9 13 11 2 15 13 9 11 9 2
7 11 7 11 13 11 9 2
9 11 11 4 13 11 9 9 11 2
8 11 11 13 11 9 9 12 2
20 15 13 3 11 11 11 9 15 13 4 13 15 9 7 11 11 9 9 12 2
12 11 9 9 9 11 11 4 13 9 7 9 2
29 11 2 11 2 11 2 13 0 9 12 11 2 11 2 13 0 9 9 2 15 3 13 11 11 11 11 11 11 2
23 15 11 9 9 13 12 9 2 15 11 4 13 12 9 7 13 12 9 7 13 12 9 2
7 9 15 4 13 12 9 2
26 11 11 9 9 13 11 4 13 12 9 2 7 13 12 9 12 9 7 12 9 2 9 13 12 9 2
12 15 13 9 9 11 11 11 11 9 11 11 2
10 11 11 9 13 0 9 11 11 12 2
16 15 13 11 11 11 9 12 2 15 11 13 15 11 9 12 2
8 9 12 9 15 13 11 9 2
8 11 11 11 13 11 13 9 2
15 15 13 11 0 11 11 11 9 3 2 16 15 13 9 2
10 9 2 11 11 2 13 11 0 9 2
11 15 13 11 3 12 9 0 3 9 1 2
8 9 9 4 13 3 12 9 2
23 9 9 13 0 9 2 15 13 9 7 9 9 0 2 9 2 7 9 0 2 9 2 2
17 9 13 0 0 11 7 9 15 13 3 9 7 9 9 9 13 2
9 3 3 9 13 9 3 0 9 2
7 9 13 3 0 9 9 2
8 15 4 13 15 0 9 9 2
5 9 13 9 13 2
9 3 0 9 13 3 9 13 9 2
5 9 9 13 9 2
18 11 9 2 13 11 2 13 11 9 9 11 9 11 9 11 9 11 2
12 9 9 11 9 13 12 9 13 11 9 1 2
6 9 13 13 3 9 2
11 9 13 0 9 2 7 3 13 3 9 2
20 9 11 9 7 9 9 11 9 13 9 2 7 0 9 13 9 0 9 12 2
11 11 9 7 9 13 3 9 11 9 1 2
18 11 0 2 9 9 2 0 9 12 2 0 9 12 2 13 11 12 2
10 9 12 11 7 9 11 0 1 9 2
6 11 13 9 9 9 2
12 9 12 7 12 15 13 9 9 11 0 1 2
12 0 9 9 15 13 11 9 1 11 7 11 2
6 11 15 13 9 9 2
20 15 13 11 12 7 13 9 12 9 11 0 9 1 2 9 7 9 9 9 2
9 0 9 12 15 13 11 11 11 2
21 15 12 9 13 2 0 11 9 11 0 11 0 2 9 9 0 11 7 11 9 11
19 11 11 11 12 13 11 11 9 9 2 15 13 0 9 12 11 11 9 2
11 9 13 9 0 2 7 15 13 11 11 2
6 9 13 11 9 0 2
14 11 11 13 0 9 9 2 15 1 11 9 13 9 2
4 11 11 9 9
13 11 11 9 0 9 11 11 13 3 11 9 9 2
20 11 11 11 9 13 9 9 2 16 15 1 13 3 0 11 13 0 9 9 2
3 11 9 12
5 11 13 3 9 2
23 9 13 13 3 9 3 2 12 12 12 9 7 12 5 15 13 9 2 15 13 9 12 2
5 9 9 13 12 2
23 11 2 11 7 11 13 15 9 0 9 2 3 16 9 13 13 2 13 9 7 3 9 2
16 3 0 12 9 9 13 3 0 9 2 3 3 9 13 9 2
18 11 9 12 13 9 1 9 13 0 9 2 11 13 0 7 9 0 2
6 15 9 9 13 0 2
15 15 9 13 9 0 9 2 15 15 13 15 9 3 9 2
10 3 9 13 12 9 3 16 0 9 2
9 15 12 0 9 13 3 3 9 2
14 15 9 13 9 1 12 12 9 3 16 12 9 1 2
8 11 9 13 13 9 9 9 2
9 9 11 13 12 7 11 12 9 2
25 11 3 13 12 0 9 2 3 9 13 12 9 11 9 0 9 1 11 2 15 9 13 3 12 2
15 11 13 3 12 9 2 16 9 13 3 3 12 9 9 2
2 11 9
9 11 9 11 13 9 0 9 12 2
18 11 9 13 13 9 7 9 2 15 13 3 12 9 7 12 9 9 2
14 11 11 1 9 4 13 12 9 9 7 3 12 9 2
9 0 9 13 9 1 3 12 9 2
7 9 4 9 1 13 3 2
11 9 9 9 12 1 4 13 9 9 12 2
16 9 9 13 3 15 9 12 2 16 9 13 11 9 13 9 2
11 9 9 13 12 2 12 9 7 12 9 2
6 3 9 13 9 9 2
19 11 11 9 1 9 13 11 9 13 13 9 13 9 2 15 9 13 0 2
15 9 9 11 11 1 15 9 13 3 0 7 9 9 0 2
6 15 4 13 15 9 2
16 9 13 13 9 9 3 9 2 7 9 1 9 13 12 9 2
12 9 9 13 3 2 7 9 13 9 13 0 2
14 15 9 4 13 0 9 7 9 9 13 9 9 9 2
11 13 9 13 3 12 9 11 11 11 9 2
21 9 4 3 3 13 9 11 9 7 11 2 15 15 4 13 9 7 9 0 9 2
14 3 9 13 9 9 4 13 2 13 9 4 3 13 2
9 9 4 3 13 0 15 9 11 2
2 9 9
9 9 11 7 9 1 13 9 9 2
15 9 4 13 9 3 3 2 7 0 9 9 13 4 13 2
11 0 9 13 9 1 9 9 13 3 9 2
23 11 9 11 11 13 13 9 9 0 9 7 15 2 15 9 9 4 3 9 13 7 13 2
13 16 9 13 13 9 2 13 9 9 3 9 9 2
15 9 4 3 13 9 2 7 0 9 9 13 9 4 13 2
13 15 2 15 9 4 13 2 13 4 13 3 13 2
6 11 4 13 0 9 2
8 15 9 13 13 12 12 9 2
6 13 9 13 13 9 2
7 11 13 11 11 1 0 9
18 9 1 13 11 11 2 15 13 3 13 11 11 7 13 15 11 11 2
9 11 13 11 11 11 0 9 9 2
7 0 9 13 9 0 9 2
17 15 9 15 4 3 13 13 3 13 13 9 9 0 9 9 1 2
7 15 13 9 9 0 12 2
3 11 13 9
6 11 9 13 3 9 2
22 9 13 3 2 16 15 9 13 13 3 13 9 7 11 4 13 9 3 3 15 9 2
27 11 9 11 11 1 9 13 9 1 0 3 9 2 9 13 0 9 1 7 13 15 2 16 9 13 9 2
35 11 9 13 9 2 3 0 2 11 9 2 2 12 9 3 12 9 2 9 9 3 3 12 9 3 12 9 7 9 12 9 3 12 9 2
8 9 13 9 0 9 0 9 2
9 11 0 9 9 9 13 9 9 2
21 12 9 9 2 11 0 9 9 2 13 3 12 9 2 16 15 3 13 12 9 2
4 11 11 13 9
11 0 9 11 13 11 11 13 0 7 9 2
9 11 13 9 11 9 11 11 9 2
10 11 13 9 11 7 11 0 9 1 2
7 9 13 11 0 11 9 2
10 11 13 9 9 12 9 11 0 9 2
9 15 13 11 11 11 9 9 12 2
15 0 11 11 9 11 13 3 13 9 9 7 9 9 12 2
12 15 4 13 3 3 3 11 2 11 7 11 2
9 11 13 13 9 11 2 11 9 2
9 15 13 9 1 12 3 0 9 2
6 11 13 9 12 9 2
5 9 13 11 7 11
14 9 13 9 9 7 9 2 15 9 13 9 13 9 2
7 9 13 9 13 9 12 2
16 9 4 13 9 12 11 12 0 9 12 7 15 1 3 3 2
13 11 9 9 13 11 1 9 12 0 3 13 9 2
21 3 11 11 13 7 9 11 11 13 11 11 7 11 9 13 1 12 9 9 11 2
23 11 9 7 9 4 13 9 12 9 3 16 11 9 12 2 16 9 13 3 0 11 13 2
13 9 12 11 13 9 9 0 9 9 7 9 1 2
6 9 4 13 12 9 2
21 9 1 9 4 13 12 9 7 13 3 12 12 9 9 2 15 4 4 13 9 2
10 9 13 11 2 11 2 11 7 11 2
11 15 9 4 13 12 12 9 9 9 9 2
20 9 4 13 9 0 9 2 11 11 2 9 2 2 11 2 11 7 11 11 2
11 9 13 9 12 9 9 13 9 11 11 2
9 15 13 9 9 11 9 9 12 2
16 11 11 2 11 11 7 11 11 4 15 12 3 13 13 15 2
19 11 9 13 12 12 9 11 11 9 9 11 9 9 12 13 9 9 9 2
11 11 11 13 13 11 11 9 9 9 12 2
12 9 9 11 11 1 12 12 9 13 13 9 2
9 9 11 13 11 11 7 11 11 2
10 11 11 13 3 11 11 7 9 9 2
6 15 13 9 11 9 2
11 11 9 12 12 9 9 2 9 13 11 1
15 0 9 1 11 11 13 9 12 0 9 9 7 0 9 2
14 3 9 12 13 3 11 9 9 0 11 9 9 12 2
20 9 4 13 11 1 2 15 4 13 9 11 3 12 12 9 2 15 9 2 2
10 9 12 9 4 13 3 3 0 9 2
10 2 9 9 2 12 9 2 2 11 9
9 2 11 2 12 9 2 2 11 9
11 2 9 9 11 2 12 9 2 2 11 9
12 2 2 9 9 9 2 0 9 2 12 9 2
24 11 9 9 4 13 9 9 2 11 2 9 2 11 2 9 2 11 2 9 2 9 7 9 2
9 12 0 9 4 13 11 13 9 2
7 11 13 4 13 15 9 2
100 12 9 9 9 4 13 2 9 9 9 12 9 2 9 9 12 9 2 9 12 9 2 9 12 9 2 11 12 9 2 11 9 12 9 2 11 9 12 9 2 9 9 12 9 2 11 9 9 12 9 2 11 9 9 12 9 2 9 12 9 2 11 9 12 9 2 9 9 11 12 9 2 9 12 9 2 9 12 9 2 11 12 9 2 11 9 2 11 12 9 2 11 9 12 9 2 9 9 12 9
9 12 0 9 4 13 11 13 9 2
7 11 13 4 13 15 9 2
4 9 13 9 11
29 11 0 9 13 0 9 9 13 0 9 12 9 11 11 9 13 9 1 2 15 9 9 1 13 11 9 11 1 2
16 9 13 11 13 11 11 7 11 11 13 9 15 1 13 9 2
22 11 0 9 2 9 11 2 13 9 2 15 13 3 3 9 11 11 7 9 11 11 2
27 9 1 9 13 9 7 9 9 13 15 2 0 9 0 9 0 9 9 13 7 9 13 9 3 0 9 2
9 9 13 9 13 9 9 9 9 2
10 9 11 11 13 9 13 9 9 9 2
16 9 1 13 9 11 11 9 3 13 9 2 11 11 11 9 2
22 9 13 11 7 11 13 9 3 9 12 9 9 11 11 2 7 3 9 7 9 9 2
5 3 9 13 9 2
15 9 9 13 9 13 11 2 7 11 11 1 11 13 9 2
15 0 11 9 1 9 4 13 13 9 9 11 2 9 2 2
13 11 13 0 11 9 9 2 16 9 13 3 9 2
10 11 13 9 9 4 13 11 11 11 2
9 15 13 0 11 9 11 9 9 2
5 11 9 13 11 9
11 11 9 13 11 11 13 9 7 0 9 2
14 0 9 11 0 9 11 13 13 9 11 11 13 9 2
18 9 11 11 13 11 9 9 13 9 2 15 9 13 13 3 0 9 2
7 15 11 9 9 4 13 2
16 9 13 11 1 13 9 11 11 13 9 13 0 9 9 9 2
7 11 13 13 11 9 9 2
16 9 11 11 4 13 13 9 11 11 1 9 1 9 9 11 2
9 9 13 11 9 13 3 9 9 2
15 15 13 13 9 2 16 11 13 9 9 9 7 9 9 2
12 0 9 13 9 4 13 3 0 7 0 9 2
11 11 13 15 9 7 9 4 13 0 9 2
10 12 9 13 11 9 12 9 9 11 2
20 9 1 9 13 13 3 7 16 15 13 11 13 3 9 7 3 9 1 0 2
18 11 9 11 11 4 13 13 9 9 9 9 9 0 9 11 11 1 2
13 9 9 13 12 0 9 2 9 2 9 7 9 2
7 15 13 9 11 7 11 2
13 15 13 9 2 9 7 9 7 13 9 11 9 2
10 11 11 2 0 9 2 13 11 9 2
10 11 11 2 9 13 9 11 11 1 2
23 9 1 9 11 13 11 9 7 15 13 11 9 13 7 9 2 9 2 15 13 9 9 2
21 9 11 11 13 2 3 13 0 13 0 0 9 2 15 9 13 9 13 9 2 2
7 9 9 13 3 13 9 2
7 11 11 4 13 11 9 2
9 11 11 9 1 11 13 0 9 2
6 11 13 9 9 9 2
7 11 13 13 0 9 9 2
9 11 13 11 9 2 9 7 9 2
10 11 13 9 3 2 11 9 9 9 0
21 11 9 9 9 9 13 2 16 0 9 3 12 5 9 13 13 9 11 11 9 2
33 0 2 9 12 9 13 9 13 13 13 9 2 12 5 13 3 9 9 9 9 13 12 5 2 2 3 15 9 9 9 13 3 2
14 9 9 13 9 0 9 3 3 13 9 7 13 9 2
15 9 9 7 15 9 2 3 0 9 13 9 13 0 9 2
17 0 9 1 9 11 4 4 13 9 12 2 3 15 0 9 13 2
15 9 1 15 9 4 13 3 3 16 15 13 13 3 9 2
20 2 3 2 13 13 0 9 2 15 4 13 9 11 15 9 0 9 0 9 2
14 2 3 2 9 3 13 9 9 9 2 9 7 9 2
11 11 9 9 13 9 13 3 0 9 9 2
35 11 9 13 3 9 9 0 9 1 3 3 3 9 2 7 12 9 1 15 13 0 9 2 3 9 13 9 9 2 13 0 9 3 11 2
17 9 13 11 9 13 9 9 7 13 9 3 11 0 9 0 11 2
6 11 9 13 3 9 2
20 11 9 11 11 7 11 9 11 11 4 15 3 13 13 9 3 9 9 9 2
11 11 3 13 9 9 12 12 9 9 12 2
3 11 13 9
10 11 13 9 0 9 11 11 9 9 2
15 11 9 11 11 11 13 9 9 12 12 9 3 13 9 2
14 11 11 7 11 11 13 9 13 9 0 9 7 9 2
7 9 13 12 9 9 9 2
15 11 11 13 9 11 7 13 12 9 11 11 11 7 9 2
12 11 11 11 13 3 4 13 15 0 0 9 2
13 11 11 13 11 9 9 12 7 13 0 11 11 2
9 9 13 9 15 9 11 11 1 2
16 11 1 11 4 3 13 13 9 11 7 13 13 9 11 9 2
13 11 13 9 9 15 13 11 11 11 9 11 9 2
14 3 11 13 11 11 11 1 9 12 0 9 11 11 2
10 13 9 13 11 11 13 11 11 9 2
5 0 9 13 9 11
9 11 9 4 13 9 0 9 9 2
20 9 4 13 9 9 2 15 1 15 9 9 11 9 13 9 11 9 13 9 2
17 9 9 13 0 11 7 11 9 13 9 9 7 11 13 9 11 2
15 9 13 13 7 0 9 2 11 2 7 3 0 9 1 2
5 11 11 0 0 9
34 11 11 13 9 11 11 11 11 9 13 1 9 0 9 16 11 11 13 12 12 9 9 8 9 9 2 11 12 11 11 11 11 2 2
6 9 13 0 11 11 2
7 9 9 13 12 12 9 2
20 11 13 15 9 11 3 13 12 9 9 9 0 7 15 9 13 3 3 9 2
10 0 11 4 9 9 13 13 9 9 2
10 9 1 11 9 13 1 12 12 9 2
3 9 13 11
10 3 0 0 9 13 9 11 15 9 2
19 9 4 13 0 9 1 11 7 11 9 15 9 16 13 9 13 9 9 2
7 9 13 9 13 3 9 2
7 9 13 9 12 9 9 2
11 9 13 3 2 0 9 13 9 0 9 2
6 15 13 3 13 9 2
5 9 13 3 9 2
8 9 13 9 3 1 12 9 2
5 9 9 13 9 13
11 9 9 13 0 9 13 12 9 9 11 2
18 9 13 9 9 13 9 1 2 16 9 4 13 9 9 0 9 9 2
24 9 13 9 9 13 3 3 12 9 2 7 9 13 15 12 9 7 13 9 3 12 9 9 2
12 15 9 9 13 9 12 9 13 9 9 9 2
11 12 9 13 9 0 9 13 3 12 9 2
5 11 9 0 9 11
7 11 13 9 0 9 11 2
6 11 9 13 9 9 2
9 0 0 9 4 13 0 0 9 2
7 15 13 13 0 9 1 2
17 0 9 11 9 11 13 9 2 15 0 9 13 13 9 7 9 2
9 9 1 9 9 13 13 7 13 2
5 11 12 0 0 9
17 0 9 11 13 9 9 1 12 0 0 9 2 13 9 13 9 2
11 0 9 13 7 9 7 9 7 9 9 2
13 0 9 13 3 11 11 2 11 9 7 11 9 2
10 15 12 13 15 9 3 0 9 9 2
10 9 12 3 12 12 9 13 11 9 2
12 3 9 0 9 13 15 9 2 13 11 9 2
3 11 9 0
12 15 0 9 9 2 11 11 13 0 12 9 2
10 15 13 9 11 9 13 9 11 9 2
5 9 13 12 9 2
23 9 9 9 13 11 9 9 9 11 11 2 15 9 0 9 13 11 11 0 9 7 9 2
16 11 9 4 13 2 16 9 13 9 15 15 15 9 4 13 2
27 0 9 9 9 13 0 9 2 16 4 13 15 9 3 7 3 7 3 13 3 2 16 13 13 9 1 2
8 9 13 3 13 3 15 9 2
9 9 11 11 13 0 9 11 9 2
7 9 11 13 0 9 12 2
16 9 9 1 15 3 3 13 9 7 3 15 13 9 9 11 2
27 9 13 11 9 3 9 9 7 15 0 9 13 9 13 3 9 0 7 15 9 9 13 3 12 9 9 2
11 9 11 13 13 3 12 9 1 9 9 2
12 9 13 11 11 9 13 3 9 1 9 9 2
7 3 13 9 9 9 9 2
16 9 3 0 9 4 13 9 2 7 3 13 13 9 9 13 2
12 11 9 11 9 13 13 3 12 9 9 9 2
15 9 1 11 11 13 13 9 11 9 3 9 11 11 1 2
15 9 0 9 9 13 3 12 9 2 15 12 9 13 3 2
35 3 2 12 2 9 13 3 3 0 11 11 2 9 9 12 2 2 0 11 11 2 9 9 12 2 7 0 11 11 2 9 9 12 2 2
4 9 9 11 9
13 13 0 9 2 9 11 11 13 11 1 11 9 2
10 9 9 13 9 7 15 13 13 9 2
14 15 9 7 9 4 13 13 9 9 2 15 13 9 2
19 11 9 4 13 2 16 9 9 13 12 9 9 7 15 0 9 0 9 2
18 9 4 3 13 2 16 9 4 13 9 9 7 13 11 11 13 9 2
13 9 13 1 15 9 2 15 9 11 13 9 9 2
22 11 11 13 9 11 11 11 11 2 16 15 13 3 12 9 1 11 9 0 9 13 2
8 9 7 9 11 0 0 9 11
15 9 7 9 11 0 13 9 0 9 9 12 11 0 9 2
27 0 9 7 9 2 0 9 7 9 2 7 9 2 9 7 9 9 13 9 13 9 9 3 12 12 9 2
9 13 9 4 3 13 0 0 9 2
12 9 13 9 1 9 3 0 9 12 9 9 2
16 9 11 0 13 0 9 9 2 15 0 9 4 3 9 13 2
15 0 9 13 3 9 7 9 2 9 7 0 9 7 9 2
20 3 9 13 3 3 9 2 9 7 0 9 7 9 7 0 9 9 7 9 2
18 3 3 9 13 3 9 7 9 2 9 7 15 0 9 9 9 9 2
11 9 13 9 7 9 9 11 11 11 1 2
14 9 1 15 15 9 2 9 7 9 13 9 0 9 2
6 11 13 3 0 9 2
30 9 4 13 9 9 3 9 2 9 12 13 0 9 9 13 3 12 2 9 12 3 12 12 7 9 12 3 12 12 2
12 9 9 9 4 13 0 9 13 12 9 1 2
13 9 13 11 9 7 15 4 13 9 11 9 9 2
4 11 9 13 9
6 11 9 4 13 9 2
20 9 12 13 2 2 11 2 2 9 11 11 2 13 9 4 3 13 3 9 2
18 9 9 9 13 11 9 2 15 13 13 0 9 9 13 9 9 9 2
13 9 11 11 13 0 9 13 9 3 12 9 9 2
11 9 9 13 0 0 11 11 11 11 11 2
20 9 13 9 13 0 9 1 0 3 0 9 9 2 15 15 13 9 11 11 2
10 15 9 13 3 4 13 0 0 9 2
17 0 9 11 11 0 9 7 0 9 9 11 11 13 15 0 9 2
18 15 9 7 9 13 0 9 13 2 16 15 9 13 3 9 0 9 2
5 11 13 9 9 9
11 9 0 11 13 13 9 9 13 9 9 2
19 0 11 9 13 9 13 9 2 3 9 2 9 2 9 2 9 7 9 2
25 3 9 4 13 11 0 13 9 2 11 9 13 9 2 7 13 3 9 9 7 15 1 13 9 2
14 9 9 13 11 11 11 1 0 9 4 13 0 9 2
15 3 11 9 9 13 9 13 0 7 0 9 13 3 13 2
5 9 13 9 3 2
29 11 11 2 11 13 9 11 11 11 13 15 2 16 11 13 9 13 7 0 9 13 0 9 15 9 16 9 9 2
28 11 0 9 9 11 11 13 0 2 16 9 15 13 13 15 9 9 4 13 13 2 3 0 15 0 9 13 2
7 15 13 0 9 3 0 2
21 0 9 11 11 11 3 13 2 13 9 13 3 3 13 9 13 9 7 9 9 2
22 15 13 3 3 9 13 9 13 9 2 7 15 16 15 13 3 9 3 3 9 13 2
10 11 9 9 9 9 4 13 0 9 2
5 15 1 9 13 2
13 3 11 9 13 13 15 9 9 9 9 9 9 2
8 11 11 7 9 9 13 15 9
14 11 0 9 9 13 9 11 11 0 9 15 9 9 2
9 3 9 11 4 13 9 11 9 2
14 9 0 9 11 11 1 11 13 0 9 9 7 9 2
11 11 7 9 11 4 13 3 9 11 9 2
18 11 4 3 3 13 11 9 9 9 2 9 0 11 11 7 9 9 2
28 9 9 11 13 9 9 11 13 2 15 15 13 2 2 11 11 15 9 13 0 9 7 9 13 3 13 9 2
7 9 13 0 9 9 2 2
6 9 13 9 9 9 2
27 9 11 1 0 9 9 9 13 9 7 9 4 13 9 9 3 16 13 13 15 15 13 0 9 9 0 2
16 11 1 2 11 11 4 9 9 7 9 13 15 9 9 2 2
22 11 13 2 16 9 0 9 13 13 9 2 15 9 11 13 13 13 9 13 13 9 2
12 9 9 13 15 4 13 9 9 7 9 13 2
11 11 1 9 9 9 1 4 13 15 9 2
24 11 13 9 9 3 15 2 13 15 4 13 15 9 9 7 16 15 4 13 9 3 9 1 2
20 2 13 15 0 2 16 13 13 9 2 15 9 9 13 2 2 11 13 11 2
19 11 11 1 15 4 13 12 9 9 9 13 9 2 7 13 4 15 13 2
15 11 11 1 11 4 13 15 9 2 15 13 0 9 9 2
3 9 13 9
12 11 11 11 13 9 0 9 13 9 9 9 2
10 9 4 13 9 12 1 3 12 9 2
5 9 12 9 13 2
16 9 4 13 3 12 9 2 7 15 1 4 4 13 3 9 2
13 11 9 4 13 3 12 9 15 1 16 9 13 2
9 1 0 9 0 9 13 0 9 2
7 3 9 13 0 9 9 2
5 11 7 11 0 9
18 11 11 2 9 2 7 11 11 2 9 2 13 0 9 11 9 9 2
11 12 9 9 13 9 9 7 9 13 3 2
13 9 9 13 9 7 9 2 7 3 13 0 9 2
18 15 9 13 13 0 9 13 2 15 9 15 9 4 13 0 9 1 2
48 2 15 4 3 13 2 16 15 13 0 9 11 11 12 9 13 7 9 11 13 13 9 2 9 2 15 1 4 13 9 7 9 7 13 0 3 7 3 7 9 3 13 0 0 2 11 13 2
7 15 13 13 11 9 11 2
11 11 3 13 11 9 9 0 2 0 0 2
7 9 13 11 13 11 9 2
13 9 15 13 15 9 2 16 11 2 13 13 2 2
30 2 13 2 13 9 11 13 2 2 2 9 11 13 13 13 2 7 2 9 11 13 3 13 2 13 15 11 13 9 2
14 11 13 9 7 15 9 3 3 3 13 9 0 9 2
15 2 13 13 2 16 9 13 12 2 2 7 9 13 12 2
19 2 3 2 15 13 2 16 15 13 0 7 0 2 11 13 13 11 9 2
28 9 11 13 13 13 2 16 13 13 11 2 11 13 7 13 2 16 9 13 9 13 2 16 13 11 13 9 2
10 15 9 13 13 9 9 0 9 9 2
22 11 13 13 9 9 2 15 13 15 13 9 11 2 16 15 9 9 13 4 13 0 2
21 11 3 13 13 9 2 15 13 11 13 9 11 2 13 15 9 4 13 15 9 2
7 11 2 9 7 9 13 11
15 9 9 9 11 11 4 13 3 9 9 9 9 13 9 2
13 15 13 2 16 11 4 13 0 11 9 7 9 2
9 3 11 13 9 9 13 9 1 2
14 3 15 13 2 16 9 9 4 13 15 9 9 9 2
16 15 15 3 13 9 9 13 9 2 7 13 3 13 0 9 2
7 11 13 11 3 12 12 9
15 9 9 4 13 2 16 9 4 13 11 3 12 12 9 2
13 3 9 4 13 3 2 16 11 7 11 13 9 2
12 11 4 13 3 12 12 9 15 9 9 12 2
4 11 9 9 13
13 11 11 11 9 13 9 12 9 9 12 9 12 2
24 11 11 13 9 9 12 9 2 15 9 15 4 4 13 4 13 12 9 9 11 9 9 1 2
17 13 0 2 16 9 9 13 3 11 11 9 7 15 9 9 13 2
7 0 9 13 3 11 9 2
7 11 11 13 15 9 13 2
7 15 13 3 13 0 9 2
7 9 13 12 9 9 0 2
7 9 13 15 7 13 9 2
12 11 1 11 11 13 0 9 9 12 9 12 2
12 15 1 11 11 9 4 13 12 9 9 12 2
3 11 11 9
15 11 9 0 9 11 11 2 12 2 4 13 0 9 9 2
13 9 13 15 11 9 2 12 2 13 13 0 9 2
8 9 11 13 9 0 9 1 2
13 3 9 11 11 13 0 9 13 9 9 12 9 2
18 11 13 4 3 13 9 13 9 2 16 9 1 3 15 0 9 13 2
14 9 4 3 13 9 2 15 4 13 3 13 3 3 2
4 11 9 9 9
13 11 9 1 15 13 13 3 13 9 9 0 9 2
16 9 13 11 9 9 9 12 9 1 2 3 9 13 12 9 2
15 9 13 3 0 9 9 2 15 1 9 13 3 12 9 2
8 9 15 13 0 9 11 9 2
10 9 13 13 13 9 1 0 0 9 2
11 3 13 11 13 12 12 9 9 11 1 2
9 9 13 9 13 11 0 9 9 2
7 11 13 9 0 9 9 2
14 3 0 9 13 11 9 2 3 15 9 13 9 13 2
15 11 4 0 9 9 13 0 9 0 9 3 11 7 11 2
18 9 0 9 4 13 0 0 0 9 9 9 7 11 13 0 9 9 2
9 9 0 9 4 3 13 0 9 2
21 11 9 4 13 3 0 11 9 11 5 11 2 16 15 13 13 13 13 9 3 2
25 11 0 9 11 4 13 9 9 2 15 1 9 9 11 11 4 13 9 16 0 9 13 9 3 2
3 11 13 9
8 9 11 11 4 13 9 9 2
9 15 13 3 11 0 9 11 9 2
7 3 11 11 13 9 9 2
10 9 9 11 11 13 9 3 9 9 2
13 15 13 12 9 7 13 12 9 9 11 11 11 2
15 11 13 12 0 9 2 7 13 12 9 9 9 9 11 2
13 9 13 9 9 1 2 7 9 13 3 0 9 2
13 11 13 12 9 2 7 13 0 9 7 13 9 2
15 3 9 11 11 13 11 9 13 9 9 12 9 9 9 2
8 0 11 11 13 9 12 9 2
15 0 13 11 11 11 13 12 9 7 9 13 11 12 9 2
4 11 0 9 13
11 11 11 9 4 13 13 9 13 0 9 2
9 9 11 9 4 13 11 9 9 2
9 9 4 13 12 9 9 12 9 2
4 11 9 9 13
15 9 4 13 9 9 2 15 13 11 9 9 12 12 9 2
11 9 13 3 9 0 9 9 12 12 9 2
11 0 9 9 9 4 13 9 3 15 9 2
20 9 13 2 16 9 9 9 13 0 9 2 0 9 11 11 9 13 3 9 2
18 11 13 3 11 11 9 9 2 7 15 13 13 3 13 9 9 1 2
13 11 9 13 4 13 15 1 16 15 13 9 12 2
5 9 13 0 9 9
13 12 0 9 9 13 0 9 11 13 9 0 9 2
11 9 13 1 9 2 15 15 13 9 3 2
16 9 1 9 13 9 1 9 13 15 9 2 15 4 13 9 2
13 9 13 3 0 9 2 7 9 13 3 15 13 2
8 0 9 1 15 3 4 13 2
11 9 12 2 0 11 13 9 2 4 13 2
14 9 13 9 7 13 9 2 13 15 4 3 4 13 2
7 9 13 3 12 0 9 2
5 9 13 13 11 9
14 0 9 12 11 11 11 11 9 9 13 11 9 11 2
7 9 0 9 7 9 13 2
12 12 9 4 13 2 12 15 13 13 0 9 2
5 9 13 9 11 9
25 9 9 13 9 13 3 9 11 11 2 9 2 9 2 15 13 15 9 13 3 12 9 0 9 2
19 9 7 9 2 15 0 9 13 3 12 12 9 2 13 9 3 0 9 2
17 3 9 13 12 9 9 7 15 13 3 15 9 2 15 13 9 2
20 9 11 11 13 9 13 15 9 13 9 15 2 16 11 9 13 9 15 9 2
11 0 9 13 9 1 9 2 9 7 9 2
6 9 13 9 9 12 2
7 0 9 9 13 9 3 2
19 11 9 9 11 11 13 13 9 2 9 2 2 16 3 11 13 15 9 2
16 9 9 9 2 11 11 9 11 11 13 9 13 0 9 9 2
26 15 9 13 0 9 13 2 13 11 0 9 9 2 7 13 0 9 15 2 13 15 11 9 0 9 2
17 9 9 9 11 11 13 2 16 9 13 0 9 9 9 9 9 2
12 11 9 11 11 13 9 9 13 11 9 9 2
13 15 13 2 16 11 9 3 9 13 15 16 9 2
20 15 1 0 9 13 11 13 9 15 9 2 15 13 15 1 4 11 9 13 2
7 9 4 13 15 9 1 2
17 9 13 9 9 1 15 2 13 9 9 7 9 7 13 15 9 2
14 9 13 9 13 0 2 7 9 4 13 3 9 9 2
5 9 11 13 3 11
19 9 12 13 2 16 9 7 9 13 11 13 9 3 13 9 0 9 9 2
6 0 9 9 13 11 2
8 9 4 13 9 11 9 1 2
4 11 13 11 9
12 11 11 11 13 9 9 9 9 9 11 11 2
15 11 11 11 13 0 1 11 11 11 2 15 13 9 0 2
7 11 13 9 3 9 1 2
25 11 13 3 9 0 2 7 13 0 16 0 9 1 3 0 13 11 11 13 0 9 7 13 0 2
14 9 12 15 9 2 11 11 7 11 11 13 0 9 2
12 11 0 9 13 3 9 0 0 9 13 9 2
15 3 11 11 2 11 11 7 11 11 13 3 9 3 3 2
5 2 13 3 0 2
11 13 3 9 11 2 7 3 15 13 3 2
19 11 0 9 1 15 13 0 9 15 9 2 15 9 4 13 2 11 13 2
15 2 3 15 0 13 2 13 15 0 9 4 9 13 9 2
11 15 1 4 13 9 7 3 15 13 9 2
17 3 13 13 3 9 7 3 9 13 7 9 13 0 2 11 13 2
4 11 11 11 9
14 11 11 11 13 0 11 9 15 13 3 9 13 9 2
15 15 13 3 3 11 3 0 9 7 12 15 0 9 9 2
12 3 3 9 13 9 12 9 13 11 0 9 2
22 9 12 15 13 13 3 9 11 11 7 11 11 2 15 13 9 0 9 0 9 1 2
11 9 9 3 13 15 13 0 9 9 1 2
11 11 9 9 9 13 15 9 16 3 11 2
15 15 13 3 13 9 0 9 2 16 9 9 13 0 11 2
18 9 13 9 9 11 11 11 13 12 12 0 9 15 13 12 12 11 2
15 0 9 9 4 13 9 1 3 9 2 7 4 13 9 2
13 3 7 0 2 7 0 9 9 9 4 13 0 2
25 15 1 9 4 13 3 9 12 2 3 9 13 3 11 11 9 7 13 15 3 9 9 12 9 2
9 9 1 9 11 11 13 9 13 2
18 9 9 1 9 13 13 9 13 15 9 2 7 13 9 9 13 9 2
15 9 9 13 9 4 3 13 13 9 9 13 9 15 1 2
12 12 9 0 3 13 9 11 11 11 9 1 2
12 11 11 11 1 4 12 9 9 1 13 9 2
34 9 13 11 11 9 13 11 11 2 11 11 7 11 11 2 7 3 9 11 11 2 15 4 9 13 11 11 9 13 11 11 11 9 2
9 9 13 9 9 9 7 9 9 2
20 3 9 9 13 2 16 9 13 12 12 9 2 12 12 9 2 13 0 9 2
10 11 1 9 4 3 13 12 9 9 2
12 11 11 9 1 9 13 9 13 3 12 9 2
17 9 11 4 13 13 9 12 9 2 12 9 7 12 9 0 9 2
10 9 15 13 9 13 9 12 12 9 2
7 15 9 13 0 11 9 2
33 7 11 2 7 11 11 11 9 9 13 2 16 1 15 15 13 9 9 3 15 13 13 9 2 16 15 9 4 13 0 0 9 2
5 12 12 11 13 9
14 11 9 13 13 12 12 9 7 9 9 13 9 1 2
22 9 4 13 9 11 7 11 7 15 4 13 9 9 2 16 9 7 9 4 13 9 2
8 9 13 9 12 7 0 9 2
11 11 9 11 11 9 11 4 13 9 0 9
12 11 9 11 11 9 11 4 13 9 0 9 2
18 15 13 3 13 9 0 9 7 15 4 13 13 0 9 9 9 9 2
12 9 12 13 9 0 9 13 0 9 9 9 2
20 3 15 0 0 9 3 11 2 11 2 11 2 11 2 11 7 11 13 0 2
9 15 15 9 13 3 9 0 9 2
13 15 9 13 1 12 9 12 2 7 13 15 9 2
59 11 2 15 3 0 11 9 2 13 3 0 9 13 9 2 7 13 0 2 16 13 9 2 9 13 11 11 13 9 2 16 15 1 0 9 9 12 13 9 2 15 13 9 12 12 5 15 9 2 13 3 0 9 12 5 15 13 9 2
10 11 9 11 13 3 3 11 0 9 2
29 0 9 9 13 11 2 15 9 9 11 11 13 12 5 13 9 2 16 15 0 9 0 11 11 13 9 12 5 2
22 9 9 4 13 7 0 11 11 11 2 12 5 2 7 9 9 2 12 5 2 9 2
8 11 13 11 7 13 11 9 9
18 11 0 9 11 11 4 13 9 7 13 9 11 11 11 11 11 9 2
16 11 13 11 13 0 9 11 7 2 11 13 13 9 9 2 2
8 11 13 15 0 9 9 9 2
10 11 13 3 11 13 3 11 9 9 2
13 11 1 11 13 9 11 4 2 13 2 11 1 2
13 15 13 13 11 9 11 11 7 13 15 0 9 2
26 11 1 11 4 13 11 9 11 11 9 1 2 13 9 0 9 7 13 9 7 13 0 7 9 9 2
13 11 11 2 13 12 2 13 11 0 9 9 12 2
9 15 13 11 9 9 0 9 9 2
4 11 13 11 9
12 9 11 11 13 3 11 9 9 12 9 12 2
16 2 3 15 4 13 9 7 4 13 9 2 13 11 9 9 2
12 9 11 11 13 9 13 0 12 9 9 11 2
16 2 11 13 0 9 2 7 13 13 15 3 3 2 13 11 2
11 0 9 13 12 9 1 11 0 11 11 2
12 11 11 11 13 9 0 7 0 9 0 9 2
21 9 13 11 0 11 11 9 2 13 9 13 9 1 0 11 11 9 15 9 9 2
17 9 0 9 9 13 3 12 9 2 15 13 9 3 3 12 9 2
3 9 12 9
10 9 4 13 9 12 0 9 7 9 2
10 2 0 9 2 9 9 11 13 12 2
17 2 0 9 2 11 2 11 2 11 0 9 9 13 0 11 9 2
7 2 0 9 2 9 11 2
10 9 0 9 13 11 15 13 12 9 2
8 9 3 13 11 3 12 9 2
27 9 9 3 9 13 12 9 2 7 15 13 3 9 13 9 3 11 1 7 13 9 9 9 9 11 11 2
20 2 0 9 2 9 11 13 0 11 9 9 9 13 11 9 11 11 9 11 2
10 2 0 9 2 11 13 3 0 9 2
13 15 11 9 9 13 2 16 9 13 4 13 9 2
13 9 13 9 13 13 0 9 9 3 9 12 9 2
10 13 3 9 11 9 11 2 0 9 2
11 2 0 9 2 0 9 13 11 9 11 2
7 13 3 11 9 11 9 2
17 2 0 9 2 11 7 11 13 11 9 2 15 13 12 9 0 2
9 2 0 9 2 11 9 13 11 2
18 2 0 9 2 11 11 13 9 9 13 0 9 9 3 9 9 9 2
12 2 0 9 2 11 11 13 11 9 0 9 2
20 2 0 9 2 11 11 9 12 11 13 9 13 9 13 3 9 7 13 9 2
5 12 9 13 9 2
7 9 9 0 9 1 9 2
15 15 9 1 9 13 9 9 9 2 7 3 11 13 9 2
8 9 9 13 9 0 0 9 2
6 3 9 13 11 1 2
14 9 11 11 1 9 13 15 9 13 3 0 16 3 2
17 9 4 13 9 3 2 7 9 4 3 13 2 3 13 9 13 2
6 9 9 13 9 9 2
9 11 9 13 3 11 7 11 9 2
8 3 0 9 13 11 7 11 2
11 11 1 9 13 9 3 0 9 13 11 2
14 11 11 9 7 0 11 13 9 2 15 9 4 13 2
16 16 11 9 13 3 9 15 9 9 2 13 9 9 0 9 2
7 9 9 13 9 3 9 2
14 0 9 9 13 13 2 16 15 9 13 3 12 9 2
24 16 9 13 0 0 2 13 0 9 9 2 16 9 13 3 3 13 15 7 9 13 3 9 2
15 11 1 9 3 13 11 3 9 9 2 3 3 3 3 2
4 3 2 9 12
11 2 9 13 9 3 0 9 9 12 9 2
14 15 13 0 11 9 3 1 0 9 13 9 9 3 2
5 2 9 13 9 2
14 11 9 9 11 11 13 0 9 13 9 9 11 11 2
30 13 9 2 15 9 0 9 11 11 11 4 13 11 9 13 2 11 13 9 11 11 13 15 9 7 13 9 9 9 2
7 11 9 13 3 13 9 2
9 11 11 13 3 4 13 13 9 2
8 2 11 9 9 12 12 9 2
17 11 11 9 11 11 13 0 9 12 12 9 9 11 11 9 9 2
9 9 13 11 9 11 13 9 11 2
5 9 13 9 9 9
19 3 12 9 9 4 13 11 13 11 9 9 2 15 9 13 0 9 9 2
9 9 13 11 3 15 9 13 9 2
13 9 1 0 9 9 13 3 12 9 9 9 13 2
15 9 1 9 9 4 13 12 9 9 12 9 9 12 1 2
16 0 9 9 13 2 16 9 9 13 12 9 2 9 2 9 2
19 9 13 0 2 16 11 9 13 9 9 12 9 9 12 9 9 12 1 2
12 9 9 13 2 13 9 9 13 3 12 5 2
9 9 1 9 13 3 3 0 9 2
17 9 13 9 13 2 16 11 9 9 13 0 7 16 0 9 13 2
13 11 9 13 2 16 0 9 4 13 9 12 11 2
14 0 9 13 9 13 11 9 9 7 9 12 0 9 2
9 12 9 0 9 9 4 13 9 5
3 0 9 11
23 11 11 4 13 0 9 16 5 0 9 2 9 5 2 13 3 9 1 9 9 13 9 2
13 9 13 9 11 11 1 12 9 7 12 9 9 2
18 9 13 9 1 9 4 13 12 9 7 9 9 13 13 3 12 9 2
15 9 11 11 1 9 4 13 9 3 1 15 9 3 9 2
7 9 5 13 9 11 1 2
16 11 9 9 11 11 4 13 9 11 9 11 11 9 9 1 2
3 11 0 9
14 3 12 9 4 13 9 12 9 13 9 11 13 11 2
6 3 13 13 3 12 2
21 9 13 9 9 9 9 13 11 11 9 2 16 9 13 9 13 9 9 0 9 2
15 16 9 9 11 13 11 11 13 9 2 13 9 9 0 2
14 0 9 4 13 9 13 7 13 7 13 9 7 9 2
4 9 13 9 11
8 0 0 9 13 9 11 9 2
17 15 9 13 12 9 2 12 9 7 12 9 9 2 4 13 9 2
7 9 9 13 13 3 9 2
3 11 9 13
11 3 9 9 13 0 3 12 12 9 9 2
8 9 9 4 3 13 12 9 2
16 3 9 9 13 3 9 9 2 16 0 0 9 9 13 9 2
32 3 0 9 11 0 9 3 9 11 2 9 11 7 9 11 13 15 1 9 12 7 15 4 13 3 11 9 3 13 9 9 2
22 3 9 11 2 15 13 3 9 2 7 4 13 0 9 13 9 2 13 9 9 12 2
9 11 13 0 7 0 9 3 11 2
7 11 13 3 11 13 9 2
4 9 13 9 9
4 11 2 11 2
32 11 11 2 11 11 11 2 11 11 11 11 11 7 11 11 11 13 3 11 9 9 1 9 13 0 11 11 12 12 9 9 2
14 11 4 13 9 13 12 9 2 7 15 13 13 9 2
20 9 13 11 15 0 9 9 2 16 3 9 4 3 13 9 9 0 9 0 2
21 11 1 9 4 3 13 9 9 9 2 16 4 3 13 9 9 0 9 13 1 2
14 11 9 13 0 9 1 2 7 9 9 13 13 9 2
3 11 13 2
16 9 4 13 2 16 11 9 13 9 0 9 9 12 11 9 2
16 9 13 13 9 0 9 9 2 7 9 9 9 13 9 9 2
7 11 11 13 11 9 12 2
32 0 9 11 11 1 0 11 11 9 9 13 11 11 11 7 11 4 13 9 11 11 1 2 15 15 13 9 9 1 0 9 2
16 11 11 1 11 4 13 3 12 12 9 7 12 12 9 13 2
20 3 9 9 9 1 13 13 9 9 9 1 2 16 11 7 11 9 13 9 2
12 0 9 1 15 13 9 9 2 16 9 13 2
19 0 11 11 13 9 0 9 9 7 13 15 11 11 11 9 7 9 13 2
8 3 9 3 13 9 11 11 2
10 11 11 3 9 1 3 4 13 9 2
13 11 13 11 9 12 13 3 9 0 7 0 9 2
4 11 0 9 9
14 9 11 4 13 13 0 9 0 7 3 13 9 9 2
16 9 13 9 12 13 0 9 9 9 13 9 7 0 0 9 2
16 9 4 13 9 0 7 3 13 9 7 9 4 13 9 3 2
8 11 9 13 12 12 9 9 2
11 9 13 13 13 9 7 9 9 7 9 2
6 9 9 13 11 11 2
4 0 9 13 9
8 0 0 9 11 11 13 9 2
16 11 9 13 0 11 11 13 9 0 9 12 7 13 0 9 2
12 9 9 13 9 9 2 15 9 3 13 11 2
12 9 13 9 9 7 0 11 9 9 12 9 2
8 15 13 3 7 12 9 9 2
10 9 4 3 13 9 11 9 0 9 2
17 15 4 13 15 9 7 9 9 7 13 12 9 9 11 9 9 2
8 9 1 13 4 13 15 9 2
5 9 13 13 3 2
12 9 11 11 13 9 13 9 7 9 9 9 2
4 9 13 9 13
22 0 9 7 9 2 9 9 11 11 11 11 2 12 2 13 13 9 13 11 12 9 2
19 9 7 9 9 13 11 13 3 9 9 7 13 9 9 13 9 9 13 2
13 11 13 4 13 0 9 2 7 15 13 9 3 2
7 11 9 9 13 3 0 2
26 15 4 9 3 13 9 9 9 2 7 15 9 15 13 4 9 13 2 3 16 15 9 13 13 13 2
15 13 9 11 13 0 15 13 9 9 7 13 15 0 9 2
10 11 1 11 4 13 9 13 9 9 2
7 2 15 13 4 13 9 2
6 15 15 13 9 9 2
13 9 9 11 7 11 9 13 3 3 9 13 9 2
8 11 1 15 13 9 0 9 2
29 9 11 11 1 11 13 4 3 13 2 7 15 15 4 12 9 3 13 9 11 2 7 15 9 15 13 4 13 2
16 9 11 1 13 13 0 2 16 9 13 9 9 7 9 9 2
32 11 9 1 9 13 15 9 9 16 9 13 12 9 2 3 3 12 9 13 11 13 3 15 9 2 15 13 9 13 0 9 2
3 11 9 0
14 12 12 9 11 13 3 12 12 0 2 13 9 9 2
5 9 13 12 9 2
15 3 3 11 9 9 13 0 9 4 13 12 12 9 9 2
7 0 9 9 13 12 9 2
10 11 9 1 9 9 13 9 9 1 2
9 11 13 0 9 3 9 9 1 2
6 9 9 4 13 3 2
8 9 11 9 2 0 9 13 9
6 11 11 13 9 11 2
5 11 9 13 9 2
6 11 13 13 3 0 2
13 15 13 3 9 2 15 1 15 9 9 13 0 2
17 11 13 0 9 9 9 11 11 7 15 13 9 2 3 15 13 2
13 9 13 13 9 2 16 15 4 13 1 9 9 2
13 11 4 13 0 9 11 9 9 9 2 12 2 2
9 11 13 9 12 11 9 9 9 2
9 3 11 13 3 0 9 13 9 2
11 11 13 11 11 11 0 9 9 9 12 2
5 0 9 13 11 9
17 0 9 4 13 9 2 15 13 9 0 9 13 15 9 11 11 2
6 9 0 13 3 9 2
13 11 9 9 11 1 9 11 11 13 9 13 3 2
14 2 9 7 9 13 3 0 9 16 0 2 13 11 2
8 11 1 9 13 13 9 9 2
8 9 13 13 9 13 9 13 2
5 9 12 9 1 2
12 9 0 9 7 9 9 4 9 1 13 9 2
9 9 1 13 3 12 9 13 9 2
24 11 11 11 7 9 2 9 0 9 2 13 0 9 12 11 7 11 9 13 11 9 9 11 2
16 11 11 11 13 9 13 13 3 3 9 9 7 3 9 13 2
15 12 9 1 13 9 4 13 7 13 12 9 9 0 9 2
13 11 11 11 4 9 1 13 9 0 0 9 9 2
22 0 9 11 11 1 15 0 9 4 12 9 13 13 3 0 2 16 15 13 11 3 2
9 11 13 9 1 13 3 11 9 2
10 11 11 11 13 9 1 11 9 0 2
8 9 13 3 13 13 11 9 2
12 11 4 11 13 1 13 11 9 13 0 9 2
8 11 1 15 13 3 13 9 2
15 11 13 11 1 3 13 13 9 15 0 9 9 13 9 2
20 3 15 9 13 9 13 0 0 9 9 13 0 7 16 11 9 13 13 9 2
4 11 13 11 11
22 0 9 12 9 11 11 13 3 13 11 11 2 15 9 13 9 0 0 9 9 11 2
6 9 13 3 12 9 2
3 11 13 3
13 11 7 11 9 4 3 9 13 9 0 11 9 2
11 3 3 11 9 4 13 9 0 0 9 2
12 11 4 13 0 9 7 13 13 9 0 9 2
25 0 11 9 9 13 0 9 7 9 9 2 16 12 9 1 11 13 11 9 13 12 9 9 11 2
8 9 11 13 9 0 9 11 2
16 3 7 9 11 9 2 7 11 9 9 13 11 9 9 12 2
9 9 1 11 9 13 9 11 9 2
14 3 11 13 9 9 2 16 9 13 11 7 11 9 2
6 9 13 3 9 9 2
14 3 4 13 2 16 0 9 13 4 13 15 9 1 2
35 15 13 13 0 0 9 16 11 9 11 11 13 2 2 7 15 2 16 0 13 15 2 0 9 2 15 9 13 3 2 13 9 15 3 2
5 9 13 13 9 11
13 9 13 9 13 13 9 15 9 9 11 11 9 2
13 9 9 13 13 9 2 7 15 13 3 9 13 2
12 9 13 9 2 16 9 13 9 9 13 9 2
10 9 13 9 9 1 7 13 3 9 2
9 9 13 9 7 13 9 13 3 2
5 9 9 13 9 9
19 9 2 5 2 0 9 11 9 7 9 9 9 0 9 4 13 0 9 2
25 0 11 2 15 13 9 9 9 7 9 2 13 15 9 9 12 9 1 11 9 3 12 12 9 2
9 9 13 9 0 9 15 9 9 2
14 0 9 13 11 2 7 3 15 13 12 5 0 9 2
16 11 5 13 12 5 9 9 2 11 12 5 7 11 12 5 2
22 0 9 9 9 13 11 2 15 15 13 9 9 12 9 7 9 3 12 9 15 9 2
10 0 9 9 11 13 3 0 1 9 2
12 15 0 9 9 13 11 12 9 11 12 9 2
16 11 2 11 2 13 3 0 0 2 3 11 2 11 7 11 2
10 11 9 4 13 3 0 3 1 11 2
17 9 13 3 15 2 16 9 13 9 11 2 15 13 12 9 9 2
14 9 13 3 2 16 15 0 9 13 9 9 9 9 2
6 11 13 3 9 9 2
17 9 9 13 9 1 0 0 11 2 15 15 13 3 12 5 9 2
10 11 7 11 9 13 9 12 9 1 2
19 9 9 3 9 13 0 9 2 16 3 9 9 13 12 5 0 9 9 2
8 3 9 0 9 13 12 5 2
1 9
10 2 0 9 12 2 11 7 11 0 9
13 2 0 9 12 2 9 11 0 9 9 11 11 9
10 2 0 9 12 2 9 13 13 9 9
11 2 0 9 12 2 11 9 13 9 15 9
8 2 0 9 12 2 11 12 9
16 2 0 9 12 2 11 9 12 12 9 9 2 9 13 11 1
9 2 0 9 12 2 9 13 13 11
12 2 0 9 12 2 11 11 9 0 9 9 1
11 2 0 9 12 2 11 9 11 11 11 9
15 2 0 9 12 2 11 11 7 11 11 9 9 13 9 9
9 2 0 9 12 2 9 2 9 11
12 2 0 9 12 2 11 13 9 2 13 0 9
13 2 0 9 12 2 9 13 11 2 9 13 9 9
11 2 0 9 12 2 9 13 9 9 11 9
14 2 0 9 12 2 11 13 9 9 2 11 13 9 9
11 2 0 9 12 2 9 13 12 9 9 0
10 2 0 9 12 2 11 11 9 13 9
10 2 0 9 12 2 9 13 0 11 9
8 2 0 9 12 2 11 9 11
10 2 0 9 12 2 11 13 9 11 9
12 2 0 9 12 2 11 9 0 9 3 3 9
13 2 0 9 12 2 3 11 9 13 11 11 13 9
12 2 0 9 12 2 11 13 11 3 12 12 9
10 2 0 9 12 2 11 13 13 11 13
13 2 0 9 12 2 11 13 0 7 9 9 9 11
8 2 0 9 12 2 9 9 11
10 2 0 9 12 2 9 13 11 11 9
10 2 0 9 12 2 11 13 9 13 13
11 2 0 9 12 2 11 11 13 9 9 9
8 2 0 9 12 2 11 9 11
8 2 0 9 12 2 9 13 11
10 2 0 9 12 2 9 11 13 3 11
15 2 0 9 12 2 11 13 11 3 12 12 9 12 9 9
8 2 0 9 12 2 11 13 9
11 2 0 9 12 2 9 7 11 11 13 9
7 2 0 9 12 2 9 11
8 2 0 9 12 2 9 9 13
11 2 0 9 12 2 11 13 13 9 11 9
8 2 0 9 12 2 9 13 9
10 2 0 9 12 2 9 13 9 9 11
8 2 0 9 12 2 11 9 12
11 2 0 9 12 2 9 11 13 9 11 11
10 2 0 9 12 2 11 11 13 11 9
11 2 0 9 12 2 11 2 9 0 9 1
12 2 0 9 12 2 9 9 7 9 13 9 9
13 2 0 9 12 2 0 9 2 11 11 9 9 12
10 2 0 9 12 2 11 0 9 9 12
11 2 0 9 12 2 0 9 11 9 9 13
7 2 0 9 12 2 9 12
10 2 0 9 12 2 9 9 9 1 11
15 2 0 9 12 2 11 13 9 3 2 11 9 9 9 0
14 2 0 9 12 2 11 9 11 9 13 13 9 0 9
8 2 0 9 12 2 11 11 9
8 2 0 9 12 2 11 11 9
13 2 0 9 12 2 11 11 7 9 9 13 9 9
14 2 0 9 12 2 2 12 9 9 2 13 3 11 9
10 2 0 9 12 2 9 13 9 11 9
10 2 0 9 12 2 11 11 13 9 9
12 2 0 9 12 2 9 2 15 13 12 9 9
13 2 0 9 12 2 11 2 9 13 13 13 11 11
11 2 0 9 12 2 11 11 9 9 0 9
9 2 0 9 12 2 11 9 12 9
10 2 0 9 12 2 11 7 11 9 9
9 2 0 9 12 2 3 2 9 12
10 2 0 9 12 2 9 11 9 9 9
9 2 0 9 12 2 11 9 13 13
10 2 0 9 12 2 9 0 9 11 9
12 2 0 9 12 2 11 2 9 9 4 13 9
8 2 0 9 12 2 11 9 9
12 2 0 9 12 2 11 2 0 9 9 0 9
9 2 0 9 12 2 3 2 9 12
10 2 0 9 12 2 9 13 11 9 9
10 2 0 9 12 2 9 13 11 9 1
9 2 0 9 12 2 3 2 9 12
6 0 9 13 9 11 9
18 0 9 13 9 0 11 1 2 16 9 13 9 11 9 11 11 11 2
16 9 1 13 9 13 9 9 9 7 9 13 12 9 7 9 2
8 9 13 12 1 9 3 11 2
6 9 9 9 13 9 2
12 15 13 11 0 9 2 15 9 13 1 9 2
4 9 9 13 11
13 11 11 9 0 9 2 11 11 2 9 13 11 2
8 11 4 13 13 12 9 3 2
7 9 13 9 9 0 9 2
13 9 1 11 4 13 9 2 7 13 13 3 9 2
11 11 11 13 0 9 0 9 2 11 11 2
16 2 15 9 1 15 13 15 9 3 2 2 13 9 11 11 2
17 11 9 2 11 11 2 13 9 0 9 2 15 13 9 13 9 2
12 9 4 13 9 3 12 9 1 2 1 9 2
12 15 1 9 13 9 13 9 7 13 15 3 2
5 11 13 9 11 11
18 11 9 9 9 11 11 4 13 3 9 11 11 9 11 11 0 9 2
7 15 9 13 3 0 9 2
11 15 11 15 9 0 9 9 13 0 9 2
28 9 1 7 11 7 11 13 15 3 12 9 9 9 7 0 13 11 11 2 15 13 9 1 12 9 13 9 2
10 9 4 13 16 11 13 11 13 9 2
16 3 3 9 12 13 9 9 11 4 13 0 9 11 11 9 2
6 9 9 13 3 13 3
21 9 9 3 13 3 2 16 12 9 13 9 13 0 11 9 9 9 13 13 9 2
11 9 13 9 2 7 9 13 4 13 9 2
18 13 9 11 11 13 9 13 9 13 7 9 1 13 9 9 1 9 2
7 9 1 9 13 1 9 2
17 9 9 13 9 13 9 3 2 16 15 13 9 13 15 0 9 2
11 9 13 4 13 9 2 16 9 13 9 2
8 9 11 1 15 13 13 13 2
7 15 1 9 9 13 0 2
16 11 13 9 7 9 9 2 16 15 4 4 13 9 9 9 2
19 2 15 3 13 2 13 9 13 13 15 3 2 7 15 9 4 4 13 2
11 15 4 4 13 9 2 2 13 11 2 2
8 9 13 9 9 9 13 13 2
7 0 9 9 0 3 9 12
11 0 9 9 13 9 12 0 3 9 12 2
25 9 0 9 12 13 11 9 9 2 11 2 2 16 9 12 9 4 13 12 5 13 0 9 12 2
21 9 9 9 13 3 9 12 12 12 9 2 16 9 13 3 9 12 12 12 9 2
9 9 13 0 3 9 12 0 9 2
9 9 9 4 13 3 12 0 9 2
13 3 9 4 13 9 2 15 9 4 13 0 3 2
17 15 4 13 3 11 9 9 15 4 13 9 12 5 13 0 9 2
21 11 13 9 3 12 12 9 7 3 13 12 12 9 9 2 15 15 13 9 12 2
19 3 11 13 0 9 2 15 13 12 5 2 7 11 9 13 3 12 5 2
35 3 0 9 4 13 9 3 3 9 7 11 9 9 1 9 2 15 13 13 3 11 7 11 2 4 13 9 0 9 9 1 0 11 11 2
4 11 9 9 13
12 11 0 9 9 13 9 4 13 3 12 9 2
9 9 4 13 15 9 3 12 9 2
27 9 13 9 13 9 9 9 9 11 11 2 11 11 7 11 11 7 9 11 11 2 11 11 7 11 11 2
15 9 9 13 9 11 11 2 9 9 11 7 9 11 11 2
19 15 0 9 13 9 9 13 9 9 12 7 15 13 0 9 11 9 12 2
12 11 9 13 12 0 7 9 7 9 9 13 2
9 9 13 12 2 12 7 12 9 2
6 3 0 9 13 9 2
12 3 0 3 13 9 9 9 13 9 11 11 2
6 9 13 9 9 11 9
8 9 4 13 9 11 9 9 2
20 9 4 13 12 11 11 2 9 2 9 7 13 12 9 11 11 2 9 2 2
17 15 4 13 12 9 9 13 9 2 15 13 12 5 9 13 9 2
8 11 13 9 3 3 12 9 2
8 9 13 3 12 5 9 9 2
8 9 9 13 11 9 11 11 2
11 9 9 11 11 13 13 9 11 13 9 2
14 9 9 13 3 15 9 0 16 9 9 13 9 9 2
3 9 9 9
15 11 2 11 7 11 13 9 11 9 0 9 13 9 1 2
13 9 11 11 13 9 13 0 9 11 11 3 11 2
7 11 4 3 13 9 9 2
11 9 13 0 9 2 7 15 13 9 0 2
10 11 4 13 9 11 9 13 9 9 2
14 9 9 1 9 9 9 13 11 1 13 0 9 9 2
9 13 9 13 13 9 9 13 9 2
3 11 9 1
15 0 9 9 13 9 4 13 12 0 0 9 1 13 9 2
11 0 9 13 11 7 11 13 9 9 9 2
11 11 11 13 0 9 1 9 4 13 9 2
24 12 9 11 9 13 9 9 13 0 2 7 9 4 13 13 15 2 16 9 9 4 13 9 2
7 9 13 13 9 9 9 2
23 0 9 2 11 11 2 13 9 12 9 1 11 7 11 0 9 1 15 13 3 9 9 2
20 11 9 13 9 9 13 9 11 9 2 11 2 11 2 11 7 11 9 9 2
9 3 9 13 3 11 7 11 9 2
24 9 9 13 11 7 11 0 9 2 15 3 15 9 1 4 13 3 7 13 3 3 11 9 2
23 11 9 13 0 9 13 3 13 15 0 9 16 9 9 7 15 13 13 9 13 15 9 2
28 3 15 9 15 9 13 13 3 9 2 7 0 11 9 13 0 9 9 16 9 13 13 3 0 13 9 1 2
6 9 13 9 12 9 13
15 0 9 13 9 7 13 9 13 12 9 11 11 11 9 2
16 9 0 9 9 13 9 9 7 9 9 7 3 0 9 9 2
27 9 4 13 0 9 9 1 9 0 11 11 11 11 11 9 2 15 4 11 11 1 13 9 15 9 0 2
8 9 13 13 13 9 0 9 2
9 9 9 13 15 9 0 9 9 2
22 0 9 13 3 3 2 16 0 0 9 13 9 1 9 2 16 13 13 0 9 15 2
5 15 4 13 9 2
4 11 9 9 9
16 9 9 9 13 9 9 9 3 3 9 7 9 13 11 11 2
33 0 11 4 3 3 13 9 9 2 7 9 12 15 13 11 2 8 8 8 2 9 0 9 2 8 8 2 11 11 9 13 15 2
16 15 13 9 7 9 7 13 9 3 3 9 12 12 9 9 2
16 0 9 13 3 3 2 7 3 11 9 13 4 13 15 9 2
21 11 11 1 9 1 11 9 13 0 9 9 7 9 15 13 3 9 1 9 9 2
30 9 13 3 16 15 13 9 13 11 13 9 9 7 11 9 13 15 3 13 2 16 15 4 13 13 13 9 9 1 2
8 11 13 9 9 9 15 1 2
13 9 9 13 0 9 1 13 0 11 9 15 1 2
17 9 4 3 3 3 9 13 9 13 9 9 9 13 9 9 9 2
6 11 9 9 0 12 9
18 11 9 9 13 0 12 9 7 9 9 9 13 12 9 2 13 11 2
16 9 4 13 9 9 12 12 9 7 3 9 4 13 12 9 2
23 3 9 9 13 3 9 2 16 9 13 9 12 12 12 9 7 9 3 13 12 12 9 2
16 9 12 13 12 9 3 16 0 9 2 7 13 13 12 12 2
18 9 3 13 9 12 13 12 9 7 9 9 13 3 3 12 12 9 2
22 9 13 3 11 2 11 7 11 7 12 15 9 7 11 2 16 15 3 16 12 9 2
14 12 9 3 9 13 7 3 13 9 13 11 7 11 2
5 9 9 9 1 11
13 11 9 4 9 11 1 13 9 9 1 9 1 2
16 11 1 0 9 9 4 13 3 11 2 0 9 7 9 0 2
22 9 13 0 9 13 9 2 15 3 13 9 2 11 11 2 7 2 11 11 2 1 2
3 13 15 2
7 15 13 15 3 0 9 2
6 9 1 13 13 3 2
7 9 13 9 9 13 15 2
7 9 13 13 11 13 9 2
2 15 13
10 0 9 9 13 9 9 13 0 9 2
13 13 9 9 7 9 2 3 3 10 9 3 13 2
6 15 13 13 13 9 2
5 11 13 0 9 2
2 15 1
9 9 13 13 9 0 9 7 9 2
5 11 13 9 9 2
7 13 13 12 9 9 1 2
21 13 15 16 15 3 11 13 3 13 15 3 3 3 3 16 13 15 13 9 9 2
9 3 15 16 9 13 2 15 13 9
7 15 13 16 13 13 3 2
14 3 10 9 15 2 15 13 2 13 8 2 3 11 2
3 13 13 2
19 9 9 13 0 9 2 16 3 0 9 13 3 9 7 3 10 9 3 2
15 11 13 2 13 13 15 9 7 13 9 10 9 9 9 2
8 16 2 13 16 9 3 7 9
5 13 11 3 3 2
5 9 13 12 9 2
5 0 9 13 0 9
3 8 8 2
28 2 10 9 9 3 9 13 3 3 2 16 3 13 15 13 10 9 2 16 15 13 13 3 13 9 9 2 2
10 13 9 7 13 9 2 15 9 13 2
4 13 13 13 2
9 3 13 13 2 3 0 9 15 2
4 13 3 9 2
7 15 13 9 13 13 9 2
3 13 3 9
3 15 13 15
16 3 13 2 13 7 13 0 2 3 13 9 9 7 13 9 2
4 13 3 9 2
5 6 6 10 9 2
3 6 3 3
15 15 13 0 2 7 16 9 13 9 2 15 0 9 13 2
14 9 13 0 13 3 13 2 12 9 2 13 9 3 2
3 13 9 9
3 15 13 11
4 0 7 0 2
3 9 13 2
6 9 13 0 7 0 2
4 9 13 0 2
9 15 13 13 3 0 15 15 13 2
7 13 11 3 13 0 9 2
12 13 11 13 9 13 9 12 12 9 1 9 2
6 9 13 3 1 0 2
2 3 3
5 2 13 15 13 2
10 9 13 3 0 9 13 13 9 9 2
6 13 11 9 0 9 2
11 9 16 13 3 2 3 13 7 13 9 2
10 9 9 13 7 15 13 13 9 9 2
16 3 3 2 3 12 9 9 1 2 13 13 9 9 12 9 2
7 11 9 13 10 9 0 2
3 9 9 2
7 15 15 15 13 13 15 2
16 13 13 3 11 9 9 2 16 13 16 9 15 13 9 13 2
7 11 13 11 1 9 9 2
13 15 13 15 3 10 10 9 1 2 7 13 11 2
15 16 9 13 0 2 0 7 0 2 3 15 13 15 15 2
2 0 9
8 9 9 3 3 13 0 11 9
12 3 15 13 3 13 9 2 7 13 13 15 2
3 9 13 13
4 16 13 15 2
2 13 0
8 15 13 10 9 1 3 16 2
11 10 9 9 13 9 9 2 3 0 9 2
12 9 9 7 9 9 13 13 3 9 7 9 2
11 3 13 9 7 9 13 3 0 9 9 2
10 15 13 15 3 0 2 15 13 9 2
8 13 13 2 9 9 2 13 2
21 15 1 13 12 15 2 15 3 13 16 15 2 0 9 7 9 2 13 13 13 2
10 7 3 13 3 3 10 0 13 15 2
16 12 0 9 2 0 9 7 9 2 13 2 0 0 9 9 2
14 13 13 9 13 9 1 12 9 2 15 13 9 1 2
9 11 9 11 11 13 0 9 9 2
11 11 9 13 9 2 7 9 13 13 3 2
5 13 13 0 0 2
7 3 9 13 13 0 9 2
10 9 13 9 13 9 0 9 13 9 2
36 16 9 13 13 15 2 16 13 13 13 3 0 9 15 13 10 9 2 16 9 13 13 13 2 13 9 2 13 9 2 16 7 16 7 16 2
13 2 13 10 11 9 0 9 2 3 13 9 2 2
9 13 13 13 9 2 13 13 9 2
6 9 13 13 13 3 2
6 15 13 13 3 15 2
12 13 15 13 13 15 0 2 16 13 15 13 2
11 0 1 9 13 0 2 0 1 0 9 2
16 13 13 2 15 3 9 9 13 2 16 3 13 13 0 9 2
4 13 13 13 2
4 15 13 0 11
4 13 7 13 2
3 0 12 9
5 15 13 0 9 2
8 9 13 13 3 12 9 9 2
4 0 9 0 9
5 3 15 13 11 2
6 15 13 9 13 9 2
9 11 13 0 2 15 13 13 13 2
4 13 15 13 2
6 10 11 0 0 9 2
7 13 9 9 13 9 9 2
6 15 13 0 10 9 2
7 13 2 16 15 13 13 2
17 11 3 0 9 11 13 13 7 11 13 13 0 9 3 12 9 2
4 13 15 13 2
16 15 13 15 13 0 9 15 8 16 16 13 13 13 7 13 2
4 2 3 13 2
2 0 9
17 9 9 1 0 3 12 9 9 13 13 3 13 9 10 9 13 2
19 0 9 13 13 9 7 13 9 2 13 3 0 9 3 3 3 16 9 2
5 15 15 13 13 2
6 0 9 13 13 9 2
6 15 13 3 3 9 2
8 9 13 2 16 11 9 13 2
2 13 13
4 6 15 13 9
10 9 13 7 13 10 9 13 9 3 2
9 9 13 3 13 12 9 3 12 2
13 3 13 13 3 2 16 3 13 0 2 13 15 2
3 9 13 9
12 10 9 16 13 15 13 9 2 13 0 9 2
6 9 9 13 9 12 9
4 0 9 13 9
4 9 13 9 9
4 13 13 3 2
6 15 13 13 10 9 2
8 15 13 9 7 9 9 9 2
8 9 13 3 0 9 16 9 2
12 16 13 3 0 2 3 3 13 13 3 13 2
9 9 13 13 9 3 16 9 1 2
4 9 13 13 13
5 0 13 9 9 2
4 13 2 9 2
15 3 13 13 13 0 9 9 2 7 13 10 9 13 0 2
5 9 13 0 9 2
16 9 13 9 10 3 16 13 13 13 3 9 7 0 9 9 2
7 15 3 13 13 9 0 2
2 9 3
5 15 15 3 13 2
3 11 11 9
10 2 6 2 2 13 7 13 13 9 2
14 13 12 9 3 9 13 13 15 16 13 13 9 13 2
10 9 13 3 13 2 3 15 13 9 2
10 0 9 9 13 9 2 7 3 9 2
4 15 13 3 2
3 13 9 2
3 13 3 2
13 3 15 3 13 9 9 7 3 10 9 0 9 2
8 3 11 0 2 0 2 9 2
14 0 11 11 13 9 11 3 2 7 9 9 13 0 2
7 0 9 13 10 9 13 2
6 9 13 2 9 3 2
5 11 13 9 9 2
7 9 13 3 10 9 13 2
8 9 13 9 1 12 12 9 2
5 15 15 13 13 2
2 0 0
8 9 2 15 13 13 1 9 2
5 9 13 13 9 9
7 15 13 7 13 0 9 2
2 11 11
15 11 9 13 9 13 3 0 9 2 16 9 13 9 13 2
9 11 12 9 13 3 12 9 9 2
9 13 10 9 13 0 7 0 3 2
9 11 9 11 9 13 13 3 9 2
9 10 11 7 11 2 13 3 13 2
4 13 15 3 2
2 13 13
7 11 15 13 13 0 3 2
7 3 9 13 3 13 13 2
6 0 2 9 13 9 2
4 13 9 9 2
4 9 13 0 2
4 15 13 0 13
4 15 13 9 9
10 15 1 11 13 3 0 3 0 9 2
6 11 13 13 13 9 2
14 15 13 16 15 13 13 15 15 1 16 15 13 15 2
11 11 13 13 13 9 13 3 11 11 9 2
5 9 11 13 12 9
9 15 13 9 1 0 9 3 15 1
8 3 15 13 16 15 3 13 2
22 0 3 13 9 13 3 9 2 3 13 3 3 9 7 9 2 7 3 9 7 9 2
9 15 13 9 3 9 0 9 1 2
8 10 9 13 3 3 3 15 2
5 15 13 0 9 2
2 3 16
8 7 15 13 10 3 13 9 2
6 15 13 13 9 9 2
8 15 13 9 15 13 15 3 2
7 11 9 13 3 12 9 2
5 11 11 13 0 9
6 13 9 7 13 9 2
8 11 13 9 9 2 9 9 2
8 9 13 3 0 2 0 9 2
9 13 15 0 9 9 7 9 9 2
7 13 3 0 13 12 12 2
2 3 3
9 15 1 9 13 13 3 9 13 2
7 13 9 0 9 9 13 2
5 9 13 9 15 2
5 3 9 13 3 3
2 10 9
4 13 15 13 2
6 15 13 13 0 9 2
5 9 13 9 0 2
5 13 13 13 9 2
6 15 13 13 9 9 2
5 3 3 10 9 13
12 11 9 2 8 2 8 2 8 2 8 7 8
3 3 13 0
8 15 13 3 3 2 13 15 2
5 7 3 9 9 2
7 15 15 13 13 13 13 2
6 9 13 2 15 13 2
13 16 15 13 10 9 13 2 10 9 13 13 13 2
4 2 13 3 2
7 9 13 13 9 13 9 2
21 15 13 3 13 9 13 3 2 13 13 2 15 13 0 9 2 9 13 13 15 2
6 13 9 3 0 9 2
9 9 13 0 2 7 9 9 0 2
9 13 3 9 2 13 15 3 13 2
14 11 13 3 13 3 12 9 7 15 13 13 3 0 2
8 11 13 9 13 9 1 3 2
6 13 3 10 9 0 2
15 9 13 13 9 1 2 16 9 13 9 13 7 13 9 2
5 9 3 9 1 2
7 9 9 13 3 0 9 2
15 3 11 12 9 9 13 10 9 16 15 13 9 12 9 2
7 3 11 13 0 9 9 2
15 3 0 9 3 13 2 16 9 13 10 9 13 15 13 2
12 0 9 13 3 2 16 9 13 13 1 9 2
18 16 13 10 9 2 3 11 11 2 15 3 13 13 9 3 9 13 2
17 2 3 13 9 2 16 11 13 13 2 2 10 9 13 9 9 2
5 13 15 1 9 2
4 13 13 13 15
4 9 13 3 2
6 10 9 15 11 13 2
17 12 9 13 10 9 2 16 13 0 13 9 3 13 13 15 9 2
2 11 2
7 9 7 9 13 3 3 2
13 15 13 10 9 2 3 3 15 13 13 3 15 2
10 3 15 3 13 13 10 9 0 0 2
8 16 13 12 3 13 13 0 2
11 0 9 13 2 16 3 13 13 3 9 2
17 3 12 12 9 12 13 13 13 10 12 9 2 15 13 0 9 2
8 13 3 9 9 7 9 9 2
7 3 9 13 13 15 0 2
11 13 2 16 0 9 9 13 13 9 9 2
4 11 13 9 2
8 13 13 13 2 16 13 9 2
16 15 13 13 9 2 7 10 9 11 0 9 13 13 3 9 2
4 2 6 6 2
3 3 13 9
4 7 9 7 9
12 13 3 15 13 2 16 9 13 0 9 1 2
8 9 15 13 13 3 9 15 3
6 9 13 9 10 9 2
7 13 9 9 13 0 9 2
6 15 13 12 3 3 12
6 13 15 13 3 15 2
5 15 13 9 9 2
14 9 13 11 2 13 13 15 3 2 13 11 9 9 2
7 15 13 0 7 13 0 2
9 15 13 9 7 15 13 13 13 2
14 3 0 9 3 9 7 9 1 7 0 9 13 0 2
5 15 13 15 9 2
11 9 13 3 13 13 12 9 1 9 9 2
12 13 15 13 9 15 2 13 9 9 7 9 2
9 12 9 13 13 7 3 9 13 2
2 6 6
6 10 9 11 13 0 2
6 10 9 15 13 13 2
3 9 13 0
6 9 13 9 13 9 2
13 13 0 9 0 9 13 2 7 3 10 15 13 2
17 10 9 13 11 9 13 3 0 9 2 15 15 13 0 9 11 2
6 9 13 10 9 9 2
8 11 9 13 13 3 16 3 2
7 11 13 3 13 0 9 2
5 3 9 13 3 2
7 10 9 13 3 16 9 2
10 9 13 9 9 13 3 3 12 9 2
15 11 11 13 3 2 16 13 9 13 13 3 10 9 13 2
6 9 13 13 13 0 2
24 16 15 3 13 10 9 3 3 3 15 3 13 1 9 7 13 7 13 16 15 13 10 9 2
23 9 9 13 3 11 0 7 9 2 15 3 13 0 13 9 7 9 13 9 9 7 9 2
7 9 13 9 2 13 9 2
5 13 15 3 3 2
5 0 9 11 9 1
4 9 13 9 2
8 13 3 9 16 15 3 9 13
11 11 13 9 9 7 9 13 0 13 12 2
2 9 9
7 10 15 13 13 0 9 2
6 9 13 9 0 9 2
13 3 9 13 10 9 2 16 9 13 13 13 9 2
4 11 13 15 9
5 0 9 13 0 9
15 11 13 12 9 2 15 13 10 9 9 9 13 3 9 9
7 16 13 13 2 13 9 9
9 9 2 15 10 12 9 13 0 9
18 11 12 9 2 0 3 13 9 7 0 9 2 13 9 9 13 9 2
4 11 13 9 2
5 15 13 9 1 2
22 9 15 13 9 3 3 2 13 9 1 7 13 2 16 13 9 2 13 3 3 3 2
12 16 15 15 3 13 2 3 15 13 3 15 2
8 9 3 13 7 13 13 9 2
4 13 3 3 2
14 3 3 11 13 11 0 9 2 16 9 13 3 3 2
13 15 13 13 15 2 16 9 9 13 9 0 9 2
3 15 13 15
7 9 13 11 1 3 9 2
5 9 13 9 15 2
5 7 13 16 9 2
9 15 13 15 16 15 13 10 9 2
10 9 0 9 2 15 9 13 12 9 2
15 13 3 13 9 11 11 7 10 9 7 9 2 16 11 2
7 11 11 2 13 15 3 9
14 13 3 13 0 2 16 9 13 13 13 9 9 1 2
5 13 9 13 9 9
7 9 13 12 9 12 9 2
9 13 15 3 9 2 9 7 9 2
8 10 9 13 15 1 13 9 2
5 10 15 13 3 2
6 15 15 13 9 3 2
19 11 9 7 11 0 9 9 12 9 1 13 0 9 9 13 13 10 9 2
19 0 9 13 2 7 3 3 13 2 3 15 0 0 9 1 13 0 9 2
6 0 7 0 9 7 9
15 9 13 9 1 15 9 2 13 0 9 13 3 3 9 2
9 9 13 13 0 16 3 3 2 2
6 10 9 13 11 0 2
7 0 13 3 9 13 9 2
9 6 13 15 13 13 3 3 3 2
11 11 2 9 2 13 3 10 9 1 3 2
6 13 15 13 13 9 2
16 16 15 13 13 3 3 3 16 15 13 15 15 3 10 9 2
8 11 13 2 16 9 13 9 2
6 11 13 13 15 9 2
6 9 13 1 10 9 2
14 15 13 13 0 13 9 1 2 3 13 9 2 15 2
4 13 9 1 2
2 13 13
12 3 13 12 9 3 2 16 9 13 13 0 2
3 13 13 13
20 0 3 13 9 15 2 16 3 13 13 3 13 9 2 13 13 3 9 1 2
6 15 3 13 9 9 2
6 9 9 13 0 9 13
8 9 13 10 0 9 7 0 9
11 2 15 13 11 13 3 0 2 15 13 2
6 15 13 3 12 9 9
7 2 6 6 2 3 13 2
10 13 10 9 13 13 2 15 13 13 2
8 9 13 9 7 11 13 9 2
17 11 9 7 15 2 13 11 15 7 13 2 13 13 15 1 0 2
10 7 15 9 13 2 13 15 7 13 2
4 3 15 15 13
4 13 9 13 9
4 0 13 13 2
14 15 3 13 3 3 13 13 15 2 3 10 0 9 2
7 13 11 10 0 9 1 2
7 9 13 3 10 9 9 2
8 11 10 11 9 13 13 9 2
12 7 15 13 13 11 2 15 13 13 3 13 2
8 15 1 13 13 0 0 9 2
14 7 12 15 9 13 2 6 9 15 13 3 13 9 2
12 9 13 3 13 13 9 0 0 9 13 9 2
11 0 15 13 0 9 1 13 0 9 1 2
3 9 13 9
7 11 13 13 15 0 9 2
12 3 13 9 3 7 9 9 13 3 9 1 2
11 15 9 2 15 13 9 9 3 0 13 2
10 13 3 3 11 13 13 2 7 13 2
5 13 15 0 9 2
2 13 15
2 0 9
3 13 3 15
5 7 15 1 9 2
19 9 13 3 3 15 1 16 9 1 2 7 15 13 7 13 3 3 9 2
16 13 15 13 15 2 15 13 2 13 15 2 15 13 13 13 2
7 15 13 3 3 3 3 16
10 0 9 7 0 9 13 13 1 9 2
4 13 15 9 2
9 12 9 10 9 11 13 9 9 2
14 13 15 3 7 13 11 2 15 15 13 10 3 13 2
5 15 13 3 9 2
13 13 13 2 13 13 2 16 13 15 3 13 9 2
8 0 9 13 3 3 16 3 2
9 13 11 2 16 15 13 9 15 2
5 3 15 3 13 2
4 13 13 3 9
10 11 11 13 0 0 9 16 9 9 2
10 13 10 1 3 2 16 13 13 13 2
10 15 13 13 3 2 7 13 3 9 2
13 9 13 9 13 9 3 3 2 9 0 9 13 2
8 11 11 13 13 3 13 9 2
9 9 13 13 1 13 9 3 3 2
4 13 9 13 9
5 9 13 9 11 2
6 13 15 13 13 3 0
9 13 15 3 9 16 15 13 3 2
5 10 12 13 13 9
14 15 13 3 13 3 10 9 10 9 9 9 9 13 2
12 15 13 13 3 13 2 15 13 13 3 13 2
13 11 11 7 11 13 9 9 13 9 9 7 13 2
12 13 9 9 9 2 13 13 10 3 0 9 2
10 10 9 13 3 3 12 12 9 9 2
2 13 13
6 0 3 10 9 13 2
4 9 11 0 9
7 9 1 13 9 9 9 2
11 13 15 13 0 16 0 9 13 10 9 2
6 11 13 3 9 9 2
21 13 9 9 2 15 13 9 10 9 15 7 11 11 2 7 13 3 13 0 0 9
7 9 13 10 15 16 0 2
10 9 9 13 2 7 3 10 9 13 2
7 2 15 13 13 13 9 2
9 9 13 13 3 16 9 13 3 2
6 9 9 0 13 9 2
12 9 13 9 12 9 2 3 16 0 9 13 0
14 15 16 13 9 9 2 3 9 13 9 13 0 13 2
2 9 9
6 15 13 10 0 9 2
8 9 13 3 3 12 12 9 2
4 9 13 9 2
7 9 13 13 13 9 1 2
12 3 13 9 0 9 16 15 11 12 9 13 2
21 13 13 9 9 9 13 9 2 0 9 2 9 7 10 9 1 0 9 13 9 2
6 9 13 9 9 1 2
6 15 13 13 9 13 2
4 9 13 0 2
13 11 11 7 11 11 13 3 0 9 13 0 9 2
8 13 13 13 15 9 7 9 13
3 13 13 13
2 10 9
10 0 9 13 9 11 1 9 11 9 1
12 0 9 3 13 9 9 3 16 13 13 15 2
15 15 13 3 16 13 3 13 2 9 3 7 9 9 1 2
8 0 0 15 13 9 9 9 2
8 13 15 3 15 3 0 13 2
12 15 13 2 16 15 13 11 9 3 12 9 2
7 13 3 15 0 9 6 2
13 15 13 3 9 2 15 9 13 13 3 1 3 2
7 9 13 9 9 1 11 2
3 13 9 2
10 9 11 11 11 13 13 3 3 11 2
6 13 3 3 13 3 2
5 9 9 13 0 9
10 9 13 13 0 2 7 13 9 13 2
18 15 15 3 3 13 9 11 13 13 15 0 13 0 7 3 0 9 2
2 3 13
14 11 13 9 7 13 11 1 3 15 13 13 9 1 2
6 11 13 11 0 9 2
11 3 9 3 7 15 13 7 13 10 9 2
10 3 9 13 9 13 9 9 13 9 2
9 12 9 9 13 12 9 7 9 2
5 9 13 15 9 9
7 9 13 9 9 9 3 2
7 9 13 13 3 0 9 2
9 9 3 13 3 9 11 7 11 2
7 13 3 3 9 13 9 2
4 9 13 3 2
4 9 13 0 9
2 9 0
10 0 9 13 11 0 9 7 9 1 2
7 13 11 13 9 0 9 2
6 6 11 13 9 3 2
6 11 13 0 9 9 2
7 3 9 13 9 13 3 2
6 11 9 13 0 9 2
10 9 7 9 0 9 13 9 0 9 2
18 15 13 9 15 7 9 2 15 15 13 0 7 3 12 9 13 13 2
16 13 13 9 2 3 7 13 9 3 2 16 13 13 9 3 2
4 15 0 9 2
8 0 9 13 0 9 7 9 2
5 3 13 13 9 2
12 9 0 9 13 9 9 3 13 11 1 9 2
20 15 13 15 11 1 2 7 10 0 9 2 15 15 9 13 0 9 9 1 2
3 9 9 1
4 9 7 9 9
10 11 13 12 9 1 0 9 0 9 2
5 13 13 3 3 2
4 13 3 9 2
4 0 11 7 9
6 15 13 3 12 9 2
4 9 13 9 2
2 0 9
5 13 0 9 11 2
4 2 13 7 2
6 3 3 9 13 3 2
7 9 9 13 9 7 0 2
6 10 9 13 9 16 9
11 9 1 9 7 9 13 13 13 9 1 2
3 10 0 9
3 6 10 9
8 9 13 3 3 9 3 3 2
7 15 13 3 9 1 3 2
5 3 15 9 1 2
4 3 3 0 9
4 13 10 9 2
3 13 3 2
15 12 10 9 10 11 11 3 15 13 13 3 13 10 9 2
10 9 13 3 13 9 13 3 9 13 2
11 11 9 0 9 13 10 9 3 3 13 2
12 6 13 13 15 2 13 11 15 3 2 13 2
13 9 13 9 9 13 9 1 3 13 3 9 9 2
47 7 3 15 3 3 0 16 13 15 15 10 9 2 0 9 7 0 9 15 13 16 13 3 2 7 3 15 0 9 15 13 10 9 3 16 15 13 3 0 3 15 3 16 13 3 0 3
3 3 13 2
9 3 9 13 12 9 9 9 3 13
7 13 11 13 10 10 9 2
7 9 13 7 3 3 9 2
6 9 13 0 7 0 2
5 9 13 3 0 2
10 0 15 13 13 9 13 0 9 9 2
4 9 13 3 9
4 15 15 13 2
2 9 2
17 11 13 11 11 2 7 0 9 13 16 9 13 3 13 9 11 2
2 9 9
19 11 13 15 11 2 13 2 7 15 0 0 9 2 15 13 0 0 9 2
5 9 13 9 1 2
4 12 9 13 15
7 3 15 13 12 9 9 2
2 13 3
10 3 15 3 13 2 3 15 13 9 2
7 15 13 3 13 13 9 2
5 13 13 10 9 2
21 11 9 13 13 2 9 13 2 9 13 2 9 13 2 12 9 13 7 0 13 2
14 3 11 9 12 12 9 9 13 3 0 9 7 9 2
10 7 9 13 13 3 9 1 13 9 2
5 3 13 7 3 2
28 13 9 3 15 1 13 9 0 9 2 16 13 9 13 3 3 9 0 7 15 2 16 15 1 11 13 9 2
11 15 13 0 2 0 2 3 2 3 13 9
7 13 3 15 13 3 3 2
5 15 13 13 9 2
6 9 13 10 10 9 2
9 9 9 13 11 11 7 11 11 2
12 11 13 13 13 9 9 2 16 15 13 0 2
5 13 3 15 13 2
11 13 15 15 2 15 9 1 13 0 9 2
13 11 13 3 15 2 16 9 0 9 13 3 3 2
9 10 15 13 13 7 0 9 13 2
6 13 15 11 10 9 2
5 9 13 1 9 2
16 15 13 3 9 13 11 9 12 2 0 15 15 13 13 9 2
11 16 9 13 0 2 3 9 13 15 3 2
3 9 13 13
8 3 13 13 9 13 3 9 2
7 3 9 13 13 12 1 2
5 3 3 9 13 2
7 13 0 13 3 1 0 9
11 6 13 13 13 3 9 16 13 13 3 13
10 12 9 9 13 9 13 0 7 0 2
9 10 10 9 3 15 15 13 3 13
14 3 3 13 9 2 13 10 9 7 13 15 3 3 2
4 15 13 3 2
10 7 13 3 12 12 3 13 11 9 2
17 9 15 13 9 13 2 7 9 11 1 13 13 10 9 13 13 2
10 9 1 9 7 9 13 13 13 9 2
12 2 13 15 3 0 2 16 9 13 3 13 2
3 11 9 9
9 13 13 11 0 2 7 13 15 2
18 12 10 12 0 9 2 0 11 7 0 11 9 11 13 13 9 9 2
6 9 9 11 13 9 2
14 16 3 13 2 16 13 13 2 13 13 9 13 9 2
6 16 13 2 13 9 2
5 2 3 3 15 2
11 3 0 9 11 13 11 2 0 0 9 2
15 15 13 13 3 2 9 13 10 9 2 7 9 13 9 2
18 15 13 9 1 7 13 3 3 2 3 3 2 3 9 7 0 9 2
6 15 13 16 11 13 0
3 6 3 2
4 9 13 0 9
6 15 13 3 9 1 2
8 16 13 10 9 9 9 9 2
6 13 15 9 3 3 2
14 15 1 13 13 10 9 2 16 9 13 10 0 9 2
9 3 3 0 9 13 13 3 0 2
13 9 13 0 7 0 2 3 15 13 13 9 9 2
12 0 9 13 9 13 0 9 7 10 0 9 2
4 13 0 13 0
9 11 0 9 13 3 3 0 13 2
6 9 13 13 7 13 2
6 13 13 13 0 9 2
6 15 13 3 0 9 2
2 0 3
2 9 9
5 9 13 9 1 2
14 10 9 9 13 0 0 9 2 15 3 0 3 13 2
7 9 13 0 13 2 7 2
3 13 15 2
7 9 2 3 3 0 0 6
11 3 9 13 3 3 3 16 9 0 9 2
26 11 11 13 0 9 2 15 1 11 13 3 9 1 2 13 3 12 3 2 13 13 12 8 7 9 2
10 0 9 2 15 3 13 3 0 13 2
2 0 9
5 3 3 0 13 2
10 0 9 3 0 9 13 0 11 1 2
22 0 9 2 0 2 13 11 7 11 11 10 11 2 15 12 9 1 13 9 11 9 2
9 15 13 15 0 9 13 9 9 2
2 9 13
14 9 13 12 9 1 12 2 7 12 13 3 12 12 2
4 15 13 9 2
10 15 13 3 0 2 16 13 3 3 2
5 9 13 13 15 9
9 7 15 13 10 3 15 3 13 2
6 13 9 3 7 3 2
3 13 9 9
10 3 9 13 12 1 10 13 2 0 2
7 11 7 11 13 9 9 2
17 15 13 2 16 15 7 11 13 13 0 11 9 7 11 0 9 2
11 15 13 3 0 9 10 9 9 3 6 2
6 3 10 9 9 13 2
6 9 13 0 0 9 2
6 9 13 3 9 0 9
4 9 13 3 2
9 11 9 13 3 0 9 7 9 2
17 3 15 13 9 1 3 9 3 7 13 12 9 9 7 0 9 2
8 15 13 13 3 3 13 9 2
6 9 13 9 7 9 2
5 15 13 9 13 2
2 9 9
4 3 13 11 9
16 9 13 3 13 2 16 13 3 3 0 9 10 9 0 9 2
19 9 10 9 2 9 7 9 1 13 3 13 3 13 12 7 3 12 9 2
3 9 13 2
4 13 3 3 2
8 9 3 13 7 15 13 9 2
4 15 13 9 1
7 13 13 9 2 3 13 9
10 15 13 16 13 2 3 13 9 9 2
4 15 13 9 2
6 13 3 9 9 15 2
14 13 15 13 15 3 13 2 13 0 9 2 16 9 13
7 9 13 13 0 0 9 2
14 13 3 2 16 15 13 10 10 9 2 7 13 3 2
12 13 10 9 2 16 13 9 2 15 13 9 2
2 9 9
12 16 0 13 9 9 9 2 3 9 13 0 2
2 0 9
7 9 13 3 3 1 9 2
3 0 9 11
5 9 13 3 9 2
2 0 9
7 9 13 13 12 9 1 2
9 11 9 13 13 3 0 9 9 2
25 13 15 13 9 13 2 13 9 13 2 13 0 9 13 0 9 2 3 0 9 15 13 16 13 2
17 15 13 13 0 9 9 3 2 16 13 9 7 13 9 3 9 2
6 9 13 15 3 0 2
33 2 13 0 9 2 13 0 9 2 9 13 13 0 9 7 11 11 13 13 15 3 3 2 16 13 13 3 13 2 2 11 13 2
4 13 13 3 2
5 15 13 13 0 2
11 3 13 9 0 2 13 11 3 11 11 2
2 0 9
11 9 0 9 1 10 9 13 12 9 9 2
6 10 9 13 3 9 2
12 13 13 0 13 0 2 15 15 13 9 13 2
3 15 13 9
3 13 9 2
11 16 12 11 9 13 9 3 2 13 9 2
9 3 9 13 9 7 3 3 9 2
6 9 13 0 12 9 2
9 13 3 13 9 16 13 13 9 2
4 13 3 13 2
7 13 2 16 13 9 13 9
9 10 9 9 13 9 9 9 9 2
6 0 9 13 9 11 2
4 9 13 3 2
7 9 7 9 13 9 1 2
19 16 9 10 9 13 9 2 13 15 13 13 2 2 15 13 0 9 9 2
8 9 13 11 0 9 9 9 2
17 9 11 11 13 9 13 13 12 9 9 2 7 13 15 0 13 2
5 9 13 9 0 9
6 9 13 12 9 9 2
3 13 7 13
4 9 13 1 9
8 9 13 9 0 9 9 9 2
14 9 7 9 15 13 2 11 13 3 13 0 9 9 2
8 3 3 13 13 13 0 9 2
13 13 13 13 9 3 13 9 13 0 7 9 0 2
14 13 2 15 13 15 0 9 2 15 13 13 10 9 2
5 13 3 3 0 2
12 15 13 0 9 16 3 13 13 9 13 9 2
7 9 13 0 7 9 13 2
12 9 13 16 9 7 3 3 12 9 13 0 2
9 9 9 10 9 13 0 16 9 2
6 13 13 9 9 3 2
11 13 3 3 16 9 13 13 9 0 9 2
4 9 13 9 2
3 9 13 9
2 10 9
4 13 3 9 9
3 13 13 0
29 3 9 13 3 0 2 15 13 13 9 12 12 7 13 2 16 13 3 13 2 3 16 13 13 12 9 3 9 2
45 3 15 13 3 0 16 3 11 13 3 3 3 15 13 11 9 15 13 3 0 9 15 13 3 13 3 13 13 15 13 3 13 16 11 3 13 3 13 3 9 7 15 13 10 9
6 11 13 11 9 11 2
4 15 13 15 2
11 9 2 15 13 2 16 15 13 3 13 2
8 11 9 13 13 3 0 9 2
10 15 13 3 2 3 11 9 9 9 2
9 13 9 9 2 15 13 10 9 2
3 2 13 2
19 12 9 13 9 12 9 7 9 3 3 7 12 9 12 9 7 3 3 2
11 0 9 13 13 0 3 15 1 2 16 2
10 9 13 9 7 13 11 9 9 9 2
11 16 13 3 2 13 12 9 1 0 3 2
9 16 9 13 11 2 11 9 13 2
10 15 13 3 9 7 9 9 10 9 2
31 9 13 2 16 3 13 0 9 13 9 2 0 9 2 15 9 13 13 9 7 10 9 1 9 13 13 10 0 9 9 2
3 13 9 13
14 15 15 13 13 2 16 9 13 0 2 0 0 9 2
13 10 9 15 13 3 3 2 16 15 13 10 0 2
2 15 13
5 9 13 3 0 2
13 3 3 13 13 9 0 9 16 13 3 13 9 2
9 16 9 13 2 13 13 3 3 2
7 13 13 2 9 13 13 2
2 13 13
9 9 13 3 13 16 15 13 3 2
3 12 9 13
15 11 9 2 2 11 0 9 2 2 13 3 0 9 9 2
7 13 13 15 15 13 11 2
8 10 9 2 15 1 15 13 3
5 15 13 13 3 2
12 15 13 0 9 2 16 15 13 3 0 9 2
28 7 3 13 3 3 3 16 3 13 3 0 7 0 10 9 3 15 13 10 9 13 10 9 16 3 3 9 2
3 13 9 2
2 9 9
16 11 13 9 9 11 9 1 7 13 3 11 2 11 7 11 2
9 9 13 13 2 3 9 9 13 2
9 9 13 3 16 9 13 3 9 2
6 3 13 13 15 3 2
10 13 13 0 7 3 0 2 13 11 2
12 13 13 2 16 0 9 2 7 15 13 9 2
5 9 13 10 0 9
3 13 11 9
13 9 9 3 13 15 2 16 9 13 13 12 9 2
3 9 13 9
16 10 9 13 3 0 9 13 13 2 16 13 3 13 9 9 2
6 11 13 13 3 9 2
17 12 9 2 15 9 13 15 2 13 16 10 9 13 0 9 9 2
13 3 9 13 0 9 2 16 9 13 13 0 9 2
9 0 13 9 13 9 3 0 9 2
16 3 0 0 9 13 13 3 13 0 9 2 15 13 9 9 2
4 9 13 0 2
6 9 13 0 9 9 2
6 9 13 12 9 9 2
7 9 0 9 9 13 9 2
4 13 15 3 2
3 13 13 9
20 9 13 12 1 0 9 2 7 9 7 9 13 9 3 3 2 3 7 3 2
7 15 15 13 15 16 13 2
12 11 13 2 16 3 13 13 0 13 9 3 2
29 3 11 11 13 9 9 11 11 13 9 13 9 12 2 13 3 13 2 7 16 13 13 13 2 13 9 3 2 2
15 11 11 9 13 13 9 1 3 0 16 0 9 9 3 2
5 9 13 13 0 2
6 9 13 13 13 9 2
7 15 13 3 0 16 13 2
8 6 16 3 15 1 2 13 2
5 15 13 13 15 2
22 6 3 2 3 13 3 13 3 10 9 3 7 9 3 13 3 16 10 0 15 13 2
9 9 2 3 2 9 7 9 0 2
18 10 9 13 13 3 12 0 9 2 15 13 12 9 3 16 0 9 2
11 3 13 13 13 3 2 16 0 9 13 2
8 15 13 13 10 9 13 9 2
6 9 13 9 7 9 2
8 9 8 7 9 13 13 3 2
14 2 3 0 9 15 13 2 15 13 13 7 9 13 2
6 3 13 9 3 9 2
3 11 0 9
9 11 13 13 15 1 3 12 11 2
14 9 13 13 0 9 2 16 15 13 13 3 0 9 2
15 9 13 2 3 11 2 2 7 9 13 3 6 2 6 2
7 9 13 10 9 10 9 2
16 0 9 13 9 3 12 12 13 9 2 15 13 9 3 12 2
10 3 11 13 3 3 9 7 11 9 2
10 13 15 13 2 15 13 7 13 0 2
5 3 13 3 13 2
12 10 10 9 13 9 3 3 0 16 10 0 2
13 9 13 3 9 12 2 16 3 9 13 10 9 2
9 13 3 3 0 9 0 9 1 2
29 3 13 1 9 0 9 7 13 9 2 16 13 2 16 13 13 3 12 9 1 2 13 13 3 9 16 13 9 2
8 13 15 3 15 2 15 13 2
9 9 13 13 15 10 3 16 15 2
12 9 13 0 13 0 9 9 1 3 9 9 2
2 10 9
8 13 13 0 9 3 9 9 2
2 0 9
6 15 13 15 10 9 2
4 15 13 9 1
5 3 15 13 13 2
7 13 15 13 9 10 9 2
17 10 0 0 7 0 9 13 9 13 15 7 9 7 13 0 9 2
2 9 9
11 16 9 13 3 3 2 13 13 9 9 2
8 3 9 13 3 10 9 0 2
4 11 0 9 9
15 0 9 9 13 13 3 2 7 0 9 9 13 3 15 2
5 15 10 9 13 2
5 0 9 0 9 13
7 0 13 9 3 9 1 2
3 13 15 3
2 3 3
5 9 13 1 9 2
17 9 13 3 3 9 3 0 2 3 1 7 1 12 9 9 9 2
2 3 16
6 13 3 7 13 3 2
10 10 9 11 9 9 13 3 12 9 2
10 9 13 0 2 0 7 9 0 0 2
13 3 13 11 12 9 2 10 9 13 3 11 9 2
4 15 13 13 13
4 0 9 13 9
19 0 9 13 0 9 1 9 2 15 9 1 13 13 0 2 11 13 3 2
11 9 13 13 10 9 2 15 13 7 13 13
3 13 3 2
3 11 11 11
8 11 2 9 2 9 2 13 13
16 9 13 3 3 2 16 15 13 7 13 3 2 15 13 9 2
6 9 13 9 9 9 2
2 13 9
3 13 9 9
9 13 15 0 9 15 13 10 9 2
4 9 13 13 9
11 3 3 0 13 13 3 0 0 13 13 2
7 12 9 13 13 3 9 2
18 9 2 0 13 0 13 2 7 13 0 2 15 3 13 10 9 9 2
11 13 12 9 9 2 16 3 13 13 3 2
16 9 13 3 2 3 3 16 9 13 13 2 9 15 1 13 2
5 9 13 9 9 2
6 10 9 13 0 9 2
9 9 1 9 13 3 3 9 9 2
8 9 0 13 3 3 0 1 2
19 15 1 0 9 13 9 9 7 9 13 13 13 7 13 0 9 15 13 2
17 0 9 1 15 13 0 0 9 2 0 2 2 10 9 13 0 2
11 3 9 13 9 3 0 3 3 9 13 2
8 15 13 0 9 2 13 13 2
5 9 13 13 9 2
9 11 0 0 9 2 0 0 9 2
15 3 10 12 9 13 15 2 7 13 3 2 11 9 13 2
14 10 9 13 13 3 2 16 9 13 13 3 0 9 2
14 9 13 13 9 2 16 13 16 13 15 13 9 13 2
16 9 11 11 7 11 11 7 11 11 13 11 9 15 0 9 2
14 11 13 3 11 7 13 0 9 1 3 3 9 9 2
12 11 1 10 9 13 3 0 2 11 13 0 2
3 15 13 3
4 13 9 13 9
2 13 9
8 10 9 13 13 3 13 13 9
5 7 2 3 3 2
7 13 13 9 3 16 13 2
2 3 2
4 13 15 3 3
6 9 13 7 15 13 2
15 9 13 9 3 2 15 13 9 3 3 3 16 9 13 2
4 15 13 9 2
4 9 13 9 9
7 9 9 9 9 13 9 2
5 15 13 9 15 9
24 9 13 13 15 2 15 15 13 13 7 9 9 2 7 13 0 2 9 13 8 7 0 9 2
6 3 13 13 0 9 2
13 13 3 0 9 3 13 2 15 13 13 3 13 2
4 13 13 9 2
16 3 13 9 2 3 12 2 7 3 3 13 12 9 9 3 2
10 13 13 13 9 3 7 16 15 13 2
5 0 9 13 3 2
6 13 15 3 3 9 2
12 9 13 12 12 2 15 1 13 16 3 12 2
8 9 13 1 9 13 0 9 2
14 0 9 13 9 15 2 16 9 13 7 13 10 9 2
12 13 9 3 15 2 15 13 0 9 10 9 2
5 9 13 0 9 2
6 13 15 10 9 3 2
6 15 15 13 13 3 2
3 9 13 15
15 3 11 7 11 13 13 3 9 2 7 11 15 13 12 2
3 10 0 9
7 13 13 15 13 10 9 2
5 3 13 13 3 2
12 15 13 3 0 2 7 13 3 13 3 0 2
3 13 13 2
6 13 15 3 11 9 2
5 2 3 13 11 2
16 9 13 0 9 1 3 3 7 3 0 9 9 9 9 1 2
12 9 13 13 2 9 13 13 3 3 7 9 2
7 0 9 13 9 0 1 2
4 9 12 9 9
8 9 11 13 13 9 9 9 2
12 0 11 9 9 13 9 2 9 13 11 11 2
6 9 13 10 3 9 2
10 11 12 9 13 13 2 12 13 3 2
9 11 11 7 11 11 13 0 9 2
7 0 16 15 13 13 3 2
4 15 13 13 3
15 9 9 9 13 0 2 7 3 13 13 0 13 15 9 2
2 3 2
8 13 2 16 15 13 13 9 2
11 0 15 13 0 2 15 13 13 3 13 2
25 3 2 15 13 10 9 3 13 10 9 13 16 9 2 9 7 9 7 3 13 15 16 9 13 2
4 9 13 3 6
4 1 9 13 9
3 0 16 13
6 9 13 0 9 0 2
11 11 1 13 3 13 2 13 9 7 9 2
8 13 2 16 9 13 13 0 2
5 15 13 0 10 9
6 15 15 3 13 13 2
11 15 13 9 3 3 13 11 11 9 11 2
3 9 9 9
8 11 13 9 3 3 3 10 9
8 3 9 13 13 13 9 3 2
3 9 13 13
11 9 9 13 9 2 16 9 13 13 9 2
8 15 13 13 0 9 11 13 2
11 11 9 13 9 13 9 13 9 7 9 2
7 15 13 13 9 9 1 2
6 9 13 0 9 1 2
7 11 3 13 10 9 9 2
6 9 13 13 13 3 2
12 11 13 0 9 13 9 2 13 9 7 13 2
8 9 13 0 2 12 9 3 2
4 13 9 13 9
5 9 3 3 15 2
4 2 3 15 2
17 15 13 3 10 9 9 7 13 16 3 13 9 7 3 15 13 2
5 0 9 13 9 2
5 9 13 13 9 2
21 15 13 13 3 13 9 7 13 3 10 9 0 9 2 15 15 13 13 0 0 2
10 16 13 0 2 13 13 13 3 3 2
5 13 9 7 13 2
3 0 0 9
7 10 9 9 13 9 9 2
4 13 0 9 2
12 9 9 13 13 9 2 15 13 0 9 9 2
10 9 9 0 0 9 13 0 7 0 2
8 9 13 7 15 13 9 3 2
15 9 13 13 13 3 2 16 0 13 0 2 16 0 13 2
4 11 13 9 9
14 9 13 15 0 9 7 10 3 15 16 0 0 9 2
9 3 2 13 15 10 9 13 3 3
7 9 7 9 13 3 9 2
6 9 1 13 13 3 2
8 9 9 9 13 3 10 9 2
10 13 3 2 16 13 9 9 15 13 2
5 0 13 9 0 2
6 9 2 10 0 9 2
4 13 12 1 2
8 12 9 0 9 13 9 12 2
8 9 13 15 13 13 9 9 2
31 9 12 13 13 9 2 12 9 7 9 2 12 9 7 9 2 12 9 7 9 2 12 8 7 9 7 3 3 12 9 2
4 9 13 15 2
12 11 13 13 11 2 16 15 13 13 0 9 2
16 0 9 9 11 11 13 11 9 12 9 7 9 11 9 11 2
11 16 9 13 3 9 2 9 13 13 9 2
5 3 3 13 9 2
7 2 6 15 15 13 3 2
14 15 16 13 13 9 3 3 13 13 9 2 3 9 2
4 3 3 3 2
8 3 13 3 13 13 9 3 3
9 11 11 13 3 13 9 9 9 2
11 10 9 9 13 9 9 3 10 12 9 2
24 15 13 13 9 13 7 13 15 2 15 10 0 9 13 0 2 3 9 7 9 7 0 15 2
6 0 9 7 0 0 2
2 13 13
8 15 11 13 9 2 13 9 2
16 11 13 11 9 3 2 16 15 13 0 7 13 15 15 13 2
9 9 13 9 2 15 13 3 3 2
11 7 9 7 9 13 9 9 9 0 9 2
9 9 13 3 2 3 10 0 9 2
18 3 10 9 15 13 13 2 16 15 13 3 13 9 7 13 3 9 2
11 13 15 13 9 7 0 2 15 13 9 2
8 13 15 10 0 7 13 9 2
7 3 10 9 3 3 13 2
10 13 2 13 11 13 11 0 9 1 2
20 15 13 13 9 9 9 2 7 15 13 15 3 2 13 9 9 15 7 13 2
7 3 0 9 9 13 13 2
8 9 1 11 13 13 13 9 2
6 13 3 0 7 0 2
5 13 3 13 9 2
10 13 13 15 13 13 13 2 13 13 2
5 16 15 13 15 2
2 3 0
4 3 3 15 2
5 13 0 13 15 2
9 16 13 13 15 2 9 13 3 2
15 9 2 9 7 10 9 13 13 3 9 9 9 7 9 2
9 9 11 7 9 11 11 13 9 2
10 9 7 9 13 12 7 12 12 9 2
4 0 7 0 9
4 13 9 3 2
19 3 13 9 7 13 11 2 16 13 15 13 10 9 10 9 16 0 9 2
2 10 9
4 11 13 3 15
18 7 15 13 3 13 3 15 13 2 3 15 13 3 3 12 12 1 2
5 13 11 13 3 2
9 3 13 2 7 13 11 9 13 2
11 9 9 11 13 3 13 2 7 13 0 2
2 10 9
13 13 15 3 0 2 13 15 3 13 0 9 9 2
14 11 13 9 7 13 9 3 3 2 16 13 10 9 2
10 15 13 10 9 3 3 13 0 3 2
8 11 7 11 9 13 12 9 2
20 15 13 3 15 13 15 13 7 15 13 3 11 7 11 9 3 3 3 13 2
10 16 10 9 13 2 15 13 13 0 2
6 13 9 13 3 3 2
9 9 13 13 13 9 2 13 9 2
8 9 7 9 3 13 9 11 2
11 0 9 13 11 12 7 0 11 12 9 2
4 9 15 13 0
4 13 13 9 2
9 10 9 15 13 0 0 16 15 13
8 13 3 15 2 16 13 9 2
5 10 9 13 13 2
7 15 13 15 3 3 3 2
19 6 13 7 13 2 9 3 13 3 0 9 7 13 2 16 9 13 9 2
3 15 13 0
21 11 9 1 11 13 11 9 1 13 3 13 10 0 9 2 15 13 13 13 13 2
7 13 11 13 3 12 9 2
3 12 9 13
11 16 0 9 9 13 2 9 13 15 0 2
10 9 15 3 13 2 7 13 0 9 2
10 10 9 9 3 15 13 15 3 9 2
3 9 13 0
10 13 9 0 9 2 15 13 3 3 2
8 11 13 9 7 11 13 9 2
8 3 15 3 9 9 15 13 2
7 9 1 13 13 10 9 2
12 10 9 11 11 13 11 13 13 9 9 3 2
5 3 15 15 13 2
20 15 13 13 9 2 16 16 9 13 9 3 9 3 2 9 13 3 9 3 2
10 0 11 13 3 10 9 13 13 0 2
3 12 9 9
8 9 9 1 13 9 9 9 2
6 16 13 15 15 13 2
2 9 13
6 15 13 15 7 3 2
9 9 13 13 9 3 12 9 9 2
14 11 13 0 9 3 13 10 11 2 15 9 13 0 2
12 10 9 7 15 9 9 9 13 3 13 9 2
5 13 9 3 3 2
12 0 9 9 9 13 9 13 13 3 0 9 2
4 8 7 0 9
7 10 9 13 13 13 9 2
9 9 13 11 12 9 0 12 9 2
2 0 9
9 15 15 13 13 3 0 3 0 2
10 15 13 9 3 0 9 1 7 13 2
4 9 13 9 2
4 13 12 1 2
7 13 13 9 3 0 9 2
8 3 3 13 11 13 9 3 2
7 0 9 13 9 9 0 9
6 9 13 2 9 13 2
5 12 13 13 9 2
7 3 3 13 9 9 13 2
11 9 13 13 3 13 3 2 13 9 9 2
9 2 3 3 3 9 9 15 13 2
5 15 13 15 1 2
9 13 15 13 10 9 16 9 13 2
5 13 9 13 9 2
6 9 9 13 10 9 2
6 3 13 9 13 15 2
2 13 13
7 11 13 3 3 13 9 2
4 11 13 13 2
11 13 3 13 3 13 2 13 9 9 11 2
3 13 13 0
4 9 13 0 2
4 13 3 3 2
13 13 13 3 3 1 12 2 13 13 3 1 12 2
9 11 11 0 9 13 3 13 9 2
15 9 9 13 3 9 2 15 13 11 9 11 11 9 9 2
7 15 15 13 0 9 13 2
9 9 9 13 13 3 9 7 9 2
13 3 10 0 9 13 13 13 3 16 13 9 13 2
7 11 13 9 3 0 3 2
14 9 13 2 16 3 13 13 0 9 13 9 0 9 2
6 9 13 0 9 1 2
7 9 13 9 12 12 0 2
12 10 9 13 10 1 9 10 9 2 11 9 2
12 15 13 0 0 9 3 13 0 2 0 9 2
9 9 9 9 13 3 3 12 9 2
8 13 13 13 10 9 2 9 2
12 11 13 11 2 16 3 13 13 9 1 9 2
14 11 13 9 13 3 9 2 7 16 15 13 1 11 2
5 13 9 13 15 2
10 0 9 9 13 13 13 3 10 15 2
2 12 9
2 13 13
7 3 15 13 15 3 3 2
15 13 3 3 13 15 3 3 3 7 13 15 3 3 9 2
9 11 13 9 10 9 2 7 3 11
12 0 0 2 13 9 11 11 7 9 11 11 2
3 13 0 2
6 9 12 9 3 9 2
3 2 13 2
4 9 13 3 9
5 9 13 9 9 2
9 9 13 13 2 15 9 9 13 2
13 15 13 3 0 9 1 2 16 15 13 9 9 2
2 13 13
6 9 13 9 13 9 2
12 9 2 15 13 0 2 3 13 2 13 15 2
7 3 13 0 7 0 9 2
14 9 13 2 16 13 11 13 13 0 9 9 7 9 2
16 0 9 13 13 13 7 13 2 13 9 7 13 9 0 9 2
4 13 3 15 2
5 15 9 13 0 2
3 9 13 3
8 9 13 13 3 3 0 3 2
8 11 2 12 2 13 9 9 2
7 9 13 11 9 7 11 2
6 9 13 3 13 9 2
9 9 9 7 0 9 13 3 9 2
4 15 13 3 2
5 15 13 11 9 2
9 11 13 13 3 3 3 16 13 2
18 16 9 13 13 2 9 13 9 13 0 9 2 16 13 13 9 9 2
5 11 13 9 9 2
13 12 12 9 11 13 0 9 3 3 2 12 2 2
7 9 13 13 3 16 3 13
4 15 13 0 13
8 11 9 13 3 3 12 9 2
7 9 9 1 13 3 13 2
6 7 3 9 3 13 2
4 6 13 13 3
5 9 13 0 11 2
13 9 13 9 3 13 2 3 16 13 13 0 9 2
6 11 13 3 13 9 2
8 9 13 13 16 13 3 3 2
9 13 9 13 3 2 9 7 9 2
5 13 3 9 9 2
7 9 9 13 13 3 13 2
4 0 9 1 13
2 13 13
11 9 13 13 12 10 9 0 9 2 2 2
8 13 9 2 9 9 7 9 2
5 3 3 13 9 2
4 15 13 15 2
28 3 13 15 16 16 9 3 16 9 3 13 13 7 13 3 3 13 3 16 15 10 9 13 0 7 13 9 2
8 13 13 2 16 9 13 3 2
4 13 13 9 2
5 9 13 12 9 2
7 9 13 3 3 3 13 2
14 13 3 10 10 9 3 3 13 16 3 13 9 13 2
4 3 9 9 2
10 11 11 13 3 9 11 2 9 2 2
11 16 13 13 3 13 10 9 13 9 1 2
4 13 0 9 2
7 13 15 9 2 11 13 2
8 9 13 3 13 9 0 9 2
6 15 13 13 0 9 2
4 15 13 9 1
2 0 9
5 15 13 9 13 2
9 2 3 13 0 9 16 9 2 2
14 13 15 3 0 10 9 7 13 13 0 9 13 15 2
7 6 13 15 13 13 3 2
17 3 13 13 11 13 3 15 2 7 3 16 15 15 13 2 13 2
26 13 9 13 13 9 2 15 13 12 2 3 13 2 16 15 13 0 13 16 9 13 9 1 16 9 2
14 3 9 13 13 3 15 2 16 15 13 0 0 9 2
7 15 13 3 3 0 9 2
6 13 9 7 0 9 2
3 13 3 2
7 15 16 13 9 9 0 2
10 9 13 0 9 2 13 13 7 13 2
7 2 8 13 15 13 13 2
5 15 13 13 9 2
8 15 1 9 9 0 13 9 2
9 3 15 13 2 16 15 13 13 2
8 9 1 13 11 13 9 11 2
9 11 13 13 13 9 15 3 11 2
5 9 13 9 9 3
4 6 3 0 9
13 11 11 9 9 13 12 9 1 2 7 13 3 2
17 9 7 3 9 13 0 9 13 9 9 7 13 15 0 9 9 2
4 3 15 13 2
16 9 13 3 15 2 13 13 0 9 2 15 13 13 13 9 2
10 3 9 0 9 9 9 13 13 15 2
18 10 16 0 9 9 13 9 13 13 13 13 10 3 9 7 9 1 2
38 9 3 13 3 3 15 3 13 7 7 10 0 9 15 13 9 6 9 9 9 15 16 0 9 13 7 7 3 15 9 6 0 9 15 13 15 6 13
11 11 13 13 9 3 3 2 16 13 13 2
4 6 3 0 2
7 9 9 11 13 9 1 2
10 15 13 0 9 2 15 13 15 13 2
2 0 9
2 13 3
17 11 13 9 2 9 2 15 13 3 0 7 15 13 3 0 9 2
3 12 9 9
18 7 16 15 13 3 2 15 13 0 0 9 2 0 9 13 3 9 2
6 9 13 13 9 9 2
8 0 9 13 13 0 9 13 2
10 15 13 3 13 10 9 15 13 10 9
12 10 9 13 15 13 3 9 3 9 13 9 2
7 2 7 13 2 11 13 2
9 0 9 9 13 3 13 0 9 2
3 9 13 9
13 15 2 13 9 13 2 13 13 3 9 7 9 2
11 3 16 9 11 13 3 3 13 2 3 2
14 9 0 9 13 9 2 7 9 15 13 13 9 9 2
6 13 15 9 9 11 2
9 11 13 13 13 3 9 11 9 2
6 9 13 11 0 9 2
2 3 0
2 11 2
3 13 13 15
14 9 13 13 9 13 7 16 9 13 13 9 13 9 2
4 13 9 3 2
5 15 13 9 3 9
7 12 9 13 3 3 0 2
6 15 15 13 3 9 2
8 15 13 9 9 15 13 9 2
4 9 13 11 2
19 9 9 13 7 3 3 2 7 13 15 3 2 13 9 2 13 3 3 2
11 16 15 13 2 15 13 9 13 9 9 2
8 13 3 9 0 9 7 9 2
9 7 13 15 10 11 9 9 9 2
13 16 13 9 2 9 7 0 9 2 13 3 9 2
8 9 13 3 9 1 13 9 2
11 3 9 13 13 12 0 16 9 13 15 2
2 9 0
2 0 9
6 9 1 13 0 9 2
19 15 13 9 1 3 15 13 9 3 7 9 9 9 3 15 13 3 3 2
5 9 9 13 3 0
6 9 13 3 3 3 2
8 15 13 13 15 2 13 15 2
8 9 13 13 9 9 13 13 2
3 15 13 2
35 7 15 13 3 0 9 3 3 13 3 16 3 15 15 13 3 3 3 3 3 15 16 16 15 13 0 3 0 9 3 13 13 9 3 2
2 9 9
10 9 13 13 13 13 9 3 12 9 2
2 9 13
34 3 16 13 16 16 13 10 0 9 15 13 3 3 10 9 3 13 10 9 3 10 9 3 10 0 9 15 15 13 3 3 16 15 13
6 15 13 13 3 13 0
14 13 9 15 2 16 9 7 9 13 0 7 10 9 2
3 9 13 2
3 13 13 3
3 0 16 9
3 11 10 9
12 9 13 9 9 13 13 0 9 9 0 9 2
10 7 9 13 0 12 9 11 0 12 2
16 9 13 3 2 7 3 9 2 11 13 3 3 12 9 9 2
10 11 13 15 1 13 10 9 0 9 2
11 3 9 13 13 3 3 9 16 3 9 2
4 15 13 13 15
19 13 10 12 9 9 9 12 3 7 13 2 15 9 13 13 9 15 1 2
8 13 13 13 9 9 13 11 2
3 13 3 2
6 9 13 15 3 9 2
15 3 3 9 9 13 3 0 9 16 15 2 15 11 13 3
4 9 13 9 2
2 9 15
4 13 0 9 2
6 0 9 11 0 9 9
10 15 13 13 13 13 9 10 9 1 2
6 9 13 2 9 13 2
2 0 9
9 15 15 3 13 2 16 11 0 2
7 13 9 15 15 13 13 2
9 9 9 13 9 9 13 9 9 2
6 15 13 13 13 9 2
4 3 0 9 2
13 9 9 13 13 3 3 2 16 9 13 3 3 2
7 15 13 13 11 1 9 2
7 11 13 13 9 9 1 2
7 9 13 9 13 13 3 2
8 9 9 13 13 9 0 9 2
7 10 0 9 7 12 0 9
5 9 13 13 3 9
10 9 9 13 9 13 9 7 3 13 2
9 3 13 9 9 0 9 3 0 2
6 9 13 13 13 9 2
10 9 9 9 13 13 9 3 3 3 2
8 13 13 0 9 7 0 9 2
4 12 9 0 9
7 9 1 15 13 13 15 2
12 16 13 9 1 9 2 3 13 3 11 1 9
17 10 9 13 0 2 15 1 15 13 0 9 0 13 7 0 13 2
11 9 13 11 2 15 13 13 11 13 3 2
4 13 15 3 2
12 15 2 16 9 13 0 9 2 13 0 9 2
4 3 13 9 2
10 9 13 9 2 16 15 13 13 9 2
8 3 13 3 15 3 0 0 2
11 13 3 0 9 2 16 13 13 13 3 2
11 13 3 9 2 9 7 9 13 0 9 2
10 10 9 9 3 3 13 11 3 13 2
2 13 13
15 10 9 13 13 3 3 13 9 2 7 3 13 13 13 2
5 3 9 13 0 2
7 15 13 9 13 0 9 2
4 9 13 13 0
2 9 11
6 15 3 9 13 0 2
5 12 13 0 9 2
2 0 9
8 9 13 11 3 13 11 9 2
8 15 13 13 3 3 9 9 2
5 9 13 13 0 2
12 3 15 9 13 15 13 16 15 13 13 1 2
7 3 0 9 9 13 9 2
9 9 13 3 11 13 3 16 3 2
6 9 1 13 9 9 2
7 15 13 0 16 15 13 2
11 6 16 10 9 13 13 2 13 15 13 2
12 9 13 3 13 0 2 7 15 3 0 13 2
5 10 9 15 13 2
7 9 13 13 2 3 9 2
2 10 9
14 9 2 0 7 9 9 13 9 3 2 9 3 3 2
8 11 13 9 7 11 13 9 2
4 13 15 13 2
6 9 9 13 3 15 2
4 9 13 0 9
14 16 11 9 13 13 2 13 16 3 3 15 13 13 2
19 9 13 9 9 13 3 13 8 2 13 13 9 13 13 9 2 8 8 2
2 13 15
10 10 13 7 3 13 9 13 13 3 2
8 10 0 7 3 0 9 13 9
10 9 13 10 9 7 9 7 0 9 2
8 3 15 13 7 13 3 3 2
9 13 15 9 2 7 13 13 3 2
3 0 9 9
13 9 9 13 10 9 10 13 9 7 13 9 9 2
10 9 13 9 13 13 9 8 7 9 2
7 13 15 3 15 3 13 2
7 11 13 0 9 13 9 2
6 9 13 13 13 0 2
22 3 15 13 3 13 16 11 13 3 9 13 3 15 1 15 13 9 9 7 0 9 2
3 13 9 9
9 3 10 9 13 3 9 0 9 2
4 13 3 0 2
5 3 3 15 15 2
3 13 3 13
7 11 11 13 9 0 9 2
3 13 9 2
14 13 15 3 0 9 16 3 2 13 3 13 0 9 2
9 13 9 13 0 9 13 15 9 2
4 13 13 3 9
4 15 13 12 9
12 13 13 12 9 2 3 16 11 13 9 3 2
3 13 9 9
12 11 13 9 9 7 13 9 13 0 11 9 2
12 9 9 13 12 9 2 15 15 13 13 9 2
2 10 9
3 6 9 2
7 10 9 13 3 7 3 0
9 9 13 3 9 7 9 13 9 2
23 11 13 12 10 10 9 0 7 12 9 0 0 9 2 15 1 0 9 0 0 9 13 2
9 9 9 13 9 7 9 9 9 2
17 13 2 16 15 13 0 7 3 0 9 13 9 13 2 13 11 2
2 0 9
4 3 12 9 9
8 0 13 9 0 2 3 15 2
6 9 13 9 0 9 2
8 15 13 9 11 0 9 9 2
2 0 9
6 11 13 3 9 3 2
10 10 9 13 15 9 9 7 11 9 2
10 9 9 13 7 9 1 13 0 9 2
6 13 9 3 9 13 2
5 9 9 13 9 11
10 11 13 0 9 3 9 0 9 9 2
4 9 13 9 2
3 15 13 2
8 11 13 3 16 13 15 9 2
6 0 16 3 13 13 2
5 15 13 15 1 2
13 7 11 13 16 15 13 13 3 9 2 13 9 2
3 13 9 2
6 9 13 9 16 15 2
9 15 15 13 13 13 3 3 9 2
9 10 9 13 15 13 3 10 9 2
8 7 3 15 13 9 1 3 2
15 13 3 0 9 2 7 13 2 16 11 9 13 12 9 2
11 15 3 13 3 11 3 13 3 9 7 2
23 13 13 0 15 9 7 9 9 9 13 11 13 13 9 13 10 9 2 15 13 13 13 2
3 9 13 13
14 15 3 13 9 2 15 3 3 13 13 3 10 9 2
6 13 11 13 3 9 2
3 9 13 2
20 15 2 3 9 13 7 9 13 2 9 13 3 0 2 9 2 2 9 9 2
4 3 13 3 2
15 13 3 0 9 16 9 13 3 0 7 3 16 15 13 2
11 13 9 13 12 9 7 0 9 9 13 2
3 10 0 2
3 15 13 9
4 11 7 11 13
17 9 13 2 7 0 9 2 15 13 11 2 11 11 2 13 0 2
10 13 15 13 13 2 13 9 13 0 2
5 9 13 3 2 2
7 15 13 9 0 9 9 2
5 11 9 13 12 2
17 10 9 13 9 9 13 3 13 2 16 13 15 10 0 9 13 2
18 0 13 9 13 9 3 8 7 9 2 9 7 9 9 12 9 9 2
2 13 13
23 1 9 13 10 9 2 15 10 9 13 2 0 9 0 13 13 9 7 3 9 13 9 2
3 6 12 9
12 10 15 13 9 3 13 13 9 0 0 9 2
10 13 9 13 0 13 10 9 0 9 2
5 13 12 9 9 2
7 10 9 9 13 13 9 2
7 12 9 11 13 15 9 2
22 10 9 2 15 10 9 13 3 0 9 9 2 13 15 3 3 2 3 13 0 9 2
7 11 7 11 13 9 12 9
4 13 11 1 2
10 9 1 11 9 13 3 0 7 0 2
2 13 11
8 10 9 15 3 13 1 9 2
14 7 3 15 3 13 9 7 9 2 7 13 9 3 2
10 10 9 13 3 9 10 9 2 11 9
12 13 9 13 3 0 9 3 9 1 2 9 2
6 9 1 9 13 0 2
5 15 13 11 1 2
3 13 13 2
6 15 13 0 9 3 2
9 9 9 13 3 3 0 9 1 2
3 1 9 9
12 7 13 15 10 0 9 13 2 15 13 9 2
10 11 9 9 13 10 0 9 16 13 2
17 9 13 13 3 0 2 15 7 11 7 9 9 13 0 9 13 2
13 0 9 13 3 9 0 9 2 7 13 3 15 2
7 11 13 13 9 9 9 2
4 9 1 13 9
3 13 9 9
13 9 13 13 13 9 2 15 13 9 9 7 9 2
7 11 15 3 3 13 9 2
4 15 13 13 2
7 15 1 13 15 9 11 2
5 15 13 15 9 2
7 9 11 13 11 0 9 2
12 13 13 0 9 16 13 13 13 9 0 9 2
10 11 9 13 11 12 9 1 0 9 2
3 15 9 2
15 11 7 11 13 9 0 9 2 15 13 13 0 9 9 2
10 0 9 15 13 2 15 13 9 13 2
3 13 9 2
8 8 7 9 13 3 0 9 2
3 13 1 9
14 13 15 3 2 16 9 9 9 7 13 15 2 13 2
3 9 13 9
16 11 13 2 16 15 13 3 9 9 2 16 11 13 13 9 2
10 13 3 3 2 16 13 13 13 9 2
10 2 15 13 15 9 2 13 3 9 2
7 9 13 10 9 12 9 2
13 9 0 7 0 2 0 7 0 9 13 3 3 2
5 15 13 0 9 2
5 9 13 9 9 2
6 11 9 13 3 0 9
10 9 9 13 13 13 0 7 0 3 2
7 11 11 13 11 11 1 2
15 13 13 9 2 15 13 2 16 10 9 9 9 13 0 2
2 13 2
4 3 9 1 13
2 3 3
2 0 9
16 9 13 13 9 9 2 7 13 2 16 9 13 13 10 9 2
43 7 15 13 3 16 15 13 13 13 9 15 3 16 16 3 12 10 12 13 0 9 15 1 0 3 15 15 15 13 16 15 3 13 3 0 3 16 15 13 13 9 9 2
18 9 13 13 3 0 2 16 9 13 13 7 13 9 9 13 9 1 2
10 9 9 9 3 13 12 9 12 9 2
13 3 9 13 13 0 13 3 0 9 1 0 9 2
3 9 0 9
15 3 0 9 9 13 13 13 10 10 9 2 15 13 9 2
2 6 2
4 2 13 13 2
6 13 15 13 16 13 2
5 6 3 13 11 6
3 13 13 2
8 16 13 10 9 9 9 9 2
9 9 7 9 13 0 9 9 9 2
9 13 13 0 13 10 10 0 9 2
5 11 13 0 9 2
12 11 13 13 9 2 7 3 9 13 13 13 2
5 13 15 13 9 2
14 16 13 10 9 3 13 3 6 15 13 13 3 15 2
5 11 9 13 9 2
6 3 13 9 1 9 2
8 12 9 1 9 13 3 9 2
11 9 11 11 13 3 9 11 11 0 9 2
5 13 3 10 9 2
16 16 13 16 9 13 13 2 9 13 16 13 3 13 3 9 2
13 16 9 13 12 9 1 2 15 13 11 3 0 2
5 3 13 9 0 9
8 13 13 3 13 10 0 9 2
7 9 13 13 3 3 12 2
3 9 13 11
9 11 13 3 12 9 11 11 9 2
5 9 9 13 0 2
2 11 9
14 15 13 2 16 9 13 2 9 13 3 2 9 13 2
20 7 3 15 13 3 10 9 16 3 13 3 0 13 0 0 13 15 3 9 2
4 9 13 9 2
7 13 15 3 2 10 9 2
2 9 9
5 9 9 13 3 2
10 13 3 2 16 0 9 9 11 13 2
6 2 15 13 9 9 2
9 9 13 3 11 7 0 9 11 2
10 3 9 2 9 13 3 13 3 9 2
14 3 13 9 2 16 0 12 9 9 13 13 11 9 2
5 2 15 13 9 2
13 13 9 2 16 3 13 11 3 13 3 3 9 2
14 9 13 9 2 15 13 3 10 0 9 2 15 13 2
16 9 13 3 15 2 16 9 13 13 13 9 0 9 11 9 2
2 0 9
16 15 13 3 0 9 13 13 2 7 13 3 9 9 2 15 2
13 2 13 13 2 3 10 9 13 15 1 13 2 2
4 13 15 9 2
4 6 3 13 2
4 13 11 1 2
3 13 9 1
4 9 10 0 9
10 11 13 10 10 0 2 9 2 9 2
5 9 13 9 13 2
5 15 13 9 13 2
5 3 9 13 9 2
15 13 9 0 9 2 3 9 2 9 2 9 2 9 3 2
4 15 13 3 3
11 3 11 11 13 9 13 13 15 9 11 2
10 9 11 9 13 9 3 1 10 9 2
27 9 7 10 9 13 13 13 9 2 3 16 13 15 13 7 13 2 9 9 2 9 11 13 9 9 9 2
11 13 3 0 2 16 13 13 3 9 9 2
12 15 13 0 15 2 16 10 9 13 3 13 2
6 13 11 3 10 9 2
8 15 15 3 13 2 15 13 2
12 9 1 11 13 13 3 0 9 7 9 13 2
5 10 9 13 0 2
6 13 3 13 10 9 2
2 9 9
15 10 9 11 13 16 13 15 0 2 0 9 15 9 13 2
2 3 3
12 3 13 9 13 13 0 13 7 9 13 9 2
9 10 9 13 0 9 13 3 13 2
9 7 3 0 12 9 13 15 0 2
6 9 12 15 13 9 2
3 13 3 2
2 13 3
7 15 2 15 13 3 0 9
8 3 0 9 3 2 13 9 2
7 0 13 13 0 9 9 2
9 15 13 10 15 2 0 0 9 2
2 9 9
15 13 2 10 13 2 7 13 2 13 10 9 2 9 1 2
8 3 9 13 3 0 9 1 2
9 10 9 13 13 9 2 3 3 2
5 15 13 3 3 2
3 15 13 9
4 2 10 9 2
2 10 9
7 9 15 13 9 9 13 9
15 9 13 13 13 2 7 9 13 13 13 3 9 9 1 2
10 7 9 2 15 13 3 13 11 9 2
5 9 7 9 13 9
15 3 13 9 2 7 13 0 9 2 15 3 13 0 9 2
7 0 9 7 3 9 13 2
7 11 13 10 9 9 9 2
10 16 15 13 13 2 15 15 3 13 2
10 13 3 3 9 3 2 13 0 9 2
9 9 13 9 3 9 3 10 9 2
4 3 13 13 2
3 13 13 13
4 15 13 3 2
2 9 9
16 13 13 13 15 2 16 13 0 9 13 0 0 9 9 9 2
5 9 13 9 1 2
6 15 13 3 10 9 2
4 15 15 13 2
10 13 13 3 13 10 9 1 7 1 2
8 11 9 11 13 3 9 11 2
12 3 3 13 9 9 2 7 6 15 13 13 2
10 13 13 15 13 2 13 13 15 13 2
6 15 13 3 9 1 3
5 9 9 13 9 2
4 15 15 13 2
3 13 0 2
12 13 0 7 0 2 13 3 3 3 3 13 2
2 13 9
9 9 12 15 13 13 3 12 12 2
21 7 16 0 9 15 15 13 3 16 2 16 15 13 15 3 0 1 13 0 0 13
7 13 15 3 13 0 9 2
4 9 9 13 11
9 13 0 9 9 9 2 13 3 2
10 9 13 2 16 9 9 13 3 9 2
11 15 13 9 2 16 13 13 15 3 3 2
5 13 13 9 11 2
8 3 13 9 9 1 13 9 2
15 9 13 3 11 13 10 9 10 9 1 2 7 13 3 2
2 3 2
7 13 9 7 9 7 15 2
12 9 7 0 9 13 3 3 10 9 7 9 2
9 13 3 13 2 16 13 3 3 2
3 9 13 9
8 3 13 9 13 2 13 9 2
12 0 9 13 13 9 7 9 9 9 12 1 2
8 10 9 11 13 9 12 9 2
6 0 9 13 0 9 2
3 15 13 15
17 3 0 11 13 3 9 3 0 12 3 9 16 0 12 3 9 2
4 9 13 0 2
6 9 9 13 13 9 2
5 9 13 0 0 2
12 3 3 15 3 13 13 13 16 15 15 9 3
15 2 13 15 3 3 13 2 2 11 13 3 13 9 1 2
7 13 15 3 1 9 13 9
3 0 15 13
9 13 13 9 9 2 16 13 13 2
2 0 2
6 11 13 10 9 0 2
19 16 10 9 13 3 0 11 2 13 10 9 13 0 2 16 3 3 13 2
14 10 9 13 13 3 15 2 16 13 9 9 3 13 2
7 10 9 9 13 3 0 2
5 3 15 13 9 2
5 15 3 0 13 2
9 3 13 3 3 9 16 13 13 2
2 0 9
7 15 13 3 9 7 10 0
2 13 13
4 3 12 9 9
5 11 13 3 9 2
3 10 9 9
10 9 9 13 3 12 7 9 9 9 2
6 3 0 13 3 0 2
5 2 10 3 9 2
6 9 13 3 0 9 2
3 0 3 2
3 3 13 11
3 13 11 2
5 11 13 9 3 2
7 3 13 13 2 11 13 2
5 9 2 15 13 9
6 11 13 9 0 9 2
5 12 9 13 0 2
3 2 0 2
6 9 12 9 13 9 2
10 9 0 9 13 3 3 13 9 9 2
7 13 9 13 15 9 3 2
8 0 0 9 13 13 0 0 2
7 12 0 9 13 9 1 2
4 11 13 9 2
20 3 13 3 9 3 9 3 15 13 3 15 13 7 2 15 13 3 9 15 2
13 3 13 2 2 6 13 2 13 15 15 13 2 2
2 0 9
6 13 0 2 0 7 13
13 11 13 3 0 2 16 11 13 13 9 3 3 2
4 3 9 13 0
5 10 9 3 13 2
5 3 13 0 0 2
10 0 13 9 2 15 13 0 16 9 2
8 9 13 0 2 0 7 0 2
4 13 13 9 2
5 9 13 13 9 2
5 9 15 13 13 2
8 3 13 13 13 9 0 9 2
17 9 0 9 9 13 13 11 9 2 16 0 9 13 15 9 11 2
15 11 13 10 9 2 15 13 15 2 16 15 13 13 13 2
15 9 2 0 9 13 3 0 2 0 9 9 0 9 13 2
4 13 15 11 2
5 3 0 9 13 2
11 9 13 13 9 3 11 7 11 1 11 2
7 10 9 9 13 9 13 2
13 3 13 3 2 9 2 13 16 13 2 13 13 2
10 2 15 13 0 9 7 13 3 3 2
17 10 2 10 9 13 0 9 2 9 13 0 16 13 3 0 9 2
3 0 12 9
10 10 13 9 13 0 9 13 3 0 2
7 15 3 10 0 1 0 2
2 13 9
6 15 15 3 3 13 2
5 11 13 9 9 2
13 13 13 2 16 3 13 13 13 3 9 9 9 2
16 13 3 2 16 3 9 9 13 3 0 0 9 13 0 9 2
5 11 13 3 0 2
13 16 15 13 12 9 2 15 13 13 13 13 9 2
11 3 9 13 13 13 2 16 9 13 9 2
9 3 13 0 9 2 9 2 9 2
11 15 13 9 9 0 9 7 15 13 9 2
6 15 13 3 10 9 2
3 13 0 2
7 3 13 9 7 9 11 2
3 15 0 2
13 9 9 13 15 2 16 9 13 13 10 9 1 2
3 12 0 9
4 9 13 9 9
14 13 10 9 13 13 10 9 9 13 2 16 15 13 2
14 0 9 9 13 15 2 16 15 13 9 9 0 9 2
17 2 9 15 13 0 7 0 9 2 16 3 10 9 13 13 9 2
6 0 9 13 9 9 2
5 15 13 3 13 2
4 15 15 13 2
15 16 15 13 13 2 15 13 9 9 9 1 7 13 9 2
9 0 9 3 13 3 9 9 9 2
16 9 13 3 9 2 13 9 9 0 10 9 7 3 9 9 2
10 3 16 15 13 3 3 13 12 12 2
9 10 3 0 9 13 13 9 9 2
5 13 15 13 3 0
6 13 13 0 13 3 2
6 9 13 11 9 9 2
12 7 16 3 13 3 15 3 0 10 9 16 2
16 16 10 9 9 13 0 2 13 15 3 9 13 3 0 9 2
10 10 9 7 10 9 9 13 3 1 2
8 3 9 13 9 3 0 9 2
6 11 13 13 13 9 2
7 9 13 0 12 9 9 2
6 9 13 3 16 3 3
5 9 1 13 13 2
9 9 11 13 9 9 0 9 9 2
6 9 13 13 0 9 2
7 9 13 13 15 0 0 2
10 0 0 9 1 13 7 13 0 9 2
10 13 13 9 2 16 13 3 3 12 2
8 11 3 3 13 0 9 9 2
10 9 13 9 9 11 7 11 9 1 2
8 15 1 0 11 13 13 0 2
15 9 13 13 9 7 9 2 9 3 13 9 2 7 9 2
4 13 0 13 2
2 9 15
9 9 13 0 2 7 13 3 15 2
15 11 13 13 3 0 9 0 9 7 9 13 0 11 9 2
10 0 0 9 1 3 9 13 13 3 2
3 15 13 0
11 9 15 2 15 15 7 11 13 3 13 2
6 13 3 3 3 0 2
17 9 1 13 9 1 13 13 0 9 3 7 16 9 13 3 13 2
6 15 13 3 0 9 2
20 16 9 13 13 3 0 9 2 13 9 3 13 9 7 9 2 15 15 13 2
10 9 15 13 9 9 7 9 13 13 2
15 0 9 12 12 13 0 7 3 0 9 9 10 9 1 2
6 9 13 3 0 9 2
16 16 15 15 3 9 13 3 15 13 3 3 3 12 12 1 2
14 7 15 0 9 13 3 2 16 12 13 9 3 0 2
3 3 3 2
8 11 7 11 1 13 0 9 2
3 13 12 9
7 9 13 0 3 1 9 2
9 13 9 0 9 3 3 13 13 2
14 0 9 13 13 3 9 2 15 13 13 9 7 9 2
4 9 13 10 9
10 11 13 2 16 13 9 3 3 13 2
9 9 13 3 13 0 12 9 9 2
14 0 9 13 13 3 9 7 13 3 13 15 13 9 2
7 2 15 13 13 13 15 2
18 9 13 13 9 2 13 9 7 2 7 7 2 9 3 9 1 7 2
7 11 13 9 1 13 9 9
17 0 13 0 2 15 0 13 13 2 13 3 3 2 7 3 3 2
4 15 13 12 12
8 3 9 7 9 3 1 9 2
4 15 13 9 2
5 13 3 3 0 2
4 9 13 13 3
4 9 0 9 11
16 3 9 13 9 0 9 2 7 12 9 9 9 13 3 9 2
4 13 0 9 9
11 3 9 9 13 9 2 15 9 13 0 2
4 13 9 0 2
5 13 15 3 13 2
5 9 13 9 9 2
4 15 9 13 2
6 11 13 0 9 9 2
12 13 3 10 0 9 2 15 15 13 13 0 2
9 13 9 7 13 0 7 0 9 2
2 10 0
2 10 9
6 3 13 13 10 9 2
10 11 13 0 9 2 15 13 0 13 2
19 7 16 13 13 10 12 2 15 1 15 13 2 13 7 15 7 10 12 2
7 16 15 13 9 13 9 2
5 6 13 13 3 2
8 13 3 15 3 13 10 9 2
22 11 13 13 13 9 1 11 9 2 7 13 15 13 13 16 13 13 3 13 13 3 2
8 0 13 0 9 15 2 15 2
13 3 3 10 9 13 9 2 3 3 9 9 13 2
13 3 15 13 9 7 0 9 1 10 9 15 13 2
6 13 15 13 3 3 2
10 9 13 9 2 13 9 7 13 9 2
17 9 13 13 15 3 15 11 13 9 3 13 7 9 13 9 2 2
10 15 13 2 9 2 13 7 13 9 2
8 15 13 9 9 3 13 15 2
15 3 13 9 2 15 13 11 0 9 13 9 12 9 1 2
18 15 13 10 9 9 1 3 0 9 3 2 16 9 13 7 13 9 2
3 13 13 0
8 9 13 13 15 15 10 15 2
3 13 3 2
4 9 13 9 2
2 3 15
23 15 13 0 9 11 9 11 12 9 7 13 13 15 9 2 15 10 9 13 13 3 13 2
13 7 3 15 13 13 16 13 0 16 15 13 10 9
9 15 13 3 9 2 13 9 3 2
8 13 9 6 2 11 11 13 2
4 9 13 13 2
4 13 9 1 2
6 13 2 16 13 13 9
6 3 0 9 13 13 2
4 9 13 15 2
20 3 15 13 13 3 0 2 16 9 13 0 13 13 13 10 9 13 13 13 2
9 11 9 13 9 3 12 0 9 2
9 13 13 2 16 15 13 9 2 2
6 13 9 10 12 9 2
7 0 9 11 13 9 11 2
6 15 13 3 3 3 2
13 13 9 2 16 9 1 13 9 9 13 13 9 2
6 0 0 9 13 9 2
14 9 3 3 13 3 2 3 13 3 7 13 7 13 2
2 10 9
8 13 13 3 0 16 15 13 2
5 3 15 13 9 2
14 11 2 9 2 13 3 9 2 8 7 9 7 9 2
8 9 13 16 15 13 13 3 2
33 12 9 9 12 3 13 9 2 9 2 9 7 9 1 12 9 2 9 2 12 9 9 2 9 2 9 2 9 7 12 9 9 2
8 9 9 9 13 0 9 9 2
12 0 9 9 9 9 13 13 13 3 0 9 2
11 15 13 3 13 9 2 15 13 0 9 2
10 15 13 15 11 2 13 13 0 13 2
12 3 3 11 3 7 11 9 13 13 9 9 2
6 9 11 13 3 3 2
21 13 13 11 15 9 3 2 13 13 15 9 2 7 15 13 13 3 0 9 11 2
5 9 13 9 0 2
6 2 3 15 15 13 2
5 15 13 10 0 2
12 9 13 13 10 9 3 3 0 9 13 9 2
4 7 15 13 2
14 9 13 11 2 11 2 11 2 11 7 11 1 11 2
7 11 13 13 15 13 9 2
3 9 13 9
17 10 9 13 13 0 9 0 9 3 13 0 13 15 13 16 15 13
4 3 15 13 2
15 16 13 9 2 3 13 13 13 10 9 3 12 9 9 2
5 13 9 11 9 2
7 13 0 9 13 3 9 2
7 13 10 15 3 13 9 2
5 15 13 9 9 2
4 13 15 0 2
15 9 13 13 9 3 9 9 2 15 13 3 16 9 9 2
3 15 13 9
17 11 13 3 0 9 13 9 2 16 13 13 10 9 3 3 13 2
6 11 9 13 9 0 9
9 9 1 11 13 13 9 3 13 2
7 9 9 13 3 0 9 2
4 9 3 13 2
9 3 13 10 9 0 9 13 9 2
2 0 9
2 13 13
2 13 15
9 15 13 0 2 0 11 13 0 2
4 11 13 9 2
12 13 0 13 2 16 13 9 13 10 0 9 2
5 13 13 3 16 13
5 3 13 3 11 2
4 11 13 11 2
8 0 9 13 9 13 9 3 2
3 13 12 1
12 9 1 13 13 11 3 0 9 13 9 9 2
12 0 9 13 9 2 16 9 13 13 9 9 2
8 9 13 0 7 3 0 9 2
11 13 13 9 3 2 7 3 15 13 15 2
7 13 0 9 9 9 1 2
20 16 9 11 9 2 12 9 7 9 9 13 13 9 2 9 13 13 0 0 2
8 7 10 9 13 13 10 0 2
9 2 3 15 13 9 9 13 2 2
6 3 3 13 13 9 2
10 9 9 13 15 2 15 15 13 9 2
8 10 9 9 13 13 2 15 2
15 13 3 15 13 9 13 9 2 7 13 10 9 13 13 2
8 9 13 0 3 9 10 9 2
7 0 9 13 2 9 13 9
4 9 13 9 1
15 9 13 9 13 7 13 9 13 3 11 9 2 13 9 2
4 13 13 3 2
9 13 13 15 2 13 9 7 9 2
3 13 9 1
11 15 13 3 9 13 9 15 2 11 13 2
6 9 13 9 9 1 2
4 9 0 11 11
2 9 9
5 13 3 0 9 2
4 13 12 9 2
11 9 13 0 13 2 7 9 13 13 9 2
15 13 0 13 9 13 10 9 7 13 15 9 10 9 9 2
4 15 13 3 2
5 15 13 9 13 9
11 13 0 9 13 9 3 3 7 9 13 2
3 3 13 2
12 9 13 3 13 13 9 2 9 9 13 9 2
13 15 13 3 0 2 15 13 3 13 2 0 9 2
5 15 13 3 3 2
9 15 13 15 2 15 13 15 9 2
14 10 11 11 9 9 13 0 9 9 1 9 13 9 2
6 9 13 13 11 13 2
29 13 3 15 13 15 13 9 3 10 13 15 3 13 3 12 9 9 16 15 3 13 7 12 7 10 9 8 6 2
4 9 13 3 2
6 13 10 9 3 13 2
15 13 15 13 3 9 3 12 9 2 13 3 10 9 1 9
7 12 9 12 9 13 13 2
4 3 15 13 2
15 11 13 13 11 0 9 7 13 13 13 11 13 3 0 9
8 16 13 11 2 13 3 3 2
12 0 9 13 10 9 2 15 10 9 9 13 2
2 13 13
11 9 9 13 9 2 15 13 10 9 0 2
9 11 13 11 0 2 0 7 0 2
8 9 13 9 0 9 13 9 2
8 13 2 16 13 9 13 9 2
17 13 13 2 16 10 9 13 13 2 7 13 13 2 15 13 13 2
6 15 13 13 0 9 2
2 9 13
15 15 15 13 3 13 15 2 3 9 13 3 13 10 9 2
9 3 13 9 2 13 15 7 9 2
4 13 3 0 9
10 13 6 9 2 11 13 0 9 1 2
2 9 9
4 13 3 0 9
9 7 3 3 15 13 9 3 13 2
22 3 13 7 3 16 15 13 13 9 2 13 13 0 9 7 9 2 15 13 13 9 2
3 10 0 15
5 9 9 15 13 2
16 11 2 3 11 13 12 9 9 3 16 15 13 3 3 13 2
21 16 11 13 3 2 15 13 13 9 13 2 13 10 0 9 9 13 9 9 9 2
9 16 13 15 2 15 13 13 13 2
26 7 16 0 9 15 15 13 3 16 2 16 15 13 15 3 3 0 15 3 0 1 13 0 0 13 2
9 7 13 15 15 0 10 9 13 2
7 9 13 11 11 13 13 9
8 9 13 3 13 13 9 9 2
5 13 15 3 15 13
4 13 13 3 2
4 9 13 9 0
16 15 13 3 3 16 10 11 1 15 2 16 0 13 9 3 2
6 9 9 1 13 9 9
17 9 9 13 13 13 10 9 2 13 3 11 9 13 9 11 11 2
12 9 13 0 7 9 13 0 2 7 13 3 2
10 10 9 0 9 11 9 13 15 2 16
4 13 9 10 9
5 15 3 9 13 2
8 9 9 15 13 12 9 9 2
9 0 9 13 9 11 9 0 9 2
3 13 3 2
3 13 3 3
9 8 8 13 0 9 0 7 0 2
14 13 15 2 16 9 13 9 9 7 9 15 13 13 2
14 15 13 13 3 2 3 3 13 13 0 2 11 13 2
6 11 9 13 9 11 2
17 3 13 3 2 7 13 15 3 3 0 16 13 9 0 9 9 2
3 9 13 9
15 9 9 13 9 0 9 7 13 13 9 16 0 9 3 2
10 2 13 15 9 3 13 16 3 13 2
2 10 3
10 3 10 11 9 9 13 15 0 9 2
7 9 1 13 13 12 9 2
11 9 13 3 2 16 15 13 0 9 13 2
7 11 13 9 7 13 15 2
10 3 2 3 6 3 10 9 9 9 2
8 9 9 13 3 15 13 13 2
11 9 13 13 9 0 7 0 13 0 9 2
7 15 13 9 7 13 9 2
3 9 13 2
10 11 0 9 13 11 9 9 12 9 2
16 11 13 15 10 9 13 9 13 3 16 13 9 13 15 0 9
11 9 1 13 13 3 16 15 3 13 9 2
3 13 9 2
11 11 13 13 16 13 13 3 3 13 9 2
4 13 9 11 2
11 13 2 13 15 13 2 10 9 15 13 2
19 9 13 0 9 15 2 16 7 0 7 0 7 0 9 13 9 13 0 2
4 15 13 13 2
9 0 9 3 13 13 3 9 1 2
4 11 13 9 2
17 3 0 9 2 3 3 9 13 9 2 3 16 3 0 13 9 2
8 15 13 3 13 9 3 3 2
8 3 13 2 3 0 9 13 2
11 15 13 12 9 9 2 15 13 13 15 13
3 15 13 15
3 12 0 9
9 15 13 15 2 16 13 3 13 2
4 10 9 13 2
18 15 13 3 13 11 9 2 16 7 3 3 16 15 13 0 16 9 2
14 13 0 9 7 9 3 2 15 13 3 13 0 9 2
19 15 13 2 16 13 2 3 15 13 15 9 2 0 9 2 9 7 9 2
12 15 13 9 2 13 9 7 13 9 3 0 2
12 16 11 13 0 9 2 10 9 13 13 9 9
2 13 13
7 15 13 13 13 9 0 2
4 15 13 13 2
7 9 13 13 9 9 11 2
11 9 9 13 13 3 0 7 0 16 9 2
7 3 11 13 10 9 3 2
7 13 13 0 12 9 0 2
7 9 1 13 13 13 0 9
5 15 9 13 13 2
6 11 13 3 9 3 2
7 9 13 9 3 16 9 2
3 13 3 3
8 6 6 16 11 13 13 3 2
11 13 0 2 16 13 11 13 13 0 9 2
2 0 9
3 13 9 2
8 3 10 9 13 3 13 9 2
6 11 9 13 9 11 9
19 9 9 13 3 1 9 2 13 12 9 11 1 7 12 11 1 13 11 2
15 10 9 9 9 13 13 2 13 15 0 9 16 9 9 2
10 3 11 13 13 15 12 9 0 9 2
11 9 16 15 13 0 15 16 15 13 2 2
7 15 13 3 9 16 9 2
7 9 9 11 9 11 11 2
13 16 15 13 9 13 13 2 0 9 13 10 9 2
4 13 9 9 2
12 15 13 3 6 13 2 15 15 13 9 13 2
10 3 2 9 13 11 1 3 0 9 2
4 15 13 3 2
13 11 13 13 11 3 3 10 11 7 11 0 9 2
5 9 13 9 11 2
9 3 9 7 0 9 13 13 15 2
9 11 0 9 9 9 13 11 0 2
7 9 13 9 3 13 13 2
2 10 9
6 11 13 3 0 9 2
3 9 13 0
13 0 13 13 3 13 3 7 10 3 15 9 13 2
5 9 13 3 9 13
14 13 15 16 11 13 3 16 15 13 15 10 15 9 2
13 13 3 13 2 16 11 13 0 9 2 7 13 2
8 9 13 3 13 9 9 9 2
12 11 9 9 7 15 11 13 9 13 9 9 2
7 11 9 13 0 9 9 2
8 11 13 13 3 11 0 9 2
7 9 3 15 13 15 13 2
10 9 13 0 10 9 2 15 3 9 2
6 15 13 13 0 9 2
15 11 13 13 2 16 13 13 3 10 0 9 16 9 9 2
13 11 11 7 11 11 13 9 0 9 11 11 9 2
6 13 15 3 3 13 2
11 13 15 11 3 2 16 10 9 9 13 2
19 16 9 13 0 9 9 16 10 8 7 9 2 13 3 13 12 9 2 2
7 2 15 13 3 0 3 2
13 13 13 2 16 3 9 13 10 3 0 0 9 2
10 3 15 15 1 13 13 9 3 9 2
7 11 13 9 9 13 11 2
8 3 3 15 2 13 0 9 2
6 9 16 15 13 0 2
12 16 9 9 13 13 11 0 9 0 9 3 2
27 10 9 11 2 15 13 13 3 9 7 0 9 2 13 9 11 0 2 11 13 0 9 13 9 9 9 2
6 15 13 13 9 9 2
9 13 0 2 16 15 13 3 3 2
2 13 13
4 13 16 13 2
12 0 9 13 11 13 3 0 9 16 0 9 2
3 10 9 16
5 3 13 0 0 2
5 0 15 13 0 2
3 13 9 2
18 15 13 3 13 2 16 15 13 9 3 13 2 16 13 13 13 9 2
11 9 2 9 7 9 13 0 0 9 9 2
5 9 9 9 11 11
4 13 13 9 2
5 15 13 13 3 0
5 15 15 3 13 2
15 3 10 9 13 9 12 9 9 2 9 7 9 0 9 2
13 13 9 3 0 7 0 3 2 9 13 3 9 2
14 15 13 3 13 9 2 15 15 7 15 13 13 13 2
2 3 15
2 0 9
3 13 3 2
5 13 15 9 9 3
2 15 13
14 9 13 13 0 7 3 0 9 2 16 13 15 3 2
8 13 13 9 0 2 15 13 2
14 7 1 9 13 3 13 9 2 3 13 3 10 15 2
6 13 9 13 7 9 2
4 15 13 0 9
11 3 12 9 0 2 0 2 0 7 0 9
5 9 13 0 9 2
5 9 13 0 9 2
4 9 13 13 11
3 9 0 9
4 15 13 9 2
2 9 13
11 3 13 2 16 13 9 15 13 3 13 2
5 13 3 3 11 2
14 0 9 13 9 9 13 13 12 9 3 7 9 3 2
4 13 9 3 2
4 11 15 13 2
19 0 9 7 3 9 13 3 9 3 9 7 10 9 13 3 3 2 16 2
3 9 13 13
6 10 9 9 13 3 9
7 15 13 9 3 9 1 2
6 9 13 9 0 9 2
6 3 9 9 13 0 2
8 9 15 13 9 9 0 9 2
5 11 13 12 9 2
13 13 3 13 9 10 9 3 2 11 13 13 9 2
7 9 2 15 13 13 0 9
5 10 15 13 15 2
5 9 9 13 9 2
4 15 13 3 13
9 9 7 9 13 2 15 13 0 2
2 0 9
10 0 12 9 7 3 13 12 9 9 2
4 13 15 9 2
14 9 9 12 11 9 9 13 3 9 9 9 9 11 2
8 11 9 13 3 7 13 3 2
7 13 16 13 13 13 9 2
11 11 12 0 9 13 11 9 7 11 9 2
14 3 11 13 9 12 12 12 9 2 0 9 3 3 2
7 9 13 16 15 13 13 9
11 16 3 13 0 9 2 13 13 9 9 2
11 15 13 10 0 9 2 13 15 10 0 2
12 9 13 3 3 2 16 13 9 3 13 9 2
2 13 3
5 15 13 9 9 2
5 3 3 15 15 13
5 0 2 0 0 9
13 15 13 3 13 3 15 2 16 13 13 15 13 2
14 13 15 13 13 3 2 16 9 9 13 3 0 3 2
10 7 3 3 3 13 6 10 0 9 2
6 11 13 0 3 11 2
5 3 15 13 9 2
5 15 15 11 13 2
12 9 13 3 12 9 0 7 3 12 9 0 2
4 11 13 13 0
5 13 10 0 9 2
15 16 15 13 13 9 2 15 13 9 7 13 12 9 13 2
7 3 9 13 13 3 0 9
4 3 9 13 2
7 9 9 2 12 9 12 9
13 9 13 13 9 9 2 9 9 2 9 0 9 2
7 3 13 12 10 9 9 2
8 10 9 9 13 13 0 9 2
7 9 2 9 7 3 10 9
4 13 9 9 3
12 9 2 11 9 12 2 13 13 9 0 9 2
39 15 13 11 9 2 7 13 16 15 13 1 9 7 15 13 10 9 7 15 13 9 7 3 15 2 13 9 1 3 10 9 2 7 13 9 16 13 10 9
6 3 13 9 0 9 2
2 13 13
21 9 13 13 13 3 9 3 2 15 13 13 0 9 3 7 13 10 9 0 9 2
9 3 13 9 3 3 9 9 1 2
4 9 13 3 9
5 9 13 13 13 2
4 9 13 13 2
11 11 13 3 10 9 9 3 0 9 13 2
10 9 9 13 9 9 9 13 16 3 2
10 9 3 0 9 9 13 9 1 13 2
18 13 2 16 16 13 13 3 13 9 2 13 0 2 16 13 13 3 2
17 10 9 13 9 9 2 15 15 13 13 9 1 3 0 2 9 2
4 13 9 13 9
5 9 13 0 9 2
15 8 7 9 12 9 13 15 2 16 9 13 3 9 12 2
4 15 13 0 2
9 16 11 13 2 13 11 13 3 2
7 9 13 0 7 3 0 2
6 15 13 9 13 3 2
7 9 13 13 10 9 9 2
13 9 13 3 10 9 2 16 3 13 13 9 9 2
4 9 9 9 11
13 13 0 9 2 3 13 0 2 16 9 13 9 2
13 13 15 3 13 13 2 3 13 9 13 13 13 2
10 13 0 2 0 0 2 9 7 9 9
10 13 11 13 2 16 9 13 0 9 2
13 3 13 0 9 2 15 3 0 0 9 13 13 2
4 15 13 9 1
5 3 13 10 15 2
9 9 10 9 1 13 3 0 0 2
12 15 13 0 9 7 0 9 2 7 3 9 2
23 3 15 7 11 13 13 9 2 11 13 13 9 9 2 15 13 3 0 16 15 3 13 2
13 13 9 13 9 9 9 2 7 16 2 3 3 2
12 13 13 3 3 3 15 1 2 16 13 9 2
6 15 13 3 9 9 2
14 15 13 3 0 2 3 15 13 13 13 3 3 9 2
4 9 13 9 1
5 11 9 13 11 2
10 7 10 9 13 3 13 13 0 9 2
15 9 11 13 13 10 9 2 0 13 15 1 9 13 9 2
10 13 13 3 3 16 13 13 9 13 2
2 9 9
6 9 13 0 12 9 2
13 0 9 9 9 13 3 9 9 11 11 9 1 2
4 12 9 3 2
8 15 13 3 3 3 3 3 16
13 9 13 3 10 10 12 9 13 3 3 15 15 2
2 3 3
6 0 9 13 3 9 2
9 11 9 13 12 9 3 12 9 2
4 3 13 9 2
5 0 9 13 3 2
6 3 0 9 13 9 2
7 9 9 9 13 3 9 2
7 9 13 9 12 9 1 2
4 15 13 11 9
16 15 13 13 3 3 2 16 11 13 0 13 13 9 9 9 2
9 9 13 13 2 16 13 9 13 2
12 6 6 2 3 13 12 0 3 0 9 11 2
8 9 13 3 3 13 11 9 2
2 0 11
4 9 13 9 2
8 13 3 10 9 13 7 13 2
6 13 3 3 0 13 2
2 9 0
3 13 9 9
5 9 13 0 9 2
9 9 13 10 9 10 9 3 12 2
5 13 9 2 3 2
9 9 13 9 9 13 15 3 9 2
7 10 0 3 13 15 13 2
5 13 3 3 13 2
12 9 13 13 10 0 2 7 15 15 13 13 2
9 9 13 9 13 15 15 3 13 2
16 11 13 13 11 0 9 7 13 13 13 11 13 3 0 9 2
6 9 13 13 0 9 2
9 15 3 13 10 9 3 15 13 13
8 9 2 15 13 3 9 13 2
2 13 3
5 15 13 9 9 2
17 9 9 13 10 0 9 2 15 0 9 9 13 13 9 10 9 2
2 9 13
3 0 9 2
3 9 9 13
16 9 2 15 13 13 13 3 11 7 10 0 9 13 0 9 2
4 0 15 13 2
2 9 9
5 9 13 0 0 2
5 9 13 9 13 2
4 15 13 9 1
6 3 13 13 10 0 2
9 15 2 16 9 13 2 13 0 2
7 15 13 0 9 13 3 9
4 15 13 15 2
18 2 7 9 13 13 0 2 16 3 3 13 13 2 2 15 13 9 2
24 16 7 9 9 7 15 9 13 0 9 2 13 15 13 13 0 9 2 15 13 9 13 9 2
6 15 13 3 12 9 2
4 8 7 0 9
12 11 13 13 9 9 7 16 9 13 0 9 2
12 13 9 3 3 10 9 7 13 9 0 9 2
7 15 13 13 3 0 15 2
20 1 10 9 13 2 8 11 11 2 9 11 0 9 16 13 3 13 9 9 2
15 11 13 9 13 2 16 9 9 9 13 0 3 12 9 2
3 13 15 13
6 9 13 3 3 13 2
10 9 1 10 9 13 13 13 10 9 2
15 13 13 3 3 13 2 16 13 13 9 0 9 9 1 2
7 13 15 3 3 10 9 2
5 9 15 13 0 2
6 9 11 9 13 12 2
7 13 15 15 13 7 11 2
11 16 9 13 13 13 3 2 3 3 13 2
20 13 0 13 2 16 11 13 11 15 1 2 16 11 13 13 13 0 0 9 2
5 12 9 9 13 2
11 7 8 7 9 13 9 13 0 9 9 2
7 13 3 13 15 2 11 2
8 11 13 13 11 9 3 3 2
7 11 13 13 15 10 9 9
4 9 9 13 9
12 13 2 16 3 12 9 13 9 0 11 9 2
2 12 9
11 9 1 13 13 9 2 15 13 9 13 2
3 9 7 9
2 3 0
8 9 13 0 0 7 3 0 2
11 11 9 9 15 16 15 3 13 13 3 2
11 9 13 0 9 2 15 11 10 9 13 2
6 11 13 11 9 3 2
23 0 7 13 2 12 13 9 13 13 2 16 9 13 3 15 13 16 13 15 15 13 15 2
12 0 9 13 9 9 2 15 13 3 9 13 2
14 16 9 13 13 9 9 12 9 9 9 13 13 9 2
14 15 13 16 3 16 15 13 3 9 3 15 15 13 2
4 15 13 0 9
7 15 13 13 9 13 9 13
21 16 10 9 13 13 9 7 9 13 13 9 9 9 2 3 3 11 13 7 13 2
3 9 13 13
6 9 9 13 13 9 2
10 11 13 13 0 0 9 9 0 9 2
14 13 3 3 13 3 13 13 0 0 9 0 0 9 2
5 3 15 13 13 2
7 9 13 0 9 9 12 2
7 11 1 11 13 9 9 2
19 9 13 15 1 3 0 0 9 3 15 1 2 16 15 13 0 0 9 2
7 9 9 13 0 9 7 9
12 9 3 0 2 7 3 0 9 13 13 9 2
24 11 13 3 0 3 3 2 3 9 9 2 9 9 2 9 2 9 7 9 13 10 0 9 2
13 9 15 13 13 9 2 15 9 13 13 3 9 2
8 10 15 13 9 13 13 3 2
3 13 13 2
3 3 7 3
5 11 13 0 9 2
9 9 9 13 3 15 16 9 9 2
6 9 9 13 13 3 2
5 10 9 13 13 2
2 3 16
6 2 15 13 10 9 2
14 9 13 9 2 15 13 11 1 13 0 9 3 13 2
14 3 15 13 13 9 2 16 13 13 10 9 3 3 2
7 0 9 9 13 0 9 2
6 13 13 3 3 9 2
3 9 13 13
12 15 13 3 13 2 16 13 3 13 11 1 2
3 9 13 11
11 2 9 9 13 3 3 9 0 9 13 2
5 9 13 9 9 2
16 9 0 9 13 13 3 9 13 8 8 2 15 3 13 9 2
5 15 13 13 13 13
13 13 13 11 3 3 12 9 2 9 13 13 11 2
3 13 12 1
13 13 13 3 15 2 7 13 3 13 13 10 9 2
9 0 9 7 13 9 9 13 13 2
6 9 13 13 0 3 2
10 9 13 9 9 9 2 3 3 13 2
7 10 9 13 13 0 9 2
10 13 15 15 13 16 15 13 10 9 2
3 0 0 9
10 13 2 16 9 13 9 1 10 9 2
28 9 9 13 13 3 13 0 2 16 0 0 9 13 13 9 1 7 13 2 2 9 2 13 10 9 3 2 2
3 13 0 9
5 15 13 9 3 13
6 15 13 9 12 1 2
5 15 15 15 13 2
4 15 13 0 9
18 7 15 13 3 2 16 9 13 15 2 15 13 9 1 0 9 9 2
10 9 13 12 9 7 13 9 12 9 2
5 9 13 3 13 2
15 9 13 9 1 13 3 0 9 13 9 0 9 9 13 2
5 15 13 15 12 9
3 9 3 13
7 0 7 13 9 7 3 13
8 0 9 11 13 0 13 9 2
11 11 13 2 10 9 9 13 2 15 13 2
7 13 3 3 13 3 9 2
6 15 13 11 1 9 2
13 15 11 3 13 2 13 13 11 11 9 11 11 2
11 9 13 2 3 12 0 9 13 13 9 2
12 9 9 13 3 12 9 0 7 3 13 9 2
11 11 13 3 9 2 7 15 13 0 9 2
11 9 13 9 13 9 9 9 7 13 15 9
4 13 9 9 2
16 10 0 9 13 11 9 11 2 15 1 13 13 9 13 0 2
2 9 13
7 3 13 12 9 9 3 2
7 0 9 13 13 9 3 2
3 13 9 2
12 16 0 13 9 1 2 9 9 13 3 3 2
6 10 9 13 0 9 2
8 11 13 0 9 0 9 7 9
7 13 15 13 15 9 1 2
5 11 13 9 3 2
2 13 13
4 13 0 9 2
8 13 15 3 13 13 9 9 2
7 3 15 13 13 9 12 2
8 15 13 3 13 9 13 9 2
13 12 9 13 3 3 9 2 12 12 13 0 9 2
5 9 13 12 12 9
14 13 3 3 12 11 7 13 2 16 15 13 0 9 2
13 11 9 13 3 0 2 16 11 13 9 11 9 2
3 10 9 9
10 9 13 13 11 9 9 9 9 12 2
13 9 13 13 9 0 9 2 10 9 13 3 0 2
2 13 13
3 2 3 2
7 13 3 10 10 9 3 2
16 9 13 16 15 13 13 15 9 15 3 2 16 15 13 9 2
11 9 13 9 13 9 7 8 16 9 9 2
4 13 9 3 2
4 15 11 13 2
6 13 13 3 12 9 2
4 6 16 13 2
6 15 13 13 1 9 2
3 13 9 0
5 3 2 0 9 2
12 0 7 0 9 13 3 13 0 11 0 11 2
11 15 13 3 3 3 13 0 9 9 9 2
9 3 12 9 9 13 15 13 9 2
9 9 13 3 2 16 13 9 9 2
10 9 13 7 3 15 13 9 9 3 2
13 15 13 13 3 9 7 15 13 7 11 7 11 2
4 15 13 9 2
8 9 13 13 9 9 9 9 2
5 2 13 13 2 2
9 11 13 9 13 3 10 0 9 2
2 9 9
2 9 13
3 13 9 2
10 11 13 9 3 0 7 0 16 11 2
14 9 13 15 2 16 13 0 0 13 9 10 9 1 2
8 9 13 3 0 16 3 11 2
6 9 9 13 3 12 9
4 15 13 13 2
6 0 9 9 11 13 9
10 16 15 13 3 0 2 15 13 3 2
15 3 11 13 13 9 10 0 2 15 15 13 9 13 13 2
14 11 13 3 10 9 1 13 9 9 11 13 11 9 2
17 9 13 13 3 9 2 9 2 16 9 13 9 7 16 9 13 2
8 9 9 13 13 13 0 9 2
16 16 15 13 9 0 9 9 2 3 15 13 3 9 3 3 2
8 3 15 13 16 13 3 9 2
7 15 13 13 16 12 9 2
17 15 13 13 13 3 13 12 9 1 2 13 11 2 7 15 13 2
2 13 3
9 3 9 3 13 9 9 0 9 2
4 13 13 12 9
11 16 0 9 13 0 9 2 15 13 3 2
10 9 13 9 12 3 9 15 13 9 2
17 13 10 9 9 0 2 15 13 9 7 9 9 3 12 9 9 2
4 3 15 13 2
7 0 9 9 9 7 9 9
9 12 9 11 9 13 12 9 9 2
6 13 3 2 3 3 2
10 3 16 15 13 9 2 13 13 13 2
10 9 13 13 13 9 2 7 11 13 2
6 15 13 13 9 9 1
3 10 13 9
11 9 13 13 13 3 3 0 9 7 9 2
2 13 11
20 11 11 13 11 9 12 2 11 11 11 12 13 9 7 11 11 11 9 12 2
3 2 13 2
3 15 13 13
14 12 9 1 0 9 13 3 12 2 10 9 3 12 2
6 15 13 13 9 3 2
2 9 9
5 15 13 0 16 3
13 6 2 13 11 13 9 7 9 2 13 9 13 2
4 12 9 13 0
7 15 13 0 9 9 3 2
19 15 1 13 0 0 9 2 9 2 0 9 2 9 2 9 2 3 15 2
20 11 7 9 11 11 13 3 13 13 9 2 3 9 13 7 13 15 1 9 2
2 13 13
14 3 15 13 3 15 15 1 13 2 3 13 13 3 2
11 11 13 7 13 13 11 0 2 0 9 2
6 9 13 15 11 13 2
2 3 15
11 11 13 13 13 2 15 9 9 13 13 2
8 9 13 3 0 9 9 1 2
5 3 15 13 9 2
5 10 9 13 13 2
6 13 13 10 9 3 2
6 11 13 9 9 9 2
13 10 9 1 9 11 11 13 2 13 11 9 9 2
10 3 7 9 11 13 13 9 3 3 2
4 9 13 3 2
10 16 3 3 13 2 13 13 3 9 2
17 3 9 13 0 2 7 3 0 7 3 10 9 9 13 11 9 2
17 0 9 13 0 9 2 16 15 13 9 3 9 7 15 13 9 2
14 10 9 13 9 2 15 13 0 9 0 9 13 15 2
12 7 3 0 9 13 11 11 2 13 11 11 2
4 13 15 0 2
6 15 13 10 3 0 2
5 3 0 9 13 2
7 3 11 13 9 0 9 2
15 0 2 15 11 13 9 13 2 16 0 9 1 13 9 2
15 0 9 1 13 3 3 13 0 13 9 2 9 7 9 2
5 9 13 1 9 2
9 9 2 15 15 13 2 13 3 0
2 3 16
24 9 9 13 9 3 12 2 12 9 2 7 15 13 9 1 13 13 3 10 9 2 11 13 2
9 13 9 2 13 9 7 13 9 2
9 7 9 13 10 9 9 0 9 2
4 13 15 9 2
13 0 9 0 9 13 13 3 3 16 15 3 13 2
4 13 15 0 2
12 9 1 13 9 7 9 13 13 3 0 13 2
3 13 13 13
5 9 16 3 13 0
6 13 13 9 9 13 2
9 11 8 7 9 13 9 7 9 2
14 15 2 3 9 13 7 9 13 2 9 13 9 9 2
14 15 13 13 2 7 3 2 15 13 2 16 15 13 2
24 9 12 9 9 13 9 15 2 16 11 9 13 13 11 13 9 0 9 11 9 11 11 9 2
9 11 9 13 13 1 9 12 9 2
4 10 9 13 0
4 9 13 7 13
7 13 16 10 9 13 13 2
5 6 16 15 13 2
6 13 3 9 10 0 9
7 0 9 13 3 9 1 2
4 9 13 9 1
2 13 13
8 3 11 9 9 13 11 13 2
18 11 1 10 9 9 13 13 13 9 2 16 9 7 9 9 13 3 2
5 11 9 3 12 9
3 15 3 2
13 3 10 9 10 9 13 2 3 15 9 13 13 2
4 13 15 3 2
5 3 13 13 9 2
12 3 15 3 13 16 9 13 7 13 12 9 2
21 15 13 0 13 15 15 1 2 16 13 13 3 12 9 2 13 3 13 13 15 2
8 12 9 13 7 13 13 9 2
6 6 15 11 13 15 2
13 11 13 13 13 0 10 9 15 0 9 3 13 2
12 15 13 13 12 9 2 13 9 11 1 9 2
2 2 13
8 9 13 9 0 7 0 9 2
2 13 13
8 11 13 13 13 9 13 9 2
5 9 13 13 0 2
16 15 16 9 13 10 9 13 0 9 2 11 13 9 0 9 2
16 16 15 13 13 9 2 9 2 15 3 13 13 9 0 9 2
15 9 13 9 13 13 9 11 11 1 13 9 13 9 9 2
13 0 9 13 2 16 13 13 0 2 3 3 0 2
9 13 0 2 16 15 13 0 9 2
13 13 9 11 11 1 9 13 13 9 10 10 9 2
6 3 15 13 0 0 2
4 0 9 13 2
10 16 11 3 13 2 15 13 0 9 2
4 15 13 0 15
18 15 13 16 3 7 3 9 13 15 7 13 3 2 7 3 15 13 2
15 9 9 9 9 1 3 12 9 9 13 9 7 9 1 2
15 7 9 13 13 15 2 16 13 0 2 7 15 16 13 0
3 13 9 2
8 16 9 13 2 13 13 9 2
6 9 13 0 9 13 2
7 9 13 9 3 16 9 2
2 13 13
11 8 7 9 11 13 3 3 16 9 13 2
5 9 13 9 9 2
2 13 13
6 3 13 3 13 9 2
2 9 2
3 9 13 9
9 9 13 3 16 9 13 3 9 2
10 15 13 3 7 3 13 7 9 1 2
14 9 0 11 9 13 15 13 9 12 9 9 1 12 2
4 15 13 9 2
7 13 15 10 9 13 13 2
6 7 13 15 0 9 2
10 13 0 0 9 2 16 9 13 13 2
15 16 9 13 12 9 9 2 13 3 13 15 2 7 13 2
11 9 13 9 13 9 2 15 9 13 13 2
5 15 13 13 9 2
2 0 2
4 9 13 12 2
6 13 13 13 3 13 2
3 9 13 0
6 9 9 13 12 9 2
8 9 13 13 13 0 0 9 2
5 13 9 0 9 2
13 11 13 0 9 16 11 7 11 7 0 16 11 2
9 0 0 9 13 13 3 12 9 2
7 9 13 9 3 13 1 2
8 3 9 13 12 7 12 9 2
11 11 9 13 0 7 15 13 10 1 9 2
5 9 13 9 1 2
7 3 13 9 1 0 9 2
16 3 15 13 9 9 9 2 3 15 13 13 9 7 13 9 2
5 13 15 3 13 2
9 3 13 9 1 15 13 13 13 2
3 9 9 11
3 15 13 15
10 3 15 13 0 2 16 13 15 13 2
14 13 13 11 2 13 9 2 15 3 13 3 16 11 2
7 3 15 13 13 9 16 2
5 9 13 13 0 2
7 3 9 13 11 1 13 2
6 0 2 3 13 9 1
21 9 13 3 15 1 16 11 9 11 13 13 2 16 11 9 13 9 13 3 0 2
5 3 3 13 13 2
5 13 9 0 9 2
5 13 3 15 0 2
9 15 13 13 10 9 10 9 1 2
7 9 13 3 3 0 7 0
3 10 9 2
11 15 13 0 9 2 16 13 0 13 13 2
11 13 0 16 11 9 13 9 3 10 12 2
9 6 2 3 11 13 13 3 0 2
2 10 9
7 11 13 9 1 11 11 2
4 13 9 3 2
9 13 3 9 3 7 13 13 9 2
10 15 13 13 9 2 11 13 9 9 2
17 13 3 0 13 2 16 13 9 13 9 2 16 13 3 9 13 2
6 3 0 0 7 0 9
25 3 3 2 3 13 13 16 15 11 11 7 11 11 13 3 0 9 9 16 11 11 7 11 11 2
10 3 16 15 13 3 12 9 2 7 2
6 13 10 9 13 13 2
7 3 15 3 13 9 13 2
3 9 13 9
5 3 15 13 9 2
2 10 3
11 0 9 15 13 0 9 3 0 16 13 2
16 9 9 11 11 13 12 7 13 12 9 1 9 7 0 9 2
8 12 9 1 9 16 13 12 2
15 13 13 10 9 9 2 16 13 13 9 9 2 15 13 2
7 3 3 13 9 7 9 2
3 9 13 13
18 11 11 7 11 9 11 13 3 9 9 1 7 10 9 11 9 13 0
13 0 9 13 11 0 9 13 9 2 9 7 9 2
11 9 13 3 7 3 3 9 13 9 0 2
9 15 13 3 3 0 7 0 9 2
14 0 9 13 3 2 16 15 13 9 0 9 13 9 2
5 9 0 15 13 2
19 0 9 9 9 13 3 13 11 9 0 0 9 2 15 13 13 13 13 2
2 13 9
9 15 13 13 13 12 9 13 15 2
11 9 1 11 13 9 13 9 11 7 11 2
5 3 13 13 9 2
6 0 9 2 11 13 2
16 13 13 13 10 9 2 7 16 13 3 9 11 9 7 3 2
8 0 9 13 0 9 9 9 2
16 9 9 13 9 2 15 13 13 13 9 10 3 0 9 9 2
12 2 2 3 16 15 7 15 15 1 13 13 2
5 3 15 13 13 2
11 11 9 9 9 13 9 9 13 0 9 2
6 13 15 0 9 9 2
6 13 13 0 9 9 2
7 11 13 10 9 16 11 2
16 15 13 15 15 13 3 3 2 7 15 13 0 9 15 1 2
20 16 11 13 9 13 3 13 13 2 9 9 13 0 9 0 11 2 9 2 2
5 3 9 13 9 2
17 9 12 9 1 13 12 9 13 13 9 13 3 12 12 9 9 2
19 13 9 13 3 0 2 13 0 0 0 9 7 13 0 9 3 13 9 2
8 13 15 3 2 15 13 3 2
4 11 13 11 2
10 3 13 0 9 13 2 2 8 2 2
5 3 13 10 0 9
2 13 13
6 15 13 3 12 9 2
6 9 13 9 7 9 2
14 9 9 13 13 9 0 9 2 15 13 9 12 9 2
6 7 15 13 13 15 2
2 7 3
8 11 13 15 13 9 9 13 2
3 2 3 2
7 9 9 9 13 3 3 2
14 13 2 16 9 13 3 9 13 7 3 3 13 9 2
7 9 13 3 9 12 9 2
10 13 2 16 9 13 0 15 15 13 2
3 9 1 9
2 13 3
3 9 13 13
5 9 9 13 9 13
10 0 0 13 15 9 1 11 8 9 2
8 13 9 2 16 13 10 9 2
3 3 3 2
15 9 11 11 7 9 11 11 13 0 9 3 9 7 9 2
15 9 13 0 13 3 2 3 3 2 7 9 13 12 9 2
2 6 9
3 15 13 2
10 13 9 3 9 7 13 0 9 15 2
7 9 13 3 9 9 12 2
8 7 16 15 13 13 10 9 2
8 13 3 3 3 2 11 13 2
7 9 13 0 9 7 9 2
6 15 13 3 9 9 2
10 13 9 2 16 9 9 13 3 0 2
14 7 9 13 3 2 16 15 13 3 0 0 13 11 2
7 10 0 13 3 3 13 2
6 3 15 13 7 13 2
12 13 9 7 13 13 9 2 3 15 9 3 2
12 9 13 13 11 2 10 9 9 0 9 13 2
5 3 15 13 9 2
9 13 0 13 10 9 0 9 1 2
13 9 13 0 9 3 3 2 16 9 15 3 13 2
4 13 15 15 2
14 9 2 15 15 13 13 9 13 2 13 13 13 9 2
9 13 10 11 3 3 9 10 9 2
10 7 3 2 13 3 13 15 1 3 2
8 9 13 3 13 9 13 9 2
3 3 3 2
4 15 13 13 9
9 13 9 7 9 13 9 13 0 2
12 11 13 2 16 15 13 3 9 3 15 1 2
17 10 9 13 9 9 13 3 13 2 16 13 15 10 0 9 13 2
14 13 0 13 3 0 2 16 9 13 15 15 3 0 2
2 13 9
17 15 13 3 13 9 0 9 2 15 9 1 13 9 0 9 9 2
13 15 13 13 2 16 10 9 13 0 10 9 9 2
9 3 13 12 9 12 13 13 9 2
3 11 3 9
19 16 11 13 9 11 13 15 0 9 9 8 7 9 2 13 3 0 16 2
10 13 13 9 2 16 10 9 9 13 2
10 0 13 3 0 9 10 9 1 9 2
13 16 3 0 9 13 0 13 10 9 0 9 9 2
4 13 9 3 2
5 11 13 0 9 2
9 3 9 13 10 9 7 13 9 2
9 9 13 3 0 7 13 3 9 2
9 9 15 13 13 2 11 9 13 2
16 9 13 9 3 2 2 11 13 15 13 2 15 15 13 2 2
6 10 9 15 3 13 2
3 13 15 2
13 3 3 15 15 13 2 13 3 3 15 15 13 2
4 6 16 0 2
15 0 9 1 13 0 2 16 9 13 7 13 0 9 9 2
11 11 13 13 9 2 3 16 3 13 13 2
4 13 13 13 2
9 15 13 9 2 15 13 9 0 2
9 0 0 9 10 12 3 13 9 2
7 9 0 9 13 10 3 2
9 10 9 13 3 13 13 3 0 2
4 9 13 2 2
5 9 13 9 9 2
3 9 9 0
8 9 9 13 0 12 12 9 2
20 15 13 3 9 9 9 12 9 1 7 15 13 3 0 9 11 9 9 9 2
4 15 13 9 2
7 15 13 11 9 11 9 2
7 15 13 0 9 12 9 2
10 9 11 11 8 8 13 13 12 9 2
11 9 13 13 13 7 13 3 3 0 9 2
8 3 3 3 6 3 3 13 2
9 10 9 13 3 0 13 16 9 2
2 3 3
13 16 3 13 2 16 13 13 2 13 13 9 13 9
5 3 10 0 9 2
10 13 3 13 0 9 13 3 15 13 2
5 13 13 10 9 2
8 11 13 10 9 10 11 9 2
6 13 9 2 16 9 13
9 9 13 9 2 7 9 13 9 2
13 10 9 2 15 3 11 9 13 13 9 12 9 2
5 13 13 0 9 2
16 9 13 0 7 0 9 2 15 9 13 9 11 3 0 9 2
6 11 9 15 13 12 2
9 0 9 9 13 13 0 0 9 2
16 9 11 13 10 9 1 10 9 15 2 16 9 13 13 9 2
9 9 13 13 3 16 9 13 15 3
10 10 0 9 9 15 13 3 9 3 2
12 3 13 9 13 0 9 9 2 9 7 9 2
5 9 15 13 13 9
6 9 9 12 11 9 9
13 0 9 9 13 13 3 9 12 9 7 12 9 2
14 11 13 3 9 1 9 10 11 9 1 13 0 9 2
5 7 15 15 13 2
9 9 13 13 2 7 9 13 13 2
5 9 9 13 3 2
6 15 13 3 13 9 2
6 9 13 3 3 13 2
10 0 9 13 13 0 9 0 0 9 2
4 9 13 15 9
5 3 12 9 9 2
7 13 3 13 3 10 9 2
9 3 2 7 3 15 13 3 9 2
9 3 13 0 13 9 9 9 1 2
5 15 13 3 0 9
9 9 7 9 13 13 13 0 9 2
6 11 13 3 9 11 2
8 11 9 13 0 0 13 15 2
9 15 13 3 16 15 13 9 15 3
6 11 13 9 0 9 2
12 0 9 9 13 1 15 13 9 8 7 9 2
2 0 9
5 13 9 3 9 2
5 2 6 13 3 2
4 9 13 9 2
5 15 13 13 3 2
11 9 13 9 12 9 9 12 1 9 11 2
11 15 13 0 12 9 13 9 13 0 9 2
13 9 15 13 3 10 0 9 9 2 15 13 15 2
5 15 15 3 13 2
3 15 13 2
11 0 13 0 9 13 13 3 11 9 1 2
6 13 9 13 3 9 2
11 9 9 13 13 13 3 3 16 9 13 2
4 13 13 13 2
17 13 0 0 9 7 15 2 16 15 7 15 13 3 15 15 13 2
6 13 13 3 9 12 1
15 0 9 13 15 16 11 11 7 3 9 13 11 9 9 2
3 15 13 2
5 2 15 13 9 2
6 11 9 13 3 9 2
2 3 9
6 13 13 3 9 11 2
14 15 15 13 2 9 1 9 1 9 2 9 7 0 2
7 9 13 3 2 0 3 2
3 13 13 13
18 9 13 3 2 13 9 13 7 13 9 12 0 9 11 7 11 1 2
4 9 13 15 13
10 11 9 9 13 0 9 0 12 9 2
8 12 9 10 12 9 13 15 2
9 16 9 13 0 2 13 13 9 2
12 13 13 13 13 9 9 13 3 9 7 9 2
8 3 13 13 13 3 9 13 2
14 15 15 1 13 9 3 16 13 9 2 15 15 13 2
9 9 2 13 3 0 2 13 0 2
9 3 11 9 13 3 3 0 9 2
8 9 13 0 9 11 9 9 2
4 10 9 13 0
8 0 9 13 9 13 9 9 13
3 15 13 2
8 13 3 0 9 13 13 9 2
9 9 13 9 13 9 13 3 9 2
8 11 11 13 3 9 7 9 2
6 15 13 13 9 9 2
4 13 13 13 9
5 15 13 0 3 0
7 9 9 13 11 13 11 2
11 3 13 13 2 16 13 13 3 15 9 2
11 9 1 9 0 9 13 13 9 2 15 2
11 9 9 13 13 12 12 7 9 12 12 2
8 9 13 9 9 7 9 9 2
3 9 7 9
6 9 13 9 13 3 2
8 15 3 13 13 9 3 9 2
3 9 13 2
23 15 13 3 2 16 9 13 3 3 3 2 16 15 13 3 13 3 3 0 13 3 3 2
8 13 3 13 15 12 9 0 9
7 10 9 13 3 0 9 2
16 12 3 13 9 13 13 3 10 9 16 15 15 13 9 3 2
4 11 3 13 11
21 3 3 10 9 13 3 2 16 13 9 13 3 10 9 2 16 15 13 9 9 2
6 13 2 16 13 3 2
11 13 3 0 2 16 9 13 15 0 9 2
10 3 13 9 13 13 11 9 7 9 2
3 9 9 2
14 9 9 13 0 9 2 3 10 9 9 13 9 9 2
16 0 9 11 11 13 3 9 12 9 0 7 3 3 3 11 2
7 9 9 13 9 7 9 2
10 0 9 13 9 13 3 3 0 9 2
9 13 9 13 13 7 3 13 3 2
8 15 13 9 13 3 9 12 2
3 13 13 9
8 9 9 13 11 7 11 11 2
10 13 3 10 9 15 15 13 13 10 9
7 0 7 0 9 13 13 2
8 15 13 3 9 3 9 1 2
12 15 13 15 3 10 10 9 1 2 3 11 2
6 9 9 13 3 13 2
18 15 13 3 3 13 13 7 13 3 13 9 15 3 15 13 3 13 2
8 0 0 13 9 11 11 9 2
4 15 13 9 2
11 11 11 11 13 0 9 7 9 10 9 2
16 15 13 2 16 10 9 9 13 3 2 16 13 9 9 1 2
9 9 13 15 9 7 9 13 9 2
9 13 3 3 2 13 3 3 9 2
13 9 13 9 0 9 2 15 13 13 9 12 9 2
7 15 1 9 13 7 13 2
12 15 12 2 3 3 12 13 13 15 16 9 2
15 15 1 11 7 11 13 9 2 3 15 3 13 13 9 2
3 9 9 2
10 13 0 9 0 11 13 13 3 13 2
2 0 9
22 7 13 3 9 2 16 13 13 9 2 16 11 9 1 13 3 13 3 9 15 1 2
5 13 9 16 13 15
11 15 13 3 3 9 0 16 10 9 3 2
17 11 13 9 12 2 7 11 13 12 0 9 2 13 9 7 9 2
3 3 7 3
2 15 1
12 9 1 15 13 13 0 13 9 10 9 1 2
6 15 13 0 9 13 9
3 13 13 2
3 15 13 13
8 9 13 3 13 2 16 13 15
5 13 13 3 9 2
3 13 11 2
8 3 13 9 7 9 0 9 2
6 15 13 3 0 9 2
7 0 9 13 0 16 0 2
6 13 15 10 0 9 2
6 11 2 0 9 15 2
5 15 13 11 11 3
6 15 13 13 15 1 2
13 3 16 15 13 10 9 2 15 13 13 13 3 2
4 12 9 0 9
11 13 13 3 3 3 13 10 9 3 3 2
8 9 15 13 9 7 12 9 2
11 9 9 13 13 12 9 2 7 12 9 2
3 13 13 2
14 11 13 3 3 3 7 3 9 2 0 9 3 13 2
10 0 9 13 0 9 0 7 0 9 2
3 11 9 9
6 9 11 11 13 11 9
4 13 9 13 9
6 11 13 9 12 9 2
3 11 13 9
21 3 13 3 9 2 16 11 13 15 2 3 3 11 13 13 7 13 2 13 3 2
12 15 15 13 0 7 15 2 13 13 10 9 2
12 11 13 3 13 9 7 13 3 9 9 13 2
10 15 13 2 16 15 0 13 0 9 2
18 16 9 9 13 9 2 9 13 13 13 9 1 2 15 13 3 13 2
13 16 9 13 0 2 15 13 0 0 9 9 13 2
8 15 13 11 13 10 9 13 2
2 10 9
16 11 13 0 9 9 8 2 8 2 8 2 8 7 9 9 2
11 7 16 11 13 9 1 2 3 13 13 2
5 15 13 3 10 0
10 11 13 3 10 9 2 13 9 0 2
3 13 9 9
9 9 9 11 2 11 13 9 3 2
9 9 7 9 13 15 1 0 13 2
6 9 13 9 1 11 2
11 9 13 2 7 3 12 7 11 1 11 2
5 15 13 3 3 13
10 11 13 13 9 0 9 0 0 9 2
2 6 0
17 11 11 13 10 9 12 10 0 9 0 9 2 3 13 3 9 2
6 6 3 0 15 13 2
12 3 3 11 2 13 2 9 7 9 13 9 2
10 0 9 13 3 12 9 2 13 11 2
11 0 9 13 13 2 16 9 13 11 10 9
13 15 13 13 3 13 12 10 9 2 13 9 9 2
3 13 3 2
3 13 9 1
8 11 9 13 3 3 0 13 2
11 11 13 10 0 3 3 7 3 9 9 2
7 9 13 15 2 11 13 2
17 9 9 7 9 9 15 3 13 9 1 9 9 3 0 9 13 2
6 15 13 9 9 13 2
4 13 13 9 3
10 6 13 15 2 13 15 13 13 3 2
11 15 13 2 7 15 15 2 9 0 9 2
6 15 13 3 13 0 2
4 13 13 13 13
9 9 13 13 10 9 9 7 9 2
3 13 13 15
4 9 13 9 2
18 9 7 0 9 13 0 9 15 10 9 2 3 13 13 9 12 9 2
8 13 9 3 9 3 13 9 2
3 0 9 9
4 9 13 9 9
3 15 13 2
9 3 11 13 0 9 7 13 3 2
5 9 13 15 13 2
23 3 15 13 2 16 9 13 13 1 9 3 16 13 2 16 9 13 0 2 9 13 9 2
5 13 9 9 0 9
14 16 13 9 2 9 13 13 2 16 3 13 10 11 2
6 9 15 13 13 3 2
11 0 9 3 13 9 0 3 3 7 13 2
3 13 12 9
6 13 3 0 7 13 2
4 9 13 11 0
3 3 13 2
7 0 9 15 13 13 3 2
12 3 2 10 3 13 0 9 2 3 3 13 2
10 11 12 9 9 12 12 9 13 0 2
2 10 9
6 9 13 13 3 11 2
5 9 1 13 3 2
2 3 3
5 13 0 7 0 2
4 11 11 13 9
8 16 13 13 10 9 7 13 2
7 9 13 2 16 9 13 2
5 15 13 3 15 2
6 15 13 3 9 13 2
10 11 11 13 0 2 0 7 0 9 2
5 9 13 13 0 9
5 3 9 9 13 2
9 16 13 9 2 13 3 3 3 2
2 9 9
8 9 2 13 13 15 9 11 2
6 9 13 7 9 13 2
18 9 1 0 9 13 9 13 3 3 10 9 16 13 0 9 7 9 2
10 3 3 13 3 12 12 9 0 9 2
7 3 13 13 9 3 12 2
9 9 13 9 9 3 13 16 9 2
9 9 3 13 13 11 7 11 3 2
11 15 13 15 13 7 0 9 1 15 13 2
5 3 0 9 0 2
3 13 9 9
2 13 13
9 9 13 3 12 9 2 3 9 2
5 15 13 15 1 2
7 16 9 13 2 15 13 2
14 2 3 10 3 15 13 13 2 2 11 13 13 11 2
13 16 11 13 2 3 13 11 9 9 13 13 9 2
2 13 9
8 12 0 9 13 3 11 9 2
23 7 3 0 13 15 9 13 10 9 3 3 2 16 9 13 13 3 13 12 12 9 1 2
13 15 13 13 3 0 16 15 11 3 13 13 13 2
6 3 9 13 9 9 2
10 11 13 13 9 7 15 3 9 3 2
15 9 13 3 0 2 9 13 13 0 2 0 15 3 13 2
3 0 0 9
10 10 9 13 0 2 0 9 13 9 2
8 3 10 9 13 13 0 9 2
8 11 13 13 3 10 9 9 2
9 0 11 13 7 13 7 13 9 2
15 15 3 13 13 0 9 1 2 7 9 13 3 0 9 2
18 9 13 3 7 3 3 2 13 9 13 9 7 3 10 9 16 13 2
11 13 13 2 3 13 2 16 13 9 9 2
5 10 9 13 9 2
18 16 9 10 9 13 0 7 9 13 3 2 9 13 11 3 3 0 2
5 9 13 9 1 2
2 13 3
13 9 9 9 9 13 9 9 7 0 9 0 9 2
2 3 12
9 11 9 13 13 0 0 9 9 2
4 9 13 9 2
29 7 3 3 13 10 3 0 9 9 7 3 13 13 3 16 13 10 9 3 3 16 16 16 3 10 10 9 13 2
12 6 3 15 2 13 11 11 7 9 11 11 2
10 9 13 9 9 13 12 12 12 9 2
7 9 13 0 12 12 9 2
11 15 13 0 0 9 7 15 13 3 0 2
20 9 9 2 7 13 15 10 9 13 3 16 13 13 10 9 0 2 3 9 2
16 10 9 9 9 13 13 1 0 11 9 11 2 11 11 1 2
19 13 13 2 13 3 3 16 15 10 9 2 0 0 2 9 7 9 13 2
10 9 13 3 3 2 7 13 9 0 2
12 15 13 3 11 2 13 15 3 13 3 3 2
4 13 9 3 2
27 15 13 12 9 9 15 15 13 9 2 9 2 9 7 9 2 15 15 13 2 13 7 13 9 1 9 2
6 9 13 9 13 9 2
3 9 13 3
7 15 13 9 13 0 9 2
7 3 13 3 13 13 0 9
3 9 3 1
10 12 9 1 10 9 13 13 10 9 2
4 13 3 0 2
7 13 15 3 13 15 9 2
7 15 13 13 13 3 3 2
19 15 13 13 9 2 16 16 9 13 9 9 3 2 9 13 3 9 3 2
11 9 13 0 13 11 1 2 3 9 11 2
1 12
6 12 13 13 13 13 9
6 11 13 13 9 9 2
3 3 13 9
2 10 9
5 13 12 12 9 2
6 0 9 13 13 13 2
9 9 13 13 9 3 1 0 9 2
1 3
4 10 12 0 9
21 11 13 9 2 16 9 13 13 2 15 13 11 1 11 2 13 11 7 13 9 2
5 11 13 13 0 9
6 13 15 13 3 0 2
2 13 3
7 2 15 13 13 10 9 2
7 7 13 15 3 3 9 2
9 15 13 13 9 9 1 13 9 2
3 3 0 9
11 0 9 13 3 13 13 9 7 10 9 2
13 16 13 0 2 0 7 0 2 3 13 9 1 2
7 13 13 9 1 0 9 2
6 11 9 2 0 11 9
12 9 7 9 13 9 2 7 3 3 0 9 2
4 9 13 15 3
17 13 13 3 3 2 7 13 9 13 9 3 0 0 8 7 9 2
13 9 7 9 13 15 7 15 1 13 13 0 9 2
4 13 15 0 2
7 16 15 13 8 0 0 13
2 0 9
13 15 13 3 13 13 15 2 16 13 3 0 9 2
13 15 13 13 10 10 9 2 13 13 3 13 0 2
2 11 11
14 3 15 13 3 7 13 13 15 2 15 13 15 13 2
5 13 15 9 3 2
6 11 13 13 3 13 2
6 9 13 13 15 9 2
14 13 9 2 9 7 9 13 9 1 3 9 7 9 2
4 9 13 9 2
3 12 9 13
11 0 13 11 7 11 10 3 16 3 9 2
8 3 13 13 3 3 13 9 2
2 13 13
18 2 0 13 3 9 2 7 15 7 12 0 13 3 2 2 15 13 2
9 13 15 13 16 0 9 13 3 2
5 3 3 12 9 1
16 15 13 9 2 16 9 13 13 9 2 16 9 15 13 0 2
16 11 13 10 9 9 2 16 10 9 13 13 3 15 13 9 2
12 9 0 9 13 13 3 13 3 9 1 11 2
10 13 3 0 2 7 13 13 3 13 2
18 13 3 11 13 15 13 2 7 15 15 13 15 2 7 3 15 13 2
5 10 9 3 13 2
10 9 13 3 0 7 13 15 1 3 2
9 15 9 13 9 2 9 7 9 2
30 15 13 15 0 2 7 13 0 0 2 15 13 15 1 9 13 13 16 2 15 9 12 13 13 3 12 12 0 11 2
14 3 9 13 12 9 1 12 9 1 7 13 0 9 2
4 15 13 0 2
7 16 9 13 13 3 3 2
9 13 13 13 9 3 16 0 9 2
7 0 9 13 9 7 9 2
15 15 0 7 0 13 3 3 2 16 13 10 9 13 9 2
6 11 13 3 13 11 2
15 16 9 11 0 9 15 13 2 3 15 15 13 9 9 2
22 3 16 9 6 16 16 15 13 13 9 9 3 15 13 16 6 15 13 13 3 15 2
11 9 2 15 13 3 9 2 13 3 0 2
8 9 12 1 9 13 9 9 2
6 9 13 3 13 9 2
17 11 9 9 11 11 7 11 9 13 11 13 12 9 9 0 9 2
5 13 9 9 12 9
10 11 13 13 2 13 15 13 7 13 2
10 11 13 11 0 7 10 11 0 9 2
3 13 3 2
14 15 13 2 16 9 13 3 2 9 13 2 9 13 2
16 12 9 1 13 9 9 1 3 13 15 16 9 9 0 9 2
17 1 9 3 13 0 0 9 2 7 15 13 0 9 7 12 9 2
10 15 13 9 3 3 12 9 3 9 2
10 10 9 15 13 13 3 0 9 3 2
5 13 9 13 9 2
6 13 3 9 3 2 13
7 15 13 9 9 12 9 2
11 9 13 13 3 2 15 13 15 1 0 2
11 9 11 13 0 7 0 2 7 3 0 2
5 13 15 9 13 2
13 16 13 13 15 0 9 2 15 13 13 3 0 2
5 15 13 9 9 2
17 3 13 9 13 3 13 0 16 13 2 7 15 13 3 0 9 2
8 15 13 13 10 9 0 9 2
7 9 9 13 3 12 9 2
6 15 13 11 13 9 2
3 9 13 9
6 13 10 11 11 13 2
6 9 13 13 11 9 2
2 9 9
4 15 13 9 2
12 11 1 13 13 13 10 9 9 15 13 9 2
5 9 13 13 9 2
13 13 0 2 16 13 9 2 9 9 7 15 9 2
4 3 3 15 2
6 3 13 0 13 9 2
14 15 13 2 16 3 13 15 13 0 13 9 9 13 2
6 15 13 0 13 9 2
2 9 1
12 9 13 13 0 13 9 7 9 3 15 1 2
9 16 3 0 9 9 2 15 13 2
14 13 15 3 2 16 0 9 0 9 13 3 13 12 2
12 11 1 13 13 13 9 1 9 13 13 0 2
13 6 15 13 13 15 3 3 0 7 13 16 9 1
6 15 13 10 0 9 2
9 16 9 13 2 15 13 10 9 2
3 3 13 9
8 11 13 13 3 0 0 9 2
12 9 13 9 12 1 11 7 11 0 9 12 2
11 15 13 2 16 9 9 13 0 9 0 2
2 13 13
8 9 13 7 9 13 15 9 2
4 3 10 13 9
8 13 9 13 3 13 10 9 9
10 9 1 9 9 13 13 9 13 9 2
10 12 9 15 13 2 15 13 0 2 2
8 9 13 3 0 2 15 13 2
3 13 3 2
3 9 13 9
13 15 15 13 9 9 2 7 15 13 3 3 9 2
11 15 13 9 9 9 9 13 0 0 11 2
14 11 9 13 3 10 9 2 15 13 9 9 7 9 2
9 11 13 13 9 7 9 16 9 2
18 9 9 13 9 13 11 9 9 9 13 9 9 9 7 11 0 9 2
11 9 13 9 13 3 2 16 13 3 7 3
2 9 9
8 15 13 13 9 2 15 9 2
7 10 12 9 13 3 9 2
8 15 13 3 16 15 13 15 2
8 13 13 3 3 3 13 13 2
6 15 13 9 9 12 2
15 12 0 9 13 12 9 7 10 0 9 2 2 9 2 2
20 16 13 15 2 16 13 12 9 13 8 7 9 1 2 3 13 15 15 13 2
8 3 10 9 13 13 9 9 2
12 3 3 13 9 9 2 7 15 3 13 9 2
8 7 3 15 0 9 3 13 2
13 3 15 13 13 9 2 15 13 9 15 13 9 2
5 15 13 9 11 2
9 15 13 3 12 9 9 9 12 2
7 9 13 12 13 9 15 2
3 9 13 3
12 10 9 13 2 10 9 0 9 13 9 9 2
7 15 13 13 9 7 9 2
15 11 13 9 13 0 9 1 2 10 9 13 15 3 13 2
7 8 2 8 7 3 10 9
2 11 9
12 9 13 0 9 3 9 9 9 0 9 11 11
4 3 15 9 2
2 0 9
5 11 12 9 9 2
8 12 12 0 9 9 13 11 2
5 15 13 16 9 2
10 15 1 9 13 0 13 9 1 0 2
5 10 0 9 13 2
7 11 7 11 13 9 12 2
7 11 13 9 2 7 3 15
11 16 15 13 10 11 1 16 15 13 3 2
12 11 13 3 13 7 11 3 13 0 9 9 2
6 13 3 13 10 9 2
20 13 13 9 9 7 13 10 9 13 3 15 15 13 2 16 15 13 13 9 2
6 9 13 3 3 0 2
7 9 13 12 9 1 11 2
13 11 13 2 16 9 11 9 13 13 3 11 9 2
11 0 2 0 9 13 13 3 9 1 9 2
18 16 11 13 11 0 9 2 15 13 3 13 15 2 16 13 13 13 2
6 3 15 13 11 3 2
29 13 13 0 0 9 2 0 9 2 15 13 10 0 2 0 2 0 7 0 0 2 3 0 2 13 0 13 9 2
8 3 13 0 13 12 12 9 2
13 10 9 15 13 15 0 2 16 9 13 9 9 2
12 3 15 13 2 3 9 9 11 13 9 9 2
5 9 9 13 9 2
2 3 9
4 13 13 3 3
8 15 13 0 7 15 13 0 2
8 0 9 13 3 12 0 9 2
6 15 13 3 3 9 2
4 9 0 0 9
3 15 13 3
11 7 15 13 13 3 0 13 15 9 7 9
3 3 13 9
10 3 13 9 9 13 3 10 9 9 2
7 13 15 10 9 13 9 2
5 11 9 9 13 9
6 13 15 3 3 13 2
10 2 16 13 15 13 15 15 13 15 2
11 11 11 13 9 3 0 7 0 9 1 2
15 13 3 9 13 13 3 9 13 2 3 9 13 13 9 2
8 9 9 13 0 10 9 13 2
14 9 13 9 9 9 2 9 9 9 7 9 3 9 2
9 9 13 13 9 2 13 0 9 2
6 9 9 13 9 0 2
12 13 3 2 16 9 8 7 9 13 3 3 2
2 13 12
11 11 9 13 0 9 13 3 13 9 11 2
8 13 13 3 3 3 7 3 2
9 15 13 3 3 11 10 11 1 2
7 9 9 9 11 11 11 3
5 0 9 13 3 2
7 10 9 7 3 0 9 2
12 11 13 10 9 2 16 7 15 7 11 13 2
11 15 16 15 13 9 9 7 9 13 9 2
23 1 0 9 2 9 9 7 0 0 9 9 12 0 12 0 13 15 1 16 9 12 3 2
5 13 3 13 10 9
6 15 13 13 9 9 2
11 3 12 0 9 13 9 13 3 0 9 2
6 9 13 13 0 9 2
3 13 0 9
6 11 13 11 7 9 2
6 10 0 13 13 0 2
8 3 13 9 13 0 0 11 2
10 3 9 13 3 16 13 9 15 1 2
7 13 9 9 7 13 13 2
5 15 13 15 13 2
5 9 13 3 9 2
5 9 13 12 9 2
14 0 13 3 0 0 9 13 2 15 3 13 9 1 2
8 3 13 9 7 3 13 9 2
7 9 13 9 9 10 9 2
10 0 9 10 15 13 7 13 9 9 2
5 13 9 3 13 2
15 9 13 13 9 2 15 13 9 3 2 3 7 3 13 2
16 9 2 12 1 13 9 9 9 2 3 9 2 13 0 9 2
6 9 13 13 13 9 2
8 13 10 15 3 13 13 9 2
13 9 9 13 13 2 9 3 13 2 13 7 13 2
3 9 13 0
11 11 11 9 13 3 9 12 9 13 9 2
7 11 7 11 13 10 9 2
8 11 9 1 15 13 15 13 2
11 3 10 9 15 13 2 15 9 13 13 2
9 11 13 9 3 9 13 9 11 2
19 0 0 9 0 9 11 1 13 9 12 2 16 9 13 9 13 9 9 2
3 13 15 2
4 8 7 0 9
5 9 13 13 13 2
5 11 13 9 9 2
8 9 13 13 9 7 9 13 2
3 13 13 13
12 10 9 13 9 9 0 9 2 9 7 9 2
2 0 9
5 0 9 13 13 2
5 15 13 13 3 2
7 3 3 13 11 7 11 2
7 15 13 13 3 0 9 2
7 16 15 13 0 0 3 2
8 0 9 0 13 9 3 3 2
5 3 0 9 13 13
11 3 9 13 9 13 2 7 3 9 13 2
10 9 13 0 9 9 9 1 13 9 2
5 0 13 3 9 2
4 13 15 3 2
14 9 11 11 13 13 11 2 7 9 11 11 13 3 2
8 15 13 13 9 3 7 3 2
11 9 13 13 3 9 12 7 12 0 9 2
22 15 13 13 10 9 3 0 9 16 13 2 15 1 2 16 10 9 11 13 3 0 2
8 10 9 13 12 9 13 11 2
5 15 13 9 13 2
13 3 9 15 13 3 9 9 9 7 13 3 3 2
10 15 13 2 3 9 13 13 3 9 2
4 15 13 0 2
12 7 3 16 9 13 3 9 13 3 7 2 2
9 15 13 3 3 3 2 3 3 2
13 9 9 13 13 3 9 7 0 9 13 3 9 2
6 9 13 3 9 13 2
8 11 7 9 13 15 12 9 2
3 3 13 2
4 9 13 3 2
17 9 9 7 9 9 13 13 3 0 16 9 9 9 9 13 13 2
7 3 9 13 9 1 9 2
7 11 2 13 15 10 9 2
4 9 13 0 2
9 9 12 13 3 9 7 9 9 2
7 15 3 13 13 2 11 2
9 11 13 12 9 9 13 3 0 2
3 0 0 9
4 13 11 9 2
7 9 13 13 3 7 3 2
11 13 3 3 2 16 13 9 13 0 9 2
15 10 9 13 9 3 15 13 3 2 16 9 9 13 9 2
8 9 13 16 13 0 3 3 0
4 13 0 16 13
11 0 9 13 13 13 2 16 9 13 13 2
13 11 9 9 13 13 3 0 2 16 13 3 0 2
11 9 1 13 3 13 13 0 9 7 9 2
6 10 9 13 0 9 2
6 10 9 13 0 9 2
12 9 13 15 9 9 2 7 15 13 0 9 2
6 15 13 16 15 13 12
10 13 2 16 9 9 13 13 11 9 2
8 11 13 11 7 11 9 1 2
2 0 9
3 13 3 2
22 7 16 3 15 13 2 16 13 9 13 10 9 2 3 3 13 0 9 9 11 9 2
5 15 13 15 9 2
5 15 13 13 9 2
5 15 13 13 3 2
4 9 13 9 2
7 3 15 13 9 10 9 2
5 3 13 11 9 2
2 13 9
5 9 13 9 13 2
6 0 15 13 13 13 2
12 13 13 13 3 0 9 7 13 13 3 9 2
6 10 9 13 10 9 2
3 12 9 0
7 12 9 13 15 13 9 2
6 9 7 9 9 7 9
10 1 9 9 11 13 11 9 9 9 2
11 0 13 13 15 13 0 9 7 9 9 2
12 15 13 2 16 3 15 13 2 9 0 9 2
12 9 13 13 9 1 9 2 16 9 13 9 2
9 15 16 13 10 9 2 3 11 2
14 13 2 16 3 15 15 2 11 13 9 0 9 1 2
8 15 13 0 16 13 9 9 2
13 15 13 9 2 15 9 9 2 15 9 13 13 2
8 0 13 13 2 15 9 13 2
9 11 9 13 3 10 11 0 0 2
2 0 9
5 9 13 11 9 2
2 13 9
6 15 13 13 11 9 2
9 15 3 13 16 16 13 3 3 13
5 15 13 10 9 2
4 9 7 9 9
3 2 6 2
3 13 3 2
4 13 1 9 2
8 9 13 9 7 0 9 13 3
5 11 13 13 9 2
15 0 9 13 0 2 0 9 2 10 9 13 3 12 9 2
10 15 13 16 13 13 9 13 9 13 2
3 13 1 9
5 9 13 3 13 9
4 0 9 7 9
13 0 9 13 9 7 3 9 9 13 13 9 9 1
17 9 13 3 10 9 15 2 13 9 3 9 2 9 7 9 1 2
25 16 9 13 3 13 3 3 15 13 2 15 13 13 16 9 3 13 9 13 3 3 16 15 13 2
7 13 13 9 13 0 9 2
3 0 12 9
15 9 13 12 9 10 9 1 13 9 2 3 13 0 9 2
5 13 3 3 13 2
7 9 13 3 13 0 13 2
11 15 13 9 7 13 16 9 15 3 13 2
9 9 13 9 15 0 7 9 0 2
6 13 3 7 13 13 2
13 9 9 7 9 9 9 13 3 9 7 9 1 2
11 3 15 13 13 16 3 3 12 9 9 2
4 9 13 3 2
7 11 1 0 15 13 9 2
10 11 13 0 9 7 11 9 0 9 2
7 11 13 13 9 9 9 2
16 9 13 3 15 2 16 9 13 13 13 9 0 9 11 9 2
8 9 13 9 9 7 9 9 2
10 9 13 13 9 1 3 9 9 0 2
2 3 2
4 15 13 13 2
2 0 9
7 9 2 15 0 9 13 9
16 13 0 2 16 9 13 10 9 1 10 9 13 9 13 9 2
4 13 3 9 0
12 15 13 2 16 15 9 10 9 13 15 0 2
6 13 13 15 3 9 2
11 9 12 9 9 13 3 12 0 9 9 2
3 11 15 13
4 15 3 13 15
11 11 13 13 15 3 9 11 3 11 1 2
16 3 3 13 3 15 13 13 3 3 15 16 11 9 7 9 2
13 9 13 13 0 9 3 16 0 9 13 13 9 2
12 13 0 3 9 2 13 9 13 2 13 11 2
17 9 13 9 1 13 3 13 9 7 13 9 13 15 9 7 9 2
2 9 9
10 10 3 9 13 9 13 3 0 9 2
18 3 13 13 9 13 2 16 11 13 13 2 7 16 11 11 13 9 2
2 0 9
7 9 13 7 13 15 9 2
12 15 13 3 3 13 7 3 3 13 0 9 2
13 9 7 10 9 9 13 10 9 3 0 9 0 2
4 15 13 13 3
2 13 13
11 9 2 15 9 13 2 13 13 9 13 2
14 10 9 2 9 11 11 2 13 3 15 9 13 9 2
2 13 13
12 9 13 13 9 2 16 9 9 13 13 3 2
5 9 13 3 0 2
10 9 13 9 11 2 15 13 9 1 2
7 15 13 7 13 1 9 2
5 10 9 13 15 2
14 13 9 7 11 7 11 7 11 7 11 9 13 3 2
8 3 9 13 9 13 9 3 2
7 6 3 0 10 10 9 2
5 13 7 13 13 2
7 15 13 0 9 2 13 2
8 13 0 9 7 9 13 9 2
16 3 9 2 0 3 13 13 9 9 11 2 13 3 12 9 2
18 13 3 10 9 13 9 3 3 2 16 13 10 13 9 13 9 3 2
8 11 11 9 13 9 11 9 2
8 9 9 13 3 9 16 9 2
9 11 1 9 13 13 13 9 1 2
2 10 9
6 13 15 2 9 13 2
9 11 13 13 11 9 3 12 9 2
6 9 13 9 9 1 2
26 12 0 9 2 11 2 11 2 11 7 8 11 2 13 9 9 9 2 7 13 13 9 3 11 1 2
11 16 13 9 3 9 2 9 13 3 13 2
7 15 13 15 3 3 13 2
3 13 9 3
6 9 0 13 9 1 2
11 15 13 9 9 13 7 3 13 3 13 2
3 12 13 9
3 13 9 2
7 11 13 9 1 11 9 2
9 9 13 3 9 1 2 3 9 2
6 3 13 13 10 0 2
11 11 13 3 13 13 15 3 16 13 0 2
2 0 0
8 9 9 13 13 7 13 3 2
7 9 0 9 13 13 9 2
3 15 13 15
4 9 13 9 2
7 13 3 13 13 9 11 2
6 10 9 13 0 13 2
6 15 13 3 9 13 2
3 9 13 13
8 10 11 13 13 10 9 13 2
3 3 0 2
4 13 9 13 2
2 0 9
8 15 13 15 0 9 0 9 2
12 15 13 13 10 9 2 13 15 15 1 13 2
9 13 0 13 15 7 13 3 9 2
10 15 13 3 9 1 13 3 0 9 2
2 0 11
8 0 9 13 3 0 0 9 2
3 15 13 9
7 10 9 11 13 11 9 2
4 6 15 13 2
8 9 12 0 9 12 9 11 11
7 15 15 13 10 0 9 2
11 9 13 3 13 3 3 7 3 16 3 2
7 15 13 3 13 13 9 2
13 9 13 13 3 3 0 9 2 7 15 1 0 0
2 0 9
9 11 9 9 13 13 9 13 9 2
11 3 13 3 12 9 13 16 16 13 3 2
10 3 11 0 9 13 16 10 3 0 9
23 16 9 13 12 9 2 15 3 12 10 9 9 2 3 13 3 9 15 2 3 9 13 2
3 9 9 9
10 13 13 9 10 9 7 9 13 9 2
2 0 9
3 3 13 9
5 15 13 13 9 9
13 11 13 13 15 2 15 13 13 13 0 9 9 2
10 13 13 2 7 3 16 13 3 3 2
6 9 13 7 13 0 2
5 9 13 10 9 2
10 11 13 13 9 1 0 9 13 9 2
9 6 2 3 9 13 3 9 13 2
18 0 7 0 9 13 13 3 9 13 9 1 11 2 11 7 11 9 2
13 13 11 15 13 15 9 7 3 3 13 0 9 2
9 11 13 13 13 11 9 13 9 2
6 13 10 15 13 9 2
7 11 9 3 13 9 9 3
16 9 9 13 3 13 2 16 15 13 10 9 13 9 9 1 2
5 15 13 0 9 2
4 11 13 9 2
12 0 9 13 9 2 15 0 9 13 13 15 2
10 13 15 3 16 15 13 3 10 9 2
6 10 0 13 9 11 2
7 9 13 3 10 9 9 2
14 11 13 13 2 7 13 2 16 9 13 3 0 9 2
4 9 1 13 9
18 9 0 9 13 13 15 2 16 13 9 9 13 15 3 9 7 9 2
16 9 13 3 12 2 15 1 9 13 9 2 9 7 9 9 2
6 15 13 15 13 0 2
9 2 13 9 2 2 13 11 3 2
14 13 9 3 7 13 16 13 3 13 13 10 3 0 2
7 15 13 13 9 9 1 2
6 9 13 3 0 9 2
5 3 15 13 3 2
6 10 9 13 11 13 2
5 3 13 15 3 13
3 3 3 2
13 11 8 7 9 9 0 9 9 13 3 13 9 2
4 13 15 3 2
10 9 2 9 7 0 9 13 9 9 2
13 3 9 9 13 3 2 16 9 13 3 0 9 2
6 15 13 9 11 1 2
4 11 13 13 2
11 15 13 10 9 2 15 1 15 13 9 2
8 0 9 10 10 0 9 13 2
8 7 11 13 2 16 15 13 2
6 9 9 13 9 1 2
9 9 13 13 3 9 13 9 9 2
5 13 13 13 9 2
3 0 9 9
11 15 13 13 3 15 16 13 15 9 9 1
3 10 11 2
8 9 0 9 13 11 9 12 2
6 15 13 9 9 3 2
4 11 7 11 9
3 0 9 2
3 15 13 11
4 9 13 3 2
3 13 13 9
4 13 3 3 2
7 9 13 13 3 12 9 2
9 9 13 9 13 0 0 11 9 2
8 13 3 9 2 3 8 8 2
17 15 13 2 16 9 13 13 9 9 2 7 15 15 3 13 9 2
22 10 9 13 9 1 13 7 15 13 9 13 2 15 1 15 13 13 9 13 9 3 2
9 1 13 9 9 13 13 13 13 2
9 3 13 3 12 9 0 12 9 2
24 13 13 3 3 3 13 10 9 3 3 3 15 13 16 2 15 1 15 3 13 10 9 3 2
4 0 9 9 2
8 7 13 9 11 0 9 13 2
4 13 10 9 2
15 9 13 13 13 2 3 2 9 2 15 13 13 0 0 2
3 2 15 2
5 11 13 11 1 2
11 15 13 9 0 2 16 9 1 13 13 2
18 9 13 11 9 7 0 9 1 3 9 9 2 0 9 9 7 9 2
3 13 15 2
11 13 9 0 9 0 9 0 8 7 9 2
3 0 9 2
6 15 13 0 3 9 2
7 11 7 11 13 9 9 2
4 9 13 16 13
8 10 9 3 3 13 10 11 2
13 11 13 9 2 9 13 9 7 13 13 10 9 2
10 13 15 3 2 16 13 13 9 9 2
10 15 13 13 10 9 3 15 15 13 2
7 15 13 3 9 7 9 2
19 7 15 13 3 3 13 2 16 13 13 3 9 2 15 13 9 3 9 2
6 15 13 3 0 9 2
13 11 13 15 13 3 0 9 2 7 3 15 13 2
8 15 13 3 9 3 0 9 2
4 13 15 3 2
5 15 13 15 9 2
10 9 7 13 13 9 10 9 2 16 2
13 9 13 3 3 0 2 16 3 13 13 3 9 2
9 9 13 2 16 0 9 13 9 2
9 9 13 13 7 9 13 13 0 2
16 0 9 9 2 15 3 13 2 13 9 9 13 13 9 9 2
9 9 13 10 0 9 2 11 13 2
4 9 13 11 2
2 13 13
7 6 3 0 15 13 15 2
3 9 13 13
9 11 9 13 13 3 16 0 9 2
4 2 13 12 2
9 15 13 10 0 9 16 15 13 2
3 15 13 15
8 11 13 13 12 1 9 9 2
9 15 13 15 16 3 13 0 9 2
7 0 9 13 13 0 9 2
14 3 9 13 13 2 16 10 9 13 9 1 13 9 2
13 15 13 3 9 2 16 13 11 0 9 13 11 2
7 9 13 13 12 0 9 2
13 10 9 12 9 13 9 13 12 9 9 13 13 2
2 13 9
7 15 13 3 0 13 9 2
15 6 7 7 3 3 11 3 13 13 13 3 9 1 3 2
14 9 13 0 9 13 9 2 13 15 9 2 15 13 2
3 13 9 2
9 15 13 2 13 15 3 13 2 2
5 9 13 9 3 2
7 9 9 13 1 12 9 2
3 9 13 13
4 13 15 12 13
7 0 9 10 0 1 12 2
4 9 13 3 2
5 3 15 3 13 2
9 15 3 13 13 3 0 9 9 2
6 0 9 13 13 0 2
5 3 3 3 3 2
7 3 9 9 13 9 9 2
15 13 13 13 13 13 9 2 13 9 10 9 9 12 0 2
2 13 15
7 9 13 13 9 12 1 2
7 11 13 13 3 0 9 2
18 11 1 9 13 3 3 12 9 1 2 7 3 15 13 13 9 1 2
10 10 9 0 8 2 8 7 9 16 9
2 9 1
7 11 13 10 9 1 9 2
8 16 9 13 2 15 13 11 2
4 13 10 9 2
6 13 9 9 9 1 2
9 0 9 13 11 9 13 9 9 2
6 9 16 13 10 9 2
15 15 2 16 9 13 2 13 15 2 16 13 13 3 0 2
6 9 9 13 9 12 2
4 9 13 0 3
8 13 13 3 3 2 9 13 2
12 9 13 3 3 3 3 9 7 3 9 3 2
5 11 13 3 9 2
10 11 9 13 0 2 10 9 9 13 2
3 9 13 9
5 3 15 0 13 9
12 9 12 9 13 13 9 13 0 9 9 1 2
13 9 13 15 7 13 0 9 2 16 9 9 13 2
4 15 13 9 2
10 9 13 13 13 9 3 10 12 9 2
17 16 11 3 3 9 9 1 13 15 13 2 9 13 9 3 13 2
19 3 15 0 3 13 9 7 15 0 0 9 9 13 13 3 13 9 1 2
12 13 9 0 3 13 15 13 3 9 1 9 2
7 0 9 13 13 9 9 2
5 13 10 9 0 9
4 13 0 9 2
20 7 3 15 13 3 11 11 0 9 13 9 9 2 15 13 9 13 9 15 2
11 15 3 11 12 13 10 0 7 0 9 2
8 13 15 13 0 16 13 13 2
14 15 13 9 2 15 9 2 0 7 0 13 13 3 2
6 13 9 11 2 16 2
7 12 0 13 7 13 9 9
5 9 13 0 9 2
10 16 13 13 9 13 2 13 0 9 2
4 9 13 0 2
3 9 0 9
5 3 3 15 13 2
7 11 13 2 7 11 13 2
3 13 3 2
4 9 13 9 9
6 13 2 16 9 13 2
5 12 0 9 13 3
6 15 13 3 13 0 2
8 0 9 0 0 9 13 3 2
2 13 9
11 9 13 3 3 3 0 16 9 13 13 2
19 13 3 2 16 10 11 11 11 3 16 13 13 3 2 10 11 11 3 2
10 15 3 3 13 13 2 9 0 9 2
6 13 3 11 1 3 2
12 15 13 9 9 2 13 15 13 13 9 15 2
4 9 13 0 2
39 7 13 13 2 16 10 15 13 13 10 0 9 2 9 3 13 9 2 10 12 9 9 9 2 16 10 1 9 7 9 9 7 9 13 7 9 13 9 2
8 13 9 0 13 9 7 13 2
7 15 13 13 13 15 9 2
21 9 13 12 7 15 9 7 9 9 13 2 3 0 2 9 7 9 13 0 9 2
6 9 13 9 3 13 9
8 11 7 15 13 10 9 0 2
14 9 13 9 2 9 2 9 7 9 7 9 13 13 2
12 3 13 9 2 0 9 2 13 3 9 1 2
8 13 9 9 3 10 9 3 2
4 15 13 11 2
9 15 13 13 0 2 0 9 3 2
10 11 13 13 16 15 13 13 13 3 2
5 13 13 3 0 13
20 15 15 13 13 2 12 9 13 2 16 3 10 15 13 13 10 9 9 9 2
12 10 9 9 13 11 2 11 15 13 13 9 2
10 0 15 3 13 7 15 13 3 0 2
12 9 9 9 13 7 9 9 7 0 9 9 2
8 9 13 13 9 12 7 12 2
10 9 13 13 2 16 10 9 13 9 2
25 11 13 12 9 0 9 2 15 9 0 9 13 9 10 9 13 9 2 16 9 13 13 0 9 2
12 9 13 3 6 2 6 13 9 1 13 9 2
4 15 13 0 2
10 0 9 9 13 13 13 11 13 9 2
10 13 13 3 13 10 9 13 10 9 2
3 13 13 13
10 9 13 9 2 13 9 3 3 3 2
4 9 13 13 3
7 9 13 12 11 0 9 2
7 13 13 9 7 10 9 3
12 13 13 2 16 13 13 3 0 0 9 9 2
2 0 9
4 15 13 13 2
4 2 13 15 2
3 10 0 9
9 13 0 13 0 9 15 2 15 2
6 15 13 3 13 9 2
12 13 9 13 9 2 16 3 13 13 13 9 2
6 9 13 9 12 9 2
7 15 13 10 9 1 13 2
4 13 13 13 13
3 8 7 9
6 9 13 13 13 3 2
13 9 1 9 13 3 9 9 1 2 9 7 9 2
4 15 13 13 2
6 0 0 2 7 3 2
13 9 9 7 9 9 13 9 3 2 15 15 13 2
8 9 13 13 3 3 0 9 2
7 11 13 3 9 13 3 3
8 13 3 9 13 2 11 13 2
16 15 13 3 9 2 16 9 13 13 13 0 2 9 13 9 2
2 0 9
6 11 13 9 9 3 2
6 10 9 13 9 10 9
5 13 0 3 3 2
3 15 13 15
5 15 13 9 3 2
21 15 1 15 13 3 0 9 3 13 13 3 3 10 9 3 3 10 10 9 13 2
10 9 11 13 3 13 9 7 10 9 2
14 9 7 0 9 13 9 9 0 9 1 13 12 9 2
11 13 13 2 16 9 13 3 2 15 13 2
7 9 0 9 11 13 13 2
5 13 15 3 13 2
14 3 13 13 9 2 16 9 0 10 9 9 13 13 2
6 9 15 13 1 9 2
16 0 9 9 13 13 2 3 0 9 3 13 3 0 9 9 2
2 13 9
6 15 13 3 12 1 2
7 15 13 13 10 3 13 2
15 3 3 9 13 13 0 9 3 2 16 15 13 3 13 2
13 9 11 11 13 3 13 9 9 3 3 9 1 2
4 9 13 9 1
7 9 9 13 11 1 11 2
8 7 11 1 13 9 9 9 2
7 9 9 11 13 9 9 2
7 9 13 0 2 15 13 2
2 16 3
3 0 9 3
9 10 9 13 3 13 3 0 9 2
19 9 13 3 2 15 13 15 2 16 10 12 9 9 13 13 7 9 13 2
11 11 1 2 11 13 15 10 0 9 2 2
9 9 13 13 13 9 7 9 1 2
10 3 9 13 3 2 16 15 13 3 2
5 9 13 7 9 2
6 9 13 15 13 13 2
11 3 15 13 13 13 9 9 2 9 9 2
6 11 13 9 3 3 2
9 15 13 3 9 0 0 9 1 2
19 9 9 13 3 3 3 0 9 9 1 2 13 15 12 9 9 2 13 2
4 9 13 9 9
26 13 13 9 9 2 7 15 3 13 15 13 2 2 13 13 2 15 13 11 2 13 11 2 9 13 2
6 15 13 9 9 12 2
11 16 13 9 13 2 9 13 3 0 9 2
2 3 9
11 9 13 9 15 13 15 0 9 13 9 2
6 15 3 13 0 9 2
19 11 13 0 2 0 9 2 7 9 15 13 9 9 13 3 9 13 9 2
5 9 13 9 9 2
21 3 12 9 1 9 13 9 7 9 10 9 12 9 0 11 1 9 7 3 11 2
15 15 3 9 9 13 3 13 9 3 16 0 9 9 1 2
8 12 9 1 13 13 12 9 2
5 13 3 3 9 2
8 11 13 3 0 9 9 9 2
10 11 13 3 9 0 7 9 7 9 2
11 9 11 13 12 3 3 0 9 2 9 2
2 9 1
2 10 9
2 10 0
3 13 9 1
2 0 9
11 9 13 15 2 16 9 13 3 0 9 2
9 15 13 9 2 15 3 9 12 2
2 0 9
5 13 9 0 9 2
12 13 13 11 3 7 3 3 13 7 13 9 2
5 3 13 15 9 2
5 3 9 13 9 2
2 3 13
12 7 13 13 13 9 3 2 16 15 13 15 2
9 10 9 13 3 3 12 9 9 2
9 9 11 13 13 0 12 9 9 2
16 9 11 11 13 13 12 7 13 13 9 11 10 9 0 9 2
8 13 9 9 13 7 13 13 2
6 13 13 11 9 9 2
8 3 9 13 13 9 9 9 2
26 13 3 15 3 15 16 3 9 7 15 13 13 16 7 10 9 3 16 9 9 3 13 15 10 9 2
11 0 9 7 3 0 9 2 15 9 13 2
10 0 3 11 13 9 9 9 9 1 2
6 15 9 13 3 3 2
5 15 3 3 13 2
2 9 9
6 15 13 3 15 3 2
17 3 16 15 13 15 13 2 15 13 13 9 9 7 13 9 9 2
3 13 9 2
16 9 0 9 2 3 9 2 9 7 9 2 9 13 3 13 2
7 9 13 9 1 13 3 2
2 9 9
6 9 15 13 15 3 2
5 2 13 15 3 2
8 0 9 13 3 13 9 0 2
3 13 9 1
5 9 1 13 9 2
6 13 3 13 15 3 2
4 9 13 12 2
8 9 13 3 0 2 7 0 2
6 9 13 3 15 0 2
11 11 13 9 0 9 2 0 13 0 9 2
20 12 13 11 3 13 9 2 16 15 1 12 13 11 13 9 9 1 12 9 2
5 9 9 0 9 9
5 9 13 3 0 2
12 9 7 9 13 13 10 9 2 3 13 9 2
5 11 13 13 0 2
6 11 13 3 10 0 2
2 9 13
5 9 13 9 1 2
20 16 9 13 13 2 7 13 13 3 13 13 9 2 0 9 13 9 13 9 2
13 13 3 13 11 9 11 9 9 2 16 9 13 2
9 13 13 2 13 15 3 0 9 2
7 10 0 9 9 13 0 2
7 9 11 9 13 0 9 2
9 15 13 13 3 9 0 9 9 2
17 9 13 13 0 0 9 2 16 11 13 9 13 0 7 0 9 2
3 9 13 3
7 3 3 13 13 9 9 2
19 13 9 2 9 2 9 2 13 9 2 0 9 7 3 3 10 3 0 2
3 13 9 2
4 13 15 3 2
10 9 13 11 7 10 9 9 3 9 2
3 9 9 9
6 15 15 13 0 9 2
3 13 9 9
22 13 15 9 2 15 13 13 3 3 13 15 7 15 2 3 16 15 3 13 15 7 2
11 11 13 11 0 9 2 15 13 3 9 2
4 0 13 0 9
14 11 13 0 13 10 0 9 2 15 13 13 11 3 2
5 15 13 9 9 9
10 9 13 9 13 9 13 9 3 3 2
7 9 13 9 9 10 9 2
10 9 13 9 7 9 9 2 3 3 2
4 9 3 9 9
7 15 13 13 3 2 7 2
11 7 13 0 13 3 13 10 9 7 9 2
16 13 3 16 13 11 13 13 3 16 13 15 13 13 0 9 2
13 9 11 9 13 2 16 15 13 3 9 13 9 2
4 13 12 9 2
2 0 9
4 15 13 13 9
4 9 13 9 1
38 15 13 3 3 0 3 10 9 16 15 13 3 0 0 7 0 7 0 3 15 3 13 7 15 3 3 15 13 0 9 16 3 15 13 3 3 7 2
11 6 3 0 9 3 15 13 12 0 0 9
7 3 3 15 3 13 13 2
3 11 9 3
2 0 9
8 15 13 9 3 0 9 9 2
5 15 10 0 13 2
4 7 13 11 2
17 0 9 3 13 7 9 13 13 3 11 2 0 9 7 0 11 2
6 13 3 12 9 10 9
8 9 2 15 9 13 0 13 0
9 2 13 13 0 2 2 11 13 2
4 9 13 12 9
13 10 9 13 13 9 2 16 3 9 13 13 9 2
8 9 13 2 16 15 13 3 2
17 15 13 15 0 0 7 15 1 13 9 3 3 7 10 9 7 2
6 3 13 9 10 9 2
5 15 15 13 3 13
5 9 13 3 1 2
8 7 13 15 13 10 9 0 2
2 10 9
7 13 3 2 3 13 9 2
5 13 15 13 8 2
4 13 9 9 2
12 1 9 9 13 9 7 3 13 13 13 9 2
5 9 13 15 9 2
23 16 9 15 13 3 3 13 7 3 3 15 13 15 3 2 15 13 3 10 9 2 13 2
2 0 9
2 9 9
8 9 7 9 1 0 13 15 2
8 8 7 9 13 1 10 9 2
4 0 7 0 9
8 10 9 13 0 16 10 9 2
12 11 9 13 10 0 0 11 2 6 2 11 2
15 15 13 13 13 0 11 9 2 13 15 13 3 0 0 2
8 9 13 13 13 16 12 9 2
6 3 13 9 13 0 2
7 11 1 15 13 13 9 2
18 3 3 13 2 3 15 13 13 3 2 3 16 15 13 3 13 15 2
8 13 0 2 13 13 7 13 2
4 13 11 9 2
4 3 13 9 2
6 13 11 9 0 9 2
9 13 0 2 16 11 13 13 0 2
14 3 15 13 3 9 1 12 9 7 13 2 16 13 2
4 15 13 13 3
20 15 13 3 0 9 7 13 9 16 9 9 2 9 0 9 2 9 9 9 2
8 16 13 2 15 13 15 3 2
10 13 13 3 15 2 7 0 0 1 2
4 13 9 7 9
2 13 2
3 13 3 9
2 9 9
11 0 9 13 0 13 13 9 15 16 9 2
6 9 13 9 13 3 2
4 15 13 0 9
2 13 13
9 9 9 11 11 13 9 13 9 2
10 0 9 9 2 9 7 9 9 13 2
12 9 7 9 9 13 13 3 13 0 9 9 2
16 13 3 3 13 13 2 16 10 9 2 13 3 10 0 9 2
6 13 9 9 7 9 2
10 9 2 15 9 13 15 0 7 0 13
14 15 13 3 0 9 2 16 9 3 13 2 9 13 2
2 0 9
8 9 13 9 13 3 12 1 2
5 13 9 7 3 2
15 11 9 13 0 2 0 9 2 0 9 13 15 3 3 2
6 9 0 9 13 9 2
3 3 15 2
18 0 9 13 13 3 9 2 3 2 7 3 15 13 13 13 0 1 2
5 15 13 9 1 2
11 9 15 13 9 9 2 3 3 2 13 2
8 13 15 2 3 15 13 9 2
6 13 3 0 9 9 2
16 13 3 3 0 15 1 7 13 15 13 9 7 13 0 9 2
16 9 13 0 9 3 3 2 16 13 9 13 9 0 9 9 2
4 9 2 9 2
7 15 13 9 13 10 9 2
5 9 13 9 1 9
11 11 13 11 9 13 13 12 9 13 3 2
6 9 13 10 9 3 2
6 15 13 0 9 0 9
6 13 9 3 7 13 2
7 0 1 9 13 3 13 2
7 9 13 9 9 3 11 2
2 13 9
10 15 13 3 16 13 13 9 9 10 9
8 7 11 13 0 7 13 11 2
12 9 13 11 9 2 15 13 15 1 13 13 9
3 9 13 11
10 0 2 9 0 7 9 3 10 9 2
7 12 0 9 15 15 13 2
3 13 3 2
8 11 13 9 3 3 13 9 2
6 10 12 13 3 9 2
3 13 15 1
5 11 2 11 13 9
5 9 13 3 13 2
2 0 9
11 9 9 13 7 13 9 7 15 13 9 2
5 2 13 15 9 2
14 13 15 10 9 13 10 0 9 7 13 15 3 3 2
4 15 13 9 2
2 0 9
16 15 13 3 3 13 11 9 2 3 3 0 9 15 13 13 2
10 3 15 13 3 13 9 7 0 9 2
6 10 9 13 3 0 2
12 9 0 9 13 15 1 2 3 9 13 9 2
15 9 9 13 2 16 9 13 0 9 9 7 0 12 9 2
19 16 11 13 9 9 2 16 15 13 13 15 3 2 13 15 3 3 13 2
6 3 13 0 13 11 2
12 15 13 0 3 2 16 9 13 9 13 9 2
4 15 13 9 2
7 10 9 13 15 1 13 2
3 11 9 9
8 13 9 11 3 11 13 16 2
5 9 1 13 9 2
13 9 13 3 13 2 16 13 13 2 16 13 13 9
8 13 3 2 16 9 13 3 2
13 11 9 13 9 2 16 13 11 3 10 9 13 2
6 9 13 3 0 9 2
6 3 15 13 2 9 2
16 9 13 9 2 13 0 2 9 13 13 9 1 7 13 3 2
18 15 7 9 13 15 1 3 3 3 9 2 13 9 9 11 2 12 2
5 9 13 0 9 2
4 16 13 3 13
7 13 0 16 13 12 9 2
8 9 9 13 13 3 9 9 2
13 11 13 9 2 13 13 3 9 2 15 15 13 2
11 7 16 0 13 11 7 0 2 13 9 2
8 9 13 9 2 13 3 13 2
5 13 9 0 9 2
5 9 13 15 9 9
3 9 13 9
8 3 0 9 13 13 0 9 2
9 9 13 3 16 16 15 0 13 2
10 6 3 9 15 13 16 10 9 13 2
20 15 13 3 0 9 13 15 15 13 12 12 9 16 15 3 13 15 1 3 2
9 6 13 15 2 11 2 15 13 2
13 9 9 9 13 9 2 9 9 0 9 13 3 2
5 9 13 0 9 2
6 11 13 9 9 13 2
4 15 13 11 2
5 3 15 13 9 2
17 9 13 13 0 9 2 15 13 13 0 9 7 0 9 9 1 2
12 9 13 3 13 9 7 9 15 16 3 9 2
5 10 9 15 13 2
5 15 13 13 9 2
6 11 13 3 0 9 2
3 13 9 2
12 9 7 3 13 3 11 9 1 0 9 13 13
4 9 13 12 9
10 13 10 9 3 6 10 9 9 13 2
10 9 13 11 2 3 13 9 1 11 2
7 9 13 9 10 9 0 9
10 2 13 9 7 3 0 9 13 2 2
4 9 13 1 9
11 13 13 3 3 2 16 15 13 15 0 2
15 11 13 13 2 7 13 0 9 3 7 13 3 3 9 2
9 10 0 0 1 13 0 9 0 2
13 9 9 13 13 13 10 9 9 0 9 10 9 2
6 12 12 9 13 9 2
6 0 9 13 13 3 3
2 9 9
9 3 9 9 13 10 9 13 3 2
9 3 0 7 0 10 9 3 13 2
5 3 15 13 9 2
13 15 13 0 7 0 2 3 9 9 13 13 9 2
4 9 9 9 9
7 9 13 3 9 0 9 9
9 11 13 0 13 7 13 9 9 2
6 6 13 3 10 9 2
9 0 9 9 13 9 0 0 9 2
5 15 13 0 9 2
8 3 11 7 11 7 11 9 2
3 8 7 9
3 0 9 9
5 3 13 10 9 2
9 11 1 9 9 13 3 9 11 2
14 11 13 11 13 10 9 9 2 16 13 9 1 13 2
5 11 13 3 0 2
12 13 0 13 2 16 0 9 13 7 0 7 0
16 11 13 13 9 2 13 3 10 9 2 15 13 9 0 9 2
3 3 13 9
11 10 9 2 16 13 15 2 9 13 9 2
16 15 13 15 1 16 13 9 1 15 13 15 1 9 7 9 2
7 9 13 0 16 0 9 2
5 15 13 0 9 2
8 0 9 15 13 3 13 9 2
2 12 12
6 15 13 13 13 9 2
12 3 0 3 0 9 13 9 9 2 13 9 2
3 9 13 13
7 10 9 15 13 3 3 9
9 6 2 15 13 3 3 3 9 2
3 13 13 2
4 13 3 9 2
8 9 9 13 9 0 7 9 2
8 15 13 0 9 3 10 12 9
5 9 13 3 10 9
11 13 10 9 15 13 9 0 0 0 9 2
8 16 3 13 3 3 10 9 2
20 6 3 6 3 12 9 16 15 13 3 15 1 13 0 9 15 13 12 9 2
5 13 10 9 3 2
17 15 1 16 9 13 13 9 2 9 9 11 9 13 13 12 9 2
2 0 9
7 0 9 9 13 13 3 2
10 9 1 13 0 9 2 13 11 11 2
13 13 15 10 0 9 9 7 3 2 15 13 13 2
3 9 9 2
8 15 13 3 2 9 7 9 2
10 9 13 9 12 9 13 3 12 0 2
12 3 16 15 13 3 13 2 16 11 13 13 2
7 13 9 15 0 11 9 2
6 10 9 15 3 13 2
3 13 9 3
8 16 15 13 9 1 7 9 2
4 0 9 15 2
6 9 13 3 13 3 2
4 9 13 9 9
10 2 15 13 0 2 2 11 11 13 2
9 13 9 13 13 9 1 9 1 2
2 9 9
7 10 9 9 9 13 13 2
4 13 3 9 2
10 15 13 3 2 3 15 13 12 3 2
10 13 15 3 2 16 3 13 9 9 2
14 9 13 7 13 13 3 15 13 2 15 13 7 3 2
7 9 15 13 0 9 1 2
12 3 10 9 3 9 13 13 12 9 13 9 2
16 3 16 15 13 13 3 3 9 2 15 13 3 3 13 3 2
4 13 15 9 2
12 11 13 7 13 9 9 2 3 15 13 13 2
6 9 13 9 11 9 2
3 9 13 13
17 13 15 13 13 3 12 9 0 2 13 9 11 9 9 11 9 2
4 9 13 3 2
4 10 9 13 2
8 16 15 13 13 0 0 9 2
10 11 13 0 9 13 0 9 9 0 2
11 10 9 1 11 13 13 13 2 16 13 9
4 3 13 15 2
5 15 13 13 15 2
6 9 13 3 12 1 2
19 15 13 3 0 2 7 13 3 2 16 13 9 13 9 2 13 15 13 2
20 11 13 15 9 2 13 2 13 11 7 13 2 13 2 16 15 13 9 9 2
4 11 13 13 13
4 15 13 15 2
14 13 9 13 9 9 7 9 9 13 12 0 9 9 2
7 13 15 13 10 0 9 2
10 13 2 13 15 13 10 10 9 9 2
4 9 11 9 13
11 3 13 16 11 7 11 9 13 15 1 2
5 11 3 9 13 2
8 6 6 16 15 13 13 3 2
13 9 9 13 9 13 3 3 9 7 0 9 1 2
8 11 13 13 15 10 0 9 2
3 9 0 9
3 13 3 2
12 11 13 9 9 2 13 11 7 13 0 9 2
20 3 3 13 9 9 13 0 15 1 2 16 15 13 13 9 7 3 13 15 2
8 10 9 2 15 3 3 3 13
17 15 13 3 3 0 9 16 16 16 15 13 3 12 9 9 10 9
14 3 9 0 9 13 11 3 3 7 13 3 0 9 2
12 9 12 15 13 0 9 11 7 9 13 9 3
6 10 15 15 13 9 2
8 9 13 0 9 13 11 9 2
10 0 13 13 3 0 3 13 9 3 2
8 15 13 9 2 13 13 15 2
4 15 13 9 9
9 3 13 13 9 2 13 13 3 2
8 0 9 9 0 9 13 3 2
4 13 3 9 2
6 3 9 13 3 3 2
8 0 1 9 13 11 13 9 2
9 11 13 11 11 13 9 0 9 2
8 13 12 9 10 12 9 9 2
5 16 15 13 0 9
13 15 13 10 9 7 13 15 2 0 16 13 13 2
14 0 1 3 13 13 0 9 2 15 3 13 15 9 2
17 3 9 13 3 3 0 2 9 2 13 9 0 9 16 12 9 2
6 9 13 3 0 9 2
3 13 9 2
5 9 11 13 0 2
6 15 13 13 9 13 2
15 3 9 13 3 3 3 16 3 2 3 9 13 13 3 2
12 11 7 11 13 9 9 10 9 7 0 9 2
8 13 13 13 11 13 9 9 2
7 12 9 9 13 9 3 9
14 9 13 15 2 16 15 12 9 9 13 9 0 9 2
6 0 13 3 13 3 2
14 0 13 2 16 13 11 9 13 3 0 9 16 11 2
9 3 15 3 3 13 16 0 9 2
8 15 13 3 13 13 13 9 2
5 3 10 9 13 2
8 9 13 7 9 13 9 1 2
5 3 9 11 3 2
11 3 3 13 9 0 9 2 10 9 1 2
7 13 15 3 13 9 16 9
3 13 15 13
8 11 13 3 9 2 11 13 2
57 13 9 9 13 9 15 13 3 15 13 9 13 2 3 16 15 13 3 3 9 13 3 7 13 9 10 9 3 16 15 13 13 15 13 2 7 16 15 13 9 10 9 9 9 13 3 9 9 2 13 15 13 15 13 9 15 2
7 13 2 16 13 10 0 2
2 13 9
8 7 13 0 16 13 9 13 2
5 13 15 13 9 2
8 13 0 7 0 0 9 9 2
8 15 13 3 0 0 9 1 2
4 0 9 15 2
13 2 11 1 15 13 3 12 9 2 2 15 13 2
3 9 7 9
25 15 13 9 3 2 15 16 13 0 9 3 3 2 15 13 12 9 13 3 15 13 10 9 13 2
20 7 15 13 3 3 9 0 8 9 15 16 3 13 16 13 3 0 13 9 2
3 13 9 1
8 13 16 13 9 15 13 3 2
4 13 3 0 2
10 9 13 9 7 13 16 13 15 13 2
2 0 9
6 9 13 9 13 9 2
8 13 16 13 13 3 13 15 2
7 7 9 13 9 9 12 2
10 15 15 13 0 9 7 9 13 13 3
13 0 13 3 9 2 15 12 9 0 9 13 3 2
11 9 13 13 9 2 15 9 13 13 3 2
4 13 9 15 2
14 9 13 3 15 15 13 2 13 13 15 10 9 13 2
9 3 9 9 13 13 9 7 9 2
4 0 13 13 2
8 9 13 3 0 0 13 9 2
7 0 13 9 2 0 12 2
6 9 13 9 7 3 0
6 15 15 13 3 13 2
8 15 13 3 13 13 10 9 2
3 10 10 9
10 2 13 13 10 9 3 7 3 2 2
2 13 15
7 0 9 13 9 0 9 2
5 0 9 13 10 9
2 13 3
2 9 9
9 13 2 16 13 15 3 3 13 2
7 13 9 3 3 13 13 2
3 9 3 11
5 15 3 13 15 2
20 15 13 13 15 10 9 2 16 13 9 7 0 2 7 16 13 0 9 1 2
7 0 9 13 9 3 9 2
7 3 0 13 9 0 9 2
16 11 9 13 0 2 0 2 0 7 0 16 10 9 10 9 2
5 9 13 12 12 2
9 15 13 2 15 16 13 13 15 3
10 9 13 9 3 1 9 13 13 13 2
6 15 13 9 7 13 3
6 3 3 0 9 13 2
3 15 13 0
18 3 9 9 13 13 9 2 15 10 9 13 0 2 15 15 13 9 2
11 9 1 15 13 3 7 13 0 9 9 2
4 11 13 9 2
7 3 15 13 3 13 13 2
8 15 13 15 1 13 3 9 13
12 11 13 15 13 3 9 7 9 9 2 16 2
16 3 13 9 13 15 2 15 15 10 9 13 13 3 0 9 2
13 7 16 11 13 2 13 9 11 2 9 9 9 2
13 9 13 13 9 10 9 2 10 9 7 10 9 2
2 13 9
7 3 9 13 9 7 9 2
3 13 13 13
7 11 9 13 9 11 0 2
8 11 7 11 13 9 11 1 2
3 9 9 11
16 9 13 9 15 2 16 13 9 13 9 9 2 13 1 9 2
12 9 13 9 0 9 7 13 15 13 9 9 2
6 9 9 9 13 3 2
17 0 11 13 3 3 0 2 0 9 13 2 16 3 13 9 2 2
9 11 13 9 2 16 13 13 9 2
3 13 9 3
14 15 15 13 2 16 15 13 15 2 10 9 15 13 2
15 9 3 13 15 13 9 9 2 3 3 3 3 13 13 2
3 15 13 13
8 9 13 9 13 9 9 9 2
6 9 13 13 13 9 2
12 3 9 13 3 3 16 10 15 13 3 13 2
15 11 13 13 3 10 9 2 15 11 13 15 3 9 12 2
2 9 9
15 9 13 3 9 1 13 9 3 13 9 9 7 9 13 2
4 13 15 15 2
6 15 13 9 0 11 2
6 9 13 9 10 9 2
11 9 13 13 10 3 9 16 9 7 9 2
11 3 15 13 3 2 16 13 13 15 0 2
12 9 2 9 2 9 7 9 13 3 2 3 2
6 9 13 0 9 1 2
7 0 9 9 13 3 11 2
16 15 15 2 0 12 0 9 3 13 9 2 13 13 3 15 2
20 9 13 13 9 1 12 12 9 1 2 16 9 13 7 13 9 9 13 9 2
7 11 13 13 9 3 9 2
10 13 3 0 2 16 13 15 13 9 2
2 0 9
8 2 3 13 2 2 11 13 2
12 10 3 9 13 3 10 16 0 0 9 9 2
5 13 13 9 1 2
6 9 13 9 3 0 2
8 13 10 9 3 15 3 13 2
11 15 2 15 13 3 13 9 0 2 15 2
10 9 13 9 2 15 3 13 9 9 9
21 9 13 3 3 0 2 7 15 13 9 2 6 2 15 13 13 3 3 9 2 2
7 10 9 9 13 9 9 2
9 9 13 9 9 2 15 15 13 2
13 3 9 3 13 3 2 13 7 13 10 9 9 2
12 9 13 9 11 11 2 9 2 13 3 9 2
15 8 8 13 7 13 16 13 9 9 9 3 9 9 1 2
11 15 13 0 7 9 7 0 9 1 0 2
2 9 13
6 13 0 9 7 0 2
4 13 9 1 9
6 10 9 9 13 13 2
6 10 9 13 0 9 2
6 3 9 2 13 15 2
4 3 15 9 2
12 15 13 9 3 13 9 2 7 15 13 13 2
17 15 2 16 9 13 13 3 9 7 10 9 2 15 13 13 0 2
5 0 9 13 3 2
3 15 13 0
7 15 13 9 3 9 9 2
8 15 3 13 2 16 13 13 2
3 13 13 13
11 1 11 9 9 0 9 13 3 9 9 2
10 9 7 9 13 13 13 3 9 1 2
9 9 9 13 3 11 9 9 1 2
5 9 13 3 9 2
8 7 15 13 13 9 13 13 2
4 10 9 13 9
8 9 1 11 13 13 12 9 2
10 3 15 3 13 13 2 16 13 11 2
5 13 3 10 9 3
7 3 3 13 9 2 3 2
3 15 13 2
5 9 15 13 12 2
10 0 13 9 9 1 13 12 9 1 2
3 9 0 9
4 10 9 13 9
2 9 9
6 9 0 9 13 9 2
4 9 13 9 2
14 11 13 13 9 15 9 3 13 9 7 0 9 9 2
12 11 13 0 11 13 11 9 10 9 0 9 2
4 0 11 7 11
8 13 13 3 13 3 10 9 2
6 15 13 11 11 3 2
6 11 13 13 9 3 2
6 9 13 3 3 3 2
9 15 13 11 9 2 15 13 15 2
10 9 13 0 9 7 3 3 9 3 9
4 15 13 9 2
6 13 2 16 15 13 2
4 9 13 9 9
12 12 9 1 3 13 7 9 13 0 9 3 2
3 13 9 2
6 9 1 13 9 9 2
8 9 7 9 13 12 0 9 2
2 3 2
3 13 13 9
6 3 13 15 11 9 2
16 16 13 13 13 9 9 2 13 13 3 3 3 2 11 13 2
10 9 13 2 16 9 13 3 3 13 2
5 9 13 9 13 2
9 13 3 13 10 9 3 13 13 2
4 15 13 13 3
2 3 3
3 11 9 11
12 9 13 13 9 9 2 3 15 13 0 9 2
12 9 0 9 13 15 2 16 9 9 13 13 2
16 3 9 13 3 13 0 9 3 2 16 13 16 13 9 11 2
11 15 2 15 13 13 13 15 3 2 13 2
6 15 9 13 13 13 2
10 9 13 9 12 9 3 16 0 9 2
4 12 9 13 9
21 3 13 16 13 13 10 9 7 3 13 13 16 13 3 13 15 13 13 10 9 2
14 9 9 13 3 0 2 16 13 9 13 13 9 13 2
3 13 9 1
5 1 9 13 3 2
9 13 3 3 9 13 9 9 9 2
5 15 13 9 12 9
9 10 0 9 13 9 7 9 0 2
4 6 16 0 2
18 9 3 15 9 13 3 12 7 12 9 2 9 9 2 3 3 12 2
6 15 13 10 10 9 2
12 3 13 3 3 0 9 2 16 13 13 13 2
14 15 13 13 3 3 2 13 13 3 2 3 9 13 2
17 13 3 3 9 13 3 6 6 9 2 9 9 2 10 9 13 2
8 9 13 3 7 3 2 9 1
6 13 9 3 16 15 2
3 13 13 9
7 15 13 13 16 11 12 2
11 9 1 0 9 13 13 9 0 9 13 2
6 15 13 0 13 9 2
13 3 9 13 9 2 10 9 7 9 0 9 9 2
20 3 10 10 9 13 3 3 3 2 3 13 3 0 13 10 9 9 10 9 2
4 13 13 9 2
3 13 15 15
10 10 9 13 9 13 0 9 3 9 2
6 0 9 13 0 9 2
6 13 13 9 7 9 2
21 9 0 9 1 13 9 13 7 3 13 16 15 13 15 2 13 15 13 7 9 2
6 3 15 15 3 13 2
9 9 13 2 13 0 9 13 9 2
7 3 9 13 13 9 1 2
12 15 13 13 9 10 3 3 9 16 10 0 2
5 11 11 12 13 9
4 9 13 0 2
6 15 13 13 9 1 2
6 9 13 10 9 9 2
9 15 13 2 16 9 13 0 9 9
6 9 13 0 9 13 2
3 13 10 9
3 10 11 9
3 11 13 9
8 15 13 12 13 11 9 1 2
3 13 13 9
10 13 0 9 9 2 15 1 15 13 2
16 9 13 3 13 0 9 2 3 9 2 15 13 15 16 9 2
12 9 9 13 11 1 0 10 9 9 13 13 2
12 10 11 9 13 2 16 12 13 11 9 9 2
7 9 9 13 3 3 11 9
7 13 13 3 0 9 13 2
9 9 2 15 13 9 7 3 3 2
8 11 13 13 3 10 9 9 2
7 10 9 13 9 13 9 2
6 15 13 3 3 9 2
7 9 13 13 13 11 9 2
40 13 15 13 13 15 16 15 13 12 9 9 16 15 13 10 0 9 13 13 16 3 3 15 13 15 7 3 7 3 13 3 11 7 10 11 7 11 13 16 2
4 15 13 3 2
2 3 3
11 9 0 0 9 13 2 13 11 3 9 2
2 13 13
9 9 9 9 13 13 3 12 9 2
10 13 0 2 16 9 13 9 0 9 2
3 15 13 3
7 13 9 9 9 9 9 2
2 13 9
8 3 12 9 13 3 3 3 2
12 15 2 15 13 3 15 2 13 13 3 9 2
16 16 0 9 13 13 3 2 13 13 2 16 13 9 9 13 2
4 15 13 11 2
5 0 0 9 13 9
3 13 9 2
7 9 13 3 12 0 9 2
5 3 0 13 9 2
5 13 9 13 9 2
6 9 9 13 0 9 2
7 11 7 11 13 11 9 2
6 13 3 10 9 3 2
12 9 9 13 3 2 16 13 9 1 13 13 2
8 9 0 9 1 13 3 13 2
7 13 0 9 0 9 9 2
9 9 13 9 9 13 9 0 9 2
9 9 13 9 13 12 2 7 12 2
5 15 13 13 3 2
4 7 6 13 2
7 9 13 13 7 9 13 2
16 9 13 9 2 15 13 9 2 16 0 9 13 9 7 9 2
5 9 13 3 13 13
6 13 13 9 13 9 2
6 0 9 0 7 0 9
4 13 3 0 9
5 9 13 0 9 2
15 0 9 13 13 3 2 13 2 13 9 7 13 3 9 2
4 9 13 9 2
16 9 13 9 7 9 9 2 7 9 13 11 1 10 9 13 2
12 11 13 0 9 12 0 9 2 11 7 11 2
15 12 9 9 9 13 11 2 15 3 13 9 11 10 9 2
6 9 9 13 3 3 2
7 9 13 0 2 11 13 2
5 9 13 0 9 2
3 13 13 9
4 9 13 3 2
5 9 13 9 13 9
6 11 13 9 9 9 2
7 15 16 13 2 13 9 2
12 9 13 13 3 10 13 2 15 13 3 13 2
9 11 13 0 9 13 9 13 9 2
22 7 16 0 9 13 13 3 3 9 7 9 16 15 1 2 3 3 15 13 0 3 2
13 3 16 13 13 9 7 9 2 13 3 3 11 13
13 9 13 3 9 1 9 12 7 12 9 9 1 2
12 11 0 7 9 13 9 13 13 0 3 11 2
6 9 9 16 13 13 2
3 9 13 2
6 9 1 9 13 0 2
6 9 13 9 13 9 2
8 13 0 2 16 9 13 9 2
3 9 11 1
13 13 3 9 9 7 15 9 7 3 9 13 3 2
19 13 3 2 16 0 9 13 9 9 2 16 0 2 0 9 15 3 13 2
11 9 13 13 10 9 0 9 1 0 9 2
9 13 13 9 1 2 7 3 3 2
20 11 9 2 9 2 0 9 7 0 9 0 9 13 3 2 15 13 13 3 2
7 13 3 3 0 0 9 2
2 13 13
6 13 3 9 1 3 2
9 13 13 3 3 0 9 16 3 2
12 0 9 3 13 15 2 13 9 3 13 9 2
3 12 0 9
8 9 12 13 13 9 0 9 2
34 15 13 0 9 3 6 3 9 10 9 7 15 15 3 13 15 9 13 13 3 0 3 15 13 9 7 13 3 15 9 9 13 11 2
4 9 1 9 9
12 13 3 0 2 13 15 13 3 15 15 13 2
7 11 13 12 11 12 9 2
3 9 9 9
10 3 9 13 0 13 15 7 10 0 2
2 3 3
9 9 13 13 9 12 9 12 1 2
8 15 13 13 3 3 15 3 15
9 13 0 2 16 15 13 3 3 2
23 15 13 9 2 9 2 9 2 9 2 9 7 9 0 9 2 15 13 3 0 9 9 2
11 10 9 3 13 9 2 3 3 13 15 2
7 9 13 13 3 12 9 2
4 9 13 9 1
10 9 9 13 9 7 9 3 13 15 2
8 15 13 15 0 9 3 9 2
9 9 13 13 9 9 13 3 13 2
10 13 9 0 9 2 13 9 0 11 2
5 9 13 11 13 2
5 15 3 13 9 2
11 11 13 3 0 2 12 9 13 9 9 2
10 13 13 13 9 3 16 15 13 9 2
15 0 9 13 3 2 16 10 9 13 3 7 16 15 13 13
5 13 13 12 0 2
5 9 13 9 13 2
9 16 15 13 15 2 11 13 11 2
6 15 13 13 13 9 2
8 9 2 9 7 9 13 13 2
10 10 9 9 9 13 3 3 12 9 2
10 13 15 13 9 9 10 15 0 9 2
4 9 13 9 2
8 3 2 6 7 13 13 3 2
4 3 13 0 9
7 9 13 3 0 0 9 2
4 15 13 0 2
6 9 13 3 0 13 2
9 16 9 13 15 2 13 9 13 2
7 9 9 13 0 13 9 2
6 9 13 13 0 9 2
9 9 13 13 3 16 0 9 1 13
3 9 1 9
16 12 0 9 13 11 9 11 2 15 1 13 13 9 13 0 2
9 3 13 0 9 16 3 0 9 2
3 10 9 2
11 9 9 13 13 3 0 2 7 15 3 2
10 9 9 7 9 13 9 10 9 9 2
5 13 15 3 13 2
9 15 13 10 0 16 13 13 9 2
14 3 15 13 3 9 15 7 13 9 9 7 9 9 2
5 9 13 3 0 2
8 15 13 13 3 3 10 9 2
5 0 9 9 13 2
9 11 9 13 3 12 9 7 9 2
6 9 1 9 11 13 9
6 9 1 15 13 0 9
4 15 13 3 2
16 9 11 3 11 11 9 13 13 9 2 16 9 13 3 13 2
8 13 15 13 9 13 10 9 2
6 15 13 13 2 13 3
7 0 9 2 13 16 13 2
13 10 15 13 0 9 2 16 9 13 9 0 9 2
3 9 9 11
2 3 0
15 15 13 15 9 3 7 13 3 13 9 9 7 13 9 2
5 15 13 15 0 2
8 13 13 10 9 7 13 11 2
6 15 13 0 9 9 2
13 13 13 3 15 16 13 15 9 6 2 9 1 7
18 13 13 2 16 0 13 2 13 13 15 13 13 9 2 16 9 13 2
2 9 13
5 2 13 10 0 2
9 11 11 13 9 9 1 0 0 2
11 16 10 9 13 15 0 2 13 9 9 2
5 3 3 3 13 2
6 10 9 13 10 9 2
9 13 2 16 13 13 13 9 3 2
5 9 13 13 9 2
6 11 13 3 3 9 2
27 3 15 3 13 13 3 0 9 3 3 0 9 16 15 11 3 13 16 3 9 13 3 13 3 12 9 2
22 13 9 3 0 16 15 7 13 3 13 2 16 3 13 3 13 7 3 13 3 13 2
9 15 13 3 13 15 0 0 9 2
14 2 11 0 13 9 13 9 11 9 2 7 3 2 2
21 13 0 9 11 15 0 0 9 7 3 9 3 0 13 9 15 13 2 13 9 2
4 16 15 3 2
19 15 13 3 16 2 3 16 16 10 9 13 13 3 12 9 9 7 3 2
13 9 13 3 9 13 3 7 13 9 13 12 9 2
6 13 9 7 15 9 2
7 9 1 15 13 9 11 2
9 11 13 9 3 13 0 9 11 2
6 13 9 3 12 9 2
4 13 15 13 2
22 2 16 15 13 0 2 2 11 13 10 9 7 9 2 2 13 15 3 13 9 2 2
7 9 13 0 13 9 13 2
10 7 15 13 3 0 16 15 13 9 2
8 3 15 13 11 16 13 15 9
5 10 9 13 9 3
11 13 9 13 15 13 9 0 2 0 9 2
4 2 6 6 2
7 3 13 10 0 9 13 2
15 13 7 3 16 13 15 3 15 3 3 13 13 12 9 2
8 9 13 0 9 9 0 9 2
8 13 9 15 9 16 13 9 2
11 13 3 13 9 2 7 15 13 0 9 2
12 9 13 13 13 13 15 13 3 3 9 9 2
13 0 9 13 12 0 11 11 9 11 7 11 9 2
8 15 13 9 1 2 9 1 2
8 15 13 9 1 2 9 1 2
14 7 3 13 11 3 1 11 2 13 3 13 9 9 2
6 11 11 13 1 9 2
7 11 2 15 13 13 3 2
6 9 9 3 13 9 2
12 13 13 10 9 7 10 0 9 11 9 13 2
6 15 13 13 3 3 2
5 2 13 15 13 2
12 9 9 13 9 13 9 7 13 0 1 9 2
8 0 9 13 13 3 16 13 2
7 11 13 3 9 9 1 2
2 10 9
14 15 13 13 10 9 9 16 15 13 15 2 11 13 2
2 10 9
5 9 13 9 13 9
10 9 7 9 13 15 0 12 12 9 2
10 9 9 13 3 13 9 0 12 9 2
10 15 13 3 13 9 3 0 9 9 2
16 9 1 15 13 9 3 2 9 9 13 13 13 3 13 13 2
9 16 15 13 9 2 13 13 13 2
16 3 16 13 9 9 9 2 3 9 13 3 0 9 9 13 2
2 13 13
5 13 3 13 9 2
7 9 13 13 3 0 9 2
4 11 13 0 9
6 11 15 13 9 9 2
8 9 12 9 1 13 10 9 2
11 9 13 13 15 2 16 15 13 13 9 2
15 0 9 13 9 9 1 3 3 3 2 16 15 3 13 2
6 13 3 13 10 9 2
14 0 9 9 13 13 0 9 2 15 9 13 13 13 2
5 9 9 13 13 2
17 11 13 16 9 2 15 13 13 13 12 9 2 13 13 13 9 2
2 13 3
17 10 9 9 2 13 10 9 0 7 0 2 13 13 3 13 9 2
10 10 9 13 9 13 3 7 15 13 2
8 11 13 13 10 9 16 15 2
3 9 0 2
6 9 13 9 11 1 9
15 11 7 11 9 13 10 9 2 15 10 3 13 3 13 2
16 3 3 13 9 2 15 13 9 11 7 13 9 10 9 3 2
11 13 15 9 2 3 13 10 0 9 3 2
5 3 15 13 13 2
7 15 13 9 3 9 1 2
4 13 13 0 2
10 3 13 9 2 16 13 9 13 3 2
9 11 9 13 3 12 9 3 0 2
2 10 9
5 13 3 13 9 3
3 3 0 9
3 15 13 2
4 13 9 3 2
2 13 13
44 3 2 3 15 13 9 2 3 15 13 12 13 9 1 10 9 2 9 1 13 9 2 13 0 2 7 3 3 0 16 15 1 13 13 9 2 16 13 9 7 10 9 9 2
4 13 13 3 2
5 0 9 13 0 9
9 13 15 3 13 2 13 15 13 2
2 9 2
11 12 0 7 3 0 9 7 9 13 9 2
3 3 13 9
8 13 15 9 9 9 7 9 2
8 9 13 15 13 13 9 9 2
8 9 3 13 13 2 9 2 2
14 12 9 9 13 3 3 9 12 9 13 9 7 9 2
6 6 3 11 7 11 2
2 13 9
7 13 3 3 13 2 3 2
10 0 7 0 13 3 0 7 3 0 2
2 9 13
5 13 3 13 13 13
9 9 13 2 15 13 13 3 13 2
10 9 13 13 9 0 9 2 13 11 2
10 7 3 13 10 9 15 13 0 9 2
2 15 13
4 9 13 3 2
8 15 15 3 13 10 0 9 2
16 9 9 13 13 9 2 16 7 16 9 13 2 3 13 9 2
6 3 11 13 13 9 2
12 15 13 3 3 9 2 15 3 3 13 9 2
9 9 13 9 9 3 15 15 9 2
9 9 13 13 9 2 7 9 3 2
7 15 13 3 3 0 9 2
10 0 9 9 11 9 9 13 0 9 2
12 13 13 3 9 3 7 13 9 2 7 3 2
3 9 13 9
5 3 9 9 13 2
3 15 13 3
10 16 13 15 13 3 13 15 13 13 2
3 9 7 9
14 3 3 13 15 10 9 3 13 15 3 0 9 7 2
4 9 13 9 2
3 13 13 9
7 9 0 9 13 3 12 2
11 16 15 13 7 15 13 3 13 13 9 2
12 13 3 3 11 2 16 13 3 15 13 13 2
6 13 2 3 15 13 2
8 11 13 0 2 7 15 13 2
8 9 1 13 13 0 7 13 2
17 13 9 9 13 11 9 12 2 3 16 11 13 2 7 9 12 2
2 9 9
9 9 1 2 3 9 13 13 9 2
10 11 13 0 9 2 15 13 9 3 2
7 9 0 15 13 0 9 2
3 12 9 9
16 9 13 13 9 9 2 7 15 13 0 9 13 0 3 0 2
3 9 9 9
6 15 13 13 13 11 2
2 9 9
8 3 13 13 3 12 9 9 2
17 0 11 9 11 11 2 9 2 13 3 11 13 9 15 2 15 2
9 13 9 2 16 13 15 15 9 2
13 13 15 9 2 11 13 2 16 11 13 9 9 2
4 13 9 3 2
12 13 15 13 2 16 15 10 0 9 13 9 2
6 6 6 2 13 13 2
12 16 0 13 2 13 10 9 13 9 9 13 2
3 9 13 3
9 9 1 9 13 0 3 1 11 2
11 9 9 13 3 13 9 13 9 0 9 2
13 12 9 1 11 13 13 2 3 3 3 9 13 2
8 9 13 3 9 3 7 9 2
2 0 9
4 13 3 9 2
8 12 9 11 13 9 9 9 2
5 10 9 13 13 2
8 0 15 13 13 16 13 9 2
10 15 1 9 10 9 11 13 11 13 2
11 7 15 13 15 3 9 9 3 3 3 2
10 11 1 0 11 13 9 2 0 9 2
17 16 15 13 3 9 3 9 3 13 13 3 0 9 16 15 13 2
11 11 13 0 2 7 16 15 13 3 9 2
9 9 9 13 13 9 8 7 9 2
9 0 9 12 9 9 13 3 9 2
16 11 9 9 13 16 15 13 3 0 2 3 12 9 2 9 2
5 13 0 13 0 2
11 9 13 13 3 2 9 2 0 9 3 2
14 0 9 9 13 3 3 15 2 15 3 11 13 13 2
2 10 9
21 13 9 2 3 9 13 0 13 10 9 2 16 15 3 13 10 9 16 13 13 2
10 9 12 1 9 13 9 1 12 12 2
5 9 13 13 9 2
3 9 13 11
9 13 0 9 16 11 13 3 13 2
11 13 15 15 13 16 13 10 0 13 2 2
7 13 9 13 13 15 0 2
3 9 13 9
11 9 9 13 13 3 2 3 9 13 0 2
4 11 13 13 2
6 0 9 15 3 13 2
3 13 3 2
8 9 12 9 13 0 9 1 2
17 7 16 3 13 2 13 13 13 3 13 2 16 13 9 7 9 2
3 13 13 2
5 9 13 9 9 13
2 0 9
7 11 1 9 13 3 9 2
9 12 9 9 9 13 13 13 9 2
7 11 11 13 9 3 9 2
4 0 9 13 9
13 9 13 3 2 3 13 10 9 2 16 11 13 2
13 13 3 13 2 16 15 13 3 13 3 0 9 2
3 9 13 0
6 13 15 10 0 9 2
3 9 13 9
6 9 3 13 0 9 2
9 13 13 9 3 16 15 13 9 2
7 9 13 13 3 3 12 2
15 9 13 3 13 9 12 3 13 9 7 13 15 10 9 2
12 12 0 9 13 0 9 13 11 9 7 9 2
9 9 13 13 2 15 9 13 13 2
8 15 13 13 9 13 15 9 2
15 11 13 3 11 9 9 12 7 12 2 15 13 0 9 2
11 9 13 3 12 12 7 9 12 12 9 2
7 11 13 3 13 9 9 2
13 11 13 12 12 9 7 9 9 9 0 0 9 2
7 13 15 2 13 9 15 2
8 10 9 13 13 9 3 3 2
7 0 9 13 3 0 11 2
13 9 13 15 9 9 2 13 15 3 2 13 15 2
4 15 13 13 2
6 13 3 9 13 13 2
11 16 15 9 12 13 11 2 9 13 0 2
18 2 3 13 3 13 13 13 9 2 16 13 13 2 2 11 11 13 2
14 7 13 3 2 16 9 9 13 3 0 9 0 3 2
7 9 13 0 7 3 0 2
9 11 9 9 13 13 3 3 0 2
16 9 13 13 3 9 12 9 2 7 0 9 13 13 15 9 2
5 13 15 3 13 2
4 9 13 15 2
17 0 9 12 15 2 15 13 0 9 2 13 12 12 9 9 9 2
16 11 9 13 0 13 3 2 16 10 9 13 9 0 0 9 2
3 13 9 2
8 9 13 0 2 15 9 13 2
7 15 13 9 9 1 9 2
11 15 9 13 13 13 9 13 9 9 9 2
25 15 13 3 0 3 10 3 13 9 7 7 3 3 3 15 13 9 9 9 11 7 13 13 9 2
2 13 9
11 16 9 13 12 12 13 7 13 13 13 2
6 15 13 7 13 9 2
2 0 9
6 11 9 13 9 0 2
6 9 13 13 12 13 2
21 3 0 13 13 15 2 10 9 13 9 2 7 15 2 13 9 9 1 2 9 2
17 13 9 10 9 12 7 12 7 3 13 9 1 9 7 13 9 2
6 9 13 13 13 9 2
11 3 13 13 0 9 2 15 13 3 3 2
8 15 13 13 9 2 15 13 2
7 9 13 3 9 9 1 2
13 13 0 13 0 7 13 9 9 2 15 13 9 2
9 16 9 9 11 13 9 3 9 2
17 9 9 13 0 9 9 2 0 9 2 13 0 3 0 1 13 2
3 3 9 13
10 16 9 13 2 15 13 13 9 1 2
5 15 13 11 9 2
4 9 13 9 2
5 9 13 13 9 2
8 10 9 9 9 13 15 9 2
17 15 13 3 9 13 13 3 0 9 2 7 3 0 15 13 9 2
12 15 13 15 2 13 15 15 16 15 13 0 2
5 15 13 13 3 2
7 10 9 15 3 3 13 2
13 0 9 13 12 3 2 16 0 9 13 12 3 2
3 13 9 1
12 13 0 9 13 3 3 0 2 11 11 13 2
5 15 13 13 3 2
8 13 9 13 3 2 13 9 2
16 9 9 13 3 13 2 16 15 13 2 16 15 3 13 13 2
4 15 15 13 2
6 9 13 9 0 3 9
6 15 13 13 9 9 2
2 9 9
3 9 9 9
8 15 13 3 13 13 9 3 2
5 11 13 13 9 2
3 13 3 2
6 7 15 13 0 9 2
9 3 13 13 12 0 9 13 9 2
7 13 13 13 3 0 9 2
13 11 13 9 9 3 2 9 7 9 13 3 3 2
7 9 15 13 3 0 13 2
5 15 13 9 1 2
4 15 13 9 9
9 7 0 7 0 9 13 0 9 2
4 13 9 0 2
6 13 13 3 9 12 1
8 0 9 9 13 13 0 9 2
18 15 13 11 9 10 9 2 16 13 2 3 9 13 13 3 9 1 2
3 9 13 0
9 15 13 3 0 9 2 13 11 11
5 9 12 9 12 2
2 10 9
14 3 2 16 13 0 9 2 13 7 13 7 13 9 2
2 3 3
5 15 13 3 11 2
8 10 9 15 13 12 10 9 2
14 9 15 13 11 9 13 9 9 13 9 8 8 8 2
8 11 9 13 16 0 9 9 2
12 9 13 3 2 7 3 15 13 13 3 3 2
4 11 9 13 2
7 11 13 9 12 11 9 2
2 0 15
5 3 9 13 3 3
6 15 13 15 13 9 2
6 13 3 2 15 13 2
16 11 13 9 9 13 3 13 12 0 9 7 10 9 12 9 2
8 9 13 2 16 13 13 3 2
2 0 9
6 0 15 13 3 13 2
32 11 13 15 3 12 9 7 2 13 10 8 15 13 13 3 3 13 13 15 13 3 3 7 2 9 13 12 7 15 15 13 2
4 9 1 9 2
17 13 15 13 13 11 7 7 15 13 13 10 9 2 7 13 15 2
5 0 9 3 13 2
5 9 13 3 9 2
4 3 0 9 2
2 13 13
5 13 15 3 9 2
2 9 13
15 11 11 2 10 9 9 13 2 13 9 9 7 13 3 2
14 9 9 13 15 13 13 9 2 9 13 13 3 13 2
7 13 0 7 13 9 9 2
4 15 13 0 0
11 0 13 13 9 12 9 7 15 13 0 2
2 3 16
5 13 9 3 9 2
7 9 13 3 2 13 3 2
20 3 9 2 9 2 9 2 0 9 7 9 7 10 0 9 9 9 9 13 2
6 15 13 3 9 3 9
4 11 13 11 2
7 3 11 13 13 3 10 9
9 9 13 0 2 16 13 13 15 2
6 9 13 9 13 9 2
8 2 12 0 9 13 12 9 2
8 9 13 3 0 16 0 9 2
2 1 9
5 9 1 13 9 2
4 3 13 0 9
4 0 13 0 2
16 9 13 10 9 3 0 2 7 3 15 13 13 3 9 3 2
3 13 13 2
11 15 13 15 9 2 3 15 13 0 9 2
13 9 9 13 12 10 9 13 10 9 1 9 9 2
6 15 13 0 9 1 2
4 13 12 9 2
8 11 13 2 16 9 13 13 2
11 0 9 9 7 3 9 9 13 13 9 2
8 13 13 13 3 1 9 9 2
7 9 9 7 9 1 13 2
10 16 9 13 9 2 13 9 9 15 2
10 16 3 13 3 13 3 7 13 15 2
2 6 6
13 3 3 0 9 9 13 9 11 11 7 9 13 2
10 9 13 13 7 13 3 7 3 3 2
9 13 13 9 11 9 9 9 9 2
10 3 13 9 9 2 13 9 9 13 2
27 9 13 3 13 2 7 9 9 2 9 9 2 9 7 9 9 2 9 9 2 9 7 9 9 13 15 2
9 9 13 9 0 7 9 13 9 2
6 15 13 9 9 9 2
7 15 10 9 3 13 10 9
7 13 11 0 9 9 13 2
13 13 12 9 9 3 8 2 8 2 8 7 9 2
8 13 9 2 16 13 3 9 2
3 12 9 9
7 3 15 13 13 0 9 2
19 10 9 3 13 13 9 7 3 10 9 9 13 3 0 9 9 7 9 2
9 0 7 0 9 13 3 0 2 2
12 15 1 13 13 13 3 16 15 13 3 0 9
6 15 13 3 9 1 3
5 9 9 13 0 2
6 15 13 13 3 0 2
10 9 13 3 2 13 9 13 9 9 2
11 3 13 11 9 2 16 9 13 13 13 2
4 3 13 0 9
9 15 13 0 7 15 13 0 9 2
2 9 11
23 11 13 3 9 2 15 0 9 9 13 3 13 13 13 15 2 16 9 3 13 3 3 2
14 9 7 0 9 13 10 9 16 13 9 9 7 9 2
5 15 13 0 9 2
16 9 13 2 16 16 9 9 13 2 15 13 13 9 9 3 2
3 9 9 2
5 0 9 13 0 2
6 3 13 9 13 9 2
5 10 12 13 9 2
4 15 13 3 13
12 11 11 11 7 11 11 9 9 13 3 13 2
10 3 3 3 9 13 9 13 9 1 2
16 9 13 13 13 13 9 2 9 3 0 0 13 13 3 13 2
8 11 15 13 9 9 12 9 2
10 15 13 13 3 16 13 3 13 0 2
22 9 13 11 9 9 9 7 13 3 10 9 2 9 9 2 3 15 13 13 10 9 2
9 10 9 9 13 13 13 9 9 2
15 8 8 9 9 11 11 1 11 13 3 13 13 3 11 2
2 13 9
11 9 9 13 9 2 15 13 13 0 9 2
5 15 13 3 0 2
9 8 7 8 8 13 9 11 9 2
10 16 9 13 0 2 13 9 9 13 2
23 3 9 13 10 9 2 10 9 13 9 11 0 12 9 15 3 2 7 13 9 3 13 9
15 16 9 13 8 11 2 3 9 13 3 0 15 9 13 2
8 3 10 9 15 13 10 9 2
2 13 9
2 13 3
10 11 11 9 13 0 9 3 9 12 2
15 10 9 13 11 2 7 3 11 13 13 15 9 9 11 2
2 8 2
11 13 15 0 9 16 15 13 13 9 9 2
3 9 13 2
8 3 0 15 13 2 11 9 2
12 9 13 13 9 0 9 2 9 13 9 13 2
4 13 12 9 2
4 9 7 9 2
7 3 15 13 13 11 13 2
7 9 9 13 3 3 9 2
17 10 12 9 13 9 0 9 3 9 1 7 3 9 3 9 1 2
5 15 13 9 13 9
11 3 13 2 16 9 15 9 13 13 0 2
5 10 11 10 12 9
13 11 9 13 11 0 9 2 15 13 3 12 9 2
8 6 16 10 9 15 13 13 2
6 9 0 13 3 9 2
11 3 13 13 3 13 13 9 13 9 9 2
6 0 13 3 3 9 2
2 0 11
7 9 13 13 0 13 9 2
13 11 11 13 9 13 13 2 16 9 13 13 3 2
7 9 13 0 0 12 9 2
5 9 13 9 1 2
6 15 13 13 15 3 2
6 3 10 9 13 13 2
9 10 9 9 13 13 3 0 9 2
3 10 9 9
4 13 3 0 2
5 13 15 9 9 2
8 0 9 13 9 13 3 13 2
3 13 9 1
5 9 15 13 9 2
5 13 13 13 15 2
14 9 13 9 11 13 2 9 15 10 9 13 13 13 2
3 15 13 0
4 13 3 9 2
10 15 13 3 3 9 13 9 3 15 2
11 9 11 2 11 2 13 13 0 3 3 2
7 9 9 13 9 3 3 2
2 9 9
5 9 13 3 3 2
7 13 2 16 15 13 11 2
5 9 13 0 9 2
9 15 13 9 13 13 9 0 9 2
6 9 13 11 3 15 2
5 3 9 16 3 9
11 11 13 0 9 1 0 9 3 0 9 2
6 11 13 15 3 9 2
7 11 7 15 13 0 9 2
7 15 15 3 13 2 16 2
11 9 13 0 13 9 2 15 13 0 9 2
16 13 13 9 13 10 9 7 9 0 9 13 13 15 3 13 2
12 9 13 2 13 13 15 2 15 13 0 9 2
6 15 13 3 3 10 9
2 9 1
14 8 11 9 13 3 13 7 13 2 9 7 9 13 2
10 3 15 0 9 13 3 3 9 3 2
9 15 13 3 0 0 9 10 9 2
5 15 13 12 9 1
7 16 15 3 13 10 0 2
10 10 9 2 15 15 13 2 13 9 2
2 9 9
13 11 13 13 9 3 3 3 12 9 1 10 9 2
10 13 15 13 9 7 13 9 9 9 2
11 3 16 9 13 9 2 9 13 10 9 2
4 9 13 12 9
5 3 15 15 13 2
5 3 13 9 9 2
4 13 3 13 2
5 15 15 3 13 2
10 7 15 13 13 13 3 3 13 9 2
6 13 11 10 0 9 2
6 9 13 9 13 9 2
9 0 9 9 9 13 13 9 1 2
10 11 13 9 3 9 7 9 9 9 2
12 9 1 9 9 2 9 3 2 13 10 9 2
7 11 9 13 15 0 2 2
14 15 1 13 3 9 11 9 2 15 13 13 9 11 2
6 13 3 13 15 15 2
4 3 13 13 2
3 10 0 9
5 11 13 3 9 2
10 13 15 13 15 16 13 15 3 3 2
39 7 16 15 13 9 9 7 15 13 10 9 7 10 9 2 7 16 15 13 10 9 2 3 16 13 9 13 2 7 15 13 13 9 2 13 15 15 13 2
7 15 13 3 0 9 9 2
2 6 9
10 11 7 11 0 9 9 13 9 13 2
8 11 9 13 9 12 9 1 2
7 3 13 3 13 13 9 2
11 15 13 13 10 11 9 9 10 10 9 2
5 11 9 11 1 2
9 3 11 13 2 0 9 9 13 2
3 3 3 2
7 9 11 13 9 11 9 2
6 11 7 11 13 15 2
7 3 13 13 3 10 9 2
18 0 9 13 7 13 13 10 9 16 9 9 2 3 7 3 7 10 9
6 13 3 13 13 0 2
8 11 3 13 0 9 9 9 2
5 15 9 3 13 2
5 13 13 0 9 2
14 7 15 13 15 7 10 15 13 15 9 13 9 9 2
32 15 13 16 6 16 15 13 13 7 15 13 16 10 9 13 3 8 9 3 3 16 3 16 15 13 3 9 3 15 15 13 2
12 3 0 15 13 13 13 0 9 0 9 11 2
3 13 11 9
4 13 15 13 2
4 9 13 3 2
8 13 9 3 7 9 3 3 2
5 9 13 9 9 2
10 15 13 9 3 12 7 13 3 9 2
8 9 13 13 11 7 9 9 2
2 11 9
14 11 11 1 11 13 13 3 13 13 9 3 0 9 2
2 13 9
11 12 9 1 0 9 13 13 9 11 1 2
9 13 0 7 13 2 13 13 3 2
11 9 13 13 9 10 9 2 15 9 13 2
13 9 15 13 11 9 9 15 13 0 9 9 9 2
10 13 0 2 16 3 0 13 15 0 2
3 13 15 13
5 15 13 9 15 2
5 13 9 3 9 2
8 13 13 3 3 10 12 9 2
11 11 2 12 2 13 9 13 3 9 1 2
8 9 1 15 13 9 9 9 2
10 13 13 2 0 9 15 3 11 13 2
4 13 3 13 13
10 15 9 13 2 16 13 13 10 9 2
3 15 13 13
3 15 13 2
3 3 13 9
18 13 3 2 16 0 9 10 9 13 2 15 9 13 2 13 3 9 2
7 9 13 13 3 12 9 2
8 16 9 13 2 13 13 0 2
11 0 9 13 9 13 13 13 13 15 3 2
3 11 13 13
4 11 13 9 2
9 13 11 9 13 13 9 0 9 2
22 9 13 13 9 0 0 9 2 15 13 0 9 13 15 2 15 13 9 3 7 3 2
7 9 13 9 1 10 9 2
34 15 13 3 3 3 3 3 7 13 13 10 10 0 9 7 3 15 13 0 9 16 3 15 3 3 3 13 16 2 15 13 9 3 2
13 3 13 9 2 1 9 2 13 3 2 13 9 2
3 9 13 2
10 15 13 3 9 2 0 9 7 9 2
7 13 2 16 13 15 3 2
6 9 13 10 9 3 2
12 9 11 11 13 2 16 9 13 9 9 9 2
9 3 9 13 11 9 9 11 11 2
13 16 11 9 13 0 9 2 9 13 13 13 9 2
5 9 2 13 13 2
14 9 13 3 13 3 15 2 16 9 13 13 3 9 2
6 11 13 9 1 9 2
8 13 13 3 13 0 13 0 2
7 13 15 15 3 3 13 2
5 10 9 13 3 2
8 9 11 11 13 11 9 9 2
18 11 15 13 3 0 9 13 9 2 16 13 13 2 16 13 13 2 2
5 3 12 9 9 2
3 13 3 2
9 15 13 2 16 15 13 9 9 2
5 15 13 3 13 2
23 9 13 12 9 2 9 12 9 7 12 9 2 9 7 9 2 7 9 13 13 3 9 2
3 13 3 9
7 13 9 7 13 3 9 2
2 9 9
7 0 9 13 13 9 13 2
6 9 13 2 16 13 2
17 13 11 11 7 13 16 11 13 9 7 13 13 3 0 9 3 2
5 15 13 0 9 2
5 11 13 13 3 2
3 13 11 2
8 9 0 9 13 9 11 11 2
4 15 13 0 2
13 9 13 13 9 2 7 15 13 13 9 0 9 2
3 13 11 9
7 11 13 3 12 9 9 2
4 13 3 9 2
19 16 13 13 3 9 2 15 13 3 0 13 3 2 16 13 13 9 9 2
3 13 9 2
21 13 13 13 2 12 1 2 15 2 15 13 9 2 9 7 9 13 0 0 9 2
9 9 3 13 3 3 16 15 13 2
4 9 13 13 2
2 15 2
4 15 13 3 15
11 11 7 11 13 3 0 9 3 9 9 2
6 11 9 13 0 9 2
10 12 0 13 11 12 9 9 13 9 2
29 0 13 2 16 13 10 9 2 15 9 13 3 2 13 13 10 0 9 2 3 3 10 9 2 7 15 13 9 2
2 10 9
2 9 9
2 0 9
14 16 9 13 9 1 2 9 13 13 9 9 0 9 2
6 15 3 3 9 9 2
6 3 10 9 13 0 2
7 11 11 9 9 13 0 2
9 10 9 9 0 9 13 9 11 2
15 15 13 2 16 13 9 3 7 13 2 16 13 13 15 2
12 9 13 9 2 15 13 3 0 12 9 9 2
15 9 13 3 13 3 0 9 2 15 13 15 9 7 9 2
5 13 3 9 16 2
4 9 9 7 9
6 0 2 0 7 0 9
12 11 11 11 13 0 9 12 9 13 9 9 2
5 9 13 9 9 2
7 9 13 9 9 12 9 2
9 13 9 13 0 9 13 15 9 2
5 9 15 13 13 2
5 13 13 3 12 2
4 13 3 9 2
20 2 15 13 0 9 2 11 13 12 9 13 9 2 13 13 3 12 9 2 2
6 13 13 9 3 13 2
8 15 13 0 2 16 13 13 2
14 13 3 15 2 9 13 2 2 3 15 13 10 9 2
10 15 13 10 0 3 2 3 9 13 2
21 15 13 16 3 3 13 13 15 13 3 3 7 2 9 13 12 7 15 15 13 2
5 15 13 13 9 1
6 9 13 0 9 1 2
15 16 15 13 13 2 9 13 0 9 2 9 13 9 1 2
7 15 13 9 1 13 9 2
9 3 9 13 9 9 7 0 9 2
9 9 13 3 10 0 9 10 9 2
8 9 7 9 9 13 0 9 2
7 15 13 13 9 9 1 2
7 9 13 3 2 13 3 2
3 15 13 13
3 9 9 15
4 9 13 9 2
22 11 13 9 13 3 2 13 9 1 15 1 2 9 15 2 16 0 15 13 9 9 2
13 9 13 9 9 2 9 7 9 1 9 7 9 2
5 9 13 9 0 2
3 15 13 2
3 3 3 2
6 15 3 13 13 9 2
5 11 13 15 9 2
13 9 15 13 13 12 9 2 15 13 9 0 9 2
5 9 13 13 11 2
4 9 13 9 2
9 16 3 13 13 2 13 13 9 2
7 9 13 13 3 12 9 2
6 6 13 15 3 0 2
6 9 1 13 3 9 2
13 16 9 13 9 2 15 13 3 13 0 0 9 2
10 13 3 9 13 2 16 13 3 9 2
8 13 13 3 0 2 3 9 2
7 6 2 13 15 0 9 2
13 16 11 13 0 10 9 9 2 13 9 0 9 2
18 16 3 9 12 0 9 9 13 13 0 9 2 13 9 3 0 9 2
8 11 13 11 9 0 12 9 2
10 13 13 3 9 7 0 9 13 9 2
20 0 9 3 13 9 15 2 16 15 13 13 9 0 2 13 7 13 0 9 2
6 11 13 3 2 0 2
16 11 13 3 0 3 15 2 15 0 9 2 3 15 9 13 2
19 9 13 0 9 3 12 12 9 9 2 16 13 8 7 9 9 11 9 2
6 13 9 13 13 10 9
10 9 7 9 13 3 13 0 9 9 2
4 15 13 0 9
8 9 9 13 9 10 12 9 2
19 13 9 16 10 9 2 9 9 12 2 9 3 9 9 1 7 3 13 2
13 13 15 13 13 16 15 13 13 0 9 7 0 9
17 11 13 2 13 9 13 2 13 9 9 13 10 9 13 9 2 2
5 3 3 9 1 2
6 6 16 15 13 3 2
7 13 9 15 3 9 13 2
2 11 9
5 13 9 9 3 2
5 15 13 13 9 2
7 9 13 12 9 13 9 2
16 9 13 3 9 9 2 13 3 10 0 12 12 9 9 13 2
4 13 9 15 2
8 13 11 10 9 9 3 3 2
9 3 9 7 9 13 9 12 9 2
7 10 9 9 9 3 13 2
11 10 9 13 13 9 9 9 2 9 13 2
4 9 13 9 2
5 3 9 13 0 2
8 9 13 13 2 16 9 13 13
5 15 13 3 3 2
15 11 13 15 13 15 10 0 9 1 2 15 15 9 13 2
10 13 13 9 7 10 0 9 9 1 2
10 9 2 3 0 2 13 15 9 9 2
14 9 13 9 3 10 2 10 9 2 7 3 0 9 2
10 0 9 9 11 11 13 3 3 13 2
9 3 3 13 3 13 9 3 16 2
11 9 13 3 3 13 3 9 7 9 9 2
9 0 12 9 13 11 11 1 12 9
9 3 15 13 15 15 15 15 0 13
3 15 13 9
14 9 10 9 13 13 9 3 9 2 16 9 13 13 2
9 15 13 9 3 7 13 9 9 2
6 15 13 15 0 9 2
4 11 12 9 9
2 0 9
9 0 9 13 2 3 9 13 0 2
6 10 9 15 15 13 2
15 11 13 13 13 2 16 0 9 7 0 13 13 3 11 2
14 3 13 9 13 9 1 2 7 15 13 3 12 9 2
10 9 13 13 0 13 3 9 13 3 2
18 0 9 9 13 3 2 16 9 0 9 7 10 0 1 13 13 9 2
4 11 13 13 2
4 13 13 0 9
8 13 13 15 9 3 0 9 2
14 15 3 13 10 9 16 8 13 3 16 3 13 13 15
4 9 3 0 9
8 13 11 3 13 13 0 9 2
5 9 15 13 15 13
5 15 13 13 9 2
4 13 3 9 2
7 10 9 13 13 9 9 2
11 15 13 13 13 0 2 10 9 15 13 2
5 9 9 13 0 9
5 9 2 9 7 9
7 9 13 3 9 2 15 2
10 13 13 16 2 16 3 12 9 9 2
14 11 13 9 12 9 2 7 15 13 7 9 7 9 2
14 13 13 16 13 15 0 9 2 16 3 15 3 13 2
6 13 3 3 13 3 2
6 10 9 13 12 9 2
7 0 2 15 13 13 9 2
10 11 13 0 7 0 9 3 3 9 2
7 3 15 13 13 3 0 2
16 9 13 3 13 9 2 15 13 13 2 15 13 13 9 2 2
5 3 3 13 9 2
3 9 13 9
4 9 13 9 2
10 9 13 13 13 2 9 13 15 13 2
16 10 9 9 15 3 13 2 9 13 2 2 16 13 13 9 2
2 0 9
4 9 13 1 9
12 9 13 0 13 2 15 13 0 7 0 9 2
5 13 9 9 11 2
10 11 7 11 9 13 11 2 11 11 2
15 9 12 9 9 13 12 7 15 13 3 12 13 9 12 2
2 13 9
5 15 13 13 9 2
11 15 13 9 9 2 11 2 11 7 11 2
13 11 7 11 13 13 3 0 9 2 15 13 9 2
6 15 13 0 16 15 2
13 15 13 13 9 9 7 13 13 3 3 3 0 2
6 11 13 9 9 9 2
8 11 9 13 3 13 9 15 2
15 9 13 0 9 7 9 2 7 12 9 13 13 7 13 2
11 9 13 9 13 3 13 0 13 9 9 2
9 13 3 13 2 13 3 7 13 2
5 13 3 13 13 2
6 15 13 9 10 9 2
3 13 10 9
4 15 15 13 2
22 3 15 13 9 9 3 15 1 2 16 11 13 9 2 13 2 16 13 15 9 13 2
6 13 3 10 0 9 2
9 16 15 13 13 2 3 3 13 2
6 13 9 7 13 13 2
8 0 13 13 3 3 16 13 2
4 6 3 3 2
3 0 13 2
6 0 9 15 13 9 2
15 11 13 0 9 2 11 9 9 2 10 0 9 9 13 2
2 0 9
6 0 9 13 3 0 2
4 13 0 9 9
5 13 0 13 13 2
7 0 9 13 9 7 9 2
5 9 1 13 9 2
10 15 13 3 0 9 7 3 0 9 2
6 13 13 9 0 9 2
12 11 9 11 9 13 0 7 13 3 3 0 2
5 15 13 13 10 9
19 16 9 12 9 13 13 12 12 9 2 3 9 12 9 13 12 12 9 2
6 15 13 9 16 9 2
8 13 15 3 15 3 9 9 2
10 9 13 13 10 9 9 3 12 9 2
9 13 9 10 0 9 10 0 9 2
7 9 13 15 1 2 9 2
6 11 13 11 9 9 2
16 0 9 13 13 0 2 16 15 13 0 2 13 3 13 9 2
7 15 13 3 13 0 9 2
8 9 13 13 9 7 3 9 2
8 9 13 13 2 13 9 13 2
9 3 9 13 9 1 3 12 9 2
6 11 11 13 16 9 2
6 15 3 13 3 9 2
3 13 0 13
2 9 9
4 15 13 0 9
6 15 13 9 13 9 2
4 13 3 13 2
6 15 13 0 9 9 2
18 3 0 9 13 3 13 9 9 9 2 3 16 9 13 0 7 0 2
15 3 3 13 13 10 9 2 16 11 7 11 13 15 9 2
8 2 13 3 15 10 9 3 2
7 9 13 3 9 1 9 2
7 13 2 16 3 13 9 2
6 9 13 13 15 13 2
5 0 9 3 13 2
8 9 13 3 9 0 9 3 2
11 15 2 16 9 13 13 9 2 13 9 2
2 0 9
10 16 13 3 13 2 13 3 12 9 2
7 13 3 9 9 7 9 2
15 16 9 13 3 0 3 3 13 13 9 7 9 13 0 2
12 11 9 13 12 7 0 2 15 13 13 9 1
5 15 13 13 9 2
11 11 13 13 9 9 13 15 3 13 15 2
10 9 9 1 9 13 0 0 13 9 2
7 15 13 9 15 7 15 2
4 3 0 11 2
8 0 13 0 9 0 9 3 2
6 15 13 3 13 3 2
19 9 7 9 13 3 11 9 0 9 9 2 16 15 3 9 1 13 9 2
5 11 13 9 9 2
4 11 9 13 13
18 16 0 9 9 13 12 9 9 2 3 13 3 2 15 10 9 13 2
10 10 0 13 2 13 3 0 13 15 2
17 9 11 9 11 11 7 9 11 13 13 9 9 2 9 9 2 2
7 3 9 13 9 3 9 2
5 15 15 13 3 2
5 3 9 9 13 2
16 11 9 13 3 8 2 15 13 16 15 13 12 9 3 9 2
9 13 9 2 13 9 3 10 9 2
7 2 15 13 13 3 3 2
16 13 13 3 15 2 16 9 13 3 2 16 15 13 0 13 2
7 0 13 13 0 9 9 2
2 9 11
17 15 13 12 9 9 2 11 11 13 7 13 12 0 2 0 9 2
4 13 9 9 1
8 9 13 0 2 15 13 9 2
7 15 13 13 13 7 13 2
4 9 9 7 9
9 0 9 13 9 7 11 13 9 2
4 15 13 13 2
7 9 13 0 9 2 0 2
13 9 7 9 13 12 9 9 2 7 3 0 0 2
12 11 9 0 9 13 0 9 3 0 9 11 2
8 9 13 10 9 11 0 12 2
7 11 2 13 15 3 9 2
6 13 13 3 9 1 2
9 13 0 13 9 2 15 13 0 2
6 13 9 13 10 9 2
19 15 13 13 9 2 16 16 9 13 9 9 3 2 9 13 3 9 3 2
9 13 13 3 15 2 15 3 13 2
10 3 9 1 13 9 1 9 13 13 2
9 9 13 13 3 16 0 9 1 13
6 7 13 15 2 11 2
9 13 3 13 16 13 15 13 9 9
3 9 13 2
3 3 13 9
3 9 13 13
4 3 13 0 9
7 15 13 13 0 0 9 2
19 16 0 9 9 13 13 2 13 9 3 2 16 15 13 0 7 0 9 2
4 9 9 9 9
17 11 9 13 3 13 11 0 9 11 2 15 0 9 13 0 9 2
6 13 3 13 0 9 2
7 13 13 3 0 16 13 2
8 11 11 13 9 0 16 9 2
13 10 9 2 16 13 9 7 9 15 13 3 13 2
6 13 13 3 9 9 2
9 15 13 0 9 2 7 9 0 2
13 13 0 9 7 3 16 9 13 3 13 16 3 2
2 0 9
8 15 13 15 2 7 10 9 2
15 10 9 1 9 9 9 13 13 11 7 11 11 9 11 2
5 13 13 15 13 2
13 0 2 13 13 9 11 13 9 9 13 9 9 2
5 3 9 9 13 2
10 15 13 13 2 7 13 3 15 13 2
8 9 13 13 7 9 13 13 2
7 15 13 9 0 10 9 2
4 9 13 3 2
15 15 13 3 9 2 16 11 13 2 13 15 13 9 9 2
11 13 2 16 15 13 3 13 3 3 16 0
6 13 10 9 9 13 2
17 11 9 9 13 0 9 13 3 9 11 11 7 9 9 1 11 2
3 3 13 2
8 13 0 13 3 3 9 9 2
6 0 3 13 12 9 2
7 3 9 13 0 9 9 2
17 13 9 9 13 12 9 2 15 13 7 9 13 13 12 12 0 2
8 11 13 9 7 9 13 9 2
5 9 13 0 0 2
13 13 9 9 7 13 9 10 9 3 3 16 3 13
3 9 13 2
4 9 13 0 2
15 16 9 1 10 9 13 10 0 9 2 9 13 3 13 2
4 13 3 9 2
11 13 9 10 9 1 10 0 9 0 9 2
4 15 15 13 2
12 11 9 13 0 9 0 9 2 15 13 13 2
8 9 9 9 13 0 0 9 2
11 11 9 13 9 13 12 11 7 11 1 2
16 9 9 13 2 16 9 3 13 6 2 16 13 9 0 9 2
10 9 13 9 9 13 10 9 3 13 2
5 15 13 9 3 2
5 15 13 9 15 2
8 15 13 2 16 15 15 3 13
3 13 9 0
6 15 13 13 9 7 9
20 0 9 9 13 15 9 1 12 9 2 16 11 15 13 12 7 11 3 12 9
14 13 3 2 16 9 9 13 2 16 9 13 3 3 2
11 9 9 9 1 13 10 9 3 12 9 2
9 13 3 10 10 6 9 6 3 2
17 9 13 13 3 2 16 16 13 9 2 13 0 9 10 9 9 2
2 3 9
11 3 13 2 13 2 13 7 13 9 13 2
4 15 13 3 9
5 15 13 10 9 2
8 9 13 13 13 13 0 9 2
3 13 0 9
21 13 13 15 2 9 7 9 2 15 13 9 9 9 2 16 13 15 9 15 13 2
9 9 13 9 1 0 2 0 9 2
4 13 16 3 2
5 13 9 9 11 2
17 9 13 13 9 9 0 12 9 2 7 9 9 13 13 11 9 2
13 3 16 0 9 13 2 13 15 13 10 0 9 2
17 0 9 13 9 9 1 3 9 2 7 9 13 9 3 1 9 2
7 15 13 3 3 13 0 9
7 15 13 13 0 7 0 2
7 15 13 0 0 7 0 2
7 9 13 13 9 7 9 2
5 3 13 0 9 2
3 15 13 9
13 9 7 9 13 3 3 13 16 15 13 10 9 2
13 13 3 13 15 2 16 13 13 13 13 13 15 2
10 13 10 15 13 0 9 0 15 13 2
5 13 3 12 9 2
5 3 9 13 9 2
10 9 13 3 13 3 0 16 9 13 2
7 6 13 3 3 10 9 3
12 11 11 13 3 2 13 3 7 13 3 9 2
13 3 11 13 9 13 3 13 12 9 9 12 9 2
9 9 1 9 13 13 3 9 9 2
8 10 9 13 0 13 3 15 2
4 9 13 3 2
3 9 13 9
2 9 1
3 13 10 0
5 13 10 9 3 2
11 11 13 1 9 2 16 15 15 13 13 2
19 15 13 10 9 16 15 13 0 9 2 3 9 13 15 13 2 11 13 2
3 15 13 9
16 11 9 9 13 3 2 16 11 13 13 9 9 13 13 9 2
6 9 13 12 10 9 2
8 15 13 13 3 0 9 7 9
19 0 9 0 7 0 9 9 13 11 1 13 9 3 0 2 0 7 0 2
18 15 13 13 0 9 7 0 9 2 9 3 7 3 3 10 7 15 9
6 15 13 3 0 9 2
6 13 11 9 0 9 2
6 0 13 0 7 0 2
10 9 9 1 15 13 13 9 13 13 2
19 13 15 10 9 13 2 16 9 13 13 0 9 3 2 16 0 13 3 2
11 10 9 13 3 9 2 13 9 10 9 2
4 15 15 13 2
6 15 13 13 10 9 2
6 11 3 3 13 9 2
2 9 1
2 0 11
12 3 13 0 9 3 16 9 9 3 13 9 2
11 9 9 11 11 13 11 13 0 9 11 2
6 15 13 9 0 9 2
2 11 15
9 13 3 3 13 0 9 9 13 2
8 13 13 13 15 2 11 13 2
18 16 0 13 13 9 0 9 1 2 3 0 9 9 9 13 13 9 2
7 9 13 9 13 0 9 2
4 13 9 13 2
18 13 9 9 11 13 3 9 9 1 3 9 7 9 2 9 7 9 2
6 12 9 13 13 3 2
2 13 9
8 15 1 9 9 13 13 3 2
5 9 9 13 9 2
5 15 13 12 9 2
7 9 13 9 9 13 9 2
6 9 13 12 9 1 2
7 9 13 9 8 7 9 2
8 11 13 11 3 13 3 9 2
6 11 13 9 3 3 2
7 13 0 13 0 13 9 2
15 0 9 9 9 11 8 7 9 13 7 0 7 13 9 2
10 7 13 3 3 0 9 10 13 13 2
5 9 13 9 13 2
10 10 9 13 11 13 9 9 9 9 2
7 9 13 9 3 11 9 2
4 11 13 9 2
2 11 9
12 13 13 9 9 7 3 13 9 13 3 9 2
11 9 13 3 3 3 15 3 2 11 13 2
16 11 13 16 2 3 15 13 3 2 16 13 13 13 3 2 2
2 3 9
12 9 13 9 7 0 2 0 9 9 13 9 2
5 9 13 9 1 2
14 0 9 13 13 0 13 2 16 9 7 9 13 0 2
5 9 13 9 12 9
11 9 9 13 0 0 2 9 9 13 0 2
4 9 13 3 2
6 7 15 13 13 13 9
14 0 9 13 13 9 2 15 13 15 1 0 9 1 2
12 16 9 13 13 2 13 15 16 15 3 13 2
14 0 7 0 13 3 9 3 2 7 15 3 13 15 2
7 15 13 13 9 13 9 2
3 9 13 9
4 11 13 0 2
11 15 15 13 9 3 0 2 0 0 13 2
3 13 13 2
11 3 13 9 13 16 15 3 15 13 3 2
3 15 13 9
4 9 7 3 9
10 9 13 0 9 7 13 3 11 9 2
7 3 15 13 13 0 9 2
7 9 13 3 13 13 9 2
6 0 12 9 13 9 2
6 15 13 10 9 9 2
10 15 15 13 13 13 2 13 3 9 2
12 9 1 13 2 16 0 13 13 3 7 3 2
2 9 9
6 3 15 3 9 13 2
11 0 9 2 9 13 9 7 9 13 9 9
10 13 0 9 13 9 3 3 13 13 2
5 9 13 9 3 2
16 12 9 3 0 7 9 2 3 11 11 13 13 3 12 9 2
2 9 11
9 9 13 9 2 9 7 0 9 2
2 15 13
13 11 0 9 10 9 13 10 12 9 16 0 9 2
6 9 13 3 10 9 9
6 3 15 13 3 9 2
4 13 15 1 2
13 11 13 3 2 16 15 1 11 7 11 13 0 2
11 15 13 0 9 3 0 7 3 0 9 2
9 15 13 9 0 2 7 9 3 2
3 9 3 2
10 9 13 3 13 9 13 3 3 0 2
5 0 9 13 9 2
15 13 3 2 10 0 9 2 7 13 3 13 3 0 9 2
4 9 13 0 2
2 13 9
6 13 3 2 15 13 2
4 9 13 9 2
10 9 7 9 13 13 3 3 9 1 2
7 15 13 13 3 0 9 2
2 15 13
8 12 9 1 15 13 13 9 2
16 0 9 0 9 13 9 9 2 15 13 9 9 9 0 9 2
3 13 15 1
11 9 13 3 10 1 9 9 7 9 1 2
7 9 13 3 3 9 9 2
13 13 13 11 16 13 15 0 9 1 9 3 13 2
3 12 0 9
3 15 13 3
8 6 16 13 13 13 15 3 2
19 16 9 13 15 2 16 9 13 13 9 0 2 3 3 13 13 3 9 2
3 9 13 9
4 9 13 9 1
5 13 13 15 1 2
6 13 16 13 13 13 2
13 9 13 3 9 13 0 9 9 0 7 0 9 2
10 9 13 3 9 3 16 15 15 13 2
9 15 13 7 13 9 9 7 9 2
2 0 9
14 16 15 13 13 13 7 13 3 2 15 13 3 0 2
7 12 9 15 13 13 9 2
8 13 13 0 9 10 9 0 9
21 3 10 0 9 13 3 2 16 11 13 3 1 11 13 13 0 9 7 13 9 2
10 9 13 0 9 3 7 3 15 1 2
7 9 13 9 13 9 9 2
14 11 9 1 9 9 2 15 13 3 9 2 13 9 2
8 13 15 9 7 13 13 0 2
11 9 0 9 13 9 11 7 13 3 3 2
5 15 13 9 13 9
10 13 0 13 3 0 2 3 7 0 2
2 13 15
3 13 15 2
10 9 7 9 9 13 9 13 0 9 2
6 13 9 0 9 1 2
2 13 0
3 13 9 9
9 15 13 3 2 15 13 9 3 2
11 16 13 0 13 9 3 2 3 3 13 2
2 0 0
13 3 15 13 3 0 9 2 16 13 13 9 0 2
12 11 13 12 13 9 1 12 9 1 0 11 2
6 9 13 3 3 0 2
6 11 11 13 1 9 2
5 15 13 8 8 2
17 9 13 3 13 3 2 16 9 9 13 0 2 7 2 0 2 2
9 13 3 0 2 7 3 3 3 2
23 15 13 9 13 9 15 2 16 15 13 13 9 7 15 13 10 9 3 3 9 9 3 2
6 9 13 9 9 9 2
11 7 9 1 13 13 0 16 13 13 9 2
8 10 12 9 13 3 0 9 2
12 13 7 13 7 13 2 13 9 7 13 9 2
11 10 11 9 13 12 9 2 15 3 13 2
9 15 0 2 9 13 3 9 1 2
7 15 13 9 2 13 9 2
8 15 13 10 9 9 16 3 2
18 13 13 9 13 9 9 2 7 3 13 3 15 13 13 2 16 16 2
5 13 15 13 15 2
6 9 13 9 3 13 2
6 9 9 13 13 9 2
7 9 1 15 13 13 3 2
10 9 13 10 0 2 16 15 13 9 2
6 13 0 13 3 0 2
14 11 13 2 16 13 10 10 9 0 9 13 9 9 2
2 13 13
3 9 13 0
14 9 13 2 13 13 3 3 3 2 13 3 0 9 2
8 11 9 11 13 9 9 9 2
20 15 1 13 0 2 16 13 13 9 2 16 16 13 9 13 2 9 13 9 2
2 3 3
7 13 3 0 13 9 3 2
4 9 13 9 2
6 9 13 3 3 3 2
8 15 15 13 2 16 13 15 2
11 3 13 3 12 9 13 16 16 13 3 2
8 15 13 9 9 2 7 15 2
14 3 10 9 13 3 3 13 2 16 9 13 12 9 2
11 11 13 9 2 16 13 3 9 9 9 2
22 15 13 9 9 15 2 16 9 13 15 7 15 13 15 1 2 13 9 3 9 2 2
17 0 13 0 2 15 0 13 13 2 13 3 3 2 7 3 3 2
11 13 13 3 13 9 16 15 13 3 10 9
3 9 13 3
10 9 13 9 13 9 9 0 9 9 2
11 9 1 13 9 1 0 9 9 7 9 2
10 9 13 13 9 2 9 7 15 3 2
9 3 13 9 7 9 7 3 15 2
12 16 0 13 9 3 2 9 13 13 3 0 2
7 9 9 13 3 3 9 2
10 16 15 13 13 3 2 13 9 9 2
5 9 13 9 13 13
13 9 13 13 13 3 10 9 2 16 9 13 9 2
5 3 9 1 9 2
9 11 13 13 3 7 13 9 3 2
10 16 13 0 9 2 13 13 15 13 2
3 10 0 9
13 3 13 15 13 9 2 7 3 13 9 13 9 2
4 11 11 0 9
4 9 13 3 0
12 11 13 0 0 9 7 9 9 0 9 0 2
15 9 9 13 9 13 9 9 9 7 9 3 9 9 1 2
9 7 3 13 15 3 13 15 1 2
7 15 13 3 3 0 9 2
4 15 13 12 9
5 15 13 9 1 2
12 9 3 9 13 9 13 3 9 7 9 9 2
15 9 11 13 2 11 9 2 2 15 13 3 3 13 9 2
10 3 9 13 13 3 10 0 0 9 2
2 13 13
3 13 9 1
5 7 15 11 13 2
13 13 11 13 13 9 3 9 12 2 12 9 1 2
12 15 13 13 0 9 3 9 2 3 9 9 2
20 3 10 0 9 13 13 3 9 9 7 9 13 7 9 2 9 7 9 0 2
8 10 9 13 15 13 0 9 2
17 15 13 3 9 2 15 13 3 12 9 2 15 3 12 13 0 2
10 3 2 13 13 9 1 9 2 15 2
5 9 13 0 13 9
12 3 13 3 3 3 15 2 15 13 13 11 2
9 15 13 3 9 2 13 9 12 2
2 0 13
13 9 7 15 13 9 2 16 9 13 13 13 13 2
12 9 9 0 9 13 15 9 3 12 9 1 2
6 3 15 13 11 11 2
16 9 2 13 15 3 15 13 10 9 2 13 15 13 3 15 2
11 9 12 11 9 13 13 7 13 9 11 2
8 10 15 13 13 9 0 9 2
16 11 13 2 13 2 13 7 13 0 9 2 15 13 9 13 2
9 0 9 13 3 13 15 0 9 2
19 15 1 15 13 2 16 13 3 10 9 15 1 9 13 7 15 15 13 2
6 10 9 13 13 0 2
5 13 15 9 9 2
2 3 3
7 15 13 13 9 1 9 2
16 13 13 15 0 15 13 3 13 13 9 2 15 13 13 0 2
5 13 13 0 9 2
2 0 9
11 15 15 13 13 9 1 3 13 3 9 2
8 9 9 13 7 9 13 9 2
9 3 10 9 13 10 9 13 9 2
3 13 6 2
10 13 3 9 13 9 7 3 3 13 2
11 15 13 13 13 15 2 3 13 0 0 2
6 9 0 9 13 9 2
2 10 9
9 11 11 13 1 15 0 9 9 2
5 3 13 3 9 2
4 13 13 3 2
20 13 3 0 2 16 9 3 13 0 9 15 2 10 10 9 3 13 13 3 2
15 3 0 9 13 13 9 2 7 0 8 2 8 2 9 2
7 9 7 9 13 0 9 2
2 15 13
6 9 13 9 9 1 2
8 9 9 13 3 3 3 3 2
6 2 15 15 3 13 2
5 8 7 11 9 9
3 11 13 2
13 12 9 9 9 13 9 2 15 3 3 13 13 2
3 13 13 2
10 15 3 13 2 16 13 0 13 3 2
5 13 0 9 1 2
6 9 13 3 7 3 2
3 13 15 13
7 3 13 9 3 9 7 9
8 9 13 3 3 13 1 9 2
3 9 13 13
8 9 13 3 3 9 9 9 2
8 13 15 15 3 13 13 13 2
9 15 13 13 3 16 15 13 13 2
6 15 15 15 3 13 2
8 9 9 13 13 12 1 12 2
12 13 9 3 13 10 9 10 9 13 7 13 2
4 15 13 15 3
11 3 10 9 13 2 16 13 2 13 9 2
16 11 8 9 13 13 3 9 16 9 13 13 13 3 15 13 2
11 7 13 13 9 9 2 16 15 13 15 2
11 0 2 0 11 13 9 13 3 11 1 2
9 11 13 11 9 9 9 9 9 2
7 0 9 13 3 9 9 2
10 3 3 2 3 3 13 13 10 9 2
8 0 9 13 3 3 9 1 2
3 9 9 9
23 16 11 7 15 13 13 9 11 7 11 9 12 2 10 9 13 13 0 16 15 13 3 2
5 9 9 7 9 9
9 9 13 13 9 7 3 3 3 2
13 9 2 13 15 13 2 2 13 11 0 9 3 2
10 11 12 9 13 13 9 11 9 9 2
5 9 13 3 0 9
17 11 13 9 9 3 0 2 16 15 13 13 3 16 3 3 13 2
3 15 13 11
14 9 9 13 0 9 9 9 2 15 13 9 10 9 2
6 15 13 3 13 11 2
9 3 9 13 9 1 3 0 0 2
8 11 13 3 13 13 0 9 2
9 15 13 9 2 16 13 0 9 2
15 13 15 3 0 9 2 7 13 2 13 15 3 0 9 2
5 9 13 9 9 2
12 3 9 13 0 9 2 15 13 9 7 9 2
15 0 9 0 9 13 13 7 13 16 13 12 9 13 13 2
8 13 3 3 13 9 13 9 2
13 15 13 15 2 13 9 7 13 2 13 3 9 2
2 13 9
9 13 3 3 2 9 11 7 9 2
7 13 9 13 9 13 13 2
10 7 16 13 2 3 3 7 10 9 2
5 13 10 9 11 2
8 9 1 15 13 13 9 0 9
8 9 9 7 9 13 0 9 2
17 13 3 10 9 2 3 15 13 9 13 9 2 16 15 13 15 2
3 9 0 9
14 13 15 3 3 0 9 9 13 9 13 12 9 9 2
9 15 13 10 9 13 15 2 7 2
4 9 13 3 2
6 15 13 15 13 0 2
6 13 9 13 3 3 2
2 13 3
9 3 9 2 16 13 9 2 7 2
16 13 3 2 16 9 13 0 9 7 3 3 3 13 9 9 2
12 11 13 13 0 9 2 7 15 13 0 9 2
4 15 13 9 1
7 13 13 13 9 13 9 2
6 3 11 9 11 13 2
5 9 13 9 13 2
11 11 13 15 0 9 2 16 15 15 13 2
10 0 9 1 9 13 3 0 7 0 2
8 9 7 15 13 9 13 0 2
4 9 13 11 2
5 15 1 13 0 2
11 9 13 9 9 13 9 9 3 0 9 2
23 13 13 13 9 15 2 15 13 2 16 15 13 15 2 16 15 13 0 9 7 0 9 2
9 3 16 15 13 3 3 0 13 2
12 3 0 9 9 13 3 3 9 0 9 9 2
3 13 15 2
2 13 3
5 15 1 13 13 2
5 15 13 10 9 2
6 9 2 10 9 0 2
4 9 13 3 2
11 11 3 13 11 13 3 10 9 11 9 2
10 11 11 12 0 9 13 3 13 9 2
2 13 9
3 13 13 13
12 9 13 13 9 9 2 9 2 9 7 9 2
17 10 9 13 13 13 0 2 7 9 7 1 10 9 13 13 0 2
2 13 11
18 9 13 9 9 2 7 13 15 13 0 9 9 7 13 15 0 9 2
5 13 9 13 9 2
11 11 13 13 12 9 3 16 13 11 13 11
9 9 13 9 13 3 8 7 9 2
3 3 3 16
5 13 3 0 9 3
15 6 10 0 2 0 7 9 13 2 0 12 3 0 9 2
14 9 9 13 13 10 9 2 16 9 13 13 9 1 2
10 7 10 9 15 13 2 3 7 9 2
6 13 3 3 0 9 2
6 0 9 9 13 9 2
15 15 3 3 13 13 2 16 13 10 0 16 9 13 3 2
15 9 13 0 9 13 13 10 9 13 3 10 9 0 9 2
14 9 11 9 7 12 9 13 13 9 7 11 9 9 2
7 0 9 3 13 0 9 2
17 9 9 13 13 13 0 2 3 16 13 0 7 9 2 13 11 2
15 9 13 13 9 15 2 16 15 3 3 13 9 7 9 2
6 15 13 15 3 3 2
10 9 13 9 2 16 15 13 13 9 9
3 0 3 13
5 9 13 9 1 2
20 16 9 13 13 9 2 15 13 15 12 9 9 2 16 13 15 2 9 9 2
11 3 15 13 13 2 16 0 9 13 13 2
3 9 13 2
4 9 15 13 13
8 11 13 13 15 7 13 13 2
6 9 9 13 3 0 2
3 9 13 9
2 0 13
4 13 0 9 9
6 13 3 3 3 3 2
2 10 0
4 9 13 0 13
5 13 9 12 9 2
10 9 13 9 9 11 1 9 3 1 2
6 3 13 9 13 9 2
9 13 3 9 2 16 13 15 13 2
8 15 13 3 3 0 9 13 2
3 13 9 11
6 13 15 3 3 9 2
5 11 1 13 9 2
19 3 13 15 2 16 13 1 9 13 15 9 3 2 3 15 13 13 3 2
4 13 9 9 2
6 3 10 3 15 13 2
10 0 15 1 13 2 16 9 9 13 2
5 3 13 3 9 2
9 10 9 0 9 0 13 9 9 2
11 3 1 9 15 13 12 0 9 13 9 2
16 12 9 1 11 13 8 8 8 13 0 9 1 0 9 9 2
13 3 10 9 13 9 9 2 3 15 13 9 9 2
7 11 7 9 13 9 9 2
5 0 9 7 9 2
15 3 3 9 13 13 9 16 0 3 13 9 13 0 9 2
13 13 13 3 16 13 3 10 0 13 2 11 13 2
4 13 13 13 2
11 15 13 11 0 9 2 7 15 13 3 2
3 13 9 1
11 11 13 3 3 16 13 3 10 11 9 2
10 9 3 0 9 13 9 12 11 9 2
4 3 13 0 2
9 13 15 3 0 7 3 15 13 2
2 13 13
6 9 13 9 9 9 2
11 15 13 3 10 10 9 2 7 9 13 2
2 0 9
12 9 13 9 12 0 9 7 11 13 0 9 2
18 3 13 13 13 0 15 2 16 9 13 3 15 2 10 9 3 13 2
3 9 13 9
11 13 15 3 13 11 2 13 3 0 9 2
11 0 9 13 13 9 3 0 9 16 0 2
26 15 1 13 0 9 10 9 3 15 13 3 2 3 15 3 3 13 2 15 13 15 9 7 10 0 2
13 13 15 13 9 2 7 13 15 15 9 10 9 2
4 9 15 13 2
11 9 9 13 13 2 16 10 9 13 9 2
7 10 9 13 15 13 0 2
4 13 9 12 1
15 3 13 13 10 10 9 2 15 9 13 9 16 13 13 2
7 3 15 13 13 9 9 2
7 3 15 3 13 9 9 2
2 0 9
7 9 13 13 12 9 1 2
23 11 9 13 13 0 9 7 9 9 11 2 3 16 9 9 0 9 13 9 7 9 1 2
13 11 2 11 7 11 13 3 2 7 9 3 0 2
5 9 13 3 9 2
2 13 0
10 11 13 13 0 9 13 0 9 0 9
12 16 9 13 0 9 2 13 3 13 13 9 2
9 11 13 3 10 9 2 11 12 2
5 3 9 7 9 2
16 3 16 15 3 13 3 3 2 16 15 13 3 9 13 16 2
7 9 13 10 9 7 9 2
3 0 9 9
3 9 13 13
10 0 9 9 13 3 2 3 7 3 2
3 9 13 3
6 10 9 13 3 12 2
9 9 13 13 3 9 1 0 9 2
5 7 10 0 0 2
2 0 9
7 10 9 13 3 0 9 2
8 13 0 13 2 15 13 3 2
17 9 2 9 7 9 13 9 2 15 1 9 10 9 13 3 0 2
5 13 15 13 9 2
2 6 2
4 15 15 13 2
4 3 13 13 2
5 9 13 9 1 2
4 0 9 13 2
21 10 12 9 1 2 16 15 13 13 3 2 13 3 15 12 9 13 2 15 3 2
18 3 9 3 10 9 13 9 13 3 2 16 13 13 3 16 10 0 2
7 11 9 13 13 9 12 2
6 15 13 16 11 11 2
8 15 15 13 9 2 13 0 2
6 15 13 3 3 9 2
4 9 13 3 2
3 13 13 2
12 9 0 7 9 3 0 9 13 3 10 9 13
2 13 9
6 0 9 13 13 9 2
12 13 3 13 15 7 15 3 2 16 9 13 2
10 9 13 13 3 3 0 9 2 16 3
3 11 13 13
11 9 13 13 9 1 0 2 15 15 13 2
3 9 9 13
7 11 13 13 9 1 0 9
13 12 0 9 13 13 11 1 7 15 13 13 3 2
7 3 9 13 13 13 13 2
3 0 9 9
9 13 13 0 9 13 9 2 13 2
7 9 9 9 13 9 12 2
5 9 13 0 9 2
5 10 9 9 13 2
5 15 13 1 9 2
4 15 13 0 13
14 15 13 3 2 16 13 15 13 13 11 7 11 9 2
6 9 13 13 9 9 2
10 15 13 9 13 13 0 9 10 9 2
7 16 13 0 2 13 0 13
7 13 3 3 3 3 9 2
5 9 9 13 3 9
5 9 13 12 9 2
9 9 9 13 13 15 3 0 9 2
2 0 0
4 13 9 3 9
7 9 13 13 0 0 9 2
9 9 13 13 9 16 9 13 9 2
7 9 11 13 9 11 9 2
10 9 13 13 13 2 16 13 13 9 2
5 13 15 15 3 2
3 10 9 9
9 11 9 9 13 9 12 9 1 2
9 13 3 9 2 15 13 15 13 2
4 0 13 13 2
6 11 7 11 13 9 2
7 9 9 13 9 0 9 2
11 9 9 13 9 11 2 11 2 11 7 11
3 15 13 13
5 13 13 3 3 2
4 9 13 9 3
6 9 13 3 13 9 2
3 15 13 3
13 13 3 3 0 2 10 9 1 9 13 9 13 2
7 15 13 0 9 1 9 2
15 16 11 13 3 3 13 9 2 13 0 9 13 13 13 2
14 10 9 16 15 13 3 2 15 13 3 13 10 9 2
4 15 13 13 2
9 11 9 13 13 10 0 9 11 1
11 13 3 15 15 2 16 13 0 9 1 2
11 0 13 13 0 12 9 9 9 11 9 2
11 0 9 9 13 0 9 9 1 0 9 2
10 11 13 9 1 3 10 9 0 9 2
3 9 13 2
6 9 9 13 9 1 2
6 9 13 13 13 9 2
5 15 13 13 9 2
7 15 13 11 9 3 3 2
13 2 6 2 15 13 13 3 2 7 3 3 13 2
11 13 0 2 3 0 2 15 13 3 3 2
30 15 13 9 13 3 16 15 13 13 9 11 2 1 11 7 3 13 10 12 9 11 2 3 15 9 13 9 9 9 2
5 7 15 13 3 2
9 10 9 13 13 12 9 11 1 2
7 9 9 9 13 11 9 2
17 0 9 13 3 3 0 9 2 15 0 9 1 3 13 13 9 2
14 16 15 13 3 9 2 13 3 10 9 2 11 13 2
15 10 9 7 9 1 2 0 7 0 2 9 13 9 9 2
11 10 13 9 13 13 9 0 2 0 9 2
10 11 7 11 9 13 11 2 11 11 2
6 9 1 13 0 9 2
4 0 9 13 13
10 10 9 9 9 13 3 3 9 9 2
6 13 13 9 7 9 2
5 15 13 9 9 2
5 9 13 9 9 9
2 13 9
10 9 13 3 2 16 16 13 3 13 2
8 0 9 13 3 9 7 13 3
6 13 9 9 1 9 2
5 9 9 13 0 2
4 13 16 13 2
7 13 16 11 13 13 9 2
13 15 13 15 2 16 9 9 13 11 0 16 11 2
10 10 9 13 13 3 13 0 9 9 2
5 11 13 9 13 9
8 9 9 13 9 13 12 9 2
12 13 15 10 9 10 9 13 7 13 13 15 2
22 16 10 9 13 2 16 13 13 9 7 3 13 3 13 9 2 9 13 9 13 9 2
4 11 9 13 2
12 11 9 13 13 9 2 3 10 9 13 9 2
3 9 0 9
11 3 9 13 9 3 3 10 9 0 9 2
7 9 13 1 9 7 9 2
6 10 9 15 3 13 2
17 0 9 0 9 1 13 0 12 9 7 15 13 13 3 12 9 2
18 16 11 13 0 9 2 9 13 9 2 16 9 1 9 13 13 3 2
30 3 9 3 13 2 8 13 9 9 7 2 13 3 3 3 2 13 2 13 3 0 2 0 9 7 13 9 15 7 2
6 11 13 11 9 1 2
6 9 15 13 0 9 2
4 3 3 15 2
7 9 13 3 9 0 9 2
7 13 0 15 2 16 13 3
7 11 7 9 13 3 9 2
11 0 7 0 13 0 11 7 11 13 9 2
2 10 9
22 7 15 9 13 13 3 0 13 13 3 9 13 13 2 16 13 3 3 1 10 9 2
9 13 3 7 3 3 13 0 9 2
15 10 10 9 3 13 15 3 16 15 13 3 12 9 9 2
24 9 13 2 13 0 9 13 9 2 7 13 15 0 9 2 15 11 13 13 3 3 12 12 2
9 15 13 3 7 15 13 0 9 2
4 13 9 3 2
4 9 13 9 2
6 9 13 13 9 9 2
2 9 9
7 7 15 13 13 0 9 2
7 9 13 3 16 13 9 0
13 3 0 2 3 9 2 13 13 3 0 2 0 2
9 9 13 9 13 9 13 9 1 2
12 15 13 3 3 7 13 9 13 9 3 3 2
8 2 6 2 11 15 15 13 2
14 11 13 7 13 12 0 9 2 9 7 9 0 9 2
6 15 15 13 3 3 2
2 9 9
9 13 13 9 9 2 0 9 9 2
9 11 9 13 9 3 16 11 9 2
3 8 7 9
14 15 3 13 9 7 12 2 7 15 13 13 9 9 2
4 15 13 12 9
6 13 15 9 15 13 2
16 3 15 3 13 16 13 10 9 15 13 16 3 12 9 13 2
7 11 13 0 9 1 9 2
6 9 9 13 9 13 13
18 15 13 2 16 13 9 13 3 3 9 2 16 13 3 12 9 0 2
6 13 16 11 13 11 2
4 0 9 9 9
14 16 15 13 9 9 2 13 9 13 10 13 0 9 2
7 11 13 3 9 9 12 2
9 13 3 13 3 0 16 3 9 2
14 9 16 13 2 13 7 3 0 9 13 9 9 1 2
9 13 15 9 7 13 15 13 9 2
11 3 13 15 13 9 9 1 7 3 9 2
8 9 9 13 13 7 13 3 2
13 15 13 13 0 0 9 3 3 10 0 9 1 2
9 9 1 11 13 13 0 0 9 2
17 13 11 13 3 9 2 3 15 13 3 3 12 12 9 0 9 2
12 3 15 1 13 9 2 16 15 13 13 9 2
11 13 3 15 7 9 7 9 2 3 9 2
2 3 13
8 15 1 9 3 13 11 9 2
13 3 11 11 11 0 9 10 9 13 3 10 9 2
12 15 13 12 9 0 9 2 16 15 13 9 2
16 10 9 15 15 13 13 3 3 3 15 13 15 10 9 0 2
16 3 16 15 13 10 9 10 9 3 3 13 3 9 13 9 2
6 9 13 13 3 9 2
4 9 13 9 11
12 13 15 3 3 13 13 10 9 16 15 13 2
17 11 7 11 9 7 9 9 11 9 7 11 1 13 11 0 9 2
9 9 0 13 9 3 13 9 9 2
6 9 13 3 13 13 2
6 13 9 2 15 13 0
13 11 9 13 10 9 16 9 2 9 13 0 9 2
12 7 9 13 13 0 2 16 3 3 13 13 2
5 9 13 0 9 2
10 10 9 9 13 13 2 9 7 9 2
6 9 13 15 0 0 2
15 9 13 9 11 11 2 9 2 9 13 13 3 9 9 2
7 15 13 13 15 10 10 9
5 0 3 13 9 2
17 3 15 13 0 9 2 15 13 13 1 9 9 13 9 3 15 2
5 15 13 11 9 9
4 15 13 13 2
21 16 3 9 13 3 7 0 9 13 13 0 9 1 2 15 13 13 9 2 16 2
8 2 13 3 2 15 13 13 2
11 11 0 9 9 9 13 9 13 3 12 2
4 10 9 0 9
3 10 9 2
6 13 13 3 3 9 2
10 9 7 9 0 9 13 3 13 13 2
13 10 15 13 13 10 9 2 15 15 3 3 9 2
12 11 0 9 11 3 11 13 13 9 0 1 2
14 15 13 9 9 7 13 11 2 13 15 3 13 15 2
12 11 1 9 13 13 15 3 0 13 0 9 2
6 3 13 13 0 9 2
8 13 11 9 16 13 9 13 2
12 3 10 11 13 6 3 9 16 13 9 3 2
6 11 11 13 10 9 2
10 16 13 3 13 2 3 13 13 13 3
7 3 13 13 9 11 3 2
8 9 15 13 13 13 2 7 2
3 15 13 9
5 0 11 13 3 2
14 15 13 2 16 9 13 12 13 9 15 9 16 9 2
7 15 13 13 9 3 3 2
2 15 1
3 11 13 13
3 10 0 9
8 10 9 13 13 12 13 9 2
15 3 10 9 13 13 15 2 16 13 13 13 10 9 13 2
3 9 13 13
5 15 13 13 13 2
5 15 13 13 3 2
3 9 13 2
4 9 9 13 3
12 0 11 15 13 13 2 16 13 13 0 9 2
14 9 13 10 9 9 13 2 7 13 9 9 0 13 2
2 10 3
17 9 13 3 9 2 15 9 13 13 9 15 15 10 9 16 15 2
4 10 9 13 0
16 3 13 13 3 2 15 1 2 9 2 13 3 3 3 13 2
6 9 13 3 12 9 2
9 13 3 13 9 3 16 10 15 2
12 10 9 13 13 9 2 7 15 13 3 13 2
7 9 13 0 9 9 13 2
10 13 13 7 13 3 9 2 3 9 2
13 2 16 13 2 3 13 3 3 3 13 3 0 2
5 13 9 0 9 2
12 15 13 13 10 0 9 2 7 3 13 11 2
3 13 3 2
6 9 13 9 3 3 2
7 13 3 9 0 0 9 2
5 13 3 16 9 2
14 12 9 13 9 3 9 1 9 2 12 9 3 9 2
10 3 9 1 13 15 0 16 0 9 2
2 0 9
3 3 0 9
6 13 9 3 12 9 2
2 9 9
9 3 0 13 13 11 11 9 1 2
9 9 7 9 13 11 12 9 9 2
6 9 13 13 3 16 13
11 9 13 15 2 15 3 9 13 12 9 2
3 9 12 9
6 9 9 9 13 13 2
16 15 13 0 9 16 3 13 9 11 16 15 13 13 10 9 2
6 15 13 3 0 9 2
4 3 13 9 2
3 13 13 2
2 13 3
4 9 13 12 9
8 15 13 9 3 15 1 9 2
10 9 13 9 9 9 7 15 1 9 2
6 0 9 13 0 9 2
14 15 13 3 1 9 2 16 13 10 9 7 13 13 2
8 7 11 9 13 0 16 9 2
16 6 2 9 3 3 2 7 0 9 13 3 13 10 9 13 2
13 10 9 9 13 13 11 2 16 15 13 0 9 2
2 6 9
18 9 11 11 1 3 9 13 9 13 3 13 10 9 13 9 13 9 2
10 11 9 13 9 13 9 7 13 9 2
15 15 1 15 13 3 13 2 16 13 3 3 7 15 3 2
9 9 13 13 3 9 16 13 9 2
4 7 9 7 9
16 15 13 13 9 2 15 0 7 9 3 13 9 13 13 13 2
7 2 9 2 2 13 11 2
5 3 13 2 13 9
11 3 10 9 7 9 13 9 3 9 1 2
8 11 9 9 9 9 13 9 2
12 10 9 13 10 9 12 9 1 3 7 3 2
7 11 13 13 9 9 9 2
4 11 13 15 13
2 10 9
8 0 7 13 2 7 9 13 2
18 9 13 2 16 9 13 9 9 1 2 3 9 13 13 3 1 9 2
6 3 11 13 13 9 2
9 9 13 9 0 13 10 9 9 2
9 9 13 13 13 12 9 10 9 2
8 15 13 2 16 9 13 0 2
5 9 13 9 1 2
11 13 9 13 7 9 13 13 16 13 3 2
11 11 13 0 9 7 13 9 1 0 9 2
4 9 13 9 1
8 11 13 10 9 9 0 9 2
10 9 13 12 9 13 13 11 9 9 2
17 10 9 13 13 15 2 13 9 7 13 9 0 0 9 9 9 2
12 0 0 2 15 13 13 9 2 16 13 13 2
4 15 13 0 2
6 11 9 7 9 13 9
5 13 3 10 9 2
7 3 13 3 13 10 9 2
2 9 13
6 11 13 15 3 0 2
5 9 13 13 9 2
7 13 3 13 13 3 9 2
7 3 11 13 9 9 3 2
14 3 13 9 9 7 9 13 2 16 13 9 9 9 2
15 3 13 9 13 0 3 2 16 13 15 13 13 0 9 2
10 9 13 9 7 13 9 9 9 9 2
6 11 13 3 0 9 2
10 10 9 15 13 9 1 15 13 13 2
11 11 13 3 12 0 9 7 15 13 11 2
12 16 9 13 3 2 11 3 13 15 0 9 2
23 9 13 16 3 13 9 2 7 9 2 15 13 13 3 13 9 7 15 3 13 11 9 2
6 13 15 0 7 0 9
11 15 13 0 9 2 16 13 9 3 0 2
19 13 9 13 9 9 7 13 7 13 9 1 7 3 3 3 3 3 9 2
7 10 9 11 11 13 3 2
7 9 13 12 9 0 9 2
14 0 9 13 2 3 13 9 2 16 15 13 13 9 1
11 7 13 9 13 13 11 0 9 13 15 2
17 9 9 13 9 1 3 10 9 13 13 2 3 16 15 13 13 2
6 15 15 3 3 13 2
3 13 13 3
6 15 13 15 3 0 9
7 9 13 15 13 3 9 2
6 9 12 7 13 9 2
13 0 9 13 13 12 9 9 2 16 13 9 13 2
7 10 9 13 9 1 0 2
3 13 3 2
4 15 15 13 2
8 13 3 13 13 3 0 10 9
15 9 13 13 10 0 16 16 13 3 2 15 9 13 13 2
11 13 0 9 3 2 16 13 0 7 0 2
16 6 15 3 13 15 13 3 7 0 9 3 3 12 3 12 2
11 11 13 9 1 3 9 16 3 3 9 2
15 11 11 13 0 2 0 9 13 9 11 9 9 12 9 2
6 15 1 10 9 13 2
6 7 3 15 13 9 2
16 9 1 13 3 13 13 3 2 15 13 13 13 3 0 9 2
3 9 13 13
10 9 9 1 9 13 13 9 0 9 2
12 13 3 9 3 10 9 16 15 13 9 9 2
2 9 9
5 9 13 3 3 2
4 9 13 9 9
7 10 9 13 0 16 10 9
5 3 3 13 13 2
11 9 13 9 2 15 13 3 9 9 1 2
5 9 9 13 9 2
6 13 13 16 15 13 2
8 11 13 13 10 12 3 0 2
5 11 3 13 11 9
13 9 13 3 9 2 13 9 7 13 9 9 9 2
7 9 1 9 13 9 13 2
3 0 13 9
3 13 9 3
11 7 15 13 0 3 7 3 15 13 3 2
5 13 3 2 11 2
19 15 7 9 13 10 9 1 3 3 3 9 2 13 9 9 11 2 12 2
12 9 13 3 3 9 12 9 13 9 9 11 2
15 13 15 13 0 9 0 2 2 11 13 9 15 13 9 2
10 3 13 13 9 16 11 10 3 13 2
7 9 13 11 9 10 3 2
8 10 9 13 9 13 0 9 2
7 15 13 9 12 9 11 2
10 15 2 16 15 13 0 2 13 13 9
8 13 11 3 7 11 3 3 2
9 13 2 16 9 13 15 9 9 2
3 9 13 13
9 15 13 3 13 9 11 9 9 2
5 13 3 9 9 2
8 15 13 3 13 12 0 9 2
5 15 13 9 1 2
6 15 13 3 12 1 2
10 9 13 10 0 9 2 3 3 3 2
4 15 13 3 3
11 16 9 13 13 9 2 15 15 13 13 2
6 9 2 9 15 13 2
3 2 9 2
8 0 9 7 9 13 9 9 2
5 9 13 13 9 2
18 16 0 9 13 13 16 13 9 13 2 3 3 13 15 13 0 9 2
12 3 9 1 13 2 9 13 9 9 9 1 2
4 11 13 9 2
12 3 11 11 9 13 9 13 3 3 9 9 2
12 15 13 10 0 16 13 13 9 2 15 13 2
9 11 7 9 3 9 13 9 9 9
16 9 11 13 0 0 9 2 11 9 2 7 15 13 15 9 2
8 11 13 13 3 7 13 13 2
10 9 0 9 13 11 13 2 3 9 2
7 3 3 3 13 9 9 2
9 9 13 3 3 2 0 2 9 2
9 9 13 3 9 0 16 9 1 2
5 10 9 15 13 2
7 11 9 13 9 13 1 2
3 9 0 2
6 0 9 13 9 9 2
3 0 13 0
21 3 15 13 13 2 16 13 2 16 9 13 9 3 13 9 7 13 9 13 9 2
9 15 15 13 13 2 13 13 9 2
7 3 15 13 2 13 9 9
2 9 9
11 9 13 13 0 12 9 1 11 13 9 2
2 10 9
9 3 15 13 13 0 9 9 13 2
10 11 13 9 9 0 0 9 13 9 2
6 0 9 13 13 9 2
4 9 9 13 9
8 9 13 13 3 12 9 9 2
15 11 9 13 3 9 9 2 11 9 13 13 3 0 9 2
5 15 13 12 3 12
10 15 13 3 0 7 15 13 10 9 2
11 0 9 9 13 9 13 9 13 3 3 2
5 15 13 3 0 2
7 9 13 3 9 9 9 2
12 11 13 9 9 2 13 15 0 0 0 9 2
12 13 13 11 2 11 2 11 2 11 7 11 2
8 11 13 10 9 12 11 9 2
8 9 13 13 12 9 12 9 2
7 9 1 13 13 3 9 2
10 9 13 9 2 16 11 9 13 9 2
5 10 9 13 9 2
6 9 13 3 12 9 2
5 13 15 0 9 2
6 10 9 13 3 0 2
14 11 13 3 9 2 16 13 9 13 3 0 0 9 2
6 3 15 10 9 13 2
7 11 11 13 12 9 9 2
15 3 13 3 13 0 9 7 9 3 7 9 7 9 3 2
7 8 8 3 13 13 9 2
10 0 0 9 13 3 3 10 12 9 0
5 15 3 9 13 2
19 15 13 9 2 3 16 13 13 15 3 15 3 13 0 9 10 9 1 2
17 16 13 13 15 2 3 3 13 15 2 3 0 9 9 13 9 2
3 10 10 11
5 15 13 3 0 2
10 9 9 13 15 13 2 16 3 13 2
8 13 13 2 3 13 0 11 2
6 3 15 13 13 9 2
10 15 13 13 0 9 0 0 10 9 2
13 9 9 13 13 3 2 16 9 13 13 3 9 2
15 15 13 2 16 13 15 13 0 0 15 1 7 11 1 2
10 15 13 15 13 3 2 15 3 12 9
7 9 9 13 9 3 9 2
10 15 13 9 2 16 15 13 13 9 2
10 13 15 15 2 13 3 3 3 9 2
7 13 9 9 2 13 9 2
15 16 13 13 9 2 13 3 16 15 13 13 7 13 0 2
8 9 15 9 13 15 9 13 2
14 9 13 9 1 2 3 1 0 9 7 0 9 9 2
6 2 9 13 3 13 2
6 7 13 15 13 9 2
8 9 13 9 13 3 0 9 2
5 13 15 13 10 9
5 9 11 7 11 2
9 0 9 13 9 2 3 13 13 2
5 15 13 13 9 2
4 9 13 9 1
6 9 9 13 9 9 3
9 3 1 0 9 13 11 11 11 2
4 2 10 9 2
7 15 13 3 13 13 9 2
7 9 13 13 2 13 7 13
5 9 13 9 9 2
14 9 9 7 9 13 13 15 2 16 15 13 13 9 2
13 10 9 13 3 13 2 16 0 9 13 15 13 2
4 9 13 13 9
15 15 13 10 0 9 2 16 9 13 0 0 2 12 9 2
9 3 13 2 16 15 13 13 13 2
15 13 0 13 2 16 10 9 9 3 13 13 9 10 9 2
6 15 13 3 3 12 2
11 13 9 3 7 9 13 3 13 9 9 2
2 0 9
7 2 3 3 13 13 2 2
6 15 15 13 0 9 2
5 10 0 9 13 3
2 0 9
6 11 13 11 9 9 2
8 10 9 16 13 15 13 9 2
12 11 13 3 0 9 7 13 3 9 9 1 2
9 11 13 11 0 9 1 12 9 2
6 11 13 13 13 11 2
9 10 9 9 13 3 0 16 0 2
4 15 13 11 3
12 15 13 13 15 3 2 3 16 13 3 0 2
11 7 9 9 7 9 9 13 15 12 9 2
12 13 9 13 2 16 9 13 0 7 0 9 2
7 3 9 13 13 9 7 9
14 16 9 13 3 13 9 2 15 3 13 13 0 9 2
14 15 13 10 9 2 16 13 15 13 13 9 13 15 2
3 6 3 0
7 13 2 16 3 13 9 2
9 9 11 13 13 9 11 9 9 2
10 15 13 2 16 15 13 11 0 9 2
9 13 13 3 2 13 15 15 13 2
9 9 1 9 1 13 3 12 9 2
9 10 0 9 13 0 12 9 9 2
11 15 13 2 16 10 9 13 13 10 9 2
8 3 9 13 11 12 0 9 2
5 0 16 10 15 2
2 9 2
8 9 11 13 12 9 9 12 2
22 0 9 2 11 2 11 2 11 2 15 2 13 3 3 0 9 2 13 9 0 9 2
10 13 3 3 12 9 7 16 9 13 0
5 15 13 9 9 2
8 13 15 2 16 13 9 9 2
5 15 13 13 9 2
11 13 13 9 10 9 2 13 15 3 13 2
8 9 1 13 9 9 0 9 2
6 9 11 13 13 15 2
10 13 9 13 2 2 13 15 9 2 2
5 9 13 9 9 2
11 9 1 13 0 9 13 3 3 13 9 2
6 9 13 13 12 9 2
3 13 9 2
15 9 10 12 13 9 12 9 2 3 16 15 13 10 9 2
11 9 13 2 16 13 15 13 3 12 9 2
5 15 13 0 13 2
10 13 13 13 9 7 9 13 15 13 2
6 9 13 15 3 1 2
2 13 9
13 9 0 9 13 9 3 3 2 15 13 3 13 9
7 15 13 3 12 11 9 2
3 9 13 9
16 11 12 9 0 9 9 13 13 0 9 7 9 9 12 9 2
12 9 9 13 3 0 2 7 13 15 9 13 2
8 9 9 2 13 7 13 13 2
21 13 13 16 10 9 16 13 16 0 9 13 9 2 13 15 0 15 2 13 9 2
6 9 13 9 13 9 2
2 13 13
3 9 13 2
8 9 13 9 7 10 9 1 2
10 9 13 13 9 9 3 3 16 9 2
6 0 15 13 13 13 2
10 9 9 11 13 13 0 2 7 0 2
10 9 13 9 9 13 2 13 9 9 2
12 9 3 15 13 13 9 15 1 2 12 9 2
8 15 13 0 9 0 0 9 2
10 9 13 3 9 2 16 13 9 13 2
4 15 15 13 2
16 16 13 9 13 12 9 1 9 13 9 9 1 3 3 13 2
17 11 13 13 9 9 13 10 0 0 9 9 0 3 9 9 9 2
14 11 11 13 13 9 10 9 1 7 13 3 0 9 2
11 15 13 3 3 16 10 9 13 12 9 2
4 9 13 9 11
4 13 9 9 2
4 0 15 13 2
6 9 13 13 13 9 2
2 9 13
6 0 9 9 13 13 2
5 15 13 3 0 2
9 9 13 13 3 0 9 13 15 2
8 11 13 3 13 0 1 13 9
14 0 9 13 2 15 13 13 2 7 13 15 9 13 2
3 15 13 3
4 13 9 9 2
4 9 2 0 2
6 9 13 7 9 9 2
16 13 13 13 9 7 9 2 3 13 3 15 7 13 0 9 2
18 13 16 13 13 15 16 16 11 13 9 0 9 15 13 3 13 13 2
5 9 15 13 12 2
17 9 13 9 9 2 9 13 13 0 0 9 7 3 0 9 13 2
6 9 13 3 13 9 2
11 1 11 11 3 0 13 13 3 3 9 2
2 0 1
5 9 13 3 9 2
11 15 13 10 9 9 2 16 15 13 3 2
2 0 9
4 13 13 9 2
11 15 13 15 3 16 15 13 13 15 13 2
8 16 9 13 9 2 13 9 2
3 13 9 2
14 10 11 13 13 9 2 7 3 15 13 13 0 9 2
4 13 15 9 2
7 3 0 9 9 13 9 2
11 9 13 10 9 11 1 0 9 9 11 2
2 13 13
7 0 10 9 3 13 9 2
2 0 9
7 13 3 0 13 12 12 2
11 13 9 10 9 1 2 15 15 15 13 2
7 13 10 0 3 3 3 2
3 13 3 2
7 7 3 13 3 3 9 2
3 3 13 2
8 9 13 3 0 16 9 13 2
7 9 9 13 9 9 12 2
7 3 11 13 9 0 9 2
6 9 13 13 0 9 2
10 10 9 13 0 2 7 13 3 0 2
10 13 9 0 9 9 1 3 13 9 2
11 15 13 13 13 9 13 0 2 0 9 2
3 11 15 2
4 13 15 9 2
9 0 9 15 13 2 13 10 9 2
8 15 1 15 13 13 3 9 2
5 9 13 12 9 2
6 13 2 16 15 13 2
11 15 13 3 7 3 13 7 9 13 3 2
7 13 3 9 9 1 1 2
13 13 13 3 16 13 9 7 13 13 3 16 13 2
18 0 9 13 11 9 13 11 9 2 15 3 12 13 9 13 9 9 2
3 0 16 15
5 9 9 1 9 13
32 11 3 13 3 15 3 13 16 15 13 13 10 9 15 16 15 13 13 3 13 10 9 7 15 13 3 0 3 3 13 15 2
7 9 13 9 13 0 9 2
11 15 13 11 9 7 9 0 12 9 1 2
14 10 9 13 13 13 2 16 10 9 13 3 0 9 9
3 12 0 9
7 0 9 9 9 13 13 2
4 13 9 9 2
33 10 15 3 3 3 3 3 13 16 15 3 3 13 16 9 13 9 3 15 2 6 15 16 0 9 15 13 7 6 15 13 15 2
13 0 9 13 9 13 2 9 15 3 9 1 13 2
4 15 13 9 2
21 13 3 16 9 9 13 13 9 2 7 15 13 13 3 13 11 11 3 0 0 2
7 11 13 13 9 3 1 2
13 9 13 0 0 2 9 13 15 9 13 9 9 2
9 10 9 15 13 13 2 10 9 2
3 13 9 0
5 13 15 13 13 2
2 10 9
7 9 13 9 0 9 13 9
6 10 9 13 13 9 2
31 15 13 3 16 15 13 13 2 13 15 1 16 13 13 16 13 7 3 13 2 13 15 1 16 15 13 3 3 7 3 2
16 15 13 3 2 16 9 13 13 9 12 0 9 15 10 9 2
12 11 15 13 3 3 3 13 9 10 9 9 2
15 9 13 9 0 0 9 2 0 9 2 3 15 13 15 2
6 3 9 13 3 9 2
6 13 9 7 13 9 2
4 11 13 3 9
9 9 13 13 13 2 15 9 13 2
5 9 13 3 9 2
2 13 9
16 9 12 9 13 13 15 2 15 3 13 10 9 10 9 1 2
6 13 15 13 3 6 2
11 9 9 13 9 7 15 1 13 0 9 2
9 9 9 1 15 13 3 0 9 2
8 9 13 9 2 7 3 9 2
31 15 13 3 9 1 16 15 13 9 15 13 3 3 3 16 15 3 13 16 6 6 16 9 15 13 12 9 9 13 9 2
14 3 11 13 3 13 13 9 3 3 3 16 15 13 2
9 10 10 9 9 13 12 9 9 2
14 13 16 13 13 3 3 10 12 9 2 7 13 9 2
7 0 11 9 13 0 9 2
16 9 9 0 0 9 13 3 0 9 2 13 9 9 15 3 2
17 9 13 9 9 7 12 9 9 13 13 3 9 9 7 11 9 2
3 11 13 3
15 15 13 13 10 9 2 7 11 1 15 13 3 3 13 2
12 15 13 11 9 12 2 15 15 15 13 13 2
8 11 1 9 13 13 10 9 2
12 0 7 0 0 9 13 9 3 10 9 13 2
13 9 13 13 13 9 2 3 15 13 13 9 13 2
6 9 13 12 12 9 2
10 0 9 13 9 2 16 13 0 9 2
4 13 9 0 2
4 0 13 9 2
16 0 9 2 13 3 13 3 2 16 3 13 15 7 0 9 2
14 13 15 13 9 13 2 16 15 13 9 13 13 9 2
12 12 0 9 2 15 13 0 7 0 10 9 2
4 11 13 13 9
3 9 7 9
9 3 9 13 9 13 9 1 9 2
6 11 11 13 9 9 2
23 10 9 13 2 12 9 1 13 13 9 2 10 9 2 15 1 13 13 15 2 9 12 2
5 15 13 11 11 9
6 9 9 7 10 9 1
5 3 9 13 9 2
18 0 9 7 9 13 0 9 2 15 13 9 7 3 3 0 16 0 2
17 15 13 13 3 9 2 16 13 3 13 13 2 3 0 9 13 2
25 9 3 13 2 16 11 7 11 13 13 11 0 9 2 13 3 13 11 10 9 16 11 9 1 2
5 13 9 0 0 9
6 13 15 13 3 9 2
4 13 15 13 2
15 16 9 13 3 7 13 9 2 9 13 7 13 3 9 2
16 11 13 13 3 15 3 2 7 9 10 9 13 3 13 0 2
11 9 9 13 9 0 2 13 15 13 9 2
11 11 1 9 13 3 3 0 15 9 13 2
6 13 13 15 9 13 2
5 15 13 12 9 2
2 15 13
2 15 1
2 0 9
15 13 9 9 13 13 2 16 9 13 3 0 9 9 13 2
10 10 12 0 13 9 13 9 12 9 2
10 3 15 13 9 10 9 2 10 9 2
3 9 7 9
9 12 9 1 3 13 3 9 9 2
19 3 15 13 2 16 15 13 13 2 7 13 15 2 3 15 13 0 13 2
9 0 9 13 13 9 0 9 9 2
2 9 0
2 13 3
3 9 9 1
3 15 13 15
9 7 3 13 9 2 13 3 9 2
5 13 15 3 13 2
7 10 9 10 9 13 13 2
4 9 0 9 2
11 15 13 15 2 3 9 9 13 0 3 2
8 11 11 13 3 0 0 9 2
5 9 13 13 3 13
10 13 3 12 9 2 3 13 13 9 2
11 9 1 13 9 3 13 9 7 10 10 9
3 9 3 2
2 13 0
5 13 16 15 13 2
2 9 3
15 3 9 1 13 13 2 3 9 0 9 13 3 12 9 2
6 15 13 3 9 1 3
4 13 13 9 2
9 11 13 12 9 3 3 11 9 11
3 13 13 2
6 11 13 3 13 0 2
4 0 7 13 2
2 0 11
14 9 9 13 3 9 15 13 9 2 7 15 13 3 2
5 15 13 9 13 2
8 13 3 13 16 15 13 3 3
13 9 1 9 13 9 0 2 9 0 7 13 0 2
8 2 0 0 9 13 12 9 2
10 13 15 10 0 13 2 9 11 13 2
7 9 9 11 9 3 13 2
2 9 13
12 16 9 13 2 9 13 16 3 9 3 13 2
6 13 9 9 9 1 2
2 0 11
18 15 13 13 9 10 9 7 10 9 3 7 9 9 11 13 3 0 2
15 15 13 0 7 0 9 2 7 12 9 3 13 13 3 2
25 9 2 9 2 9 2 9 7 9 9 13 11 3 12 10 9 2 15 1 9 9 13 9 11 2
8 9 13 3 0 2 0 9 2
2 0 9
3 13 9 9
13 13 15 3 3 0 13 2 16 13 9 9 9 13
2 11 0
5 15 13 9 3 2
2 9 9
9 11 3 13 3 0 13 13 9 2
6 15 13 3 13 3 2
6 9 13 12 3 12 2
4 9 13 3 2
6 13 9 9 12 1 2
7 11 13 3 13 11 9 1
6 11 9 13 0 9 2
15 9 9 2 3 15 13 13 3 3 13 2 13 9 9 2
6 9 13 11 13 13 2
6 7 3 13 3 13 2
5 13 15 3 3 2
9 13 9 2 3 9 3 9 9 2
5 13 0 9 9 2
6 9 13 13 3 9 2
7 9 13 13 3 0 3 2
5 13 3 3 9 2
8 9 11 11 13 12 9 9 2
4 15 13 9 2
9 10 9 9 15 13 9 2 16 2
2 10 9
8 10 9 13 11 9 9 12 2
17 11 13 13 11 9 0 9 1 13 9 13 13 12 9 9 9 2
6 1 9 2 7 9 2
4 15 13 9 2
11 10 9 16 9 13 2 15 13 10 9 2
12 3 13 10 9 2 16 3 3 9 13 3 2
6 15 13 13 10 13 2
8 9 13 3 12 9 12 9 2
14 9 13 0 9 13 2 16 13 13 13 3 9 9 2
4 13 13 9 2
14 13 13 7 3 11 11 0 9 2 15 9 13 3 2
5 15 13 9 3 2
7 13 13 9 13 3 9 2
10 10 9 13 3 12 13 11 11 11 2
8 9 13 11 2 11 7 11 2
12 9 13 7 13 9 0 9 0 9 13 9 2
1 12
7 9 13 9 13 9 9 2
6 9 13 9 13 0 2
8 9 9 13 3 3 16 0 2
6 9 13 0 10 9 2
2 9 9
9 15 13 3 0 2 13 7 13 2
5 9 13 12 3 12
14 15 13 9 9 7 13 3 9 7 13 2 16 13 2
7 15 13 13 13 13 9 2
3 9 9 2
5 10 9 15 13 3
6 9 13 13 13 9 2
8 3 15 13 12 13 11 3 2
7 13 15 3 15 3 0 2
12 11 13 13 3 13 7 13 3 0 7 15 2
7 9 13 7 3 3 9 2
5 13 10 15 3 2
6 15 13 13 0 9 2
10 9 13 13 9 2 16 13 15 13 3
4 2 13 15 2
5 10 9 3 13 15
12 10 9 13 0 9 2 13 0 7 13 0 2
5 13 15 15 13 2
6 15 13 0 10 9 2
5 13 9 7 13 2
11 0 9 1 0 9 9 9 13 13 9 2
5 0 13 3 9 2
8 3 15 9 1 9 13 15 2
19 0 9 1 13 11 0 9 2 0 11 9 9 11 11 9 0 9 9 2
11 13 9 9 7 13 0 0 9 10 9 2
5 9 13 9 13 9
6 15 0 9 13 13 2
8 11 13 9 3 7 9 3 2
14 13 13 2 16 10 0 9 13 13 13 0 12 9 2
7 3 0 9 13 9 15 2
4 13 12 9 2
7 11 11 13 3 0 9 2
2 9 1
7 15 13 13 9 7 9 2
6 16 15 13 10 11 2
7 13 9 13 13 11 9 2
9 13 9 9 13 10 0 7 0 2
7 13 9 9 3 13 9 2
5 9 13 10 9 2
7 0 9 13 13 15 9 2
11 9 13 13 9 2 10 9 13 13 9 2
15 10 9 9 2 9 7 9 13 9 13 13 13 13 9 2
12 11 9 13 15 9 2 15 15 3 13 11 2
5 13 15 3 9 2
4 13 3 9 2
9 13 2 9 9 2 2 9 13 2
9 11 9 13 9 11 0 9 9 2
5 15 13 13 9 2
4 13 12 1 2
10 15 13 3 0 9 2 15 13 9 2
10 15 13 0 9 16 13 2 9 1 2
6 9 13 13 13 9 2
4 0 13 0 2
9 9 13 0 16 15 13 9 1 2
14 11 13 13 9 9 7 13 13 3 13 10 9 15 2
9 3 13 9 2 13 11 13 9 2
6 3 9 13 9 0 2
3 9 3 2
11 10 9 13 3 0 15 15 2 11 13 2
7 9 13 9 7 9 13 2
13 10 9 15 13 3 0 2 16 9 13 9 9 2
11 6 6 2 3 15 3 13 2 9 13 2
4 15 13 0 2
5 9 13 9 3 2
11 12 9 12 9 13 3 13 13 3 11 2
3 13 10 9
18 9 13 0 2 9 0 7 0 2 9 0 2 1 7 1 12 9 2
10 15 13 15 7 15 13 0 13 9 9
2 10 9
15 11 13 9 13 13 9 9 13 9 0 9 13 9 1 2
16 3 15 3 13 13 2 16 13 9 13 10 12 9 3 9 2
6 9 11 13 11 9 2
5 13 9 13 9 2
8 0 9 10 10 9 13 13 2
19 6 15 10 9 2 3 11 9 13 2 13 7 13 13 11 1 0 9 2
3 9 13 13
9 3 16 15 13 3 3 13 12 12
5 15 15 13 13 2
8 3 16 15 13 3 3 15 13
6 9 13 10 9 9 2
15 15 13 9 9 2 7 15 11 13 9 13 9 0 9 2
10 9 3 9 2 9 3 7 0 9 2
6 0 9 13 12 9 2
5 9 13 13 0 13
11 13 3 13 3 9 0 9 12 9 9 2
11 11 13 13 2 13 15 0 0 13 9 2
7 11 13 9 2 12 2 2
4 11 13 9 2
2 13 3
5 13 13 3 13 2
15 0 9 13 9 9 7 13 12 0 11 2 11 7 11 2
7 13 13 10 12 9 13 2
13 15 1 9 13 0 9 9 9 3 12 12 9 2
12 11 7 10 9 13 13 9 10 9 9 1 2
4 9 13 3 9
4 11 13 11 2
6 11 13 9 3 13 2
16 11 1 10 11 9 9 7 12 10 9 13 11 9 9 9 2
13 9 13 13 9 3 10 9 2 16 11 13 13 2
5 9 13 11 9 2
7 9 9 9 13 12 9 2
8 9 13 13 0 0 2 3 2
7 15 13 13 10 9 3 2
18 3 9 1 9 13 9 9 11 13 3 9 9 11 9 9 9 9 2
6 0 9 13 9 9 2
7 9 13 13 0 12 9 2
13 11 13 0 9 9 2 16 10 9 13 9 9 2
11 11 13 9 9 7 13 15 13 9 9 2
5 13 13 10 9 13
9 16 13 0 13 10 9 13 9 2
13 16 15 13 3 0 9 2 13 13 9 3 9 2
19 13 9 13 2 16 15 13 9 9 2 7 13 13 13 2 16 15 13 2
14 15 13 13 9 2 7 13 15 9 13 7 0 9 2
13 9 10 9 13 13 9 2 3 0 13 11 9 2
6 3 9 1 9 13 0
8 0 10 9 13 10 3 13 2
7 11 9 13 3 3 9 2
8 3 13 13 13 9 13 9 2
26 16 3 11 9 3 13 13 13 15 15 13 3 3 15 3 3 13 3 15 15 3 13 10 0 9 2
2 13 13
9 9 13 9 13 13 11 0 9 2
3 13 13 3
7 13 9 9 9 7 13 2
3 9 10 9
3 2 13 2
8 13 0 16 9 13 13 3 2
4 15 13 13 2
2 10 9
14 11 13 3 0 9 2 16 0 0 9 13 9 9 2
6 9 13 3 15 3 13
8 3 0 9 16 9 13 13 2
6 9 13 9 13 0 2
2 13 0
9 15 13 0 9 7 3 0 9 2
22 10 0 9 2 3 9 2 13 3 13 3 12 9 9 0 12 2 13 15 15 13 2
5 9 13 16 9 2
12 3 9 11 9 13 13 9 13 9 2 15 1
18 3 15 13 13 9 3 15 1 2 16 11 11 13 9 9 9 9 2
7 13 3 3 13 10 9 2
6 11 16 13 13 3 2
4 13 3 3 9
8 13 13 0 13 0 9 9 2
3 13 15 13
15 9 9 11 11 13 9 11 2 16 9 13 2 3 13 2
10 12 0 13 9 7 13 15 9 3 2
2 0 9
6 13 3 3 9 15 2
13 9 11 12 9 11 11 0 9 13 3 13 9 2
5 15 13 13 9 2
11 13 2 16 9 13 0 9 13 0 9 2
3 11 13 9
4 9 13 9 2
7 9 13 13 3 0 9 2
9 0 8 7 9 13 15 1 3 2
10 13 11 0 9 7 13 0 9 15 2
4 11 9 12 13
10 0 9 1 11 9 13 13 0 9 2
7 10 9 13 9 1 9 2
8 15 13 9 7 13 15 9 2
15 9 13 3 13 2 16 9 1 9 9 13 3 12 9 2
13 9 13 3 13 13 9 2 7 15 13 9 1 2
10 15 13 0 9 15 13 12 0 9 2
10 9 13 3 12 7 3 12 9 9 2
15 16 13 13 3 3 3 2 13 15 3 3 0 9 15 2
8 3 0 9 13 9 13 9 2
2 13 9
5 13 15 13 0 2
5 11 13 13 9 2
13 3 9 13 13 2 13 3 16 3 9 13 13 2
3 0 9 9
5 9 13 0 13 2
4 6 16 3 2
10 15 16 13 9 13 2 3 13 13 2
10 11 13 9 9 12 1 13 9 1 2
12 3 3 10 9 13 7 10 9 1 13 13 2
6 13 13 3 10 9 2
3 9 9 9
6 15 13 0 9 0 2
12 3 3 2 0 9 15 13 13 7 3 3 2
16 13 3 13 2 3 13 9 13 2 3 3 13 13 13 9 2
6 13 9 9 7 9 2
11 15 15 13 15 13 13 13 0 9 3 15
2 9 9
7 13 3 13 2 11 13 2
18 11 3 13 13 13 2 16 13 3 0 7 0 9 9 15 1 13 2
12 9 13 13 2 16 9 13 9 3 0 13 2
7 10 9 15 13 13 0 2
12 15 3 13 13 13 2 13 10 3 9 13 2
5 11 7 11 13 9
6 9 9 13 9 9 2
4 16 13 15 2
4 15 13 13 2
6 16 13 3 2 16 2
7 15 13 12 7 12 1 2
9 9 11 13 9 13 13 15 13 2
16 9 7 9 13 3 2 3 13 7 13 7 3 3 13 13 2
28 3 15 13 13 16 15 15 3 9 13 16 13 10 11 6 6 6 9 13 3 9 1 6 13 9 0 9 9
6 9 12 9 13 0 2
8 9 9 13 3 0 2 13 2
7 13 13 10 9 11 11 2
14 9 9 13 13 2 3 9 13 13 3 3 0 9 2
12 13 3 9 9 11 2 15 13 13 11 9 2
7 13 11 15 13 9 1 2
4 9 9 9 0
6 9 13 9 0 9 2
6 13 15 13 3 15 2
2 13 3
7 13 9 9 2 13 15 3
11 9 13 12 9 12 9 7 12 9 9 9
4 3 13 3 2
13 13 3 3 0 9 2 3 9 13 0 9 9 2
15 13 0 9 9 2 0 9 13 10 9 2 13 9 9 2
2 9 13
8 3 10 11 9 15 13 13 2
16 15 13 11 13 9 3 0 9 10 10 9 16 11 9 9 2
18 13 13 9 9 2 9 2 13 0 9 3 9 7 9 9 9 1 2
13 7 3 13 9 13 3 7 13 9 2 9 0 2
10 13 13 2 16 9 13 3 10 9 2
6 15 13 13 3 13 2
11 11 11 13 9 9 7 11 16 11 9 2
9 15 13 13 0 9 15 13 13 3
14 13 9 13 3 0 9 1 7 13 3 13 1 9 2
7 9 13 0 9 2 16 2
5 15 13 11 11 9
4 15 3 13 2
5 9 13 9 13 2
6 15 13 12 9 9 2
5 15 13 13 13 2
9 0 9 2 13 13 13 13 0 2
5 13 3 3 9 2
7 0 15 13 2 9 9 2
10 3 13 13 15 3 0 7 13 9 2
11 9 13 9 13 2 16 0 9 13 13 2
13 2 11 11 9 13 3 13 2 2 15 13 3 2
7 12 9 13 13 0 9 2
6 15 13 13 15 13 2
3 10 9 2
2 13 13
3 9 13 9
4 15 15 13 2
3 13 13 13
5 9 13 9 1 2
8 13 9 2 15 13 3 3 2
15 11 13 3 0 9 7 10 0 9 13 13 9 0 9 2
5 9 9 13 13 11
3 9 9 9
2 3 9
11 11 13 9 3 2 3 3 3 0 9 2
8 13 0 2 16 13 3 9 2
4 13 9 13 2
6 13 3 10 10 9 2
3 10 0 9
12 6 2 3 13 13 9 2 15 13 0 13 2
13 3 13 3 3 2 13 3 13 3 13 13 3 2
4 10 9 9 9
15 13 0 16 3 15 13 3 3 7 15 13 2 13 3 3
7 13 15 13 13 9 12 2
5 0 9 7 9 2
10 9 1 13 9 7 13 15 13 9 2
9 15 13 0 2 7 15 13 9 2
2 11 2
6 15 15 3 3 13 2
6 15 13 9 13 13 2
6 11 13 2 13 9 2
4 13 10 9 2
4 13 3 13 2
2 13 13
5 15 13 3 9 2
2 13 9
3 9 13 13
7 3 15 13 10 0 9 2
5 9 9 13 12 12
8 16 15 13 13 2 13 3 13
9 3 3 9 13 13 9 9 13 2
10 9 13 9 7 9 9 13 9 7 9
3 15 13 0
25 11 9 13 3 3 13 9 2 9 9 2 15 13 13 9 9 1 7 15 13 9 3 9 9 2
5 13 13 15 13 2
30 15 13 3 9 9 16 15 13 3 9 16 15 13 9 13 3 3 9 13 3 7 2 0 3 10 9 13 9 3 2
7 15 13 3 0 9 9 2
13 9 13 9 2 9 7 9 13 7 13 9 13 2
7 0 9 9 13 9 9 2
15 9 9 13 3 2 16 9 9 13 3 3 13 7 13 2
3 15 15 2
15 9 13 0 13 9 9 2 15 13 7 9 13 9 13 2
7 9 15 13 3 12 9 2
12 9 13 11 11 13 2 16 15 13 9 3 2
3 9 0 11
4 0 9 13 0
7 3 0 13 10 0 9 2
18 9 13 3 12 2 9 0 9 2 10 15 0 9 7 15 13 9 2
6 9 13 3 11 9 2
15 9 13 2 9 13 7 0 9 13 2 15 13 9 9 2
11 13 13 0 3 2 7 13 3 9 1 2
17 15 13 3 13 10 9 10 11 2 15 15 7 11 13 0 9 2
10 15 13 2 16 13 13 3 13 9 2
26 16 3 9 13 0 2 13 11 7 11 13 13 0 9 9 2 15 13 9 7 13 0 9 9 11 2
9 10 12 0 9 9 13 12 9 2
11 11 1 3 12 10 9 13 9 0 9 2
4 9 15 13 9
17 11 11 9 12 9 1 9 13 13 9 1 7 3 0 9 1 2
23 10 0 9 2 0 9 2 13 11 9 2 16 13 13 3 9 2 3 13 9 9 13 2
5 13 9 10 9 2
11 0 9 13 13 0 7 3 3 0 13 2
15 11 13 9 15 2 16 0 0 9 13 13 0 9 9 2
9 3 0 13 9 3 0 12 9 2
9 9 13 9 13 3 9 9 1 2
10 9 15 1 13 3 0 7 0 9 2
9 3 9 13 9 11 13 3 12 2
12 13 15 2 3 13 9 2 15 11 13 0 2
2 0 9
12 11 13 13 3 3 0 16 9 9 13 13 2
5 15 13 13 9 2
4 10 9 9 2
11 16 15 13 13 9 2 9 13 9 13 2
2 0 9
6 13 9 7 9 9 2
7 13 15 13 10 9 3 15
9 11 7 15 13 16 9 7 9 2
7 9 11 13 11 0 9 2
6 12 12 0 13 9 2
21 16 15 15 3 13 16 16 15 13 3 9 9 13 16 16 15 13 3 9 13 2
5 10 9 13 0 2
7 0 9 13 13 3 9 2
4 13 13 9 2
7 9 9 13 12 9 1 2
5 9 9 13 9 2
30 13 2 16 12 9 13 10 9 3 13 2 16 9 13 3 13 2 16 13 3 9 3 7 16 9 3 15 13 3 2
4 3 15 13 2
5 9 13 1 11 2
18 15 13 3 3 15 2 16 11 13 13 13 10 9 2 11 13 9 2
2 13 3
4 13 15 3 2
12 0 2 0 12 9 9 13 13 9 3 3 2
8 0 7 0 9 13 9 3 2
4 3 13 13 2
13 9 9 13 0 2 16 8 7 9 13 13 0 2
10 9 1 9 13 8 2 8 7 0 2
8 10 15 13 13 7 13 9 2
9 15 13 13 3 2 3 15 9 13
11 2 15 13 3 2 16 3 15 3 13 2
11 15 13 13 2 13 0 9 7 13 9 2
9 0 9 15 1 13 3 0 9 2
9 0 9 13 13 9 12 9 1 2
6 13 9 9 3 9 2
11 9 13 9 13 13 9 13 9 0 9 2
4 13 7 13 2
4 13 0 9 2
12 15 7 11 13 13 11 3 3 3 2 16 2
3 0 9 11
7 3 13 0 13 7 13 2
5 13 15 13 9 2
6 9 1 9 13 0 2
7 13 9 7 13 9 3 2
8 9 9 13 0 7 9 0 2
12 12 9 2 0 3 12 1 2 13 3 9 2
8 15 13 0 15 15 13 13 2
12 11 11 13 15 3 16 15 13 15 7 15 2
22 16 9 13 13 2 13 13 3 9 2 15 13 9 13 10 9 2 15 15 9 13 2
12 16 13 9 2 13 16 13 13 9 10 9 2
9 0 9 11 13 15 1 9 9 2
10 9 13 3 9 13 10 13 9 1 2
3 13 13 9
17 15 13 15 3 9 9 15 15 13 16 15 13 11 3 3 9 2
3 9 13 13
4 0 0 0 9
2 13 13
10 15 13 13 9 3 0 2 9 13 2
9 2 7 3 3 16 13 9 0 2
6 13 9 7 9 9 2
3 13 15 1
12 9 9 3 13 3 12 9 9 1 9 9 2
3 13 0 2
5 9 13 0 9 15
5 15 13 13 13 15
14 9 9 11 13 13 3 13 2 16 13 9 12 9 2
4 13 13 13 2
8 0 9 13 13 11 13 9 2
17 15 13 9 9 0 9 2 15 9 13 9 9 9 11 9 9 2
4 2 13 13 2
2 0 9
16 10 9 13 15 2 15 13 9 16 15 13 7 13 7 13 2
4 3 13 11 2
8 9 15 13 3 9 7 13 2
14 7 11 13 9 13 3 0 2 16 15 13 3 11 2
11 16 11 13 3 2 3 13 13 3 3 2
6 3 13 9 13 9 2
3 13 10 9
6 15 13 13 15 3 2
4 15 13 0 9
11 0 13 3 2 13 3 12 0 9 9 2
6 13 7 13 9 7 15
3 13 3 3
6 9 13 13 13 9 2
3 15 13 13
5 9 13 2 3 13
4 13 16 13 13
2 13 13
7 15 13 9 13 9 1 2
8 10 9 9 9 13 13 3 2
7 9 15 1 13 0 9 2
8 13 15 0 10 0 9 9 2
3 3 3 16
1 11
8 2 13 3 15 13 0 2 2
13 15 13 13 7 15 13 13 3 7 3 0 9 2
16 13 9 2 13 13 3 2 13 13 9 2 13 7 13 0 2
18 0 9 13 13 3 3 12 9 2 15 3 12 13 13 0 9 9 2
4 3 13 13 2
7 2 13 9 2 7 9 2
5 9 13 13 13 9
2 13 13
5 10 9 13 13 2
7 9 9 13 13 13 9 2
8 10 9 13 13 9 12 9 2
21 11 13 9 12 12 9 13 9 13 0 9 2 15 13 13 3 9 9 13 9 2
6 3 13 9 13 9 9
20 11 13 13 11 9 9 2 7 13 15 1 2 16 9 13 13 3 16 9 2
9 13 15 2 16 15 13 3 0 2
6 0 9 13 9 9 2
11 15 13 9 9 13 13 9 9 3 3 2
11 9 13 3 9 9 2 15 13 13 9 2
5 3 13 0 9 2
4 13 15 15 13
9 3 13 13 3 11 2 13 9 2
7 10 9 13 13 0 9 2
6 15 13 13 9 3 2
4 9 13 0 2
4 6 9 10 9
12 9 13 9 3 2 3 9 13 3 3 3 2
19 15 13 3 3 15 13 16 15 13 13 16 3 15 13 3 16 6 9 2
9 11 3 13 11 13 3 12 9 2
9 15 13 16 15 15 15 3 3 13
5 13 15 9 3 2
4 9 13 12 2
11 11 13 13 9 1 9 12 9 9 0 9
10 13 3 0 13 7 13 3 9 1 2
3 13 11 1
19 9 13 9 13 3 9 3 9 2 3 9 13 3 10 12 9 9 1 2
3 13 11 2
17 9 9 13 8 2 8 7 9 2 15 13 9 2 9 7 9 2
16 0 9 13 9 2 16 9 7 9 13 13 3 3 3 3 2
9 9 10 9 13 3 3 7 3 2
12 10 9 9 13 13 12 9 7 12 9 9 2
13 15 13 16 13 3 3 9 16 13 3 3 9 2
14 13 11 11 11 7 15 13 3 3 3 13 10 9 2
5 11 13 9 9 2
4 13 3 9 2
11 16 0 9 13 13 13 2 13 15 13 2
7 0 9 11 13 0 9 2
6 3 13 13 3 9 2
13 9 13 13 13 9 2 15 13 10 9 13 3 2
7 15 13 3 13 9 3 2
7 13 3 3 10 9 13 2
6 9 13 9 3 0 2
6 15 13 16 13 0 9
4 9 13 15 2
7 15 13 9 0 9 1 2
6 13 13 11 9 3 2
12 15 13 0 9 2 13 15 13 3 12 9 2
2 0 9
12 2 6 13 15 10 12 9 15 10 9 13 2
10 9 13 3 16 3 13 13 10 9 2
5 12 0 9 13 9
4 9 13 3 9
2 9 13
8 9 13 9 2 15 13 0 9
8 11 7 11 11 13 13 0 2
6 11 13 9 13 13 15
13 16 13 11 2 13 9 3 9 7 13 0 9 2
4 15 13 13 13
15 9 13 2 3 11 7 9 11 9 13 2 0 9 2 2
4 9 13 3 2
7 0 9 15 13 13 9 2
11 13 10 9 13 0 13 9 9 9 9 2
9 12 9 13 16 13 13 9 9 2
8 16 15 13 2 13 13 0 2
20 11 13 3 0 2 0 7 0 11 9 2 15 1 11 13 3 3 13 9 9
10 15 13 13 9 9 15 3 16 9 2
13 9 8 13 0 9 2 13 11 13 13 3 3 2
2 0 9
14 11 2 3 13 11 2 13 9 7 13 9 11 11 2
6 9 13 0 0 13 2
4 9 13 9 2
15 11 2 12 0 9 15 13 9 0 9 2 13 15 9 2
19 10 13 9 13 0 9 9 2 15 13 3 13 3 0 16 3 9 9 2
8 13 16 13 13 9 9 1 2
11 12 10 0 9 13 9 9 3 0 9 2
6 13 3 13 9 3 2
4 9 13 9 2
6 3 13 3 9 9 2
7 13 10 9 3 13 9 2
7 15 1 13 3 3 9 2
5 15 15 3 13 2
12 0 11 11 13 11 13 9 9 9 11 11 2
6 11 13 13 0 9 2
9 15 13 3 13 9 10 3 9 2
12 13 13 15 2 13 13 2 3 3 10 9 2
11 7 13 9 3 2 10 0 9 13 9 2
14 11 13 3 9 9 1 11 2 15 10 9 3 13 2
3 13 9 13
8 15 10 9 13 9 15 15 13
7 9 13 3 7 13 9 2
7 13 3 13 13 15 9 2
3 13 13 13
6 0 9 13 12 9 2
13 9 9 13 13 9 9 7 9 13 10 9 0 2
4 9 13 3 2
5 13 13 13 15 2
4 3 15 13 13
3 9 0 9
6 9 9 7 0 9 2
5 13 13 15 0 2
6 9 13 9 0 9 2
3 13 3 2
5 13 15 3 3 3
3 0 9 9
6 9 1 13 13 9 2
5 11 13 12 0 2
10 9 13 0 2 16 15 13 13 15 2
4 9 13 9 2
6 13 9 7 13 9 2
9 9 13 2 16 13 13 10 0 2
4 15 13 13 15
19 9 13 13 15 2 7 3 13 2 3 2 16 13 9 13 13 0 9 2
5 15 13 3 13 2
4 13 0 9 2
13 16 13 9 13 12 0 9 2 7 13 13 9 2
7 11 9 13 0 0 9 2
6 3 15 13 13 15 2
13 11 9 3 13 3 0 9 13 0 3 11 9 2
19 3 13 0 7 0 9 11 2 16 3 9 13 13 9 2 16 3 13 2
17 3 15 3 13 16 13 15 3 15 3 13 10 9 15 15 13 13
8 9 9 13 13 9 9 9 2
3 9 13 13
8 11 11 13 0 9 9 9 2
2 13 15
6 9 1 9 13 0 2
8 13 10 11 2 15 3 13 2
5 9 13 3 3 2
8 9 13 13 3 3 9 1 2
4 2 13 3 2
5 15 13 13 15 2
10 9 13 3 9 9 7 0 9 1 2
17 16 13 13 10 0 9 2 11 0 9 13 3 13 9 9 1 2
8 3 13 13 3 9 12 9 2
8 13 15 13 3 16 10 9 2
2 13 9
6 0 9 13 0 9 2
3 9 13 13
6 12 9 11 13 12 2
11 10 9 15 13 11 1 13 2 15 13 2
4 9 13 0 2
5 9 13 12 3 12
7 9 9 13 13 13 9 2
9 9 13 3 3 0 16 0 9 2
11 11 13 3 13 11 7 13 3 13 9 2
14 9 13 7 13 11 11 2 16 15 13 13 11 9 2
4 0 13 9 2
13 10 0 9 9 13 3 1 15 13 11 11 9 2
8 13 3 9 7 9 13 13 2
12 7 16 9 13 9 1 2 9 13 13 0 2
3 13 0 2
3 9 13 2
13 3 9 13 3 0 9 0 12 9 9 11 11 2
7 3 9 13 3 0 0 2
12 11 13 9 9 0 1 3 3 16 13 13 2
2 10 11
4 15 13 9 2
2 13 13
11 9 11 11 13 13 9 0 9 12 9 2
6 10 9 15 3 13 2
2 9 13
5 13 15 9 0 2
5 13 13 15 15 2
8 9 9 13 13 12 9 13 11
7 9 0 9 13 13 0 2
5 9 9 0 0 9
8 15 15 13 13 3 0 9 2
5 15 13 15 9 2
4 3 13 9 2
3 10 0 9
3 12 0 9
2 9 9
10 9 13 3 0 9 2 15 13 9 2
4 15 13 0 2
9 0 9 13 13 9 13 13 9 2
12 9 1 12 0 9 9 13 9 13 9 9 2
14 3 10 9 13 9 9 1 0 13 9 3 0 9 2
12 16 9 13 9 9 2 15 13 9 9 1 2
4 9 13 9 2
9 3 13 10 11 7 10 10 9 2
6 13 3 0 13 9 2
13 0 9 13 13 9 2 13 11 13 3 0 9 2
5 15 13 13 9 2
9 9 13 13 3 0 13 15 9 9
14 10 10 0 11 13 9 9 3 7 13 3 10 9 2
3 13 3 2
8 9 7 9 13 12 0 9 2
22 16 11 12 9 1 13 0 9 2 15 13 13 9 1 12 11 9 0 11 0 9 2
2 13 13
13 3 11 13 7 13 3 13 10 0 7 0 9 2
4 9 9 13 9
8 2 13 15 16 15 9 13 2
4 13 11 9 2
7 0 0 9 13 12 0 2
7 7 12 9 13 13 3 2
9 13 13 7 13 13 7 13 15 2
9 9 13 15 3 9 1 13 9 2
12 13 13 9 7 10 0 9 12 9 1 9 2
5 15 13 10 0 9
5 15 13 13 3 9
3 12 9 9
7 13 16 15 13 0 9 2
7 13 2 16 3 13 9 2
19 9 9 9 13 2 3 2 0 9 2 0 3 2 9 7 9 9 1 2
9 11 13 13 0 7 11 0 9 2
11 15 13 10 9 15 13 0 9 3 12 2
3 0 9 2
7 13 9 12 9 13 9 2
9 3 13 13 3 15 2 11 13 2
19 3 0 9 9 9 3 9 13 3 15 1 2 16 9 9 3 13 9 2
8 11 13 9 3 9 0 9 2
17 9 7 3 9 13 0 9 13 9 9 7 13 15 0 9 9 2
4 3 0 0 9
8 3 9 13 3 9 13 9 2
2 13 3
8 9 2 3 0 15 13 13 2
7 9 9 7 9 13 9 2
7 11 13 3 0 16 15 2
6 13 2 16 6 9 2
3 13 9 3
13 9 1 3 12 9 9 13 0 13 9 9 1 2
2 6 9
2 13 9
18 13 15 13 15 2 3 10 9 13 3 16 11 11 13 2 11 13 2
6 15 3 13 9 9 2
6 11 13 9 13 9 2
5 11 13 3 9 2
6 0 9 13 3 9 2
13 9 13 13 0 9 2 15 13 3 0 13 3 2
12 15 13 0 7 0 2 0 2 7 3 0 2
16 11 9 13 9 0 2 16 10 9 13 9 9 13 9 9 2
5 15 13 0 13 15
5 11 13 10 9 2
15 11 12 11 13 0 9 3 9 2 9 11 12 2 1 2
22 2 15 11 13 2 9 13 9 13 12 9 2 15 13 3 0 9 13 3 0 9 2
1 12
11 0 9 9 13 12 9 2 16 15 13 2
6 9 1 13 0 9 2
6 3 13 10 9 9 2
2 13 2
21 9 13 9 9 13 15 2 16 12 9 13 13 9 7 0 9 1 12 9 9 2
8 13 16 9 13 13 3 0 9
24 13 13 3 13 9 10 0 9 9 15 13 3 9 7 3 13 3 9 9 7 10 0 9 2
6 15 13 3 0 9 2
21 7 16 15 13 13 13 13 3 3 10 10 9 16 10 10 9 15 13 13 13 2
12 0 9 13 15 2 16 13 9 13 0 9 2
6 13 9 3 13 3 2
3 9 13 13
17 7 3 15 13 0 9 16 11 11 11 15 3 9 1 13 10 9
5 11 13 3 13 2
6 15 11 9 13 3 2
8 0 9 13 2 13 15 9 2
13 9 1 9 11 13 13 10 9 3 0 0 9 2
3 11 13 11
4 11 3 11 9
19 9 13 15 3 3 9 9 15 1 2 16 9 13 13 16 9 13 9 2
3 15 13 11
16 15 1 15 13 9 16 15 13 13 13 3 13 10 0 9 2
8 15 13 16 13 13 15 15 2
2 9 0
10 3 10 13 9 9 2 7 15 13 0
2 0 9
4 3 9 13 2
14 15 1 15 9 13 2 16 15 13 2 9 13 9 2
6 9 15 13 3 11 2
5 9 9 13 0 2
5 9 13 0 9 2
15 13 15 13 15 15 13 2 13 15 15 13 2 0 9 2
4 11 9 13 9
8 9 13 9 13 13 3 9 2
11 6 13 15 9 3 13 2 16 15 13 2
6 3 13 9 9 9 2
5 9 13 11 11 2
3 13 3 2
6 15 13 3 10 0 2
14 7 13 13 9 2 16 9 13 9 2 3 13 9 2
6 3 13 0 13 9 2
2 9 9
11 3 15 7 10 15 1 9 13 0 9 2
15 9 7 3 9 13 13 13 9 0 7 0 9 9 1 2
15 9 13 10 11 2 15 13 13 9 3 9 11 11 1 2
4 9 13 9 2
9 11 9 13 13 2 16 9 13 2
6 13 13 11 7 11 2
4 13 0 9 2
9 9 13 3 3 9 3 9 9 2
7 13 13 0 9 13 9 2
5 15 13 9 3 2
8 13 15 13 9 2 10 9 2
11 13 7 0 7 0 2 13 13 13 15 2
2 9 9
4 13 9 13 2
9 9 1 9 13 9 1 13 13 2
8 13 2 16 9 13 10 0 2
5 9 1 13 9 2
6 9 13 0 16 9 2
20 3 9 13 3 0 2 7 0 7 0 9 13 3 2 16 0 9 13 2 2
5 16 13 13 3 2
14 13 9 10 11 12 9 13 9 9 9 3 3 13 2
12 13 2 16 13 0 9 13 0 10 0 9 2
12 11 13 2 16 9 2 3 2 13 15 9 2
9 13 9 9 7 13 0 9 1 2
4 15 13 9 2
11 3 13 13 9 2 3 13 3 12 12 2
20 9 12 9 11 11 9 11 2 15 13 11 11 2 15 13 3 11 9 2 2
19 15 13 15 9 11 0 9 2 15 13 13 9 15 1 7 11 9 9 2
9 13 15 13 10 9 2 15 13 2
6 12 9 13 13 9 2
14 13 3 0 13 2 16 3 13 9 2 15 13 3 2
3 0 9 15
2 0 9
12 2 9 13 13 13 2 2 9 13 9 12 2
5 9 13 3 0 2
3 13 13 2
9 11 13 13 13 9 9 7 9 2
10 10 9 7 11 7 15 13 10 9 2
12 11 3 9 9 13 3 0 13 10 0 9 2
8 6 0 9 15 3 13 13 2
12 11 13 9 2 7 13 9 13 10 9 13 2
10 7 12 7 0 9 13 9 0 9 2
10 9 13 0 9 0 9 9 9 9 2
6 9 9 13 3 0 2
8 3 3 12 12 9 13 13 2
9 9 9 13 9 13 9 9 9 2
18 0 9 9 13 10 3 0 2 16 0 9 13 3 13 13 15 3 2
8 9 9 0 9 13 9 12 2
4 3 7 3 2
13 9 13 3 10 9 2 16 11 13 13 10 9 2
6 13 16 15 13 3 0
9 13 0 9 0 9 3 3 1 2
3 13 13 9
7 7 16 15 13 12 0 9
6 16 13 3 13 3 2
9 15 15 15 13 16 15 3 13 2
8 15 13 0 9 9 16 15 2
7 11 13 3 16 13 9 2
9 11 9 13 9 9 13 13 9 2
5 3 15 9 13 2
10 15 13 13 0 9 9 7 9 9 2
2 0 9
6 3 12 13 9 3 2
20 0 9 13 9 9 12 2 7 10 9 13 13 0 12 9 12 0 9 1 2
15 11 13 3 12 0 2 15 10 9 13 3 13 9 9 2
9 9 7 9 1 13 13 13 9 2
13 9 9 1 2 9 13 3 3 9 0 9 9 2
11 3 15 13 3 2 7 15 13 13 9 2
20 10 9 2 9 7 9 7 10 9 9 2 13 3 16 13 9 9 13 3 2
11 15 13 9 13 15 2 7 13 13 9 2
18 10 0 9 7 9 13 2 10 9 7 15 1 13 15 13 0 9 2
8 10 9 13 13 9 7 9 2
16 16 3 0 13 2 11 13 3 0 2 3 9 7 9 9 2
3 2 15 2
12 9 13 13 3 9 0 9 2 13 15 9 2
13 9 2 15 13 13 13 9 10 3 0 9 9 2
8 10 9 13 13 3 9 9 2
10 9 13 3 9 0 12 9 9 1 2
8 9 15 13 9 7 9 9 2
10 13 13 15 13 2 16 13 9 9 2
14 13 11 9 9 9 13 2 15 15 13 9 9 11 2
2 13 13
15 13 3 13 9 9 2 16 3 13 9 7 16 15 13 2
6 15 13 16 13 9 2
6 3 3 9 13 13 2
2 0 9
6 3 13 3 10 0 2
5 6 15 15 13 2
12 0 13 13 3 2 13 11 7 13 0 9 2
5 9 13 9 9 2
14 0 13 13 9 11 2 15 9 13 0 16 9 9 2
10 3 16 9 9 13 13 13 3 13 2
10 9 13 2 7 16 13 2 3 9 2
11 0 11 9 13 2 9 7 9 9 2 2
7 11 13 0 9 0 9 2
7 15 13 3 9 13 3 2
17 0 1 13 3 0 13 2 7 0 9 13 13 13 0 9 9 2
10 3 11 15 9 13 2 15 13 13 2
15 3 9 13 13 9 13 9 12 9 0 9 0 9 1 2
10 11 13 13 9 10 9 10 9 0 2
12 9 13 9 2 15 13 7 3 7 3 1 2
6 15 13 3 0 9 2
3 15 13 9
9 15 2 9 9 2 13 13 15 2
7 9 13 13 9 7 13 2
6 13 9 13 7 13 2
6 15 13 13 13 9 2
10 9 9 13 0 9 2 7 13 15 2
19 3 13 13 9 9 3 15 1 13 0 9 1 2 13 15 9 7 9 2
7 15 13 0 13 3 9 2
2 0 0
11 3 13 13 2 13 9 13 8 7 9 2
20 11 9 13 13 1 11 9 2 13 13 10 9 2 15 13 3 13 7 13 2
3 13 13 13
26 11 11 13 11 2 16 13 11 11 9 3 13 2 16 13 15 13 2 7 3 2 16 13 9 13 2
6 13 3 9 11 1 2
3 9 9 0
8 15 13 3 16 13 9 13 2
6 12 9 13 11 10 9
16 10 9 13 13 0 9 9 2 15 13 2 15 15 3 13 2
5 9 13 13 13 2
13 0 9 13 15 2 13 0 0 9 0 7 0 2
7 9 9 9 3 13 13 2
8 3 9 9 2 15 13 3 2
2 9 1
16 16 9 3 13 11 1 2 7 3 13 2 11 13 9 13 2
9 13 13 13 10 9 3 15 13 2
8 11 1 9 13 11 11 1 2
4 13 3 13 9
2 0 9
11 15 9 13 2 11 9 9 9 11 11 2
9 3 9 13 3 0 16 12 9 2
6 9 13 9 13 9 2
28 7 13 3 2 3 15 13 3 3 15 13 3 13 15 13 3 3 13 16 15 13 3 3 15 1 15 3 13
6 11 9 13 12 9 2
8 15 13 9 13 0 9 1 2
4 13 13 9 3
8 9 13 3 13 0 9 9 2
6 9 13 13 1 9 2
4 15 13 13 2
8 3 10 9 13 3 9 13 2
19 16 15 13 9 7 9 12 9 2 3 13 15 9 9 0 0 9 9 2
3 9 13 9
9 13 13 2 13 13 2 13 13 2
4 11 11 13 9
5 3 13 9 13 2
7 13 0 16 13 13 9 2
4 3 15 13 2
3 11 13 0
2 3 11
9 9 9 13 3 13 11 7 11 2
2 3 3
16 3 13 2 16 13 2 16 9 13 0 9 7 9 13 9 2
12 15 13 13 3 0 2 3 15 13 3 0 2
18 16 9 3 13 15 2 15 3 15 7 9 13 10 9 13 9 13 2
10 11 13 3 0 9 2 0 13 0 2
10 16 13 13 1 9 2 3 0 9 2
7 16 13 2 13 1 9 2
4 7 15 13 2
11 11 13 15 9 13 2 3 16 13 3 2
9 9 0 2 9 0 2 12 9 0
6 13 13 9 3 9 2
10 7 9 9 7 9 9 13 13 9 2
6 15 13 9 9 1 2
3 9 13 13
12 9 13 9 2 16 13 13 9 13 13 3 2
7 13 9 13 11 1 13 2
12 10 11 13 3 3 11 9 16 13 13 9 2
14 9 13 3 3 0 9 9 2 15 13 3 12 9 2
9 9 9 13 3 13 3 0 9 2
8 9 13 9 13 13 15 3 2
8 13 15 13 12 7 10 3 2
18 9 1 9 9 13 13 13 9 9 0 9 2 16 9 9 13 9 2
9 11 13 1 9 11 11 9 9 2
23 9 7 9 13 3 3 9 13 9 7 13 15 7 3 13 9 2 9 2 9 7 9 2
6 13 3 3 0 15 2
4 9 3 13 2
16 16 10 9 13 15 1 13 2 15 13 3 13 13 15 0 2
10 13 0 9 2 15 13 13 12 9 2
7 13 15 3 15 3 13 2
8 9 9 13 10 9 3 7 3
8 0 9 13 9 9 3 3 2
3 0 9 1
15 9 13 13 3 0 2 3 16 15 13 13 2 13 11 2
17 13 13 9 7 13 13 13 9 1 9 2 15 13 15 0 9 2
13 13 13 3 10 3 15 9 3 13 3 13 3 13
7 15 13 3 13 9 9 2
13 13 13 9 2 7 13 16 13 11 13 13 3 2
2 13 9
8 9 11 9 13 10 9 11 2
12 9 13 9 9 2 15 13 0 16 11 15 2
4 0 13 9 2
20 13 13 15 9 3 9 2 7 13 2 16 13 11 3 13 13 15 9 13 2
4 8 13 9 2
6 13 15 15 10 9 2
7 15 13 3 13 9 9 2
5 3 15 13 13 9
13 13 2 16 15 13 15 15 15 7 10 15 13 2
7 9 10 9 7 9 15 2
7 13 15 12 9 0 9 2
9 10 15 13 11 9 1 13 9 2
13 9 13 13 13 3 0 2 7 13 3 3 0 2
20 11 9 13 13 3 2 7 3 16 11 9 9 13 9 13 9 13 9 9 2
6 9 13 9 9 13 2
4 9 13 13 2
5 9 13 13 9 9
6 11 13 0 7 0 2
7 3 13 3 13 9 13 2
9 3 3 3 15 1 2 11 13 2
7 10 0 9 13 13 13 2
3 9 0 9
9 9 13 3 9 7 15 9 0 9
3 0 9 9
6 0 9 3 1 13 9
12 9 0 9 7 9 13 3 3 13 9 9 2
14 9 3 13 15 13 2 7 15 13 9 9 7 9 2
16 10 2 9 13 9 13 9 7 0 9 3 9 16 0 9 2
8 10 9 13 0 7 0 2 2
2 0 9
17 16 9 13 3 9 2 13 9 9 13 3 3 16 10 10 9 2
12 11 11 10 0 9 9 13 11 11 13 11 2
8 15 1 15 13 13 9 9 2
12 15 13 0 13 2 16 9 13 13 3 3 2
14 0 9 9 13 13 10 13 9 9 2 9 9 9 2
9 9 16 9 13 2 9 13 9 2
4 13 15 9 2
11 11 13 9 15 2 15 13 13 0 9 2
13 13 3 0 16 10 9 9 9 13 9 3 9 2
4 9 9 13 3
6 13 11 13 10 9 2
2 10 9
6 9 13 9 9 9 2
2 3 13
5 15 13 13 0 2
5 9 15 13 9 2
10 13 0 13 3 2 7 16 13 13 2
5 9 13 15 13 9
2 0 9
6 3 15 1 13 9 9
10 11 11 11 13 3 1 11 11 9 2
2 0 9
5 11 13 11 9 2
3 13 9 2
11 13 0 13 2 16 11 9 13 3 9 2
11 11 13 13 9 9 2 7 9 13 3 2
4 15 13 15 2
5 13 9 13 9 2
10 9 9 13 10 9 0 16 13 9 2
11 15 13 13 12 7 15 13 3 13 0 9
5 15 13 9 9 2
5 9 13 0 3 2
4 10 9 13 2
9 9 9 11 13 0 9 0 9 2
2 9 9
7 10 9 13 13 0 9 2
7 13 13 3 15 2 13 3
7 9 13 13 2 13 9 2
5 10 9 13 0 9
9 9 13 9 9 13 13 13 3 2
5 0 3 0 9 2
6 9 1 9 13 0 2
8 10 9 13 3 0 7 0 2
7 9 13 3 0 7 9 2
5 13 15 15 13 9
7 3 15 13 13 0 9 2
3 9 13 9
11 7 3 15 13 2 16 9 13 9 9 2
13 0 9 1 9 9 13 13 13 3 12 9 9 2
14 13 13 13 0 0 0 9 2 15 13 3 3 3 13
4 13 0 9 2
8 11 7 11 13 9 11 9 2
2 0 9
15 9 15 13 13 2 13 11 9 13 0 9 13 9 1 2
7 10 9 9 9 13 11 2
11 9 13 15 2 13 9 11 7 10 9 2
5 0 9 13 9 2
3 9 0 9
6 13 9 11 9 11 2
4 15 13 3 3
7 11 9 13 3 12 9 2
2 9 13
8 9 15 1 3 13 0 9 2
5 11 11 13 9 2
15 3 13 3 9 9 9 2 7 3 13 3 3 0 9 2
13 9 9 13 11 13 9 2 7 13 3 0 9 2
8 9 11 13 13 9 9 11 2
14 9 7 0 13 3 7 3 3 9 13 9 13 9 2
10 11 13 13 13 15 7 9 13 9 3
10 15 3 13 2 16 13 3 0 9 2
9 13 3 13 13 9 0 9 9 2
7 16 13 15 3 9 13 2
7 13 9 2 3 9 9 2
6 15 13 9 9 3 2
9 9 3 15 2 15 13 3 9 2
7 3 13 13 10 9 13 2
5 15 13 3 0 2
8 11 13 9 11 9 2 16 2
4 9 9 10 9
3 9 15 13
2 9 9
17 16 15 13 3 9 3 9 3 13 13 3 0 9 16 15 13 2
2 0 9
7 9 13 9 1 12 9 2
9 0 9 15 13 15 2 0 9 2
19 9 13 2 16 9 13 13 9 9 13 9 9 15 3 16 15 15 13 2
6 15 15 13 9 13 2
15 11 11 13 0 9 11 12 7 13 7 11 7 11 9 2
6 11 13 13 9 9 2
6 15 13 3 12 1 2
6 13 3 16 3 13 2
9 3 9 11 13 13 16 3 13 2
4 13 9 3 2
11 13 13 3 0 9 2 16 9 9 13 2
8 11 13 13 13 9 9 13 2
10 3 13 9 2 3 13 9 13 3 2
6 7 9 9 8 8 2
6 13 3 2 12 9 9
6 7 13 3 9 3 2
2 13 13
5 15 13 10 9 2
7 15 13 3 12 9 9 2
9 9 0 9 9 13 3 0 9 2
7 9 9 13 13 9 9 2
4 9 3 9 2
17 0 9 9 13 15 2 16 16 13 13 9 2 13 9 13 3 2
8 9 13 3 9 13 9 9 2
13 9 13 0 13 2 15 13 13 7 13 10 9 2
5 13 15 11 9 2
7 15 13 3 9 13 9 2
5 9 13 13 13 9
7 13 3 2 16 13 9 2
10 15 13 3 2 16 13 13 15 0 2
9 13 13 13 9 2 16 13 9 2
9 15 13 15 2 16 9 13 15 2
8 9 1 9 13 3 13 9 2
2 13 13
10 9 13 3 3 3 0 15 9 13 2
14 3 0 9 13 0 9 13 2 16 3 13 0 9 2
3 0 9 2
29 9 13 3 12 12 9 7 15 10 9 13 3 0 3 15 2 16 11 13 3 12 3 9 2 15 13 10 9 2
15 3 0 9 13 0 2 16 15 13 3 15 3 0 9 2
11 9 13 0 9 0 9 11 2 11 2 11
14 9 9 11 9 12 9 9 13 9 9 9 13 3 2
9 3 13 9 10 9 13 9 9 2
6 16 3 13 2 3 2
7 3 11 13 3 13 15 2
4 9 15 13 2
23 16 15 13 13 10 9 11 9 2 13 15 9 3 7 10 0 15 13 2 15 13 9 2
11 10 9 9 13 3 9 9 9 13 9 2
5 9 13 3 9 2
5 9 9 13 13 2
6 11 13 9 1 9 2
16 11 13 13 2 13 9 9 3 13 0 13 16 0 9 9 2
8 13 15 9 1 13 7 13 2
8 15 3 13 13 9 15 13 2
3 9 0 9
6 9 13 9 13 9 2
5 3 15 3 13 13
3 9 13 2
9 7 9 13 0 9 3 9 9 2
11 9 13 9 13 12 9 13 13 9 3 2
6 13 3 13 15 15 2
4 0 13 15 2
17 9 9 1 13 0 9 13 11 2 15 13 9 2 3 2 9 2
8 9 12 9 13 10 0 9 2
14 9 13 3 13 2 15 13 9 9 9 11 11 13 2
12 9 13 9 13 10 9 2 15 13 9 9 2
23 15 2 16 11 13 3 3 3 13 9 2 11 13 13 9 7 9 2 9 9 7 9 2
10 9 13 2 16 9 15 13 13 9 2
5 10 9 13 3 2
7 11 13 11 9 13 13 2
4 9 15 13 2
8 3 10 9 13 10 9 3 2
3 13 9 2
13 11 11 13 2 16 9 13 13 9 3 10 9 2
10 9 13 3 9 7 9 7 9 9 2
3 11 13 9
6 13 3 0 0 9 2
18 11 11 13 9 2 13 0 12 9 9 9 9 7 13 3 9 9 2
6 9 13 13 9 9 2
6 0 9 13 12 9 2
9 11 16 3 13 13 3 3 9 2
2 3 9
11 13 15 9 1 9 2 0 9 7 9 2
6 9 13 9 9 9 2
17 11 13 2 16 9 13 13 11 11 7 15 0 9 9 7 9 2
5 6 13 13 3 2
3 0 13 9
14 0 9 11 13 3 13 13 9 9 15 16 10 9 2
13 3 11 7 11 13 0 11 9 2 15 13 13 9
6 9 13 10 9 9 2
6 11 7 11 13 13 9
5 13 11 3 7 3
12 10 9 2 9 7 9 10 13 0 9 13 2
6 9 13 13 1 11 2
10 6 3 15 13 12 9 10 11 3 2
2 9 9
5 3 9 13 9 2
15 3 9 13 0 9 9 13 2 7 9 13 15 15 3 2
4 9 13 3 2
7 3 11 3 13 13 3 2
2 10 3
7 9 2 0 9 2 9 2
8 15 13 9 9 1 12 9 2
7 9 13 13 15 13 9 2
16 0 9 13 0 2 16 13 15 3 13 15 13 0 10 9 2
12 3 13 3 3 0 9 9 13 11 2 3 3
8 13 9 3 3 13 13 13 2
12 9 0 9 13 15 2 16 0 9 13 13 2
11 9 13 2 16 3 9 9 13 9 3 2
6 15 13 3 13 9 2
10 3 13 0 9 2 15 9 13 9 2
15 15 13 13 0 9 7 9 9 2 7 12 15 0 9 2
3 13 3 9
13 15 13 2 16 13 15 0 13 13 2 13 0 2
8 11 3 13 9 13 11 9 2
6 10 9 10 15 13 2
7 9 9 13 9 11 9 2
8 9 9 13 9 0 0 9 2
10 13 9 2 13 9 9 7 13 9 2
9 10 9 9 13 3 12 9 1 2
12 15 13 0 9 2 16 9 13 9 16 9 2
4 9 13 3 2
20 9 1 2 15 13 9 12 9 2 13 13 3 12 9 9 3 16 13 9 2
8 10 9 13 9 13 0 9 2
9 7 15 13 13 0 9 7 9 2
23 15 13 10 11 2 9 3 7 15 13 16 15 3 13 15 16 13 3 13 13 15 3 2
13 11 13 2 16 11 13 9 9 3 12 9 1 2
11 13 2 10 9 9 13 13 2 10 9 2
9 3 9 13 12 12 12 9 9 2
4 6 10 9 2
7 9 11 11 13 13 9 2
13 7 3 13 3 0 2 16 0 9 13 0 0 9
2 9 9
2 11 2
6 3 9 13 10 9 2
17 0 9 13 13 13 11 3 9 2 7 9 11 13 9 13 0 2
7 9 9 13 13 3 0 2
6 15 13 9 3 9 2
4 6 16 0 2
2 13 9
9 9 13 11 1 13 10 9 0 2
6 13 3 3 16 13 2
4 3 13 13 2
9 9 13 11 3 13 3 9 13 2
8 10 9 13 3 13 1 15 2
11 15 13 9 2 9 2 9 7 11 9 2
8 9 9 11 9 13 3 9 9
7 9 9 13 0 0 13 2
13 9 11 11 13 10 9 9 9 1 13 0 15 2
9 13 9 13 11 7 9 13 9 2
6 10 9 0 13 13 2
6 10 12 0 3 13 2
3 9 13 3
4 13 9 3 2
9 11 13 9 13 9 3 7 3 2
4 2 13 3 2
20 9 7 9 1 13 3 13 13 9 7 3 10 9 2 3 3 9 7 9 2
9 15 13 3 9 16 10 9 13 13
7 15 13 13 9 13 9 2
11 11 13 0 9 2 15 13 9 1 9 2
5 9 13 13 0 2
7 13 15 13 15 1 13 2
7 9 9 13 9 11 9 2
8 2 0 9 15 9 9 13 2
15 11 13 3 13 13 9 7 9 2 16 15 13 13 15 2
27 16 10 9 13 0 9 2 11 13 9 13 2 7 15 13 3 10 9 2 15 10 9 13 2 9 1 2
14 13 13 15 2 7 15 3 13 13 13 10 0 9 2
8 9 9 9 13 0 16 3 2
3 3 13 2
13 3 9 13 9 12 2 3 9 13 13 12 9 2
6 9 13 9 9 1 2
10 13 9 3 12 9 3 16 13 9 2
4 7 9 13 2
8 3 12 13 7 13 13 9 2
10 9 9 9 7 9 9 13 9 9 2
18 0 9 9 13 13 13 2 10 9 3 3 13 2 7 3 13 13 2
6 15 13 9 13 0 2
4 13 0 9 2
10 0 9 9 13 9 12 9 9 13 2
4 3 7 3 2
5 3 3 13 3 2
5 13 13 9 3 2
7 9 9 2 9 7 9 2
10 9 13 13 13 9 9 13 9 9 2
8 3 9 15 1 13 0 9 2
2 3 0
11 9 13 0 7 0 2 11 13 0 9 2
6 9 1 9 13 13 2
4 9 13 13 2
6 9 13 3 0 9 2
10 13 0 2 16 13 13 2 10 9 2
4 13 9 9 2
6 15 13 3 9 13 2
2 10 9
11 9 13 9 1 9 13 9 9 12 9 2
9 13 15 3 9 15 9 13 9 2
7 15 13 9 3 3 9 2
9 9 13 0 0 9 3 0 9 2
14 7 10 10 9 3 13 13 3 3 13 7 13 15 2
14 3 9 0 7 9 13 13 13 9 3 9 9 9 2
15 10 9 7 9 13 11 3 13 2 15 13 7 3 13 2
7 11 13 9 11 9 9 2
6 3 10 9 13 9 2
8 13 13 13 3 3 10 9 2
4 9 1 9 2
12 9 9 13 3 3 9 2 3 3 16 13 9
7 13 3 15 3 3 9 2
6 15 15 13 13 2 2
17 16 9 1 3 13 2 9 13 13 13 9 11 11 1 1 9 2
20 9 15 13 13 9 13 0 9 7 10 9 13 3 0 9 7 3 0 9 2
6 0 9 13 9 1 2
4 9 13 9 13
4 10 9 12 9
6 3 15 13 3 9 2
4 13 15 3 2
9 15 13 12 9 9 3 13 7 2
5 15 13 3 0 2
7 9 13 13 9 9 9 2
5 9 13 0 9 2
6 13 15 13 9 0 2
7 15 13 9 3 7 13 2
7 15 13 15 9 7 9 2
8 13 3 13 12 9 9 0 9
13 7 16 15 13 13 9 2 3 13 13 13 9 2
29 7 0 10 9 3 15 16 16 13 3 0 9 7 13 3 13 9 3 13 15 13 3 15 16 15 15 9 13 2
13 9 9 13 9 2 16 15 15 13 2 13 3 2
15 9 9 13 9 2 16 13 9 13 13 0 9 13 9 2
5 10 9 13 9 2
3 11 13 13
7 13 13 9 2 7 9 2
7 11 13 9 9 13 11 2
22 15 13 3 0 9 10 10 9 13 9 15 13 15 2 3 16 3 10 9 13 3 0
7 9 13 3 3 13 9 2
9 13 3 2 15 9 13 3 13 2
6 9 13 13 11 9 2
15 11 9 9 13 9 13 0 9 2 0 13 9 12 9 2
6 13 13 3 9 1 2
4 0 9 13 9
5 3 3 13 13 2
3 0 0 9
2 10 9
3 11 0 9
9 9 13 13 9 7 0 9 9 2
11 3 15 13 15 2 16 13 11 7 13 2
8 10 9 13 0 9 13 9 2
8 0 0 9 9 13 3 3 2
9 15 13 9 2 9 7 12 9 2
8 9 13 2 16 13 15 0 2
6 9 9 13 0 9 2
2 3 9
4 9 13 7 13
16 11 13 13 13 3 2 7 13 3 2 3 2 15 13 0 2
12 15 16 9 7 9 13 3 13 3 0 9 2
10 11 13 3 13 9 2 15 13 13 2
10 9 13 7 11 13 7 13 9 9 2
4 15 13 3 13
11 9 13 9 2 12 9 0 9 7 9 2
21 3 3 11 7 11 7 11 13 13 3 16 0 2 16 13 3 13 15 7 13 2
3 13 3 13
3 3 9 2
6 11 13 3 13 3 2
5 7 10 9 3 2
16 9 9 13 3 3 9 13 2 3 9 9 13 3 13 9 2
13 0 7 0 9 2 9 1 2 13 10 11 0 9
8 11 13 16 15 13 13 9 2
17 0 9 2 15 0 9 13 13 9 2 13 16 9 13 0 9 2
13 11 9 13 11 11 2 15 13 0 9 9 9 2
5 13 3 2 9 2
8 3 15 13 15 2 9 13 2
16 15 13 13 13 15 10 9 13 13 13 15 15 13 10 9 2
5 13 3 0 3 2
5 9 13 9 13 2
6 9 13 3 3 3 2
12 11 13 0 2 15 13 13 12 9 0 9 2
20 9 13 11 9 3 3 2 16 9 13 11 9 9 13 3 12 12 9 0 2
33 15 13 13 3 3 3 13 0 0 9 3 15 13 3 3 9 6 9 13 16 13 15 13 16 3 13 13 15 13 3 0 13 2
4 15 3 13 2
16 13 0 13 9 0 8 7 9 2 3 9 13 0 9 13 2
6 9 13 3 0 9 2
17 13 3 2 13 10 0 9 0 9 2 16 13 3 9 12 9 2
9 15 13 2 16 13 3 16 13 2
3 9 13 2
6 13 15 10 3 3 0
3 15 13 9
2 11 9
9 9 9 13 10 9 3 12 12 2
7 11 7 9 13 1 9 2
15 9 13 9 15 13 15 0 9 13 9 3 1 9 9 2
8 13 3 13 13 9 9 3 2
5 9 13 0 9 2
6 15 1 15 13 13 2
8 16 13 0 2 13 13 13 9
21 0 9 9 13 9 13 15 3 3 16 13 12 10 11 9 13 13 9 7 9 2
17 16 13 0 9 9 2 13 15 9 0 9 7 9 13 3 3 2
4 9 13 0 2
11 3 9 13 0 9 2 16 13 3 9 2
7 7 3 13 11 7 11 2
16 3 15 13 3 13 2 16 9 13 3 9 12 13 15 13 2
17 15 13 3 13 9 10 10 9 2 7 9 7 9 13 3 3 2
4 9 9 13 2
9 11 13 13 0 9 12 9 12 2
3 9 13 9
5 9 13 3 15 9
5 9 13 3 9 2
10 9 13 13 13 3 13 13 13 13 2
8 11 9 13 3 12 9 1 2
17 9 13 9 11 2 9 11 2 15 7 12 9 2 11 7 11 2
4 8 7 0 9
7 15 13 3 7 9 3 9
5 9 13 3 13 2
14 11 2 11 2 11 2 11 7 11 13 3 9 0 9
4 3 15 13 9
8 3 13 9 13 7 13 9 2
12 11 13 13 16 13 15 15 13 3 13 3 2
19 9 11 13 9 2 2 3 15 13 13 9 9 2 9 13 13 15 2 2
19 10 9 13 2 16 15 13 9 3 2 16 13 13 3 7 3 10 9 2
6 9 3 13 13 9 2
3 13 3 2
14 13 13 9 9 7 13 2 16 13 3 13 13 9 2
5 9 13 0 9 2
4 13 13 13 2
7 9 11 13 9 9 1 2
9 9 13 9 9 1 7 3 9 2
4 3 9 13 2
12 3 0 7 9 0 9 0 13 0 9 13 9
5 13 13 11 13 2
5 0 9 13 15 2
8 9 11 13 11 9 1 9 2
5 13 13 9 11 2
10 2 13 1 9 2 2 13 15 13 2
7 13 13 3 2 7 13 2
5 9 13 3 9 2
4 13 9 9 2
13 16 9 13 3 11 2 13 9 0 9 9 9 2
13 2 3 3 13 13 7 15 13 2 2 13 9 2
5 9 13 3 0 2
6 15 13 2 13 9 2
5 9 13 3 0 2
8 3 13 9 1 2 3 9 2
4 10 9 13 15
12 11 13 9 3 0 9 2 16 13 13 9 2
11 10 9 15 13 7 13 11 13 9 13 2
20 3 11 13 9 3 9 7 9 2 7 15 13 12 11 9 12 9 12 9 2
13 9 11 11 7 11 11 13 9 3 11 11 1 2
5 13 0 9 13 9
10 15 13 13 9 2 7 9 15 13 2
12 0 7 0 9 0 9 13 13 12 12 9 2
7 9 13 13 7 9 13 2
6 6 2 0 2 3 2
5 15 13 11 3 3
22 9 13 13 13 0 9 9 2 3 3 1 15 2 16 10 9 13 13 9 3 3 2
2 16 3
8 3 13 3 9 7 10 0 2
20 9 13 13 3 2 16 13 9 13 13 9 13 9 9 7 13 0 9 9 2
5 11 13 9 0 2
10 0 9 13 13 2 15 13 13 9 2
3 9 13 9
11 11 13 9 9 1 11 7 9 1 11 2
5 9 13 13 9 2
5 15 13 13 9 2
2 0 9
7 9 13 13 3 9 3 2
5 9 13 9 0 2
5 9 13 13 9 2
10 3 15 13 13 13 7 9 7 9 2
4 9 13 0 2
3 0 15 13
10 9 13 9 7 9 10 12 9 1 2
7 9 13 0 16 13 13 2
13 9 9 13 9 2 7 9 1 9 13 3 0 2
11 13 9 9 11 7 11 13 3 9 9 2
6 15 13 3 0 15 2
4 9 1 13 2
14 11 9 13 7 13 2 16 15 13 16 13 0 9 2
9 3 10 9 13 3 15 15 9 2
5 15 13 10 9 2
8 13 13 0 9 2 16 13 2
6 9 9 13 3 13 2
16 9 13 13 9 2 15 13 3 13 7 13 3 0 7 0 2
14 9 3 11 13 3 3 2 15 1 11 13 13 13 2
5 15 13 9 3 2
3 9 13 9
15 9 13 9 9 2 3 16 10 9 13 13 13 9 9 2
7 13 13 13 1 9 9 2
13 15 3 11 13 9 3 13 9 13 12 9 9 2
12 3 9 2 3 9 2 13 9 2 16 9 13
2 0 9
8 6 3 2 13 15 9 9 2
19 9 9 1 13 9 9 1 2 7 15 13 15 2 16 13 15 3 9 2
2 3 9
5 13 16 15 13 2
2 9 13
7 13 15 10 9 2 9 2
4 13 15 13 2
2 13 9
8 7 3 9 9 13 15 13 2
10 9 9 13 9 12 7 13 3 9 2
4 0 9 13 11
8 9 0 9 0 9 13 9 2
9 16 13 3 3 1 12 3 11 2
12 9 2 9 9 7 3 9 13 0 3 9 2
9 11 1 9 13 13 9 3 3 2
18 15 2 16 3 13 13 9 9 9 7 2 9 2 13 9 11 9 2
5 9 13 0 0 9
3 13 13 2
4 13 3 3 2
4 11 13 3 9
16 9 1 9 9 13 15 2 16 9 9 13 9 11 9 9 2
12 11 13 11 11 13 9 9 8 7 9 9 2
22 0 9 13 15 2 15 13 3 13 9 2 7 13 13 2 3 13 3 7 13 3 2
7 13 3 13 3 9 9 2
9 15 3 13 2 7 13 3 9 2
8 15 13 9 7 13 10 9 2
5 15 13 9 13 15
9 2 9 2 1 9 2 13 2 2
10 15 13 3 0 2 0 7 9 9 2
14 11 7 11 13 3 2 7 3 3 13 3 3 13 2
4 3 13 3 2
8 11 9 11 13 9 0 9 2
4 15 15 13 2
14 11 13 3 15 13 13 13 9 13 0 9 9 1 2
16 13 3 13 11 9 1 3 2 7 15 13 13 9 13 15 2
5 9 13 12 9 2
15 16 11 13 2 13 15 9 9 2 11 7 11 3 9 2
8 9 13 15 2 16 13 9 2
14 15 13 13 9 3 9 2 16 13 13 7 13 13 2
3 13 13 2
6 9 9 13 10 9 2
14 15 13 3 13 16 13 3 0 15 13 2 11 13 2
3 3 13 15
12 9 13 2 16 15 1 9 13 3 7 13 9
4 9 13 9 3
5 10 9 11 13 2
2 9 9
7 15 13 3 10 3 13 2
3 11 9 9
9 15 13 13 9 13 9 13 9 9
11 9 13 3 13 10 0 9 0 9 2 2
4 0 9 7 9
4 15 13 13 2
3 9 13 13
6 9 9 13 13 3 2
4 12 15 13 9
2 0 9
13 9 0 9 3 15 13 9 9 2 0 9 13 2
8 9 13 9 3 7 3 9 2
11 9 13 10 9 2 16 9 9 13 13 2
12 15 13 6 13 15 7 13 15 3 9 1 2
2 0 9
7 16 15 3 9 13 13 2
3 15 13 3
12 13 15 11 9 13 2 16 13 13 9 0 2
5 9 15 1 13 2
15 10 9 9 13 3 9 13 11 11 11 9 12 9 12 2
13 15 0 9 13 10 9 13 9 0 9 1 9 2
4 13 15 15 2
4 13 15 3 2
13 9 3 13 9 13 3 13 0 9 0 3 9 2
8 3 15 13 13 9 13 9 2
3 0 9 15
5 13 3 15 0 9
8 13 15 2 16 13 13 13 2
4 9 0 13 2
6 9 13 9 7 13 2
3 9 13 9
5 13 13 15 3 2
3 6 3 2
13 13 3 13 2 16 0 0 9 15 13 3 9 2
10 9 13 13 3 13 2 9 13 0 2
6 11 11 13 3 9 2
9 0 3 13 9 2 10 3 13 2
10 13 10 9 7 9 3 15 3 13 2
14 0 9 13 13 9 3 9 2 16 3 13 3 9 2
11 15 13 12 3 0 9 2 9 7 15 2
3 9 3 2
16 12 9 13 9 1 3 12 9 13 0 9 9 12 12 9 2
17 8 8 8 2 13 7 13 2 15 10 9 7 9 9 9 13 2
5 15 13 13 9 2
5 3 9 9 13 2
5 13 0 9 3 2
7 9 13 9 12 9 1 2
7 3 0 9 13 0 9 2
11 13 9 3 2 16 13 13 3 13 9 2
4 6 15 15 2
12 13 3 0 2 16 15 13 13 13 0 9 2
14 11 11 13 13 9 2 15 15 13 7 13 9 9 2
2 9 9
5 15 13 3 9 2
10 9 13 3 0 13 3 16 13 3 2
5 0 9 13 3 11
4 13 11 9 2
5 9 13 11 9 2
4 9 13 9 1
17 9 13 3 9 9 15 13 15 0 16 15 2 13 3 16 15 2
5 3 13 9 0 2
18 0 13 9 0 9 2 0 15 13 3 13 10 9 13 2 11 13 2
8 11 13 3 10 0 0 9 2
15 13 11 3 3 13 9 3 3 16 13 15 13 9 0 2
4 13 13 13 2
4 15 13 0 13
9 15 13 3 0 3 10 9 9 2
2 9 9
7 9 13 0 0 7 13 2
15 2 3 13 2 16 2 2 10 9 9 13 9 13 9 2
5 11 7 11 9 13
13 9 13 15 9 9 2 13 15 3 2 13 15 2
24 15 13 16 15 7 13 13 9 10 9 7 16 10 11 13 13 3 13 3 3 13 15 3 9
4 13 3 3 2
5 15 13 0 9 2
12 10 9 16 11 13 13 0 9 2 13 11 2
10 15 13 9 9 2 15 1 13 9 2
20 9 13 13 3 10 9 2 3 9 13 13 7 15 13 13 3 3 12 9 2
17 13 13 13 3 10 10 9 16 13 3 13 3 3 0 9 3 2
5 9 13 13 13 2
16 11 9 13 13 9 9 2 16 11 9 3 12 9 13 9 2
5 11 13 13 11 2
14 11 11 11 12 13 0 9 13 11 11 9 1 12 2
5 0 13 13 13 2
13 11 13 0 9 13 0 0 7 0 9 0 9 2
11 13 13 3 13 7 13 2 13 3 3 2
11 11 13 3 11 2 3 9 9 9 9 2
7 9 15 13 3 0 9 2
14 16 9 15 1 13 13 1 9 2 13 9 11 9 2
9 9 13 0 13 3 3 0 9 2
13 11 13 9 9 0 9 2 15 9 9 13 13 2
8 15 13 13 13 15 3 3 2
5 15 1 13 9 2
6 13 3 16 0 13 2
5 15 13 9 9 2
8 15 13 9 13 0 0 9 2
6 13 9 2 9 13 2
5 9 13 0 9 2
15 13 15 13 3 2 2 3 9 13 13 9 9 9 2 2
5 13 13 9 3 2
6 9 13 10 10 9 2
4 3 12 13 11
4 9 13 9 2
9 16 9 13 9 2 13 0 9 2
8 10 0 9 11 9 11 13 2
6 13 3 12 9 9 2
2 0 9
6 16 13 10 10 9 13
3 13 9 2
5 13 3 9 15 13
9 3 13 3 3 10 0 3 3 2
7 9 8 7 0 9 7 9
6 9 10 9 2 13 2
7 9 13 9 9 0 9 2
6 15 13 16 13 9 2
13 16 9 13 13 3 2 15 9 9 13 9 1 2
6 9 7 11 13 9 2
6 3 15 13 13 11 2
39 15 13 10 11 0 9 3 10 9 16 15 13 11 3 11 13 15 13 3 3 3 10 0 3 0 9 10 0 3 9 1 16 15 13 15 13 10 9 2
4 0 0 0 9
11 0 9 13 3 0 2 3 15 15 13 2
8 9 13 9 9 11 11 11 2
12 9 9 13 9 13 3 13 13 9 7 9 2
7 3 9 13 13 12 9 2
8 9 13 0 16 8 11 13 2
14 16 15 13 9 9 2 3 15 13 13 15 0 9 2
6 15 13 9 12 9 2
7 10 15 13 9 10 9 2
5 15 13 11 1 2
10 9 13 9 9 9 13 9 10 9 2
22 11 13 3 2 7 13 13 3 2 9 13 9 2 7 13 9 16 10 9 13 9 2
11 13 9 9 13 2 16 15 13 9 1 2
11 9 13 3 0 9 2 15 13 3 3 2
11 3 9 1 13 9 13 11 3 3 12 2
5 12 9 13 9 2
11 15 13 3 3 12 9 3 16 13 15 2
13 10 9 13 3 9 1 7 3 9 13 9 12 2
6 9 13 9 1 0 2
5 13 3 3 13 2
10 0 9 3 11 13 9 9 13 9 2
7 9 13 9 3 9 9 2
5 13 0 13 0 2
16 16 9 13 9 13 13 13 3 2 9 13 9 13 13 9 2
11 16 13 3 13 2 16 3 13 13 11 2
10 9 13 9 1 11 11 13 9 1 2
10 13 9 2 16 13 13 15 9 13 2
4 9 13 9 13
12 13 16 9 7 9 13 0 7 13 0 9 2
8 11 9 13 9 7 9 3 2
3 15 13 2
5 15 13 0 9 2
5 13 3 3 9 2
6 6 9 9 16 15 13
5 3 13 13 13 2
8 10 12 9 11 13 11 9 2
2 0 9
2 6 9
6 9 13 9 13 9 2
7 11 9 13 3 0 9 2
8 9 11 13 13 3 0 9 2
4 9 13 3 2
3 9 13 0
4 9 13 9 2
8 13 0 9 12 9 15 1 2
12 9 9 13 12 9 13 9 9 1 3 0 2
5 15 3 13 9 2
5 15 13 9 0 2
2 9 9
10 3 3 0 9 0 9 7 3 13 2
3 13 13 13
9 10 0 9 15 13 3 9 13 2
4 13 15 7 2
4 9 1 13 9
3 3 1 9
6 3 13 7 3 13 2
6 10 9 15 13 9 2
9 13 11 9 2 15 13 3 9 2
19 10 9 11 13 13 9 9 9 3 9 2 16 9 9 13 13 13 3 2
15 9 13 13 2 16 13 9 13 7 15 13 13 13 9 2
3 9 13 13
3 9 13 13
19 16 9 13 10 9 10 9 13 9 9 7 10 3 9 13 0 0 9 2
6 0 13 3 3 9 2
9 13 3 15 2 15 13 9 3 2
12 3 2 15 3 13 13 16 13 10 9 13 2
6 13 3 2 13 13 2
8 13 16 15 13 3 3 0 2
12 10 9 15 13 9 9 12 9 12 9 1 2
9 11 16 13 11 9 3 13 9 2
9 13 3 9 2 9 13 13 9 2
10 9 11 13 9 9 13 11 13 9 2
8 9 13 3 0 13 0 9 2
4 10 12 0 9
12 3 13 3 13 9 9 7 13 0 9 3 2
3 9 0 9
4 15 15 13 2
8 9 13 9 7 9 13 3 2
9 15 13 13 0 9 13 15 0 2
10 8 7 9 13 13 9 11 1 9 2
9 3 3 0 9 13 13 0 9 2
7 9 9 13 9 0 9 2
3 0 0 9
4 13 10 9 2
7 11 11 13 11 10 9 2
11 3 15 13 13 11 12 9 10 9 9 2
5 9 13 9 13 9
5 15 13 11 1 2
7 16 9 0 13 15 13 2
5 13 15 0 15 2
9 9 13 13 9 10 9 13 9 2
14 10 15 9 13 15 2 16 15 13 13 3 0 9 2
9 9 13 9 0 9 3 13 9 2
2 9 1
5 9 1 9 13 2
8 0 13 2 16 9 13 9 2
4 9 13 0 2
19 9 13 3 0 9 2 12 9 9 13 13 13 2 3 9 13 13 9 2
9 3 9 13 13 13 9 9 3 2
5 13 13 0 3 2
5 6 2 13 15 2
7 9 1 13 13 10 9 2
9 9 1 13 9 3 13 13 9 2
7 10 9 13 13 3 13 2
10 12 9 9 13 13 13 12 9 9 2
8 0 9 9 9 13 3 11 2
2 10 9
3 0 0 9
8 13 13 12 11 9 0 9 2
5 12 13 3 13 9
14 11 9 13 13 10 0 2 0 2 7 3 10 0 2
6 9 13 3 9 2 9
9 0 9 13 13 9 9 3 3 2
5 9 13 0 9 2
4 13 3 13 2
6 9 13 15 13 3 2
10 15 13 16 15 13 3 3 3 13 2
7 9 9 13 3 3 0 2
8 13 15 13 2 15 13 13 2
2 13 9
10 6 3 3 3 16 13 15 0 3 2
20 13 9 12 2 12 7 10 15 2 15 13 2 16 9 13 0 2 11 13 2
10 13 10 9 13 13 9 2 11 13 2
4 15 13 3 0
14 11 15 13 13 2 7 3 2 15 13 13 0 9 2
3 9 12 9
10 11 13 13 9 2 13 10 10 9 2
4 13 15 3 2
5 13 11 13 3 2
6 9 13 13 15 13 2
10 13 9 0 9 2 16 13 15 3 2
12 9 2 11 7 9 13 9 13 9 2 16 2
5 9 13 13 9 3
10 3 9 7 10 10 9 13 13 9 2
5 9 13 3 13 2
11 13 3 0 2 16 0 9 13 3 3 2
4 11 13 9 0
7 9 15 13 3 9 1 2
12 9 9 13 13 3 3 11 9 13 9 1 2
14 9 13 10 0 9 2 15 15 13 13 9 1 13 2
4 15 13 3 2
3 0 0 9
10 13 15 13 10 0 9 3 13 3 9
9 13 13 9 9 9 13 10 0 2
7 9 13 9 7 13 9 2
7 15 13 15 9 9 1 2
10 10 9 1 9 13 0 9 13 9 2
17 3 0 2 15 13 3 3 13 2 13 13 3 10 9 9 1 2
7 11 13 2 9 15 13 2
2 0 9
7 7 3 15 13 15 13 2
19 3 13 10 9 2 15 13 0 7 0 2 13 10 9 13 13 3 15 2
37 15 13 9 7 9 2 15 13 13 15 7 15 13 9 1 15 2 13 15 9 2 9 2 9 2 9 2 9 2 9 2 9 7 0 9 9 2
8 13 11 3 7 3 2 15 13
6 9 13 9 0 9 2
8 9 13 9 16 9 9 9 2
11 10 9 13 13 0 2 7 15 13 0 2
18 9 13 9 9 7 9 1 2 15 1 15 13 0 13 13 9 9 2
7 13 2 13 15 13 3 2
15 2 13 13 0 0 9 2 16 9 13 13 3 0 2 2
11 15 13 9 9 9 2 13 11 9 9 2
5 15 15 13 3 2
15 15 3 13 13 9 7 12 2 7 15 13 13 9 9 2
11 16 0 9 13 3 9 7 13 9 9 2
16 3 11 13 13 9 9 0 9 2 3 13 2 16 13 9 2
16 15 13 13 11 1 10 9 16 15 13 2 13 15 3 3 2
13 11 9 13 12 7 0 2 15 13 13 9 1 2
7 15 15 13 0 0 9 2
16 9 13 0 9 13 13 3 9 9 13 15 13 3 0 3 2
16 16 15 3 13 13 10 12 9 9 1 2 15 13 3 13 2
9 15 13 15 15 13 2 9 9 2
18 16 15 9 3 13 10 9 3 9 13 2 11 2 9 7 15 3 2
9 11 9 11 13 9 13 13 9 2
3 13 15 2
9 13 3 9 1 7 15 13 3 2
24 16 3 9 13 2 3 3 2 12 9 9 3 2 3 15 2 3 13 3 2 0 9 0 9
5 15 13 9 9 2
12 3 0 13 2 16 9 9 9 13 9 9 2
3 15 13 15
9 3 9 13 11 9 13 9 9 2
5 3 15 13 3 2
12 15 13 13 9 9 1 9 2 13 3 9 2
6 9 0 9 13 9 2
8 9 0 9 13 13 3 0 2
13 13 13 2 16 10 11 9 3 0 9 13 9 2
4 11 13 11 9
2 9 11
3 8 7 9
18 3 3 13 3 2 13 16 9 13 3 13 7 13 9 2 3 9 2
5 13 3 10 9 2
12 9 13 13 9 13 3 2 16 15 13 9 2
4 9 13 9 3
12 12 9 15 13 13 9 3 7 13 9 3 2
4 7 10 9 2
4 10 12 0 9
3 11 11 9
7 7 13 10 9 13 9 2
8 9 13 3 12 9 1 9 2
6 15 13 9 0 9 2
21 11 11 9 13 9 1 2 7 11 13 0 9 10 0 2 16 13 13 9 1 2
3 15 13 13
18 11 9 13 13 2 3 9 2 3 0 9 2 7 11 13 3 0 2
3 13 12 9
8 11 13 2 16 13 13 9 2
5 15 13 3 13 2
5 15 13 15 9 2
3 9 13 3
5 9 13 9 9 2
9 13 3 13 10 9 2 11 13 2
3 13 3 0
2 13 13
2 13 13
4 9 13 0 9
21 15 13 7 15 13 2 13 13 2 7 15 13 3 0 9 16 13 13 12 9 2
4 2 13 3 2
15 9 9 13 15 0 2 16 15 13 0 9 3 16 0 2
5 9 13 3 13 2
5 6 2 13 10 9
4 9 13 0 2
9 9 13 3 0 3 10 0 9 2
10 9 0 9 13 3 0 9 11 13 2
15 0 9 9 13 9 9 2 3 9 7 9 13 13 9 2
8 15 13 13 3 13 9 9 2
3 9 13 13
7 15 13 3 9 9 9 2
6 13 10 9 3 0 2
4 3 3 9 2
15 11 13 3 2 15 13 9 0 2 9 2 9 7 9 2
4 15 13 3 0
4 13 13 9 2
7 13 13 3 12 9 9 2
12 9 1 9 13 13 10 15 3 9 13 1 2
2 13 9
8 7 3 3 13 13 15 3 2
5 9 13 9 9 2
6 9 13 13 7 9 2
9 13 15 3 13 9 2 11 13 2
14 13 13 0 9 2 15 13 13 13 13 9 7 9 2
11 11 9 13 3 13 12 7 11 3 12 2
7 9 13 3 12 9 3 2
24 10 9 13 13 2 16 3 0 9 13 0 13 9 3 7 9 3 2 16 3 9 13 13 2
10 15 13 2 16 9 13 3 3 9 2
23 9 13 13 13 2 13 7 13 2 16 15 15 1 13 9 2 9 7 10 9 13 9 2
8 15 13 9 2 9 7 9 2
28 16 9 13 3 12 9 2 0 2 0 2 0 2 11 11 13 0 2 16 2 0 13 0 16 10 15 2 2
3 15 13 0
17 11 11 9 1 13 3 9 15 2 15 13 9 9 7 10 9 2
12 16 9 9 13 9 9 2 3 9 13 0 2
8 13 13 13 2 16 13 9 2
15 7 15 13 13 2 16 9 15 15 13 13 15 3 13 2
10 9 13 13 9 10 9 2 13 11 2
10 9 11 9 9 13 3 12 9 12 2
8 3 15 13 3 3 13 15 2
14 8 8 8 8 8 8 8 2 11 13 0 0 9 2
5 7 3 13 9 2
9 11 9 13 3 13 3 3 0 2
13 16 9 9 13 3 2 13 9 7 9 3 9 2
18 16 15 13 13 13 16 15 13 3 9 2 3 15 13 3 3 3 2
13 15 13 13 9 13 9 2 7 9 9 3 3 2
10 9 11 11 15 1 13 9 1 9 2
7 15 13 3 16 15 13 3
3 15 13 11
11 9 13 9 1 13 3 7 3 1 11 2
4 9 9 11 11
15 11 13 11 9 16 13 9 0 16 13 11 9 13 9 2
11 13 9 7 15 13 15 13 9 7 9 2
9 9 9 13 7 15 13 9 1 2
6 9 13 13 13 9 2
13 0 9 13 3 0 2 16 13 0 7 9 13 2
4 9 13 9 2
11 11 9 9 9 9 9 13 3 9 13 2
2 0 1
11 13 11 7 13 3 9 9 3 10 9 2
20 9 9 11 13 3 15 2 13 15 3 3 0 9 16 3 11 9 3 13 2
3 15 13 2
12 9 13 13 9 2 3 3 13 10 9 9 2
6 11 13 13 13 3 2
13 2 13 13 2 15 13 13 3 15 2 11 13 2
19 11 13 9 11 2 7 13 3 3 13 11 2 7 9 13 13 0 9 2
11 13 15 13 11 2 15 9 13 9 9 2
4 13 15 13 2
5 10 12 9 13 3
11 9 9 13 3 0 2 16 13 3 0 2
15 15 1 16 13 9 0 9 2 13 9 12 13 0 9 2
13 15 13 3 3 3 9 1 12 13 3 10 9 2
14 0 13 13 15 2 16 11 13 9 13 0 9 9 2
14 9 13 3 0 2 9 13 13 0 16 15 3 13 2
11 9 1 9 13 15 2 15 13 9 3 2
4 9 13 13 9
7 11 13 9 3 9 3 2
8 13 15 3 2 9 13 13 2
5 9 13 9 0 2
11 0 13 15 2 16 13 9 9 9 13 2
11 15 15 13 13 2 13 13 7 13 9 2
8 13 16 13 3 9 9 13 2
6 0 9 13 3 9 2
7 3 13 3 13 11 9 2
13 9 13 9 2 15 3 12 0 13 3 9 9 2
30 11 13 9 1 0 9 9 2 15 15 13 9 13 2 15 13 13 15 9 2 15 15 2 0 9 2 13 0 9 2
26 9 3 13 2 13 10 3 9 2 16 0 13 2 16 11 9 13 10 9 2 10 9 9 1 13 2
2 13 9
9 9 13 0 7 9 13 13 3 2
42 3 15 13 10 0 2 9 2 16 12 3 13 3 16 10 9 2 10 3 0 16 12 9 13 0 9 13 9 9 7 9 9 9 2 16 3 15 13 10 9 13 2
12 11 9 9 13 9 9 9 11 11 9 1 2
12 15 13 11 11 9 13 12 9 9 0 9 2
11 3 13 9 9 13 2 3 13 9 11 2
21 11 11 2 3 2 7 11 11 13 9 13 10 1 9 2 9 2 9 7 9 2
10 9 13 15 3 13 2 0 9 3 2
4 15 13 13 2
17 3 13 13 13 0 15 2 13 10 9 9 9 9 7 9 9 2
7 9 13 9 1 9 9 2
5 13 13 9 9 2
2 10 9
7 9 9 13 13 9 0 2
14 13 0 9 7 3 9 3 13 10 9 7 0 11 2
13 3 10 9 13 13 9 2 7 15 13 13 11 2
7 15 13 0 9 9 13 2
5 13 11 12 9 2
2 9 13
6 3 9 13 15 13 2
4 6 3 0 2
4 9 13 3 3
6 15 13 3 3 9 2
4 3 13 9 2
6 9 11 13 0 9 2
4 0 9 9 13
2 11 9
16 9 2 9 7 9 13 13 3 2 16 10 0 9 13 9 2
10 9 13 2 16 13 15 13 9 2 2
12 9 13 3 3 9 13 7 9 10 9 13 2
8 0 11 9 13 13 9 12 2
14 16 9 13 7 13 2 15 13 9 2 13 13 11 2
3 9 0 9
11 15 15 13 0 9 2 15 15 13 0 2
10 15 13 15 2 16 9 13 13 0 2
4 13 15 9 2
6 10 9 15 9 13 2
11 3 9 13 13 9 2 13 0 3 13 2
6 3 0 13 0 9 2
10 9 13 3 0 9 2 3 0 9 2
5 15 13 9 1 2
3 3 13 2
11 9 12 11 13 7 9 16 0 9 9 2
30 6 2 3 7 3 13 13 0 9 16 15 13 13 9 2 3 2 6 3 2 16 9 1 13 3 10 0 9 7 2
5 13 3 9 1 2
16 7 11 13 11 0 0 9 2 0 2 15 11 13 3 13 2
16 3 16 15 13 0 9 16 13 15 13 15 15 13 10 15 2
10 13 15 0 9 2 15 13 10 9 2
5 9 13 13 9 2
4 3 9 13 2
3 13 9 12
17 16 13 15 2 3 13 15 3 2 16 9 13 3 3 13 9 2
4 9 13 15 9
6 6 15 15 3 13 2
10 11 0 9 13 3 12 12 9 13 2
2 11 9
9 9 13 9 7 9 13 16 9 2
8 15 13 0 7 0 0 0 2
12 10 9 13 13 11 0 9 9 13 9 9 2
2 0 9
10 9 13 9 13 9 9 1 0 9 2
7 0 9 13 9 9 9 2
7 9 7 9 13 0 13 2
10 9 13 10 9 12 9 7 15 3 3
14 2 9 2 13 0 13 2 16 10 9 13 13 3 2
8 13 2 7 11 3 13 9 2
10 9 9 9 13 13 3 15 3 9 2
5 2 6 15 15 2
12 3 3 9 13 2 3 0 9 13 7 13 2
6 15 13 3 9 9 2
5 9 13 9 0 2
7 9 13 9 1 10 0 9
7 15 13 3 9 7 9 2
9 3 13 0 9 9 2 13 11 2
5 13 9 13 9 2
6 10 9 9 15 13 2
7 9 13 13 3 12 9 2
28 3 9 9 13 13 3 0 9 2 7 16 15 13 10 9 13 2 13 15 3 3 3 13 2 3 0 9 2
13 9 9 3 13 2 7 9 13 13 12 9 11 2
3 13 13 2
15 11 13 13 13 9 15 13 9 9 9 9 12 11 9 2
17 15 13 0 9 16 3 13 9 10 11 16 15 13 13 10 9 2
6 9 13 3 9 1 2
14 9 13 13 3 0 3 2 10 9 13 0 13 3 2
5 15 13 0 13 15
12 13 3 0 9 9 7 16 13 13 0 9 2
3 3 3 3
2 0 9
12 13 9 13 3 13 7 13 3 9 13 9 2
3 13 13 2
5 11 13 11 3 2
10 9 13 9 7 13 9 13 0 9 2
11 9 0 0 9 13 9 11 13 13 9 2
6 15 3 3 13 10 9
11 3 9 9 9 13 13 3 15 9 13 2
10 9 13 13 13 9 2 7 3 9 2
13 15 13 9 2 15 3 0 7 0 9 13 9 2
11 9 13 9 13 13 13 3 3 9 1 2
3 2 11 2
12 9 2 3 0 9 13 13 9 13 9 9 2
6 9 9 13 0 9 13
14 13 3 15 2 16 13 0 0 9 9 2 7 3 2
14 16 10 9 13 2 16 9 13 12 3 2 3 13 15
17 13 13 3 0 13 2 3 7 3 0 9 13 0 13 0 9 2
8 3 13 0 9 16 13 13 3
4 13 10 0 2
10 11 9 13 9 9 16 13 0 9 2
13 16 13 3 13 2 13 8 8 3 0 0 9 2
10 13 13 1 9 2 15 1 7 1 2
8 16 11 13 0 2 15 13 2
3 9 13 2
2 13 13
5 15 13 10 9 2
6 13 9 3 0 9 2
9 9 9 13 3 3 0 16 13 2
6 11 13 3 10 9 2
3 13 9 1
4 13 9 13 2
10 13 0 16 13 13 3 0 9 13 2
5 13 3 0 11 2
6 9 13 13 3 9 2
7 10 9 9 13 12 9 2
11 0 13 13 13 2 16 9 13 3 13 2
3 12 9 13
4 15 13 3 2
4 12 9 9 11
4 15 11 13 2
10 15 13 13 3 0 3 10 9 9 2
8 15 13 10 9 3 12 9 2
8 9 9 9 9 13 13 9 2
2 10 9
12 11 1 10 9 9 13 3 12 12 9 9 2
7 13 3 9 7 13 0 2
3 9 9 2
10 0 13 0 9 3 3 10 9 1 2
14 0 15 13 2 7 13 3 10 9 16 10 9 13 2
4 9 13 13 2
4 11 9 0 9
11 13 3 3 2 16 9 13 3 3 3 2
21 7 9 13 10 9 3 3 2 16 9 13 13 9 2 16 15 13 9 13 9 2
6 9 13 0 9 9 2
5 13 9 7 13 15
11 13 9 9 2 3 9 2 9 13 13 2
13 10 9 2 9 11 2 9 13 13 10 0 9 2
9 15 13 3 9 2 13 9 3 2
7 13 15 2 15 7 15 2
5 11 9 13 15 2
12 13 13 10 9 9 13 2 7 3 15 13 2
15 9 13 9 3 3 7 15 1 13 9 2 13 9 9 2
10 3 0 9 13 3 13 13 13 9 2
6 13 9 13 3 9 2
6 13 9 0 9 13 2
6 15 13 13 13 9 2
2 9 9
7 3 9 7 9 13 9 2
22 9 9 9 11 13 7 13 0 9 2 13 9 7 13 9 2 15 9 13 9 11 2
7 3 15 13 3 13 15 2
11 11 9 13 13 9 13 16 12 9 11 2
14 15 13 13 11 2 11 2 11 2 11 7 3 3 2
12 15 13 13 13 7 13 3 9 7 10 9 2
9 11 13 13 2 7 15 13 15 3
6 11 13 0 0 9 2
15 13 3 3 0 9 2 15 13 3 2 16 13 13 9 2
6 15 13 3 0 9 2
8 13 13 9 7 10 10 9 2
3 0 9 2
7 9 13 3 3 3 9 2
6 15 15 13 3 9 2
10 13 9 1 2 15 13 9 10 9 2
12 11 13 9 3 7 13 0 9 9 9 16 9
7 2 3 3 13 3 2 2
20 11 7 11 0 9 13 0 9 15 2 3 12 15 13 9 13 13 15 15 2
6 9 9 9 13 0 2
2 10 9
14 13 3 0 10 9 13 13 0 9 9 0 9 9 2
4 15 13 3 3
24 10 9 9 9 9 3 3 7 11 13 13 3 13 3 15 13 3 7 13 16 13 15 13 2
5 13 9 13 9 2
8 11 13 16 9 13 3 9 2
12 9 13 9 7 9 0 2 0 2 0 9 2
3 13 9 9
13 9 9 13 9 2 16 3 8 7 0 9 13 2
10 15 13 15 2 15 7 9 7 9 2
13 15 13 15 2 16 9 7 11 9 13 3 3 2
7 9 13 13 12 9 9 2
14 15 13 9 7 13 2 6 9 1 2 11 15 3 2
3 15 13 13
5 15 15 13 9 2
5 13 3 10 9 2
12 3 16 11 13 2 3 13 0 9 13 9 2
4 9 13 9 2
13 16 9 13 3 16 9 2 9 13 9 0 0 2
8 13 13 11 2 10 9 9 2
13 15 13 3 3 9 7 13 3 3 3 3 3 9
5 9 13 9 9 2
8 13 3 10 9 13 15 1 9
14 9 13 9 9 7 15 9 2 13 9 7 13 9 2
10 15 13 0 13 2 13 0 16 9 2
16 11 13 9 2 13 9 0 9 13 11 9 7 13 9 11 2
6 3 10 9 13 13 2
13 9 13 2 16 11 13 13 3 0 9 13 3 2
5 13 11 0 9 2
8 9 3 13 13 13 10 9 2
15 9 13 9 3 9 1 7 13 9 7 13 16 13 3 2
9 11 13 13 3 9 7 9 3 2
14 3 15 3 9 9 9 2 15 3 13 0 0 9 2
7 15 13 9 3 13 9 2
17 10 0 9 13 13 13 2 16 11 15 13 10 9 13 0 9 2
9 10 9 11 13 13 9 9 1 2
7 11 13 2 13 13 9 2
7 9 16 13 15 13 13 2
29 7 3 15 13 3 3 3 1 10 0 0 9 3 3 3 13 0 9 7 9 7 9 3 16 15 13 13 3 15
5 11 13 15 9 2
4 9 13 9 9
18 9 13 2 16 8 7 9 13 3 15 2 15 13 3 12 9 9 2
7 9 13 3 0 13 9 2
13 9 13 0 9 2 16 13 0 13 13 3 3 2
3 9 13 9
3 3 13 9
16 13 11 1 7 13 9 3 3 16 9 2 9 7 9 3 2
16 3 13 13 13 3 2 7 13 13 13 16 9 13 3 3 2
7 3 15 13 13 13 13 2
2 9 9
2 0 9
9 15 9 13 2 13 9 3 3 2
11 6 3 2 10 15 13 13 9 0 9 2
13 15 13 13 13 15 2 15 13 13 13 3 15 2
20 7 3 3 2 13 12 9 3 3 7 3 13 10 9 9 1 2 3 7 2
6 3 3 9 13 0 9
10 15 13 13 13 9 2 7 13 13 2
8 10 12 9 13 13 0 9 2
10 13 0 2 0 9 10 9 9 1 2
2 6 0
6 13 15 15 7 11 2
14 9 13 13 13 9 13 0 9 13 13 3 0 9 2
12 3 9 13 15 9 1 13 15 1 13 9 2
8 15 13 16 15 13 10 9 2
7 11 13 13 0 10 9 2
6 9 13 0 12 9 2
2 13 3
5 2 7 13 13 2
14 11 11 13 9 3 3 2 13 9 13 3 9 0 2
17 15 13 3 10 9 2 16 9 13 13 3 10 12 9 3 3 2
9 11 13 9 7 13 9 11 3 2
3 11 13 11
12 15 13 13 2 3 9 13 15 2 0 0 2
5 15 13 13 9 2
9 11 13 3 13 13 3 11 11 2
15 9 13 11 9 7 13 15 9 2 10 9 13 0 9 2
6 9 13 13 3 0 2
17 9 13 3 9 7 3 13 2 16 13 13 0 0 9 11 9 2
12 9 15 13 15 9 2 3 15 3 9 13 2
7 3 15 13 9 1 3 2
4 9 13 0 2
17 16 13 13 9 9 13 7 13 9 2 13 13 9 13 3 9 2
17 11 2 12 2 13 0 9 10 15 2 15 13 1 9 9 9 2
7 15 13 9 3 15 13 2
6 9 13 13 2 9 2
4 2 9 0 2
8 9 11 13 12 0 9 9 2
7 12 9 13 9 1 9 1
16 13 13 2 16 15 13 9 12 9 1 2 16 9 13 0 2
18 7 9 13 3 2 7 3 13 2 7 3 9 13 2 7 15 13 2
6 11 13 3 0 13 2
8 13 0 2 11 2 13 13 2
6 9 13 7 13 0 2
15 13 13 2 16 10 9 13 13 2 7 13 13 2 15 2
2 13 9
6 11 1 13 13 9 2
4 13 3 3 13
3 13 3 13
3 13 15 2
6 13 9 9 13 9 2
3 9 13 13
2 0 9
9 11 13 10 9 13 3 0 9 2
16 15 13 3 15 13 13 15 7 15 1 7 13 9 7 15 2
3 13 15 2
23 9 2 9 2 13 3 9 0 9 2 15 3 13 3 12 2 16 3 0 9 0 9 2
6 15 13 12 9 9 2
6 3 15 13 13 13 2
5 15 13 13 13 9
6 3 9 13 3 9 2
4 9 13 9 2
6 11 13 9 1 9 2
16 13 13 2 16 13 13 2 7 15 13 15 13 3 9 9 2
6 7 13 15 13 13 2
6 15 13 3 9 3 2
13 9 13 13 3 3 2 1 9 15 13 13 15 2
11 7 16 10 9 3 13 2 3 15 3 2
12 11 9 13 13 9 2 0 11 13 3 3 13
6 15 13 9 3 0 2
4 13 3 9 2
4 0 9 15 1
5 13 15 11 3 2
12 15 15 13 13 0 9 2 13 3 3 9 2
19 10 9 13 2 16 13 15 13 10 9 2 16 15 13 13 15 1 9 2
6 15 13 3 3 3 2
7 3 2 11 13 13 9 2
4 15 3 13 2
9 15 13 3 0 0 3 0 9 2
5 15 13 3 9 2
5 3 0 15 13 2
7 13 11 9 7 13 3 2
4 15 13 13 2
13 0 9 13 13 0 2 13 10 9 3 0 13 2
5 9 9 13 9 2
11 10 9 9 1 13 11 11 13 11 9 2
4 13 13 1 9
15 15 3 13 10 9 3 3 16 15 13 16 13 0 13 2
3 15 13 2
7 15 13 13 3 10 9 2
22 3 13 13 11 0 9 7 3 15 1 13 13 0 9 2 16 15 10 9 3 13 2
7 0 9 13 13 0 9 2
6 11 0 9 13 11 2
9 9 9 13 9 13 9 3 9 2
8 9 7 9 13 13 0 9 2
7 13 13 0 9 13 9 2
9 9 13 13 0 3 16 9 1 2
6 11 13 3 13 9 2
8 9 13 13 13 3 10 12 2
15 9 13 9 9 0 9 0 7 13 15 9 7 9 1 2
2 11 9
13 6 15 15 13 2 16 13 15 13 10 0 3 2
4 13 13 13 2
5 15 15 13 13 2
9 6 2 13 15 3 13 2 7 2
3 0 15 13
7 13 13 10 13 9 1 2
7 11 7 11 9 13 15 2
10 9 13 9 1 3 13 0 13 9 2
16 9 13 13 10 9 7 10 9 9 2 7 9 13 13 0 2
5 0 9 13 3 2
2 9 9
11 11 1 13 0 9 16 15 15 15 13 2
2 13 3
10 15 13 13 9 9 0 2 0 9 2
16 9 9 13 0 9 2 15 9 9 1 13 9 7 9 9 2
9 13 2 16 9 13 0 13 13 2
4 9 13 0 2
16 9 15 13 0 2 3 15 13 13 13 13 9 7 9 1 2
14 3 2 9 11 2 13 11 13 2 16 11 9 13 2
7 13 9 3 12 9 7 2
7 3 3 13 0 9 15 2
8 10 9 1 9 13 3 0 9
4 0 8 7 9
6 13 15 13 15 15 2
2 13 9
16 7 15 16 13 0 9 13 3 15 16 9 13 9 0 9 2
3 3 13 9
11 10 0 13 13 9 15 13 13 10 9 2
11 9 13 3 3 2 7 9 13 0 3 2
12 16 13 13 9 2 13 15 0 3 9 1 2
7 15 13 3 13 13 15 2
2 9 9
11 0 9 9 13 9 13 3 9 0 9 2
11 9 9 1 0 9 13 9 13 2 16 2
6 10 9 13 13 9 2
3 11 0 9
15 0 9 11 11 13 3 2 9 15 1 13 15 0 9 2
13 15 13 9 13 13 9 2 15 13 13 9 3 2
7 9 11 13 3 0 9 2
8 7 3 13 10 9 15 15 13
15 0 13 2 16 0 9 11 13 12 9 9 1 0 11 2
22 9 2 16 9 7 15 13 13 7 13 9 2 9 2 9 2 9 2 2 13 0 2
20 15 1 11 9 13 9 13 2 13 7 9 13 3 11 3 11 7 11 13 2
16 16 13 0 9 13 9 2 13 15 13 15 13 2 11 13 2
10 11 9 13 9 2 11 13 9 13 2
5 11 13 13 9 2
11 10 9 16 15 13 0 9 2 7 13 2
10 11 13 13 11 3 9 15 0 9 2
2 0 9
2 13 13
4 15 13 0 9
5 9 9 7 9 1
12 16 9 13 0 2 15 13 13 9 7 9 2
15 13 9 3 2 13 9 9 2 7 9 13 13 3 9 2
7 11 7 11 13 0 9 2
4 9 13 9 2
15 15 13 7 3 13 9 0 9 2 2 13 2 0 9 2
15 9 13 11 13 2 16 9 13 3 9 0 9 9 9 2
14 15 13 13 9 2 3 9 9 9 13 3 9 1 2
6 3 13 15 0 9 2
8 13 13 3 16 13 13 13 2
3 3 13 2
4 9 13 3 2
2 3 0
5 13 3 0 9 2
6 9 9 13 9 0 2
5 13 15 3 9 2
6 15 13 0 9 0 2
14 13 2 9 3 13 16 2 15 15 3 13 0 9 2
9 0 9 13 3 13 9 13 9 2
7 13 15 13 9 13 9 2
4 15 13 9 2
11 9 9 13 16 15 3 13 13 15 3 2
5 16 3 13 15 2
25 9 9 13 13 2 16 9 13 13 7 16 9 13 3 9 7 16 9 13 3 0 2 3 0 2
7 3 10 9 13 13 13 2
14 16 9 1 13 10 0 2 0 15 2 0 9 13 2
15 9 13 9 0 9 9 2 7 15 13 13 3 12 9 2
2 6 15
2 0 9
2 0 13
10 13 15 13 3 0 9 7 9 9 2
10 0 9 1 9 13 0 9 0 9 2
12 16 0 13 2 9 13 3 13 12 9 3 2
7 9 13 9 3 0 9 2
6 0 9 13 15 3 2
5 9 7 9 13 9
4 9 7 9 9
10 0 12 0 0 9 13 3 0 8 2
9 13 3 3 2 16 9 13 0 2
3 13 9 9
5 13 9 9 13 2
6 13 15 3 16 11 13
26 11 2 11 11 13 12 11 9 9 2 3 15 13 11 9 2 13 3 2 16 0 9 13 3 9 2
9 13 0 13 2 15 0 13 13 2
11 11 13 13 9 2 13 15 3 13 9 2
5 9 13 9 13 2
9 13 3 13 2 16 9 15 9 2
14 13 2 16 13 15 7 10 15 13 9 0 1 9 2
6 0 9 13 9 9 2
15 16 0 9 13 3 3 9 2 16 15 13 13 9 9 2
13 13 9 2 13 9 9 9 2 16 15 13 9 2
22 13 16 3 15 13 12 0 9 16 15 3 13 3 9 15 15 13 13 3 8 10 9
10 9 13 9 13 2 13 7 13 9 2
9 7 2 15 13 3 2 3 3 2
8 13 13 9 9 2 3 9 2
11 11 13 9 0 9 2 7 3 0 9 2
18 9 13 2 16 9 13 13 9 7 13 10 3 0 9 2 3 9 2
11 9 13 2 16 10 9 13 15 3 13 2
7 9 9 13 9 0 9 2
8 11 13 3 9 3 0 9 2
7 11 9 13 3 9 11 2
7 11 13 9 9 3 3 2
7 9 13 3 3 11 9 2
8 13 9 2 3 0 2 13 2
5 13 15 3 3 2
19 16 13 13 3 2 16 9 9 13 2 13 9 9 9 7 9 13 3 2
5 9 13 9 11 2
10 9 2 16 0 0 9 13 3 10 15
11 13 3 2 16 13 13 13 15 1 9 2
6 15 13 13 3 13 2
7 9 13 7 13 13 9 2
21 16 9 13 13 3 2 3 10 3 0 9 9 13 9 13 13 10 0 9 0 2
3 13 3 3
8 3 13 15 13 9 13 9 2
4 9 13 15 1
8 10 9 9 7 9 13 9 2
8 3 11 13 12 9 13 9 2
10 15 13 9 11 7 15 9 11 9 2
10 15 13 13 2 16 15 13 10 9 2
4 13 13 13 2
10 3 15 13 13 16 3 9 13 3 2
5 10 10 9 9 2
10 15 13 10 0 3 2 3 9 13 2
12 9 13 13 9 2 7 15 13 3 13 9 2
4 6 15 7 2
11 9 3 0 9 13 8 2 8 7 9 2
5 13 15 0 9 2
5 11 13 3 9 2
11 11 13 13 13 9 2 7 13 15 13 2
11 9 3 13 9 9 9 2 15 3 13 2
4 13 3 13 2
10 9 13 9 2 10 9 13 15 13 2
6 11 11 13 10 9 2
6 3 15 3 9 13 2
3 0 9 11
7 15 13 9 13 0 9 2
4 15 13 3 2
4 9 13 0 9
11 3 13 0 9 13 2 9 13 9 0 2
10 3 13 13 9 0 9 2 3 0 2
8 11 13 13 9 9 1 9 2
7 13 12 9 9 9 13 2
9 13 13 9 2 13 9 3 3 2
8 15 13 3 9 3 0 9 2
5 9 13 13 9 2
13 15 13 13 9 13 9 2 16 13 0 9 9 2
7 9 13 7 9 13 3 2
12 15 13 3 0 9 2 16 13 13 15 0 2
7 9 10 9 13 13 9 2
7 9 15 13 3 10 11 2
6 15 13 13 13 9 2
7 9 13 0 9 11 11 2
8 9 13 9 10 9 0 9 2
10 15 13 3 9 7 15 13 3 9 2
12 9 9 13 9 2 3 9 13 12 11 9 2
16 13 9 12 9 1 2 15 1 13 9 13 9 3 0 9 2
4 13 12 1 2
7 9 13 12 9 3 16 13
10 13 15 2 15 9 13 3 13 0 2
7 9 13 13 9 13 9 2
7 15 15 3 13 3 9 2
18 2 11 2 12 7 2 11 2 12 9 9 13 13 15 3 9 9 2
32 16 15 13 9 9 2 15 13 8 8 1 7 13 11 3 9 2 3 3 3 1 12 2 16 15 13 13 11 1 3 9 2
13 9 13 13 3 15 2 16 9 9 9 13 9 2
7 10 9 13 9 13 11 2
5 13 13 0 9 2
3 9 0 9
14 9 11 11 1 0 9 9 13 0 13 3 0 9 2
7 9 13 13 11 0 9 2
5 9 13 10 9 2
7 11 13 3 0 9 9 2
8 9 13 9 13 9 0 9 2
6 3 11 9 13 0 2
12 12 9 13 13 12 9 7 3 12 9 9 2
11 3 13 3 9 2 16 9 13 9 1 2
14 10 9 13 10 9 2 16 15 13 8 7 15 9 2
3 12 0 2
4 11 13 9 2
9 9 0 9 13 2 16 13 9 2
15 0 2 0 7 13 9 13 7 15 13 2 16 9 13 2
10 0 9 13 9 9 7 0 9 9 2
5 10 9 13 13 9
4 15 13 9 2
4 11 12 9 1
12 3 11 7 15 13 2 16 15 13 0 9 2
8 3 3 2 16 15 13 15 2
3 13 9 2
8 15 13 9 13 13 0 9 2
7 16 3 0 9 9 13 2
8 10 10 0 13 9 13 13 2
15 3 16 9 13 0 9 2 10 9 13 3 3 13 9 2
3 13 13 9
5 9 13 13 12 2
3 9 13 13
6 15 13 9 7 9 2
5 15 13 16 3 2
13 10 9 2 15 13 13 3 13 13 3 9 3 2
7 9 9 13 7 9 13 2
8 9 0 9 13 9 9 1 2
14 0 9 13 0 0 9 2 15 13 3 3 9 3 2
7 3 3 15 13 13 3 2
9 15 13 3 9 9 9 9 9 2
9 11 13 3 9 2 15 1 13 2
8 13 3 9 9 10 9 13 2
7 15 13 13 9 9 9 2
9 13 9 9 13 9 0 16 3 2
6 13 13 15 9 11 2
10 9 13 3 13 9 9 9 13 0 2
23 13 15 15 13 16 15 13 11 2 7 15 15 13 13 13 13 16 13 15 13 15 3 2
7 13 15 3 3 13 15 2
12 7 3 3 13 9 3 0 9 2 9 9 2
8 7 3 15 13 10 9 13 2
15 9 13 9 3 3 9 7 9 13 9 9 7 3 9 2
2 0 9
15 15 13 13 13 0 9 9 9 7 3 13 13 15 9 2
6 9 13 9 9 1 2
7 13 11 13 3 3 3 2
18 11 11 9 9 13 10 9 9 3 9 2 16 9 13 13 9 9 2
5 15 13 15 1 2
3 9 9 13
23 16 11 7 15 13 13 9 11 7 11 9 12 2 10 9 13 13 0 15 15 13 3 2
6 0 12 12 9 11 2
12 3 13 9 13 0 7 0 2 7 13 0 2
22 9 9 9 9 13 13 0 2 0 9 15 13 9 9 11 13 9 2 9 9 2 2
6 9 13 15 3 3 2
14 13 16 15 13 3 9 1 13 9 2 9 13 13 2
4 15 3 13 2
11 3 16 9 0 9 13 3 3 9 9 2
8 13 13 0 9 2 3 13 2
5 15 13 9 1 2
7 13 3 0 16 13 3 2
13 9 13 3 3 2 11 3 13 9 3 10 3 2
12 13 3 13 9 2 16 15 13 13 9 9 2
7 3 15 13 0 7 0 2
6 11 9 13 10 9 13
8 9 15 13 13 12 0 9 2
7 10 9 13 11 9 9 2
9 11 2 11 2 11 2 11 7 11
5 15 13 0 9 2
2 11 9
17 11 2 11 2 7 11 2 11 2 13 0 9 9 2 9 1 2
6 13 10 9 9 9 2
12 11 13 11 9 3 9 9 11 13 0 9 2
12 11 9 13 3 0 13 9 16 9 3 9 2
11 9 13 9 7 11 13 3 9 7 9 2
24 0 9 13 9 2 13 9 1 7 3 3 9 9 1 10 0 9 1 2 0 16 13 3 2
66 15 13 3 0 16 2 15 9 13 13 3 15 13 0 9 0 8 2 9 9 16 3 0 9 2 9 9 7 3 2 3 3 3 15 15 13 10 9 15 13 13 13 3 10 12 9 7 15 13 13 3 2 3 10 0 9 16 2 16 13 13 3 3 3 13 15
7 9 13 9 13 13 2 2
16 9 13 13 13 9 3 2 7 15 13 13 2 9 7 15 2
19 15 3 0 9 9 13 2 0 9 0 9 11 13 13 15 15 9 9 2
17 10 9 3 13 9 1 10 9 3 11 7 11 1 13 0 9 2
9 6 13 15 13 3 16 11 9 2
24 9 9 13 3 0 0 9 2 15 13 10 9 0 9 2 15 1 9 13 13 3 13 15 2
6 9 9 13 0 9 2
5 0 9 13 13 9
8 9 9 10 9 13 9 0 2
10 11 15 13 9 9 11 1 3 9 2
6 9 13 13 12 9 2
2 12 9
3 9 13 13
3 13 15 2
15 11 9 2 3 15 2 13 13 3 0 9 11 9 13 2
10 11 13 13 7 11 7 11 0 9 2
11 11 9 13 9 13 9 13 9 0 3 2
3 15 13 13
16 9 13 3 9 0 9 2 15 13 3 13 11 0 9 1 2
5 9 13 12 9 2
9 10 9 9 13 12 12 12 9 2
9 0 0 9 1 11 13 13 0 9
5 13 15 3 13 2
6 10 9 13 3 11 2
5 13 10 9 3 2
8 3 9 13 13 2 3 13 2
2 13 13
6 3 13 13 9 7 9
11 9 1 13 9 13 13 9 3 9 12 2
4 15 15 13 2
6 9 9 13 13 13 2
7 11 13 10 9 0 9 2
8 13 15 3 10 9 10 11 2
5 15 13 9 1 2
6 6 16 13 15 3 2
14 7 13 13 9 7 13 3 2 16 9 13 0 13 2
8 10 9 9 9 13 9 0 9
8 9 13 13 0 9 0 9 2
12 9 9 13 0 9 3 16 15 13 0 9 2
17 10 9 13 15 2 13 13 12 2 12 2 12 7 15 9 9 2
6 12 15 13 16 15 13
6 0 13 3 0 9 2
17 3 0 9 13 13 13 3 0 9 7 15 13 3 13 0 9 2
11 16 13 3 2 16 13 13 12 9 0 2
5 13 9 13 0 2
9 9 13 13 9 13 15 3 9 2
8 3 3 13 9 9 13 0 2
4 13 9 9 2
6 9 11 13 13 9 2
14 9 13 2 16 11 13 10 9 9 7 13 15 15 2
8 11 1 11 13 3 9 9 2
8 9 13 13 9 0 0 9 2
6 6 13 9 3 9 2
6 9 10 9 9 13 2
22 9 13 9 2 15 13 0 2 10 9 13 13 2 15 13 9 7 15 13 13 9 2
8 6 10 15 15 13 9 13 2
21 15 3 13 13 3 10 9 2 7 10 0 9 13 3 11 2 3 2 3 3 2
8 9 11 13 13 9 9 9 2
8 10 9 13 13 9 13 15 2
7 13 9 13 13 0 3 2
7 10 13 9 13 10 9 2
9 13 15 13 15 7 13 3 13 2
3 6 11 2
7 9 13 3 3 9 9 2
10 0 9 13 3 13 0 9 13 16 0
10 3 0 13 9 13 0 3 9 9 2
17 13 3 2 3 15 13 3 3 15 13 3 13 15 13 3 3 13
6 3 9 13 15 13 2
11 11 13 9 3 7 13 15 3 3 3 2
5 13 2 16 13 2
6 13 7 13 9 9 2
4 10 9 13 15
23 15 11 13 13 9 0 9 9 2 3 3 0 7 0 9 13 13 2 9 2 0 9 2
8 9 13 3 0 9 2 11 13
8 15 13 9 7 13 3 9 2
5 13 15 15 13 13
13 12 11 9 13 15 2 16 11 13 9 11 13 2
6 9 13 13 13 3 2
8 3 0 13 9 3 9 15 2
9 1 11 9 0 9 9 13 9 9
2 13 13
15 3 15 13 9 9 2 15 13 3 13 16 15 13 3 2
5 15 13 13 9 2
11 15 1 9 13 13 7 0 7 3 0 2
12 9 13 2 16 9 9 13 3 10 9 1 2
11 10 9 13 0 2 16 15 13 9 13 2
10 12 9 9 13 13 9 13 9 13 3
6 9 13 13 9 1 2
6 15 13 3 12 1 2
13 9 1 9 9 7 9 3 13 11 9 12 9 2
12 13 15 13 13 13 15 15 1 16 11 13 9
14 15 13 13 3 0 9 1 7 3 10 0 9 1 2
13 13 13 9 3 16 13 13 15 9 7 9 1 2
6 0 9 9 13 0 2
12 9 13 9 13 13 9 0 7 0 13 9 2
17 9 13 0 9 9 2 7 15 13 13 3 15 13 13 3 3 2
12 3 15 13 2 16 13 15 3 9 13 13 2
9 9 13 9 2 16 13 9 13 2
8 3 11 9 13 13 13 9 2
10 16 11 13 15 2 15 13 16 9 2
8 13 15 13 7 16 3 3 2
6 6 3 2 0 9 2
4 9 13 9 2
3 13 13 2
11 3 15 13 9 9 0 2 0 7 0 2
3 0 9 2
10 15 13 0 13 2 16 13 13 9 2
2 9 1
2 11 9
5 3 13 13 9 2
6 15 13 13 13 9 2
8 9 13 3 13 11 9 9 2
6 9 13 9 7 13 2
8 13 13 3 13 0 13 0 2
12 13 15 15 0 9 9 9 2 15 13 3 2
8 11 7 11 13 13 9 9 2
7 3 0 9 13 13 9 2
2 13 9
3 13 3 2
8 9 13 12 12 3 0 9 2
12 3 13 9 2 9 2 9 7 9 10 9 2
14 3 9 9 13 3 0 2 16 9 13 13 3 13 2
18 9 13 9 2 13 13 3 9 7 13 0 9 2 15 15 3 13 2
6 11 13 9 9 1 2
12 11 11 13 9 2 15 13 9 0 9 11 2
12 11 13 9 2 15 9 13 9 0 9 9 2
6 13 3 13 15 13 2
13 0 9 13 13 2 3 16 9 13 13 1 11 2
9 3 13 11 9 13 9 11 9 2
11 9 13 13 3 9 3 10 10 3 9 2
18 0 9 0 9 13 9 2 7 3 9 7 9 9 0 13 13 0 2
6 9 11 7 11 9 1
6 15 13 13 0 9 13
18 13 2 16 9 9 7 12 9 13 3 2 7 9 13 9 3 12 2
13 13 3 3 2 16 11 13 13 0 13 0 11 2
5 3 15 13 13 2
9 15 13 3 9 15 7 15 13 2
6 13 15 13 9 0 2
4 15 13 13 13
2 9 9
2 0 0
2 13 3
17 13 9 3 2 16 13 9 13 9 7 9 7 3 15 0 9 2
5 3 13 0 9 2
3 15 13 2
7 0 9 13 3 13 3 2
2 9 1
3 10 0 9
7 13 0 2 16 13 10 9
7 9 13 12 3 3 0 2
5 9 13 0 9 2
5 9 1 15 13 2
15 3 0 16 10 9 13 2 15 13 13 9 10 9 1 2
9 11 13 9 9 1 9 0 9 2
5 13 13 13 9 3
8 3 15 13 7 3 15 13 2
14 3 9 13 9 1 9 2 15 9 1 13 9 9 2
16 11 2 15 0 9 9 13 9 13 2 13 3 3 3 9 2
9 13 15 13 9 2 11 13 3 2
7 13 15 9 2 13 13 2
7 3 13 10 0 3 3 2
6 13 9 7 9 3 2
6 9 1 13 13 9 2
12 3 10 9 9 13 11 13 13 9 0 9 2
3 13 13 9
9 9 13 0 9 11 13 0 9 2
18 15 13 13 10 9 2 15 9 13 2 13 15 13 9 15 15 13 2
8 11 11 13 3 3 3 13 2
15 10 9 11 13 13 11 7 13 9 9 9 0 9 9 2
3 13 9 3
7 12 9 13 3 9 13 2
5 13 15 15 9 2
11 11 13 3 16 11 13 7 13 9 3 2
21 3 9 13 9 7 11 13 7 13 16 13 13 0 13 7 13 7 13 3 3 2
18 9 9 2 16 13 9 2 16 9 13 2 16 9 13 3 3 9 2
12 3 15 13 2 3 15 3 13 13 9 9 2
6 9 13 0 3 9 2
4 13 9 9 2
16 6 15 3 13 15 13 3 7 0 9 3 3 12 3 12 2
23 7 16 12 9 13 3 3 13 9 2 10 10 7 15 15 9 2 3 15 13 10 9 2
11 3 15 13 0 9 9 2 15 13 3 2
11 9 13 10 9 2 7 9 13 13 9 2
28 16 15 13 16 13 3 16 9 1 3 7 15 3 6 13 15 13 3 16 15 3 8 15 13 15 7 13 15
7 11 13 13 9 10 9 2
8 9 16 13 15 13 13 3 2
4 15 13 13 0
2 15 13
7 0 9 13 3 10 9 2
10 9 9 11 13 13 9 3 3 3 2
10 11 3 13 2 16 13 13 9 3 2
4 0 9 11 11
13 3 10 9 13 13 10 10 9 3 0 9 9 2
8 13 13 9 9 2 15 13 2
10 3 11 13 11 9 12 0 9 7 2
2 0 9
10 9 13 13 3 16 0 9 1 13 13
5 9 13 9 1 2
7 6 3 2 13 9 3 2
11 3 3 15 13 13 2 15 3 13 13 2
4 15 13 9 1
12 9 11 7 9 11 13 13 3 11 10 9 2
24 3 13 9 3 13 3 2 13 13 11 3 2 9 13 0 11 11 2 16 15 13 13 9 2
16 9 7 9 13 13 2 13 11 9 9 2 0 9 11 11 9
10 0 13 12 12 7 0 9 12 9 2
11 9 9 12 11 3 13 11 9 0 12 2
14 0 7 9 9 13 10 9 3 9 13 7 9 9 2
11 9 13 3 0 2 13 3 0 13 0 2
9 15 13 0 9 3 16 13 9 2
3 12 9 0
3 9 13 13
9 13 13 13 9 9 2 3 9 2
4 15 13 9 2
21 9 13 13 9 9 2 7 9 9 15 13 13 3 2 16 13 15 13 3 13 2
2 9 9
3 13 9 2
5 0 9 13 9 2
3 10 0 9
10 11 13 13 15 9 2 9 7 9 2
10 11 9 13 12 13 9 13 9 9 2
5 9 13 9 1 2
8 10 3 9 13 13 9 9 2
8 9 9 13 13 13 13 0 2
7 10 0 13 16 13 9 2
15 3 16 13 3 13 2 13 13 3 0 9 13 3 3 2
9 3 13 0 9 9 13 13 3 9
28 9 13 9 13 9 9 7 13 15 13 2 3 8 7 9 9 13 9 10 9 2 15 13 13 3 10 9 2
2 8 13
8 13 3 16 13 13 9 9 2
10 9 11 9 9 12 9 9 11 9 1
2 9 13
9 13 9 13 3 10 0 9 9 2
11 9 13 13 9 2 16 9 13 3 13 2
4 13 9 13 2
3 15 13 2
19 11 13 3 3 3 0 9 2 16 3 11 0 9 9 13 0 10 9 2
14 3 15 13 2 16 9 13 3 2 11 13 0 9 2
5 13 3 3 9 2
8 9 13 0 7 0 16 9 2
11 3 13 0 13 9 15 16 13 15 3 2
11 11 13 9 13 8 7 9 0 0 9 2
14 13 9 3 13 7 13 15 13 2 16 15 13 9 2
11 13 13 11 13 2 0 9 1 13 9 2
20 3 0 11 13 13 13 9 13 15 3 9 11 7 11 9 0 9 0 1 2
12 15 15 3 0 13 2 13 9 3 0 9 2
14 9 1 10 9 13 13 13 11 2 15 13 9 9 2
14 3 13 13 3 2 16 9 7 9 9 13 3 9 2
6 13 13 15 13 15 2
11 13 2 3 9 13 9 2 3 9 13 2
5 3 3 13 9 2
21 7 3 3 2 3 13 10 0 9 6 3 13 10 9 7 10 9 13 10 9 2
4 13 3 3 2
2 3 13
6 15 13 13 10 0 2
2 3 2
8 15 13 2 16 15 13 9 2
21 9 13 13 0 9 9 9 7 9 0 9 13 9 13 9 2 15 13 13 9 2
9 9 9 13 3 0 2 11 11 2
15 10 9 9 9 13 3 13 2 7 0 9 15 13 13 2
12 15 13 13 9 2 16 9 13 3 0 9 2
9 15 13 13 9 15 1 13 9 2
16 13 13 15 2 9 7 9 2 15 13 9 9 9 2 16 2
4 11 7 11 13
7 13 10 9 13 0 9 2
7 13 15 2 16 13 9 2
20 9 13 13 2 16 13 10 9 13 9 13 9 2 16 9 13 0 15 13 2
16 16 9 13 9 2 13 13 13 15 2 16 13 10 9 13 2
7 9 13 3 9 7 9 2
11 13 9 9 2 7 3 13 13 3 9 2
3 2 9 2
5 0 9 3 3 13
16 9 13 15 2 16 9 11 1 13 9 2 0 7 0 2 9
9 3 3 15 13 3 0 9 13 2
24 11 13 11 11 2 11 9 2 13 3 3 2 7 13 16 2 0 13 13 15 3 3 2 2
8 9 12 13 0 9 11 9 2
9 7 15 13 3 13 15 12 9 2
2 15 1
7 11 13 7 13 9 9 2
8 12 9 13 9 0 9 11 2
2 0 0
10 9 9 13 3 13 0 9 0 9 2
7 9 13 2 16 13 9 2
4 9 13 15 2
14 15 2 15 13 2 13 13 3 9 2 9 7 11 2
27 12 0 9 13 13 15 16 2 16 16 11 0 0 8 0 0 0 9 13 13 10 3 16 15 13 10 9
10 0 9 11 9 13 9 9 9 9 2
4 15 16 13 15
7 0 9 9 13 16 13 2
4 9 13 9 2
8 12 13 11 11 11 9 12 2
5 9 13 9 1 2
7 0 9 13 9 11 9 2
13 13 13 9 10 9 2 16 15 15 13 13 9 2
6 10 9 13 13 15 2
28 10 9 3 16 15 13 9 3 2 7 10 9 7 15 3 2 15 13 2 9 1 0 2 15 13 0 9 2
3 15 13 13
22 16 15 13 1 15 8 2 15 15 13 9 3 2 3 15 13 16 15 13 12 15 13
12 7 3 16 13 2 10 9 13 0 9 9 2
4 15 13 9 1
10 9 13 0 9 0 9 7 0 0 2
10 9 13 13 2 7 13 2 16 13 2
7 9 13 13 13 3 9 2
12 9 11 2 9 2 13 3 16 12 10 9 2
10 13 9 2 15 13 0 13 7 13 2
7 9 15 13 9 3 9 2
14 3 11 13 10 9 2 16 9 13 0 9 9 13 2
4 13 13 9 2
5 15 13 15 1 2
11 11 11 7 11 9 13 3 10 9 1 2
6 9 13 0 9 9 2
6 3 9 13 13 9 2
5 9 13 0 9 2
22 11 0 9 7 10 9 13 3 10 9 16 11 9 7 9 7 3 13 12 9 1 2
8 13 9 13 1 9 13 3 2
6 9 13 10 0 9 2
9 9 13 11 1 3 12 9 9 2
8 13 11 15 15 13 13 15 2
4 0 9 7 9
2 13 3
17 7 16 13 15 3 10 9 13 9 3 3 15 13 13 0 9 2
6 0 9 13 9 9 2
4 10 9 3 9
10 13 15 7 9 7 15 13 3 3 2
14 15 2 15 13 0 9 13 9 2 15 13 0 13 2
8 13 16 9 13 0 9 13 2
5 11 13 12 9 2
11 11 13 11 9 13 11 2 9 9 2 2
4 3 12 9 11
9 0 9 9 13 11 9 11 11 2
8 11 13 3 3 0 13 9 2
5 15 13 13 11 2
14 3 9 11 7 9 11 13 9 0 9 0 9 9 2
10 0 9 13 3 9 9 10 9 9 2
26 11 2 13 16 9 13 13 2 13 13 9 2 3 3 16 13 2 13 3 2 2 3 15 9 13 2
10 13 10 15 16 13 13 13 0 9 2
5 3 13 7 13 3
6 11 13 0 9 9 2
6 3 13 15 13 9 2
8 0 9 13 3 10 9 13 2
18 13 3 12 7 12 9 9 7 9 16 13 13 13 13 9 9 13 2
15 9 7 9 9 13 9 1 7 9 9 3 13 0 9 2
8 15 13 9 2 7 13 9 2
12 3 13 0 13 9 9 16 13 15 3 9 2
48 12 9 9 3 11 13 13 3 2 7 15 13 11 13 3 3 3 15 13 3 9 2 3 13 3 13 2 10 9 13 13 15 3 3 2 16 16 2 15 13 3 0 9 7 9 13 13 3
7 3 11 9 9 13 9 2
9 9 13 2 7 3 3 0 13 2
10 15 13 3 12 10 0 9 1 9 2
14 0 13 3 3 0 7 13 3 0 11 7 11 9 2
5 15 13 9 13 9
16 9 13 16 16 9 3 13 2 3 15 13 9 7 13 9 2
8 3 2 13 3 0 3 13 2
10 12 9 13 9 2 16 9 13 9 2
8 15 13 15 0 2 10 0 2
4 9 13 9 2
6 9 9 13 3 13 2
7 15 13 0 13 13 9 2
3 13 15 2
13 13 13 9 10 9 2 16 15 15 13 13 9 2
4 13 9 15 2
15 11 13 10 1 9 9 2 16 13 15 3 0 13 13 2
3 3 9 1
17 13 13 9 13 9 3 13 2 16 3 13 13 9 2 13 2 2
13 11 13 9 12 13 3 15 2 3 9 13 9 2
16 9 1 13 9 13 3 0 9 2 15 13 9 3 12 9 2
5 9 13 12 9 2
15 15 13 9 9 2 15 13 13 15 3 13 2 0 13 2
10 15 13 16 10 9 13 15 7 15 15
3 9 13 0
5 11 13 9 9 2
11 13 9 9 13 13 3 12 9 9 9 2
2 9 13
10 11 0 9 13 0 2 9 7 0 2
12 15 1 15 13 9 2 16 9 13 9 9 2
4 9 13 9 9
11 15 2 15 13 13 13 15 3 2 13 2
6 10 9 15 3 13 2
12 11 13 3 12 11 9 2 15 12 13 0 2
10 6 13 10 9 2 3 15 13 9 2
3 0 9 2
6 9 1 9 13 0 2
5 9 13 9 9 2
10 15 13 13 9 2 16 15 13 9 2
9 15 13 16 15 13 3 0 9 2
4 15 13 13 2
3 10 9 2
8 9 15 15 13 2 9 13 2
7 9 9 13 11 9 1 2
6 3 9 9 13 13 2
12 15 1 9 13 13 9 9 9 7 9 9 2
12 13 2 16 11 9 13 9 11 1 13 9 2
6 9 13 13 1 9 2
11 9 13 9 13 9 2 9 13 3 9 2
3 9 13 9
13 15 13 13 13 9 2 7 11 13 15 10 9 2
5 0 9 10 9 13
9 13 15 13 16 13 13 9 9 2
5 15 13 9 15 2
2 13 3
7 0 9 13 13 3 13 2
5 9 13 3 9 2
4 3 13 13 2
11 9 15 13 13 2 7 9 13 13 13 2
14 9 11 13 13 3 0 9 2 15 13 3 0 9 2
10 13 10 9 15 13 16 2 6 2 2
2 13 13
10 13 13 9 9 9 12 2 12 9 1
13 9 13 3 9 9 7 13 13 2 9 7 9 2
6 9 13 0 0 9 2
2 10 3
10 9 13 9 3 3 16 0 9 13 2
19 11 9 9 9 13 3 2 13 9 2 9 1 9 9 13 3 12 9 2
6 9 9 13 13 9 2
8 9 13 0 9 16 10 9 2
11 0 13 9 9 3 13 9 13 0 9 2
9 7 15 13 9 3 13 2 15 2
10 9 13 9 13 2 9 13 3 3 2
6 15 13 3 9 1 3
4 15 13 13 2
5 9 13 13 11 2
5 15 15 13 13 2
3 0 9 9
2 9 13
6 15 13 3 12 1 2
8 3 13 13 0 9 13 9 2
19 16 13 0 9 11 13 0 2 0 13 9 2 15 13 2 2 3 2 2
6 9 13 0 16 15 2
2 10 9
18 7 3 15 3 13 1 9 9 9 7 9 13 2 9 13 16 9 2
5 15 13 13 11 2
2 10 9
9 9 13 3 11 11 9 0 9 9
6 11 9 13 12 9 2
6 11 13 9 3 0 2
2 9 9
7 11 13 0 0 16 9 2
13 11 11 13 2 16 13 0 9 13 3 3 0 2
6 12 3 12 13 12 2
11 13 15 2 16 3 15 13 3 10 9 2
16 11 13 9 0 9 2 3 9 13 7 11 9 13 9 9 2
18 9 13 2 11 13 9 9 2 13 7 13 11 1 9 1 2 12 2
13 11 9 13 12 1 1 13 8 2 8 7 9 2
11 15 13 13 3 11 2 15 0 9 13 2
4 13 13 9 2
7 15 15 3 13 3 13 2
3 3 13 9
9 3 13 3 3 2 7 3 0 2
3 3 13 3
3 11 9 11
24 3 15 13 3 10 9 9 11 11 12 9 13 0 8 11 8 8 7 3 13 9 9 11 2
4 13 9 0 2
19 15 13 15 9 11 0 9 2 15 13 13 9 15 1 16 11 9 9 2
4 9 13 9 2
8 9 13 13 13 3 12 9 2
11 11 13 11 9 7 13 9 9 13 9 2
11 11 9 13 13 12 9 9 0 9 1 2
2 13 9
10 9 13 13 3 3 0 16 9 13 2
8 2 7 9 2 2 11 13 2
6 3 9 9 13 9 2
2 0 9
3 9 13 9
12 9 13 9 9 15 2 16 15 13 13 11 2
23 13 16 13 2 16 0 9 7 9 13 13 13 15 16 15 13 13 0 3 0 2 7 2
11 9 13 0 9 3 0 9 13 13 3 2
4 15 13 0 2
7 11 13 3 2 13 2 2
8 0 13 13 13 13 0 9 2
12 11 1 13 9 13 3 3 7 13 13 9 2
5 0 9 3 13 13
4 9 1 9 2
3 0 3 13
7 9 13 3 9 9 9 2
3 13 13 13
8 11 13 13 0 9 9 9 2
5 9 13 12 12 2
5 13 13 10 9 2
2 0 9
11 15 13 13 3 3 13 3 9 13 13 2
12 3 9 13 3 0 2 16 15 13 13 9 2
9 10 15 13 3 9 1 3 9 2
2 0 9
10 9 1 9 13 13 9 9 7 9 2
5 11 13 3 9 11
7 11 13 3 12 9 9 2
4 9 13 9 2
15 9 0 7 0 9 13 3 2 7 3 3 2 9 9 2
8 3 13 3 3 0 13 15 2
9 9 9 1 9 13 15 0 9 2
5 15 13 13 9 2
13 9 13 0 7 0 0 2 16 13 15 0 9 2
4 8 7 0 9
6 9 11 9 13 12 2
8 9 13 13 0 9 1 9 2
8 13 2 16 13 13 9 0 2
5 11 13 0 9 2
8 3 11 11 13 13 2 16 2
4 15 13 0 2
12 9 2 15 6 2 16 15 13 13 1 9 2
7 11 13 15 12 9 0 2
6 15 13 13 0 9 2
5 15 13 13 11 2
9 10 9 9 13 3 15 11 1 2
9 15 1 9 13 11 9 0 9 2
8 13 15 9 7 13 15 9 2
17 3 12 9 9 12 13 9 13 9 9 13 3 10 9 9 9 2
12 13 13 13 0 9 2 16 9 13 10 9 2
7 9 13 3 0 0 9 2
5 13 13 13 3 2
4 11 13 9 2
10 9 13 9 13 13 9 9 9 1 2
7 15 13 11 2 12 11 1
4 3 0 9 2
10 9 13 3 0 7 3 3 13 9 1
15 3 9 13 13 9 13 9 9 7 9 2 13 9 9 2
6 9 9 13 13 9 2
6 13 9 3 9 9 2
13 9 0 7 0 2 0 7 0 1 13 13 13 2
6 13 13 13 9 9 2
2 0 11
5 11 13 3 3 2
6 15 13 13 13 9 2
4 9 13 9 3
4 9 13 13 9
17 9 13 15 2 16 9 13 3 0 9 2 16 15 13 15 0 2
10 11 9 13 12 9 13 3 9 1 2
13 9 13 13 9 7 9 7 9 7 0 0 9 2
23 9 9 13 0 2 15 13 12 9 7 0 2 3 13 9 2 7 15 13 3 0 9 2
15 9 1 3 13 0 9 13 9 2 0 13 9 1 13 2
15 0 9 9 13 13 15 2 16 15 3 13 13 9 9 2
2 13 3
17 9 0 9 13 2 16 13 13 2 7 9 13 0 13 13 3 2
11 13 3 7 3 2 3 15 13 3 13 2
7 9 13 13 13 9 9 2
12 13 13 10 13 16 13 9 7 9 9 13 2
10 3 9 13 15 1 3 3 9 3 2
4 11 15 13 2
10 3 0 13 13 13 9 3 13 9 2
6 15 13 10 0 9 2
6 15 13 9 3 0 2
4 15 13 9 2
8 15 13 13 11 9 12 1 2
4 9 13 9 2
4 3 13 3 2
6 9 15 13 11 9 2
10 11 9 13 0 2 3 12 12 9 2
5 13 7 13 13 2
14 16 13 13 3 2 3 11 9 13 3 13 0 9 2
10 10 9 13 0 2 16 13 3 15 2
7 3 13 9 13 12 9 2
4 13 0 9 2
24 3 3 13 10 9 3 3 3 16 13 0 9 3 15 13 13 8 7 3 9 1 10 9 2
5 10 9 13 13 2
6 9 13 13 13 9 2
14 7 10 10 9 3 13 13 3 3 13 7 13 15 2
14 9 13 9 9 9 3 13 9 9 9 13 9 1 2
7 0 9 9 13 3 0 2
12 9 13 9 3 13 3 13 9 13 9 3 2
23 15 3 13 11 13 10 9 2 16 12 9 13 13 0 9 9 2 15 13 13 15 0 2
4 13 13 0 2
8 9 13 3 13 2 11 13 2
5 10 9 13 13 2
7 15 13 11 3 16 11 2
7 11 9 13 3 3 3 2
8 9 11 0 9 7 9 13 9
17 15 13 11 7 13 9 2 16 9 13 2 13 11 13 15 3 2
2 0 9
14 9 13 3 3 2 16 15 1 13 13 13 3 9 2
4 15 13 3 2
4 0 13 13 13
5 13 15 3 9 2
13 3 0 13 9 13 13 9 13 0 9 0 9 2
9 11 13 9 13 16 9 13 9 2
25 11 13 9 2 15 13 15 0 9 2 7 3 3 0 15 13 2 16 3 9 9 13 10 9 2
5 15 13 9 9 2
19 13 9 9 3 7 3 13 9 2 16 3 3 9 13 13 2 13 11 2
4 9 13 0 2
4 9 13 13 2
2 9 9
29 11 9 9 2 9 7 9 9 9 2 13 9 0 1 0 0 9 2 15 3 13 13 13 9 9 7 9 2 2
17 15 15 13 2 16 9 13 3 0 13 13 3 0 2 0 9 2
6 13 13 15 3 2 2
9 9 13 13 2 16 15 3 13 2
17 13 13 13 2 16 10 15 13 13 11 9 9 11 9 3 3 2
8 10 9 13 3 10 12 9 2
9 9 13 11 3 3 3 9 13 2
3 13 9 2
15 9 13 13 9 7 13 0 8 2 8 2 8 7 9 2
5 6 13 13 0 2
3 13 9 2
4 13 9 9 2
3 13 13 13
10 15 13 0 9 2 15 13 3 13 2
8 9 3 12 3 9 13 9 2
7 0 9 11 13 13 13 2
18 8 11 13 9 2 15 13 12 9 1 0 9 2 12 9 1 11 2
8 13 9 10 3 16 9 15 2
9 11 15 13 11 9 9 1 9 2
16 16 3 13 2 3 13 13 3 0 7 0 0 16 9 1 2
4 6 3 0 2
4 9 9 13 9
5 15 13 9 3 2
12 10 9 9 7 3 9 13 9 1 0 9 2
9 11 7 11 13 13 10 9 9 2
6 7 15 13 0 13 2
2 0 9
4 15 13 9 2
11 2 9 13 3 13 3 2 16 3 13 2
8 9 9 13 13 13 9 11 2
6 13 13 10 9 3 2
6 15 13 9 9 1 2
10 9 9 13 15 2 3 15 13 13 2
4 15 13 13 3
6 9 13 11 0 9 2
10 13 13 10 9 2 16 15 13 13 2
2 13 13
5 9 13 3 9 2
2 0 9
3 0 15 1
16 11 11 2 15 9 12 15 3 3 13 11 9 13 9 9 2
8 7 15 13 9 9 9 13 2
9 11 7 11 11 13 11 3 3 2
10 15 13 0 9 7 15 13 0 0 2
6 9 13 13 3 3 13
4 9 13 13 9
4 11 2 9 9
2 9 13
10 0 9 9 13 2 16 15 13 9 2
2 9 11
10 3 11 9 13 3 0 7 3 0 2
3 13 9 2
3 13 15 15
6 3 15 15 15 13 2
3 9 11 9
5 13 11 10 9 2
15 3 3 9 9 13 3 0 9 16 15 2 15 11 13 3
2 13 13
3 15 13 9
7 13 9 1 13 10 9 2
12 0 9 13 15 2 16 13 13 9 3 3 2
3 10 9 2
4 9 13 3 12
9 13 15 15 13 2 3 3 3 13
6 15 13 13 9 13 2
12 9 7 9 0 9 1 13 3 13 9 9 2
7 13 9 3 13 9 11 2
2 13 13
2 3 3
4 9 13 15 2
8 9 9 13 0 3 12 9 2
7 2 13 15 13 0 9 2
4 15 15 13 2
22 3 9 1 15 2 16 11 13 13 3 11 11 9 2 13 9 9 0 0 9 9 2
9 11 9 13 13 3 3 9 1 2
6 9 13 13 3 3 2
12 11 13 9 3 13 2 15 11 10 9 13 2
4 9 13 3 9
4 15 13 3 0
5 13 3 9 1 2
16 11 13 9 0 9 16 0 9 13 13 11 2 11 7 11 2
7 9 15 13 2 15 13 2
6 15 13 3 1 9 2
7 13 15 13 3 15 1 2
11 10 15 13 2 0 9 0 9 3 13 2
2 0 9
2 0 9
9 13 9 9 13 13 9 9 9 2
10 3 13 13 9 9 9 9 0 9 2
6 9 13 3 3 9 2
7 10 9 13 9 1 0 2
5 11 13 9 13 2
3 10 9 15
8 15 13 13 15 9 10 9 2
5 11 13 9 1 2
10 13 13 3 13 2 15 9 3 13 2
5 9 13 11 11 9
7 11 13 9 3 13 9 2
5 15 13 13 3 3
8 12 15 13 2 9 2 11 2
3 9 13 0
15 9 13 12 9 3 9 7 15 1 0 9 11 9 11 2
4 13 9 13 3
3 13 3 13
7 11 11 13 9 0 9 2
8 15 1 15 13 9 13 0 2
7 11 13 13 0 9 9 2
4 15 13 9 2
3 12 9 13
10 13 0 2 16 11 13 15 13 11 2
15 3 12 9 9 13 13 3 9 16 0 9 12 0 9 2
4 11 9 11 9
4 13 11 7 13
2 13 13
6 16 15 13 3 3 2
7 10 0 9 13 13 9 9
7 10 0 9 13 3 0 2
11 3 13 9 2 9 9 2 7 9 1 2
14 0 9 9 13 9 2 7 13 15 9 9 13 9 2
7 0 9 13 9 9 9 2
10 15 13 9 10 3 16 13 13 15 2
13 9 13 13 9 0 9 7 3 15 13 3 9 2
9 0 2 0 9 13 9 16 9 2
4 15 13 11 9
8 15 13 13 13 15 11 15 2
12 13 15 13 16 13 9 2 11 13 13 3 2
12 9 13 9 9 9 7 3 13 15 0 9 2
6 15 13 13 13 15 2
11 15 15 13 11 2 3 16 13 13 15 2
15 3 13 9 3 13 9 2 15 11 9 3 13 9 12 2
4 15 13 9 2
11 11 3 3 13 16 13 13 9 0 9 2
11 9 9 9 9 12 9 13 3 3 0 2
3 3 9 2
10 15 13 13 9 2 16 9 13 3 2
26 15 13 15 0 2 7 15 13 10 10 9 7 15 13 3 13 15 3 7 13 16 13 0 15 13 2
6 3 0 9 13 13 2
7 15 13 0 12 9 11 2
9 9 13 3 16 13 13 9 0 2
9 7 15 13 13 2 16 13 15 2
5 15 13 0 0 2
10 11 9 13 13 3 2 15 15 13 2
11 16 13 3 9 12 2 9 13 3 0 2
4 15 13 12 12
5 9 13 9 9 2
13 10 9 13 9 13 13 9 9 9 9 2 9 2
3 13 9 15
9 16 15 13 13 2 13 15 3 2
3 13 15 2
4 3 13 13 2
15 15 13 2 13 9 9 2 13 3 9 2 15 9 13 2
11 13 15 13 10 9 13 9 3 12 9 2
10 13 15 9 2 16 9 13 13 3 2
13 15 3 2 0 9 2 13 11 16 11 9 13 2
2 3 3
8 10 9 13 13 3 0 9 2
7 9 13 13 3 0 9 2
13 0 13 0 9 3 3 3 15 13 13 2 9 2
6 3 9 13 0 9 2
3 13 9 12
9 15 13 15 13 3 13 15 13 2
2 13 11
8 9 9 11 13 13 3 13 2
12 9 13 0 13 0 9 11 7 9 0 9 2
6 15 13 13 10 0 2
12 9 9 13 0 9 2 9 9 13 10 9 2
4 9 13 3 3
2 9 1
5 11 9 11 9 1
3 9 13 2
6 9 13 9 7 9 9
8 7 10 9 15 13 3 9 2
5 9 13 3 1 2
5 3 11 13 3 2
3 9 3 9
3 13 3 2
9 13 10 9 13 0 7 0 3 2
8 3 9 13 13 11 3 13 2
3 3 13 13
10 16 9 13 9 2 13 9 0 13 2
9 3 3 13 3 0 9 10 9 2
7 15 13 13 9 9 1 2
3 13 15 3
9 15 9 3 13 3 3 0 9 2
6 11 13 13 9 9 2
36 7 3 11 7 11 7 11 7 9 9 11 11 7 10 9 13 15 9 16 13 13 9 9 7 9 8 13 9 15 13 13 9 1 13 3 2
5 11 7 11 13 2
3 13 15 2
11 10 9 15 13 0 9 9 9 1 11 2
8 9 13 3 3 7 0 0 2
7 10 15 0 9 13 13 2
11 3 9 9 13 13 13 3 3 16 9 2
2 13 3
3 10 9 2
4 3 13 9 2
6 9 13 10 9 9 2
14 9 9 13 11 2 9 11 7 9 9 11 7 11 2
10 15 13 2 16 13 2 16 13 9 2
2 3 13
7 2 6 13 13 15 13 2
7 11 13 3 0 9 9 2
13 10 9 13 3 3 0 9 2 16 13 3 15 2
9 13 3 2 9 3 13 11 1 2
9 3 15 13 12 9 1 12 9 2
4 15 13 9 9
5 13 13 12 3 2
11 11 9 13 9 13 3 0 9 9 9 2
5 15 13 3 13 0
13 0 9 1 13 3 0 9 2 9 13 3 0 2
6 15 13 3 3 3 16
13 6 16 15 3 13 3 16 15 13 3 3 6 2
6 10 10 9 9 13 2
13 13 13 3 13 0 9 15 2 13 11 13 9 2
5 9 13 12 12 9
5 15 13 13 9 9
6 3 15 13 16 9 2
9 0 9 10 9 9 13 3 9 2
12 10 10 9 9 13 3 13 1 9 0 9 2
10 3 13 13 15 13 9 13 13 9 2
6 15 13 13 13 9 2
12 13 3 13 2 3 15 13 13 10 10 9 2
7 10 9 13 15 9 9 2
8 16 13 13 2 13 9 9 2
5 9 13 0 9 2
14 0 9 13 13 3 3 2 13 9 3 13 7 13 2
5 13 3 9 9 2
12 0 9 13 15 2 13 15 13 7 3 15 13
2 3 13
3 9 13 2
4 11 13 11 2
10 13 10 9 13 9 13 10 9 9 2
9 13 15 13 16 15 2 3 12 2
2 13 15
18 9 9 13 13 3 3 9 9 2 7 15 13 3 3 8 7 9 2
7 12 9 9 13 9 1 2
9 9 9 13 13 13 12 9 1 2
8 9 9 13 12 9 9 1 2
9 7 3 10 12 9 13 13 9 2
6 3 13 13 0 9 2
5 11 13 9 0 2
16 11 13 9 13 3 3 13 2 16 13 15 13 13 0 9 2
21 16 15 13 13 13 3 9 2 13 13 9 9 1 2 15 3 13 13 13 15 2
4 9 13 3 2
5 13 15 0 0 2
8 0 0 9 9 9 13 13 2
9 9 13 0 2 7 13 3 15 2
10 9 9 2 9 9 7 13 16 13 2
10 13 16 13 3 13 13 7 13 15 2
11 15 13 13 3 0 16 9 2 3 9 2
14 15 13 13 9 7 15 13 3 0 9 9 10 9 2
4 15 13 9 2
10 15 9 13 2 13 1 10 0 9 2
6 9 13 11 13 9 2
4 11 3 3 2
7 3 13 9 7 13 3 2
6 0 9 13 0 11 2
24 9 13 13 13 12 9 0 9 9 2 7 10 9 16 13 13 9 7 9 2 9 13 13 2
11 3 11 13 3 9 12 7 12 12 9 2
3 13 13 13
5 15 13 15 0 9
10 15 13 13 0 2 0 3 9 13 2
14 9 13 9 13 15 1 2 16 0 9 13 3 13 2
7 9 2 9 13 0 9 2
15 11 11 9 13 9 11 2 10 15 13 10 0 0 11 2
13 13 13 10 9 2 16 13 13 13 9 1 15 2
2 9 9
8 3 3 13 15 12 9 0 9
9 13 0 7 13 2 10 9 13 2
4 9 13 15 2
10 15 13 13 0 9 3 9 11 9 2
12 13 9 9 13 9 3 2 16 15 13 13 2
5 9 13 9 1 2
8 15 15 13 3 13 0 9 2
3 12 9 13
5 13 15 3 9 2
7 13 15 3 13 3 13 2
6 13 3 10 0 9 2
9 9 11 13 11 9 13 12 9 2
13 9 9 13 3 0 2 16 15 13 13 9 3 2
14 9 9 13 9 11 11 13 3 13 9 13 9 9 2
6 11 13 9 7 13 9
7 9 9 1 9 13 0 2
17 11 1 3 13 0 9 13 9 9 9 3 2 16 9 13 9 2
2 9 9
15 11 13 9 9 9 13 9 1 13 12 9 9 9 9 2
3 9 9 9
8 13 13 0 2 16 13 13 2
16 16 15 13 2 13 13 9 2 7 10 9 15 13 13 13 2
4 9 15 13 2
11 0 9 9 13 13 2 13 9 9 9 2
16 15 13 3 13 10 0 9 9 2 3 16 0 3 15 13 2
15 11 15 13 13 0 2 16 13 3 9 9 7 9 13 2
4 15 13 3 2
9 9 13 13 3 10 9 13 9 2
20 3 15 15 13 2 16 15 13 3 0 10 9 2 16 13 13 13 3 9 2
9 0 9 1 9 13 3 12 9 2
9 11 3 0 9 13 15 2 16 2
2 9 13
16 9 13 13 3 9 3 0 9 2 3 16 13 0 9 1 2
2 9 9
10 13 13 13 2 3 0 9 15 13 2
14 10 9 13 9 2 7 9 13 13 3 12 9 1 2
13 9 7 13 3 13 7 13 3 13 9 1 9 2
11 16 13 9 9 3 3 16 13 3 13 2
12 9 13 3 13 2 0 9 13 13 0 9 2
11 7 9 3 13 2 16 3 10 9 13 2
6 11 13 15 9 9 2
11 15 13 9 13 2 16 13 10 9 3 2
7 9 13 9 3 13 9 2
9 15 13 9 2 15 3 13 12 2
15 0 13 13 11 2 16 15 13 10 7 15 9 2 7 2
17 3 0 9 2 3 3 9 9 13 10 10 9 16 0 7 9 2
4 9 13 9 2
8 15 13 9 13 0 9 9 2
6 15 13 13 1 9 2
11 9 13 13 15 15 7 3 15 13 13 2
5 12 9 1 12 9
5 0 9 9 9 1
2 10 9
4 3 13 13 2
5 15 13 9 1 2
12 13 13 2 13 3 7 16 3 3 9 13 2
12 13 10 9 2 15 9 13 13 13 9 9 2
6 15 13 3 11 11 9
4 10 9 13 13
18 13 13 3 13 2 3 13 3 1 9 9 2 15 13 13 9 9 2
2 13 13
9 9 13 9 13 3 9 13 9 2
23 11 11 15 9 3 13 13 3 3 3 13 3 13 7 10 9 15 13 15 13 3 0 0
12 6 16 13 15 13 3 13 3 13 10 10 9
8 0 9 3 13 7 13 15 2
2 13 13
2 13 9
11 15 13 13 15 10 9 2 16 13 9 2
9 10 0 9 13 13 13 9 3 2
23 15 13 13 9 9 13 9 1 7 13 0 9 2 7 13 3 9 13 9 7 13 9 2
2 0 9
4 11 12 0 9
4 13 9 9 2
6 15 15 13 7 13 2
3 13 16 13
3 0 0 9
4 13 15 13 2
3 0 13 2
7 9 13 13 3 12 9 2
8 7 3 3 2 15 13 9 2
7 13 2 16 15 13 9 2
7 15 10 9 13 3 13 2
14 0 9 13 13 12 9 9 2 0 9 9 13 9 2
20 7 16 11 13 9 2 15 13 13 12 2 7 12 9 7 15 13 11 1 2
9 15 13 9 11 13 8 11 9 2
6 9 13 13 9 3 9
7 7 3 3 13 12 9 2
9 9 13 3 0 9 10 9 9 2
12 13 9 3 3 2 3 9 9 13 13 9 2
5 9 13 3 0 2
4 13 9 13 9
10 3 10 9 13 10 9 3 9 1 2
7 9 13 3 3 9 1 2
11 11 11 13 12 9 7 13 9 3 9 2
5 13 16 13 13 9
7 0 9 2 9 9 11 11
4 7 9 3 13
6 9 13 13 13 13 2
14 15 13 13 9 7 12 2 7 15 13 13 9 9 2
3 13 15 3
5 9 9 3 9 9
7 3 3 13 3 0 9 2
14 15 13 2 16 9 13 13 0 9 7 15 13 13 2
13 11 9 7 11 13 0 9 1 13 9 9 13 2
7 11 9 13 3 13 3 2
5 9 13 3 9 2
4 9 13 13 2
3 15 13 3
10 3 0 13 13 9 13 9 0 1 2
7 9 9 13 3 9 0 2
8 9 13 0 9 2 13 13 2
4 15 13 3 2
5 15 13 9 9 2
6 9 13 13 3 9 2
9 11 9 13 0 9 13 9 13 2
5 12 9 9 13 2
7 9 13 9 13 15 15 2
5 11 7 11 13 2
9 15 13 9 2 3 11 13 9 2
6 12 9 13 10 9 2
10 9 13 13 15 16 13 15 13 15 2
11 3 13 3 12 9 13 16 16 13 3 2
2 13 13
10 3 13 13 3 0 9 16 16 16 2
8 9 13 9 2 9 7 9 2
3 13 13 2
2 13 0
22 15 13 3 13 13 15 13 9 0 9 2 13 3 13 3 3 13 9 9 11 13 2
11 12 9 13 9 9 13 9 11 9 9 2
9 9 9 13 3 0 9 2 9 2
15 9 9 13 11 9 2 0 2 0 2 0 2 0 9 2
2 8 2
9 9 9 13 13 9 7 13 9 2
6 11 11 11 13 9 2
5 9 13 9 9 2
7 9 13 9 13 9 12 2
12 15 13 7 13 9 11 0 9 11 11 13 2
8 0 9 1 13 13 10 9 2
12 15 13 13 13 2 0 13 12 9 3 9 2
5 10 9 13 0 2
8 9 9 0 9 13 10 9 2
7 9 13 10 9 13 13 2
4 10 9 0 9
3 13 9 2
7 2 15 15 13 3 3 2
9 13 9 2 16 9 9 13 9 2
16 13 11 7 9 11 7 3 13 3 0 2 16 3 13 13 2
8 13 16 15 13 12 13 12 2
5 9 13 13 9 2
7 15 15 3 13 13 9 2
6 2 9 13 13 13 2
7 10 9 7 9 15 13 2
10 9 9 13 3 3 0 0 16 0 2
7 2 3 3 9 13 9 2
9 15 13 13 9 11 9 7 9 2
17 0 13 2 16 13 11 9 13 3 0 9 16 11 2 13 11 2
7 13 3 7 13 9 9 2
11 9 0 9 13 3 0 7 13 7 13 2
16 9 13 13 15 2 15 11 13 2 15 13 2 15 7 3 2
11 13 3 0 2 16 13 13 3 13 15 2
8 13 15 13 2 15 15 13 2
14 11 9 13 9 3 13 9 1 12 9 1 13 11 2
13 13 3 0 3 2 16 9 1 13 3 3 9 2
9 15 13 9 9 15 9 13 9 2
10 0 11 11 9 0 9 13 10 9 2
8 15 13 9 13 13 3 9 2
7 15 1 13 12 0 9 2
2 9 9
13 9 11 11 2 3 10 9 13 3 13 0 9 2
5 15 13 9 9 2
13 11 0 9 13 13 3 9 2 16 13 3 9 2
17 3 13 9 11 2 3 9 13 13 0 11 0 9 13 0 9 2
19 11 11 13 7 13 9 9 11 2 15 13 9 9 11 2 7 13 3 2
4 9 13 9 2
15 0 9 13 13 9 2 7 3 0 9 13 9 3 13 2
13 16 15 3 13 10 9 9 2 3 13 15 15 3
13 3 3 15 15 13 2 16 10 9 13 3 13 2
4 9 13 3 2
2 9 12
5 11 13 1 9 2
8 9 13 2 16 13 13 9 2
4 6 13 13 3
5 13 15 3 15 2
4 9 3 0 2
21 15 13 3 9 13 13 3 0 9 2 7 3 0 15 13 0 7 15 13 9 2
10 13 3 3 9 3 2 13 0 9 2
12 10 9 13 13 15 13 7 9 3 7 9 2
21 9 13 13 9 3 0 9 2 3 9 13 0 2 2 9 2 7 9 9 13 2
5 9 13 13 0 2
6 10 9 13 3 3 2
27 15 13 9 13 9 1 0 9 3 2 16 3 13 13 9 9 13 9 11 2 15 9 13 15 3 11 2
2 13 9
8 9 1 3 9 13 9 9 2
7 15 15 13 16 9 13 2
20 10 9 13 13 12 9 7 3 13 9 7 13 3 9 2 3 13 13 0 2
10 16 9 13 0 9 2 9 13 13 2
2 3 2
2 10 9
15 3 13 15 16 10 15 9 13 13 10 0 16 0 9 2
5 15 13 15 0 2
5 3 15 13 13 2
6 15 13 3 13 11 2
3 13 15 3
9 9 3 13 11 7 11 9 3 2
5 15 13 3 13 2
10 16 13 3 0 2 13 13 3 13 2
9 15 13 9 2 3 13 13 13 2
17 9 13 13 2 16 9 13 9 1 3 9 0 2 12 9 1 2
12 15 13 9 7 3 3 9 3 13 13 9 2
18 3 3 12 9 13 9 7 9 15 0 9 13 13 3 9 0 9 2
12 11 9 13 0 3 0 9 13 9 0 9 2
6 13 15 13 16 13 2
15 3 0 9 13 3 2 0 9 9 13 3 13 13 0 2
11 9 13 13 11 8 7 11 9 9 12 2
10 15 13 10 9 3 16 10 9 13 2
4 9 13 0 2
6 13 13 10 0 9 2
7 9 13 13 3 11 9 2
4 2 15 3 2
8 13 15 13 0 16 15 13 2
9 9 13 13 16 13 15 13 9 2
8 9 13 9 1 7 13 9 2
13 13 15 13 13 13 9 9 3 7 13 15 9 2
2 0 9
2 13 9
6 13 13 13 13 15 2
8 13 15 13 3 2 15 13 2
6 9 13 13 11 11 2
5 13 3 13 3 2
2 10 9
6 9 13 9 9 12 2
5 15 13 0 9 2
9 0 9 1 3 13 3 0 9 2
21 15 13 13 3 9 3 12 9 9 0 9 2 15 13 13 13 9 1 3 13 2
6 9 2 13 11 11 9
9 10 11 13 0 9 3 0 9 2
3 9 13 13
10 10 9 13 2 0 2 0 2 0 2
10 9 1 11 13 13 13 3 3 9 2
3 13 9 3
4 15 15 13 2
17 3 0 9 13 13 9 0 7 9 0 16 11 9 9 0 9 2
6 9 13 9 9 13 2
13 3 15 13 13 9 2 3 0 9 2 10 9 2
9 11 13 13 10 9 9 16 11 2
4 9 0 9 9
16 3 13 3 0 9 2 16 15 13 13 2 13 0 9 9 2
3 13 13 9
3 10 9 9
6 11 15 3 9 13 2
10 3 15 13 3 16 16 13 9 3 2
3 15 13 9
11 11 0 9 11 11 13 0 9 2 16 2
19 11 1 0 13 9 15 2 16 9 13 13 0 2 16 3 0 13 0 2
12 15 1 16 13 3 0 2 13 13 3 13 2
12 11 3 13 0 9 2 15 13 10 9 1 2
14 9 11 13 3 0 9 13 2 16 15 13 10 9 2
15 6 2 6 2 13 3 2 11 13 7 13 9 12 9 2
11 15 13 9 0 9 3 16 9 13 3 2
28 15 13 3 13 11 2 16 11 13 3 9 2 11 10 9 13 13 13 11 2 15 13 13 13 0 9 9 2
9 0 9 0 9 13 3 9 13 2
19 15 13 9 7 9 13 2 7 16 13 9 13 13 2 3 13 9 3 2
6 11 13 3 13 9 2
14 3 0 9 9 13 13 3 7 13 2 9 7 9 2
5 9 13 15 9 2
17 13 13 3 15 2 16 13 13 3 10 9 15 10 9 13 9 2
8 0 9 13 11 10 9 10 9
5 7 9 15 13 2
3 9 13 2
2 0 9
8 11 11 13 13 0 9 9 2
6 9 13 3 9 1 9
16 13 3 13 2 3 13 9 13 2 3 3 13 13 13 9 2
7 15 13 9 9 13 11 2
7 15 13 3 12 9 13 2
9 9 13 0 13 2 16 15 13 2
3 3 3 2
13 15 13 3 0 2 15 13 3 13 3 9 9 2
15 15 13 9 2 13 9 3 0 3 7 13 9 7 13 2
7 10 9 13 12 0 9 2
4 15 13 9 2
3 9 0 9
15 15 13 3 11 2 16 15 2 3 3 2 13 9 9 2
7 13 13 15 13 9 2 2
8 12 9 11 0 13 3 9 2
4 13 9 9 2
6 0 9 9 13 9 9
18 11 9 13 0 9 9 13 3 3 0 9 9 9 8 8 8 8 2
2 3 13
8 13 3 0 9 7 0 9 2
15 9 9 13 0 9 13 9 9 7 13 9 2 11 13 2
6 9 13 3 13 3 2
3 15 13 9
9 13 13 0 2 16 9 13 9 2
5 13 13 15 15 2
4 9 13 13 13
4 3 13 13 2
4 0 9 7 0
9 11 9 13 9 16 15 13 3 2
17 15 13 13 9 2 15 13 11 9 9 2 7 13 9 15 1 2
15 15 13 13 0 3 2 13 10 9 13 9 1 9 1 2
2 13 3
4 9 13 0 2
9 10 9 13 2 15 13 0 9 2
17 9 13 11 10 9 1 3 13 9 9 13 11 7 11 0 9 2
7 3 0 9 9 13 13 2
2 10 9
3 15 9 2
12 13 9 2 16 13 10 3 3 3 11 9 2
11 13 3 13 13 11 11 9 9 0 9 2
15 7 15 13 7 13 9 7 13 3 3 3 16 15 13 2
12 13 9 3 9 7 15 1 2 13 13 13 2
3 15 13 9
17 11 0 9 13 3 9 2 15 15 13 9 9 9 13 11 11 2
6 15 13 13 15 15 2
12 13 15 3 2 7 15 13 16 10 9 13 2
26 15 13 3 2 16 0 9 2 9 7 9 13 13 3 7 13 2 15 9 1 2 2 0 9 13 2
7 9 9 13 9 9 1 2
16 13 0 9 2 3 9 9 9 13 13 2 8 8 3 11 2
9 9 13 13 0 9 13 9 1 2
4 9 9 13 9
5 15 10 9 13 2
19 0 9 3 2 10 9 3 9 13 15 2 15 13 16 3 13 0 9 2
6 11 13 12 0 9 2
23 0 9 13 13 15 13 9 2 15 13 15 0 7 13 10 9 2 15 15 13 0 9 2
6 7 13 3 3 9 2
3 13 9 9
7 9 13 13 9 0 9 2
5 9 13 3 9 2
11 13 0 2 16 13 7 16 13 3 9 2
6 13 15 3 7 3 2
8 15 13 13 3 3 9 9 2
12 11 13 11 9 3 3 16 15 15 3 13 2
10 9 13 15 3 13 9 7 11 9 2
4 13 3 3 2
5 9 13 3 3 2
7 3 13 9 13 9 9 2
7 13 10 0 9 7 9 2
11 9 13 0 3 13 7 13 10 3 15 2
4 13 9 0 2
14 6 2 9 13 3 0 7 13 3 3 0 9 1 2
9 0 9 13 3 13 3 9 9 2
5 9 1 13 11 9
4 13 13 15 9
7 9 13 13 3 15 9 2
6 13 9 3 9 13 2
10 15 13 13 9 2 0 9 7 9 2
8 13 11 2 15 13 3 0 2
18 15 13 3 3 13 0 2 16 9 13 9 2 9 2 9 7 0 2
3 9 13 9
7 9 9 13 15 13 13 2
7 15 13 13 0 13 9 2
7 0 9 13 0 16 0 2
14 15 13 13 3 9 12 2 13 15 3 13 10 9 2
2 13 9
24 16 9 13 12 9 2 15 3 12 10 9 9 2 3 13 3 0 9 15 2 3 9 13 2
11 13 9 13 9 2 7 13 15 9 9 2
4 16 13 10 9
2 0 9
9 9 13 0 13 3 9 13 0 2
8 9 15 13 12 9 2 3 2
4 9 3 9 13
3 15 13 9
10 10 9 13 13 12 9 0 9 9 2
12 13 10 9 3 13 16 9 13 0 9 3 2
12 3 13 9 13 3 9 7 9 0 9 1 2
8 9 13 2 16 13 1 9 2
4 13 9 11 2
14 9 13 3 12 9 2 7 13 9 7 3 13 13 2
12 9 13 9 13 3 2 3 15 13 13 9 2
6 15 13 2 7 11 13
6 10 9 13 13 0 2
11 15 13 9 1 0 9 2 3 15 1 2
15 13 13 16 9 13 13 9 2 16 3 13 12 0 9 2
6 13 13 16 9 13 15
3 15 13 13
7 9 13 8 7 9 9 2
13 9 9 13 9 13 3 9 2 9 9 7 9 2
8 13 13 3 2 13 13 9 13
8 9 11 13 11 9 9 13 2
7 0 13 9 7 9 1 2
21 13 9 13 2 16 15 13 9 9 2 7 13 13 13 2 16 15 13 9 9 2
6 13 3 9 11 13 2
6 9 13 9 0 9 2
14 16 13 13 2 16 10 9 13 9 2 13 3 3 2
8 2 13 15 13 13 3 9 2
2 9 9
2 0 11
7 13 13 13 15 2 11 2
9 15 13 9 1 2 13 7 13 2
18 15 13 11 7 13 9 2 16 9 13 2 13 15 3 13 15 3 2
4 9 13 9 13
9 13 9 7 13 3 7 13 15 2
3 9 13 13
2 0 9
7 11 9 13 9 9 9 2
4 9 13 3 0
7 9 13 13 13 10 9 2
7 9 2 15 13 3 11 11
9 13 3 3 0 9 13 16 15 2
14 3 13 13 0 9 7 9 13 13 7 13 9 9 2
20 11 0 9 11 7 11 11 13 11 11 9 2 3 15 13 3 13 9 9 2
11 3 13 9 2 7 15 0 13 0 9 2
8 8 7 9 11 13 0 9 2
2 10 9
13 11 13 15 9 11 11 7 11 9 13 9 11 2
11 15 3 13 13 15 2 13 9 7 13 2
6 3 13 3 3 9 2
20 0 9 13 9 9 2 13 13 2 13 9 2 13 2 7 13 16 13 9 2
15 9 13 3 0 7 0 9 9 2 15 13 13 9 9 2
3 9 13 2
9 9 13 13 9 9 3 13 9 2
9 9 13 9 13 0 9 9 9 2
10 9 13 9 0 0 9 7 0 9 2
7 15 13 3 3 10 9 2
9 13 11 11 3 16 13 11 11 2
7 13 13 0 16 15 13 2
8 9 9 9 13 15 13 9 2
6 11 13 11 0 9 2
13 13 0 9 13 3 9 7 9 2 15 13 13 2
13 15 13 3 9 13 15 13 15 16 15 13 13 3
8 3 0 9 15 13 10 9 2
12 9 13 3 0 9 2 7 3 13 0 3 2
5 13 9 13 9 2
8 1 9 11 13 13 0 9 2
6 13 15 13 3 3 3
8 11 13 11 9 11 11 13 2
6 9 13 11 3 0 2
8 9 12 9 13 9 12 9 2
13 0 9 13 13 9 9 2 9 2 9 7 9 2
4 9 1 13 2
9 15 13 13 9 9 15 3 16 9
7 11 9 9 9 2 9 11
6 9 13 13 10 0 2
2 9 9
8 9 13 3 13 1 11 9 2
7 15 13 15 13 9 9 9
19 11 13 0 2 13 9 9 7 13 9 0 16 13 3 2 11 9 13 2
6 16 13 15 13 15 2
4 13 9 1 9
6 9 13 9 12 9 2
8 9 9 13 3 0 16 9 2
5 13 3 3 13 2
4 3 9 13 2
10 13 9 13 9 16 9 13 13 3 2
14 3 13 16 9 13 0 0 2 13 15 3 3 3 2
2 3 16
10 9 13 13 2 7 15 13 13 0 2
15 15 13 3 13 2 16 13 10 9 1 13 9 0 9 2
13 9 13 3 0 2 16 13 8 9 13 15 3 2
12 0 9 13 9 9 13 0 9 2 11 9 2
16 9 9 13 9 13 2 9 13 0 9 2 9 15 3 13 2
22 3 12 9 9 9 2 15 13 9 9 2 15 13 0 9 9 9 16 11 11 3 2
17 11 13 0 9 2 15 13 3 13 9 2 7 10 9 1 3 2
8 9 9 13 9 13 13 13 2
4 3 0 0 9
12 2 11 9 2 7 0 9 9 0 9 13 2
4 3 16 13 2
18 11 13 2 16 9 13 13 9 9 2 15 13 13 13 9 15 1 2
14 9 9 9 9 1 13 13 10 9 13 3 0 9 2
6 13 0 7 0 9 2
4 15 13 15 2
18 13 3 0 9 10 9 9 7 9 7 13 10 0 9 0 9 13 2
7 3 15 13 15 3 11 2
2 13 9
15 3 16 15 13 13 13 13 10 0 2 16 15 3 13 2
10 9 11 11 13 3 13 3 0 9 2
5 11 13 9 0 9
14 15 13 9 7 9 2 3 3 2 9 7 9 9 2
8 12 9 13 12 9 9 3 2
18 9 13 13 3 0 9 13 9 2 7 9 9 13 0 9 10 11 2
5 9 13 0 9 2
13 0 9 13 9 9 13 3 3 13 9 13 9 2
7 13 15 3 10 9 3 2
6 3 13 10 1 9 2
5 0 13 0 9 2
6 0 9 10 10 9 2
7 6 16 15 3 13 10 11
13 11 9 13 13 9 2 16 9 9 13 15 3 2
9 13 15 15 2 16 13 9 9 0
3 15 13 9
7 9 2 12 2 13 9 2
12 15 13 16 15 13 10 9 3 3 3 10 15
4 9 9 13 9
4 16 3 13 3
9 0 9 13 0 9 13 0 9 2
9 16 13 3 9 2 13 3 9 2
4 13 9 9 2
13 16 9 13 0 9 3 13 2 13 16 9 13 2
13 7 11 13 3 10 9 13 3 12 12 12 9 2
16 13 13 15 2 16 13 3 9 7 9 9 9 13 10 9 2
2 9 11
18 3 0 9 3 13 0 2 16 15 13 9 9 7 13 3 13 9 2
5 13 13 13 9 2
7 13 13 9 2 13 0 2
6 13 13 3 13 11 2
5 15 13 0 3 2
3 0 0 9
8 3 15 13 15 3 16 13 2
5 11 13 13 9 2
5 9 13 12 9 2
3 3 13 9
4 9 13 11 1
3 9 13 13
6 13 16 13 15 9 2
12 9 13 9 3 2 3 9 13 8 7 9 2
6 11 13 12 0 9 2
11 7 10 9 13 9 10 12 9 3 9 2
25 16 15 13 13 0 11 11 15 13 13 3 15 3 2 0 9 13 15 13 13 13 15 0 9 2
15 10 9 13 9 2 7 15 13 0 9 0 9 13 15 2
4 13 15 13 2
12 15 1 13 9 13 15 16 3 15 15 13 2
6 9 9 9 13 9 2
2 9 1
12 9 7 9 13 0 0 9 0 9 9 9 2
15 9 13 0 9 2 9 0 9 7 13 15 12 9 3 2
2 9 13
9 3 0 9 13 10 9 16 0 2
3 15 13 13
7 6 13 15 13 0 3 2
4 15 13 13 9
20 11 13 9 11 2 3 13 3 0 7 0 16 10 11 7 11 2 7 3 2
5 9 13 9 3 2
12 15 13 9 2 9 2 9 9 7 9 9 2
8 9 13 13 9 13 9 11 2
4 15 13 3 13
8 0 9 11 13 3 3 0 2
6 9 13 9 13 9 2
6 3 3 11 13 3 2
10 9 13 9 2 15 13 9 0 9 2
3 3 13 9
3 10 9 9
6 7 0 9 3 9 2
5 15 13 0 9 11
5 3 9 9 13 2
7 11 13 0 7 11 0 2
6 3 13 9 12 9 2
9 11 11 13 9 3 3 12 9 2
6 13 3 9 0 9 2
10 13 13 3 15 16 13 15 9 9 1
15 15 13 13 15 2 15 15 13 3 3 13 6 0 9 2
3 13 9 2
4 13 13 0 2
17 16 9 13 13 9 2 3 0 15 3 13 2 16 13 9 3 2
8 15 3 13 3 15 2 16 2
5 9 15 15 13 2
14 9 13 3 9 9 7 13 9 3 7 10 9 3 2
6 3 15 13 3 3 2
10 3 11 9 2 0 9 9 13 9 2
5 12 9 13 9 2
19 0 9 9 13 10 9 3 12 9 9 2 7 10 9 13 3 3 9 2
13 9 13 3 3 15 2 7 13 15 13 3 13 2
19 16 15 3 13 13 3 9 7 13 3 3 2 15 13 9 9 13 15 2
7 3 13 0 9 16 13 2
10 15 13 10 9 7 15 13 10 9 2
13 9 13 13 3 9 1 2 7 15 13 0 9 2
14 16 9 13 9 2 3 11 11 9 13 3 15 13 2
4 15 13 9 2
4 11 13 9 2
10 13 3 13 2 11 13 2 13 9 2
4 13 9 9 2
11 13 9 13 9 13 9 3 13 9 9 2
6 15 13 0 1 15 2
5 13 11 11 10 9
16 9 13 7 9 7 9 0 9 7 3 15 13 13 0 9 2
2 0 9
12 9 9 13 13 10 9 7 3 13 12 9 2
6 16 9 13 3 13 2
3 12 0 9
3 13 13 13
11 9 13 13 13 9 2 13 9 7 9 2
14 0 9 7 15 1 13 9 9 13 9 9 9 12 2
3 3 1 9
2 13 12
11 9 3 13 9 13 3 13 3 0 9 2
7 13 3 3 16 15 13 2
6 13 13 13 13 9 2
4 9 13 3 2
19 15 13 9 9 3 9 9 7 9 2 9 7 9 2 9 7 0 9 2
10 15 13 13 10 9 2 13 0 3 2
19 9 13 3 13 9 0 9 7 9 13 13 0 9 1 2 16 13 9 2
9 9 1 13 13 10 9 9 13 2
14 3 13 3 13 10 9 2 16 9 13 13 0 3 2
10 0 11 10 0 9 13 10 9 9 2
7 15 13 13 11 10 9 2
5 15 13 9 13 3
5 15 13 3 3 2
5 0 9 15 13 2
4 13 13 10 9
3 9 13 9
2 0 11
16 8 2 8 2 8 2 8 7 0 9 13 0 1 3 0 2
9 9 13 13 3 9 7 3 9 2
4 13 9 13 2
9 3 15 13 10 9 13 15 13 2
6 9 13 13 12 9 2
3 13 13 13
2 9 9
16 15 13 3 10 0 9 15 13 3 3 7 3 15 13 15 2
8 11 13 3 3 16 9 11 2
3 13 13 9
7 15 13 3 3 3 3 2
10 11 9 9 13 9 7 9 13 9 2
4 15 13 11 2
2 9 3
8 15 2 13 2 13 0 9 2
10 6 15 13 13 15 3 13 0 9 2
5 9 13 9 3 12
5 15 15 3 3 13
17 9 13 13 2 7 9 13 3 3 2 16 9 13 0 7 9 2
3 9 13 13
5 3 15 13 13 2
2 13 9
11 15 1 0 9 9 9 9 0 13 9 2
5 13 13 9 0 2
7 11 13 9 1 13 9 2
8 11 13 10 9 10 11 9 2
5 15 13 15 3 2
17 0 9 13 15 2 13 9 13 3 9 3 12 9 9 1 9 2
6 9 13 9 13 9 2
3 10 12 9
5 3 13 15 9 2
5 13 13 11 9 2
13 10 15 10 9 9 3 13 2 13 10 0 9 2
12 13 3 9 13 9 15 13 7 15 13 9 2
15 12 9 13 9 7 9 2 7 15 13 3 13 3 15 2
9 9 9 13 3 3 3 16 9 2
3 13 13 2
9 10 9 13 3 0 9 10 0 9
9 0 9 13 3 9 7 3 9 2
14 16 9 13 2 3 13 3 13 15 9 3 13 9 2
11 9 13 13 0 2 16 13 13 3 9 2
4 10 9 11 2
6 15 13 3 0 10 9
5 0 0 13 13 2
8 2 10 9 13 13 9 9 2
9 2 7 9 13 2 2 15 13 2
13 9 7 9 11 13 9 13 2 7 13 1 9 2
2 13 9
14 11 13 3 13 0 2 16 9 13 11 9 13 9 2
8 9 0 9 11 13 0 3 2
8 9 13 9 13 13 0 9 2
9 11 13 9 1 13 13 13 9 2
6 11 9 13 3 0 2
5 10 9 13 3 2
18 9 11 11 13 3 1 9 9 2 16 13 9 9 3 13 13 3 2
4 15 15 13 2
9 11 1 0 9 13 3 0 9 2
13 0 9 13 13 2 15 9 13 12 9 9 1 2
11 13 9 0 0 9 2 15 13 9 9 2
5 2 13 13 3 2
7 13 13 3 9 7 9 2
6 15 13 0 9 13 15
15 9 13 10 9 3 2 16 13 9 3 13 10 0 9 2
7 9 9 13 13 0 9 2
5 15 13 9 3 9
6 9 13 12 12 9 2
7 3 13 7 13 9 9 2
4 15 13 9 2
8 9 13 13 0 9 9 9 2
12 15 13 3 13 9 2 15 13 13 9 9 2
3 15 13 15
3 13 9 1
17 15 13 11 0 9 2 11 11 11 9 2 16 9 13 9 12 2
7 13 3 2 16 13 9 2
18 11 11 13 13 2 16 13 0 13 9 2 7 3 0 13 13 0 2
6 13 13 0 2 16 13
7 15 13 3 16 3 3 2
5 9 13 3 0 2
6 9 13 2 16 15 13
2 0 9
12 9 9 13 3 2 1 9 2 9 7 9 2
4 15 15 13 2
9 0 9 9 13 13 3 16 3 2
9 16 13 0 13 2 15 13 13 2
23 13 13 3 9 12 2 15 13 3 0 2 9 12 13 15 3 13 2 15 10 9 13 2
31 15 13 9 2 16 9 9 9 13 13 3 0 16 0 3 2 13 10 9 7 13 9 2 16 10 9 13 13 10 0 2
4 13 3 3 2
6 15 13 3 13 9 2
10 11 9 3 0 13 9 13 13 11 2
4 2 13 3 2
8 3 15 9 1 9 13 15 2
19 0 9 9 0 9 13 13 0 0 9 2 10 9 13 9 7 9 3 2
3 3 0 9
17 13 13 3 13 9 1 9 0 9 7 16 2 3 10 0 9 2
15 13 3 2 13 10 9 3 7 13 3 15 1 10 9 2
12 10 9 13 13 0 2 7 15 13 3 0 2
5 15 15 13 13 2
5 15 13 9 13 2
3 8 8 0
5 16 13 9 13 2
3 13 3 2
10 13 9 13 2 3 13 15 13 13 2
11 15 9 11 13 13 9 3 2 7 15 2
2 9 13
4 9 15 9 13
5 13 3 9 13 2
13 15 13 9 0 9 2 0 2 0 9 0 9 2
12 15 13 10 11 3 13 15 13 3 3 11 2
6 15 13 15 9 13 2
5 9 13 9 1 2
6 15 13 13 15 0 2
6 13 9 11 2 16 2
8 15 13 9 1 0 9 1 2
8 15 3 13 13 3 13 15 2
4 11 13 9 2
13 3 15 13 13 3 9 2 7 15 13 13 15 2
8 2 11 2 13 9 9 11 2
2 9 2
13 16 9 3 13 2 15 13 13 9 3 9 1 2
17 7 13 9 9 9 2 3 13 13 9 9 13 1 9 2 7 2
12 9 9 13 13 9 2 16 9 13 10 9 2
11 13 0 13 2 16 13 9 13 10 0 9
12 9 13 3 13 9 2 7 9 13 13 13 2
7 9 13 9 9 9 0 2
3 13 9 13
17 16 13 2 16 13 11 3 0 9 9 1 2 9 13 13 9 2
12 16 15 13 9 15 2 15 13 15 3 15 2
13 3 13 0 3 3 3 12 2 12 7 12 9 2
6 3 3 13 13 9 2
8 13 9 13 9 13 11 13 2
8 13 13 2 16 15 13 9 2
11 9 7 10 9 13 9 13 3 9 13 2
3 12 9 0
4 9 13 9 2
21 9 13 9 7 9 13 15 1 2 13 13 13 9 15 1 2 0 2 7 13 2
5 0 13 11 9 2
13 3 10 9 9 9 13 3 9 13 3 0 9 2
3 9 3 2
34 3 3 13 10 9 2 3 3 3 16 13 0 9 3 3 3 3 13 9 6 3 6 3 15 13 13 8 7 3 9 1 10 9 2
7 0 1 13 0 13 13 2
5 15 13 13 9 2
8 3 13 9 7 3 9 1 2
25 9 13 9 3 3 2 3 9 13 13 7 3 15 1 13 2 9 7 13 9 9 7 9 9 2
5 9 13 9 9 2
2 3 15
19 13 9 11 13 9 3 10 9 16 11 2 13 13 7 13 0 0 9 2
7 15 1 13 0 9 9 2
17 15 3 9 13 13 0 9 1 13 2 9 10 9 13 0 9 2
11 9 7 9 13 13 0 9 13 9 9 2
22 15 3 13 16 13 13 0 9 16 15 13 3 13 7 3 15 3 13 16 13 15 13
15 11 13 9 9 9 9 9 0 9 13 11 0 9 9 2
3 9 13 13
13 11 15 13 13 13 16 3 13 13 0 3 9 2
5 15 15 15 13 2
13 15 13 13 15 13 15 9 7 13 15 3 3 2
6 11 13 16 13 0 2
9 3 13 3 13 2 3 9 13 2
9 15 13 2 7 13 13 15 11 2
6 13 13 3 12 9 2
8 15 13 13 11 2 10 9 3
7 15 13 13 9 12 9 2
3 9 13 9
7 3 13 3 13 13 0 2
11 9 13 13 13 9 7 13 15 9 9 2
3 3 9 2
8 10 9 1 11 9 13 11 2
11 13 10 9 9 3 10 3 0 9 13 2
5 15 13 10 9 2
6 9 13 0 9 13 2
5 11 13 11 9 2
11 15 3 13 13 2 16 9 13 13 9 2
8 3 9 9 13 13 0 9 2
7 13 12 9 13 9 3 2
4 6 13 15 0
15 13 15 13 3 0 9 3 9 2 7 15 2 11 13 2
6 15 13 3 3 9 2
3 9 9 2
15 15 2 13 9 9 7 10 9 13 2 13 13 13 9 2
5 15 13 15 13 2
4 15 13 3 2
4 3 13 9 2
5 9 9 13 3 2
15 16 13 13 10 0 9 2 3 13 9 9 10 13 9 2
7 13 9 13 9 7 9 2
4 13 12 11 2
14 3 13 13 3 2 16 9 7 9 9 13 3 9 2
27 11 9 11 13 9 9 2 16 3 10 9 13 9 10 9 1 2 3 10 0 9 7 9 13 7 3 2
2 0 15
15 3 0 13 10 9 2 16 9 9 13 0 7 0 9 2
7 13 3 13 12 9 9 2
15 7 3 13 3 13 9 2 3 9 13 15 1 0 9 2
8 10 9 13 9 7 9 9 2
5 11 7 11 13 15
4 9 13 9 2
8 15 13 13 7 13 9 9 2
5 13 9 0 9 2
17 9 9 13 9 13 9 9 3 1 9 7 15 13 12 9 9 2
10 11 9 13 13 9 9 13 3 9 2
7 9 13 3 16 13 13 2
7 9 13 9 3 9 9 2
16 15 13 0 9 3 2 3 13 2 15 15 13 10 9 3 2
9 9 1 11 13 2 16 9 13 2
13 9 13 9 9 7 9 2 3 13 3 0 9 2
16 11 13 13 0 13 9 2 15 1 15 13 13 9 11 9 2
9 9 9 9 13 13 9 9 8 2
12 13 3 9 13 3 0 9 16 3 2 0 3
9 11 9 13 2 15 3 3 9 2
16 3 3 16 11 13 13 9 2 10 9 1 13 3 0 9 2
7 0 9 9 7 12 9 2
9 13 15 13 13 15 15 3 3 13
4 13 11 11 2
6 15 13 13 3 11 9
7 9 13 3 12 9 9 2
7 13 15 10 9 16 3 2
17 13 15 2 16 15 13 10 7 9 9 16 9 13 16 0 9 2
7 11 9 13 13 0 9 2
16 7 1 0 15 13 13 9 2 7 3 15 3 13 3 9 2
16 15 13 0 9 2 3 0 7 0 2 7 15 13 13 13 2
5 3 11 13 15 2
9 9 13 2 9 13 13 3 3 2
13 3 13 11 2 3 13 0 9 2 9 2 9 2
5 11 13 9 9 2
4 9 13 9 2
6 13 13 0 9 11 2
8 9 13 9 13 9 0 9 2
17 15 13 3 9 2 15 7 13 9 7 13 9 13 9 0 9 2
5 9 9 13 10 9
6 11 9 13 13 10 0
4 3 13 3 0
5 12 9 1 13 11
15 3 15 13 15 15 1 2 16 15 13 9 3 9 13 2
4 9 13 13 2
7 3 13 3 13 13 9 2
9 15 13 0 16 9 13 13 9 2
5 15 3 15 13 2
17 16 15 13 0 9 7 9 7 9 2 15 13 10 9 9 1 2
4 9 13 9 2
22 9 0 9 9 7 9 2 0 9 13 12 9 0 9 7 13 15 9 9 9 1 2
6 9 13 3 0 9 2
10 9 2 9 0 9 2 13 15 13 2
13 15 13 13 7 13 9 7 15 13 9 9 9 2
10 9 13 3 3 2 7 13 9 0 2
20 3 13 13 3 11 2 15 10 0 0 9 13 13 9 7 15 9 9 1 2
9 9 9 9 11 13 9 15 1 2
6 0 9 9 11 13 2
10 9 13 9 13 15 3 3 10 9 2
13 11 9 13 3 3 0 9 16 3 11 9 9 2
10 12 11 13 9 9 13 11 9 9 2
5 13 3 3 3 2
3 0 0 9
2 3 11
5 15 13 10 9 2
3 0 9 2
3 13 3 3
5 13 9 9 1 2
6 13 3 13 12 9 2
9 9 1 3 13 3 3 0 9 2
2 0 9
6 11 13 15 13 0 9
16 9 9 9 9 15 13 15 2 16 9 13 3 13 9 9 2
4 3 13 15 2
10 15 13 0 7 15 13 13 0 9 2
11 0 9 13 3 12 9 13 9 11 9 2
12 9 13 13 7 9 13 3 15 2 13 3 2
2 13 0
12 9 9 2 11 2 13 3 9 3 12 0 2
4 15 13 13 3
14 9 7 9 13 9 1 3 15 2 15 13 13 9 2
10 9 13 9 9 1 9 15 10 9 2
7 10 9 9 13 3 15 2
9 9 13 15 15 1 2 6 6 2
5 15 13 9 9 2
7 3 15 13 2 13 13 2
3 9 0 9
13 9 13 9 2 9 2 15 13 0 7 0 9 2
5 9 13 0 9 2
6 15 13 10 0 9 2
4 15 13 15 1
6 3 13 13 0 9 2
10 16 11 13 3 0 9 13 11 9 2
3 0 9 9
11 11 13 11 2 16 11 9 9 13 9 2
11 3 12 0 13 3 0 9 9 9 9 2
13 3 9 9 13 3 2 13 11 0 9 13 9 2
3 9 13 13
10 13 13 0 9 2 15 9 13 13 2
17 9 13 3 3 2 16 9 13 13 13 9 2 13 13 15 13 2
6 13 3 10 0 9 2
3 13 9 1
6 9 9 1 13 0 2
10 15 13 9 9 10 9 2 1 9 2
6 13 13 15 12 9 2
2 13 13
7 9 13 0 9 0 11 2
14 9 13 3 11 7 3 11 3 3 8 7 9 11 2
12 3 13 13 10 9 2 15 15 13 10 9 2
13 0 7 0 9 13 3 0 9 16 0 0 9 2
4 15 13 3 0
9 13 9 9 1 13 9 9 9 2
9 2 15 13 13 15 3 12 1 2
2 0 9
8 9 13 3 0 16 3 3 2
15 9 13 15 15 7 13 3 9 0 9 13 7 13 13 2
15 13 3 15 2 16 3 0 9 2 10 0 13 13 9 2
11 7 15 13 3 9 2 3 15 13 15 2
18 13 2 15 13 2 13 2 15 13 2 7 3 13 13 15 10 9 2
12 11 13 9 1 3 0 9 9 16 10 9 2
11 13 13 9 2 16 13 13 13 3 3 2
3 11 0 9
9 0 0 9 2 15 13 13 9 2
5 3 15 3 13 2
5 11 13 13 9 2
10 10 9 13 2 7 3 10 9 13 2
7 13 9 3 3 9 9 2
2 9 2
7 3 13 13 0 0 9 2
8 13 15 9 16 13 3 10 9
15 11 9 11 13 12 10 0 10 9 2 15 13 9 3 2
7 3 3 3 9 13 13 2
11 3 13 13 2 7 3 9 13 15 13 2
15 10 9 3 3 13 0 9 15 16 3 3 10 0 13 3
3 0 13 3
15 9 2 9 2 9 2 9 2 9 2 12 0 9 13 15
10 9 11 11 13 12 9 9 9 11 2
4 12 9 13 0
11 9 11 9 13 0 2 7 9 13 0 2
12 13 9 9 13 3 0 2 16 13 0 13 2
5 2 15 13 9 2
6 10 9 13 13 9 2
5 11 13 9 9 2
31 13 13 9 0 9 15 2 3 3 2 12 9 1 0 11 13 9 9 9 13 13 9 3 13 0 2 9 2 9 1 2
4 10 9 9 13
16 11 0 9 13 11 2 15 13 3 0 16 11 7 12 0 2
9 11 13 13 11 9 7 13 13 2
12 3 13 13 3 15 9 2 7 13 13 13 2
11 13 13 13 7 13 2 3 0 15 13 2
9 9 13 3 3 2 3 15 13 2
2 9 9
6 3 3 13 13 9 2
24 9 15 13 3 3 2 11 3 13 10 11 9 7 2 9 15 13 11 3 3 13 10 2 9
6 9 13 13 11 11 2
6 13 11 12 0 9 2
3 3 3 2
9 13 15 3 9 9 13 2 3 2
4 13 9 13 2
13 0 9 9 13 9 13 0 12 9 11 11 9 2
5 13 15 13 9 2
18 3 3 10 9 12 13 11 13 9 2 7 13 13 15 0 9 12 2
4 13 15 11 2
17 12 9 2 9 2 3 12 9 2 13 15 1 9 0 9 1 2
5 13 13 10 9 2
3 13 13 2
8 3 13 13 9 1 13 9 2
2 13 9
5 9 15 3 9 13
4 9 13 9 2
19 13 2 16 13 7 13 3 13 9 7 9 3 7 13 0 9 7 9 2
19 15 13 3 0 2 3 3 3 9 13 2 9 16 13 9 15 3 13 2
9 9 13 3 13 12 3 3 12 2
6 13 15 10 10 9 2
8 3 15 13 13 9 7 13 9
6 3 0 0 0 0 9
15 9 9 1 13 0 9 2 8 7 9 7 0 9 9 2
6 9 9 13 3 15 2
8 13 10 9 1 13 15 9 2
7 15 3 13 3 0 9 2
7 9 9 13 0 9 9 2
4 3 9 9 2
2 9 9
9 9 13 15 13 13 0 9 9 2
7 13 15 3 9 7 9 2
4 15 13 3 3
2 9 11
10 13 9 2 16 13 3 13 13 9 2
14 12 13 0 9 11 13 9 13 0 9 9 0 9 2
3 3 0 2
6 9 0 9 13 9 2
11 9 13 2 16 9 13 0 9 3 9 2
15 6 2 6 2 13 3 2 11 13 7 13 9 12 9 2
8 15 9 1 13 13 9 9 2
8 3 3 9 15 13 0 9 2
4 10 9 13 15
12 9 13 3 9 2 10 9 13 11 7 9 2
33 16 15 13 10 11 7 11 9 3 3 15 3 13 9 1 3 3 3 10 11 10 9 3 0 9 13 3 13 12 11 13 9 2
3 13 9 2
5 15 13 3 3 2
5 15 13 15 13 2
12 11 13 0 9 2 15 13 9 7 9 13 2
5 2 13 16 15 2
2 9 11
8 3 16 15 13 13 9 9 2
9 3 13 15 2 15 3 13 9 2
3 9 3 2
5 3 13 9 0 2
8 11 9 13 3 13 0 9 2
6 9 13 9 13 9 2
4 9 13 13 2
8 15 13 13 2 15 3 13 2
4 6 16 0 2
10 15 13 0 9 7 13 15 9 1 2
6 9 1 9 13 0 2
2 0 3
15 7 9 9 13 13 0 2 3 9 13 13 3 9 1 2
10 13 9 13 13 9 9 7 13 9 2
9 11 1 11 13 9 1 0 9 2
10 12 9 9 13 9 9 2 15 0 2
10 3 11 13 2 16 10 9 13 3 2
8 9 13 9 9 7 13 9 2
5 15 13 3 9 2
2 13 9
11 3 0 0 9 13 13 13 13 15 9 2
9 0 13 9 13 9 13 7 13 2
11 13 13 2 3 13 0 13 13 10 9 2
5 11 13 15 3 2
4 0 13 13 2
5 2 6 15 13 2
9 9 13 3 16 9 13 9 9 2
7 15 13 13 0 0 9 3
3 13 15 13
7 15 13 3 9 9 9 2
2 13 13
15 3 16 13 16 16 13 10 0 9 15 13 3 3 10 9
16 9 13 9 1 9 3 13 9 13 15 9 13 9 7 13 2
18 7 15 13 13 2 16 10 3 0 13 9 3 15 1 16 13 0 2
14 9 13 3 10 9 0 16 10 9 3 2 11 13 2
8 9 9 13 0 2 0 9 2
12 9 13 9 2 16 9 13 9 12 12 9 2
6 10 9 13 10 9 2
4 9 13 3 0
8 13 3 3 13 9 13 9 2
3 13 3 2
5 9 13 13 9 2
2 3 3
2 13 9
17 13 13 3 0 9 2 10 9 13 2 16 13 9 2 13 9 2
19 9 9 9 13 9 11 13 13 15 0 7 0 7 3 0 7 0 9 2
10 13 9 2 7 15 13 11 11 9 2
7 10 9 9 13 15 9 2
5 13 15 9 6 2
14 16 11 13 9 9 2 13 10 9 9 13 3 0 2
13 7 13 3 3 15 2 16 9 13 0 13 3 2
10 15 13 13 2 16 9 13 9 1 2
9 11 13 15 15 13 3 9 1 2
12 16 11 9 13 9 2 11 13 13 9 13 2
23 3 15 13 11 7 11 7 10 11 7 2 11 7 2 15 3 13 11 7 3 2 13 3
2 15 13
3 13 15 2
6 15 13 3 9 7 9
3 13 13 13
13 0 9 10 15 2 15 3 13 13 9 7 9 2
18 15 13 3 0 9 15 2 16 3 7 0 9 13 3 13 10 9 2
12 9 13 13 0 9 2 16 13 9 13 9 2
3 9 13 13
14 3 13 3 0 9 3 16 16 9 13 13 3 13 2
9 0 0 9 13 13 9 0 9 2
8 9 13 12 2 12 7 12 2
4 10 10 0 9
18 16 3 3 13 0 9 13 9 2 13 16 9 13 7 0 9 13 2
10 11 13 13 2 3 13 13 3 3 2
15 0 9 11 7 10 9 1 13 13 3 11 0 9 1 2
2 3 0
13 11 9 11 11 9 9 9 13 9 13 3 9 2
13 11 0 9 9 13 3 0 9 0 0 7 0 2
10 9 13 9 2 15 13 13 7 13 2
8 9 13 13 2 16 13 3 13
14 7 15 2 15 1 10 9 13 2 13 10 0 9 2
13 15 13 13 2 11 13 2 16 9 13 13 9 2
2 13 13
6 2 13 3 0 9 2
10 9 13 9 1 13 13 12 12 9 2
4 9 13 9 2
7 15 13 3 11 9 9 2
13 3 13 1 0 9 7 3 13 13 3 0 9 2
6 0 10 10 9 3 2
5 9 13 9 1 2
16 13 11 13 3 13 3 11 2 3 3 2 3 0 15 13 2
11 9 13 3 13 2 16 9 13 9 9 2
2 13 9
6 10 9 9 13 11 2
6 3 15 15 3 13 2
11 0 9 11 7 10 9 11 13 0 9 2
5 0 9 13 0 2
6 10 9 13 9 9 2
11 11 9 13 13 9 2 16 3 9 13 2
3 9 13 9
2 0 9
9 13 13 12 9 13 9 9 13 2
3 11 9 0
17 13 13 3 12 9 13 15 3 13 11 3 7 16 13 3 3 2
8 3 13 13 13 9 13 15 2
15 13 15 13 15 2 2 3 9 13 13 9 9 9 2 2
11 12 9 13 15 0 2 9 2 7 9 2
2 10 9
9 3 3 0 9 13 13 13 13 2
4 9 9 2 12
11 0 9 13 13 3 13 9 13 2 16 2
8 9 9 13 13 2 13 9 2
19 11 9 13 13 9 9 2 9 13 9 7 9 7 9 13 0 0 9 2
10 9 11 3 13 11 13 13 0 9 2
5 0 9 13 9 2
6 9 11 7 11 13 11
18 3 3 9 9 13 11 9 13 11 0 2 16 15 13 11 10 11 2
5 13 3 9 3 2
3 13 9 2
12 11 13 13 13 10 9 9 1 9 9 9 2
8 11 13 13 15 13 0 9 2
15 9 13 9 9 13 9 13 9 1 3 9 3 0 9 2
11 15 13 9 2 7 15 13 3 3 9 2
4 13 9 12 2
12 3 10 11 0 9 13 13 9 9 13 11 2
8 11 13 12 0 9 9 9 2
2 9 1
11 13 3 10 9 16 15 13 9 3 13 2
14 15 13 0 9 3 3 2 16 13 9 13 0 13 2
6 13 3 13 3 0 2
17 13 0 9 13 9 7 9 2 16 13 10 9 3 3 3 0 2
4 13 15 9 2
17 15 13 13 3 0 13 15 13 13 16 15 13 0 0 7 0 2
6 11 13 0 9 9 2
10 9 13 13 10 12 0 9 13 9 2
5 11 13 9 9 2
6 10 15 13 3 9 2
3 12 9 9
10 13 13 3 9 2 15 10 9 13 2
5 0 9 9 6 2
3 3 3 0
3 3 13 9
5 13 7 13 13 2
5 13 0 13 10 9
13 3 12 9 1 13 0 2 16 13 9 13 3 2
9 3 11 0 9 13 13 3 9 2
8 9 11 13 13 0 1 9 2
8 9 13 3 9 11 9 9 2
6 6 13 3 13 13 2
9 9 1 11 13 7 13 13 3 2
20 7 3 13 13 13 9 9 3 7 3 13 3 2 13 9 7 13 9 9 2
9 11 9 7 11 13 11 16 15 2
5 9 13 3 0 2
6 9 13 12 0 9 2
11 16 9 13 13 3 3 3 2 16 15 13
10 10 9 15 13 12 9 9 3 9 2
12 0 9 7 0 3 13 9 13 13 3 9 2
9 11 13 10 9 15 3 9 9 2
4 10 9 13 2
6 3 13 8 13 3 2
13 9 9 9 12 13 12 9 9 9 9 9 11 2
10 11 9 11 1 9 13 13 13 13 2
9 13 15 13 10 9 7 9 13 2
3 12 9 0
4 0 9 7 9
10 13 15 9 2 15 13 3 13 9 2
9 9 13 9 13 13 13 0 9 2
6 9 13 9 13 9 2
17 13 3 13 2 16 15 13 13 9 13 13 13 9 9 0 9 2
10 13 15 9 13 7 13 2 13 11 2
5 3 13 12 9 2
4 9 13 3 13
6 3 15 13 3 9 2
20 13 13 15 2 16 9 13 13 3 16 11 9 7 13 16 13 3 15 9 2
8 9 7 10 9 13 3 9 2
7 13 13 9 3 9 9 2
6 9 9 13 3 9 2
14 9 13 0 9 2 10 9 13 13 2 13 3 9 2
7 3 10 9 13 9 3 2
6 13 9 3 13 13 2
12 13 15 3 3 3 13 13 2 10 9 13 3
12 11 9 13 12 11 7 3 11 9 9 9 2
8 12 9 13 0 9 11 9 2
15 9 13 13 13 2 16 9 13 0 9 9 9 3 11 2
6 15 1 13 13 3 2
7 13 3 11 9 13 0 2
2 0 9
10 9 1 7 9 1 15 13 13 9 2
8 9 13 0 9 11 11 9 2
13 3 13 0 13 2 16 11 9 13 3 3 0 2
17 3 11 7 3 11 13 0 9 2 7 13 13 9 9 13 11 2
8 15 13 13 3 0 0 9 2
16 11 7 11 9 13 3 9 9 13 11 2 15 9 13 13 2
18 9 0 9 13 0 2 3 3 9 2 9 2 11 7 11 3 11 2
3 13 3 2
3 9 13 9
6 9 13 15 13 9 2
11 9 13 15 13 11 2 7 13 3 9 2
14 9 9 13 13 9 13 9 9 2 9 7 9 9 2
7 13 15 3 12 9 13 2
4 13 0 9 2
13 10 15 13 13 13 9 15 13 3 7 13 9 2
3 13 0 9
9 9 3 9 13 9 13 0 3 2
5 3 13 0 9 2
13 3 9 15 13 2 16 13 3 13 15 15 1 9
5 2 0 13 9 2
6 9 1 9 9 13 2
4 3 13 0 9
7 6 3 15 13 13 3 2
15 11 13 13 2 16 3 3 11 13 3 13 9 11 11 2
3 12 9 13
15 11 13 0 2 15 13 13 7 13 9 2 13 13 15 2
5 13 15 15 13 2
3 0 9 2
3 9 13 13
16 13 15 16 13 0 9 9 13 2 16 9 15 13 13 9 2
4 13 3 3 2
2 3 9
2 13 13
4 15 13 3 2
7 13 15 13 13 3 13 2
14 15 13 2 16 13 13 9 2 16 0 13 9 9 2
7 13 0 7 13 15 9 2
8 0 9 13 13 9 16 0 2
6 15 13 13 3 0 2
5 13 3 0 9 13
15 10 9 1 0 9 13 13 9 2 3 16 15 13 3 2
2 10 9
11 9 13 9 0 9 13 15 9 0 9 2
5 15 13 0 9 2
6 9 1 13 9 9 2
4 13 15 9 2
9 13 9 9 13 12 9 9 9 2
15 16 15 10 9 13 13 9 2 9 9 13 11 0 9 2
6 11 13 9 3 9 2
14 3 15 13 0 16 9 2 16 3 10 9 13 9 2
22 9 12 13 11 9 11 13 9 1 9 0 9 2 16 9 13 9 11 1 0 9 2
2 13 13
5 15 13 9 12 2
6 15 13 2 15 13 2
14 15 13 3 13 3 3 2 15 2 13 9 9 2 2
4 3 0 9 2
14 9 13 9 7 9 9 2 3 13 3 11 9 9 2
4 9 13 10 12
3 13 13 15
5 0 9 13 9 2
9 12 9 9 11 11 13 0 9 2
7 3 15 15 15 0 13 2
15 10 9 9 9 2 9 2 9 2 9 13 11 11 9 2
5 15 1 15 13 2
10 15 13 13 0 3 3 11 13 11 2
6 15 13 9 11 11 2
3 9 7 9
3 9 15 13
12 10 9 16 9 13 2 3 15 13 10 9 2
13 10 9 13 13 9 11 13 9 0 0 9 9 2
7 9 13 9 12 9 1 2
8 12 9 1 9 13 9 1 2
6 13 9 13 9 1 2
11 11 13 13 9 2 7 3 10 3 0 2
8 15 13 0 2 16 13 11 2
7 0 9 9 11 7 11 11
8 0 9 13 3 0 9 9 2
2 15 13
9 15 13 0 2 3 16 13 13 2
2 10 0
18 9 10 9 13 0 11 2 0 9 13 0 11 8 7 0 8 9 2
12 9 13 0 9 2 13 10 0 9 9 3 2
16 3 3 15 13 9 0 9 7 15 9 9 2 15 13 15 2
15 15 13 3 0 9 7 10 9 13 13 9 9 1 9 2
16 11 11 13 13 3 10 10 9 2 0 15 9 13 13 13 2
9 9 1 9 13 0 9 7 9 2
13 9 13 9 9 2 3 9 9 7 0 9 9 2
4 15 3 13 2
9 3 13 11 3 0 9 7 0 9
9 11 13 9 9 3 3 2 16 2
9 3 13 3 13 7 13 0 13 2
12 7 15 15 9 13 2 13 2 0 9 2 2
12 9 13 13 9 9 2 15 15 13 0 9 2
7 3 13 2 16 13 9 2
8 9 13 9 9 7 15 9 2
14 9 7 9 7 12 9 13 13 0 9 3 11 11 2
4 3 13 13 9
15 9 9 13 12 9 2 10 9 3 10 0 9 13 0 2
6 13 13 9 3 9 2
13 13 7 13 0 9 13 9 9 12 9 9 2 2
6 15 13 2 13 9 2
4 13 3 15 2
4 13 13 15 2
7 13 13 3 9 12 1 2
10 13 13 13 7 13 0 0 9 9 2
10 9 13 9 11 13 12 0 9 1 2
3 9 9 9
10 9 13 0 9 13 3 9 9 9 2
7 3 15 13 15 0 9 2
5 9 13 12 9 2
5 3 15 13 9 2
5 11 11 13 13 2
11 13 13 15 7 2 13 9 0 0 9 2
2 13 2
4 13 9 12 2
8 13 13 9 9 9 9 3 2
8 15 13 9 9 9 7 13 2
7 12 9 0 12 9 13 9
9 16 13 13 3 3 2 13 13 3
11 0 13 3 13 2 16 9 13 0 9 2
5 13 15 11 10 9
7 9 12 9 13 0 3 2
3 13 13 9
8 3 9 13 9 13 3 9 2
8 11 11 13 11 9 12 9 2
8 13 16 13 0 9 0 9 2
4 13 15 13 2
3 9 0 9
4 13 15 9 2
7 11 7 11 13 11 9 2
3 3 10 15
4 13 13 0 2
2 9 1
9 2 3 13 2 15 13 3 3 2
16 0 9 1 13 3 0 9 0 9 2 0 9 7 0 9 2
11 2 15 13 3 9 0 2 7 0 2 2
4 0 9 9 9
16 3 0 9 13 13 12 9 3 2 16 13 13 13 3 3 2
7 13 3 2 3 13 13 2
3 9 0 9
12 9 13 3 13 13 9 12 0 9 11 9 1
7 15 13 2 16 13 9 2
13 15 13 13 9 0 9 1 2 15 11 13 13 2
16 13 13 2 7 15 13 13 15 16 13 13 13 7 3 13 2
16 9 13 13 9 9 12 2 7 0 9 13 13 13 9 12 2
11 9 13 9 13 13 12 9 9 9 1 2
5 15 13 3 9 2
5 11 13 11 9 9
3 13 13 2
5 9 13 13 9 2
3 11 11 1
13 16 7 16 9 13 9 2 9 13 0 9 9 2
6 15 1 15 13 9 2
4 3 13 9 3
13 3 0 9 13 3 13 16 11 9 13 9 9 2
11 13 15 2 16 9 13 13 3 3 3 2
7 9 1 15 13 13 3 2
4 13 13 3 2
5 15 13 0 13 2
52 9 1 2 15 13 13 0 0 8 7 9 9 2 13 2 16 15 1 13 9 13 0 3 3 9 13 7 9 3 0 9 3 9 9 7 9 2 13 9 2 10 9 9 1 13 9 3 9 13 0 9 2
3 9 13 13
3 13 13 9
2 13 9
7 13 9 9 9 1 9 2
9 13 13 10 9 3 9 7 3 2
7 15 13 13 9 13 9 2
18 13 3 3 0 2 16 15 13 3 13 9 9 2 16 13 13 0 2
5 9 13 9 0 2
6 13 15 0 15 13 2
8 15 15 13 13 15 13 15 2
5 11 13 9 1 2
6 11 0 9 13 9 2
16 13 9 9 13 13 2 7 3 10 9 13 3 13 9 9 2
5 15 13 15 9 2
7 13 0 7 0 9 1 2
11 9 13 3 12 9 7 9 13 9 9 2
11 13 11 9 11 7 3 15 1 11 11 2
13 7 13 0 2 15 13 16 13 15 3 0 13 2
5 0 9 13 13 2
11 3 16 0 9 3 13 10 15 7 15 2
18 11 13 13 0 2 16 3 15 15 3 13 13 15 13 13 15 9 2
13 13 15 2 16 11 13 3 13 2 0 2 9 2
5 11 13 3 3 2
4 13 15 9 2
7 15 1 13 3 9 9 2
3 10 9 0
9 0 11 11 9 9 13 9 11 9
7 9 13 15 13 9 13 2
7 13 9 3 11 9 9 2
8 10 15 13 13 10 9 9 2
3 9 3 2
17 3 1 0 11 13 11 9 13 2 15 3 15 13 9 9 12 2
4 13 11 13 2
4 15 13 11 2
5 13 10 3 9 2
5 13 15 13 9 2
11 13 9 13 15 13 0 9 11 11 9 2
9 3 15 3 3 13 3 3 3 2
10 3 9 13 0 2 10 9 3 0 2
13 13 3 3 11 7 13 2 16 15 13 0 9 2
3 13 3 9
3 13 9 9
8 3 15 13 0 16 3 3 2
16 9 13 2 16 0 13 3 9 0 9 16 10 11 9 9 2
12 15 13 13 9 2 16 12 9 13 13 15 2
7 10 9 13 11 0 9 2
4 13 13 13 2
3 9 13 2
17 15 13 3 0 9 2 15 13 0 7 0 9 2 9 7 9 2
7 13 10 9 1 3 9 2
17 9 13 3 13 12 12 9 1 12 9 13 3 12 9 0 9 2
16 9 13 0 9 7 15 13 13 3 3 16 11 13 9 13 2
6 9 13 0 13 9 2
6 10 9 13 9 13 15
8 15 13 9 2 9 2 9 2
4 9 13 15 2
4 13 13 9 2
4 9 9 13 9
6 10 15 13 3 9 2
4 10 10 0 9
9 10 9 9 9 13 0 11 11 2
7 15 13 13 9 9 1 2
12 3 11 13 15 2 15 13 9 9 9 11 2
5 13 15 3 3 2
13 11 7 11 13 9 9 13 9 3 16 13 9 2
14 13 2 16 11 3 13 2 7 0 9 13 3 13 2
6 15 13 3 1 15 2
10 9 13 2 16 9 13 15 13 3 2
5 13 15 15 13 2
8 11 9 9 13 3 13 13 2
60 3 3 3 13 3 15 13 3 2 3 10 10 9 2 9 1 7 2 7 3 13 3 16 16 3 3 10 0 9 9 3 13 13 3 2 3 3 2 3 10 10 9 3 3 3 16 11 16 3 2 16 3 15 13 13 13 15 13 16 2
7 9 9 13 3 13 9 2
8 9 13 0 7 9 9 13 2
13 3 13 3 10 9 15 13 13 13 15 2 16 2
2 13 3
5 13 3 9 9 2
9 15 13 16 11 9 13 10 9 2
10 16 9 13 2 9 13 0 9 13 2
13 13 3 0 16 9 13 9 7 13 16 10 9 2
11 10 9 13 13 9 2 15 13 15 0 2
6 9 13 9 9 3 2
11 15 13 13 10 9 2 15 9 13 0 2
9 2 7 16 13 2 2 9 13 2
5 16 13 11 13 2
6 12 9 13 13 13 2
8 11 7 11 13 9 0 9 2
2 10 9
6 3 13 9 7 9 2
7 15 13 9 11 12 9 2
5 13 15 10 0 2
6 15 13 13 13 13 2
3 15 13 0
9 15 13 9 9 13 0 12 9 2
4 11 9 0 2
9 2 3 3 13 2 6 15 0 2
7 9 13 13 9 3 3 9
6 9 13 9 1 3 2
5 15 15 15 13 2
14 13 9 1 13 0 9 10 0 9 16 10 9 9 2
3 13 3 2
15 7 15 13 13 3 3 2 16 15 13 3 9 10 9 2
5 9 13 13 0 2
12 11 1 9 13 13 10 9 9 7 9 13 2
7 9 13 9 13 3 9 2
4 13 15 0 2
2 0 9
8 6 3 9 15 13 13 13 2
11 3 10 0 7 0 9 13 9 13 15 2
8 13 9 7 9 9 8 8 2
4 9 0 9 9
15 9 13 15 2 16 9 13 9 9 1 13 9 3 11 2
6 15 13 3 0 13 2
24 7 11 13 3 10 10 9 13 9 2 15 3 13 15 0 9 13 15 9 3 7 9 9 2
10 13 15 13 10 9 3 2 11 13 2
5 11 13 13 9 2
10 10 0 0 13 9 10 10 9 13 2
11 9 13 0 2 16 13 3 2 11 13 2
10 15 13 13 2 16 13 13 9 9 2
7 9 8 7 0 9 7 9
12 3 9 13 0 13 13 0 7 0 9 15 2
10 11 13 3 0 9 9 7 10 9 2
4 13 9 9 2
14 9 13 13 2 7 13 9 13 9 12 9 1 9 2
4 11 9 0 9
3 9 13 13
10 3 15 13 10 9 3 12 9 3 2
10 15 13 2 16 9 13 13 9 9 2
5 13 15 15 13 2
5 3 12 0 9 2
3 15 9 2
3 9 11 1
10 7 15 15 13 3 10 9 13 3 3
8 15 13 3 3 3 10 9 2
16 7 15 9 3 3 16 15 13 2 13 3 3 16 13 9 2
9 15 13 13 16 9 9 13 13 2
6 9 13 3 3 9 2
10 15 13 3 13 7 9 13 9 1 2
11 9 9 2 15 15 13 10 0 0 9 2
3 15 13 9
4 15 13 3 2
7 15 13 9 9 3 3 2
20 15 13 0 9 9 2 3 13 9 2 0 15 2 11 13 2 13 10 9 2
5 9 13 9 0 2
11 15 13 3 3 7 13 9 2 13 11 2
6 15 13 3 9 1 3
15 9 13 2 7 3 13 9 13 0 2 16 13 3 13 2
10 11 13 13 16 0 9 7 9 13 2
10 11 13 2 3 10 9 13 13 13 2
11 15 13 9 1 7 13 3 9 0 9 2
20 10 3 0 15 13 13 3 2 9 9 2 9 2 9 2 9 7 0 9 2
8 11 13 9 3 7 9 9 2
9 3 9 9 9 9 13 3 0 2
6 13 3 9 11 11 2
13 15 13 3 13 9 7 9 7 15 13 9 3 2
4 13 15 13 3
24 15 13 9 2 9 2 9 2 9 2 9 2 9 13 2 9 13 2 9 13 2 9 13 2
14 13 13 2 16 0 13 0 2 16 0 13 13 0 2
5 15 13 13 13 9
14 2 13 3 0 9 13 2 13 13 9 2 13 9 2
8 16 13 9 1 9 9 13 2
10 15 1 15 13 2 16 15 13 15 2
7 9 9 13 7 9 13 2
12 11 13 13 15 9 2 16 13 9 9 9 2
2 13 9
10 15 13 9 2 15 13 3 9 9 2
16 0 13 2 16 0 9 7 9 13 3 9 13 13 15 13 2
8 15 15 13 2 9 7 9 2
4 15 13 16 9
4 15 13 12 9
7 9 13 13 13 9 13 2
16 13 15 2 13 13 2 11 11 13 0 7 0 9 0 13 2
5 9 9 2 11 13
5 3 13 9 9 2
14 9 1 11 11 13 13 2 16 15 13 3 3 11 2
10 11 9 13 9 0 12 12 9 9 2
13 12 7 12 9 13 13 2 13 2 13 2 13 2
7 3 0 1 9 13 13 2
7 3 10 11 9 13 9 2
8 9 13 3 9 9 12 9 2
14 16 3 13 9 13 13 13 2 16 0 9 11 13 2
10 9 9 13 9 13 9 2 7 3 13
10 9 13 9 2 16 13 13 11 9 2
12 3 0 16 15 13 2 9 13 13 13 9 2
3 11 13 9
2 9 9
2 6 2
7 9 13 3 13 9 9 2
6 15 13 3 1 9 2
15 3 15 9 13 16 9 2 13 9 9 13 0 9 9 2
8 9 13 10 9 11 11 1 2
3 13 15 2
2 13 9
7 9 15 1 13 3 13 2
5 13 9 0 9 2
5 9 3 3 0 9
8 15 13 13 9 13 13 9 2
10 9 13 0 2 7 13 3 10 9 2
2 9 13
5 13 15 13 9 2
8 13 13 9 13 13 0 13 2
3 9 3 2
7 7 13 13 10 9 9 2
3 0 9 2
14 15 3 16 9 13 9 13 13 3 9 9 13 9 2
8 11 13 3 13 3 3 9 2
3 9 13 9
5 10 9 15 13 2
3 0 11 11
16 13 13 9 3 9 2 9 2 9 9 2 9 7 1 9 2
7 9 13 9 13 9 12 2
3 15 13 9
31 11 9 10 0 9 3 13 12 9 9 10 0 9 13 0 13 9 9 13 10 9 13 13 7 13 0 9 9 9 11 2
7 11 13 3 13 9 9 2
8 3 13 2 15 9 13 13 2
12 13 3 2 9 2 11 13 3 7 13 11 2
3 9 9 3
7 13 11 9 2 9 13 2
11 10 9 13 13 13 9 9 7 9 9 2
12 15 13 3 9 2 13 9 13 3 0 9 2
15 13 3 2 13 15 13 2 13 3 9 7 13 0 0 2
7 9 9 13 3 12 9 2
7 13 9 13 7 9 13 2
7 15 15 3 13 13 13 2
11 11 13 13 2 16 13 10 9 13 0 9
5 0 9 15 13 2
7 9 13 13 12 9 1 2
24 16 13 9 13 2 3 10 9 13 2 7 3 13 13 2 0 9 2 2 3 9 13 13 2
13 13 13 9 11 9 3 2 16 15 13 3 13 2
9 13 3 9 7 3 3 16 15 2
2 0 0
16 0 9 13 0 2 16 9 7 15 9 9 13 3 9 9 2
10 13 3 3 13 11 7 15 0 9 2
9 9 9 9 9 13 11 9 11 2
6 13 3 13 15 3 2
4 15 3 15 13
30 16 3 13 3 7 13 15 15 2 13 9 2 10 2 3 15 9 15 2 3 15 13 3 2 15 13 15 9 9 2
15 3 0 9 13 9 2 15 15 13 13 9 13 9 9 2
6 15 3 13 0 9 2
8 10 9 13 3 0 9 9 2
5 15 13 9 15 2
24 3 15 13 3 10 9 3 7 10 10 9 13 10 9 15 13 16 16 15 13 9 0 9 2
4 3 3 13 2
8 9 13 13 9 9 2 7 2
14 15 9 9 13 13 16 15 13 3 2 0 7 0 2
9 9 9 13 9 13 11 11 12 2
8 15 13 10 11 7 11 9 3
4 15 13 9 2
9 15 3 13 10 9 16 15 13 13
11 13 13 2 16 11 13 9 0 9 1 2
2 6 3
5 3 15 3 9 2
10 13 0 2 16 9 13 2 3 13 2
4 15 13 3 2
11 7 0 13 13 2 7 3 15 13 0 2
11 11 13 13 9 9 13 0 9 11 9 2
6 13 10 9 12 9 2
5 13 15 13 13 2
11 0 9 13 13 13 9 13 9 9 9 2
15 9 13 3 2 16 10 13 13 9 13 13 15 15 9 2
3 3 0 2
17 16 13 9 9 9 2 9 13 16 3 3 13 15 15 13 13 2
5 9 13 9 13 9
9 13 13 3 2 7 15 13 15 2
4 13 13 9 2
16 9 9 9 13 13 2 7 10 9 9 13 3 10 12 9 2
7 15 3 13 9 3 9 2
20 12 0 9 0 9 2 16 15 13 13 3 3 0 9 2 7 3 3 3 2
10 9 13 9 2 16 15 13 3 3 2
4 9 13 9 2
3 10 12 9
2 0 9
19 9 13 0 13 9 2 7 15 13 0 0 13 2 16 13 7 13 9 2
13 15 13 3 3 16 15 13 7 13 11 15 3 2
9 11 9 13 9 12 7 12 9 2
4 15 13 9 2
6 13 9 7 13 15 2
11 9 13 13 0 0 2 16 15 13 3 2
12 9 13 9 1 9 13 0 2 7 13 0 2
10 3 13 13 13 0 0 9 3 9 2
11 9 13 3 9 9 2 15 13 7 13 2
5 13 13 13 13 2
6 3 15 13 10 3 2
8 3 15 3 13 16 0 9 2
12 15 13 13 15 7 13 9 9 10 0 9 2
4 9 13 9 2
6 13 9 9 7 9 2
10 3 13 3 3 1 9 10 0 9 2
5 3 13 3 9 2
2 3 0
4 13 3 3 2
6 15 13 3 13 0 2
13 11 7 10 9 13 9 3 7 13 11 1 9 2
5 13 13 9 12 2
10 11 9 13 13 3 9 2 11 13 2
6 9 13 9 9 11 1
8 2 7 13 9 9 10 9 2
10 10 10 9 0 9 7 9 0 9 2
16 9 0 9 11 13 13 13 13 9 2 16 15 13 15 13 2
7 11 13 3 0 11 9 2
5 11 13 11 0 9
5 10 9 13 0 2
3 9 13 13
16 9 9 7 9 9 9 13 3 3 2 16 11 13 3 0 2
9 13 9 13 3 3 0 9 1 2
10 13 9 9 1 3 2 16 15 13 2
14 9 13 3 13 3 9 2 9 2 9 9 7 9 2
10 13 3 13 10 9 2 7 13 3 2
12 9 13 9 3 3 16 15 13 9 7 9 2
10 7 16 15 13 13 2 3 10 0 2
3 13 9 1
19 13 15 16 15 13 9 7 9 7 9 7 9 7 9 7 9 7 9 2
3 12 9 9
13 16 13 3 9 2 3 15 13 10 9 1 9 2
7 13 15 9 7 15 9 2
7 3 3 11 13 0 9 2
7 9 7 9 13 13 3 2
8 11 9 13 9 9 13 0 2
5 13 13 0 9 2
4 9 3 13 9
7 13 3 13 13 3 9 2
4 0 15 13 13
14 15 3 13 13 9 9 2 7 1 10 10 0 9 2
5 15 13 0 9 2
10 0 11 13 9 13 9 9 9 9 2
4 13 13 13 2
5 3 3 9 13 2
20 15 13 9 10 0 9 2 15 13 13 2 16 10 9 9 0 9 13 0 2
11 9 13 3 13 9 2 15 13 9 13 2
4 3 9 13 2
12 3 9 13 13 13 2 15 13 13 0 9 2
12 13 15 1 2 16 13 15 13 13 0 9 2
4 3 9 13 2
5 3 9 13 0 2
2 9 0
15 15 13 9 7 9 7 13 16 15 13 3 10 9 9 2
6 9 9 13 3 0 2
8 9 13 3 16 13 3 13 2
10 0 9 9 13 11 13 9 9 1 2
13 3 3 3 9 9 13 3 3 0 16 0 9 2
6 15 13 3 9 1 3
10 13 13 9 9 3 3 12 9 1 2
8 10 9 13 3 12 9 1 2
7 3 0 9 3 3 13 2
7 9 13 3 3 10 9 2
7 3 9 13 10 9 13 2
6 11 13 9 9 9 2
3 12 9 0
5 13 3 13 9 2
14 3 15 13 13 15 9 7 9 2 16 13 0 9 2
11 11 13 0 10 12 2 15 13 3 3 2
2 9 1
6 10 9 15 3 13 2
7 11 13 13 3 11 9 2
6 0 9 13 0 9 2
9 13 3 13 9 2 15 13 9 9
2 0 9
2 9 9
5 15 13 3 9 2
6 3 13 13 13 15 2
5 9 13 0 12 2
13 9 13 0 7 0 9 9 2 9 7 3 13 9
6 15 13 16 13 15 2
5 3 15 13 9 2
16 10 9 13 9 2 9 3 7 9 3 2 15 13 3 3 2
5 9 13 13 3 2
6 3 13 13 13 3 2
9 11 9 13 9 7 9 13 9 2
3 11 3 13
11 9 13 0 0 9 9 13 3 0 9 2
13 15 13 13 10 9 1 2 3 0 16 15 13 2
3 9 13 9
14 10 9 13 2 16 9 13 13 13 13 13 9 9 2
8 13 13 10 10 9 13 9 2
5 9 9 13 0 2
7 9 13 3 11 1 11 2
20 11 9 11 2 15 13 9 9 0 9 2 13 15 13 13 3 3 0 9 2
11 13 0 2 16 15 13 10 9 2 13 2
3 15 13 0
4 9 13 3 2
4 13 3 3 13
16 13 0 9 9 15 15 13 10 9 2 13 15 15 13 9 2
9 3 3 3 9 13 13 3 9 13
13 12 9 13 3 9 1 9 2 12 9 3 9 2
13 2 15 13 13 7 13 7 13 9 7 3 13 2
3 12 0 9
4 6 15 13 2
9 9 9 13 9 7 11 7 11 2
8 9 13 13 9 0 0 9 2
2 9 9
7 13 13 0 3 16 9 13
7 0 9 2 13 0 9 0
12 9 9 11 11 2 2 9 9 13 13 9 2
11 10 0 9 13 2 3 0 9 13 9 2
5 3 15 15 13 2
4 13 13 15 3
9 9 13 9 12 9 13 3 12 0
2 6 6
2 0 11
4 13 15 3 2
5 9 13 15 0 2
12 11 9 13 12 9 1 3 0 11 11 9 2
21 15 13 13 11 2 16 3 15 10 9 13 2 13 7 13 2 16 13 9 3 2
4 9 13 15 1
7 15 13 9 13 10 9 2
11 0 9 13 2 16 9 13 9 9 9 2
10 9 13 13 0 2 7 3 0 9 2
15 3 11 11 13 9 11 11 0 12 9 1 11 13 9 2
12 10 9 13 3 9 9 13 9 9 9 1 2
6 15 13 3 12 1 2
9 3 0 9 13 9 7 9 9 2
10 9 13 9 9 13 13 3 10 9 2
13 0 9 11 3 13 2 16 11 13 15 13 3 9
9 3 11 7 10 12 9 13 9 2
8 9 13 9 9 7 9 9 2
11 15 1 11 13 3 0 7 0 9 9 2
3 9 13 15
19 9 1 15 13 15 12 0 9 2 15 13 9 1 11 9 7 11 9 2
11 15 13 3 16 13 0 9 2 9 13 2
17 12 9 12 13 12 9 2 15 11 7 12 10 9 13 9 1 2
12 13 15 15 15 13 16 15 13 10 9 9 2
3 0 9 1
2 0 11
7 9 13 13 3 0 9 2
16 3 13 13 16 0 0 9 2 3 10 9 0 9 13 3 2
9 11 13 7 3 0 7 0 0 2
7 13 12 9 9 13 9 2
14 15 13 0 9 7 13 3 13 2 16 15 13 13 2
6 9 2 3 12 12 2
12 9 13 3 2 7 13 9 7 13 9 3 2
21 9 1 15 13 9 2 13 0 9 0 7 13 9 2 15 13 3 13 0 9 2
10 9 0 9 11 9 9 13 15 3 2
3 3 13 9
25 10 11 13 0 9 9 16 15 13 10 9 13 9 7 3 9 9 2 7 15 15 13 3 0 2
11 11 9 9 13 9 2 3 9 9 13 2
9 7 3 13 13 11 13 3 15 2
9 7 9 13 3 2 3 10 9 2
19 11 13 3 13 0 2 7 10 9 15 13 13 9 3 16 13 0 9 2
9 10 9 9 13 15 0 9 9 2
5 13 12 0 9 2
4 9 13 9 15
7 13 15 3 13 3 9 2
4 9 13 13 2
11 9 13 13 2 16 11 9 13 9 9 2
7 9 10 9 0 13 9 2
4 3 13 9 9
4 15 13 9 2
8 13 9 0 9 3 0 9 2
4 13 0 9 0
4 13 13 9 2
15 11 12 9 13 0 11 1 11 7 11 9 13 3 0 2
12 7 3 15 3 13 0 9 2 16 3 13 2
4 0 13 0 2
8 13 3 9 13 0 9 9 2
7 3 13 9 13 9 0 2
5 15 13 11 1 2
8 13 3 9 15 3 13 9 2
8 15 13 10 9 12 0 9 2
5 15 0 11 8 8
10 9 13 16 9 13 3 3 1 9 2
3 9 13 3
15 3 15 13 9 2 7 15 15 13 3 9 7 9 9 2
7 13 15 15 13 7 13 2
9 15 13 13 15 10 7 15 0 2
12 9 13 0 9 9 13 7 13 16 9 9 2
9 9 13 13 9 9 7 15 9 2
7 13 11 13 9 7 9 2
8 11 9 9 12 7 9 9 12
4 15 13 3 6
11 9 13 3 9 1 13 0 2 0 9 2
14 15 13 13 11 7 13 10 9 9 12 7 13 3 2
2 0 9
6 11 9 13 0 9 2
14 3 10 3 13 9 13 3 9 2 13 9 13 9 2
7 15 7 15 13 3 9 2
7 13 12 9 9 7 9 2
10 0 9 13 9 9 3 9 13 3 2
7 10 12 11 9 13 9 2
5 11 13 9 9 2
6 9 1 9 13 0 2
6 11 13 9 3 9 2
8 3 15 13 0 0 2 11 13
5 13 3 3 0 2
4 9 13 13 2
4 11 13 11 2
8 13 9 9 2 13 15 3 2
13 13 15 3 2 3 16 15 13 10 9 1 9 2
2 13 13
5 13 9 13 9 2
7 3 10 0 9 13 13 2
9 9 13 0 9 2 15 9 13 2
6 11 13 13 3 11 2
6 3 13 9 13 15 2
18 13 13 9 2 16 9 13 0 9 7 9 2 15 15 3 9 13 2
6 0 9 13 3 3 2
9 15 13 13 3 13 0 9 9 2
12 11 9 13 13 9 13 9 3 3 0 9 2
13 12 9 3 11 13 13 3 11 12 9 0 9 2
17 9 13 3 15 2 16 10 12 9 13 9 1 13 10 9 9 2
12 11 13 11 3 12 2 3 15 13 3 0 2
3 9 0 9
10 0 12 9 13 13 12 9 12 9 2
3 9 13 9
3 15 13 11
13 9 1 11 13 13 7 13 9 3 9 7 9 2
8 9 13 13 13 9 9 13 2
11 13 0 2 16 9 0 9 13 13 0 2
15 11 11 13 3 9 11 2 15 13 9 9 7 9 1 2
12 12 9 13 15 15 2 7 15 3 13 15 2
15 13 2 16 3 3 3 15 13 10 0 9 7 0 9 2
7 11 13 13 9 9 9 2
12 7 13 13 3 2 15 13 10 9 3 9 2
12 13 13 12 12 9 3 16 9 9 13 13 2
6 11 13 11 9 9 2
8 9 13 0 2 13 9 9 2
11 15 13 0 13 16 10 9 10 9 13 2
11 9 13 13 2 16 13 10 9 13 9 2
13 3 13 13 2 16 10 9 9 13 13 1 9 2
10 15 13 9 3 9 2 0 15 13 2
11 2 11 13 3 15 13 13 9 3 15 2
10 9 13 13 2 7 9 9 13 13 2
7 9 9 13 9 0 9 2
3 13 7 13
14 9 13 9 2 16 9 13 9 9 11 0 11 9 2
8 10 9 16 13 15 13 9 2
5 13 13 3 9 2
2 13 13
2 12 9
11 9 13 9 2 15 13 13 9 0 9 2
9 15 13 13 15 1 16 15 13 15
4 9 13 9 9
11 13 15 13 2 3 13 13 10 0 9 2
9 11 13 0 2 16 9 13 9 2
28 3 10 9 9 13 13 0 9 16 16 3 3 11 13 10 0 9 7 15 3 13 0 3 8 0 0 9 2
7 2 15 13 3 13 15 2
8 9 13 9 13 0 12 0 2
12 13 15 13 2 16 11 13 3 9 9 1 2
14 16 3 13 13 16 15 13 3 9 7 10 10 0 2
3 9 13 0
4 13 15 0 2
5 10 0 9 13 6
5 15 13 0 9 2
27 15 2 15 9 13 3 13 2 13 13 2 16 3 15 3 13 2 16 3 13 9 13 13 15 0 9 2
23 2 3 13 13 11 9 2 2 11 13 3 2 2 16 13 9 2 15 3 13 13 2 2
11 13 9 13 9 13 9 9 9 13 9 2
19 3 9 3 10 9 10 9 13 9 11 3 3 0 9 2 12 13 9 2
16 10 9 13 13 9 2 16 3 9 13 13 9 2 11 13 2
10 13 3 9 9 2 16 13 13 3 2
2 9 9
10 15 15 13 15 13 16 15 13 15 2
8 9 9 3 9 13 0 9 2
4 15 13 13 2
6 0 11 2 11 7 11
6 9 13 9 13 3 9
12 11 9 13 9 13 13 9 2 7 13 9 2
2 13 9
10 7 10 9 13 9 7 9 0 9 2
3 10 0 9
6 15 9 13 9 9 2
5 13 3 13 9 2
8 12 0 9 13 13 9 9 2
6 9 13 13 0 9 2
31 16 3 10 0 3 0 0 9 13 3 3 3 7 3 10 9 15 13 3 15 13 3 15 13 16 15 13 3 3 3 2
12 3 3 13 13 3 13 2 3 10 0 9 2
10 0 9 15 3 13 13 2 13 11 2
10 9 9 13 11 2 11 7 9 9 2
4 15 13 0 2
5 15 13 13 0 9
8 15 3 13 2 16 15 13 2
3 15 13 15
12 6 2 3 3 15 9 13 3 3 9 1 2
8 9 13 11 13 3 12 9 2
18 13 9 13 2 16 15 13 9 9 2 7 13 13 13 2 16 13 2
11 16 10 9 13 13 2 13 15 3 3 2
3 13 9 2
7 9 7 11 13 13 0 2
9 13 9 9 0 9 9 13 9 2
7 15 13 13 3 0 9 2
9 9 13 9 2 9 2 7 11 2
13 11 13 13 10 0 9 2 7 3 15 3 13 2
5 10 9 1 13 2
2 13 9
8 9 9 13 11 3 0 9 2
16 16 9 9 13 3 13 2 9 9 2 12 9 2 13 9 2
1 13
9 11 9 13 9 0 9 11 11 2
15 11 13 15 2 16 11 9 13 0 9 9 9 0 9 2
4 13 12 1 2
6 13 9 7 9 12 2
12 13 15 13 2 15 13 12 9 3 9 9 2
6 9 13 3 12 9 2
6 9 13 13 13 9 2
24 15 1 13 13 0 9 10 9 2 13 3 0 9 2 13 9 7 9 2 13 16 0 9 2
8 11 9 9 13 3 3 13 2
5 15 13 3 13 2
7 3 15 13 13 9 9 2
4 0 9 11 11
7 9 13 3 9 3 9 2
2 13 13
14 3 11 7 11 9 2 10 12 9 2 13 9 9 2
15 9 13 3 9 9 15 13 15 15 0 2 13 15 3 2
13 9 9 13 15 2 16 0 13 9 9 13 9 2
3 9 1 13
6 15 13 13 11 9 2
2 9 9
13 11 7 11 11 13 13 15 13 15 3 13 7 9
8 11 0 9 13 13 13 13 2
3 13 15 0
7 15 13 13 0 0 9 2
6 3 9 13 0 3 2
6 13 15 13 3 3 2
17 9 11 11 13 10 9 2 16 9 13 7 13 13 9 13 3 2
7 3 3 13 13 10 9 2
2 13 13
12 6 3 2 16 3 13 2 13 11 0 9 2
5 0 13 9 1 2
12 9 0 9 13 3 9 0 7 3 0 9 2
3 13 9 2
7 13 9 3 7 13 9 2
11 13 15 3 3 13 3 15 3 13 3 2
3 0 9 13
8 11 13 0 9 0 9 9 2
4 9 13 0 2
10 13 9 7 3 13 9 7 13 9 2
4 15 15 13 2
5 15 13 13 9 2
7 9 1 13 13 2 16 2
2 9 13
6 13 2 3 13 9 13
5 9 13 13 0 2
7 3 15 13 9 2 3 2
4 15 13 3 0
5 15 13 13 9 2
8 13 3 3 13 0 9 9 2
7 10 0 9 13 13 0 2
7 15 13 3 15 13 9 2
5 9 13 9 13 2
4 11 9 0 9
4 13 13 3 2
14 9 13 11 9 13 2 7 15 13 13 9 3 9 2
7 9 13 9 1 9 12 2
4 13 13 3 2
14 3 13 0 9 9 2 16 3 15 13 0 9 9 2
15 15 13 13 3 12 9 9 1 2 15 13 13 13 3 2
5 9 13 3 13 2
5 15 13 3 13 2
6 9 9 9 13 9 2
6 9 13 9 9 0 2
24 15 13 3 15 13 13 15 3 3 15 3 15 13 0 9 3 15 13 13 15 3 0 3 2
2 0 11
2 9 3
19 12 9 9 9 9 9 13 3 13 13 9 2 16 15 13 13 9 9 2
2 0 9
9 11 13 9 9 2 16 13 15 2
8 13 9 2 15 3 13 9 2
4 13 9 1 2
14 9 9 13 9 1 13 11 9 12 9 11 9 1 2
7 0 13 13 15 11 9 2
16 9 7 0 9 13 9 3 9 9 2 0 9 9 7 9 2
4 15 13 13 2
6 13 13 13 10 9 2
6 3 13 10 0 9 2
6 13 3 15 3 13 2
13 11 9 9 11 11 1 9 13 9 13 0 9 2
5 13 3 9 0 2
16 9 13 13 11 2 11 2 11 2 11 2 11 7 11 9 2
2 0 9
11 2 9 2 2 15 13 9 9 9 9 2
13 11 13 3 0 13 9 2 9 3 12 12 9 2
17 9 13 3 9 9 2 9 7 9 2 13 3 10 10 9 13 2
21 11 13 10 9 7 13 13 10 9 2 15 1 0 7 0 9 13 9 0 9 2
10 15 13 15 13 13 9 9 9 9 2
6 3 13 9 1 9 2
5 13 15 10 9 2
8 13 3 13 15 2 11 13 2
5 9 13 15 9 2
6 9 9 13 0 9 1
3 13 0 9
8 3 13 7 13 10 9 9 2
2 10 9
8 9 13 13 0 9 9 1 2
7 10 9 13 3 9 13 2
5 13 9 13 9 2
4 6 15 13 0
7 12 9 13 13 0 9 2
5 6 16 13 0 2
4 9 13 15 2
5 9 13 9 0 2
5 15 13 9 13 2
5 15 13 13 9 2
4 9 0 9 2
11 3 13 13 13 9 11 2 13 0 9 2
4 6 13 13 2
5 9 13 1 9 2
16 9 9 13 3 9 2 16 9 13 13 12 9 9 9 13 2
19 13 3 13 9 9 7 13 0 9 2 16 12 9 13 3 11 9 1 2
12 11 9 11 2 9 11 2 13 0 9 13 2
3 13 0 9
8 0 9 2 15 13 13 11 2
9 13 15 13 9 2 16 13 3 2
5 15 13 0 9 2
10 11 13 13 2 16 13 13 13 9 2
9 0 10 9 13 13 13 9 1 2
11 13 13 13 13 9 0 2 16 15 13 2
5 11 13 13 12 2
2 15 1
8 9 9 7 9 9 13 9 2
6 12 9 13 9 9 2
13 9 9 13 13 9 2 7 15 13 9 10 9 2
5 6 2 10 9 2
5 9 13 9 13 2
8 3 3 13 9 3 7 13 2
11 9 9 13 16 15 3 13 13 10 3 2
6 15 13 0 13 13 3
7 9 13 3 0 16 9 2
5 15 15 13 3 13
5 13 3 13 9 2
2 13 13
13 15 13 13 13 2 16 2 15 13 3 3 2 2
6 10 9 13 13 9 2
4 10 12 0 9
11 10 9 13 9 2 15 13 3 0 9 2
3 11 13 9
6 9 13 12 12 9 2
6 15 13 13 13 13 2
10 15 13 3 3 13 10 11 11 2 9
13 9 13 12 9 13 9 2 7 3 13 0 9 2
5 9 15 13 9 2
13 9 1 11 13 1 11 2 7 13 13 15 9 2
11 3 0 9 13 11 7 11 9 11 1 2
7 0 9 9 13 9 9 2
16 3 9 13 9 16 13 0 9 2 16 10 0 15 3 13 2
9 13 9 1 2 1 7 15 1 2
4 15 13 9 2
2 9 9
11 3 16 10 9 13 3 13 3 3 3 2
8 11 13 9 1 0 9 1 2
19 3 13 13 13 15 2 13 15 2 13 9 13 9 2 13 9 13 9 2
4 3 13 3 2
18 0 9 15 13 10 9 13 2 7 13 3 3 15 13 0 9 13 2
17 9 13 13 11 2 3 15 13 13 2 2 3 11 13 13 2 2
10 11 9 13 9 13 9 3 1 9 2
7 11 13 13 7 13 9 2
8 9 9 13 12 9 9 9 2
16 11 13 9 12 9 3 2 7 13 15 3 3 3 9 13 2
3 3 15 1
3 9 13 9
3 10 9 2
16 9 13 9 3 3 2 16 9 13 0 9 7 9 13 3 2
6 13 3 0 10 9 2
18 3 15 13 2 15 15 13 2 15 13 7 13 16 15 13 13 3 2
6 9 13 9 1 9 2
6 9 11 11 13 9 2
3 3 9 2
12 3 2 15 13 9 0 2 7 3 7 3 2
3 11 13 15
8 3 9 13 3 10 9 3 2
3 3 9 2
2 13 3
12 3 13 3 10 0 9 2 13 15 7 13 2
3 13 3 2
5 11 13 9 3 2
6 9 1 9 13 0 2
12 15 13 3 7 9 13 3 9 1 9 1 2
3 12 0 9
9 9 9 13 3 13 10 9 9 2
5 11 13 3 9 2
9 13 7 13 7 3 13 13 9 2
3 3 13 9
7 9 7 9 13 13 11 2
10 3 13 12 0 9 2 15 13 9 2
4 10 13 9 9
4 3 9 13 2
4 9 9 12 2
9 3 15 13 3 0 16 15 13 2
9 3 3 13 3 0 9 10 9 2
10 13 3 13 9 2 16 9 13 3 2
6 15 15 3 3 13 2
4 15 13 9 2
29 13 16 3 15 13 9 9 9 7 3 15 3 15 13 3 12 7 3 13 10 9 3 13 3 13 13 3 3 2
11 15 13 10 9 2 3 0 9 7 9 2
4 13 13 9 2
4 11 15 13 2
10 15 13 13 2 13 15 15 7 13 2
4 0 0 9 2
10 11 13 3 2 10 15 3 9 2 2
10 9 10 9 13 0 9 13 9 9 2
6 11 12 9 13 9 2
5 9 13 9 1 2
6 15 15 13 13 3 2
7 9 13 16 13 9 3 2
8 15 9 9 13 10 0 9 2
10 2 15 13 3 13 9 2 13 15 2
8 13 3 13 13 9 3 3 2
8 11 13 13 2 7 15 13 13
4 15 13 0 13
4 3 15 13 2
5 9 9 13 0 2
5 9 11 13 12 2
8 0 9 15 13 2 15 3 13
5 9 7 9 13 2
15 11 13 13 13 3 12 9 1 2 7 9 13 9 13 2
8 11 12 9 13 0 9 9 2
7 11 9 13 15 16 11 2
3 13 9 0
7 9 7 9 13 3 13 2
13 13 15 9 9 2 7 3 9 7 9 13 9 2
10 15 13 7 13 2 16 9 13 13 2
5 15 13 13 9 2
9 13 0 2 16 3 0 13 0 2
3 9 13 13
10 15 13 16 13 9 3 15 13 13 2
5 15 13 11 9 2
11 0 9 13 9 2 0 7 3 9 9 2
15 11 9 13 3 0 2 16 3 7 3 13 13 9 9 2
4 11 13 12 2
11 13 10 9 0 3 3 2 13 10 9 2
5 15 13 1 9 2
10 13 13 13 2 16 0 9 13 3 2
9 13 13 3 3 16 15 13 9 2
15 13 13 9 2 15 13 0 9 7 13 11 13 9 3 2
14 15 13 3 13 13 2 16 13 13 9 9 11 9 2
10 15 13 13 13 15 10 11 3 7 2
8 15 13 13 3 3 12 9 2
7 9 2 9 2 10 9 2
13 12 9 9 7 0 9 13 13 11 13 9 11 2
10 15 13 2 16 15 13 13 0 9 2
9 9 13 11 13 11 11 12 9 2
13 13 13 9 3 0 2 16 9 13 3 3 0 2
3 9 13 13
12 11 9 9 13 13 2 16 15 13 3 9 2
9 13 2 16 13 13 3 3 13 2
5 9 13 11 11 9
2 0 9
15 10 9 13 13 13 0 2 7 9 7 1 10 9 13 2
15 16 13 11 9 2 15 13 3 3 2 13 9 9 11 2
4 15 13 13 2
11 15 13 2 16 0 9 13 1 10 9 2
4 3 3 9 2
5 9 13 9 13 2
2 11 9
7 13 9 13 7 9 3 2
3 13 9 3
3 9 13 9
2 13 9
13 15 13 9 7 9 2 15 3 13 9 7 9 2
6 13 9 7 13 9 2
3 13 9 9
12 11 13 2 16 9 3 13 13 9 7 9 2
8 13 15 13 9 15 13 3 2
7 9 11 13 13 9 1 2
18 3 10 11 3 13 13 10 9 16 15 3 3 13 10 9 10 9 2
4 15 15 13 0
2 12 9
2 15 1
3 13 13 2
8 9 13 3 0 13 0 9 2
7 13 0 9 3 10 9 2
7 15 13 11 16 9 13 2
11 0 9 13 3 2 16 9 9 13 9 2
11 16 15 0 13 2 13 9 3 10 9 2
9 9 13 3 13 9 2 13 9 2
6 15 13 3 0 9 2
12 9 13 3 0 2 16 3 13 9 13 15 2
4 3 13 9 2
3 8 7 9
5 15 13 0 9 2
8 15 13 13 3 3 3 12 9
7 6 15 13 13 15 3 2
4 9 13 15 9
2 3 11
14 15 13 0 9 2 7 0 9 13 9 0 2 0 2
13 9 9 13 9 11 11 7 9 13 12 12 12 2
6 13 2 16 9 13 0
15 11 9 13 13 13 2 3 10 9 3 12 9 9 13 2
9 7 15 1 15 13 13 3 9 2
3 13 0 9
4 13 15 11 2
6 3 7 13 9 3 2
9 3 9 13 13 12 9 9 1 2
3 13 13 9
2 9 15
11 11 13 13 9 7 15 13 13 9 3 2
7 13 3 3 13 3 15 2
8 13 0 13 0 7 13 15 2
10 13 3 15 2 16 9 13 3 13 2
5 9 13 3 0 2
2 11 9
4 9 12 10 9
7 3 3 13 13 3 0 2
2 0 9
2 11 9
6 9 13 9 3 3 2
9 0 9 15 13 13 12 9 11 2
7 9 9 13 1 10 9 2
5 13 0 13 9 2
5 9 13 9 9 2
13 0 12 7 3 12 9 1 9 13 13 11 0 2
4 13 13 15 2
4 2 13 9 2
3 13 9 9
4 9 7 10 13
6 13 3 3 12 9 2
9 15 13 10 9 13 13 0 9 2
3 9 13 13
5 15 13 9 0 3
6 13 13 9 0 11 9
5 6 16 13 0 2
9 13 3 9 3 7 3 0 9 2
11 9 7 9 2 9 12 9 2 0 9 2
12 15 3 15 13 15 9 2 16 13 0 9 2
2 10 9
4 13 0 16 13
10 9 13 13 0 9 3 0 9 1 2
3 9 13 3
3 15 13 3
5 13 13 9 0 9
12 11 13 13 3 9 2 7 13 10 0 9 2
4 9 3 13 9
8 13 0 3 2 16 3 13 2
3 13 13 13
17 16 15 13 3 3 15 1 13 3 2 13 9 7 13 9 3 2
4 15 13 13 11
5 9 13 15 13 9
4 9 13 9 2
11 10 9 13 3 2 16 13 3 3 9 2
6 9 13 9 13 9 2
15 13 2 16 3 13 13 10 9 2 13 3 9 7 13 2
7 9 13 0 9 3 13 2
4 13 15 13 2
4 0 9 0 9
3 13 0 13
7 13 3 16 15 13 9 2
25 1 15 2 13 11 9 9 7 9 2 1 9 11 0 9 13 0 9 2 11 9 13 0 0 2
11 9 11 11 13 13 3 13 3 13 9 2
10 15 7 10 9 13 10 0 0 9 2
1 12
5 9 13 7 13 3
12 11 11 2 3 11 2 13 11 12 9 12 2
4 11 13 13 2
12 13 3 0 13 9 7 3 13 9 13 13 2
8 3 9 13 7 13 0 9 2
3 13 3 2
6 15 13 0 15 15 13
7 10 15 13 15 13 9 2
16 16 13 15 13 0 13 2 3 9 1 13 13 9 7 9 2
15 11 7 0 15 13 13 15 3 2 16 15 13 13 9 2
3 13 9 2
4 2 13 13 2
4 9 13 0 2
12 10 9 13 3 12 9 2 10 9 13 13 2
5 15 13 3 9 2
8 9 1 3 9 13 3 11 2
10 3 13 3 0 13 15 0 9 1 2
4 15 13 9 2
9 3 13 9 7 15 13 3 0 2
8 7 15 13 2 15 13 13 2
4 15 13 9 2
17 10 10 3 9 16 13 16 15 3 3 15 13 3 16 13 15 13
21 9 13 3 2 16 9 13 9 9 2 7 13 15 13 2 16 9 13 3 3 2
15 3 0 9 7 0 9 1 13 13 13 9 9 12 9 2
7 7 15 13 3 9 0 2
9 11 13 9 2 16 9 13 13 2
4 13 0 13 9
19 9 1 9 3 13 13 9 0 9 13 15 2 13 9 11 11 3 11 2
7 11 13 13 12 9 13 2
6 13 3 15 0 13 2
6 3 13 9 13 9 2
5 9 13 3 12 2
9 9 13 3 2 16 13 13 9 2
14 3 15 13 10 10 9 7 13 16 13 15 9 9 7
9 9 15 13 2 15 9 9 13 2
20 10 9 13 9 3 3 13 9 2 16 13 9 15 13 10 0 9 2 7 2
4 11 13 9 2
15 15 13 3 13 16 15 13 3 13 2 3 13 3 13 2
13 13 9 15 13 11 9 13 9 2 0 11 2 2
2 13 13
4 15 13 9 11
4 3 9 13 2
8 11 13 0 9 9 1 7 13
4 9 9 13 2
7 10 9 13 3 9 9 2
9 9 9 3 12 9 7 12 9 2
8 13 3 2 16 15 13 13 2
18 11 9 13 2 16 9 13 13 3 12 9 9 2 15 13 3 0 2
5 9 13 0 9 2
6 3 10 3 13 9 2
5 11 15 13 7 2
7 13 3 16 9 13 13 2
10 9 13 12 1 9 2 9 12 9 2
4 13 3 9 2
6 13 3 16 0 9 2
4 9 13 9 2
6 3 13 9 0 9 2
10 9 13 13 9 9 7 3 13 0 2
4 11 13 9 2
7 9 16 13 3 13 9 2
5 9 9 9 11 11
4 9 13 3 9
6 3 13 3 3 0 2
8 10 0 13 0 0 9 9 2
3 9 13 9
2 9 9
5 9 13 3 9 2
5 15 13 0 9 2
8 11 13 9 9 13 9 1 2
8 9 13 13 2 7 13 13 2
5 11 13 3 0 2
4 9 13 3 2
4 13 15 3 13
8 9 0 9 3 12 9 9 2
13 10 9 13 3 13 2 16 15 13 9 0 9 2
7 9 13 3 3 10 9 2
5 13 3 0 9 2
7 9 13 3 13 9 9 1
9 7 13 10 9 13 13 11 9 2
11 11 13 13 11 0 9 7 13 15 3 2
2 9 1
5 6 6 2 9 2
10 9 13 3 11 3 0 9 13 11 2
4 9 7 0 9
9 13 13 13 10 9 2 13 0 2
14 3 0 9 11 13 13 11 9 11 7 11 9 11 2
8 7 9 1 15 3 13 13 2
11 9 7 3 9 1 0 13 9 9 0 2
6 3 15 3 3 13 2
10 15 15 3 3 13 2 0 0 9 2
9 11 13 9 2 7 9 13 9 2
4 0 9 9 3
9 15 13 0 9 9 7 9 0 2
8 0 9 13 9 0 9 1 2
5 15 13 12 12 2
3 9 13 9
10 11 13 11 9 7 13 3 0 9 2
6 3 0 9 13 3 2
24 13 11 11 11 12 9 2 9 9 2 2 2 15 13 3 3 0 9 2 9 7 9 2 2
10 9 13 3 9 7 15 13 9 0 9
16 10 9 15 13 2 15 13 9 9 9 7 9 9 9 9 2
9 9 13 2 13 3 3 0 9 2
7 9 13 0 12 9 9 2
4 3 15 13 2
7 13 13 2 15 13 9 2
8 9 9 13 13 9 1 0 9
6 9 13 10 9 3 2
6 13 3 9 13 9 2
3 13 13 3
7 9 13 9 15 13 9 2
6 15 13 3 3 0 2
6 13 9 0 0 9 2
2 15 15
4 9 9 0 9
10 15 13 0 7 3 3 0 7 0 2
12 7 12 9 13 7 13 9 9 12 7 12 2
17 7 15 13 16 15 15 3 13 0 9 7 0 7 9 13 7 2
4 13 9 3 2
3 13 3 13
15 0 0 9 13 15 2 16 9 9 13 9 3 0 9 2
4 11 13 11 2
6 15 3 3 13 15 2
16 11 13 3 3 9 9 3 16 13 13 2 16 9 13 13 2
2 13 9
6 13 13 3 13 9 2
5 9 13 9 9 2
4 0 10 9 2
14 9 13 9 0 9 0 9 7 9 0 9 9 1 2
8 10 9 9 13 9 13 9 2
5 9 13 12 1 12
12 9 9 13 2 16 9 13 13 3 13 9 2
19 3 3 9 9 2 15 3 13 13 13 11 9 9 2 13 11 9 3 2
6 3 3 15 13 13 2
9 13 11 0 9 7 11 0 9 2
11 15 1 11 3 13 3 10 9 9 9 2
7 13 2 16 13 10 0 2
12 15 3 13 13 10 9 3 10 9 1 9 2
9 3 3 13 12 9 13 11 9 2
11 7 13 13 3 2 16 9 13 13 9 2
4 13 9 13 2
22 3 12 13 9 13 13 0 0 9 2 16 0 9 9 7 9 9 13 13 0 9 2
8 13 15 0 16 15 13 13 2
7 11 13 0 9 3 0 2
4 13 15 9 2
8 3 15 13 3 3 0 9 2
4 15 15 13 2
7 3 15 13 2 13 9 2
13 15 13 9 1 13 3 9 9 0 9 0 9 2
8 13 13 9 9 9 3 3 2
11 3 9 13 3 3 2 15 15 3 13 2
6 9 9 13 13 9 2
9 9 13 13 3 13 13 3 9 2
3 15 13 9
8 9 0 13 0 15 0 9 2
12 3 15 7 13 9 7 15 13 7 13 9 2
5 9 13 13 0 2
5 15 13 15 15 2
10 7 16 9 13 3 2 15 13 3 2
12 11 9 7 9 9 13 15 13 3 12 9 3
13 11 11 9 7 11 9 2 13 13 9 12 1 2
2 11 9
4 13 0 3 2
2 13 9
5 9 13 12 3 12
21 0 9 13 10 3 0 9 2 16 15 13 13 13 7 0 7 0 2 3 15 2
4 13 15 13 2
10 15 13 2 13 13 13 3 9 9 2
9 16 15 13 15 2 13 13 0 2
5 9 13 0 3 2
8 9 9 16 13 2 6 9 2
2 13 11
21 16 13 13 2 13 13 10 9 9 12 9 1 9 9 2 7 9 0 9 9 2
9 13 13 10 9 7 3 15 13 2
4 9 10 9 2
6 13 13 13 0 9 2
6 3 12 9 13 13 2
11 9 9 9 13 3 9 2 9 7 9 2
11 16 0 13 2 0 9 13 13 0 9 2
7 9 13 9 0 7 0 2
4 9 13 13 2
8 11 13 15 13 15 9 9 2
5 15 15 3 13 2
16 3 0 13 2 16 11 2 15 13 13 9 2 13 9 13 2
2 10 9
17 11 13 2 16 13 9 9 3 7 13 15 15 1 13 0 9 2
2 13 9
10 3 11 13 13 10 9 9 2 7 2
18 9 13 13 9 15 1 2 16 3 13 13 3 13 3 0 13 0 2
10 2 15 13 13 13 3 15 16 9 2
8 15 13 3 13 3 9 1 2
9 13 10 15 13 0 9 16 15 2
4 15 13 3 9
3 13 15 13
8 13 3 2 9 13 3 3 2
3 13 13 2
5 0 9 10 9 2
13 9 13 0 2 9 3 0 16 15 3 13 9 2
10 9 11 13 9 2 9 9 1 2 2
6 15 9 10 9 13 2
11 9 13 3 3 3 9 1 15 2 16 2
16 16 13 9 9 7 9 1 9 3 13 9 13 13 9 9 2
18 15 3 13 11 9 3 10 9 7 7 3 10 9 3 13 13 9 2
13 11 0 8 8 8 13 9 7 3 3 13 13 2
2 13 9
13 9 11 13 9 9 9 9 2 3 9 9 13 2
9 16 9 13 11 2 11 9 13 2
4 13 0 2 16
8 7 9 1 13 9 7 9 2
2 3 13
8 10 9 11 11 13 9 9 2
57 7 3 10 9 0 9 13 13 15 16 10 9 13 13 13 13 10 9 15 15 13 2 7 10 9 13 13 9 2 7 3 16 3 3 13 3 10 9 13 10 9 1 15 16 10 9 13 9 2 15 13 3 0 9 9 1 2
6 3 13 9 3 13 2
4 15 3 13 9
17 16 15 13 3 9 0 9 2 15 13 3 13 3 0 2 0 2
12 9 13 9 9 7 1 0 9 13 9 0 2
13 16 9 13 9 11 2 13 15 3 13 13 11 2
14 0 9 11 13 9 9 1 13 0 9 2 9 9 2
4 11 13 9 2
12 3 11 13 10 0 9 9 2 16 13 9 2
2 7 3
5 13 3 13 3 2
11 13 3 3 9 2 15 10 9 13 13 2
3 2 3 2
2 0 9
7 9 13 13 0 9 9 2
5 3 13 3 9 2
11 13 9 13 3 0 9 13 9 0 9 2
6 2 13 13 16 13 2
10 11 9 13 9 13 3 13 13 13 2
8 13 2 16 15 13 3 9 2
7 15 13 3 15 15 13 2
10 3 11 13 2 16 10 9 13 3 2
8 13 3 9 13 3 13 9 2
16 7 15 13 13 15 3 16 15 3 13 3 16 15 13 3 13
10 3 13 3 9 9 13 9 0 9 2
9 9 2 15 9 13 13 3 9 2
12 9 13 9 13 9 12 9 9 9 12 1 2
2 3 3
7 9 13 12 9 9 3 2
4 15 3 9 2
7 15 13 13 9 3 9 1
9 13 13 16 13 15 13 0 9 2
24 9 2 10 9 0 9 3 9 0 9 2 3 9 13 0 1 13 3 3 7 13 9 9 2
10 8 8 9 9 13 3 0 9 9 2
7 15 13 0 9 9 12 2
5 13 3 3 3 2
6 3 11 13 13 9 2
12 16 9 3 13 9 2 9 13 13 12 9 2
7 15 13 3 12 9 9 2
14 2 13 3 15 3 3 13 2 7 13 3 13 15 2
8 9 1 9 13 9 12 9 2
13 9 9 13 9 9 3 2 9 9 7 9 9 2
7 12 0 9 13 3 9 2
12 9 13 9 13 0 13 2 16 9 9 13 2
2 13 9
3 13 9 2
4 13 13 3 2
11 15 16 13 11 1 9 13 7 13 3 2
6 9 13 0 9 9 2
4 13 3 13 2
2 13 9
5 15 13 9 3 2
12 3 15 3 13 3 2 16 13 13 15 0 2
16 15 13 3 16 10 9 13 3 13 3 16 15 3 13 9 2
4 0 16 9 1
6 10 9 13 3 11 2
2 13 13
9 3 16 9 13 2 9 13 9 2
6 13 0 0 7 0 2
8 13 13 15 2 15 13 13 2
2 9 1
6 9 11 7 9 11 2
7 9 9 13 9 12 9 2
5 9 13 11 13 11
8 15 13 3 3 13 9 3 2
4 0 3 13 2
2 0 3
3 13 15 1
8 9 7 9 13 0 1 9 2
3 0 9 9
17 10 9 9 13 9 2 12 0 9 2 15 13 13 13 9 9 2
9 13 15 13 16 15 2 3 12 2
2 16 13
9 9 13 9 0 7 3 15 13 2
20 11 9 1 11 13 13 13 13 9 2 7 9 2 15 11 13 13 3 3 2
23 11 13 3 3 3 0 9 2 16 3 13 10 9 13 9 2 15 13 3 0 7 0 2
11 11 11 13 0 11 9 11 0 9 1 2
13 11 13 16 9 13 3 3 3 16 15 13 13 2
4 0 13 11 2
12 9 13 3 0 9 2 16 15 13 15 0 2
4 9 13 13 2
2 0 3
6 3 13 3 10 15 2
8 13 13 13 15 9 0 9 2
12 0 9 1 9 13 11 7 11 11 0 9 2
8 13 15 13 11 1 13 9 2
9 13 12 9 9 7 13 15 9 2
7 9 3 13 2 15 15 13
12 11 13 2 13 9 7 13 9 10 9 2 2
13 9 13 7 3 11 9 3 3 13 7 3 3 2
4 3 3 13 2
6 9 9 13 0 13 2
3 13 9 9
10 0 9 9 13 3 13 12 0 9 2
6 3 15 13 15 13 2
8 9 13 3 0 9 16 9 2
4 3 9 9 3
16 11 11 13 13 13 3 10 9 3 13 16 11 9 9 1 2
7 13 3 13 9 2 7 2
5 13 15 3 0 2
13 7 3 3 15 13 15 13 16 15 13 3 3 2
4 3 13 3 2
4 11 13 13 13
6 15 13 3 13 3 2
9 13 3 13 10 9 3 7 15 2
7 13 9 3 7 13 9 2
13 16 9 13 9 13 3 13 2 13 9 0 9 2
4 15 13 9 15
20 13 9 3 0 2 16 15 9 1 13 13 9 9 9 2 9 9 7 9 2
10 7 2 6 2 15 13 0 9 15 2
8 9 13 3 3 0 9 9 2
9 15 13 13 9 2 13 13 9 2
8 13 2 0 13 13 0 9 2
11 13 13 15 2 15 13 7 13 9 9 2
10 13 13 3 0 9 2 13 2 0 2
11 0 9 9 13 9 7 7 9 7 9 2
6 11 13 13 0 9 2
18 15 13 3 3 16 15 13 10 9 16 10 15 15 13 3 13 16 2
8 9 13 0 7 0 10 9 2
13 9 13 2 16 13 9 9 13 10 9 16 9 2
4 9 13 3 2
4 3 9 13 2
2 10 9
7 3 13 16 12 9 9 2
2 9 2
3 9 13 9
3 10 0 9
3 13 9 2
2 13 13
11 9 13 12 9 2 9 13 3 13 3 2
14 3 15 13 2 16 0 9 2 0 9 13 9 9 2
7 15 13 2 3 15 9 13
9 9 13 0 2 16 3 13 13 2
12 9 13 13 9 9 1 9 2 7 3 9 2
2 6 6
5 15 13 9 13 9
6 11 13 13 9 9 2
15 9 13 0 9 2 16 13 12 9 2 3 13 15 3 2
3 12 9 0
2 6 2
19 11 13 13 0 12 9 1 7 13 3 13 0 9 2 15 13 13 9 2
9 3 15 13 13 3 3 16 11 2
6 9 13 13 0 11 2
5 15 13 9 9 2
16 11 13 0 0 9 2 16 3 13 3 13 13 9 9 9 2
6 11 13 11 0 9 2
11 0 9 1 9 13 13 13 9 3 13 2
9 9 9 13 13 3 1 9 9 2
4 15 13 10 9
12 11 1 9 13 13 13 2 13 3 10 9 2
10 15 13 3 10 9 15 13 3 3 9
5 13 10 11 9 2
23 3 15 13 3 0 13 16 13 15 15 13 13 15 13 13 3 3 16 13 13 0 9 2
13 3 10 9 13 13 3 7 3 15 13 13 9 2
5 15 13 15 9 2
2 3 13
10 0 11 11 13 13 0 9 0 9 2
7 9 13 13 12 9 1 2
3 13 3 11
14 13 13 10 9 2 16 9 10 9 9 9 3 13 2
6 9 9 15 13 9 2
16 0 9 2 16 15 13 15 2 16 13 7 13 7 13 15 2
17 10 0 9 13 9 1 13 13 9 9 2 15 3 13 9 9 2
5 9 15 13 0 2
6 9 2 15 13 13 9
2 13 13
9 13 13 9 2 11 13 1 9 2
18 9 9 7 3 3 13 9 1 11 13 3 9 7 9 7 3 9 2
7 13 13 9 7 9 7 9
14 13 13 2 16 15 13 10 0 9 0 12 9 1 2
10 9 13 3 0 9 13 10 9 9 2
13 15 11 9 13 3 0 7 10 9 13 9 0 2
2 0 9
2 0 13
6 15 13 11 7 11 2
8 11 13 9 9 11 9 9 2
15 0 9 13 0 7 0 13 2 7 10 9 13 9 9 9
22 15 13 13 2 15 15 13 15 15 13 13 2 7 3 13 11 13 16 15 13 15 2
8 10 9 15 13 12 9 15 2
5 15 15 13 15 2
7 15 16 15 13 0 9 2
5 9 13 9 13 2
16 3 2 16 13 9 2 15 13 13 3 9 9 0 9 1 2
6 15 13 13 7 13 2
2 9 9
10 15 13 9 9 13 7 13 13 9 2
11 9 11 7 11 11 13 0 13 9 3 2
9 10 12 13 13 13 9 3 9 2
9 15 13 0 9 2 15 13 0 2
4 13 3 9 2
14 0 3 13 0 9 0 9 2 13 15 13 9 3 2
5 15 13 3 3 2
7 3 15 13 13 9 15 2
4 9 13 9 2
4 15 13 13 11
4 11 13 9 0
26 9 13 15 1 0 9 2 3 0 7 0 2 0 7 0 16 13 15 0 9 13 0 9 0 9 2
12 13 0 2 16 9 13 2 9 13 3 3 2
5 15 13 0 9 2
6 9 13 2 9 13 2
5 11 13 13 9 2
6 13 9 13 15 3 2
8 15 13 9 9 7 13 9 2
9 16 9 13 9 2 11 13 9 2
3 13 15 1
12 3 9 13 9 2 16 11 13 13 0 9 2
14 16 11 13 9 2 9 2 2 13 11 15 10 9 2
8 3 15 13 10 0 0 9 2
19 0 9 13 10 11 9 13 9 2 7 0 0 9 15 13 9 13 13 2
3 13 13 2
6 0 13 11 13 9 2
3 13 11 2
7 9 2 3 0 9 15 2
7 0 9 13 3 3 3 2
5 15 1 13 9 2
4 9 3 3 2
10 3 12 9 1 13 9 3 13 9 2
6 9 13 3 0 9 2
17 3 9 13 9 2 0 9 2 7 9 9 13 0 9 0 9 2
18 9 2 16 9 13 3 3 3 9 9 9 2 16 9 9 3 13 2
7 0 9 9 13 3 9 2
6 9 13 3 0 0 2
7 13 9 7 9 10 9 2
21 11 13 13 2 16 11 1 13 13 9 2 2 15 9 0 9 13 13 13 2 2
5 9 13 9 13 2
6 9 13 16 13 13 2
12 15 13 9 9 2 9 2 9 7 10 15 2
3 13 3 15
9 11 13 11 9 9 0 7 0 2
5 11 13 11 1 2
9 10 9 13 9 1 9 9 3 2
10 3 9 13 3 3 16 9 9 0 9
11 9 13 13 0 3 9 7 3 0 15 2
10 9 13 9 13 0 9 9 9 9 2
8 10 9 16 15 13 13 9 2
2 12 9
9 15 13 9 2 3 0 7 3 0
5 9 13 1 9 2
2 15 13
2 13 13
5 15 13 15 3 2
32 3 15 13 15 13 10 9 9 0 16 16 15 13 13 15 9 3 15 13 3 13 3 9 3 3 3 16 9 13 16 9 9
13 9 9 13 9 9 2 15 13 9 1 13 9 2
4 9 13 13 2
6 9 13 13 13 0 2
10 13 11 2 15 15 13 9 9 9 0
10 13 13 15 3 3 13 10 9 9 2
12 3 0 2 15 13 16 9 13 3 9 13 2
4 9 13 0 2
4 15 13 0 9
11 15 3 13 9 2 15 13 13 15 13 2
9 9 13 9 13 9 0 16 9 2
6 15 13 2 15 13 2
2 0 9
2 0 11
16 9 9 13 13 9 1 13 9 2 10 9 13 13 10 13 2
21 9 2 10 9 9 9 9 13 2 13 3 3 2 9 9 2 2 3 9 13 2
21 13 3 0 16 0 9 9 13 15 15 13 0 2 16 3 9 13 13 3 3 2
8 13 13 9 9 15 13 3 2
9 15 3 13 2 16 13 9 13 2
5 9 9 10 9 1
7 13 9 13 3 9 1 2
8 9 13 3 10 9 9 9 2
15 9 15 3 13 7 13 15 2 16 13 13 3 9 9 2
5 13 15 9 0 2
3 15 13 3
7 0 9 0 9 13 9 2
19 3 15 13 0 2 16 9 13 15 9 15 13 7 13 9 3 16 13 2
8 13 3 3 15 13 10 9 2
2 9 11
5 13 15 13 13 11
5 9 13 3 3 2
8 10 9 15 13 13 1 15 2
6 15 13 13 13 3 2
5 15 13 9 3 2
12 15 3 15 9 2 9 13 0 7 9 9 2
8 9 13 13 0 9 12 9 2
8 13 3 0 2 13 0 0 2
9 3 15 13 13 13 9 3 3 2
7 9 9 13 3 12 9 2
4 9 13 9 9
2 0 9
12 0 9 13 3 13 2 16 9 13 13 0 2
17 13 9 7 9 13 10 9 2 15 13 15 3 2 16 9 13 2
3 0 0 11
13 9 10 9 3 13 2 16 9 13 9 0 9 2
10 11 0 9 13 3 0 2 15 13 2
14 15 9 15 13 3 0 9 2 0 15 15 3 13 2
17 9 15 13 11 1 11 2 9 13 15 10 9 7 9 13 3 2
2 0 11
10 9 13 0 13 2 7 3 0 13 2
11 13 11 7 11 13 11 13 11 11 9 2
7 9 13 9 7 9 9 2
14 12 3 9 13 11 2 15 13 9 3 9 7 9 2
22 0 9 1 12 9 13 9 12 9 9 0 11 9 13 13 9 11 7 9 11 11 2
10 15 13 15 15 13 16 11 13 13 2
9 11 9 13 3 3 13 3 0 2
5 15 13 13 9 13
7 9 9 9 7 3 0 9
11 3 15 13 3 0 7 15 13 3 10 9
7 6 2 15 13 3 9 2
61 3 3 2 3 15 9 11 7 13 0 9 7 3 15 13 13 13 3 7 3 15 13 16 11 7 11 13 3 3 7 3 7 3 16 8 16 11 13 3 9 7 13 16 13 9 6 3 15 13 7 15 13 3 11 9 7 3 11 13 16 2
10 13 0 15 2 16 10 9 13 13 2
12 9 13 9 2 7 15 13 3 3 9 1 2
5 13 10 9 3 2
8 13 0 2 16 15 13 13 2
9 0 9 13 3 0 3 9 13 2
10 9 2 9 2 9 13 3 9 15 2
6 10 9 13 9 13 2
9 11 13 3 9 9 7 9 9 2
11 10 9 10 9 13 9 2 15 3 13 2
4 2 13 9 2
3 3 9 3
3 13 3 2
6 9 13 9 3 3 2
10 9 13 3 3 3 16 9 9 13 2
10 9 13 13 12 9 13 9 3 9 2
9 0 9 15 13 9 0 0 9 2
10 13 13 13 10 0 16 15 3 13 2
4 13 3 9 2
6 11 7 11 13 15 2
2 9 13
3 9 9 1
4 3 15 13 3
4 9 13 3 2
7 11 9 13 15 0 3 2
20 0 9 9 13 13 9 2 7 15 13 15 2 16 3 3 9 13 9 0 2
2 9 13
15 15 1 12 9 9 13 13 3 15 3 13 3 7 3 2
4 10 9 13 2
8 13 9 7 0 0 9 9 2
7 9 1 15 13 3 3 2
7 3 10 9 9 13 9 2
9 15 13 13 2 16 9 3 13 2
12 9 3 13 9 9 7 9 13 13 15 3 2
5 3 9 13 0 2
6 11 2 15 13 9 2
9 10 9 13 9 10 9 9 9 2
8 15 13 0 2 16 9 13 2
2 3 0
8 11 13 2 9 13 3 13 2
7 9 13 3 13 9 3 2
6 15 13 9 3 13 9
7 9 9 13 9 11 11 2
11 13 3 11 11 2 15 13 9 3 9 2
15 15 13 3 0 9 2 16 13 12 9 13 3 0 9 2
4 9 13 3 2
6 3 13 3 3 3 2
2 0 9
12 15 13 9 9 1 2 15 13 3 12 12 2
2 6 6
14 0 13 13 3 9 2 16 13 13 9 13 0 9 2
2 9 0
16 3 16 13 3 3 7 3 13 12 9 3 2 3 3 15 13
17 7 3 13 10 0 3 6 0 3 15 3 13 9 9 10 15 2
6 15 13 13 16 15 13
5 15 13 9 1 2
5 11 13 13 9 15
6 9 13 13 3 16 13
5 9 13 13 9 2
3 15 15 13
14 10 9 13 15 13 2 16 9 13 10 15 16 9 2
15 11 11 9 13 0 13 12 9 2 15 13 0 0 9 2
15 15 3 13 10 9 2 7 3 13 9 7 9 7 9 2
13 9 13 3 13 13 2 15 13 2 16 13 9 2
15 6 3 2 16 9 13 15 16 15 13 12 9 9 9 2
6 3 10 10 0 9 13
24 0 9 2 16 15 13 3 2 13 2 16 9 13 13 13 3 10 9 2 16 9 13 9 2
4 9 13 12 9
7 13 13 3 9 13 3 2
7 3 15 13 9 0 9 2
5 0 9 15 13 2
3 3 9 2
6 11 13 15 13 3 2
10 9 13 13 15 0 9 1 0 9 2
8 15 13 10 9 15 13 9 2
12 9 9 13 3 0 2 15 13 13 7 13 2
5 15 13 9 3 2
10 7 3 13 3 12 9 3 10 9 2
14 16 9 13 13 9 3 13 1 9 2 13 3 13 2
4 15 13 10 9
2 0 9
11 9 9 13 13 13 9 7 13 0 9 2
3 9 13 0
8 9 11 2 13 3 0 9 2
7 13 9 2 13 15 13 2
7 3 13 9 7 9 9 2
18 7 3 9 13 13 11 11 7 3 10 9 2 16 13 9 9 13 2
3 3 0 2
3 9 0 9
3 9 13 0
8 3 13 9 2 13 3 9 2
6 11 15 13 9 1 2
10 3 10 9 13 13 3 9 0 9 2
7 9 13 9 0 3 9 2
9 0 7 0 11 13 13 9 9 2
4 13 15 15 2
15 12 7 12 1 15 9 9 13 13 9 9 2 0 9 2
14 9 13 0 2 12 9 2 2 13 9 13 9 9 2
10 15 13 9 15 9 13 9 13 9 2
17 11 7 11 13 3 0 9 2 16 15 13 3 3 3 9 15 2
11 15 13 13 3 1 15 13 3 0 9 2
6 9 15 13 3 0 2
4 9 0 0 9
7 3 13 9 13 16 15 13
11 10 0 7 3 0 9 7 9 13 9 2
17 11 0 0 9 11 11 1 11 11 11 9 13 9 11 11 9 2
16 11 13 9 9 13 0 13 2 16 11 13 0 9 1 9 2
7 11 11 13 9 0 9 2
15 13 13 9 2 16 13 3 9 13 7 13 0 9 9 2
5 9 13 15 3 9
4 13 9 3 2
7 9 13 3 12 12 9 2
11 16 15 13 13 9 3 2 13 13 15 9
11 13 9 13 9 2 16 15 13 0 9 2
6 15 13 11 7 11 2
6 15 15 13 15 13 2
20 13 13 13 10 9 16 13 7 13 16 15 3 3 9 13 13 13 15 7 2
5 9 13 13 9 2
18 9 13 13 13 3 2 16 13 3 13 9 13 0 9 0 9 1 2
4 13 0 9 2
5 3 9 13 13 2
8 9 13 2 16 9 13 9 12
7 15 13 9 1 9 1 2
2 0 9
9 15 13 15 3 9 7 10 9 2
8 9 9 3 0 16 10 9 2
18 11 13 13 11 2 3 7 11 11 9 9 3 3 13 7 13 9 2
15 15 13 2 16 15 13 11 1 3 2 13 15 3 9 2
8 9 13 13 3 3 0 9 2
11 10 9 9 9 1 13 13 3 0 9 2
4 13 15 13 2
17 16 15 13 10 0 0 15 15 13 16 13 13 13 2 9 13 2
14 3 9 13 9 13 9 7 11 13 2 7 3 3 9
2 0 9
7 10 12 9 13 9 1 2
8 9 13 9 9 13 3 9 2
9 0 0 9 13 0 9 0 9 2
19 9 2 15 13 0 10 9 13 3 2 13 10 9 3 13 3 13 9 2
4 9 13 9 2
13 11 11 2 11 7 11 0 9 13 3 13 9 2
11 3 13 16 3 13 9 7 15 13 3 0
7 0 9 13 9 9 3 2
7 15 13 3 11 9 15 2
4 13 3 0 2
11 0 9 13 3 11 9 2 15 13 13 2
3 9 13 9
10 13 15 13 3 0 16 9 3 13 2
9 11 9 13 0 16 2 3 0 2
9 10 9 13 16 13 9 10 9 2
10 0 9 13 9 2 15 13 9 1 2
3 11 13 2
2 0 0
12 9 13 0 2 16 9 2 0 9 13 0 2
19 9 9 11 11 13 13 13 0 9 2 16 15 13 13 15 9 1 13 2
2 0 9
5 3 15 13 0 2
11 6 2 15 13 13 3 2 15 13 0 2
12 10 9 13 0 9 7 13 15 1 13 9 2
17 15 13 13 3 12 9 9 2 7 3 15 13 3 13 9 9 2
2 0 9
16 15 13 9 7 13 0 9 2 7 3 0 9 13 13 13 2
12 3 16 9 13 9 0 2 15 13 0 9 2
14 13 9 3 7 13 3 10 9 3 9 1 7 9 2
17 16 15 13 10 0 2 0 2 0 7 9 13 2 15 3 13 2
14 11 11 13 9 7 13 13 15 7 13 15 3 0 2
2 9 1
6 15 13 3 0 9 2
11 15 13 13 0 12 9 0 0 9 1 2
2 13 13
7 10 0 0 9 9 9 2
4 9 7 9 0
6 13 3 13 13 9 2
2 0 9
2 9 13
18 15 13 3 0 0 3 13 15 10 9 13 7 15 13 0 9 3 2
4 15 13 9 2
5 10 15 15 13 2
6 13 3 13 10 9 2
8 0 9 1 9 13 3 9 2
7 15 10 9 13 0 13 2
7 9 13 13 7 9 13 2
6 15 11 9 3 13 2
4 13 3 9 2
8 13 13 13 7 13 13 13 2
3 9 13 2
8 9 13 13 13 11 9 1 2
21 3 15 13 0 13 2 16 15 10 9 13 9 13 2 16 13 13 13 10 9 2
10 11 11 13 2 16 9 13 9 9 2
6 15 13 11 0 9 2
4 15 13 11 1
8 11 11 13 9 0 9 9 2
3 9 13 2
11 3 9 13 9 2 7 3 13 3 9 2
3 9 13 2
5 11 7 11 13 2
5 3 3 13 13 0
7 9 13 0 9 0 9 2
3 13 3 15
3 13 13 9
4 13 9 9 2
13 9 13 0 9 13 0 9 2 16 9 13 13 2
10 16 13 9 9 2 13 13 3 9 2
5 10 9 13 0 2
10 9 13 13 15 3 13 9 0 3 2
9 15 13 3 0 9 13 10 9 2
6 13 3 13 13 13 2
9 3 3 12 9 13 3 0 9 2
20 11 9 9 13 3 1 9 0 2 15 10 9 13 13 10 9 11 9 1 2
8 6 2 3 3 13 13 13 2
18 15 13 11 1 9 9 2 7 3 10 9 3 0 13 13 3 13 2
24 7 10 9 15 13 3 16 13 10 0 7 13 9 10 9 13 3 0 16 15 15 13 10 9
4 13 3 11 2
8 9 13 3 12 9 9 13 9
3 11 9 9
3 9 13 9
13 9 13 3 0 9 2 16 13 3 9 10 9 2
7 11 13 16 9 13 13 2
10 9 13 13 9 2 9 13 3 3 2
16 13 10 0 9 15 15 13 13 3 13 2 13 10 0 3 2
6 11 9 15 13 13 2
2 9 13
7 15 13 0 9 3 13 9
9 3 11 13 13 0 13 9 0 2
6 9 13 0 7 0 2
7 9 3 3 3 13 9 2
16 3 13 13 15 2 15 13 13 9 7 13 2 3 9 3 2
4 13 11 9 2
8 9 13 0 9 13 13 9 2
27 15 13 9 7 9 2 15 13 13 15 7 15 13 9 1 15 2 13 15 9 2 9 2 9 2 9 2
4 13 15 9 2
12 7 3 13 3 9 3 16 3 13 13 13 2
5 9 13 9 12 2
8 3 3 15 13 2 3 9 2
8 0 2 15 13 13 0 9 2
7 15 13 15 2 15 15 13
10 0 9 13 9 2 9 9 10 0 2
14 3 13 9 9 7 9 13 2 16 13 9 9 9 2
2 9 9
5 9 13 13 13 2
7 13 13 13 3 15 3 2
3 9 13 13
6 15 13 0 13 9 2
11 3 15 11 13 12 12 9 1 0 9 2
4 9 13 9 2
4 13 3 11 2
9 11 9 11 13 9 13 9 9 2
9 11 12 9 9 13 13 0 9 9
28 11 13 9 2 3 9 11 11 1 13 13 0 7 3 9 13 0 9 9 13 2 7 9 13 15 15 3 2
14 0 7 0 9 2 9 1 2 13 10 11 0 9 2
6 15 13 15 15 13 2
5 15 13 13 9 2
7 13 15 13 13 13 15 2
6 9 7 9 13 9 2
4 3 13 9 2
4 0 8 7 9
5 15 13 3 9 2
16 3 9 13 2 3 9 13 9 13 9 7 3 0 15 13 2
22 7 9 9 13 3 1 9 13 3 2 16 13 13 16 15 13 3 9 9 13 9 2
4 15 13 11 2
9 11 13 13 15 1 3 12 11 2
6 9 13 9 13 9 2
5 9 1 13 9 2
3 13 9 1
5 2 13 16 9 2
3 15 13 9
11 11 13 13 9 3 2 7 11 13 3 2
4 15 9 13 2
6 0 13 2 0 13 2
3 13 11 2
7 9 13 13 15 13 3 2
3 3 13 2
3 3 13 2
17 3 10 15 13 0 13 9 9 1 2 7 15 13 13 0 9 2
7 11 13 3 13 9 13 2
3 11 13 9
6 9 0 9 13 11 2
2 13 3
11 11 9 1 13 3 3 0 7 0 9 2
4 9 13 0 9
8 10 9 2 0 2 9 2 9
7 9 13 13 9 11 1 2
2 0 0
3 9 13 2
7 6 2 13 3 3 13 2
6 13 3 7 3 13 2
5 15 13 9 9 2
3 13 9 9
15 13 0 9 2 15 13 9 1 13 13 9 11 0 9 2
21 15 15 13 13 11 9 2 3 16 13 13 2 16 13 3 13 10 9 10 9 2
11 13 9 3 2 16 15 13 13 9 9 2
13 9 13 13 9 10 3 0 9 2 7 13 0 2
4 13 15 15 2
5 3 0 15 13 2
5 13 15 13 15 3
9 9 9 13 0 9 2 3 3 3
22 0 9 13 12 1 2 16 1 0 9 9 13 12 2 15 13 0 9 9 13 11 2
25 0 9 1 9 13 2 16 9 13 3 2 7 9 7 9 13 9 2 7 9 13 13 9 9 2
18 9 13 2 16 13 3 0 9 13 13 3 2 16 13 0 9 13 2
4 15 13 9 2
7 10 9 13 13 13 9 2
9 11 13 9 9 13 0 9 9 2
13 15 13 13 10 3 0 9 15 13 3 13 9 2
6 13 3 13 1 9 2
16 11 9 13 0 9 2 15 3 13 0 9 2 15 9 13 2
10 9 13 9 0 9 2 16 13 0 2
17 15 15 13 13 2 7 15 13 13 13 15 2 15 13 13 15 3
5 9 13 13 3 2
19 9 2 15 13 13 9 9 2 13 15 12 9 1 10 9 9 0 9 2
9 10 9 13 13 13 0 9 9 2
7 7 15 1 13 10 9 2
4 13 15 11 2
10 3 13 0 9 9 15 13 16 9 13
3 9 13 9
6 15 13 3 3 0 2
8 11 13 15 13 9 0 9 2
3 3 13 2
6 16 15 13 10 9 2
8 16 15 3 3 13 9 9 2
7 16 13 2 13 13 13 2
5 3 11 13 0 2
3 9 13 0
2 13 13
4 9 12 1 9
14 15 13 16 16 15 13 13 13 16 15 13 3 9 2
14 11 13 10 11 3 11 9 2 15 13 13 9 13 2
4 13 15 0 2
8 9 13 13 9 3 16 9 2
13 13 15 13 3 7 13 9 15 10 9 9 13 2
29 9 13 11 1 3 0 3 0 9 2 7 15 13 3 10 9 2 16 15 1 13 15 9 3 13 9 0 9 2
8 16 13 3 13 13 7 13 2
8 3 13 9 13 0 9 3 2
6 15 15 13 3 9 2
3 15 13 15
11 0 13 2 0 13 2 9 13 2 9 13
10 9 13 15 0 3 0 9 13 9 2
8 15 13 9 2 13 0 9 2
6 11 7 11 13 3 2
14 9 2 15 13 9 9 9 9 1 2 13 13 0 2
18 9 9 13 3 3 13 9 9 7 13 15 2 16 13 13 9 9 2
7 15 13 2 16 15 13 9
2 0 9
4 13 15 13 2
8 11 13 13 3 10 0 9 2
9 9 13 13 3 16 0 9 1 13
4 9 13 9 2
4 13 9 1 2
9 15 13 12 9 10 9 0 9 2
13 3 15 13 3 3 0 0 16 11 13 10 9 2
7 15 13 13 9 9 11 2
8 2 13 13 15 2 11 13 2
13 9 12 13 11 12 9 2 0 9 9 13 12 2
15 9 13 13 9 9 9 12 7 12 9 3 3 2 16 2
9 13 13 3 13 10 9 3 9 2
5 10 0 3 13 9
6 16 15 13 3 13 9
14 11 13 0 9 2 7 3 9 13 13 15 15 1 2
2 13 9
20 9 13 9 1 3 0 3 2 16 13 3 13 15 15 1 13 13 15 1 2
5 9 13 13 9 2
15 2 3 3 13 2 13 15 3 10 9 13 13 13 15 2
8 13 3 3 15 2 15 13 2
12 9 13 9 0 9 2 13 16 13 11 9 2
13 15 13 13 15 13 2 13 15 13 15 13 3 2
8 9 9 9 13 13 3 11 2
11 0 13 13 15 9 3 16 15 13 0 2
6 15 13 7 13 15 2
4 9 9 12 9
13 9 9 13 13 15 13 0 2 3 10 0 9 2
7 15 13 3 9 0 9 2
11 0 1 13 3 15 2 16 9 13 9 2
7 9 13 3 12 0 9 2
5 13 15 6 9 2
7 9 13 13 3 16 3 13
6 0 0 13 9 3 2
7 2 13 13 12 12 1 2
11 9 13 0 9 2 10 9 13 13 3 2
12 11 13 9 13 9 9 13 13 3 0 9 2
8 3 3 13 0 9 9 11 2
2 13 13
4 15 13 9 13
13 9 9 13 9 9 7 13 9 2 15 13 3 2
11 9 9 0 9 9 13 13 3 1 9 2
13 15 2 13 9 0 7 0 9 2 13 13 15 2
3 8 7 9
8 9 13 7 13 9 7 9 2
13 13 15 13 3 0 2 7 13 9 3 3 13 2
7 0 7 0 9 13 9 2
23 0 0 9 13 15 2 16 15 13 13 0 9 3 12 9 2 15 1 15 13 9 9 2
4 3 13 13 2
6 11 13 0 9 11 2
4 13 9 9 2
5 15 13 10 0 2
7 9 13 3 2 3 3 3
15 3 2 9 9 13 9 0 9 0 9 1 1 9 9 2
9 15 13 13 9 3 9 7 9 2
9 0 12 9 0 11 13 16 9 2
2 0 9
5 9 13 13 9 12
12 11 13 9 2 13 9 13 7 9 13 13 2
9 16 13 3 2 13 3 13 9 2
5 9 13 13 15 3
2 11 9
4 3 3 9 2
10 13 11 13 2 15 10 9 13 13 2
1 11
6 11 13 0 9 0 2
12 15 2 15 13 9 9 9 1 2 13 9 2
12 3 13 10 9 15 13 15 2 10 11 11 2
10 9 9 13 0 7 0 0 9 1 2
14 9 13 9 13 0 9 2 7 15 9 13 10 9 2
5 15 13 15 13 2
10 9 13 10 9 9 7 12 0 9 2
7 13 9 9 13 9 1 2
21 9 13 13 3 2 16 15 13 3 2 7 3 10 9 2 16 15 13 9 13 2
14 15 13 9 2 13 9 7 15 13 15 3 13 13 2
19 15 13 3 0 2 0 2 9 7 9 15 13 9 3 16 11 10 9 2
6 15 13 10 9 3 2
4 6 9 9 2
4 11 13 0 9
4 13 13 15 2
3 13 3 13
10 15 13 9 2 15 13 9 7 9 2
9 15 13 13 0 2 3 0 9 2
4 13 3 3 2
7 13 2 16 13 13 3 2
8 9 13 9 9 13 0 9 2
19 11 9 13 0 9 2 7 11 13 9 13 0 9 11 2 3 11 2 2
5 9 13 9 15 2
6 13 15 13 3 9 2
6 9 13 13 9 7 9
3 2 13 2
10 13 13 13 9 13 9 9 9 9 2
12 0 9 9 11 9 13 0 3 12 9 1 2
12 15 13 3 13 2 16 9 9 13 13 9 2
5 11 9 13 9 2
10 15 13 0 9 9 11 9 13 9 2
7 3 13 0 9 13 9 2
11 16 9 13 2 3 10 9 15 13 9 2
9 12 9 9 1 13 9 12 9 2
9 0 9 13 9 13 3 3 13 2
5 13 9 13 9 2
10 9 13 13 3 9 2 7 3 15 2
24 11 13 15 2 16 9 13 13 9 9 1 3 9 2 16 9 13 13 2 16 9 13 13 2
10 2 15 15 13 3 7 15 13 9 2
7 11 13 9 1 13 9 2
8 11 13 13 9 11 9 1 2
7 0 2 16 13 0 3 2
15 15 13 3 15 10 0 9 2 13 0 13 9 3 13 2
8 13 0 16 3 13 13 13 2
15 9 13 9 13 3 2 16 10 9 13 3 3 9 1 2
6 13 9 3 3 9 2
4 0 7 9 0
7 11 13 9 9 0 9 2
11 11 13 9 0 2 3 3 13 3 9 2
7 0 9 15 13 13 9 13
13 9 13 13 13 9 2 15 13 10 9 13 3 2
8 10 9 13 10 9 13 9 2
17 9 9 9 13 13 3 9 9 9 2 15 13 13 9 3 3 2
12 11 9 12 9 9 8 7 9 9 13 13 2
3 3 0 13
5 15 13 15 9 2
2 3 9
4 9 13 13 3
8 0 9 9 13 0 9 9 2
10 3 11 10 9 13 9 1 9 13 2
6 11 9 13 9 1 2
4 0 9 7 9
10 9 13 0 9 15 9 13 3 13 2
2 9 9
15 15 13 9 2 13 9 3 0 3 7 13 9 7 13 2
2 13 13
5 9 13 3 3 2
2 0 9
4 0 9 15 2
5 0 9 0 13 2
15 0 9 11 9 13 9 1 11 9 2 15 13 0 9 2
5 9 11 13 9 2
3 3 3 2
9 13 2 16 13 15 9 3 15 2
6 9 9 13 3 3 2
14 15 1 13 9 11 11 9 9 2 13 9 13 12 2
10 9 13 9 9 13 9 7 15 13 2
7 7 13 10 9 3 9 2
18 3 13 9 3 13 9 9 11 13 9 13 13 15 13 9 11 9 2
6 9 13 16 9 13 2
7 13 3 3 13 9 13 2
11 9 12 11 13 7 9 16 0 9 9 2
11 15 13 3 15 1 16 13 13 15 0 2
9 9 1 9 1 13 3 12 9 2
4 15 13 15 13
2 3 3
16 7 9 13 10 9 2 9 7 9 9 16 9 13 13 9 2
19 11 7 11 9 13 0 3 3 2 16 10 12 9 13 3 0 9 1 2
4 11 13 9 9
9 3 15 13 13 9 2 7 9 2
13 9 7 9 13 0 13 13 9 15 1 13 9 2
7 15 13 3 0 12 9 2
7 13 9 7 13 15 9 2
10 1 9 9 13 9 2 13 10 0 9
5 13 13 13 0 2
7 12 9 13 13 9 1 2
11 15 13 3 13 9 10 9 2 13 11 2
5 3 0 9 13 2
11 9 13 13 3 1 2 16 9 13 13 2
20 7 3 15 13 0 9 10 0 3 0 15 13 3 2 3 13 12 9 9 2
2 9 9
5 0 13 13 13 2
12 15 13 13 15 9 2 16 13 10 9 9 2
8 11 13 11 9 13 0 9 2
5 15 13 9 1 9
16 9 13 13 13 0 13 3 2 7 3 15 13 3 3 0 2
6 10 9 13 11 1 2
8 11 13 9 9 9 3 9 2
3 9 9 9
3 15 13 15
8 9 13 3 15 13 7 13 2
6 9 13 9 9 1 2
9 15 13 9 2 7 13 13 3 2
5 15 13 0 3 2
7 10 11 3 13 0 0 2
10 3 15 13 3 2 13 15 3 13 2
5 3 3 13 6 2
10 16 13 13 15 0 2 13 13 3 2
5 0 8 7 10 9
5 15 13 13 0 2
2 10 9
13 0 11 9 13 9 9 9 10 9 11 11 1 2
4 16 13 0 2
2 9 13
30 15 13 13 13 3 2 7 9 7 9 0 13 9 3 2 0 9 13 0 9 2 0 16 0 9 9 15 13 9 2
6 11 13 0 0 9 2
9 13 13 0 2 7 13 3 0 2
12 9 10 3 0 9 9 13 13 0 0 9 9
15 15 13 13 3 15 13 3 13 10 9 13 3 12 12 2
6 15 15 13 13 3 2
19 8 13 3 2 7 3 9 13 2 3 13 3 10 2 9 3 9 7 2
5 0 9 13 3 2
8 9 11 2 11 2 11 2 11
2 0 9
9 9 13 13 3 0 13 10 9 2
18 11 11 13 9 3 0 0 9 2 15 9 13 13 3 9 7 9 2
7 3 15 3 13 3 3 13
6 9 13 1 0 9 2
5 9 13 13 3 2
4 15 13 3 13
19 7 11 9 7 9 13 0 9 7 8 7 9 2 7 8 16 9 9 2
7 15 13 13 0 9 9 2
7 13 3 13 9 13 15 2
7 3 13 13 11 10 0 2
4 9 13 13 13
5 13 15 9 3 2
9 9 9 9 9 13 3 12 9 2
5 13 3 0 13 3
7 9 9 10 9 13 9 2
9 12 9 13 9 2 16 13 9 9
15 13 2 16 9 13 15 0 9 3 16 15 13 9 13 2
5 9 13 13 9 2
13 13 13 3 15 16 13 15 9 9 1 7 13 3
9 3 9 3 13 3 15 16 11 2
5 15 13 0 9 2
3 9 13 13
15 0 9 13 9 13 2 16 9 13 13 7 13 3 13 2
2 9 13
14 3 9 13 9 9 9 1 2 7 3 9 13 9 2
9 10 9 9 9 13 12 9 9 2
4 13 7 13 2
8 15 13 13 3 7 13 15 2
12 12 9 13 9 11 7 0 12 9 9 11 2
9 13 9 9 13 12 9 9 9 2
11 9 13 13 9 0 9 9 9 7 9 2
11 13 0 7 10 9 0 9 10 0 9 2
2 10 9
7 9 13 12 9 12 9 2
8 15 13 2 13 15 3 3 2
2 13 9
3 9 13 0
6 0 13 13 13 9 2
10 12 9 9 13 2 16 13 10 9 2
2 10 9
3 13 0 9
6 9 13 13 9 9 2
7 15 13 3 0 13 9 2
9 10 9 9 13 9 10 9 9 2
2 9 2
4 9 13 3 3
16 11 1 12 9 1 13 9 13 15 2 16 9 13 9 13 2
8 3 0 9 9 13 13 9 2
7 13 13 15 13 13 13 13
11 12 2 9 2 13 3 9 9 9 12 2
8 13 15 9 2 7 11 9 2
12 3 9 13 9 2 15 13 3 9 13 9 2
4 11 9 12 1
10 13 9 2 16 13 13 15 9 13 2
17 3 15 3 13 10 9 9 2 9 13 9 9 16 15 13 9 2
9 15 1 13 11 3 13 0 9 2
14 3 9 13 9 13 9 3 2 13 9 13 10 9 2
4 11 9 11 1
14 11 13 13 11 2 7 9 13 9 1 13 9 1 2
3 9 13 9
9 15 13 3 3 10 9 2 13 2
16 11 7 11 11 13 16 0 9 7 9 13 13 10 0 9 2
7 0 9 13 7 13 13 2
2 13 15
3 10 0 9
3 9 0 9
7 9 3 13 13 3 9 2
6 9 13 12 9 1 2
4 15 13 9 2
8 11 9 0 13 9 7 9 2
10 13 13 13 7 13 0 0 9 9 2
14 15 13 13 11 11 9 2 13 13 13 13 10 9 2
3 13 3 13
5 13 15 15 13 2
12 2 15 9 13 13 13 13 15 13 13 13 2
3 9 13 9
11 3 0 0 9 13 13 0 9 11 9 2
10 3 13 2 16 9 9 13 3 13 2
5 12 13 9 1 2
8 13 15 0 13 2 7 0 2
7 13 10 9 13 3 9 2
2 0 15
4 13 0 9 2
22 3 9 13 13 3 0 2 16 13 15 3 13 9 2 7 15 13 9 13 9 9 2
18 9 9 13 0 0 9 11 2 15 10 9 9 13 9 3 3 3 2
7 9 13 10 12 12 9 2
13 3 3 9 9 13 3 0 9 16 15 11 13 3
6 9 13 13 0 9 2
10 15 1 9 13 13 9 1 0 9 2
5 2 10 9 13 2
16 9 0 9 11 11 2 12 2 13 13 9 1 9 7 9 2
9 7 15 13 3 3 9 16 15 13
11 16 9 13 13 3 3 3 2 16 13 15
19 11 13 12 9 9 2 7 15 13 3 13 2 16 11 9 13 13 9 2
4 13 1 9 2
9 13 3 9 10 0 0 9 11 2
5 13 9 7 9 2
5 15 13 0 0 9
12 3 9 11 13 3 2 16 13 12 9 11 2
3 7 16 13
17 15 13 13 3 0 0 13 9 3 3 2 16 9 13 0 0 2
4 13 13 13 13
2 0 9
12 11 13 13 3 9 13 15 13 13 0 9 2
12 0 9 7 9 9 13 9 2 9 7 9 2
9 3 0 9 2 16 13 13 15 13
11 11 13 3 13 2 16 13 15 13 9 2
7 15 13 0 7 15 0 9
6 15 13 13 9 13 2
17 3 13 9 15 15 1 13 3 0 9 3 3 9 12 9 9 2
18 11 13 13 9 13 0 9 0 10 9 2 16 3 11 9 13 13 2
6 11 13 9 9 12 2
11 13 3 13 2 16 13 10 9 13 13 2
4 3 9 13 2
6 7 9 9 13 9 2
10 11 13 3 13 9 2 7 3 13 2
2 3 11
10 9 0 13 3 0 11 13 11 9 2
8 10 10 9 13 3 3 11 2
15 9 9 13 3 13 0 9 2 15 9 11 11 13 13 12
9 9 13 3 3 7 13 9 9 2
6 13 2 16 3 13 2
2 0 9
19 9 13 2 16 16 15 13 3 2 9 13 13 9 15 2 15 3 13 2
7 9 11 2 13 9 3 2
3 13 3 2
5 9 13 13 0 2
3 9 7 9
21 3 9 13 2 16 13 15 10 3 13 9 13 13 7 0 2 7 15 13 3 2
5 15 13 16 0 0
11 9 13 2 15 13 0 9 13 13 9 2
7 13 13 3 2 13 9 2
9 0 9 3 13 9 13 3 9 2
2 13 9
15 3 15 3 13 2 16 3 3 13 3 16 15 13 3 2
11 15 13 10 9 0 2 16 9 13 3 2
11 9 9 13 13 13 11 11 9 0 9 2
24 11 13 11 9 9 2 15 3 10 11 9 13 8 7 9 13 13 3 11 11 7 11 11 2
20 7 3 13 2 3 16 10 9 7 9 7 9 13 13 9 0 7 9 0 2
21 16 10 9 13 10 9 13 2 15 13 3 3 10 9 0 9 16 13 13 9 2
15 10 9 13 3 9 9 13 15 13 10 7 10 9 9 2
5 3 3 3 13 2
5 10 0 9 13 3
4 10 10 0 9
12 13 13 13 15 2 16 9 13 9 11 3 2
11 11 9 13 9 13 9 2 3 7 3 2
8 15 7 15 13 13 9 1 9
7 13 2 16 13 10 0 2
4 10 9 13 13
7 11 13 3 0 16 15 2
10 13 3 2 16 3 13 3 12 9 2
17 11 13 3 9 2 16 11 13 13 0 9 2 16 13 9 13 2
9 9 2 3 0 2 13 9 1 2
7 11 9 13 0 9 3 2
6 3 15 15 3 13 2
10 3 11 9 11 1 13 9 0 9 2
20 10 11 13 13 9 2 16 15 13 9 1 13 15 2 11 2 9 13 9 2
14 11 2 15 13 3 10 9 15 13 3 3 9 13 2
8 13 9 2 3 11 13 11 2
21 7 3 13 13 3 3 16 2 12 9 2 15 13 2 11 2 16 3 13 13 2
3 3 10 0
15 10 9 13 3 15 16 15 9 13 13 9 10 1 9 2
9 13 15 13 9 10 9 9 13 2
7 3 15 9 13 15 15 2
9 11 13 9 15 2 15 13 9 2
19 9 13 16 12 9 9 2 15 3 13 13 12 9 9 2 13 3 3 2
8 3 9 13 2 16 13 9 2
4 11 7 9 13
10 15 13 3 7 3 9 9 0 9 2
10 9 13 13 9 0 7 12 9 0 2
4 6 15 13 2
2 11 9
4 13 9 3 2
11 3 9 0 0 9 13 3 3 9 1 2
4 15 9 13 2
3 9 13 9
7 11 13 12 9 0 9 2
5 9 13 3 3 2
11 9 15 13 13 13 0 9 7 9 9 2
5 13 10 9 11 2
20 0 9 13 13 0 13 3 3 12 1 2 16 0 9 9 1 13 0 9 2
13 9 13 3 13 13 9 3 3 0 0 9 13 2
16 3 0 0 9 9 13 3 13 8 8 8 1 13 9 12 2
13 0 9 13 0 0 2 15 13 3 15 0 9 2
9 11 13 11 9 13 11 11 9 2
21 16 11 13 13 3 10 0 9 7 2 3 10 10 10 9 2 13 9 15 11 2
2 0 15
11 0 9 13 13 9 13 9 9 9 9 2
5 15 13 0 13 3
5 11 13 9 11 2
7 15 13 2 13 7 13 2
3 15 13 2
9 9 13 9 3 0 9 13 0 2
6 0 9 1 15 13 9
10 9 13 0 7 15 13 3 3 12 9
3 16 11 13
6 0 9 9 13 11 2
15 9 13 9 7 13 0 2 16 3 11 13 3 0 9 2
6 10 9 13 3 3 2
7 15 16 15 13 15 13 2
6 11 9 13 9 13 2
7 9 13 0 0 0 9 2
16 0 9 9 13 13 13 3 12 9 2 15 13 15 0 9 2
4 9 13 9 2
5 13 15 3 3 2
9 3 13 15 2 16 15 13 9 2
12 13 3 15 13 3 13 0 16 2 3 3 9
4 9 7 9 9
2 9 0
4 11 13 3 13
10 11 13 13 10 9 1 9 9 9 2
6 9 13 15 0 3 2
3 2 3 2
11 13 13 2 13 3 7 16 3 3 9 13
4 11 13 9 0
14 0 11 13 9 15 2 16 0 9 1 9 13 0 9
5 15 13 9 13 2
4 9 13 15 1
9 9 13 13 2 7 13 9 3 2
4 15 13 3 11
2 10 9
3 9 13 0
13 13 3 0 0 9 9 2 15 13 13 11 9 2
2 13 3
5 11 13 11 9 2
7 13 13 3 15 2 15 13
23 7 2 13 3 3 2 15 13 3 9 2 16 15 13 13 9 3 9 9 2 13 9 2
9 13 3 9 9 15 13 9 9 2
4 13 3 13 2
5 13 15 15 13 2
5 13 13 9 3 2
16 13 13 10 9 13 2 16 13 9 13 0 13 3 0 9 2
7 9 10 9 13 0 11 2
10 9 9 1 11 9 13 3 12 9 2
5 10 9 13 3 2
4 7 15 11 2
14 13 9 16 3 3 9 9 2 3 0 9 13 9 2
13 13 13 3 0 2 16 13 3 13 3 9 13 2
2 13 9
5 13 9 13 13 2
9 13 9 2 3 13 11 11 9 2
5 13 13 13 15 2
10 15 13 15 3 9 2 15 13 9 2
11 9 0 8 2 8 7 9 13 3 13 2
8 9 13 3 13 13 13 9 2
2 13 13
3 0 9 9
7 9 13 3 9 9 9 2
5 13 13 3 15 2
2 3 9
10 0 13 9 2 13 9 9 7 9 2
3 13 3 3
6 15 13 13 15 13 2
11 11 9 1 13 13 2 16 9 13 3 2
10 9 13 9 13 15 13 15 10 9 2
4 13 15 13 9
11 15 13 2 16 9 13 15 13 15 1 2
9 13 0 2 10 9 9 13 9 2
8 0 11 13 13 9 9 1 2
14 16 0 9 13 10 9 1 3 2 13 3 0 9 2
11 0 9 13 0 2 15 3 0 13 0 2
9 16 15 13 3 13 9 13 3 2
7 3 3 15 13 15 13 2
8 0 9 15 15 1 13 15 2
8 15 13 13 13 11 12 9 2
6 9 13 15 16 12 2
3 15 13 9
4 13 3 9 2
17 3 15 13 2 16 13 0 2 16 13 10 10 9 13 13 0 2
3 0 9 9
16 9 9 13 0 0 1 15 2 16 10 9 13 3 3 3 2
6 6 15 15 13 3 2
2 13 13
14 9 13 7 13 11 11 2 16 15 13 13 11 9 2
5 9 0 13 3 2
11 9 9 13 13 0 9 2 7 0 9 2
9 15 13 15 10 15 3 13 9 2
10 3 10 9 13 7 13 0 13 3 2
17 16 13 3 13 10 9 2 15 15 7 10 9 13 3 3 13 2
8 10 10 9 3 13 15 15 2
15 9 1 13 9 2 13 15 7 16 13 2 3 10 9 2
8 15 13 3 13 7 13 9 2
10 15 13 10 9 3 12 10 9 9 2
15 9 13 3 2 16 9 13 3 3 7 9 13 0 9 2
8 16 11 13 0 2 11 13 9
7 3 13 9 11 13 13 9
4 9 13 3 2
11 8 7 9 13 13 3 7 3 9 1 2
6 15 3 13 0 9 2
5 15 13 9 1 2
4 9 13 9 2
9 16 13 13 0 2 13 13 9 2
7 11 13 9 1 1 9 2
6 9 9 13 3 9 2
5 9 13 9 1 2
6 11 0 9 13 0 2
2 11 9
6 13 9 9 7 13 2
11 16 9 0 13 2 10 9 13 13 13 2
2 1 9
8 10 9 15 13 9 13 9 2
8 11 13 12 9 3 0 9 2
9 0 2 15 13 9 9 7 9 2
18 15 13 3 13 2 15 13 3 2 16 13 0 9 7 13 3 9 2
7 3 16 15 13 0 9 2
6 13 2 16 13 3 2
9 0 9 13 13 3 12 9 3 2
8 9 13 3 13 16 0 9 2
4 15 13 0 2
6 9 13 13 12 1 2
8 13 2 16 13 9 13 9 2
13 16 15 13 3 0 16 13 0 9 2 12 9 2
4 3 13 9 2
2 9 9
2 9 9
6 11 13 13 13 9 2
7 15 13 13 9 7 9 2
8 9 13 3 0 9 1 9 2
3 13 9 2
7 9 13 9 1 12 9 2
9 9 9 13 3 3 0 13 9 2
12 13 3 13 3 9 3 3 0 2 13 11 2
10 16 9 13 2 3 9 13 3 13 2
22 15 13 3 9 10 1 9 2 7 3 12 9 13 3 10 0 9 1 2 3 9 2
7 2 13 15 13 13 3 2
4 0 2 0 9
11 11 9 13 13 12 9 12 13 0 9 2
16 11 13 13 9 2 16 13 0 9 13 0 9 13 0 9 2
6 9 13 13 3 16 13
6 10 9 9 13 3 2
5 3 13 13 9 2
18 9 13 3 11 9 7 3 3 9 13 13 0 2 13 0 11 11 2
8 15 3 13 0 13 13 15 2
9 3 9 13 2 9 0 9 13 9
48 3 13 3 3 0 9 15 13 2 13 2 3 15 2 13 2 13 3 3 2 3 2 3 2 13 3 6 10 9 15 13 3 15 2 15 13 9 2 15 3 10 11 13 7 15 13 16 2
11 9 13 9 0 9 1 12 9 1 9 2
11 15 13 9 9 1 13 9 7 9 9 2
2 9 13
5 3 13 9 12 2
2 9 0
6 9 15 13 0 9 2
15 3 12 9 15 3 3 2 3 13 15 3 3 10 9 2
9 16 13 15 9 2 3 15 13 2
6 10 9 15 13 9 2
6 10 9 13 11 9 2
27 9 13 15 1 3 0 9 2 15 9 1 13 16 9 13 10 11 2 15 13 16 9 13 13 7 13 2
9 9 11 13 11 9 12 0 9 2
6 13 10 0 0 9 2
8 9 13 9 9 13 13 3 2
16 9 7 0 9 13 9 9 3 2 16 9 13 3 3 13 2
13 11 9 7 9 13 13 12 9 1 3 7 3 2
2 13 11
13 16 7 16 15 3 13 3 2 13 1 13 9 2
3 13 13 15
9 0 9 13 3 0 0 9 1 2
12 9 13 13 0 9 1 2 3 13 3 9 2
13 3 13 0 2 7 3 3 0 7 3 7 3 2
5 9 13 9 3 2
9 10 9 13 9 13 9 13 9 2
7 11 9 13 7 13 13 2
18 9 13 3 9 2 3 13 13 2 13 15 3 7 3 13 13 15 2
4 11 13 9 2
15 9 7 9 13 13 9 2 3 13 9 13 13 15 0 2
12 16 9 9 13 2 9 0 9 13 13 9 2
14 11 13 3 0 10 9 16 15 13 13 9 0 9 2
15 11 13 13 9 2 16 15 13 13 3 12 0 9 9 2
4 3 13 13 2
5 9 13 15 1 2
6 11 11 13 9 0 2
2 9 13
7 15 13 13 3 0 9 2
4 9 13 13 2
7 0 9 13 0 9 9 2
7 3 15 15 2 13 0 9
5 9 3 13 3 2
10 9 1 11 11 13 11 3 11 9 2
8 9 13 13 3 9 1 11 2
6 16 13 2 13 9 2
13 13 15 13 3 9 2 9 7 9 16 13 3 2
16 9 13 13 0 9 9 2 15 13 3 3 8 7 9 11 2
15 3 9 7 11 13 10 9 2 7 9 7 9 13 9 2
5 0 0 2 0 9
10 3 9 2 9 9 7 9 9 9 2
5 13 3 13 15 2
14 10 9 13 0 9 1 13 9 13 9 9 12 1 2
2 13 13
6 15 3 9 10 9 3
3 13 12 9
9 3 9 13 12 9 13 10 9 2
6 15 13 9 12 9 2
20 9 13 3 0 2 16 13 9 3 3 13 2 16 15 13 9 9 9 1 2
6 13 13 9 12 1 2
6 13 15 13 11 9 2
13 9 7 9 9 9 3 13 2 15 13 13 9 2
6 0 9 13 12 9 2
8 15 13 13 3 9 9 12 2
14 9 7 9 3 13 3 9 2 3 7 9 7 9 2
9 13 13 10 9 2 15 13 15 2
10 10 9 13 3 0 0 7 3 9 2
5 10 9 13 0 2
7 16 15 3 13 15 15 2
11 0 3 13 13 9 0 9 7 0 9 2
12 13 0 7 13 9 0 3 0 9 13 11 2
8 11 9 13 11 11 9 9 2
5 9 13 0 9 2
6 15 13 12 9 9 2
9 10 9 1 13 3 10 12 0 9
3 9 13 9
5 12 13 3 9 2
8 16 9 13 2 15 13 0 2
2 10 9
13 9 13 9 3 9 12 9 3 9 9 9 12 2
14 0 9 3 13 2 3 13 13 13 9 9 7 15 2
4 9 15 13 2
5 13 3 11 13 2
5 15 3 13 0 9
2 0 9
7 13 9 9 2 2 9 2
10 11 1 0 9 13 13 3 0 9 2
22 3 13 9 1 13 9 13 9 0 9 2 13 2 9 2 0 9 13 13 0 9 2
2 13 13
6 15 3 2 0 9 2
7 9 9 13 9 9 1 2
3 9 13 2
2 0 9
4 2 13 15 2
68 3 10 0 15 13 13 3 2 15 3 13 10 2 9 9 7 9 16 2 8 2 15 13 3 0 16 15 8 2 13 3 3 15 13 3 15 2 15 2 15 13 3 10 9 13 7 9 7 2 0 0 9 15 3 3 13 8 2 15 13 10 9 13 3 12 12 7 2
7 15 1 15 13 13 13 2
8 7 13 3 11 13 3 0 2
16 9 7 9 10 9 3 13 9 9 3 9 13 3 9 3 2
3 13 3 2
7 13 13 13 15 0 9 2
20 3 13 9 3 7 3 3 13 2 10 9 13 3 13 13 2 13 11 9 2
10 7 15 9 13 2 13 15 7 13 2
19 13 13 2 16 0 9 13 13 3 13 15 2 3 0 9 9 9 13 2
11 15 13 7 13 9 2 16 15 13 9 2
5 13 15 3 9 2
2 0 9
4 9 0 0 9
8 15 13 13 13 13 9 9 2
6 6 9 13 9 3 2
11 0 9 9 3 9 1 2 0 0 9 9
8 10 9 13 3 13 1 9 2
5 9 9 1 9 2
4 9 13 9 2
17 9 13 0 13 9 9 9 1 2 16 15 13 13 9 9 9 2
5 13 15 13 13 2
3 13 15 2
5 9 9 13 3 9
14 11 13 9 13 9 2 7 3 9 13 13 9 1 2
21 16 13 13 10 9 3 3 9 2 13 9 0 9 3 7 9 13 15 13 3 2
2 0 9
8 9 9 13 3 3 3 9 2
10 15 13 9 1 7 13 9 9 3 2
4 9 13 9 2
7 3 11 13 15 1 9 2
3 9 0 9
5 9 9 13 13 2
11 9 13 9 7 9 13 3 3 3 2 2
5 13 10 9 13 3
5 9 13 13 15 2
7 3 9 9 13 3 0 2
11 9 13 3 12 0 9 2 15 15 13 2
18 11 13 13 13 13 9 11 2 11 13 13 2 16 13 9 9 13 2
10 11 13 9 10 0 9 12 9 1 2
11 16 3 3 13 3 9 15 12 9 3 2
32 13 3 10 11 11 15 13 6 15 13 9 7 13 15 9 15 15 13 13 7 9 13 10 11 15 13 0 3 9 9 11 2
13 3 12 9 9 2 15 13 13 3 3 16 13 2
13 2 13 13 13 3 10 9 7 12 0 9 2 2
13 12 9 13 9 9 13 0 9 9 9 7 9 2
6 13 11 9 7 9 2
10 3 9 13 2 9 13 3 9 9 2
2 13 3
14 13 15 3 9 7 2 9 7 9 16 15 13 3 2
5 3 15 3 13 2
14 9 9 13 0 9 3 16 13 13 3 3 13 15 2
13 0 3 13 9 9 1 2 16 15 13 3 3 2
7 9 13 13 12 9 1 2
15 3 16 13 3 2 0 9 2 9 7 9 13 10 9 2
15 9 9 13 9 13 9 2 15 13 3 13 9 15 13 2
4 15 13 9 1
14 11 13 9 13 3 12 3 13 12 9 13 12 1 2
13 9 13 9 7 3 13 9 9 9 13 9 9 2
4 9 13 9 2
4 15 13 0 9
7 9 11 9 13 3 0 2
14 13 13 3 9 13 2 16 13 13 16 13 9 9 2
6 13 13 9 13 13 2
4 13 3 3 2
5 11 13 13 9 2
17 11 13 13 9 2 7 3 0 2 16 15 13 13 0 9 13 2
3 15 1 16
5 11 13 13 13 9
10 11 13 13 9 9 7 13 0 9 2
12 13 15 13 13 13 9 9 3 7 13 9 2
4 3 3 13 2
10 16 9 13 3 2 13 3 13 9 2
6 9 13 3 9 0 2
6 13 13 3 9 12 1
5 3 3 9 13 2
18 13 10 0 9 10 9 2 16 13 9 7 9 1 13 15 13 3 2
9 10 10 9 9 13 3 13 9 2
3 13 9 2
6 10 9 13 3 6 2
7 3 9 13 13 0 3 2
17 15 13 2 16 11 9 13 3 3 3 10 9 16 15 13 9 2
10 9 9 7 15 9 1 9 13 9 2
5 7 15 10 0 2
5 0 9 3 13 2
10 3 9 2 15 13 13 3 3 13 2
5 11 7 11 13 9
8 15 13 3 13 13 11 1 2
7 13 3 9 9 15 1 2
5 2 13 16 15 2
3 9 13 2
6 3 13 12 0 9 2
6 0 9 15 13 0 2
6 9 13 3 9 9 2
2 10 0
14 12 0 9 13 7 13 3 9 9 3 3 12 9 2
9 9 2 15 9 9 13 3 13 2
9 9 9 9 13 3 10 0 9 2
7 13 15 13 13 15 9 3
8 11 13 3 13 13 9 9 2
12 9 13 9 2 16 9 9 13 9 13 12 2
12 9 13 0 12 9 0 9 16 10 0 9 2
2 3 11
6 9 13 9 13 9 2
3 9 3 11
12 3 16 9 13 9 2 13 2 9 9 2 2
8 9 13 13 3 3 15 1 2
2 6 9
3 9 13 9
15 9 9 13 15 2 13 9 13 9 9 13 7 13 9 2
6 6 2 6 3 3 2
9 15 13 9 9 3 16 9 11 2
3 13 9 2
3 13 3 2
2 9 13
13 13 3 13 0 9 7 15 13 13 2 9 13 2
14 0 9 11 13 13 2 16 15 13 13 9 1 9 2
11 11 9 1 13 13 9 0 9 9 9 2
4 9 0 9 9
4 9 13 3 2
9 15 13 9 9 7 13 13 9 2
18 16 10 9 13 13 9 3 15 13 9 16 15 13 7 3 3 13 2
14 9 13 9 2 3 3 13 9 1 9 2 3 9 2
7 15 13 15 7 15 9 2
15 16 10 9 9 13 13 2 15 13 10 3 9 9 9 2
8 15 13 13 15 13 0 9 2
15 7 3 6 11 11 2 15 13 3 13 0 3 9 3 2
11 10 9 13 3 13 13 15 9 0 9 2
11 15 13 9 0 9 2 7 13 15 13 2
12 13 9 13 0 9 2 9 7 9 7 9 2
9 13 3 2 9 3 13 11 1 2
5 9 1 13 9 2
9 10 9 13 11 7 15 9 11 2
4 15 13 3 2
3 13 3 2
5 9 13 12 9 2
25 13 15 0 9 2 16 13 7 13 2 3 9 13 9 2 15 13 13 10 9 2 13 3 0 2
3 15 13 2
16 15 13 9 13 9 3 7 13 9 10 9 2 16 15 13 2
21 9 13 13 9 9 9 1 2 7 16 13 13 9 9 13 3 10 9 13 9 2
3 15 13 15
3 9 13 15
10 3 15 13 15 13 2 16 13 13 2
9 13 13 15 2 16 15 13 13 2
16 12 0 9 13 9 1 9 2 9 2 9 2 9 7 9 2
3 15 3 2
2 13 9
5 9 13 9 1 2
5 13 13 16 9 13
14 9 13 13 2 15 13 9 2 0 9 7 9 1 2
2 12 12
4 11 13 9 2
7 0 9 9 15 3 11 2
7 13 2 16 15 13 3 2
6 15 13 0 9 13 2
11 9 9 13 9 11 1 3 11 7 11 2
7 9 0 3 12 9 13 9
12 0 9 13 0 13 9 16 13 15 0 9 2
25 13 13 9 13 2 3 2 0 9 2 13 13 2 3 7 3 2 3 7 3 2 3 7 3 2
4 16 3 13 13
16 9 9 13 9 2 15 1 11 9 13 3 11 13 9 9 2
11 13 10 0 9 2 15 13 13 9 9 1
5 9 13 3 0 2
8 13 0 9 2 15 3 13 2
11 13 0 13 2 13 10 9 13 0 9 2
11 9 13 10 0 9 13 9 0 7 9 2
3 10 9 9
13 3 12 0 9 12 9 2 7 3 13 0 9 2
2 12 12
12 15 13 3 0 13 2 7 15 13 3 9 2
2 9 9
13 11 11 13 13 15 9 2 9 2 9 7 9 2
6 9 7 9 13 3 2
5 0 9 13 9 9
3 13 9 9
10 9 13 3 13 2 7 15 13 9 2
15 15 13 9 0 15 13 13 2 15 13 11 7 13 15 2
6 15 13 16 15 15 13
15 13 3 12 9 15 13 9 13 2 13 2 13 7 13 2
14 13 15 3 13 2 16 13 9 11 7 13 9 3 2
3 13 13 2
9 9 7 9 13 15 3 0 9 2
17 9 13 2 16 11 13 9 9 2 16 9 10 9 13 3 0 2
5 9 13 16 9 2
21 11 9 13 9 2 11 9 2 11 9 7 9 2 11 9 7 11 7 11 11 2
2 6 16
9 3 15 3 13 13 3 9 3 2
8 13 9 7 3 9 13 9 2
7 3 0 13 0 0 1 2
8 15 13 9 9 11 7 11 2
15 11 15 13 2 16 13 9 13 13 9 9 13 3 13 2
4 13 9 3 2
9 12 0 9 13 9 9 1 11 2
8 13 9 9 9 7 13 9 2
10 13 9 0 9 13 13 0 9 9 2
7 3 15 13 3 13 3 2
3 9 13 2
8 9 13 16 13 9 13 9 2
6 10 9 15 13 13 2
2 13 3
12 11 13 11 11 13 13 10 9 9 0 9 2
5 10 9 3 13 2
8 13 9 3 3 3 16 9 2
2 9 9
11 16 11 13 13 3 2 15 13 13 9 2
9 16 3 13 13 2 13 13 9 2
13 10 9 15 13 2 16 0 9 13 9 0 9 9
2 15 13
16 11 13 0 9 13 3 9 2 7 11 11 13 13 15 15 2
12 11 13 3 12 9 1 13 3 0 16 3 2
5 0 9 7 9 2
11 16 15 13 9 13 3 15 13 16 13 15
2 9 9
5 15 13 3 13 2
10 16 13 13 15 2 3 15 13 13 2
5 13 9 10 9 2
13 15 13 3 2 3 3 2 16 15 13 13 9 2
13 13 9 7 9 13 7 13 11 8 7 9 1 2
8 13 15 13 2 16 13 15 2
6 13 12 9 9 9 2
12 11 9 13 9 13 9 0 9 7 9 9 2
16 9 13 13 3 9 2 7 3 9 9 2 15 13 13 13 2
14 6 15 13 9 3 9 7 15 3 13 0 12 9 2
6 10 9 13 12 9 2
9 9 13 3 13 3 3 9 0 2
3 9 7 13
12 15 13 3 15 2 13 11 0 7 0 9 2
13 15 13 13 2 11 11 2 7 2 11 11 2 2
2 13 9
6 13 3 9 13 9 2
13 15 15 2 15 13 3 13 13 3 9 9 0 2
11 15 15 13 3 16 13 15 13 13 13 9
9 16 9 13 0 2 13 9 3 2
9 9 9 13 0 0 13 9 13 2
9 9 11 1 9 13 0 0 3 2
13 0 9 9 13 9 2 16 3 9 13 9 9 2
9 3 3 13 16 11 13 13 9 2
8 13 13 2 16 13 13 13 2
8 9 13 7 13 9 12 9 2
18 15 13 15 3 0 7 3 0 2 0 0 2 0 9 7 0 9 2
6 12 9 13 9 1 11
12 13 13 0 9 15 1 2 16 13 13 9 2
12 11 13 9 13 15 2 15 13 9 13 2 2
6 3 9 13 0 3 2
3 9 9 2
7 15 13 13 3 12 9 2
5 0 9 13 0 2
7 0 9 9 9 9 3 2
5 13 9 9 9 2
12 15 13 15 13 9 15 2 15 15 13 13 2
17 9 13 13 9 3 13 2 15 13 13 9 7 15 13 15 15 2
7 3 13 13 9 9 15 2
5 9 13 13 15 2
3 9 9 9
4 13 15 0 2
18 3 10 9 13 13 3 3 2 7 13 3 15 1 2 16 15 13 2
11 10 9 0 9 9 9 9 13 9 9 2
12 7 3 13 3 13 2 7 15 13 15 9 2
7 9 13 13 9 13 9 2
14 11 2 11 7 11 9 13 13 12 9 0 9 9 2
6 3 15 13 13 3 2
6 9 13 9 13 11 2
13 9 1 13 3 9 2 9 2 9 7 9 9 2
8 15 13 9 2 7 13 9 2
14 11 13 16 13 15 0 2 0 9 10 15 9 13 2
14 6 15 13 3 3 10 9 16 9 13 3 3 9 2
8 15 13 3 0 16 9 13 2
12 15 13 13 2 15 15 13 15 15 13 13 2
8 15 10 9 13 13 13 3 2
10 15 3 13 3 2 9 3 3 3 2
4 15 13 9 1
7 11 11 13 13 10 0 2
2 13 3
14 3 9 13 13 2 16 10 9 13 9 1 13 9 2
5 9 13 13 0 2
2 13 9
12 13 15 10 9 2 3 15 13 3 13 9 2
4 15 13 15 3
8 13 9 9 3 16 9 13 2
6 13 9 3 15 13 2
9 3 9 13 13 13 3 0 9 2
5 15 13 15 0 9
12 13 3 13 2 16 11 13 9 7 13 9 2
12 9 1 13 9 2 16 10 9 13 13 13 2
19 3 13 13 9 15 2 3 9 9 13 2 9 7 9 7 9 7 9 2
6 11 13 11 10 9 2
4 0 15 13 2
3 0 10 9
11 15 13 13 15 9 3 16 15 13 13 2
2 9 9
11 3 9 9 13 9 13 9 3 0 9 2
9 3 15 13 9 9 9 7 9 2
8 13 3 3 2 3 13 3 2
18 16 13 13 7 13 0 9 13 13 13 9 11 7 13 13 13 9 2
22 7 15 13 10 9 13 7 16 13 10 10 9 13 2 10 9 3 15 13 3 13 2
7 16 13 2 3 13 2 2
5 13 2 15 13 2
10 13 13 9 7 9 13 15 0 9 2
15 9 10 9 13 9 2 9 7 9 13 2 3 9 13 2
3 9 13 9
10 9 13 0 2 16 15 13 13 13 2
6 11 9 13 3 0 2
9 8 7 9 13 13 3 13 3 2
9 9 13 9 13 9 8 8 8 2
12 10 9 13 0 9 2 10 10 2 9 9 2
5 0 9 13 0 2
7 9 11 13 0 9 11 2
14 3 10 2 12 3 16 3 3 3 7 2 3 3 0
5 13 9 9 9 2
4 13 15 15 2
3 9 13 9
11 9 13 13 9 2 9 2 9 7 9 2
6 15 13 13 9 9 2
12 13 15 2 16 9 9 13 11 9 13 0 2
13 11 1 13 12 9 3 9 16 10 9 1 3 2
5 13 10 9 3 2
8 13 13 2 15 15 13 13 2
12 16 9 13 13 9 2 9 15 13 7 13 2
2 9 9
14 13 16 3 15 3 3 13 10 9 13 3 9 3 2
6 9 1 9 13 9 9
3 9 9 9
10 9 13 3 9 7 9 13 0 9 2
7 13 3 3 13 0 0 2
13 15 1 3 15 3 3 13 2 15 15 13 9 2
16 0 0 9 9 2 15 13 9 15 9 2 13 3 0 9 2
8 13 9 3 2 7 13 9 2
10 15 3 13 2 16 0 9 13 13 2
7 15 13 0 13 3 9 2
14 13 13 3 15 13 2 15 13 13 9 12 9 9 2
5 15 13 0 9 2
11 9 9 2 9 11 11 13 0 9 11 2
5 15 1 13 0 13
7 13 15 3 13 9 13 2
10 9 9 13 0 2 15 13 15 9 2
3 0 0 9
9 9 0 9 9 13 0 9 9 2
8 9 13 13 10 0 13 9 2
12 3 9 13 0 7 9 13 0 9 13 0 2
9 3 9 13 13 3 9 7 9 2
5 3 0 15 13 2
4 3 13 0 9
10 15 13 0 9 15 13 3 0 9 2
10 9 13 3 13 2 10 9 15 13 2
3 13 15 1
3 9 7 9
14 7 10 9 7 9 15 13 9 2 16 13 13 9 2
15 7 13 13 9 1 2 7 13 3 2 15 9 13 9 2
11 9 9 7 9 13 13 10 9 10 9 2
6 15 13 13 13 13 2
9 13 3 0 9 3 2 13 11 2
20 3 3 3 15 13 3 13 13 16 13 3 13 13 3 16 0 9 13 3 2
7 9 13 9 7 9 9 2
8 9 11 2 3 13 13 9 2
3 13 9 1
9 3 13 3 0 12 9 0 9 2
10 11 13 0 1 3 3 16 13 13 2
9 3 13 13 2 15 11 13 13 0
10 13 9 2 16 13 9 13 13 3 2
4 11 13 13 0
6 9 13 3 9 1 2
4 9 13 3 2
3 13 9 9
11 13 9 13 12 9 2 15 13 3 12 2
5 15 13 13 3 2
2 13 13
6 9 7 9 13 3 2
6 10 9 15 15 13 2
5 9 13 9 1 2
13 16 3 13 0 13 3 13 13 13 15 7 15 2
5 3 3 0 9 2
9 9 2 15 13 0 9 7 13 9
8 10 9 13 13 0 7 0 2
2 10 9
14 11 9 13 3 0 2 7 9 15 13 0 16 9 2
5 9 13 3 9 1
3 9 9 1
11 9 9 9 13 3 15 16 11 11 9 2
7 13 9 9 13 13 9 2
4 9 13 0 2
6 13 16 15 13 9 2
6 13 13 13 3 3 2
22 16 11 12 13 11 11 2 11 9 7 3 10 9 13 0 7 0 9 13 9 9 2
4 13 15 13 9
7 9 11 9 12 13 9 12
9 10 10 9 13 13 10 9 15 2
7 15 13 3 0 13 0 2
13 3 15 13 13 9 13 13 15 16 13 15 11 2
10 15 13 13 15 3 2 13 3 3 2
4 15 13 1 9
8 15 13 9 3 3 8 9 3
7 0 9 13 9 3 9 2
12 11 7 10 9 13 13 0 9 2 0 9 2
5 0 0 7 0 9
10 13 3 3 13 2 15 13 7 13 2
5 0 9 2 0 9
4 13 3 3 2
13 9 1 13 9 9 3 9 7 0 9 9 11 2
9 11 11 9 9 13 3 12 9 2
7 13 13 9 13 3 13 2
7 0 15 13 16 9 9 2
11 10 15 13 9 13 0 9 13 3 0 2
5 0 9 13 9 2
8 10 9 9 13 3 15 13 2
2 0 11
6 15 13 0 9 13 2
4 9 1 13 2
5 3 11 13 3 2
10 3 9 13 0 13 9 0 9 1 2
16 13 13 13 2 13 9 3 0 9 2 9 9 13 11 13 2
7 9 15 13 3 10 11 2
6 13 3 3 10 11 2
6 9 13 2 13 7 13
8 13 3 15 2 15 13 13 2
9 0 3 2 8 11 13 0 9 2
9 7 3 3 1 9 13 3 13 2
11 9 11 9 11 9 13 13 11 9 9 2
9 15 13 0 7 0 9 9 7 9
13 3 15 13 13 9 2 16 9 13 3 9 1 2
8 15 13 9 7 13 13 9 2
3 9 13 3
14 13 15 3 3 0 13 16 3 13 0 3 9 13 2
22 11 9 13 3 11 2 15 15 13 9 2 15 11 2 11 7 11 9 13 15 9 2
11 9 13 3 12 9 0 2 0 7 0 2
16 2 16 15 13 7 13 10 9 16 15 13 13 2 6 13 2
2 12 9
12 15 13 13 9 0 9 9 13 7 9 11 2
5 10 9 9 13 9
9 11 9 13 3 3 0 7 13 2
13 11 13 2 16 15 13 0 9 10 9 9 9 2
16 9 13 13 10 3 3 9 13 7 9 13 3 0 9 1 2
8 11 13 11 9 0 12 9 2
11 15 13 0 9 16 13 15 13 10 9 2
8 9 9 13 9 3 9 12 2
9 11 9 13 9 2 7 11 13 2
12 9 2 8 8 2 13 13 3 7 11 7 11
8 9 9 13 3 3 0 9 2
9 10 10 9 3 15 13 3 0 2
5 9 13 3 9 2
2 13 3
3 0 9 2
3 15 13 9
10 13 13 9 2 16 13 13 11 9 2
11 9 13 9 12 3 12 9 0 9 9 2
15 9 13 13 3 0 2 7 9 9 11 11 13 9 9 2
5 15 15 13 9 2
10 13 9 13 9 13 0 1 0 9 2
6 15 13 3 0 9 2
5 9 2 13 3 2
6 13 13 3 9 12 1
13 15 13 13 10 15 2 15 13 13 7 15 13 2
15 11 9 13 0 2 16 3 11 9 13 13 9 15 0 2
5 13 3 3 15 2
11 9 11 11 9 13 11 0 7 0 9 2
5 15 13 3 9 2
5 15 13 3 9 2
10 0 9 9 13 9 12 9 1 9 2
4 13 10 9 3
15 16 15 13 13 15 2 16 15 13 9 2 11 13 3 2
3 13 9 2
23 11 11 13 13 9 3 2 16 15 13 9 9 0 2 15 13 13 3 13 13 9 9 2
4 13 7 13 2
13 9 13 9 0 9 2 10 9 9 12 9 9 2
7 3 10 9 13 15 15 2
7 16 13 0 2 13 0 13
2 9 13
8 3 16 9 13 3 15 3 2
14 3 3 9 9 13 15 2 16 9 13 9 3 0 2
5 11 15 13 9 2
5 10 9 13 9 2
4 3 13 1 9
13 15 13 9 2 16 13 3 3 9 9 10 11 2
17 10 9 0 9 13 9 0 9 2 15 13 13 13 7 13 15 2
5 15 13 3 3 2
5 15 13 9 0 2
12 9 13 0 0 13 0 9 13 9 0 9 2
5 9 1 13 9 2
14 11 13 15 13 9 9 2 16 9 13 3 9 1 2
9 9 13 11 0 9 1 0 9 2
4 11 13 13 2
5 15 13 13 9 2
8 9 9 13 3 3 9 9 2
3 3 15 13
10 13 13 13 2 16 15 13 0 9 2
9 0 13 2 13 2 11 3 0 2
2 3 2
4 9 13 0 2
3 10 9 2
12 3 0 7 3 0 9 9 13 10 9 3 2
11 9 9 13 3 9 9 9 2 9 13 2
15 11 13 10 9 2 15 13 11 11 12 0 0 9 9 2
6 9 13 13 7 9 2
15 15 1 9 13 15 2 16 9 0 9 9 13 13 3 2
13 11 9 13 12 13 13 3 9 2 13 13 13 2
38 7 13 0 9 9 9 2 11 11 9 2 16 9 13 11 9 2 11 11 9 2 16 9 13 9 2 11 11 0 0 9 2 16 9 13 0 9 2
5 6 13 13 3 2
4 15 13 9 2
5 13 3 10 9 2
16 13 3 0 2 16 13 0 9 11 2 15 13 0 9 9 2
4 6 15 9 2
15 3 13 9 13 13 9 1 2 15 13 13 12 9 9 2
7 15 13 15 0 0 9 2
11 11 13 3 0 9 1 8 7 3 9 2
6 9 13 13 3 9 2
16 15 13 13 2 13 15 0 9 7 13 15 3 3 9 11 2
9 13 2 16 0 9 13 3 15 2
5 9 15 13 9 2
6 15 13 13 9 1 9
25 9 11 12 13 11 11 9 9 7 13 15 11 2 3 9 11 7 0 0 9 2 9 2 11 2
8 9 9 13 13 10 9 9 2
12 13 2 16 0 9 13 15 9 9 9 11 2
9 11 9 13 9 0 0 7 0 2
5 9 9 9 1 13
10 15 13 9 0 9 11 7 9 9 2
9 15 13 15 0 9 13 9 9 2
8 16 13 2 13 15 0 3 2
7 11 13 13 7 13 13 2
10 11 9 13 11 13 9 7 0 9 2
7 9 13 9 0 9 11 2
12 15 13 13 9 2 0 13 13 3 13 3 2
18 9 9 15 15 1 15 1 13 13 9 2 16 9 13 0 9 9 2
10 15 9 1 13 13 15 9 12 9 2
7 0 9 13 3 15 1 2
18 9 9 9 13 2 3 13 9 12 9 2 2 16 15 13 10 9 2
13 11 8 7 9 9 9 13 9 13 10 9 9 2
6 9 13 0 13 9 2
2 9 9
4 15 13 9 13
2 0 13
5 9 13 0 9 2
28 15 13 13 9 0 9 15 13 3 11 11 9 15 13 9 7 9 15 9 7 3 3 13 6 6 7 9 2
9 9 1 13 0 9 0 9 1 2
11 9 13 3 0 2 0 16 15 13 13 2
10 0 3 3 13 9 9 13 10 9 2
7 13 13 3 9 9 3 2
14 16 0 9 9 9 13 11 13 2 3 3 9 13 13
8 3 13 3 9 0 3 9 2
10 9 13 9 9 7 3 3 9 1 2
5 9 1 13 9 2
3 9 7 9
18 9 13 12 9 0 0 12 9 1 2 3 9 13 13 3 9 13 2
6 11 9 13 13 0 2
4 12 13 9 2
11 9 13 13 9 2 7 15 13 9 13 2
9 13 13 2 16 0 13 0 9 2
3 9 0 9
14 13 15 3 13 13 2 3 16 10 9 13 0 9 2
2 0 0
6 7 3 15 13 15 2
5 12 9 0 9 9
6 9 13 3 0 9 2
3 9 13 0
10 9 0 9 1 8 8 7 11 9 2
6 15 15 13 2 13 2
3 9 13 0
2 0 9
7 9 13 13 13 13 1 9
6 13 9 9 7 13 9
12 3 9 13 0 9 2 15 13 9 7 9 2
3 13 13 13
6 15 13 0 9 13 2
4 15 13 9 11
8 15 13 15 2 3 9 13 2
7 9 9 13 13 0 9 2
3 3 9 2
4 13 13 3 2
12 10 9 13 12 9 3 16 10 0 9 13 2
5 11 13 11 1 2
7 12 9 9 11 0 9 1
10 9 9 13 10 12 9 9 3 9 2
6 9 9 13 13 3 2
3 9 9 9
2 3 0
8 9 7 13 9 1 7 1 2
5 9 13 3 9 2
6 0 9 13 3 3 3
4 9 13 13 9
4 9 13 0 2
10 3 15 15 13 2 16 15 9 13 2
5 9 13 12 12 2
4 3 15 13 2
8 3 2 15 13 13 10 0 2
19 13 13 2 16 9 13 3 3 13 10 9 13 9 7 13 0 9 9 2
12 15 13 11 13 3 9 15 3 13 0 9 2
7 11 13 9 3 1 9 2
23 7 16 9 13 13 3 9 2 13 15 13 9 2 16 9 9 13 13 13 13 7 13 2
7 3 9 13 3 9 9 2
14 2 16 13 13 10 9 2 7 15 13 12 9 3 2
3 9 3 9
6 9 13 13 13 9 1
6 15 13 8 3 9 3
4 10 9 13 0
6 13 9 13 13 9 2
12 9 9 1 13 13 12 16 13 3 12 12 9
16 0 9 13 9 11 2 10 0 9 9 13 13 9 0 9 2
8 7 3 13 3 16 9 9 2
16 11 13 0 9 9 2 16 15 13 13 9 9 7 9 9 2
7 9 13 13 9 7 9 2
4 13 6 3 3
3 9 15 9
7 13 2 16 15 13 3 2
12 9 13 3 0 0 9 2 0 11 3 13 2
7 9 9 13 10 9 0 2
12 15 13 3 3 15 3 15 13 13 10 10 9
6 9 0 9 13 9 2
6 15 13 9 13 9 2
2 9 9
17 15 1 13 3 13 2 16 13 15 15 12 9 13 7 15 13 15
4 9 13 15 2
5 10 9 13 15 2
3 15 13 15
13 15 2 13 9 7 13 2 13 11 7 11 1 2
9 9 13 9 13 2 15 15 13 2
11 11 13 9 9 9 7 15 13 9 3 2
4 0 9 9 13
2 9 9
11 11 9 7 9 13 3 0 9 0 9 2
6 3 9 13 9 3 2
8 3 13 15 13 13 15 9 2
15 9 13 13 9 3 2 16 15 13 0 9 10 9 1 2
4 9 13 13 9
6 7 13 13 9 9 2
20 3 15 13 3 0 9 2 16 13 15 15 3 13 2 3 15 15 3 13 2
2 3 3
9 9 9 13 13 13 3 12 9 2
7 3 0 9 9 13 9 2
14 0 9 3 13 9 2 16 3 13 13 15 13 9 2
5 1 9 13 9 2
12 13 15 3 9 13 2 16 9 13 13 0 2
12 13 3 0 9 9 2 16 13 0 9 13 2
3 13 13 13
3 9 9 9
2 0 9
17 9 9 13 9 9 0 9 13 9 9 2 9 2 9 7 9 2
7 15 13 13 13 10 9 2
12 15 13 9 3 3 3 2 16 13 13 9 2
14 9 13 3 13 9 2 15 13 13 13 13 0 9 2
7 9 13 0 9 11 11 2
12 9 13 13 3 2 16 3 13 13 13 13 2
5 15 13 3 3 2
16 9 13 11 11 11 11 2 15 13 9 2 16 13 9 1 2
4 15 13 9 1
5 9 9 13 13 0
4 12 9 13 3
7 12 9 13 13 9 13 2
19 11 2 12 2 11 7 11 12 9 0 2 13 0 9 0 11 11 1 2
7 15 13 13 0 2 0 2
10 9 13 3 13 13 11 9 9 9 2
9 9 13 9 7 15 1 13 9 2
7 13 13 9 0 11 1 2
10 13 2 11 2 13 13 12 9 9 2
3 9 13 0
4 9 13 9 2
8 16 13 9 3 2 9 13 2
4 9 13 9 2
7 15 13 3 3 0 9 2
3 0 9 2
17 9 13 9 7 9 13 15 2 16 2 13 3 15 15 13 2 2
6 0 9 9 13 9 2
13 13 9 13 9 10 9 1 2 16 9 13 13 2
6 3 3 13 9 1 2
12 7 3 15 13 2 16 9 1 13 0 13 2
12 12 9 9 9 13 2 16 15 13 9 13 2
5 15 13 9 13 9
3 9 0 9
5 2 13 15 9 2
20 15 13 9 2 13 9 7 13 9 9 2 15 11 11 13 11 12 9 12 2
11 9 9 13 9 13 9 13 11 3 9 2
3 11 9 2
10 3 13 0 9 13 9 2 3 9 2
6 10 9 13 10 0 2
8 9 9 9 9 13 0 9 2
5 3 3 13 3 2
3 9 13 9
13 9 9 1 13 13 12 16 13 3 12 12 9 2
11 13 13 13 10 9 7 3 13 13 15 2
7 7 9 13 9 0 9 2
3 9 13 15
19 13 3 10 9 13 13 2 7 3 13 13 13 0 9 3 9 7 9 2
7 11 13 0 9 13 9 2
13 16 9 13 13 9 3 13 9 7 13 9 3 2
7 13 15 15 3 2 3 2
7 0 9 13 9 10 9 2
10 6 3 15 13 0 0 2 9 3 2
4 13 15 0 2
8 9 9 13 0 9 13 12 2
16 3 10 12 9 7 3 10 12 9 0 9 13 3 9 13 2
5 16 13 0 0 2
4 13 15 9 2
8 15 13 15 13 3 9 11 2
7 9 9 13 3 3 9 2
4 9 13 3 2
4 9 13 9 2
4 15 13 15 9
3 3 13 2
6 13 13 3 0 9 2
11 6 2 3 15 9 13 2 9 13 9 2
14 9 13 9 13 9 13 2 16 15 13 13 9 9 2
4 3 15 3 9
7 13 3 13 3 15 13 2
5 9 13 11 9 2
2 3 3
12 9 13 3 13 2 16 0 7 9 13 0 2
8 11 13 3 13 2 3 13 2
22 3 12 13 9 13 13 13 0 9 2 16 0 9 9 7 9 9 13 13 0 9 2
2 0 9
2 0 9
7 15 13 10 9 13 9 2
4 13 9 7 9
22 13 13 3 9 10 9 2 10 9 15 1 2 15 15 13 10 9 1 2 15 3 2
10 15 9 13 2 16 13 3 0 9 2
9 0 9 15 3 13 2 11 13 2
8 0 9 13 9 1 12 9 2
3 13 13 2
9 6 3 2 15 13 10 9 15 2
2 12 9
7 11 13 10 9 11 9 2
7 10 9 10 9 13 13 2
3 9 13 9
5 13 0 9 11 2
4 10 9 2 16
13 15 3 13 3 2 6 6 16 15 13 3 9 2
14 6 6 2 13 3 0 16 13 9 9 2 16 13 2
6 9 13 9 12 9 2
9 16 15 13 3 3 3 13 15 2
2 9 9
11 9 13 9 2 16 3 9 13 13 3 2
6 9 13 9 13 9 2
2 9 1
4 3 10 0 2
12 9 2 15 13 13 10 9 2 13 15 0 2
7 9 13 13 13 9 0 2
4 9 13 0 9
3 13 15 13
8 0 9 13 13 0 16 0 2
10 13 2 16 11 9 13 9 12 9 2
12 15 1 9 13 13 9 9 9 3 13 9 2
3 15 13 9
7 9 13 13 9 13 9 2
3 3 9 13
31 3 13 13 2 16 11 13 10 9 9 3 9 1 7 9 13 9 10 9 2 16 10 10 9 13 3 3 7 9 3 2
8 15 15 13 0 2 15 9 2
10 7 3 13 15 2 16 13 9 13 2
4 15 13 0 9
3 9 13 13
4 9 16 11 9
5 13 9 7 9 2
29 15 13 13 2 3 3 0 2 0 9 3 16 13 2 10 9 7 2 0 2 3 10 9 15 13 13 7 2 0
4 13 15 9 2
12 11 15 13 3 3 0 16 15 13 3 3 2
6 15 16 13 10 0 9
4 13 13 3 2
19 10 0 13 9 16 10 11 9 3 0 7 10 0 9 13 9 9 13 2
3 9 13 9
10 9 0 0 9 13 9 9 13 9 2
9 9 13 0 9 13 9 3 3 2
2 3 3
5 9 1 13 3 9
19 11 13 15 2 16 15 13 13 2 16 13 13 13 3 16 9 13 13 2
9 9 13 9 13 0 11 0 9 2
11 15 13 13 9 13 9 2 7 0 9 2
4 13 9 1 2
3 9 13 13
6 11 13 3 13 9 2
6 2 11 15 9 13 2
10 0 11 9 12 11 9 13 12 9 2
3 9 9 15
14 3 3 13 3 3 9 2 3 16 9 13 3 9 2
7 3 15 13 3 16 3 2
1 12
14 9 13 12 9 1 11 12 9 2 9 13 13 9 2
6 10 0 9 13 9 2
6 9 13 9 9 13 2
10 11 9 13 3 0 9 13 0 9 2
6 15 13 9 3 9 2
10 11 13 13 11 3 7 3 0 9 2
19 0 9 9 3 2 13 2 9 3 2 3 16 15 3 13 13 15 3 2
5 9 13 13 3 9
4 3 13 13 9
3 9 0 9
10 13 13 13 2 16 13 3 3 3 2
4 10 11 13 9
5 9 7 9 13 2
7 9 13 9 13 9 1 2
13 0 9 13 13 3 0 9 2 13 0 7 0 2
12 9 13 0 9 13 9 9 12 9 1 1 2
5 15 13 9 9 2
5 15 13 3 9 2
7 11 13 9 7 13 9 2
11 11 11 13 3 3 7 11 11 3 3 2
5 13 0 9 9 2
6 10 9 13 13 9 2
9 15 13 3 2 16 15 13 0 2
5 13 15 12 1 2
17 11 9 13 9 13 9 10 9 13 9 2 15 13 13 13 13 2
4 0 13 0 9
4 13 9 9 2
14 3 13 11 11 2 11 9 9 13 9 13 3 3 2
8 13 10 9 3 7 13 13 2
5 15 13 13 10 9
10 11 9 13 9 0 9 9 3 9 2
13 9 9 13 11 13 12 0 9 13 0 9 11 2
3 13 0 9
14 13 10 9 9 9 2 13 2 3 13 13 9 3 2
7 13 15 13 13 15 3 2
5 3 13 9 13 2
17 13 10 11 13 16 15 13 3 16 15 13 9 9 3 13 13 3
12 16 9 10 9 3 13 2 13 9 13 3 2
6 3 9 13 3 9 2
14 11 11 13 13 9 9 1 2 7 9 16 9 9 2
14 13 15 13 10 0 9 13 13 9 13 9 3 3 2
2 0 9
10 3 3 12 9 1 13 0 9 13 2
10 0 9 1 13 13 15 9 0 9 2
2 11 9
9 3 15 3 3 13 16 0 9 2
10 9 13 13 3 0 9 16 9 9 2
10 9 13 3 13 2 3 15 13 9 2
9 0 9 13 13 11 11 11 9 2
16 0 9 13 9 7 13 13 15 13 0 9 13 15 0 9 2
6 13 13 3 9 9 3
15 15 15 3 13 9 16 15 3 13 7 13 7 13 9 2
4 9 13 3 9
5 10 9 13 11 9
14 0 9 13 11 11 13 0 9 0 9 9 3 3 2
13 9 15 13 13 0 9 2 15 9 13 13 9 2
9 9 13 9 1 7 9 13 9 2
4 9 13 0 9
4 16 13 9 2
6 9 13 0 0 9 2
10 15 13 13 13 13 16 3 13 13 2
6 15 13 13 13 9 2
2 9 1
12 15 13 3 13 10 9 15 15 13 10 9 2
12 15 13 9 7 13 3 2 16 13 3 0 2
6 15 13 3 3 3 2
3 9 9 9
8 11 9 0 9 13 9 0 9
6 9 13 0 0 9 2
10 13 13 2 7 11 13 13 13 13 2
7 9 9 13 3 0 9 2
8 15 13 13 3 13 15 13 2
12 10 9 13 9 2 16 9 13 13 13 9 2
14 0 7 0 2 3 13 7 3 13 9 13 3 12 2
22 15 13 13 9 9 9 2 7 15 13 2 15 3 15 3 7 13 3 13 3 2 2
4 13 0 9 2
5 15 13 13 15 2
4 10 0 0 9
7 9 13 3 3 11 7 11
2 9 9
5 13 3 3 3 2
3 9 7 9
24 9 13 9 9 3 12 9 9 2 15 9 9 1 13 9 2 7 3 11 1 3 0 9 2
3 0 9 11
5 9 3 1 11 11
5 13 9 9 9 2
14 13 0 9 2 13 9 2 13 9 2 15 13 0 2
12 9 13 1 13 13 9 13 12 9 9 0 2
7 0 9 1 9 9 13 2
5 13 15 13 3 2
8 9 13 9 13 7 13 0 9
6 3 15 13 3 13 2
5 15 9 13 13 2
13 7 6 2 13 3 13 2 16 15 3 3 13 2
11 15 13 9 11 11 1 13 3 11 7 2
6 13 0 9 2 0 11
17 7 15 2 15 9 9 3 13 2 13 9 7 15 13 9 9 2
12 11 9 11 9 13 10 13 9 11 9 9 2
5 9 13 3 11 2
4 15 13 12 9
12 13 3 12 9 3 0 9 1 10 9 9 2
5 15 9 15 15 2
8 0 9 15 13 10 9 13 2
15 9 9 13 13 3 2 16 11 13 13 0 9 0 9 2
7 15 1 15 13 0 9 2
10 15 13 13 9 12 9 2 3 9 2
5 13 13 3 3 2
6 15 13 13 15 9 2
2 13 13
8 9 13 3 13 9 7 9 2
6 15 13 0 9 9 2
14 15 13 3 11 13 2 7 9 13 9 13 3 3 2
12 9 13 0 2 16 9 13 3 9 0 9 2
7 12 0 9 13 0 9 2
16 9 9 13 3 13 9 2 3 16 9 13 11 7 10 9 2
8 15 15 13 2 16 13 9 2
14 9 9 13 9 2 15 13 9 9 7 13 3 3 2
9 0 0 9 13 3 13 13 3 2
7 11 9 13 3 13 3 2
12 11 13 11 3 9 12 7 3 0 9 12 2
8 11 9 11 13 13 10 9 2
11 9 0 9 9 9 9 13 13 0 9 2
15 3 15 11 1 10 9 13 2 16 9 2 7 15 11 2
3 9 13 13
16 3 13 0 9 7 9 2 3 0 16 15 13 13 15 13 2
13 12 13 3 11 2 12 15 15 13 13 9 13 2
15 7 15 13 13 3 0 2 16 13 13 13 11 9 1 2
21 11 9 13 11 0 9 2 7 13 9 13 15 3 2 16 9 3 13 13 0 2
2 9 9
6 13 3 7 13 3 2
3 9 13 13
5 9 13 3 13 9
15 13 3 3 13 13 3 10 9 2 15 10 9 15 13 2
9 0 9 13 9 13 9 12 9 2
2 13 9
11 0 9 9 12 9 13 13 9 0 9 2
5 15 13 3 15 2
4 0 9 13 2
7 13 15 13 13 3 16 13
7 7 3 15 13 15 13 2
20 9 13 3 9 2 10 9 2 9 7 9 13 9 2 13 9 7 13 9 2
17 9 9 9 13 9 11 13 9 2 15 15 13 11 13 0 9 2
14 9 13 9 2 3 3 0 2 16 9 9 13 13 2
7 15 13 9 7 9 9 2
6 9 9 7 9 3 2
5 3 13 9 9 2
7 9 7 9 7 3 9 2
6 9 13 3 0 9 2
10 11 9 13 3 13 3 9 7 9 9
3 15 13 9
7 9 13 3 13 3 0 2
14 9 9 1 13 9 2 16 9 13 0 7 0 9 2
10 9 13 13 9 2 3 2 15 13 2
4 3 13 0 9
4 13 13 0 2
10 3 0 9 16 9 13 10 9 13 2
6 3 13 10 12 9 2
3 6 13 2
10 13 15 9 2 13 15 0 13 15 2
10 13 0 2 16 9 13 13 9 13 2
11 9 13 10 9 9 13 10 9 3 13 9
14 10 9 13 13 3 2 16 13 13 9 10 0 9 2
19 0 13 9 12 9 0 9 7 3 13 11 3 13 13 9 13 11 3 2
13 9 13 13 0 2 7 9 1 15 13 13 9 2
14 16 3 0 9 9 9 9 13 3 0 9 13 9 2
14 9 9 13 9 2 10 9 13 3 13 13 10 9 2
7 9 9 13 0 0 13 2
8 11 9 13 9 1 9 9 2
8 13 12 13 0 0 0 9 2
5 3 9 9 13 2
6 3 10 9 13 13 2
8 13 3 3 12 9 9 9 2
7 15 13 16 15 13 13 2
13 3 15 15 3 13 2 13 13 9 3 16 13 2
2 7 16
11 3 15 13 13 0 2 16 13 13 9 2
6 15 13 13 9 3 2
11 11 9 13 9 3 16 13 13 10 9 2
5 13 0 13 0 2
9 9 1 13 9 0 9 7 9 2
11 0 9 9 1 2 9 7 9 13 9 2
6 13 15 15 9 13 2
4 3 11 13 2
6 13 3 3 13 13 2
9 9 13 3 10 9 1 13 3 2
8 11 13 9 2 13 3 13 2
4 11 13 9 2
10 11 13 15 3 13 9 1 3 9 9
5 15 13 3 3 2
8 13 9 13 9 9 1 11 9
14 10 9 13 10 9 13 9 2 16 13 3 3 9 2
11 9 7 9 13 0 9 13 0 9 9 2
11 9 9 15 13 9 16 15 13 3 9 9
12 13 13 3 16 0 13 13 13 7 13 9 2
7 13 15 3 13 3 9 2
7 13 0 9 13 9 9 2
6 3 9 13 9 0 2
2 13 9
16 15 13 2 16 11 13 3 0 7 16 10 9 13 13 9 2
7 3 15 13 0 10 9 2
8 11 1 9 13 9 0 9 2
9 11 13 0 7 3 0 11 11 2
6 9 13 13 1 9 2
17 15 3 13 2 2 3 15 10 9 13 2 15 13 3 9 2 2
7 11 13 0 8 7 9 2
6 15 13 3 13 9 2
11 15 13 11 1 7 13 13 15 9 9 2
2 0 9
10 9 1 10 9 13 13 13 10 9 2
8 13 15 10 9 3 9 13 2
19 16 13 13 9 13 7 13 0 9 9 0 11 9 2 13 3 0 9 2
19 8 8 13 13 11 11 13 9 9 2 13 0 9 13 3 13 3 3 2
4 15 13 0 2
7 13 13 13 3 13 9 2
11 0 9 13 1 15 3 0 0 2 15 2
5 15 13 0 9 2
16 15 13 0 7 0 2 0 2 12 9 2 15 3 13 13 2
10 13 9 3 9 7 13 0 9 15 2
5 9 13 9 11 2
9 9 2 13 13 0 9 9 2 2
2 13 9
11 9 13 11 9 0 9 3 9 11 9 2
13 11 13 9 7 9 11 9 13 13 13 9 9 2
14 0 2 15 11 13 9 13 2 16 9 1 13 9 2
5 11 13 15 13 2
4 9 13 9 2
10 3 15 3 3 13 2 16 13 9 2
19 7 10 0 13 9 13 3 9 2 15 13 13 9 12 9 0 9 11 2
5 9 13 13 3 9
8 11 12 9 13 12 13 9 2
7 11 9 13 3 13 3 2
2 9 13
3 2 3 2
8 13 0 16 15 13 3 9 2
7 13 15 9 13 13 13 2
3 13 13 2
3 11 13 2
4 9 9 11 11
4 9 13 0 9
8 0 9 9 13 3 3 9 2
8 0 9 9 13 0 9 9 2
5 10 10 12 11 9
10 9 1 7 1 13 9 2 7 9 2
7 9 2 16 13 9 9 2
3 13 3 2
4 15 13 9 1
7 7 11 15 13 13 9 2
20 16 15 13 3 3 2 13 15 9 9 2 11 1 3 16 15 13 11 3 2
5 9 13 9 9 13
2 9 9
11 0 12 9 9 13 13 0 3 13 9 2
20 9 3 15 13 0 7 0 13 9 3 2 7 3 15 1 0 9 13 9 1
3 9 13 13
7 0 9 9 13 15 13 2
3 15 13 9
9 13 13 9 7 13 13 13 15 2
8 13 3 3 0 9 10 9 2
12 11 13 13 11 11 9 11 0 11 0 9 2
6 0 9 13 3 9 2
3 9 13 9
4 15 13 15 2
5 13 15 10 9 2
5 3 9 9 13 2
10 9 13 3 9 3 9 9 7 9 2
6 15 13 13 13 15 2
12 13 3 13 2 13 10 0 9 1 13 9 2
5 9 13 9 12 2
9 11 13 16 11 13 9 0 9 2
11 0 9 13 15 1 15 13 9 0 9 2
7 2 13 16 9 13 3 2
4 13 0 9 2
9 11 2 9 10 9 13 0 9 2
17 16 3 13 9 10 9 13 3 13 2 13 0 9 3 13 12 2
12 9 9 13 12 9 9 12 1 0 9 1 2
9 15 13 10 0 9 15 3 13 2
6 9 13 13 9 3 2
9 3 9 13 3 3 9 7 9 2
3 15 13 2
20 9 13 9 9 3 13 3 10 9 13 15 7 10 9 9 3 16 11 1 2
17 15 13 12 3 0 7 0 9 2 7 13 3 0 2 9 13 2
11 9 13 0 7 0 2 7 3 0 0 2
15 15 3 13 13 9 2 3 2 9 7 0 13 13 2 2
12 11 13 0 9 13 3 13 2 0 7 0 2
6 3 3 15 9 13 2
21 0 9 15 13 11 9 13 0 0 3 13 1 9 9 7 9 3 15 2 16 2
7 13 3 2 9 13 9 9
12 9 9 13 2 16 9 9 13 12 0 9 2
4 9 15 13 3
8 6 2 10 9 15 13 9 2
6 10 9 13 0 9 2
10 11 13 3 9 2 16 15 13 9 2
16 13 13 9 1 0 9 7 0 13 2 3 3 16 9 13 2
16 16 15 13 9 13 2 13 1 15 0 2 16 15 13 13 2
3 9 13 2
4 15 15 13 2
6 9 13 12 9 9 2
5 13 9 15 1 2
3 9 13 13
10 15 1 9 13 13 3 11 13 9 2
9 15 13 13 0 2 7 0 3 2
3 9 9 2
6 3 13 13 3 15 2
3 9 13 13
8 13 3 9 15 3 13 9 2
11 9 7 3 3 12 9 13 9 1 0 2
12 11 9 12 9 9 8 7 9 9 13 13 2
14 9 3 9 13 15 2 16 0 9 1 9 13 0 2
15 9 13 9 7 16 15 13 13 13 0 9 2 13 9 2
8 3 9 9 13 13 0 9 2
11 11 9 13 9 11 2 11 7 12 9 2
4 13 3 3 2
5 9 13 9 9 2
26 13 3 15 2 16 16 9 13 9 9 9 7 10 10 0 9 13 9 2 3 0 13 13 9 9 2
8 15 13 3 13 13 9 9 2
15 9 9 0 9 13 2 16 13 0 9 13 9 0 9 2
3 9 13 0
10 9 13 13 9 3 13 10 12 9 2
2 9 13
5 3 3 13 0 9
9 9 13 0 9 7 11 7 11 2
7 9 13 3 3 3 9 2
9 0 9 11 11 13 9 9 9 2
2 11 9
4 15 13 9 2
4 3 15 13 2
11 11 13 2 16 11 13 0 9 3 9 2
3 13 0 2
13 15 13 3 12 9 9 7 3 12 9 3 9 2
8 9 9 9 13 10 9 9 2
5 15 13 9 3 2
19 9 13 9 2 1 10 9 2 15 15 13 3 3 2 0 2 0 9 2
9 13 13 13 0 9 3 9 1 2
4 13 15 3 3
8 9 13 0 13 9 13 9 2
8 11 3 13 15 13 3 12 2
5 16 15 13 13 9
6 9 11 13 12 9 2
9 13 9 2 9 7 9 0 9 2
2 3 3
4 9 13 3 9
8 3 11 0 9 9 13 13 2
5 3 15 3 13 2
8 11 13 3 12 7 11 12 2
5 15 13 12 9 9
8 9 9 13 13 13 9 9 2
4 3 15 13 2
6 13 13 13 0 9 9
5 13 15 13 9 2
12 9 9 1 9 13 3 3 3 0 16 9 2
5 15 1 3 15 2
25 7 3 3 13 3 3 3 13 10 0 2 10 2 9 9 7 2 10 9 3 13 3 3 3 7
6 9 9 13 13 3 11
9 10 9 2 15 9 13 13 9 3
4 13 11 13 9
2 15 1
6 9 13 9 13 9 2
3 9 3 2
7 9 13 3 13 0 9 2
5 9 13 3 9 2
5 13 15 13 9 2
9 3 9 12 9 13 11 3 12 2
14 15 3 13 2 7 9 9 13 13 13 3 0 9 2
11 15 13 0 9 13 2 3 15 13 9 2
14 15 0 9 3 13 10 9 16 13 3 11 7 11 2
3 15 13 2
24 2 11 2 13 15 0 2 16 11 13 13 15 9 2 12 2 7 13 15 9 2 12 2 2
7 9 1 13 15 13 3 2
12 0 9 2 15 13 2 13 16 9 13 9 2
8 3 13 9 13 2 3 9 2
6 9 13 9 9 13 2
5 13 15 13 13 2
13 9 9 13 3 13 12 9 9 13 10 13 9 2
22 3 16 16 13 0 9 13 3 3 3 12 9 3 3 13 8 7 9 10 11 9 2
7 9 13 3 9 0 15 1
6 2 15 13 9 13 2
7 11 13 15 7 13 9 2
9 13 9 7 9 9 0 9 9 2
4 0 9 13 11
9 16 13 13 2 3 15 13 9 2
4 9 13 13 2
17 11 13 13 2 16 15 1 11 13 0 2 7 15 2 11 13 2
11 9 13 2 3 3 13 9 9 13 9 2
4 15 13 3 11
11 9 13 3 9 9 13 9 0 12 1 2
12 9 2 15 13 3 9 2 13 13 9 9 2
2 6 2
9 13 9 1 7 13 1 0 9 2
2 3 9
8 9 1 13 13 10 9 9 2
9 0 9 13 9 7 3 0 9 2
11 1 15 9 13 13 15 0 13 9 9 2
14 16 9 13 0 9 2 9 13 3 13 12 9 9 2
5 9 13 13 3 2
11 10 9 2 15 13 9 9 2 15 13 2
10 13 13 15 3 3 13 3 11 9 2
3 0 9 11
6 11 13 9 9 11 2
6 9 15 13 12 9 2
6 3 15 13 15 13 2
3 9 13 0
5 15 13 0 9 2
12 3 10 10 9 13 13 13 13 3 9 1 2
4 13 13 3 2
4 13 9 9 9
8 9 13 13 9 9 11 9 2
13 13 13 15 10 9 2 11 13 13 16 9 13 2
27 15 13 9 7 9 13 9 9 2 9 9 7 9 7 13 9 9 7 9 2 9 9 2 9 7 9 2
3 9 13 13
5 3 0 9 13 13
2 10 9
6 15 13 3 13 13 2
6 2 3 3 15 13 2
10 15 13 13 2 13 10 10 9 0 2
9 15 13 9 9 2 9 13 13 2
4 2 15 3 2
11 9 13 13 9 12 13 9 11 9 1 2
6 9 13 11 13 0 9
15 7 13 3 9 2 3 13 0 2 16 9 13 3 3 2
5 9 13 9 1 2
7 0 9 13 13 3 9 2
6 0 9 13 15 3 2
12 16 13 13 9 0 9 2 13 13 15 3 2
12 3 15 13 13 13 2 16 9 13 15 13 2
5 9 13 13 0 2
8 9 9 13 2 9 13 9 2
3 13 12 9
12 9 1 13 13 3 0 9 9 2 7 9 2
2 3 9
5 3 15 15 13 2
19 9 13 9 9 2 13 9 2 13 9 2 13 2 13 2 13 7 13 2
15 9 15 13 9 11 2 9 9 2 7 15 15 13 0 2
2 9 9
9 11 13 3 13 0 1 13 9 2
8 15 13 3 12 11 0 11 2
7 6 7 15 13 3 0 2
8 13 3 0 10 0 9 13 2
7 11 13 9 9 1 11 2
26 13 10 9 13 2 16 9 2 16 9 13 0 2 3 0 9 9 13 13 9 9 7 10 0 9 2
8 13 13 3 16 13 13 9 2
3 9 11 9
6 9 13 9 9 1 2
8 13 3 7 15 13 0 9 2
11 3 9 13 13 9 3 12 9 9 13 2
10 7 3 2 13 9 16 13 3 13 2
3 3 13 3
4 15 13 0 9
6 15 13 3 1 9 2
13 3 3 12 12 9 9 13 11 9 11 9 9 2
5 10 9 13 0 2
5 11 3 3 9 2
12 11 9 9 13 11 9 9 13 10 9 11 2
6 13 15 3 10 9 2
8 13 9 2 15 13 3 13 2
4 13 2 13 9
9 3 11 13 0 9 2 3 0 2
5 3 13 10 9 2
6 15 13 15 9 3 2
2 13 13
16 13 15 13 3 9 12 0 2 15 15 9 13 13 9 11 2
17 0 13 13 3 0 15 2 7 13 3 2 15 15 13 10 9 2
3 15 13 2
5 13 3 9 9 2
13 12 9 9 2 9 13 0 9 2 3 13 9 2
8 9 13 3 2 15 13 3 2
14 12 9 9 13 3 0 7 0 9 13 9 12 9 2
5 11 3 13 9 2
23 0 9 13 3 15 2 16 9 13 13 0 9 3 0 9 1 2 7 9 13 3 3 2
5 15 13 0 11 2
4 2 13 13 2
11 13 3 9 0 9 9 7 3 9 3 2
9 9 13 3 0 9 2 3 3 11
26 7 3 10 3 0 0 9 7 15 13 3 13 3 15 16 13 3 16 13 16 13 13 9 7 15 2
2 10 9
2 10 9
7 11 13 3 13 3 9 2
14 13 0 9 13 2 15 11 7 11 13 13 13 9 2
4 13 13 13 2
7 15 15 9 13 13 13 2
17 3 3 13 9 9 12 9 0 9 2 3 3 9 9 9 13 2
6 10 9 13 3 15 2
2 13 9
13 15 13 10 9 2 15 9 9 9 9 13 13 2
2 9 9
6 9 15 13 3 3 2
8 9 9 13 11 7 9 11 2
4 3 9 0 2
4 15 13 9 2
11 13 11 0 9 12 9 9 1 7 1 2
8 13 3 13 0 13 16 9 2
2 9 9
3 9 9 13
13 3 3 13 2 16 9 7 9 13 13 3 9 2
17 15 13 13 12 9 15 13 9 2 3 16 15 13 3 0 9 2
17 10 9 0 9 13 13 15 2 16 11 9 9 13 3 9 0 2
8 15 13 13 3 6 0 9 2
7 13 0 7 3 13 0 9
5 15 13 9 3 2
15 11 11 11 13 9 3 12 9 0 2 13 9 13 9 2
2 0 9
25 11 13 9 1 0 0 7 0 0 2 2 13 15 3 3 2 16 13 3 13 3 10 9 13 2
8 3 3 15 13 2 13 15 2
9 9 13 0 9 13 15 13 9 2
3 13 9 2
10 9 13 9 9 9 13 3 10 9 2
4 15 13 13 13
20 7 6 16 15 13 9 9 9 7 13 7 13 9 2 15 13 0 0 9 2
19 12 9 13 8 8 2 8 8 2 15 13 0 9 9 3 9 9 1 2
11 13 9 13 2 16 9 13 15 3 13 2
15 16 9 9 13 3 9 0 9 2 0 9 9 13 13 2
3 12 9 2
6 15 13 3 0 9 2
3 13 9 2
17 9 13 0 2 10 9 13 13 9 2 3 0 9 3 13 13 2
4 11 11 13 2
13 13 13 9 9 7 13 2 16 13 3 13 13 2
2 0 9
5 9 13 3 3 2
12 13 15 15 3 13 16 15 13 10 9 9 2
7 13 10 9 3 0 13 2
3 2 13 2
4 9 13 0 2
14 3 0 15 13 13 10 0 9 2 15 15 13 3 2
2 10 0
8 13 15 15 13 2 9 13 2
14 0 13 2 16 13 11 9 13 3 0 9 16 11 2
5 13 3 13 13 2
2 0 11
3 9 13 9
17 9 13 0 3 2 3 9 13 3 9 3 9 3 13 9 9 2
3 13 9 2
10 11 13 7 13 13 9 9 13 9 2
3 15 13 11
3 13 9 2
2 3 3
11 9 9 9 13 3 9 2 0 0 9 2
7 11 11 3 13 0 9 2
6 9 13 13 3 9 2
6 9 9 13 9 3 2
19 10 9 2 12 2 13 3 12 9 9 2 15 13 9 2 16 13 9 2
9 13 13 2 16 13 9 13 0 2
2 3 9
11 10 9 15 13 2 16 11 13 15 9 2
13 9 9 9 13 2 16 9 13 13 1 9 9 2
6 0 9 13 0 9 2
9 15 3 13 13 7 3 3 13 2
4 13 11 9 1
4 13 0 13 2
10 13 9 13 0 7 9 1 13 9 2
10 16 9 13 3 2 9 13 3 13 2
3 9 13 9
7 9 13 13 10 9 1 2
9 15 13 15 13 13 16 13 0 2
9 13 15 2 7 13 13 13 3 2
4 15 13 13 9
7 0 9 13 0 12 9 2
2 10 9
6 11 13 15 3 9 2
6 9 13 9 9 9 2
6 15 13 0 9 9 2
12 0 9 9 13 9 9 13 7 15 1 9 2
13 13 15 3 13 13 10 9 2 15 13 13 9 2
6 9 9 13 3 0 2
7 0 9 13 3 9 9 2
6 9 9 9 13 3 2
17 9 3 13 7 13 3 3 3 3 10 9 7 9 3 3 0 9
14 16 15 13 2 16 15 13 3 2 15 13 3 3 2
20 13 13 3 3 13 0 2 3 15 13 13 12 9 3 16 13 9 0 9 2
20 3 13 12 9 15 13 0 9 3 16 15 7 15 13 3 3 13 15 3 2
14 16 15 13 9 2 15 15 13 2 9 13 13 3 2
4 13 0 9 2
7 15 13 15 9 9 9 2
16 9 3 13 2 12 2 3 12 9 2 7 15 0 7 13 2
3 15 13 2
3 9 9 11
21 13 9 13 9 2 13 9 2 9 2 9 2 9 2 13 9 2 9 7 9 2
10 15 13 0 13 2 7 13 13 15 2
6 12 9 13 9 0 2
16 3 13 3 9 15 2 7 3 8 0 9 16 3 13 7 2
7 0 0 9 13 1 9 2
8 2 11 2 3 13 11 9 2
15 11 13 13 11 13 9 0 2 7 15 13 3 9 1 2
8 11 13 9 2 7 9 13 3
4 9 13 13 13
18 11 11 13 9 13 13 12 9 7 9 15 13 13 13 9 7 9 2
5 3 13 9 9 2
9 3 15 13 13 0 2 15 13 2
12 15 13 9 13 0 9 9 13 7 9 13 2
6 13 10 9 13 9 2
9 11 9 13 13 0 9 15 1 2
10 9 13 3 9 2 15 9 13 9 2
6 15 13 13 9 0 2
15 3 9 13 9 1 13 2 3 9 13 9 13 9 1 2
2 13 13
14 9 13 3 0 2 9 2 9 7 9 9 7 9 2
2 13 3
13 9 13 3 3 0 2 16 0 13 9 9 9 2
3 13 13 13
4 0 9 7 9
11 13 15 3 15 16 11 9 13 9 1 2
3 15 13 9
2 2 13
14 16 13 10 9 7 9 2 7 3 3 3 13 9 2
2 0 9
8 9 0 9 9 13 16 9 2
10 9 2 16 15 13 13 2 13 0 2
6 13 15 9 11 1 2
51 9 13 13 2 7 15 13 0 3 11 2 16 13 10 0 9 2 3 9 2 13 13 2 3 3 16 13 9 2 3 15 13 2 9 13 13 13 9 7 9 2 7 15 13 9 15 2 16 13 13 2
9 9 13 0 9 2 16 13 3 9
10 0 9 13 3 9 0 13 9 9 2
18 9 13 9 2 15 3 15 13 13 13 2 7 15 15 13 13 13 2
13 10 9 15 3 16 9 13 13 9 1 3 13 2
18 3 10 9 13 2 13 3 3 9 2 7 10 9 15 13 13 9 2
7 15 13 9 13 10 9 2
15 15 15 13 2 16 10 9 13 13 9 7 13 3 3 2
5 3 9 3 13 2
19 6 3 13 13 3 13 9 16 15 13 9 9 16 15 13 13 13 15 2
12 9 15 13 13 0 13 0 8 7 9 1 2
