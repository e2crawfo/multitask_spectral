298 17
29 15 13 16 1 15 7 10 9 1 9 7 9 0 15 15 4 3 13 2 15 4 13 10 0 9 1 10 9 2
16 15 4 3 13 1 9 1 11 1 2 9 1 10 9 2 2
60 2 15 4 4 3 13 16 10 9 0 1 10 9 3 0 1 10 11 0 13 10 9 1 0 9 1 10 9 0 2 1 10 9 0 2 10 9 7 10 9 2 2 13 10 9 0 2 13 1 12 9 2 13 1 10 9 1 9 0 2
42 12 2 9 1 10 9 0 1 10 11 1 10 11 7 10 11 1 11 2 11 2 2 1 1 10 12 9 2 2 1 10 11 2 12 2 7 10 11 2 12 2 2
38 7 3 2 3 1 10 0 9 1 11 0 2 10 9 12 2 15 13 10 9 1 10 9 13 1 10 11 2 13 1 10 9 11 11 11 1 11 2
11 10 9 1 1 10 9 13 1 10 9 2
34 15 14 13 3 10 9 2 3 16 1 10 9 15 14 13 3 10 9 1 10 9 0 2 7 15 13 1 15 15 15 15 15 13 2
48 15 15 15 13 15 13 3 16 15 4 13 1 10 9 1 10 9 1 9 7 13 10 7 10 9 2 0 7 0 9 2 1 10 9 2 3 16 10 9 13 1 10 9 2 12 9 0 2
15 10 9 2 13 1 10 9 1 10 9 2 4 13 9 2
29 1 15 2 15 13 3 16 10 9 13 3 2 1 10 9 1 10 9 1 10 9 0 1 10 9 15 15 13 2
25 13 15 10 9 1 10 9 7 1 10 9 16 10 10 9 13 1 10 11 7 10 11 13 0 2
35 3 2 1 10 3 1 0 9 15 13 16 15 15 4 13 0 7 0 2 7 16 10 9 14 13 3 10 9 1 10 9 2 7 3 2
18 0 3 2 10 9 1 9 4 3 13 1 4 13 2 13 7 13 2
33 1 4 13 1 9 10 9 0 2 10 9 0 13 9 1 9 0 1 13 10 2 9 0 2 13 1 10 9 1 10 11 0 2
18 0 2 0 2 0 2 0 1 9 2 15 13 3 3 1 10 9 2
32 7 16 3 10 11 14 13 3 10 9 0 2 0 2 1 11 2 15 14 4 3 13 10 9 1 15 13 1 10 9 0 2
13 12 9 3 3 2 15 13 10 9 1 10 9 2
4 15 13 0 2
51 1 15 2 10 9 4 13 1 9 1 13 10 9 1 10 9 1 10 9 1 9 2 2 3 16 10 9 0 2 1 10 9 13 1 10 11 0 2 1 10 9 3 1 10 9 13 1 10 9 0 2
28 10 12 9 2 10 11 0 1 10 11 11 11 4 4 13 1 11 1 10 9 11 7 10 0 9 11 9 2
21 15 15 13 1 10 10 9 13 10 9 7 10 9 1 10 9 7 1 10 9 2
21 1 10 9 2 10 9 1 11 11 13 10 9 1 9 7 1 9 1 10 11 2
7 9 1 9 2 9 2 2
12 3 3 13 0 7 1 9 1 10 9 0 2
13 3 13 1 10 9 0 1 10 9 1 10 9 2
9 10 9 1 9 13 0 1 9 2
35 1 15 2 15 13 16 10 0 9 1 11 14 13 3 1 10 0 9 0 7 2 1 3 2 14 13 3 1 10 9 1 10 0 9 2
11 3 3 1 15 13 13 3 1 1 15 2
9 15 15 13 10 9 13 11 11 2
6 12 2 10 9 0 2
9 15 13 12 9 12 1 9 0 2
32 7 10 9 0 13 10 9 0 15 10 9 0 13 1 10 9 0 15 13 1 9 1 9 13 13 10 10 9 7 3 3 2
16 10 9 15 4 13 2 7 3 1 10 9 13 1 10 11 2
26 3 16 10 11 2 11 0 1 10 9 0 2 2 13 1 9 1 2 0 9 2 1 2 13 2 2
7 10 9 13 15 10 9 2
7 15 13 10 9 1 11 2
24 16 1 10 10 9 0 2 15 15 13 10 9 2 13 10 9 2 13 10 0 9 1 9 2
20 3 1 9 14 13 15 16 0 2 7 14 13 15 3 3 9 1 10 9 2
8 0 15 13 0 1 10 9 2
35 3 2 10 11 13 1 13 10 9 1 10 9 0 1 10 9 1 10 11 2 3 16 1 10 9 1 9 0 1 10 9 1 10 9 2
18 1 10 9 1 10 9 0 2 10 9 1 10 11 0 13 3 0 2
12 10 9 0 14 4 13 16 13 7 15 13 2
33 1 9 2 10 6 9 4 13 0 7 4 13 3 3 1 12 9 13 1 10 9 1 10 9 7 1 10 9 1 10 9 0 2
12 15 14 13 10 9 1 9 1 10 9 0 2
16 7 10 9 13 16 10 11 14 13 3 10 11 7 10 11 2
27 1 11 2 15 13 10 9 16 10 9 4 3 13 3 2 16 15 15 13 7 14 13 10 9 1 13 2
14 15 13 15 10 9 1 13 10 9 13 3 1 11 2
10 15 13 0 2 15 15 13 10 15 2
36 13 1 11 11 1 10 9 1 2 10 11 1 10 11 2 10 11 11 2 2 10 12 12 9 1 10 9 0 13 0 1 10 12 9 0 2
31 3 10 0 9 13 1 10 9 1 10 9 2 15 15 13 16 10 9 1 10 9 1 9 14 13 3 3 0 16 15 2
30 13 1 10 2 11 2 1 10 11 2 11 0 15 13 3 1 10 9 1 10 9 2 0 2 0 7 3 0 2 2
11 13 10 9 2 16 15 15 13 1 3 2
13 15 13 1 10 0 9 1 10 9 2 9 0 2
4 12 9 12 2
91 10 0 9 13 1 10 9 4 13 10 9 1 10 10 9 0 2 1 10 9 0 7 0 2 1 15 13 1 13 10 9 0 2 3 1 10 9 0 7 13 10 9 1 10 10 9 13 1 10 9 1 10 9 0 1 10 9 2 13 10 11 0 1 13 10 9 1 9 0 7 1 13 10 9 1 10 9 2 1 10 11 2 1 10 9 0 1 10 11 0 2
24 15 15 13 1 9 2 2 15 13 3 3 10 9 1 9 1 10 9 1 10 9 1 11 2
11 1 10 9 2 15 14 13 3 1 3 2
62 11 11 11 11 7 11 11 11 2 12 9 0 1 10 9 0 1 11 11 2 15 4 15 13 13 9 0 1 10 9 1 11 2 10 9 0 1 10 11 0 2 3 16 15 13 10 9 15 15 4 13 1 10 9 1 11 2 1 9 1 9 2
17 1 10 9 16 15 13 10 9 2 10 11 13 15 1 10 9 2
14 10 9 0 2 11 11 7 11 11 2 4 4 13 2
6 15 4 13 10 9 2
51 10 9 12 13 3 10 9 2 11 2 2 7 16 10 9 1 9 0 4 3 13 1 9 1 10 9 2 10 9 13 1 10 9 1 10 9 1 9 4 4 13 1 10 9 1 10 9 2 9 2 2
50 3 4 3 13 1 13 3 1 12 12 12 9 2 10 9 2 15 13 0 15 15 15 13 1 13 10 9 0 2 13 16 10 9 14 13 16 10 9 0 14 13 3 3 3 10 9 1 10 9 2
27 10 9 1 0 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 8 2 2
46 15 13 1 11 2 15 15 15 13 9 1 2 9 2 15 4 13 1 15 13 1 3 16 2 9 2 2 1 15 13 1 9 1 10 9 1 9 0 2 16 10 9 4 13 9 2
38 4 3 13 1 10 9 2 10 9 1 10 9 0 13 1 11 2 3 1 11 1 10 9 2 1 11 2 1 10 11 2 1 11 7 1 10 11 2
23 9 2 3 10 9 14 13 3 10 9 0 2 3 3 10 9 1 15 15 15 4 13 2
57 7 10 9 1 9 0 13 3 2 15 13 10 3 0 9 1 10 9 2 15 13 10 15 1 10 12 9 9 2 15 13 0 1 10 9 1 10 9 2 1 10 9 2 15 13 10 9 0 7 15 4 13 1 10 9 11 2
8 15 15 13 1 2 9 2 2
54 10 0 11 15 13 1 14 13 3 1 15 13 2 1 3 16 0 9 1 10 9 2 1 13 10 9 0 1 10 9 0 1 10 9 1 10 9 0 7 1 10 9 1 10 9 7 1 13 10 9 1 10 9 2
16 11 11 1 11 14 13 3 3 1 13 10 9 3 3 0 2
19 1 3 16 10 9 13 1 13 10 9 15 13 3 7 1 9 2 0 2
9 15 13 10 11 1 10 9 0 2
9 7 15 13 2 3 2 15 13 2
34 1 15 13 10 9 1 10 9 1 10 9 0 2 15 15 13 1 13 10 9 1 10 9 1 3 13 10 9 0 1 10 11 3 2
40 1 9 1 10 9 2 10 9 12 7 12 1 10 9 0 1 10 9 0 2 9 2 13 10 9 1 9 1 9 1 9 1 9 1 10 11 7 10 9 2
29 13 2 15 2 10 9 1 10 9 7 1 10 9 3 1 10 0 9 0 13 1 13 10 9 1 10 0 9 2
29 1 4 13 10 9 1 10 9 0 2 10 12 9 1 9 4 13 10 9 1 13 1 10 9 7 1 10 9 2
24 15 13 1 10 9 16 10 9 0 3 0 2 9 2 4 4 13 1 10 9 12 1 12 2
21 15 15 13 16 15 15 13 10 9 1 15 15 4 13 10 9 1 10 9 0 2
76 3 1 13 16 2 10 11 13 1 9 0 2 2 1 10 13 1 10 9 0 1 10 9 1 10 9 0 2 15 4 13 10 9 1 10 11 1 10 11 1 9 1 10 11 2 6 13 10 11 1 10 9 1 10 9 1 10 11 1 13 10 9 7 10 9 1 10 9 1 10 9 1 10 9 0 2
41 13 10 9 1 10 9 2 13 15 13 1 10 9 1 15 15 14 13 3 15 2 13 1 10 9 0 1 10 9 7 1 10 9 15 15 13 2 13 10 9 2
49 3 2 13 15 10 9 2 2 2 3 2 10 11 13 16 10 9 13 9 1 10 9 10 12 9 2 10 9 2 7 16 15 15 4 13 15 0 2 9 1 10 9 2 15 14 3 13 3 2
33 1 10 9 2 3 3 13 2 2 1 10 9 1 11 11 7 10 9 1 10 9 1 11 11 2 10 9 4 13 1 10 11 2
25 1 9 2 10 11 0 4 4 13 1 10 11 1 12 7 12 9 1 10 9 0 1 10 9 2
18 3 2 1 10 9 1 9 2 10 9 0 13 3 16 10 9 0 2
10 15 15 15 4 13 1 10 11 2 2
28 10 9 1 10 11 2 11 11 2 13 2 1 10 9 13 1 10 11 2 10 9 0 1 10 11 0 2 2
49 10 9 0 11 11 4 13 2 10 9 0 2 1 10 9 1 10 9 2 15 4 13 16 10 9 15 4 13 1 13 10 9 1 10 9 2 0 2 0 2 7 3 0 2 1 10 9 0 2
68 13 12 9 1 10 0 9 0 1 10 11 2 11 2 2 10 0 9 15 13 1 10 9 1 10 9 0 1 10 9 0 1 10 11 0 1 10 11 0 2 9 11 11 2 1 9 1 10 9 1 10 12 9 7 10 9 1 10 12 9 0 2 10 11 7 10 11 2
9 10 9 13 0 2 10 9 0 2
16 1 10 9 2 1 10 9 7 1 10 9 16 15 15 13 2
25 15 4 1 3 13 10 9 1 10 9 1 13 7 13 10 9 0 1 10 12 9 1 10 9 2
28 1 9 2 10 11 1 10 9 7 9 1 10 9 9 1 9 2 9 2 4 13 1 11 2 1 9 12 2
17 3 13 3 1 15 13 9 7 0 9 1 10 9 0 2 5 2
23 1 1 16 10 11 0 13 15 10 9 1 10 9 1 10 9 1 10 9 1 10 9 2
7 15 14 15 15 13 3 2
42 9 11 13 15 1 13 13 10 9 0 1 10 9 2 11 13 1 10 9 2 1 9 2 1 10 9 0 1 10 11 1 9 1 10 11 2 10 11 1 10 9 2
21 16 15 13 10 9 1 13 10 9 10 9 2 15 13 10 9 3 0 1 15 2
14 10 9 1 9 1 11 13 1 10 9 1 15 13 2
34 10 9 13 1 9 1 12 9 1 10 9 1 10 9 1 10 9 1 9 15 13 10 9 0 1 12 9 1 12 9 10 9 0 2
31 15 3 15 13 10 9 1 10 9 2 3 15 15 13 16 11 12 13 10 9 1 10 0 9 15 15 13 1 10 9 2
29 10 9 7 10 9 1 10 9 1 9 11 2 3 13 2 4 13 1 11 2 9 1 11 1 10 9 1 9 2
31 3 2 16 10 9 4 13 10 9 1 10 9 1 10 9 1 13 13 11 1 10 11 2 16 15 15 15 13 13 2 2
12 15 15 13 7 10 0 9 4 13 2 11 2
51 1 10 9 9 1 10 9 0 7 0 2 10 9 1 10 0 9 1 10 9 4 13 1 8 2 16 1 10 9 7 10 9 1 9 2 10 9 0 13 10 0 9 2 7 3 10 9 7 10 9 2
45 1 10 9 1 10 9 2 15 15 13 1 10 9 16 16 10 12 9 15 14 13 3 10 9 1 12 8 9 10 12 8 9 12 4 13 10 0 9 2 12 9 4 4 13 2
11 13 1 12 2 10 9 2 11 8 2 2
19 1 10 9 2 15 10 9 13 1 10 9 0 1 10 11 14 13 3 2
27 10 9 2 3 16 0 2 13 0 2 2 15 15 4 13 3 2 15 13 9 1 15 13 10 9 2 2
8 9 0 1 9 2 9 2 2
17 10 9 13 13 1 10 9 1 13 10 9 2 1 3 0 9 2
21 1 15 2 10 9 11 2 13 1 13 1 10 9 1 9 1 12 2 13 0 2
23 7 15 14 13 3 3 16 10 9 14 4 3 4 13 2 2 4 13 10 15 1 15 2
35 1 9 11 2 13 1 15 1 11 1 10 9 2 15 13 9 11 15 4 13 9 9 10 9 13 7 10 9 13 2 1 10 9 9 2
36 10 9 4 4 13 1 11 1 13 10 0 9 1 10 9 1 11 11 2 9 2 9 7 9 1 10 9 0 2 10 12 9 12 1 11 2
33 1 10 9 1 10 9 0 2 15 13 0 7 13 10 9 1 13 1 13 1 10 9 1 10 9 1 11 7 1 10 9 0 2
52 10 11 2 9 1 11 1 9 2 13 3 0 1 11 8 7 10 9 3 0 2 1 15 2 1 9 9 1 10 9 1 9 1 10 11 1 10 9 2 7 13 10 9 2 1 10 9 16 1 10 9 2
23 12 9 3 3 2 15 13 15 13 1 10 9 1 10 9 1 10 9 2 12 9 2 2
23 10 0 9 13 10 9 1 9 2 15 15 13 1 10 11 1 10 9 1 9 1 9 2
30 13 10 9 2 11 11 11 4 13 10 9 0 1 1 13 1 10 9 13 2 13 16 10 9 0 3 4 4 13 2
23 10 9 9 2 15 15 4 13 1 10 9 13 1 11 2 10 9 1 10 9 1 11 2
58 1 10 9 1 10 9 2 10 9 1 10 9 1 10 11 2 1 9 1 10 9 1 0 9 1 10 9 2 13 3 1 9 7 9 1 9 2 13 10 9 1 10 9 2 2 9 11 2 3 10 9 1 11 4 13 2 2 2
63 10 9 2 14 13 3 3 10 3 0 1 10 9 2 15 13 3 10 3 0 2 1 10 9 2 13 7 13 2 1 9 2 3 1 13 1 9 9 1 10 9 0 2 2 13 9 10 11 11 2 0 9 1 10 9 2 13 3 0 1 10 11 2
24 9 2 9 2 9 2 15 15 13 1 10 3 0 9 1 10 9 7 9 1 9 1 9 2
46 15 4 13 16 10 9 1 10 0 9 13 10 9 0 1 10 9 1 12 9 5 7 16 10 9 3 0 13 10 9 1 12 9 5 2 15 13 3 0 1 13 10 15 1 9 2
37 11 11 11 15 15 13 13 2 10 9 1 10 11 2 2 4 13 12 9 1 9 1 13 13 1 10 9 16 15 4 13 10 9 1 10 11 2
8 1 15 13 1 10 0 9 2
35 10 9 0 1 9 13 12 12 1 9 2 1 9 1 12 9 2 7 10 9 0 0 13 10 9 1 12 9 2 1 12 12 1 9 2
7 1 3 2 15 4 13 2
28 10 9 1 12 9 1 9 13 10 0 1 10 9 4 13 1 10 3 12 9 10 9 2 4 13 10 11 2
21 10 9 1 10 11 11 13 3 2 7 3 2 16 10 9 4 13 1 10 9 2
40 0 9 2 11 11 2 11 2 15 15 4 13 2 12 2 2 16 11 11 7 11 11 2 10 12 1 11 11 7 13 1 3 1 12 1 9 1 10 9 2
38 1 10 9 2 10 9 1 10 9 1 10 9 9 14 13 3 10 0 9 1 10 9 1 10 11 2 15 13 1 3 1 3 9 9 1 10 11 2
20 15 15 13 10 9 3 0 3 1 10 9 1 10 9 2 10 2 9 2 2
4 13 10 9 2
37 16 11 14 13 16 10 9 14 4 3 13 1 3 1 12 9 2 10 9 14 13 3 10 0 1 10 11 0 2 15 10 9 4 13 12 9 2
32 9 1 9 15 2 3 2 13 1 10 0 9 10 9 1 9 1 10 9 13 3 10 9 1 10 9 1 9 1 9 0 2
22 15 13 3 1 9 2 7 1 10 9 0 2 15 13 0 1 12 9 1 10 9 2
6 15 13 10 9 0 2
24 3 2 10 9 2 1 1 10 9 7 10 9 2 4 13 10 9 1 10 9 1 10 11 2
22 15 15 13 1 10 9 13 1 10 11 11 1 13 10 9 1 10 9 1 10 9 2
27 15 15 4 13 2 2 16 15 13 10 12 9 1 13 2 15 15 13 10 3 3 2 2 4 13 11 2
27 15 13 3 13 16 15 13 3 1 0 9 1 10 9 13 1 10 9 0 2 1 13 10 7 10 9 2
22 15 13 15 16 12 9 16 15 15 13 7 16 15 15 13 12 10 10 9 1 11 2
16 1 12 9 1 12 9 7 12 9 1 12 9 9 1 9 2
29 1 12 2 4 15 13 2 15 4 13 10 9 1 11 1 4 13 10 9 0 1 10 9 1 9 1 10 9 2
13 10 9 12 2 1 11 2 1 10 9 1 11 2
23 3 2 15 13 15 13 10 9 7 15 13 10 9 2 2 4 13 10 9 1 10 11 2
12 3 13 15 10 9 1 9 1 10 9 0 2
23 10 9 0 0 2 11 2 13 3 10 9 13 10 3 1 12 9 1 10 9 1 9 2
50 15 13 10 0 9 1 9 1 11 1 10 9 9 2 10 9 1 10 9 1 11 1 10 9 2 1 3 1 3 13 1 10 9 7 10 9 3 3 10 0 9 0 15 10 9 15 13 1 0 2
39 3 13 2 12 12 1 9 9 12 2 2 10 11 4 13 10 9 12 1 9 1 10 9 0 1 12 9 1 10 9 7 10 9 1 3 1 12 9 2
33 3 10 11 4 15 13 1 10 0 9 1 10 9 0 2 15 1 10 9 0 1 10 11 1 10 9 1 10 11 2 12 2 2
49 10 11 4 13 10 0 9 1 10 11 1 9 1 10 9 2 12 9 1 10 12 9 1 12 2 1 13 10 11 1 11 12 1 12 2 9 2 12 2 1 9 9 1 10 11 11 1 11 2
16 15 4 13 10 9 1 13 2 10 9 0 1 15 13 2 2
29 1 10 9 2 10 9 1 9 0 0 14 4 3 13 10 9 1 10 9 1 10 9 1 11 1 10 9 12 2
15 3 10 9 1 9 2 15 13 2 13 7 13 10 9 2
48 9 9 2 10 9 4 13 10 9 0 1 10 9 1 10 11 0 2 11 11 2 3 16 10 12 9 0 13 1 0 1 10 9 7 15 13 1 13 10 9 0 1 10 9 1 10 9 2
15 3 1 10 9 1 10 9 2 11 11 13 10 9 0 2
14 4 15 13 1 15 13 1 10 9 1 10 9 0 2
24 15 4 3 13 1 10 9 1 10 9 2 10 11 2 11 13 12 9 1 15 13 1 12 2
23 2 15 4 13 2 1 10 9 1 10 9 1 11 2 16 10 11 13 3 10 3 0 2
17 13 10 9 1 10 0 11 11 15 13 10 9 1 9 1 9 2
35 3 1 12 9 4 1 3 4 13 2 15 12 3 2 3 1 9 13 1 10 9 0 1 10 9 1 10 9 2 11 2 1 10 9 2
20 16 2 1 10 9 2 12 0 9 4 13 1 13 1 10 9 7 3 9 2
9 1 9 9 1 9 13 1 11 11
21 1 15 2 15 13 3 1 12 9 1 9 15 4 4 13 1 13 10 9 0 2
49 10 9 4 1 3 4 13 3 1 10 9 11 11 1 10 9 1 10 9 1 9 0 1 10 9 1 10 9 0 1 10 9 7 1 10 9 2 16 15 4 13 16 15 14 4 13 1 9 2
18 1 3 2 15 4 3 13 10 9 1 10 9 1 10 9 1 9 2
18 1 10 9 2 12 9 1 12 7 12 9 13 1 11 2 11 2 2
8 15 4 3 15 13 10 9 2
39 9 1 10 9 0 0 1 10 9 13 1 10 9 1 10 9 7 10 9 13 2 13 2 10 9 9 13 3 10 9 7 10 9 1 10 9 1 9 2
26 10 9 13 10 9 1 9 2 1 10 9 13 1 12 1 12 9 1 9 2 1 10 9 1 9 2
32 11 11 11 2 15 10 9 4 13 10 9 1 9 1 11 0 2 4 13 10 9 9 2 16 10 9 13 1 15 13 2 2
34 10 9 1 10 9 3 0 13 3 0 2 7 15 15 13 1 15 1 10 9 1 10 11 2 7 13 3 10 9 1 10 9 2 2
31 2 15 13 10 9 0 1 10 9 2 7 10 9 1 10 9 13 10 9 9 2 2 13 11 11 2 9 1 11 11 2
9 15 13 10 9 1 10 0 9 2
33 10 9 2 15 13 10 9 1 0 9 1 9 7 10 9 1 10 9 0 2 4 3 13 13 10 9 1 12 9 1 12 9 2
32 1 13 10 12 9 1 10 9 1 10 11 2 10 9 0 11 11 4 13 1 13 13 10 0 9 1 10 9 7 10 9 2
12 9 9 2 10 9 13 3 1 9 1 9 2
19 1 10 0 9 2 10 9 4 13 10 3 3 0 16 10 0 9 0 2
13 3 2 15 4 13 1 13 10 0 9 1 9 2
10 15 13 10 9 2 1 13 1 2 2
23 1 11 2 10 0 9 4 3 3 13 10 9 3 1 9 1 11 11 1 13 10 9 2
28 2 10 9 1 9 2 15 13 3 10 0 9 1 15 2 15 13 12 9 1 10 9 1 9 2 13 15 2
57 13 9 9 2 1 10 9 1 10 11 2 3 10 9 0 1 10 9 1 11 11 15 15 13 1 13 11 1 10 9 1 10 9 0 2 15 13 1 10 0 9 2 2 15 15 13 3 10 10 9 2 7 15 13 1 9 2
32 13 10 9 2 11 2 13 1 10 9 1 10 12 12 12 2 12 9 1 9 1 9 1 10 9 2 7 13 1 10 9 2
39 11 11 15 4 13 9 1 10 9 0 1 11 13 16 10 10 9 1 10 9 1 10 11 13 0 7 13 1 13 10 9 1 10 9 0 13 1 11 2
13 3 13 15 3 0 1 13 3 3 2 6 2 2
48 10 9 0 1 9 0 7 10 9 1 10 9 4 13 1 10 9 2 1 10 9 2 1 13 13 10 9 0 1 12 9 1 12 1 12 12 1 9 2 1 12 9 1 9 1 9 0 2
26 12 9 4 4 13 9 2 7 15 1 10 9 1 10 9 1 10 9 1 10 0 9 1 10 9 2
36 2 15 14 15 13 3 10 9 1 9 7 10 9 2 15 14 13 3 15 15 15 13 2 2 14 4 13 1 13 10 9 13 1 11 11 2
29 11 2 12 2 13 3 1 10 9 11 2 12 2 2 15 10 9 1 11 11 2 12 2 14 4 13 1 15 2
15 7 9 9 2 11 11 14 13 3 1 10 9 1 9 2
26 1 10 9 1 9 2 1 10 9 2 15 2 16 15 15 13 13 2 13 16 15 15 13 1 15 2
63 1 16 10 9 1 9 9 11 11 13 10 9 1 10 9 13 1 10 11 1 10 9 1 10 9 0 1 11 2 10 9 0 2 12 2 12 2 9 13 1 1 10 9 13 10 9 1 9 13 1 10 9 11 11 2 1 10 12 1 9 1 3 2
14 2 3 15 15 13 2 7 15 13 16 15 15 13 2
17 10 0 9 1 10 11 1 10 9 0 15 13 10 9 1 11 2
28 2 10 9 13 1 10 9 0 3 16 0 1 9 2 15 14 13 16 13 1 10 9 1 3 1 12 9 2
9 1 12 9 1 9 1 10 9 2
32 9 0 1 11 15 13 10 3 0 9 7 10 9 1 9 0 13 1 9 0 2 10 9 1 9 7 1 10 9 3 0 2
2 3 2
40 3 15 13 3 1 10 11 2 10 9 13 3 3 1 15 13 1 13 10 9 2 10 9 13 3 0 7 15 13 3 10 0 9 2 13 7 15 3 13 2
22 11 11 2 13 10 9 15 10 9 1 9 1 9 7 9 0 14 13 3 1 13 2
23 1 10 9 1 9 2 15 13 3 0 7 3 15 14 13 3 9 1 10 9 3 13 2
25 1 10 9 2 1 9 2 10 3 0 9 2 1 10 1 9 3 2 7 10 9 1 9 0 2
22 1 10 9 1 10 9 1 9 2 15 4 13 1 10 9 0 2 10 9 1 13 2
26 3 1 10 9 15 15 13 10 9 1 10 9 2 1 15 13 13 16 15 13 9 1 13 10 9 2
18 1 3 1 12 9 2 15 4 13 1 10 9 0 1 10 10 11 2
13 6 2 13 2 15 4 13 1 13 0 7 0 3
13 6 2 15 4 13 10 9 1 10 11 9 12 2
12 9 9 0 7 15 13 10 9 2 10 9 2
18 6 2 10 9 1 10 9 1 11 15 13 1 9 1 13 3 3 2
5 6 2 1 13 2
10 9 2 10 9 1 10 9 1 9 2
12 15 13 10 9 1 10 9 1 9 1 11 11
14 15 13 3 0 1 4 13 1 10 9 1 10 9 2
21 15 13 10 9 0 2 7 15 13 1 13 10 9 1 10 9 15 13 10 9 2
22 15 3 2 15 4 13 16 15 13 1 10 9 0 7 0 2 16 13 1 10 9 2
14 7 6 15 4 13 3 3 10 9 0 1 10 9 2
25 15 13 12 9 16 15 13 10 9 0 7 15 13 10 12 9 16 15 13 1 10 9 3 0 2
9 10 9 13 3 3 0 7 13 3
18 15 13 1 13 2 13 2 13 2 13 2 9 1 10 9 0 0 2
12 9 0 1 15 4 4 13 15 1 10 11 2
14 1 12 9 2 9 7 9 2 15 13 3 10 9 2
26 1 13 16 10 9 1 9 0 7 0 13 13 1 10 15 15 13 1 10 9 1 9 1 10 9 2
19 1 3 15 13 0 2 1 10 9 7 15 13 16 15 13 3 10 9 2
17 3 2 13 10 9 15 4 3 13 1 10 9 1 10 9 13 2
24 3 10 9 1 11 15 6 15 4 13 10 9 7 10 9 0 15 14 13 3 1 1 9 2
13 7 10 9 1 10 9 13 3 3 3 2 0 2
5 7 10 9 0 2
5 13 10 9 0 2
9 0 2 7 1 3 15 13 0 2
6 3 15 13 3 0 2
7 15 4 13 1 15 13 2
14 15 13 3 13 7 10 0 9 1 11 13 3 0 2
10 15 15 13 3 10 9 1 10 9 2
15 15 13 10 9 1 9 2 7 13 10 9 1 10 9 2
35 15 15 4 13 16 15 13 10 9 1 9 16 15 13 10 9 1 10 9 2 3 13 15 2 1 1 2 15 13 0 1 2 13 2 2
6 15 4 13 10 0 9
7 15 13 1 11 1 12 2
18 15 3 13 3 3 2 7 16 15 13 15 13 3 10 9 15 13 2
8 15 13 10 9 7 10 9 2
13 15 4 3 13 1 14 13 16 10 9 5 9 2
18 15 4 13 10 9 1 9 1 10 9 2 3 13 1 10 9 0 2
22 15 4 13 1 9 11 1 13 1 11 10 9 1 9 2 10 9 13 3 10 9 2
19 15 3 4 13 12 9 1 10 9 1 9 7 15 14 4 3 4 13 2
15 15 13 3 10 9 1 10 15 15 4 13 10 0 9 2
45 15 13 9 1 11 1 12 9 2 7 1 16 15 15 4 13 1 13 10 9 13 1 10 11 0 7 1 10 9 0 2 9 2 9 0 2 9 2 2 15 4 4 15 13 2
45 15 13 3 16 15 13 10 9 0 2 12 9 10 9 15 1 3 2 7 15 13 16 10 9 14 4 3 4 13 1 10 9 2 10 9 14 4 3 3 4 13 1 10 9 2
12 10 9 13 1 9 3 1 9 16 1 9 2
32 10 9 1 10 0 7 10 0 4 13 1 3 9 1 3 1 10 9 2 15 15 14 13 3 10 12 9 3 0 1 3 2
18 10 9 11 4 13 1 10 2 12 2 9 11 11 2 11 2 8 8
28 10 9 13 3 0 2 7 10 9 14 13 3 1 10 9 1 15 1 10 9 0 2 1 9 1 9 0 2
19 10 9 13 13 1 9 1 14 3 13 10 9 1 10 9 1 10 9 2
27 10 9 15 14 13 3 2 10 9 3 2 10 9 1 9 14 13 16 10 9 2 7 10 9 13 0 2
15 10 9 0 13 16 15 13 3 1 9 7 13 10 9 2
16 10 9 13 0 1 10 9 1 10 9 7 10 9 1 9 2
20 10 9 13 3 3 0 16 1 10 0 9 7 15 13 10 9 13 10 9 2
8 10 9 1 9 13 1 9 2
6 10 9 0 13 0 2
11 9 11 13 10 0 9 15 15 13 3 2
10 9 1 9 1 9 2 9 3 0 2
15 7 1 13 16 3 10 9 14 13 10 9 1 10 9 2
5 6 3 1 15 2
25 10 9 13 3 0 2 9 9 2 9 7 9 1 9 2 7 13 0 1 10 9 7 10 9 2
31 10 9 1 10 9 1 10 9 15 13 10 9 1 10 9 1 10 0 9 0 3 1 13 10 9 7 10 9 1 9 2
22 15 4 13 1 10 9 12 9 1 10 9 2 10 9 7 10 9 2 1 9 2 2
22 15 4 13 9 1 12 9 9 13 10 9 1 0 2 9 7 9 13 1 10 9 2
6 15 3 13 10 9 2
15 1 1 2 16 15 13 0 13 10 9 15 13 3 0 2
20 1 1 10 9 13 0 7 3 0 2 10 9 0 7 10 0 9 3 0 2
30 0 9 1 9 1 13 1 10 9 2 1 12 9 2 9 1 10 11 13 10 9 0 15 15 13 3 1 10 9 2
24 1 13 10 9 2 10 9 1 10 9 14 13 3 0 2 7 0 2 15 13 3 3 0 2
60 1 10 12 9 2 15 13 9 1 10 9 1 9 7 15 4 4 16 16 10 9 13 1 13 1 10 0 7 0 9 10 9 9 1 10 3 0 9 7 1 0 9 3 0 7 3 9 7 3 1 10 9 10 9 6 10 3 3 0 2
17 1 13 15 13 16 15 13 9 0 2 7 15 14 13 3 3 2
11 9 3 0 7 15 13 3 1 10 9 2
11 9 2 10 9 0 15 3 13 1 9 2
6 16 15 15 15 13 2
19 15 13 1 3 16 15 4 3 13 1 10 9 3 0 7 3 0 2 2
26 16 15 13 1 9 0 2 1 10 9 2 7 1 9 0 1 15 2 15 13 1 11 11 11 11 2
23 16 15 13 10 9 1 3 13 16 10 9 13 0 15 13 9 1 10 9 1 10 9 2
13 16 15 13 13 2 10 9 2 14 13 3 3 2
12 10 9 13 0 7 1 10 9 1 10 9 2
17 9 1 9 10 3 0 7 3 16 1 10 0 9 15 4 15 13
13 3 0 2 15 15 13 10 9 0 7 3 0 5
22 10 9 0 2 0 7 3 0 2 10 9 0 2 10 9 0 1 10 9 1 9 2
31 13 2 15 13 16 10 9 4 13 10 3 16 11 13 10 9 15 15 13 2 15 15 13 7 3 10 9 15 15 13 2
5 15 13 3 0 2
15 15 4 13 2 13 1 10 0 9 16 10 9 4 13 2
34 15 4 13 9 1 13 13 10 9 1 10 9 1 9 0 7 0 2 7 2 11 11 2 4 2 1 10 12 9 13 1 10 9 2
12 15 14 4 15 13 1 10 9 1 10 11 2
14 3 1 12 9 12 9 1 3 0 12 9 12 9 2
24 1 13 1 10 9 10 9 0 1 10 9 2 15 4 13 9 1 15 7 10 9 13 0 2
14 3 0 9 10 9 13 3 0 7 0 0 9 9 9
5 10 9 12 9 2
11 15 13 10 9 1 13 10 2 9 2 2
