5241 17
15 10 9 13 9 9 9 7 9 13 1 15 1 9 9 2
13 9 9 13 1 10 9 7 13 1 15 9 0 2
25 10 9 13 7 3 7 3 16 13 10 9 13 12 1 10 9 7 1 10 9 1 9 10 9 2
24 9 7 9 13 1 9 10 9 2 1 9 15 1 10 9 2 1 13 1 10 9 10 0 2
24 16 13 10 9 13 2 13 10 9 14 9 10 9 2 13 7 13 14 9 15 1 10 9 2
6 15 13 14 9 15 2
9 3 10 9 3 13 14 10 9 2
22 1 10 9 16 1 9 10 9 16 1 9 10 9 13 1 9 10 9 14 9 11 2
22 11 11 2 9 11 2 13 1 9 15 9 7 13 1 10 9 3 13 1 10 9 2
16 1 10 9 13 9 2 1 10 9 13 13 14 9 10 9 2
6 9 15 1 9 12 2
15 9 1 10 9 2 9 1 10 9 2 9 1 11 11 2
26 4 13 14 10 9 1 9 10 9 11 7 3 1 9 7 9 13 9 15 14 11 11 1 10 9 2
12 3 13 14 10 9 2 7 10 9 13 9 2
5 13 9 10 9 2
5 13 9 10 9 2
6 2 13 9 7 3 2
17 3 9 13 3 1 10 9 2 13 9 11 1 9 9 10 9 2
6 9 3 13 13 15 2
35 3 10 9 16 13 1 9 2 3 9 1 10 9 10 15 2 16 1 9 9 10 9 13 9 3 13 1 9 3 1 10 9 10 0 2
36 9 2 10 9 2 1 10 9 2 13 2 9 13 3 1 9 12 1 10 9 1 11 2 0 1 9 15 14 9 10 9 2 11 11 11 2
4 9 3 13 2
28 9 9 0 2 1 9 9 9 10 9 2 3 2 9 11 11 2 13 1 9 7 1 9 0 1 10 9 2
35 1 10 9 1 11 13 9 2 1 16 9 13 16 13 1 9 0 1 9 2 11 2 2 13 9 9 0 2 16 13 13 1 10 9 2
54 11 11 2 16 13 3 1 9 9 9 10 9 10 0 1 11 2 13 16 10 9 13 1 9 15 7 16 1 9 11 11 13 14 15 10 9 16 0 9 16 9 0 13 13 1 9 9 0 1 10 9 10 0 2
34 10 9 13 3 9 2 11 0 7 9 9 0 1 10 9 10 0 2 16 13 1 9 10 9 2 16 0 9 1 9 9 1 15 2
10 15 13 13 1 10 9 1 9 15 2
39 9 13 2 9 13 1 9 9 7 0 13 1 9 15 2 12 13 2 1 9 0 2 7 3 13 12 9 11 7 9 12 1 9 10 9 1 10 9 2
20 12 9 11 13 1 9 0 1 9 0 16 13 1 9 10 9 1 9 11 2
10 15 13 1 9 10 13 11 1 11 2
24 1 9 0 16 13 1 10 9 3 7 3 13 11 11 11 11 2 9 12 2 9 9 9 2
26 12 13 1 9 0 7 12 13 2 1 9 0 2 12 1 15 1 9 9 0 2 9 9 7 9 2
21 10 9 13 1 9 2 1 15 9 0 1 9 12 7 12 7 12 9 1 9 2
15 9 9 11 1 9 9 13 13 1 15 9 13 10 9 2
17 9 0 1 9 9 13 16 12 9 13 7 12 13 1 9 15 2
20 10 9 16 13 3 1 10 9 9 9 7 1 9 0 1 10 9 13 3 2
14 9 0 0 13 16 10 9 13 1 10 9 10 0 2
27 10 9 13 3 1 16 13 9 9 15 14 9 0 1 11 2 16 13 0 1 9 10 9 1 9 11 2
11 9 16 13 13 1 9 9 1 10 9 2
16 9 0 13 16 10 9 13 1 10 9 9 3 1 9 11 2
21 12 9 13 14 9 11 1 9 7 1 9 9 7 13 9 7 9 1 9 9 2
11 15 13 14 9 9 9 11 1 9 15 2
25 9 0 13 16 9 10 9 13 3 1 9 9 9 2 16 3 13 12 9 2 1 15 12 3 2
5 1 10 9 9 2
33 3 13 16 10 9 13 1 10 10 9 10 0 1 9 11 7 3 1 9 10 9 11 2 9 11 2 9 11 7 10 9 11 2
12 3 13 12 9 9 1 9 14 11 1 11 2
9 10 9 13 2 7 3 13 9 2
14 10 9 10 0 13 1 9 1 9 9 1 9 9 2
22 11 11 11 2 16 13 1 9 9 1 10 9 2 13 1 9 9 7 9 15 13 2
15 1 9 10 9 11 13 9 14 11 9 11 2 9 12 2
29 3 13 1 9 9 0 1 9 9 11 11 2 9 12 2 16 13 1 9 0 7 13 1 9 9 2 10 9 2
46 1 9 9 10 9 1 11 13 14 9 9 15 14 11 11 11 11 11 2 9 12 2 9 1 9 9 2 0 7 9 1 12 9 2 16 13 0 3 1 9 15 16 1 9 11 2
11 9 0 13 16 11 13 1 9 14 9 2
12 9 0 16 13 1 10 9 13 14 9 15 2
17 1 10 9 13 1 9 11 9 0 1 9 10 9 1 9 11 2
28 3 13 11 14 10 9 1 10 9 10 9 10 0 2 16 13 1 9 0 1 9 9 11 7 1 9 0 2
25 9 0 13 16 1 9 10 9 13 1 9 11 12 9 0 1 9 11 2 13 1 9 10 9 2
36 1 9 11 1 9 9 9 13 12 9 9 1 9 9 0 9 11 11 2 9 12 2 16 13 1 9 0 1 9 10 13 11 11 1 11 2
38 9 0 13 16 1 9 11 13 9 9 1 9 9 10 9 1 9 9 10 9 1 9 9 2 7 15 13 1 13 7 1 13 1 9 7 1 9 2
28 1 9 1 9 9 1 9 0 1 9 2 13 1 9 11 0 9 1 9 15 2 7 15 13 1 10 9 2
30 9 10 9 11 11 13 3 9 0 1 9 11 7 13 9 1 10 9 3 2 16 13 15 10 9 10 12 1 9 2
19 11 13 1 9 11 1 10 9 1 9 15 3 1 9 2 9 1 13 2
28 1 9 10 9 13 10 9 9 1 9 9 10 9 7 1 9 11 1 10 9 2 7 13 1 9 2 11 2
25 3 13 10 9 10 0 1 9 11 7 15 13 3 1 9 10 9 1 9 10 9 7 1 11 2
11 9 0 13 1 12 9 2 3 1 11 2
28 1 9 15 2 13 9 1 11 1 9 0 1 1 9 10 9 10 0 2 16 12 9 9 13 9 1 9 2
17 9 0 13 14 16 13 1 10 9 1 10 9 10 0 1 9 2
8 9 11 13 1 12 9 3 2
14 10 9 10 0 13 16 9 11 13 13 1 10 9 2
12 3 13 12 9 9 1 9 14 11 1 11 2
11 10 9 13 2 7 3 13 1 10 9 2
22 1 10 9 13 16 1 10 9 13 3 7 3 1 10 9 9 0 1 9 1 9 2
26 9 0 13 16 1 9 9 1 13 9 1 9 9 13 9 0 2 16 13 13 9 1 12 10 9 2
14 10 9 13 1 9 15 7 13 14 15 1 9 0 2
14 10 9 13 1 9 10 13 11 9 2 9 1 11 2
21 1 9 9 3 1 11 13 9 0 1 9 9 9 0 2 16 13 1 9 9 2
41 9 0 13 16 9 2 16 13 1 9 0 1 9 11 1 11 2 13 1 9 9 9 14 9 13 14 9 0 2 1 15 3 14 9 9 15 14 13 11 11 2
23 9 0 13 16 1 9 14 9 1 10 9 2 13 16 10 9 3 13 1 2 9 9 2
28 9 14 11 13 3 9 9 1 9 9 2 16 13 1 9 11 1 9 9 0 2 1 9 11 16 1 11 2
16 9 10 9 13 1 9 9 14 11 7 13 1 9 11 0 2
15 9 11 13 16 10 9 13 1 9 7 3 13 1 9 2
22 15 10 9 12 1 10 9 10 0 2 16 9 14 11 13 1 9 0 1 10 9 2
15 1 9 9 0 2 13 7 13 10 9 13 1 9 0 2
24 12 9 1 9 9 9 13 3 2 9 15 1 9 0 2 1 9 14 9 3 13 9 0 2
37 10 9 13 16 9 14 11 13 9 14 9 1 9 9 9 7 13 14 15 1 9 16 0 1 12 9 1 10 9 9 9 2 13 1 9 11 2
13 10 9 13 1 9 10 9 7 1 1 3 13 2
16 12 1 15 13 1 9 9 1 9 10 13 10 0 1 11 2
58 11 11 11 11 2 9 1 9 2 9 10 9 11 2 13 1 9 15 7 9 15 13 2 11 11 11 11 2 9 12 1 11 2 9 1 10 9 1 11 13 12 1 9 15 2 12 9 0 13 1 9 0 7 13 1 9 15 2
19 9 11 13 1 9 2 2 9 14 11 13 9 14 12 9 1 13 9 2
9 9 15 13 7 0 13 1 9 2
16 12 1 15 16 13 1 10 9 13 1 1 9 10 9 2 2
34 9 0 13 3 16 1 9 11 1 11 13 9 9 12 2 11 11 2 1 9 9 1 9 15 2 7 13 1 9 10 13 1 11 2
24 9 13 16 10 9 13 1 9 1 9 0 2 16 13 1 9 9 9 10 9 1 10 9 2
17 1 11 13 16 9 9 0 3 13 9 7 16 3 13 9 0 2
20 12 9 9 13 3 1 9 9 11 1 10 9 2 16 13 1 10 9 11 2
18 9 0 13 16 12 10 9 13 2 7 3 13 10 9 7 13 9 2
15 1 9 9 0 13 3 1 10 9 1 9 11 12 9 2
15 10 9 13 1 9 1 9 10 9 7 1 10 9 11 2
22 9 9 11 1 9 10 9 13 7 1 9 7 1 12 9 16 13 1 9 10 13 2
32 1 9 10 9 1 11 13 3 12 9 1 9 9 2 1 16 13 1 9 9 0 7 9 15 1 9 9 15 1 9 9 2
63 3 16 16 15 13 0 10 2 3 16 13 1 9 14 16 13 9 15 2 13 9 15 14 11 11 1 3 16 13 1 9 9 10 9 1 11 2 2 10 9 2 2 12 2 9 0 0 1 10 9 16 13 7 13 9 1 10 9 10 0 1 11 2
17 16 16 15 2 9 15 13 3 9 0 13 9 0 1 15 9 2
58 15 13 1 10 9 10 0 2 7 0 3 10 13 2 16 7 9 10 9 3 13 7 13 10 10 9 2 1 10 9 10 0 2 1 9 10 9 14 10 9 2 7 1 9 15 1 9 13 2 7 3 1 10 9 10 0 15 2
30 15 3 13 9 0 16 13 1 10 9 3 11 4 7 3 4 13 1 9 11 2 7 1 10 4 16 13 1 15 2
63 15 9 16 13 1 9 0 2 0 3 7 0 2 3 3 11 13 14 15 2 9 0 2 2 2 7 15 9 0 1 9 10 9 10 0 1 9 0 2 1 16 13 1 9 1 9 0 0 14 10 9 2 9 2 10 9 7 9 1 9 0 2 2
48 7 3 2 1 9 13 0 16 16 4 1 3 16 0 1 15 1 9 9 7 1 10 9 10 9 2 13 11 7 9 15 13 10 9 1 9 0 2 1 9 0 2 1 9 2 9 0 2
31 10 9 13 16 7 9 13 14 10 9 2 9 16 15 0 1 10 9 2 7 1 15 4 13 0 7 0 1 9 15 2
24 9 2 9 2 11 2 10 9 7 9 15 2 9 1 10 15 13 1 10 10 3 9 0 2
5 7 13 1 15 2
3 3 3 2
46 10 9 1 10 9 2 1 2 9 9 15 2 13 3 9 0 7 3 0 2 7 15 13 1 2 9 0 2 2 16 9 15 10 0 13 3 3 16 15 1 11 2 9 7 11 2
27 2 9 7 9 2 2 13 11 14 3 16 13 2 1 16 15 13 1 15 1 9 0 7 0 14 9 2
30 1 3 13 9 11 11 14 10 9 10 0 10 15 1 9 1 12 1 9 15 2 15 13 0 1 10 9 10 0 2
31 7 16 9 15 10 0 14 11 0 3 2 7 13 16 7 0 1 9 15 2 1 10 9 10 0 16 13 1 15 9 2
29 11 13 1 9 10 9 10 0 1 10 9 10 0 14 10 9 16 1 10 9 2 16 14 15 13 2 9 2 2
40 15 13 1 10 9 2 9 7 9 2 1 13 14 10 9 16 1 10 9 10 0 10 0 14 10 9 10 0 1 10 9 10 0 14 10 9 10 0 15 2
20 3 1 15 1 9 0 1 10 9 16 1 15 9 10 9 13 1 9 15 2
29 7 9 13 2 10 9 2 9 7 9 2 13 13 1 10 9 10 0 10 0 3 14 9 10 9 1 10 9 2
36 4 13 14 15 1 9 1 9 9 7 9 1 9 10 9 1 9 11 2 1 9 1 10 9 16 13 1 9 1 9 9 2 7 1 0 2
34 13 3 9 2 3 13 10 9 10 0 10 15 16 10 9 16 13 13 9 0 2 1 2 1 9 15 13 1 15 14 10 9 2 2
35 9 1 9 2 7 7 1 9 15 2 9 7 9 2 2 1 9 15 10 0 14 9 9 2 3 13 10 9 1 9 1 2 9 2 2
45 1 10 9 10 0 10 15 0 2 16 3 9 15 7 0 13 16 13 1 11 2 7 1 9 15 13 9 9 7 9 2 16 13 13 3 1 15 2 2 7 10 9 9 15 2
23 13 16 10 9 2 10 9 0 1 10 9 10 0 10 15 2 13 1 9 15 1 9 2
24 1 9 2 15 3 13 16 13 2 13 7 13 13 14 10 9 16 13 14 10 9 10 0 2
25 15 3 13 13 1 9 9 2 7 3 16 13 15 9 0 2 0 2 3 3 9 14 9 0 2
41 1 9 15 2 7 3 1 9 9 15 10 0 7 10 0 2 15 13 16 10 9 13 0 1 10 9 2 7 3 4 13 7 13 14 15 1 9 0 2 0 2
2 3 2
24 3 1 16 10 9 0 1 10 15 3 13 4 13 14 10 9 15 2 14 10 9 10 0 2
19 15 0 2 3 2 7 3 11 3 13 16 10 9 13 4 1 9 0 2
22 1 16 13 9 0 2 3 3 13 9 16 13 9 7 13 9 9 1 9 9 15 2
17 10 9 2 7 3 2 13 1 9 10 9 13 1 9 10 9 2
34 7 16 1 9 10 9 2 1 1 10 16 13 1 10 9 1 9 11 1 9 0 2 13 1 10 9 9 0 2 7 3 3 0 2
42 7 15 3 16 13 14 11 1 10 9 10 3 2 0 10 0 2 2 10 9 13 9 16 9 15 9 7 9 2 7 9 0 3 1 9 2 1 9 7 1 9 2
17 15 13 14 9 15 1 12 9 2 10 12 0 7 10 0 0 2
15 13 1 15 9 0 0 2 9 15 10 0 13 3 2 2
33 7 3 13 12 9 10 9 2 9 14 2 9 16 9 15 9 7 9 2 13 3 7 3 16 2 9 15 10 0 13 3 2 2
11 7 3 13 13 16 1 10 9 13 9 2
11 13 13 16 9 7 9 0 13 3 0 2
28 16 10 9 10 9 10 0 7 13 9 10 9 2 7 13 1 9 7 13 9 0 0 2 13 3 9 9 2
35 13 13 16 13 1 10 9 10 15 10 9 16 0 12 9 1 9 0 2 7 1 10 15 9 0 2 3 9 15 2 3 13 14 15 2
36 13 13 16 9 0 13 12 10 9 3 0 7 0 1 10 9 2 3 1 9 15 1 9 9 0 1 9 2 9 9 2 9 7 1 0 2
50 13 13 16 9 1 9 7 9 2 3 9 9 2 0 1 10 9 2 10 9 2 10 9 2 7 3 1 10 9 0 1 9 15 2 7 16 1 15 3 3 2 10 9 13 10 0 7 10 0 2
12 1 9 12 2 11 2 1 9 15 2 13 2
60 15 7 9 15 1 10 9 7 13 7 13 14 10 9 1 15 2 3 13 7 13 1 15 10 9 0 2 1 2 15 13 13 1 10 9 10 0 14 10 9 16 9 0 2 7 3 10 9 1 15 2 0 1 9 0 7 13 1 15 2
37 7 1 16 9 1 10 15 3 13 1 9 0 3 14 10 9 2 3 10 9 16 3 16 13 13 7 13 1 9 0 13 0 1 9 0 0 2
27 3 3 9 0 1 9 15 14 11 2 1 0 1 15 14 13 0 2 3 13 9 2 10 9 1 11 2
24 11 13 16 15 13 2 1 13 9 1 9 2 2 7 15 13 3 15 4 13 15 3 3 2
43 15 9 0 0 2 3 16 2 3 1 15 9 2 2 7 3 9 10 9 10 15 2 2 1 9 2 9 3 13 0 1 15 2 7 3 16 13 13 3 13 14 15 2
13 7 3 16 13 1 11 13 3 15 4 13 3 2
31 9 13 13 14 15 13 2 7 15 13 1 16 3 16 15 4 13 3 4 1 15 3 3 2 14 15 13 1 10 9 2
63 3 2 7 3 2 15 13 1 11 3 16 16 13 1 9 15 9 0 0 2 7 15 13 1 15 9 7 9 2 7 1 16 9 9 1 11 13 3 13 14 10 9 10 15 1 9 1 10 3 16 13 2 9 9 2 1 10 15 3 1 10 9 2
31 3 13 2 1 10 13 2 3 1 9 0 1 11 7 9 11 2 11 2 7 1 9 10 9 14 10 9 7 10 9 2
63 10 9 10 0 14 9 2 10 9 13 16 7 9 10 9 2 10 9 7 10 9 10 0 4 1 9 2 3 16 13 7 3 2 0 2 13 13 1 9 10 9 1 13 1 15 15 9 9 7 9 0 2 3 0 2 2 16 13 3 9 10 9 2
22 3 2 1 11 2 7 3 4 13 2 7 3 3 1 9 15 14 10 9 2 2 2
26 3 13 16 9 15 10 0 14 10 13 1 10 9 2 1 9 1 11 2 13 1 15 3 1 3 2
29 15 13 1 1 11 7 1 11 2 1 13 1 16 13 13 9 0 2 7 13 14 9 15 1 9 0 7 0 2
31 3 2 13 2 13 9 0 1 10 9 3 9 15 3 16 3 11 13 9 0 2 16 4 13 9 14 9 7 9 0 2
37 7 16 1 1 10 9 16 11 7 9 15 0 1 15 1 9 10 9 1 9 0 1 9 0 2 10 9 16 15 13 13 9 14 9 2 9 2
10 3 13 7 10 9 10 0 3 13 2
23 9 1 9 10 9 1 11 7 1 9 9 15 3 13 14 10 9 1 9 15 10 0 2
19 10 9 2 7 10 9 3 2 13 9 3 2 0 1 10 9 10 0 2
40 7 1 9 1 10 15 2 3 10 9 16 10 9 10 0 3 16 15 13 13 10 9 1 9 0 2 16 1 9 15 13 10 9 13 0 7 13 1 15 2
40 0 16 13 1 10 9 15 3 9 14 9 0 1 9 0 1 9 2 7 1 9 1 9 0 9 10 9 2 7 9 1 9 3 0 1 2 10 9 2 2
36 7 10 9 10 0 13 16 9 0 3 15 13 1 9 9 0 3 2 13 1 2 9 10 10 9 10 0 2 7 3 16 4 13 1 15 2
53 7 16 9 9 1 11 13 9 0 14 15 13 14 9 2 10 9 1 15 9 14 9 10 9 10 0 16 15 0 2 1 9 13 14 10 9 10 0 15 2 14 9 15 7 14 9 15 2 7 13 1 15 2
40 10 9 16 11 13 13 3 10 9 1 10 9 16 13 7 13 14 0 1 9 2 10 9 1 9 0 2 2 7 2 13 14 9 15 10 0 3 1 9 2
25 1 9 9 15 13 11 2 2 3 7 3 13 1 10 9 16 10 9 13 1 15 13 1 11 2
67 3 13 1 9 15 16 15 13 14 15 13 14 10 9 2 3 9 1 9 0 2 3 9 10 9 10 0 1 3 2 16 11 15 13 1 10 9 1 9 9 1 10 15 8 2 2 13 1 9 2 13 1 9 7 1 9 10 9 2 13 1 9 9 3 0 2 2
44 11 13 13 1 9 15 16 9 9 2 10 9 1 9 10 9 10 0 2 0 13 15 9 1 10 9 10 3 0 14 2 10 9 1 9 2 1 10 9 10 0 2 0 2
47 13 3 1 9 0 13 16 7 9 10 9 7 9 10 9 13 13 1 9 0 7 0 1 10 9 10 0 1 10 9 10 0 2 9 1 10 15 13 13 13 3 1 10 9 1 11 2
43 16 13 9 1 9 0 7 15 13 1 9 0 2 13 10 9 0 2 9 16 4 13 1 10 9 10 0 1 13 0 1 9 9 10 9 7 10 9 16 13 14 15 2
31 7 10 3 16 13 1 9 0 13 1 10 9 10 0 2 1 9 0 14 10 9 2 13 3 0 14 13 1 10 9 2
34 3 0 13 14 2 9 10 9 2 2 7 3 13 10 9 9 0 0 2 16 3 13 3 9 0 7 9 0 0 2 7 9 0 2
30 1 12 1 9 15 10 0 3 2 13 9 11 1 11 1 9 2 9 16 13 1 9 7 13 16 15 9 2 11 2
54 9 3 13 13 14 15 2 1 16 13 15 9 16 13 1 15 1 1 10 9 2 13 9 2 7 1 9 0 7 0 13 14 15 16 3 9 2 11 4 13 1 10 9 2 13 7 13 2 1 9 2 9 2 2
41 13 1 9 15 9 0 0 7 0 3 2 3 2 4 13 1 9 7 1 9 13 14 9 15 10 0 1 9 0 14 9 7 9 1 10 9 16 13 15 9 2
44 1 9 14 9 1 11 2 11 13 1 9 14 11 11 3 13 3 1 12 9 2 7 12 9 13 1 10 9 10 0 16 9 15 13 1 15 1 9 10 9 1 10 9 2
24 3 3 13 1 11 13 12 9 9 1 9 7 9 15 2 7 1 9 15 1 11 13 9 2
42 9 9 15 1 9 15 10 0 3 14 10 9 10 0 1 9 10 9 10 0 16 13 3 1 9 2 13 9 3 7 13 16 3 13 10 9 1 13 1 10 11 2
45 13 15 0 13 16 11 10 0 0 2 10 9 15 2 1 9 2 11 2 2 7 9 9 9 15 1 9 15 14 11 11 13 1 9 10 9 16 13 10 9 1 11 2 11 2
26 10 9 16 13 9 1 9 9 16 13 1 2 9 9 2 13 1 9 15 14 10 9 1 10 9 2
22 10 9 10 15 13 13 2 3 7 10 9 14 9 9 15 14 11 11 13 1 9 2
77 7 1 10 9 1 10 9 2 1 11 7 1 9 9 13 9 13 14 9 16 10 9 13 1 9 0 7 15 13 13 14 9 10 9 1 9 10 9 1 9 1 10 9 10 0 2 4 16 15 16 13 14 11 11 13 13 14 10 9 10 0 13 14 10 9 16 13 1 15 1 10 9 10 0 2 0 2
29 3 1 10 9 13 12 1 9 10 9 2 11 11 2 2 15 3 13 1 9 2 7 4 16 15 13 1 9 2
25 15 3 13 3 13 2 7 0 16 13 9 14 0 1 9 2 7 16 9 13 1 2 15 2 2
21 13 13 9 1 10 9 2 11 11 13 1 9 14 9 16 15 13 16 3 13 2
44 15 13 1 13 1 9 14 9 9 2 11 2 2 7 4 16 15 3 13 9 1 13 9 9 2 16 4 13 14 10 9 1 10 9 16 13 1 9 10 9 7 10 9 2
24 7 9 15 1 15 1 9 1 10 11 11 2 13 7 13 14 9 11 1 9 7 15 9 2
48 7 10 9 13 4 13 0 3 1 10 9 2 9 2 11 2 13 2 3 7 3 2 1 9 0 2 14 10 9 2 10 11 2 9 10 9 7 10 9 1 2 9 9 2 14 11 11 2
18 8 8 2 9 13 3 1 10 9 16 9 10 9 13 1 9 15 2
42 1 10 9 10 15 3 13 16 2 9 10 9 13 3 9 9 9 9 16 13 1 9 10 9 11 11 10 12 1 2 9 10 11 2 10 9 7 10 9 10 0 2
6 9 15 1 15 2 2
62 7 11 11 2 11 13 1 9 15 16 2 3 13 9 10 9 1 10 9 3 2 10 9 7 1 10 9 9 2 2 7 16 9 2 11 2 13 2 3 2 10 9 1 9 2 1 9 11 7 1 9 16 9 13 16 13 1 9 15 1 11 2
68 13 9 16 9 10 9 10 0 13 13 14 10 9 10 15 2 7 16 4 13 9 1 10 9 16 2 4 16 9 1 10 9 13 2 7 13 1 10 9 10 0 2 9 14 9 2 9 9 7 9 7 13 14 15 1 9 1 9 2 2 2 10 9 2 2 12 2 2
28 13 16 9 2 3 7 13 1 15 10 9 1 10 9 2 13 1 15 9 1 15 16 0 1 12 10 9 2
56 10 9 16 13 9 1 10 9 7 1 11 7 13 13 12 9 1 9 9 13 3 15 1 9 15 2 1 15 9 4 2 13 2 9 1 13 9 1 9 15 10 0 2 1 9 9 16 9 2 11 2 3 13 7 13 2
21 10 9 13 16 10 9 10 0 13 13 1 10 9 16 4 13 14 9 9 15 2
30 7 15 3 13 3 1 13 10 12 13 9 9 2 16 4 13 1 10 9 3 3 7 3 7 3 7 1 10 9 2
12 7 9 15 13 2 13 3 1 9 9 9 2
16 15 10 9 2 7 1 10 9 13 9 0 1 13 14 15 2
23 16 13 11 11 7 11 11 9 1 10 9 16 9 2 11 2 13 14 15 1 10 9 2
28 9 15 2 7 9 10 10 0 16 13 1 11 11 2 0 2 0 16 13 13 14 10 10 9 4 3 13 2
32 9 11 13 9 0 1 13 14 10 9 16 13 1 9 10 9 1 11 2 15 13 13 1 9 15 2 7 3 3 1 11 2
16 9 1 10 9 13 3 3 3 9 7 9 2 7 3 9 2
51 1 10 9 3 2 7 1 9 10 9 3 2 13 10 9 13 14 9 15 14 10 10 9 1 9 10 9 16 1 15 13 1 9 1 10 3 16 13 14 10 9 12 15 7 13 1 9 7 1 9 2
49 9 10 9 0 13 1 9 9 9 15 1 9 14 9 1 9 10 9 1 12 10 9 2 16 16 13 14 15 9 10 9 2 9 10 9 10 0 13 4 13 0 3 1 9 9 16 13 0 2
16 1 10 9 13 9 13 9 1 9 11 16 13 1 10 9 2
34 15 16 13 14 9 15 14 11 11 2 1 10 0 16 13 14 9 15 1 10 9 2 7 4 1 15 13 13 1 9 15 10 0 2
37 4 13 9 0 16 13 9 1 9 15 14 9 2 11 2 2 7 16 13 14 10 9 16 9 13 1 9 16 11 11 2 11 13 1 9 15 2
14 4 13 9 16 1 15 2 11 13 1 10 9 11 2
14 15 4 13 3 1 9 1 11 2 11 7 1 11 2
49 10 9 10 0 16 9 11 13 1 9 15 9 9 15 10 0 14 10 9 1 10 9 10 13 13 13 15 1 9 9 1 11 7 1 9 1 9 2 16 13 13 1 9 10 9 9 14 9 2
21 10 9 4 13 9 16 13 3 3 14 10 9 7 3 14 15 1 9 10 9 2
14 15 4 13 1 9 10 9 13 9 0 1 10 9 2
12 10 9 1 10 9 10 0 13 1 12 9 2
47 13 10 9 2 10 0 7 10 0 2 14 9 7 14 3 2 9 1 9 11 10 0 2 14 11 16 13 3 14 10 9 10 0 2 7 14 11 11 2 9 9 13 1 9 9 0 2
53 7 13 10 9 2 10 13 7 10 13 2 16 13 1 15 9 9 16 13 1 9 9 0 14 9 0 7 0 7 14 3 16 13 3 9 0 2 14 9 9 9 9 7 14 9 9 11 16 13 1 9 15 2
41 13 9 0 1 9 10 12 1 10 9 3 2 7 10 9 13 1 9 0 1 10 9 2 1 15 10 13 7 13 13 1 10 9 1 3 16 3 13 9 0 2
34 9 13 1 9 9 15 2 16 7 7 3 13 14 10 9 10 0 7 10 0 16 13 1 10 9 1 15 2 13 16 13 10 9 2
68 7 16 9 3 2 4 13 2 7 1 10 9 15 3 13 14 10 9 1 10 9 2 9 13 14 10 9 3 2 1 9 1 11 3 13 10 9 2 9 15 14 9 11 13 1 10 9 1 9 9 0 1 14 15 2 7 10 9 1 10 9 13 9 10 4 13 13 2
22 1 10 9 16 1 10 9 2 10 9 2 13 10 9 7 10 9 1 9 1 9 2
6 7 13 3 9 12 2
7 15 13 0 7 13 0 2
19 15 13 0 2 0 7 0 2 7 7 3 9 1 10 9 1 10 9 2
33 1 9 9 15 13 13 16 10 9 10 0 2 0 2 16 13 12 9 7 3 7 3 2 13 1 10 9 3 12 0 14 9 2
33 3 9 0 1 10 9 16 15 2 0 16 16 13 2 13 16 13 1 9 10 9 2 7 3 3 9 0 2 0 16 16 13 2
33 15 13 13 1 9 15 14 3 10 9 2 9 2 3 3 1 9 15 14 10 2 7 3 13 3 1 9 15 7 1 9 0 2
10 3 13 13 1 9 15 14 10 9 2
11 9 10 9 1 10 9 10 12 13 0 2
15 13 1 15 9 9 16 13 1 10 11 1 9 9 15 2
45 9 4 13 9 0 7 0 2 7 9 2 1 10 9 7 1 10 9 2 0 1 15 1 9 15 10 0 2 16 13 16 7 3 13 10 9 1 15 9 13 13 1 9 15 2
12 10 9 13 9 14 15 7 14 10 10 9 2
40 3 3 13 1 9 10 9 13 1 10 9 10 12 2 16 4 13 13 10 9 10 0 10 0 2 16 9 15 10 0 2 0 16 16 13 2 1 10 9 2
33 10 9 13 1 10 9 2 13 13 16 10 9 1 12 1 12 10 9 1 10 11 2 7 3 3 12 1 12 9 10 11 13 2
54 1 7 16 10 9 13 3 9 0 7 0 16 3 13 1 15 1 13 9 12 0 9 2 16 13 1 10 9 7 13 13 1 9 15 3 9 0 2 13 16 13 1 15 3 3 9 12 9 9 11 2 11 11 2
47 4 16 11 13 0 1 10 9 10 15 16 16 13 1 9 10 9 2 1 10 9 14 10 9 2 7 13 13 3 1 11 10 0 1 9 15 10 0 2 16 15 13 1 9 10 9 2
45 15 13 16 1 9 13 9 2 7 10 10 9 10 0 13 1 10 9 16 4 13 1 9 11 9 15 7 1 9 10 9 2 0 1 9 15 2 13 13 1 9 1 10 9 2
22 4 16 13 1 10 9 10 12 16 16 13 13 1 3 16 13 7 13 1 10 11 2
27 1 1 10 15 15 13 1 13 9 0 2 1 13 13 1 12 1 12 10 9 16 13 16 13 4 13 2
30 15 13 13 13 9 2 7 1 9 9 13 1 10 9 13 3 7 3 1 9 0 2 1 3 2 9 16 13 0 2
25 7 3 11 13 9 10 9 10 15 1 3 16 13 1 10 9 14 10 9 1 10 9 1 11 2
9 1 10 9 10 0 13 1 9 2
35 9 10 9 2 1 10 9 2 13 1 9 0 2 16 15 4 13 1 9 1 9 0 3 2 3 10 0 3 2 16 9 0 14 15 2
14 11 13 13 1 3 16 13 1 10 9 10 12 3 2
7 4 16 3 3 13 3 2
17 9 10 9 2 16 13 14 15 3 7 3 2 13 13 14 15 2
66 1 10 9 14 9 1 9 7 1 9 2 16 9 13 1 9 10 9 7 9 13 9 7 13 3 14 10 9 16 13 4 1 9 7 13 4 13 2 11 13 7 13 1 3 9 3 0 14 2 13 1 15 3 3 2 2 16 10 9 10 15 13 3 10 9 2
7 15 13 13 14 9 11 2
32 12 9 13 1 3 13 10 9 10 0 1 10 9 2 7 3 12 9 1 3 13 14 9 10 9 2 16 1 15 3 13 2
30 10 9 10 0 2 16 15 3 9 9 10 9 16 13 1 11 7 13 1 10 9 2 13 13 16 11 13 1 3 2
18 10 9 2 10 9 10 0 2 1 15 2 13 13 1 11 10 0 2
18 11 13 13 3 15 10 9 9 12 9 16 4 16 13 3 9 0 2
22 15 13 14 10 9 1 9 11 2 16 13 14 9 15 1 9 10 11 1 12 9 2
31 1 12 12 10 9 15 2 0 1 9 15 7 1 9 15 16 13 7 13 2 13 1 9 15 2 7 10 9 13 13 2
8 1 11 10 9 3 0 9 2
27 1 10 12 10 12 2 1 3 13 10 9 10 0 1 10 9 15 1 10 9 2 13 12 9 1 9 2
26 9 15 10 0 10 0 14 10 9 1 9 15 1 10 9 13 14 10 9 2 7 3 13 14 15 2
21 1 10 9 16 13 13 10 9 13 14 9 15 10 0 7 10 0 16 13 0 2
43 15 7 1 11 2 1 11 2 1 11 10 0 7 1 9 0 1 11 2 15 1 11 2 1 9 11 2 1 11 7 1 9 0 1 11 2 7 15 1 10 9 11 2
22 1 9 15 14 11 13 3 9 0 2 0 7 13 9 2 9 2 16 13 9 0 2
26 15 10 9 10 3 2 0 2 16 13 1 12 10 9 16 13 15 1 15 1 9 10 9 10 13 2
30 9 0 16 13 13 13 11 2 7 3 3 13 7 13 9 0 1 9 15 9 0 0 2 16 13 1 12 9 0 2
38 10 9 13 1 9 16 13 1 12 10 9 10 0 1 9 15 14 9 2 10 9 13 9 2 7 16 13 3 1 9 7 13 9 3 2 0 0 2
23 1 9 10 9 9 10 9 2 16 1 15 13 9 1 12 12 9 9 2 13 10 9 2
15 9 0 13 1 9 2 7 9 0 13 1 10 9 15 2
16 10 9 16 16 13 0 1 9 13 4 1 9 9 1 9 2
53 12 9 13 1 15 9 9 2 1 10 12 9 10 9 10 0 7 10 0 2 9 9 1 10 9 2 7 9 7 9 3 2 13 13 1 9 10 9 16 13 1 15 1 10 9 7 9 13 13 13 1 15 2
16 9 15 13 0 3 1 9 15 2 1 9 15 13 1 9 2
13 9 15 13 14 15 1 0 10 9 1 9 15 2
25 10 16 13 13 9 2 9 1 9 2 10 9 10 0 2 16 13 1 9 11 10 9 1 11 2
15 10 16 13 13 15 2 15 13 2 3 13 13 1 15 2
20 15 13 16 13 9 7 1 16 13 7 1 16 10 9 13 1 9 9 15 2
28 11 11 13 13 14 15 1 9 15 10 0 14 10 9 10 0 2 3 13 3 14 10 9 10 0 1 15 2
32 13 1 10 9 9 0 2 15 13 1 9 15 1 9 10 9 2 7 1 9 1 15 13 3 9 1 9 10 9 10 0 2
29 1 9 15 14 9 15 13 10 2 9 2 16 10 1 9 10 9 10 0 13 1 15 9 0 3 1 10 15 2
12 10 9 2 1 9 0 2 13 1 9 0 2
11 11 13 9 1 9 0 2 0 2 0 2
9 15 10 9 10 0 1 9 15 2
16 1 13 1 10 11 13 13 1 13 16 15 13 14 10 9 2
21 3 2 3 13 7 14 10 9 16 1 15 13 14 9 15 2 1 10 9 3 2
15 12 1 10 9 13 13 1 9 9 16 13 1 9 11 2
38 1 10 9 16 13 13 1 15 2 13 3 1 9 9 10 9 7 0 0 12 16 13 13 1 9 10 9 1 9 7 1 15 9 9 1 10 9 2
13 7 16 13 1 11 2 11 13 11 9 0 3 2
17 15 13 1 9 0 0 2 13 1 9 15 7 13 1 9 15 2
20 3 13 13 1 9 15 9 0 7 13 14 15 1 9 2 1 13 9 11 2
34 15 13 1 10 9 16 1 9 10 9 15 13 1 9 10 9 2 7 10 9 13 1 15 16 16 13 1 10 9 10 9 10 15 2
36 1 11 3 13 3 2 9 2 14 3 2 7 1 9 9 15 3 10 9 16 13 13 14 15 13 3 3 9 14 9 2 3 2 9 2 2
20 7 11 10 9 13 3 3 0 1 9 16 13 2 7 7 3 3 3 0 2
43 9 7 13 3 9 0 1 10 9 16 13 1 15 10 11 14 15 2 7 7 3 1 12 1 15 15 13 14 9 10 9 7 13 3 1 9 10 9 10 0 14 15 2
59 1 9 0 13 11 9 0 1 10 9 10 0 2 10 3 13 13 16 13 1 15 9 1 10 9 13 14 10 9 2 3 13 10 9 4 1 9 0 3 1 10 9 0 16 9 13 1 9 15 10 0 14 10 9 1 9 9 0 2
47 1 10 9 10 0 13 11 14 10 9 10 15 2 7 10 9 13 9 0 1 9 2 13 10 9 1 9 10 9 2 13 10 9 14 10 9 2 9 1 9 9 10 9 1 9 9 2
33 1 15 10 9 14 11 11 2 15 13 2 0 2 3 1 15 14 11 2 2 0 2 3 2 0 2 9 15 10 0 0 3 2
36 11 10 0 4 3 1 11 14 10 9 16 10 11 13 1 9 15 2 7 10 9 13 9 13 15 1 9 15 2 1 13 12 1 14 15 2
12 3 11 4 14 9 15 1 10 11 1 11 2
3 3 3 2
30 10 9 14 11 13 1 10 9 2 1 15 1 15 9 0 16 13 3 1 10 9 10 0 14 10 9 2 10 9 2
30 10 9 13 1 15 16 10 9 10 0 1 9 10 9 13 13 3 1 9 1 15 2 1 10 9 1 10 9 15 2
19 10 9 10 0 13 13 1 10 9 2 7 1 9 9 15 1 9 0 2
19 14 13 9 15 1 3 0 4 13 13 14 9 15 1 11 1 9 0 2
16 13 13 7 11 13 13 1 0 14 10 9 10 0 10 15 2
36 3 7 3 2 3 1 9 9 15 10 0 2 1 10 9 7 1 10 9 2 15 4 3 13 1 11 11 1 11 11 1 15 13 1 15 2
52 1 12 1 9 10 9 11 2 11 2 3 3 1 10 9 16 13 1 15 2 1 9 10 9 10 12 2 9 10 9 14 10 9 10 0 2 13 9 0 16 10 9 13 14 15 13 3 1 10 0 3 2
29 7 15 13 16 3 3 13 9 1 10 9 10 0 2 7 13 13 3 1 10 9 16 13 3 1 11 14 15 2
28 3 13 1 15 9 0 1 9 15 15 2 13 1 11 9 7 1 15 2 14 13 14 15 3 1 9 15 2
42 15 13 0 2 3 13 1 15 9 13 1 10 9 7 1 10 9 7 1 10 9 2 13 1 15 2 7 11 11 13 1 9 14 9 2 9 2 13 2 9 9 2
7 3 3 13 1 15 12 2
16 3 15 13 3 1 10 9 2 15 4 1 15 14 9 15 2
40 13 3 2 1 11 2 1 11 7 1 9 10 9 2 13 9 13 9 16 13 7 9 15 2 9 9 1 9 11 2 2 1 9 2 9 7 9 2 2 2
13 9 10 9 13 3 1 9 2 11 13 10 9 2
19 1 9 10 9 10 0 15 13 1 10 9 2 7 1 9 2 12 13 2
20 1 9 7 9 1 1 3 13 10 9 16 13 1 10 9 13 1 10 9 2
19 10 9 16 13 3 13 13 14 9 15 7 14 9 2 10 9 14 15 2
34 3 11 13 13 2 10 9 13 16 4 13 1 10 9 13 9 9 2 1 10 9 1 9 16 13 1 10 9 10 0 1 9 9 2
17 1 9 0 13 11 10 9 10 3 2 0 10 0 1 10 9 2
51 9 10 9 14 15 13 1 1 9 9 0 2 9 13 13 2 1 10 9 10 9 7 10 9 2 3 12 13 1 9 10 9 2 1 9 16 13 1 9 15 7 13 1 9 10 9 10 0 2 11 2
22 11 13 1 15 9 7 9 9 16 13 13 1 15 14 9 10 11 2 11 2 11 2
13 13 13 1 15 9 1 9 15 7 1 9 15 2
21 9 11 3 13 0 3 2 13 16 13 9 13 1 10 9 1 9 1 9 15 2
19 11 13 13 1 0 1 15 9 16 13 1 15 13 1 9 1 10 9 2
60 1 3 16 13 1 9 15 14 9 10 9 15 2 13 9 3 1 9 10 9 2 15 13 13 1 9 9 10 9 14 15 2 13 1 9 10 9 1 10 9 2 3 10 9 10 0 7 10 9 2 7 10 3 16 13 13 1 9 15 2
20 1 1 10 9 15 15 12 1 9 10 9 10 3 2 0 10 0 16 13 2
35 9 11 13 1 15 14 10 9 2 9 9 10 9 2 2 7 15 13 13 9 9 1 10 9 16 1 9 2 9 7 9 2 1 11 2
35 1 3 16 13 1 9 10 9 7 10 9 1 10 9 2 13 11 1 9 15 9 9 0 14 9 7 9 16 13 1 15 1 10 9 2
59 12 1 15 13 14 15 3 13 9 1 9 9 2 15 13 14 15 1 9 10 9 14 15 13 1 9 2 7 1 15 13 9 12 1 9 2 1 9 13 16 15 13 2 13 14 15 1 9 1 9 10 9 7 13 1 15 9 0 2
29 3 2 3 2 13 3 1 9 10 9 2 1 10 9 10 0 2 13 14 15 2 7 11 13 1 15 1 9 2
25 3 15 13 3 2 13 1 10 9 2 7 15 9 10 9 16 13 9 15 2 1 9 10 12 2
85 15 13 9 0 2 13 9 10 9 10 0 2 11 13 1 9 1 9 2 9 13 1 15 9 1 15 2 7 13 9 11 2 7 13 10 9 7 13 14 10 9 1 16 13 2 7 3 13 10 9 7 13 14 10 9 2 7 11 11 13 9 0 1 10 9 2 9 13 7 13 2 9 13 7 13 2 7 9 1 9 7 9 4 3 2
41 9 10 9 14 15 2 9 0 14 9 7 9 1 9 10 9 16 13 14 11 1 9 10 12 2 13 3 1 9 10 12 2 14 15 2 11 13 13 14 15 2
17 13 14 15 1 10 9 2 3 13 13 3 1 16 13 1 15 2
19 11 13 16 10 10 9 16 15 13 3 13 14 15 14 10 9 10 15 2
14 7 10 9 13 0 10 3 2 15 3 13 13 9 2
11 3 15 13 13 7 13 13 1 9 15 2
8 13 13 1 15 1 10 9 2
20 15 13 9 1 10 15 2 14 13 1 9 10 9 14 15 2 1 10 9 2
16 13 1 10 9 2 3 13 13 3 1 16 13 1 10 9 2
7 11 13 16 13 10 11 2
20 12 1 10 12 1 9 9 10 9 3 13 0 2 1 9 9 3 1 12 2
50 13 1 15 1 11 9 1 14 15 2 7 1 9 9 15 9 10 9 16 13 1 9 13 1 3 12 12 2 7 10 10 9 16 13 0 1 15 2 3 1 9 7 9 2 13 1 3 12 12 2
30 7 1 10 15 2 13 14 11 2 3 13 14 10 9 1 3 16 13 9 1 3 16 13 13 15 7 3 13 15 2
10 11 13 16 15 0 1 9 1 9 2
20 7 3 15 0 1 10 9 2 3 1 10 9 10 0 2 3 1 10 9 2
11 1 1 9 15 0 9 0 14 10 9 2
9 15 3 13 14 15 13 1 15 2
25 10 9 3 3 13 3 11 13 14 15 2 13 2 7 3 3 13 1 15 2 1 9 3 0 2
19 15 13 1 9 1 10 9 10 0 16 13 1 15 2 9 15 13 9 2
13 3 15 13 3 10 12 13 3 7 10 12 3 2
7 0 16 9 13 13 3 2
7 3 15 13 4 13 3 2
22 1 10 9 15 13 14 15 1 16 3 13 3 2 13 1 15 7 13 1 9 0 2
25 15 13 1 9 9 0 16 13 1 9 15 14 9 0 7 1 15 9 0 16 1 9 15 9 2
11 1 16 13 13 13 9 9 0 7 0 2
11 13 9 0 1 10 9 2 7 3 9 2
8 3 9 10 9 13 9 0 2
25 11 11 13 16 1 10 3 3 13 3 2 7 13 9 9 1 10 3 16 3 13 14 15 3 2
19 13 16 13 1 15 9 1 9 10 9 2 15 13 14 15 3 2 13 2
9 11 11 13 9 0 7 9 11 2
16 15 9 0 7 9 9 2 1 9 9 10 12 1 9 15 2
11 11 13 9 0 2 0 2 9 10 9 2
19 9 14 15 2 16 13 9 9 9 1 11 2 13 14 15 1 10 9 2
19 16 16 15 13 3 13 1 15 9 0 2 1 15 9 3 13 1 9 2
16 7 11 13 1 9 15 9 0 7 13 3 14 9 14 15 2
10 1 9 13 14 11 7 13 1 11 2
11 15 13 16 13 1 11 7 13 1 9 2
15 3 13 13 1 9 14 15 2 7 3 12 9 13 13 2
16 3 13 2 1 9 12 10 9 2 16 9 1 11 4 13 2
4 3 15 13 2
6 9 14 15 3 13 2
11 3 15 13 14 15 3 9 11 14 15 2
14 9 15 13 16 3 1 10 9 4 13 13 14 15 2
37 11 13 9 0 16 13 1 15 1 10 9 2 7 3 1 15 15 13 9 1 9 0 1 9 9 10 9 16 3 9 15 1 9 2 11 2 2
17 12 10 9 16 14 9 15 13 13 3 13 1 9 15 7 0 2
18 7 10 9 10 0 16 14 15 13 11 13 13 16 13 14 9 15 2
15 1 16 9 7 9 3 13 1 10 9 15 13 9 0 2
30 13 4 3 13 1 15 16 15 13 1 10 9 9 3 1 9 15 14 9 10 9 10 0 16 14 15 15 13 13 2
31 10 9 16 13 9 15 1 11 15 9 16 13 9 1 9 10 9 10 0 13 0 2 7 10 9 13 3 1 10 9 2
11 11 13 3 13 1 10 9 1 9 15 2
46 13 4 3 13 1 9 15 1 9 12 1 9 10 9 14 10 9 2 2 10 9 13 9 16 9 15 9 7 9 2 2 2 7 9 0 3 1 9 2 1 9 7 1 9 2 2
11 15 10 9 1 10 9 7 1 10 9 2
10 3 10 9 13 9 1 2 11 2 2
25 3 9 9 10 9 1 9 11 16 13 1 9 10 9 1 9 10 9 13 9 1 9 0 15 2
39 9 12 1 9 10 9 2 16 13 1 9 0 1 14 0 11 2 13 1 9 15 15 2 9 9 11 0 2 15 9 1 10 9 14 15 1 10 9 2
59 7 7 7 16 13 1 10 9 10 0 2 0 7 0 2 7 10 9 14 3 13 10 9 14 3 2 3 10 9 0 10 9 10 0 7 9 10 9 7 9 10 9 1 9 10 9 7 9 7 3 3 7 3 9 13 1 9 0 2
12 11 2 13 14 15 9 0 7 9 12 0 2
18 3 16 12 10 9 1 10 9 1 15 13 16 13 1 10 9 9 2
21 13 1 9 15 10 0 10 9 16 13 2 10 9 16 13 2 10 9 16 13 2
29 3 16 1 9 13 1 3 16 13 1 10 9 10 0 16 13 1 15 1 16 13 1 9 15 14 9 9 15 2
31 1 10 9 16 13 1 10 9 13 1 10 9 7 1 9 10 9 7 13 1 0 2 16 15 13 13 14 12 10 12 2
13 3 0 1 15 16 10 10 9 3 13 1 15 2
38 10 9 10 0 16 13 1 15 13 1 11 2 7 15 13 9 0 3 2 3 14 15 2 9 9 10 9 10 0 2 10 9 13 13 1 10 9 2
7 9 1 15 13 1 11 2
11 15 13 10 9 10 0 3 1 9 15 2
12 13 13 3 10 9 10 0 1 2 9 2 2
7 1 9 15 15 3 9 2
24 9 13 9 0 2 7 15 3 13 1 9 16 13 14 9 15 7 1 9 16 13 14 15 2
5 3 0 1 15 2
25 13 0 16 13 1 15 9 7 9 13 1 15 2 3 2 2 13 3 16 13 2 15 13 3 2
32 7 3 13 1 10 9 10 15 2 3 0 2 2 3 10 9 14 15 7 10 9 14 15 1 10 9 10 0 14 15 13 2
32 15 3 13 3 16 1 9 10 9 10 0 4 13 9 0 3 1 10 9 10 0 2 9 10 9 2 9 10 9 7 3 2
14 15 9 16 3 7 1 9 13 1 9 7 1 9 2
21 15 4 13 9 1 10 15 7 13 1 10 9 14 9 7 9 1 9 10 9 2
37 3 2 1 9 10 9 2 15 13 9 16 3 11 11 2 12 1 12 9 8 16 13 1 15 2 13 3 1 9 9 0 16 13 1 10 9 2
18 15 13 3 16 13 9 13 1 10 9 10 15 9 1 11 14 3 2
7 4 13 14 15 3 3 2
30 15 13 3 16 13 14 15 2 3 4 13 9 1 10 9 7 13 1 15 2 7 3 13 9 1 3 16 13 3 2
9 10 9 14 15 4 13 0 3 2
20 15 13 13 1 15 1 3 16 13 2 13 14 15 3 13 1 9 0 3 2
21 15 13 14 15 1 9 0 2 7 1 16 13 1 11 13 9 0 1 9 0 2
32 1 9 0 13 1 15 9 2 16 16 9 15 13 13 1 11 2 11 7 9 15 1 10 11 13 13 1 10 9 9 9 2
21 3 1 15 13 1 10 9 10 0 16 0 1 15 2 3 3 7 1 10 9 2
28 14 13 1 11 14 10 9 16 13 1 9 15 13 1 15 4 13 9 1 15 2 9 2 3 2 0 2 2
13 3 13 1 9 15 14 9 15 16 9 13 9 2
27 0 16 16 13 1 15 12 9 2 1 11 2 2 13 9 2 1 9 15 2 16 16 13 1 10 9 2
25 7 14 13 1 15 1 15 2 13 1 10 9 16 15 13 3 9 0 16 3 13 9 7 9 2
13 12 1 12 10 9 10 15 13 10 9 11 11 2
53 3 13 1 15 10 9 16 1 10 10 9 16 13 1 15 2 7 1 10 9 1 10 9 10 0 2 15 4 13 16 9 15 9 1 15 9 2 3 9 15 7 3 9 2 9 15 10 0 13 1 10 9 2
6 13 3 9 1 15 2
11 1 9 15 13 9 7 13 1 15 9 2
27 4 1 15 13 14 15 7 13 1 15 3 1 15 16 13 13 1 10 9 2 7 13 4 13 14 15 2
17 15 4 13 14 16 13 1 9 15 7 13 1 15 9 1 3 2
25 3 1 15 4 1 15 13 1 10 9 10 0 14 10 9 10 0 16 0 1 10 9 10 0 2
71 1 10 9 13 1 12 9 9 16 1 15 4 13 9 15 14 10 9 10 0 2 1 10 13 2 13 1 10 9 2 2 9 11 2 9 11 2 7 10 9 10 0 1 10 9 7 10 9 16 1 15 2 7 14 12 10 9 10 0 13 1 9 15 1 16 3 13 1 9 15 2
56 1 9 9 15 2 13 16 3 12 13 1 9 10 9 16 13 9 1 15 1 11 2 7 16 13 9 1 13 16 13 16 1 15 13 14 10 15 16 13 2 16 16 15 13 1 15 3 13 1 10 9 16 13 14 15 2
54 3 13 9 7 9 0 2 16 1 0 7 1 0 2 13 16 1 15 13 1 2 9 9 2 7 1 11 2 1 9 15 2 16 13 1 10 9 2 7 3 1 9 2 1 9 15 9 10 9 1 9 11 2 2
48 2 11 14 15 2 16 16 13 7 13 2 7 16 16 13 1 9 15 0 7 1 15 16 13 14 15 9 0 16 13 1 10 9 1 15 1 10 9 2 14 15 9 0 3 13 2 3 2
44 7 13 1 9 14 9 9 15 2 2 11 11 13 1 10 9 16 13 9 2 2 2 4 13 13 16 13 7 13 2 16 4 13 9 9 16 3 13 1 15 9 1 9 2
23 13 1 9 0 2 0 2 14 3 9 10 9 1 9 15 15 13 1 9 1 10 9 2
28 15 13 2 2 1 10 9 16 13 10 9 13 1 15 1 9 10 9 2 3 1 9 0 7 3 1 9 2
7 11 13 1 10 9 2 2
88 3 9 7 3 9 15 2 7 3 13 1 10 9 1 9 10 9 2 1 10 9 16 13 1 10 9 2 1 2 9 11 2 2 1 9 10 11 7 9 15 10 0 2 1 9 10 9 13 10 9 16 13 10 9 2 1 9 9 16 13 1 9 9 15 2 7 3 13 10 9 10 0 1 10 9 2 7 15 13 3 9 0 1 10 2 9 2 2
52 3 0 13 10 9 7 10 9 14 13 14 10 9 10 0 14 15 2 2 15 13 1 10 9 2 15 9 2 15 13 13 1 3 15 13 2 3 2 13 1 1 12 1 12 9 14 16 13 1 15 3 2
15 1 10 9 13 7 13 2 2 3 15 1 10 9 2 2
18 3 13 9 1 10 9 2 1 1 13 14 10 9 1 9 10 9 2
22 1 10 9 10 0 16 13 2 13 3 2 7 13 16 3 3 2 13 2 1 9 2
28 3 3 2 1 9 15 2 13 13 1 9 15 10 9 2 7 6 1 13 1 15 2 13 9 2 14 3 2
20 13 2 13 2 13 7 13 2 13 1 9 7 13 1 9 9 1 10 9 2
19 7 2 10 9 0 3 1 3 16 9 15 0 7 9 15 13 7 13 2
50 1 3 16 13 2 13 7 13 10 9 0 2 0 2 2 9 9 13 1 11 2 2 15 13 2 2 9 2 2 2 9 2 2 2 9 2 2 7 13 3 2 9 2 2 2 0 2 7 3 2
15 9 15 9 0 2 16 13 2 1 9 15 9 0 2 2
17 10 11 13 9 10 9 2 7 13 9 7 9 0 1 9 15 2
13 1 13 15 4 9 2 9 15 13 13 1 15 2
24 15 13 16 1 9 10 11 13 1 10 9 3 9 16 9 15 10 0 2 11 14 15 2 2
5 3 2 7 3 2
7 3 15 13 1 10 9 2
17 10 9 10 0 14 15 13 2 13 1 9 7 13 1 9 2 2
37 1 10 10 9 13 3 13 14 10 9 2 1 9 0 2 7 13 14 10 9 15 13 9 15 2 7 15 13 1 15 2 7 15 9 9 15 2
8 13 16 9 15 13 1 9 2
58 7 1 9 15 13 9 7 9 2 13 13 9 16 9 15 13 12 9 9 1 1 13 1 10 9 16 13 1 15 9 2 7 1 1 3 13 9 1 11 2 13 1 15 10 9 2 2 2 7 13 1 9 0 3 1 10 11 2
28 3 4 9 0 0 1 9 10 9 2 16 13 13 14 10 9 1 9 10 9 1 9 10 9 1 9 11 2
63 15 13 16 0 12 9 2 10 9 10 12 2 16 1 15 15 13 14 10 10 9 2 13 16 1 15 9 16 10 9 11 13 12 1 10 9 10 0 3 1 9 15 2 3 13 10 9 2 7 4 13 9 16 1 9 15 13 9 7 3 3 13 2
36 10 9 13 16 9 1 10 9 10 0 14 10 9 10 13 4 13 13 1 10 9 1 9 10 9 2 9 16 13 1 10 9 14 10 9 2
26 13 1 15 0 16 3 13 10 9 16 13 14 10 10 9 3 2 7 9 13 10 12 1 9 15 2
27 1 12 9 13 16 13 9 2 16 1 15 10 9 11 13 1 9 0 2 7 10 9 1 9 13 13 2
15 13 1 15 9 16 3 15 3 0 1 10 9 10 15 2
26 3 2 7 13 9 16 13 1 9 1 9 2 14 13 14 10 9 2 10 9 13 13 15 1 15 2
38 1 9 1 15 13 9 15 2 7 10 9 4 13 2 10 12 13 1 15 14 9 10 9 14 15 2 7 3 13 16 3 15 4 13 14 10 9 2
6 15 3 1 10 13 2
48 10 9 10 12 2 10 3 0 1 9 15 2 13 16 1 10 15 13 9 16 13 16 15 9 10 9 16 13 13 1 10 9 7 1 10 16 13 1 15 2 7 3 7 13 14 15 3 2
19 7 1 10 9 15 3 13 9 1 10 15 16 9 13 13 1 9 15 2
31 1 9 1 10 9 13 3 9 16 1 10 9 13 1 15 2 7 3 15 13 3 13 1 9 7 16 13 13 14 15 2
16 13 1 9 1 11 11 2 7 1 9 1 10 9 11 11 2
18 1 10 3 16 15 13 3 2 11 11 9 13 10 9 10 3 0 2
26 15 0 1 10 10 9 1 10 9 2 13 1 15 3 9 2 7 15 13 7 15 13 0 1 9 2
16 9 0 13 1 9 15 14 10 10 9 10 0 7 13 3 2
24 7 13 4 13 9 1 9 2 13 13 16 1 9 2 1 9 0 2 10 9 3 13 13 2
2 3 2
14 11 13 14 10 9 7 3 14 10 9 13 14 15 2
22 13 9 9 9 16 13 9 9 1 10 9 14 10 9 7 1 10 9 14 10 9 2
9 1 10 9 13 3 4 13 9 2
13 11 13 13 1 2 15 10 9 1 9 1 9 2
11 15 13 13 1 15 12 12 9 1 9 2
6 0 14 3 15 13 2
46 13 1 15 9 2 16 13 9 3 0 14 9 16 9 15 3 13 1 10 9 7 1 10 9 2 7 9 1 15 3 3 13 1 10 9 10 9 14 10 9 2 7 15 1 15 2
13 3 16 13 14 15 13 10 9 10 0 14 15 2
33 13 1 15 9 16 10 9 14 15 1 9 10 9 1 12 9 13 3 3 1 10 9 16 15 13 1 15 7 3 1 10 9 2
83 9 2 16 1 12 9 10 9 10 0 10 9 13 0 2 10 9 13 1 10 9 10 0 2 7 10 9 13 1 9 10 9 3 2 1 12 9 10 9 10 15 3 13 11 14 9 10 9 2 7 7 1 9 10 9 14 12 2 15 13 1 9 0 3 3 9 10 9 1 10 9 16 9 15 13 2 7 13 3 1 12 9 2
3 15 13 2
12 10 9 11 13 3 2 2 9 2 9 2 2
11 3 13 1 15 9 1 10 9 14 15 2
15 0 16 13 13 16 13 14 10 9 1 9 1 10 15 2
14 7 1 9 15 15 3 13 13 7 3 9 9 0 2
18 15 13 14 15 1 9 10 9 1 9 12 13 1 9 1 9 11 2
48 9 1 10 9 13 14 15 3 2 7 13 1 15 9 1 9 2 7 11 3 13 13 2 7 15 13 9 15 9 1 9 2 2 3 2 13 1 15 9 1 9 2 7 9 1 9 2 2
9 15 13 9 9 15 1 9 12 2
30 15 13 16 3 1 9 9 16 3 3 13 16 15 13 1 9 15 14 9 9 15 3 1 12 9 13 11 1 13 2
35 13 1 15 1 9 0 3 1 10 9 10 0 3 7 3 1 10 9 10 3 10 2 3 0 16 15 3 3 13 9 1 9 1 9 2
6 15 13 16 15 13 2
18 15 13 12 10 9 10 0 1 10 9 16 9 15 7 9 15 0 2
9 15 13 1 9 1 9 12 3 2
11 1 9 9 10 12 13 11 1 9 0 2
29 1 9 10 9 10 0 16 13 1 10 9 10 15 2 3 13 9 10 9 7 10 9 16 1 15 13 14 15 2
7 7 1 10 9 13 13 2
44 3 3 1 9 9 16 15 13 13 1 15 13 1 10 9 9 9 2 16 1 15 13 16 10 9 11 13 13 1 15 9 1 15 9 13 14 10 9 16 1 9 10 9 2
23 15 13 9 10 9 2 11 11 2 7 15 13 14 10 9 2 14 15 13 1 9 0 2
53 10 9 10 0 1 15 1 9 9 10 9 13 3 1 9 12 2 16 13 1 15 1 12 9 3 2 16 13 1 15 9 1 10 9 10 15 2 7 16 10 9 13 1 9 15 14 10 9 11 11 11 0 2
24 13 1 15 2 7 15 1 13 3 10 9 16 13 9 13 13 1 15 7 13 14 9 15 2
37 13 3 9 2 16 1 9 15 14 9 15 1 10 9 2 13 1 9 15 14 10 9 1 9 15 7 0 2 7 10 12 3 13 13 1 15 2
12 15 13 16 15 13 3 1 9 1 9 0 2
35 15 13 1 15 3 2 16 12 1 10 9 16 13 14 15 13 1 15 3 14 10 9 16 15 4 13 1 9 15 9 9 1 10 9 2
19 15 3 13 2 16 15 3 3 13 9 1 9 16 4 13 1 15 9 2
47 13 1 15 3 1 9 10 9 11 2 1 9 16 13 13 15 1 10 11 2 7 13 1 15 13 9 0 3 1 10 9 10 15 2 7 13 13 9 1 10 16 13 1 9 1 9 2
13 15 13 2 1 9 3 0 14 9 2 15 13 2
6 3 13 1 15 13 2
10 3 13 13 9 1 10 9 10 15 2
17 15 13 10 9 10 0 16 13 14 15 13 1 9 1 10 15 2
11 3 2 15 13 9 3 0 1 9 15 2
24 10 9 14 15 13 2 3 13 3 16 15 4 1 10 9 10 15 2 7 3 9 1 9 2
69 15 13 1 9 16 1 9 12 2 16 13 1 10 11 7 13 9 10 9 10 0 1 15 1 9 2 13 2 3 1 9 15 2 9 11 2 9 0 1 11 11 2 16 1 15 13 10 9 11 13 1 9 14 9 1 10 9 16 15 13 13 1 9 0 14 12 9 11 2
57 7 13 1 15 2 1 15 9 9 10 9 13 16 3 2 13 2 1 11 2 16 15 13 7 9 2 7 1 10 15 13 10 9 10 0 10 15 1 11 2 1 9 16 13 0 1 10 9 16 15 13 1 9 15 14 11 2
15 10 9 1 9 2 3 13 1 11 7 3 13 1 15 2
14 15 10 9 10 0 10 0 1 3 13 9 1 11 2
11 15 13 13 2 3 3 1 15 10 9 2
6 10 9 7 9 15 2
17 11 11 13 1 9 12 10 9 10 0 3 1 10 9 10 0 2
42 9 15 2 9 15 7 9 15 13 1 9 0 1 9 10 9 7 11 2 7 10 9 10 0 3 13 1 13 1 15 3 1 16 10 9 10 0 13 13 1 15 2
16 1 12 13 11 10 9 10 0 16 13 1 9 9 2 0 2
29 9 15 14 2 11 2 9 2 3 2 11 11 2 13 16 4 1 9 15 13 1 10 9 10 0 9 14 9 2
9 9 15 1 11 3 13 0 3 2
22 15 13 13 1 11 1 9 1 9 11 2 7 1 10 9 0 10 9 14 15 9 2
21 1 11 4 13 2 3 2 13 14 3 16 13 13 1 10 9 10 0 14 11 2
54 9 15 13 3 9 9 2 7 7 3 1 9 0 14 15 1 9 11 2 1 10 9 2 11 2 11 2 2 13 10 9 16 11 13 1 9 9 10 9 1 9 10 9 2 2 15 13 14 3 16 9 13 2 2
20 2 11 2 11 2 13 7 13 3 2 1 10 9 2 14 10 9 10 0 2
14 11 13 1 15 1 10 9 16 15 13 13 14 15 2
30 15 13 9 7 13 3 16 10 9 13 14 10 9 2 7 13 1 15 9 16 13 13 1 9 15 7 1 9 15 2
27 2 1 9 13 15 13 14 3 16 13 1 15 10 9 7 14 3 16 13 1 15 9 2 2 13 11 2
18 7 10 9 10 0 13 1 15 2 2 7 3 1 15 13 9 2 2
20 7 11 13 1 9 2 2 7 7 15 4 13 14 15 1 9 1 3 2 2
18 11 13 1 9 15 13 1 9 2 12 7 13 3 13 1 9 15 2
16 15 13 13 14 9 9 10 9 7 13 1 15 1 9 0 2
16 9 15 1 10 9 7 1 9 10 9 1 11 13 3 9 2
11 7 1 9 0 0 13 1 9 15 9 2
47 3 13 1 15 9 0 3 1 9 9 15 14 10 9 10 0 2 1 1 15 16 10 1 9 10 9 10 0 10 0 9 10 9 13 1 10 9 13 1 15 1 10 9 1 10 11 2
20 1 9 15 4 13 9 15 13 1 9 0 3 14 10 9 10 0 10 0 2
14 9 0 14 9 1 12 10 9 16 13 15 14 15 2
38 1 10 9 10 0 7 1 10 9 11 13 15 3 16 10 9 14 15 13 16 16 13 9 11 9 15 14 11 2 7 9 15 14 10 9 10 0 2
39 7 2 1 1 9 14 9 1 9 10 9 2 9 10 9 1 10 9 1 10 9 13 14 9 2 9 1 9 10 9 16 10 9 10 0 3 4 13 2
33 9 1 9 15 14 11 2 1 9 7 1 9 9 1 10 9 10 0 2 16 9 15 0 7 3 0 7 10 9 13 14 15 2
33 3 16 13 3 14 10 9 1 10 9 10 0 13 10 9 2 16 1 10 9 10 0 10 0 9 1 9 13 9 0 1 11 2
43 1 9 11 13 15 3 1 9 15 10 0 3 14 11 11 1 10 9 2 1 16 3 2 13 9 0 0 13 14 15 1 9 0 1 9 10 9 1 9 2 10 9 2
25 9 10 9 2 16 4 1 10 9 10 0 1 11 2 13 4 13 16 9 1 9 11 13 3 2
14 3 9 9 0 2 3 9 9 2 7 3 9 9 2
30 10 9 3 13 15 2 7 10 9 16 13 1 9 11 1 9 10 9 7 1 9 10 9 1 10 9 13 0 3 2
26 7 9 13 1 12 9 16 9 1 11 13 1 3 2 3 3 4 11 13 9 1 16 9 3 13 2
32 10 9 14 9 9 1 10 9 2 16 15 3 10 9 10 0 1 10 10 9 16 13 9 10 9 13 1 9 1 9 15 2
34 1 10 9 13 1 10 9 10 0 10 9 0 2 1 9 15 9 0 10 3 10 9 1 10 9 1 9 1 9 1 11 7 11 2
71 9 12 13 9 0 0 2 2 11 13 1 15 3 3 10 9 9 2 2 7 9 0 12 13 13 14 9 15 14 10 9 1 10 9 0 2 10 9 7 13 1 10 9 10 0 2 2 1 10 3 10 9 13 9 7 1 11 14 15 2 3 13 14 15 1 9 0 1 9 2 2
35 9 10 9 15 13 1 10 0 7 1 10 0 1 9 0 2 14 15 13 14 9 10 9 3 1 9 15 7 1 9 15 14 10 9 2
33 9 0 2 3 9 2 13 3 16 1 10 9 2 3 1 9 15 10 0 2 13 1 10 9 14 15 3 10 9 0 1 9 2
21 13 16 11 9 13 14 10 9 1 9 9 1 9 1 13 1 9 15 10 0 2
31 7 3 10 9 2 13 16 15 13 9 0 7 9 0 3 2 13 1 10 9 15 1 13 9 7 9 2 3 0 3 2
71 9 10 9 1 9 0 13 3 9 0 2 3 0 2 3 13 14 9 10 9 1 9 12 2 11 11 2 16 13 1 15 3 1 11 9 9 1 10 9 14 10 0 13 16 15 13 13 14 10 9 1 10 9 16 13 14 10 9 14 9 11 1 9 11 9 0 1 2 1 3 2
16 1 9 9 1 9 16 13 1 15 12 9 0 4 3 13 2
31 3 1 10 9 2 16 12 1 15 13 9 3 0 1 9 10 9 1 9 16 9 15 13 2 9 9 2 10 9 2 2
26 3 10 9 10 0 10 15 13 13 1 9 15 14 9 10 9 1 10 9 1 9 15 13 10 9 2
80 1 10 9 0 10 9 16 15 13 1 9 15 2 1 9 9 10 9 14 2 11 10 9 2 2 3 15 9 13 2 2 2 3 13 1 9 16 15 13 3 1 16 15 0 2 2 7 4 13 2 1 9 10 9 10 0 2 7 13 2 2 7 9 3 13 1 15 7 3 2 1 0 9 2 7 1 13 9 2 2
31 3 0 3 13 14 10 9 15 1 9 16 13 1 9 11 2 7 16 13 3 10 9 1 10 9 16 13 10 9 11 2
6 7 1 15 3 13 2
66 10 16 9 10 9 10 15 2 7 16 9 10 10 10 9 7 15 2 13 0 7 13 1 15 16 10 9 13 3 1 15 7 1 3 16 15 13 2 3 13 15 16 3 13 2 7 3 3 13 0 1 15 16 10 9 13 1 10 9 10 0 7 1 9 3 2
6 9 13 1 10 9 2
18 1 3 13 9 15 13 11 9 4 13 0 1 9 13 2 7 0 2
29 15 7 15 2 10 9 16 15 13 1 10 9 2 7 3 10 9 1 10 9 2 13 9 10 9 7 10 9 2
15 9 9 9 13 9 10 9 2 10 9 7 9 10 9 2
35 3 3 13 13 11 11 2 7 1 9 15 13 13 13 7 9 0 7 3 13 10 3 1 11 11 2 9 9 9 1 9 1 9 15 2
22 3 1 9 15 3 13 2 3 3 1 9 10 9 2 3 3 16 16 13 1 9 2
43 1 11 1 9 0 2 9 16 13 3 16 16 13 2 9 0 1 15 7 1 11 2 2 2 4 13 9 1 10 9 2 15 9 2 1 9 10 9 10 3 2 0 2
47 15 16 13 14 9 15 10 0 7 10 9 4 13 1 15 2 7 16 15 13 14 10 9 10 0 14 15 1 9 9 15 16 15 2 1 9 9 2 15 16 13 14 15 1 10 9 2
47 7 16 13 15 9 15 1 9 9 3 2 0 2 1 9 9 2 10 9 16 13 3 2 7 1 10 9 10 0 1 9 2 10 9 10 0 10 0 14 10 9 10 3 2 0 2 2
9 13 15 9 3 13 2 13 2 2
32 7 3 4 3 13 3 2 13 9 13 7 1 10 9 1 10 15 2 14 10 13 1 9 9 2 7 1 10 9 0 15 2
65 13 1 15 9 15 14 10 9 10 0 11 9 2 9 15 14 11 9 2 16 3 13 2 3 2 1 9 9 1 9 2 2 1 9 15 14 11 11 2 2 10 9 16 9 14 9 0 13 15 10 9 10 0 10 0 3 1 9 15 13 14 9 15 2 2
18 1 15 4 13 13 2 3 7 3 9 14 9 0 13 1 9 15 2
39 7 10 9 10 0 3 13 2 7 13 1 9 15 14 10 10 9 2 10 9 16 0 9 1 2 10 9 10 0 3 2 14 9 0 13 1 9 15 2
28 3 2 3 3 13 13 10 9 16 9 0 12 13 3 1 10 10 0 2 7 3 2 1 10 9 10 0 2
47 9 0 2 0 14 15 13 1 9 15 14 11 1 9 9 1 9 1 9 15 2 2 3 2 3 3 13 14 15 3 1 11 11 2 2 10 9 2 3 2 1 10 9 2 3 2 2
29 7 13 1 9 10 9 2 16 1 15 9 9 10 9 13 1 9 0 2 1 10 13 7 1 10 9 1 12 2
20 10 9 4 13 0 7 0 2 7 13 1 9 15 3 1 10 9 10 0 2
42 3 9 1 10 9 10 0 1 9 0 1 10 9 10 0 11 11 10 0 2 16 7 13 1 2 10 9 10 0 0 2 10 9 3 13 1 15 14 10 9 2 2
39 10 9 15 7 9 14 10 9 10 3 2 0 2 7 10 0 2 7 3 13 9 2 0 2 3 1 11 2 2 13 16 15 13 14 10 9 10 15 2
46 7 16 3 13 15 13 3 10 9 13 1 15 16 9 10 9 1 10 9 10 9 13 4 13 1 9 13 11 1 2 9 9 9 0 12 3 13 13 1 15 7 13 1 15 3 2
14 2 9 0 2 2 13 11 2 2 13 0 2 2 2
14 3 13 10 9 10 0 7 9 15 3 1 9 15 2
75 7 2 9 0 1 9 15 13 1 10 9 10 0 1 10 9 10 0 1 11 2 16 13 3 10 9 16 1 15 13 1 9 10 9 2 15 9 1 10 13 10 9 10 0 10 0 4 1 15 2 2 3 13 9 12 14 15 1 15 16 1 10 9 13 1 15 1 9 16 11 13 1 10 9 2
35 2 3 13 1 15 7 13 15 2 7 15 13 15 1 9 15 7 7 13 2 10 9 13 13 1 9 16 3 13 1 15 11 2 2 2
25 3 7 3 2 9 15 14 11 13 3 1 10 9 10 0 14 10 9 16 10 9 13 1 15 2
58 3 13 16 9 15 0 3 1 9 13 1 15 11 2 11 7 11 1 15 16 13 9 1 11 11 11 7 11 11 2 3 13 9 0 0 16 3 13 1 9 2 7 3 3 16 16 13 1 15 9 2 1 9 9 9 15 0 2
22 7 1 9 12 13 3 15 1 9 1 10 9 10 0 15 2 2 10 0 3 2 2
25 10 9 13 16 13 2 0 3 2 7 3 16 15 0 1 10 9 10 0 2 10 3 2 0 2
33 3 2 10 10 9 10 15 14 9 13 0 2 0 2 7 0 1 9 15 14 10 9 2 1 9 0 3 16 0 1 9 15 2
39 13 14 10 9 16 13 16 9 16 13 1 9 9 13 4 13 0 3 2 7 16 13 1 10 9 9 0 3 1 1 10 9 10 0 2 10 0 3 2
34 7 1 9 12 3 2 4 1 10 9 3 2 7 1 9 9 3 2 16 9 15 13 9 3 1 10 9 10 11 11 11 7 9 2
19 4 9 2 0 1 15 2 7 16 13 1 9 15 7 13 1 9 15 2
14 7 7 3 13 13 2 3 3 3 9 14 9 0 2
30 7 13 9 0 2 3 2 0 2 1 9 1 9 2 9 15 14 9 15 3 1 10 9 10 0 16 1 10 9 2
20 13 2 3 2 1 10 15 16 13 9 0 1 9 15 14 10 9 10 0 2
71 9 12 14 15 2 16 9 15 13 13 1 15 9 1 9 9 2 15 13 1 9 0 0 1 9 0 0 2 7 3 13 10 1 3 13 15 1 9 15 2 2 13 1 9 9 9 2 9 2 2 10 9 10 0 10 0 3 2 1 13 14 10 9 10 0 16 13 1 10 9 2
14 2 3 13 1 9 2 2 15 13 1 15 3 9 2
5 2 3 3 13 2
5 2 2 15 13 2
13 2 7 7 13 13 1 9 0 15 13 3 0 2
16 2 2 13 9 15 10 0 2 1 10 9 16 13 3 9 2
28 15 15 9 1 10 9 16 7 3 11 13 14 9 11 3 13 14 15 9 0 16 9 15 13 1 10 15 2
21 3 7 3 2 9 10 9 3 3 13 13 14 10 9 1 11 7 3 3 3 2
8 7 1 9 9 11 13 0 2
17 11 1 9 9 0 1 9 11 2 3 3 1 10 9 10 0 2
28 1 9 10 9 13 9 2 16 1 9 1 9 10 9 10 9 2 0 13 13 9 1 11 1 9 1 9 2
29 13 3 9 1 9 1 11 16 13 9 1 9 2 9 2 7 9 9 1 11 16 13 1 9 9 1 9 0 2
11 12 1 12 10 9 16 13 3 1 11 2
25 1 9 9 15 10 0 15 13 1 10 9 10 0 1 13 1 10 9 2 16 13 14 10 9 2
20 2 3 1 16 13 11 11 2 2 13 11 11 1 9 15 1 1 12 9 2
33 11 2 16 13 1 11 1 12 9 2 7 3 9 15 1 12 9 13 1 11 7 1 9 15 2 13 1 9 15 1 9 0 2
35 3 12 9 9 13 1 15 3 1 11 2 7 1 9 10 9 13 3 1 10 9 12 1 9 15 2 2 13 14 10 9 10 12 2 2
14 10 9 1 2 11 2 11 11 9 11 2 13 0 2
35 10 9 2 1 12 0 2 1 9 9 15 2 2 2 9 1 11 2 7 2 13 1 15 1 11 2 13 1 9 15 14 11 1 11 2
32 10 9 13 13 1 10 9 14 10 9 10 0 2 14 9 10 9 14 11 2 7 3 14 9 2 9 14 9 9 10 12 2
47 3 16 13 11 11 1 11 2 11 7 11 11 1 11 14 9 15 2 13 13 1 10 9 10 0 1 11 3 9 0 2 0 1 9 2 16 13 1 10 9 10 9 2 0 14 3 2
33 1 10 1 9 15 14 11 13 9 16 13 1 15 9 0 16 4 13 15 7 1 10 15 13 13 15 2 9 10 9 2 0 2
54 9 2 9 14 9 10 9 10 0 1 11 2 14 9 10 9 7 10 9 1 11 2 14 10 9 1 9 2 14 10 9 10 0 7 10 9 2 14 9 10 9 14 10 9 7 10 9 10 0 1 9 10 9 2
30 10 15 13 3 1 2 13 14 10 9 10 12 2 2 9 0 1 12 9 0 16 13 1 11 1 9 9 10 12 2
21 10 12 13 13 9 7 9 2 7 10 9 9 13 1 10 9 2 9 1 11 2
42 10 12 2 16 13 4 7 13 13 13 1 9 0 2 13 14 9 15 1 9 1 9 0 0 1 9 10 9 14 9 2 9 7 11 7 1 9 10 11 1 11 2
18 10 9 10 0 13 14 10 9 2 7 9 15 10 9 13 14 15 2
9 1 9 10 9 15 13 1 9 2
61 2 13 14 10 9 10 12 2 2 7 1 9 1 10 9 10 0 2 13 14 10 9 1 10 12 2 2 2 13 1 9 0 14 9 2 3 15 13 1 9 0 2 1 7 16 10 9 13 14 9 9 2 3 13 1 10 9 9 14 9 2
56 10 9 2 13 1 2 9 9 0 1 9 10 9 10 12 7 1 9 15 1 9 0 2 13 1 9 0 9 16 13 15 13 1 10 9 10 0 10 0 2 16 1 15 7 1 15 2 13 1 15 9 1 10 12 2 2
33 15 3 10 9 16 3 16 15 13 1 9 9 9 15 15 13 4 13 1 9 15 13 14 15 2 7 13 13 1 9 10 9 2
24 1 1 10 9 15 14 11 11 2 3 1 10 9 10 15 13 1 10 10 9 9 0 0 2
50 15 13 1 12 1 11 2 2 9 9 15 2 2 2 16 3 13 1 9 2 2 13 1 9 1 9 1 9 16 13 1 12 1 9 15 2 2 7 16 1 9 15 13 9 7 9 10 9 2 2
15 1 9 0 15 13 13 1 9 13 7 13 14 9 15 2
28 1 9 12 13 3 14 9 10 9 7 13 13 1 9 9 2 13 9 2 13 9 1 10 9 7 9 9 2
21 1 9 3 0 13 1 9 2 1 9 10 9 14 10 9 7 1 9 10 9 2
18 10 15 0 13 9 9 16 13 14 15 1 9 7 13 1 9 15 2
24 1 15 2 11 13 13 7 13 3 2 7 1 9 15 10 0 4 13 9 14 9 0 0 2
26 1 9 12 13 11 11 1 10 9 10 0 14 11 2 1 9 9 1 9 16 13 3 1 10 15 2
47 15 13 1 10 9 10 0 3 1 11 10 0 2 7 13 1 10 9 14 2 11 2 11 2 2 1 9 7 3 1 10 9 2 2 9 0 16 13 1 9 15 1 9 0 2 9 2
26 11 11 13 3 1 9 0 2 16 13 14 9 15 3 3 1 9 0 7 3 1 9 9 7 9 2
73 9 9 15 10 0 2 2 9 0 1 10 9 2 2 7 10 9 10 0 14 15 2 2 10 9 10 12 14 10 9 2 2 16 13 9 1 12 2 9 0 9 7 9 1 11 10 3 2 0 2 13 9 1 9 10 9 7 1 10 9 10 0 14 10 9 10 0 1 10 9 10 0 2
29 9 0 7 0 13 0 3 1 10 9 16 13 1 10 9 10 0 2 7 13 13 1 9 9 15 7 1 9 2
43 1 10 9 13 1 15 14 10 13 10 0 1 10 9 14 10 9 2 10 0 10 13 2 1 11 2 16 13 1 9 9 7 9 3 2 0 14 10 9 16 16 15 2
34 2 10 9 10 12 14 10 9 2 13 1 12 9 2 7 1 9 2 1 12 2 13 1 9 0 16 13 1 9 10 9 1 11 2
8 1 11 3 13 3 12 9 2
32 10 9 10 0 2 10 9 7 10 9 1 9 10 9 10 0 14 11 13 13 2 7 1 1 9 10 9 13 13 9 0 2
49 9 10 2 9 2 10 0 2 16 1 11 12 13 1 10 9 14 11 11 2 3 13 9 0 2 7 10 9 7 10 9 14 10 9 10 0 13 7 13 14 9 15 10 0 1 9 10 9 2
10 10 9 13 9 15 1 9 7 9 2
54 1 7 16 1 10 9 15 1 15 9 3 13 11 14 10 9 10 0 7 14 10 9 14 10 9 10 0 2 7 13 13 1 10 9 10 0 2 3 4 13 10 9 13 14 9 15 10 0 7 10 3 2 0 2
64 9 15 10 0 2 9 15 10 0 7 9 10 9 10 0 14 15 1 10 9 2 16 13 1 15 14 9 10 9 2 13 3 16 13 1 15 14 9 9 15 14 10 9 10 0 7 3 14 10 9 10 0 2 16 13 15 13 9 10 9 14 10 9 2
67 11 10 9 7 10 9 2 11 10 9 10 13 2 16 13 14 9 10 9 1 9 10 9 10 0 7 14 9 10 9 1 9 10 9 10 0 2 13 1 3 1 9 1 10 9 14 11 2 7 14 13 1 12 1 9 1 10 9 15 13 14 10 9 13 1 15 2
26 10 9 10 0 1 9 13 14 15 2 9 0 2 2 7 13 14 15 1 2 9 9 7 0 2 2
53 7 3 1 10 13 1 15 9 15 14 10 9 7 10 9 13 1 9 12 9 0 2 2 10 9 2 7 2 10 9 10 0 9 11 2 2 1 7 10 9 16 12 1 15 13 3 3 1 10 15 1 9 2
38 1 10 9 15 7 9 15 13 11 14 12 10 9 1 9 2 10 9 0 10 9 2 11 2 2 9 3 0 14 10 9 10 3 2 0 1 11 2
25 1 9 10 9 13 9 1 9 1 10 9 2 7 3 1 9 10 9 10 0 2 9 0 9 2
16 15 13 13 14 9 10 9 14 15 2 7 13 16 13 3 2
16 11 13 16 7 13 2 15 13 7 13 1 15 13 7 13 2
33 1 7 16 13 16 2 10 3 16 3 13 1 11 7 13 13 1 15 13 13 14 15 2 2 13 13 1 10 9 1 13 9 2
32 7 10 9 3 13 2 7 15 13 15 13 1 11 1 11 2 1 11 2 1 9 11 2 7 3 2 1 9 12 1 11 2
7 3 13 13 3 1 3 2
8 10 9 1 9 1 15 0 2
25 10 12 13 16 15 13 1 2 9 9 15 11 11 2 9 9 7 9 0 16 13 1 10 9 2
50 11 2 9 9 2 10 9 2 1 9 2 9 7 3 9 1 9 11 2 11 2 13 1 15 16 2 11 13 1 10 9 1 16 1 10 9 13 9 11 2 10 9 10 0 14 15 1 11 2 2
39 9 0 13 11 11 2 16 13 9 15 14 11 1 9 9 1 11 7 12 1 9 15 10 0 1 11 2 2 11 13 1 11 16 13 1 2 9 11 2
32 10 9 1 9 0 11 11 13 1 15 9 9 2 7 13 1 11 16 13 1 10 9 2 7 1 10 9 10 9 13 2 2
24 3 7 3 2 11 10 3 2 0 13 13 1 11 9 0 1 10 9 10 0 1 9 15 2
24 12 12 9 13 1 10 9 12 14 11 1 9 0 2 7 13 3 9 9 0 1 9 0 2
30 9 2 9 2 9 2 9 7 9 16 13 1 11 13 14 10 9 10 0 1 9 11 1 9 15 10 0 2 0 2
15 7 10 9 16 13 11 11 1 15 3 13 1 9 15 2
16 15 13 15 13 9 3 2 7 13 13 7 13 1 9 13 2
31 15 13 1 11 1 9 0 14 9 15 11 11 1 10 9 14 11 1 11 9 2 1 9 1 9 9 7 1 9 9 2
30 15 7 4 13 13 1 2 11 2 1 10 9 1 10 9 10 0 2 7 7 1 9 15 3 13 1 9 10 9 2
16 1 9 15 13 13 1 9 7 13 3 2 7 10 9 13 2
21 7 13 1 10 9 16 13 2 2 0 9 10 12 2 2 15 13 3 9 9 2
17 2 15 3 0 16 1 11 15 13 9 9 2 2 13 11 11 2
45 9 0 13 11 1 9 15 14 11 2 7 3 1 2 15 2 14 13 13 1 9 2 11 2 7 1 9 2 11 2 1 11 2 13 10 12 13 9 1 9 9 7 1 9 2
8 2 11 13 3 9 14 9 2
7 15 13 13 16 15 0 2
4 16 15 9 2
11 15 13 9 7 3 3 13 1 10 9 2
26 3 1 16 13 14 10 9 9 1 11 11 13 1 3 11 13 14 10 9 7 14 10 9 14 15 2
7 15 13 13 14 11 11 2
16 15 13 0 2 0 2 0 9 7 9 13 2 13 1 15 2
9 7 11 13 13 0 7 13 2 2
34 12 1 15 9 1 9 15 3 10 9 16 1 9 15 13 11 11 2 9 1 9 11 11 2 16 1 9 15 13 12 1 9 15 2
14 10 9 1 15 13 1 9 9 1 9 1 12 9 2
30 14 13 11 14 11 2 13 11 14 10 9 7 13 1 9 1 2 11 2 9 2 1 16 4 13 15 3 1 9 2
9 3 1 11 13 1 9 14 9 2
34 15 13 14 15 1 9 2 7 3 1 9 7 1 9 2 1 9 14 9 9 2 9 16 13 1 9 10 9 10 0 7 9 0 2
50 3 10 3 16 13 1 15 13 11 1 9 1 9 15 2 10 9 16 1 9 15 2 9 15 11 11 7 9 15 2 9 10 9 1 9 2 11 2 2 9 9 2 9 9 2 9 0 7 9 2
28 1 7 10 9 16 13 7 13 1 9 15 1 9 2 9 2 13 9 15 1 9 15 14 9 9 2 9 2
52 10 9 7 10 9 10 0 9 10 9 1 2 11 2 7 10 9 16 3 12 9 14 15 13 1 11 2 2 10 9 10 12 1 10 9 2 7 9 1 9 1 2 10 9 10 15 2 2 13 14 15 2
17 1 9 14 9 2 1 9 15 14 15 2 2 13 1 15 2 2
16 15 13 1 9 15 14 11 11 2 7 1 12 13 14 11 2
35 14 11 2 9 0 2 13 3 1 11 1 12 14 13 1 10 9 10 0 1 9 1 9 9 15 2 10 9 10 12 14 10 9 2 2
13 2 15 13 9 1 9 0 2 2 13 11 11 2
13 2 1 10 9 10 0 1 9 13 11 1 11 2
25 11 2 16 3 13 11 2 13 1 10 9 2 13 1 15 16 15 13 13 1 15 1 10 9 2
6 10 9 13 7 13 2
18 11 13 1 9 15 7 13 14 15 1 10 9 1 9 10 9 2 2
13 1 15 13 9 15 2 7 10 9 1 15 13 2
37 14 13 1 11 11 1 9 15 10 0 14 9 15 15 13 1 11 2 13 1 10 9 2 11 2 2 7 1 1 9 9 13 14 15 1 15 2
15 11 2 16 13 9 2 13 9 2 15 3 13 1 11 2
27 10 9 13 1 9 1 11 2 7 14 9 15 2 1 9 15 14 11 2 15 13 1 11 11 1 11 2
11 7 10 9 7 10 9 3 13 9 0 2
32 14 10 9 15 1 16 13 1 10 9 10 0 7 1 10 9 14 9 10 9 7 14 9 15 1 11 2 13 1 9 15 2
16 13 15 7 0 7 0 1 9 15 16 10 9 3 13 9 2
20 10 12 13 2 7 1 3 13 11 11 13 7 10 9 13 3 1 9 0 2
8 11 13 13 14 15 7 13 2
32 3 2 1 9 9 15 14 9 15 1 11 2 10 9 7 10 9 11 11 2 13 1 9 2 10 9 7 13 1 11 11 2
14 1 11 13 9 0 16 4 13 1 11 1 9 9 2
9 7 3 13 10 9 1 9 15 2
24 9 9 0 16 11 13 9 9 1 9 15 13 1 11 9 2 15 7 10 9 7 9 15 2
15 11 13 1 10 9 2 7 3 9 15 13 1 9 15 2
23 3 2 1 9 15 2 2 9 1 11 2 2 13 10 9 2 9 14 9 15 1 9 2
28 3 10 9 10 0 7 11 13 14 11 2 13 1 15 7 13 1 10 2 11 9 2 14 15 13 7 13 2
11 9 15 10 0 7 10 0 13 7 13 2
33 1 9 15 13 13 1 9 9 2 7 1 3 1 3 13 9 1 9 0 1 9 0 16 2 13 15 2 1 11 2 11 11 2
23 10 15 9 15 13 7 13 16 13 1 15 2 11 2 11 2 2 16 4 13 1 11 2
15 15 7 13 9 1 9 1 11 7 1 9 0 1 15 2
53 1 9 15 10 0 1 11 11 16 3 13 14 15 13 16 13 1 15 3 9 1 15 2 7 15 13 12 12 9 7 13 9 1 10 9 1 13 14 10 9 1 9 9 1 9 15 7 9 15 14 10 9 2
24 2 3 10 9 2 2 13 10 9 2 9 0 16 13 1 9 2 10 9 2 14 11 11 2
8 2 13 10 9 2 2 13 2
11 1 9 10 12 13 11 1 11 12 9 2
19 1 10 9 10 12 2 1 12 2 13 1 15 9 13 1 15 1 9 2
26 15 13 3 1 9 14 9 2 1 13 1 9 2 1 9 9 15 2 1 2 9 10 9 10 0 2
10 10 9 10 0 13 13 9 7 0 2
20 1 10 9 13 1 15 9 9 1 11 11 16 13 3 15 2 1 11 11 2
11 3 13 11 16 13 13 14 11 1 9 2
20 15 13 1 11 13 9 0 1 9 1 10 9 2 7 13 13 3 1 11 2
21 7 1 12 1 11 12 15 13 0 1 9 15 1 9 15 14 10 9 10 0 2
7 9 12 13 1 9 15 2
9 1 9 15 13 9 9 1 11 2
14 1 9 15 13 9 14 9 11 16 13 9 7 13 2
15 2 9 2 2 13 11 11 2 2 11 13 1 9 9 2
6 9 15 13 13 9 2
11 15 13 9 7 3 9 9 1 9 2 2
32 15 13 1 9 9 0 1 11 2 7 1 9 15 13 9 15 13 2 11 11 9 13 9 0 7 9 13 1 15 9 2 2
14 9 13 1 15 9 13 9 12 1 9 15 10 0 2
50 11 11 2 9 9 11 2 11 2 11 16 13 3 1 3 1 9 15 2 13 1 9 15 2 16 13 9 1 9 1 10 9 2 7 13 16 9 2 9 13 13 3 7 16 13 1 15 10 9 2
14 7 1 15 13 3 10 10 9 16 15 4 1 15 2
25 10 9 3 13 1 10 3 16 10 9 10 0 4 13 2 3 1 9 10 9 10 0 14 15 2
22 1 9 16 1 15 9 2 9 11 7 9 9 13 14 9 15 2 3 4 1 9 2
27 15 3 12 10 9 16 3 9 7 9 0 7 3 0 16 13 13 1 9 1 9 0 0 10 2 3 2
36 13 1 15 10 9 10 0 11 11 2 16 1 9 9 3 15 13 9 2 0 1 10 9 2 1 10 9 2 9 9 7 9 7 9 9 2
24 1 9 15 13 1 9 0 11 11 2 16 13 2 3 1 11 2 3 9 1 9 10 9 2
23 7 3 12 15 13 3 2 7 9 15 13 9 10 9 10 0 2 10 0 7 10 0 2
45 3 10 9 13 1 9 15 2 13 1 15 9 15 10 0 2 9 15 7 9 10 9 10 0 14 15 2 7 10 9 16 1 10 9 0 7 0 7 0 2 15 13 9 0 2
21 10 9 13 3 13 9 2 3 3 1 10 9 16 13 1 15 9 14 9 0 2
95 1 10 9 0 9 0 1 9 9 2 7 15 16 13 2 7 2 11 11 2 10 9 10 0 2 16 13 1 15 7 1 9 15 1 9 0 2 13 9 0 2 0 9 2 13 1 9 16 13 14 9 10 9 7 3 14 9 10 9 2 9 16 3 13 1 9 14 10 9 10 0 2 14 10 9 2 14 10 9 2 16 13 14 10 9 1 9 16 13 1 10 9 10 0 2
36 3 3 16 13 10 9 0 1 9 0 2 7 10 12 13 9 1 9 2 9 2 7 16 16 13 0 3 2 3 13 9 15 13 1 9 2
26 11 11 7 11 11 9 0 7 0 7 9 9 9 0 2 16 13 1 9 9 10 0 13 1 0 2
24 1 10 9 16 13 7 1 10 9 16 13 14 15 2 0 16 13 10 9 7 9 1 9 2
14 15 13 13 1 15 9 16 13 1 15 14 10 9 2
44 11 13 1 9 1 10 2 9 2 2 16 15 3 9 1 11 11 2 7 1 9 0 0 1 9 0 2 7 11 13 13 10 9 10 0 2 10 9 2 10 9 10 0 2
10 3 15 13 13 1 9 0 2 0 2
23 1 10 9 10 0 14 15 15 13 1 10 10 9 14 10 9 10 0 7 10 0 3 2
31 1 16 10 0 7 10 13 13 7 13 1 9 15 14 9 0 2 3 9 15 13 15 2 7 9 15 0 9 7 9 2
16 7 7 13 3 7 3 15 3 1 10 9 7 9 10 9 2
39 4 13 13 16 10 9 2 9 11 2 10 0 10 2 3 2 13 9 9 7 9 9 0 1 10 9 10 0 7 10 0 2 7 10 9 0 7 0 2
37 11 11 16 13 13 14 9 10 9 13 1 9 0 2 7 13 10 9 16 15 13 1 2 9 9 0 3 2 7 13 1 9 15 1 9 0 2
3 0 3 2
19 11 11 13 3 3 15 13 14 13 16 2 3 9 0 1 10 9 2 2
10 3 16 9 15 14 11 13 1 15 2
20 1 9 10 9 13 13 1 9 15 3 9 0 7 0 1 10 9 10 0 2
27 3 13 1 9 15 14 11 11 2 9 10 9 2 7 13 3 13 1 15 10 9 0 16 13 1 15 2
11 3 13 9 15 1 9 2 15 3 13 2
36 7 7 1 13 1 9 2 9 11 4 13 11 13 13 1 9 0 0 2 9 9 0 7 9 0 2 0 7 9 14 13 1 9 9 9 2
24 7 3 15 13 14 11 11 16 13 9 0 7 0 2 7 13 1 0 9 7 9 2 9 2
12 4 13 16 13 3 16 16 4 1 10 9 2
12 1 10 9 10 9 13 11 11 7 11 11 2
29 12 9 10 9 1 9 11 16 3 13 4 13 16 13 13 1 15 9 1 14 15 3 13 1 10 9 7 13 2
21 10 9 10 0 14 15 1 10 9 10 12 13 1 9 0 2 0 7 0 9 2
21 13 16 3 14 15 13 10 9 10 0 10 0 2 7 7 15 13 1 15 9 2
33 3 10 9 13 1 9 9 2 1 10 15 16 4 13 13 3 1 11 11 2 7 11 11 2 7 3 13 3 1 9 10 9 2
24 3 7 9 10 9 13 14 10 3 16 13 14 15 1 15 2 3 13 1 15 9 0 3 2
16 3 1 9 15 14 2 9 9 2 13 14 15 9 14 9 2
31 7 3 15 13 7 10 9 13 11 11 2 16 13 14 9 15 10 0 2 7 11 11 16 13 13 3 1 9 9 15 2
22 10 9 10 15 13 9 0 16 3 13 14 15 2 7 9 14 9 1 9 0 0 2
30 3 0 10 9 10 0 2 16 13 1 0 1 9 7 1 9 2 7 10 9 15 13 1 9 1 9 1 10 9 2
23 7 16 3 10 9 10 0 2 10 0 2 1 2 9 10 9 2 13 3 14 10 9 2
23 9 11 1 10 9 10 12 13 9 13 1 10 9 1 9 2 7 16 1 9 14 9 2
51 13 16 10 9 13 2 1 9 9 2 0 1 9 7 3 3 1 9 2 9 0 1 9 15 14 10 9 2 7 1 10 9 16 1 15 11 11 2 16 13 13 14 10 9 1 9 9 3 2 0 2
21 7 3 15 4 13 13 7 9 15 10 0 14 10 0 1 9 16 1 10 9 2
17 3 3 16 15 13 14 9 15 2 7 15 3 9 9 9 0 2
27 7 7 7 13 9 0 2 10 9 10 0 7 9 10 9 13 1 15 9 0 16 13 1 9 14 9 2
26 10 9 2 3 3 16 15 13 13 14 10 9 2 9 2 2 13 7 15 13 14 10 9 10 15 2
24 13 1 15 3 9 13 14 15 1 9 0 2 1 16 10 9 13 1 9 0 7 13 9 2
19 3 7 2 9 11 10 0 16 9 15 13 9 16 13 9 0 7 0 2
11 9 16 13 1 9 14 9 0 2 0 2
33 9 15 13 1 0 3 3 1 15 2 7 3 1 10 9 10 0 2 10 0 2 16 9 15 9 0 1 10 9 7 10 9 2
37 1 11 13 13 1 9 0 9 0 2 0 16 0 1 9 1 9 15 1 10 9 0 2 7 1 15 13 14 15 1 0 2 7 7 1 0 2
25 13 4 13 1 10 9 10 0 16 13 9 16 13 1 9 1 11 2 7 13 16 3 15 3 2
12 7 3 3 13 1 13 7 13 9 1 15 2
31 10 9 14 15 0 1 9 10 9 10 0 2 15 13 1 9 0 14 9 9 2 7 1 15 15 13 1 10 9 15 2
22 10 9 13 1 10 9 10 0 7 10 0 16 9 15 0 2 7 15 3 4 13 2
23 4 13 1 9 16 13 1 9 7 9 15 13 1 10 9 2 14 15 13 14 9 15 2
11 13 3 10 9 10 0 7 9 10 9 2
51 1 9 0 13 1 9 15 10 0 16 13 1 15 1 9 14 9 9 1 9 0 0 2 7 10 9 13 1 9 10 9 15 13 1 9 15 14 11 2 11 2 11 2 7 1 10 9 14 11 11 2
16 13 16 13 9 0 7 9 9 0 1 13 9 0 2 0 2
28 7 1 15 9 10 9 13 1 9 10 9 2 7 10 9 10 0 10 0 16 15 13 13 15 14 10 9 2
14 3 16 15 15 13 10 9 0 3 0 1 9 9 2
16 11 13 13 1 11 2 9 2 1 9 9 1 9 10 9 2
24 11 7 11 13 1 11 11 1 10 9 10 3 0 1 9 2 16 13 1 11 2 11 12 2
21 3 13 11 1 9 0 9 1 9 9 14 10 9 10 0 1 10 9 10 0 2
31 9 10 9 2 9 11 2 11 11 13 3 2 2 13 1 15 3 13 1 15 2 16 3 3 13 1 15 9 9 2 2
24 10 9 10 0 1 9 15 14 11 13 3 10 9 1 9 1 15 9 10 9 10 3 0 2
27 11 13 4 13 14 10 9 2 7 11 13 16 1 10 9 1 10 9 13 3 1 11 3 13 10 9 2
22 10 9 11 13 2 16 9 9 10 9 13 3 1 16 13 7 10 9 13 1 11 2
30 10 9 11 13 16 9 10 9 13 1 10 0 14 11 2 7 10 9 3 13 1 10 9 1 9 9 1 10 9 2
23 3 13 3 9 15 14 11 13 1 11 1 13 1 9 10 9 2 11 2 14 9 15 2
16 10 9 13 14 11 1 2 12 1 11 1 9 3 9 11 2
14 11 13 1 9 10 9 1 9 15 1 11 12 12 2
7 1 9 15 13 3 11 2
40 11 13 4 13 1 9 9 1 9 11 7 11 1 9 10 9 2 7 13 1 9 11 16 13 1 11 1 9 2 7 13 16 9 11 3 3 13 1 11 2
42 3 2 1 9 11 1 10 9 2 10 9 1 16 13 1 9 14 11 11 2 13 9 9 9 9 0 1 9 10 9 14 9 2 11 2 1 11 7 13 9 13 2
80 1 9 10 9 14 11 11 16 13 1 9 9 2 1 9 0 16 13 1 9 9 1 9 10 9 7 1 10 9 16 13 1 15 1 9 9 0 16 13 9 14 9 16 4 13 1 9 15 2 1 15 16 1 3 7 3 4 1 10 9 13 3 1 15 2 12 7 12 9 1 9 2 16 16 9 4 13 1 15 2
8 9 0 14 9 13 1 15 2
25 15 13 1 9 2 13 1 9 15 9 1 10 9 2 13 3 3 14 9 15 2 7 3 13 2
9 12 9 0 13 1 15 9 9 2
14 15 3 13 2 7 15 13 1 3 16 13 9 0 2
36 16 13 1 10 9 16 13 14 10 9 7 13 14 9 15 2 13 10 9 1 15 9 7 9 2 2 9 1 15 2 14 15 4 13 2 2
24 10 12 13 1 9 1 10 9 16 3 2 7 13 1 9 9 16 13 0 1 9 10 9 2
21 3 2 1 10 9 10 12 14 10 9 2 1 9 2 11 2 2 13 9 9 2
16 9 13 14 15 13 1 15 14 9 10 9 2 7 13 3 2
8 13 1 15 16 13 1 9 2
24 1 10 9 3 13 13 9 7 1 15 9 9 10 9 16 4 13 1 9 15 14 10 9 2
29 12 10 9 13 9 9 9 2 3 1 9 10 9 10 0 2 16 16 13 9 15 14 10 9 11 1 9 15 2
27 7 3 13 10 9 11 1 9 15 14 9 15 1 3 16 13 1 9 12 1 0 9 15 14 9 11 2
20 7 3 2 11 13 1 10 9 7 0 9 0 1 10 9 16 13 1 15 2
21 15 13 1 15 3 9 2 9 2 9 16 13 14 9 15 1 9 9 10 9 2
57 3 13 11 1 9 11 11 2 16 13 1 15 1 12 9 1 9 9 15 14 10 9 10 0 1 10 9 2 16 10 9 10 0 16 1 15 15 13 9 13 11 10 9 2 1 15 15 13 1 10 9 7 13 1 10 9 2
9 1 9 15 11 11 13 3 9 2
32 1 9 15 13 1 9 11 1 10 9 2 2 9 15 2 13 1 15 9 2 2 7 14 9 9 15 13 1 9 10 11 2
52 11 13 16 16 13 1 11 1 9 9 15 10 0 2 13 1 15 9 2 11 2 1 9 14 3 16 10 9 10 0 0 1 15 2 2 15 9 15 2 3 15 13 2 15 3 16 0 1 9 15 13 2
15 3 16 15 13 15 10 9 10 0 3 14 10 9 2 2
39 1 9 15 2 9 3 0 1 9 0 2 13 3 3 7 3 3 2 16 7 9 9 11 13 13 3 2 13 15 2 11 2 10 9 10 0 14 11 2
22 15 13 16 1 9 15 4 13 1 1 9 11 11 11 1 9 16 13 14 10 9 2
20 1 9 2 11 2 13 9 9 0 2 7 13 14 15 1 9 0 1 9 2
15 15 13 7 13 1 9 10 9 1 9 10 9 10 0 2
35 10 9 10 13 13 9 10 9 2 13 2 7 3 7 15 15 13 1 9 10 9 13 9 0 1 9 11 7 9 15 3 13 1 9 2
71 11 13 14 9 10 9 1 9 0 13 7 13 2 1 10 9 10 0 16 1 15 15 13 1 10 9 2 9 11 13 14 15 1 1 9 9 15 2 1 9 15 14 10 2 9 11 7 11 13 7 13 1 9 11 2 10 9 13 1 9 15 2 13 1 9 7 13 1 9 0 2
30 1 16 13 2 3 3 16 15 4 13 9 1 9 2 9 7 13 1 9 15 9 16 1 15 15 13 1 9 11 2
13 15 7 13 13 1 9 1 10 9 1 9 15 2
17 1 9 0 3 13 11 11 14 15 1 13 9 15 14 11 11 2
18 9 15 13 1 10 9 2 13 10 9 2 7 3 1 9 10 9 2
16 3 3 13 13 1 9 15 14 10 9 16 1 15 13 13 2
11 1 9 15 10 0 7 10 0 13 0 2
12 1 9 15 7 1 9 15 13 14 11 11 2
36 16 13 11 1 10 9 1 12 13 11 2 2 3 3 13 1 15 9 9 0 2 2 7 13 14 10 9 10 0 1 2 9 10 9 2 2
18 1 9 2 16 13 9 11 2 11 2 13 1 15 9 15 9 0 2
50 15 13 1 11 9 16 13 1 9 15 7 1 9 15 2 7 1 9 1 2 11 11 2 13 16 9 10 9 13 1 2 9 10 9 2 1 15 16 10 9 14 15 1 10 9 13 1 9 10 2
23 11 13 1 10 9 10 3 0 14 10 9 10 0 1 13 1 15 14 9 15 10 0 2
56 1 15 13 1 10 9 16 13 1 9 0 2 9 9 9 9 7 9 0 13 1 9 15 14 9 10 9 13 9 1 9 0 16 13 1 9 15 9 1 9 1 10 9 10 0 2 7 1 9 9 0 1 9 9 0 2
30 10 9 2 13 10 9 11 9 2 13 1 10 9 9 16 13 1 15 9 1 9 10 9 7 1 10 9 1 9 2
30 11 13 1 9 14 9 10 9 1 10 9 2 7 13 1 15 9 16 13 1 15 9 1 9 0 7 0 0 3 2
22 3 13 1 9 15 9 9 7 9 0 3 13 1 15 14 9 15 7 14 9 15 2
21 9 15 1 10 11 1 12 13 1 9 9 15 1 9 1 9 1 9 9 15 2
38 1 10 9 14 11 12 2 16 9 9 10 9 13 1 15 9 14 12 1 12 9 2 13 9 15 16 9 9 13 14 9 15 1 9 9 10 9 2
64 15 13 13 16 9 10 9 13 14 9 15 14 2 11 2 1 10 9 2 7 16 11 13 1 9 9 16 13 1 15 13 9 0 3 1 10 9 2 1 11 7 1 10 9 2 11 7 9 15 3 13 9 1 15 2 2 7 2 13 14 9 10 9 2
25 9 9 16 13 14 9 9 15 14 11 13 9 1 10 9 2 7 13 9 0 1 2 11 2 2
16 10 9 13 1 9 15 14 10 9 7 9 15 10 0 13 2
32 9 15 13 7 13 3 1 9 14 13 9 2 0 2 4 13 2 1 9 2 1 9 7 1 9 1 9 9 0 1 9 2
15 11 11 13 1 2 11 2 16 13 1 15 9 14 9 2
14 11 13 10 9 10 0 16 1 9 15 13 10 9 2
20 15 13 10 9 2 9 10 9 2 10 9 7 10 9 10 0 14 10 9 2
12 15 13 9 14 9 7 9 1 9 10 9 2
35 15 2 7 9 0 2 13 16 2 11 2 3 13 3 3 9 14 10 9 1 11 2 7 9 3 2 0 1 9 15 7 1 9 15 2
14 11 13 0 7 13 14 9 15 10 0 1 9 0 2
37 7 13 1 10 9 10 0 1 15 9 1 11 11 2 11 11 7 11 11 2 16 13 9 0 0 1 15 16 1 15 13 10 9 2 11 2 2
25 7 7 15 13 9 9 15 2 3 13 1 15 13 9 2 7 1 9 13 9 2 11 2 3 2
36 1 2 11 2 3 9 9 9 9 9 1 9 15 14 9 10 9 10 0 2 7 13 1 15 9 9 9 0 1 9 15 14 9 9 9 2
28 13 1 10 9 9 0 14 3 2 7 10 9 15 13 0 1 9 12 7 0 1 15 7 1 9 9 15 2
10 1 9 15 13 11 9 0 7 13 2
22 15 13 9 0 2 7 13 13 16 16 13 9 15 13 9 9 1 10 9 16 13 2
21 13 1 15 9 0 2 15 13 14 9 15 1 10 9 10 0 16 1 10 9 2
11 3 13 3 1 10 9 1 9 1 11 2
42 1 10 9 13 9 1 9 10 9 2 7 13 13 1 10 9 9 16 3 9 1 10 9 13 1 15 2 7 13 13 13 14 15 2 1 1 10 9 10 0 2 2
11 15 13 1 9 0 1 10 9 10 0 2
30 1 9 14 15 1 9 11 2 7 2 13 1 9 0 1 15 16 10 9 13 1 15 14 10 9 1 9 15 3 2
10 15 13 9 1 9 10 9 3 0 2
11 3 9 0 1 9 15 13 14 9 15 2
33 3 3 13 9 10 9 14 9 15 10 0 2 9 9 10 9 13 9 1 9 9 15 1 9 16 9 15 13 1 9 9 15 2
6 11 13 1 9 15 2
29 1 12 9 13 1 9 15 10 0 2 2 10 9 2 2 14 10 9 2 7 13 16 10 9 10 0 13 3 2
40 3 13 1 15 1 10 9 10 0 9 16 13 13 1 9 3 0 7 13 14 9 10 9 14 15 2 7 13 14 9 9 15 2 7 3 3 14 9 15 2
38 3 2 3 1 3 2 3 2 4 9 0 2 1 9 13 7 13 2 13 14 9 15 14 11 11 2 2 0 1 9 15 15 13 16 15 13 2 2
15 1 9 11 3 13 9 15 14 9 11 11 1 9 0 2
57 1 9 10 9 10 0 14 10 9 2 1 9 10 9 14 9 10 9 10 0 2 13 9 11 11 7 9 0 9 11 1 9 9 7 1 9 2 7 13 1 15 9 0 7 9 1 9 14 12 9 9 2 1 12 9 2 2
15 7 9 15 10 0 13 10 9 13 14 10 9 1 9 2
48 9 15 14 9 11 11 3 13 1 9 10 9 16 1 15 13 10 9 2 7 3 13 1 9 15 14 10 9 3 2 9 11 11 2 9 13 11 11 2 9 2 7 9 2 9 11 11 2
76 1 9 9 9 1 10 9 2 9 11 11 2 1 10 9 2 9 11 11 7 9 11 11 2 13 1 9 10 9 10 0 10 9 16 1 9 16 1 15 13 12 10 9 1 9 10 9 1 9 13 9 2 9 9 12 2 9 1 12 2 16 13 1 15 9 14 9 10 9 10 0 1 9 9 11 2
24 3 1 9 10 9 10 0 3 13 3 16 1 9 1 10 9 14 10 12 13 9 11 11 2
13 13 3 16 15 13 1 9 0 7 16 9 13 2
25 12 10 9 10 0 7 10 0 14 11 7 11 13 1 9 9 1 10 9 10 0 1 10 9 2
55 15 13 13 14 10 9 1 9 15 10 0 2 7 13 1 10 9 16 9 9 11 13 16 3 2 4 13 14 12 10 9 1 9 0 1 9 2 16 16 13 9 13 16 10 9 16 13 1 15 13 16 13 14 11 2
56 1 9 3 0 14 9 2 16 1 15 13 10 9 14 9 15 2 13 12 10 9 1 9 2 9 10 9 13 13 1 15 10 9 16 13 14 9 15 14 11 7 13 16 10 9 16 13 10 12 3 13 1 9 9 9 2
16 3 13 9 16 13 14 10 12 1 3 2 9 1 10 9 2
37 3 13 9 13 1 9 10 9 7 10 9 10 0 16 3 13 9 16 3 13 13 14 10 9 16 1 15 9 11 11 2 13 14 9 15 2 2
43 13 10 9 1 9 9 15 14 10 9 2 16 13 9 1 9 13 1 9 9 1 9 9 10 9 16 13 1 10 9 2 7 1 9 0 1 9 10 9 7 10 9 2
14 11 13 1 2 9 10 9 2 2 12 1 11 12 2
32 16 13 2 13 9 11 16 13 0 1 9 1 9 10 9 16 13 1 9 9 1 9 9 15 2 7 16 9 9 15 13 2
21 16 13 1 9 15 2 1 9 2 13 9 11 1 10 9 16 9 9 15 13 2
33 3 9 7 9 1 1 3 2 9 10 9 10 0 1 2 10 9 2 1 10 9 2 13 9 11 13 16 11 13 14 10 9 2
15 16 13 13 1 10 9 2 13 16 9 11 13 9 0 2
21 11 3 3 13 14 10 9 16 16 13 0 1 15 9 9 10 9 7 3 9 2
13 3 13 9 11 16 9 15 1 9 15 13 9 2
23 13 1 9 9 10 9 7 15 13 2 1 9 2 16 10 9 13 1 9 9 10 9 2
31 16 13 9 9 9 10 9 2 13 9 9 10 9 13 2 10 9 14 15 3 13 14 10 9 7 13 13 1 15 3 2
19 9 9 10 9 13 9 0 2 10 9 13 1 9 9 10 9 10 0 2
7 1 10 9 13 9 0 2
85 13 9 16 10 9 16 13 1 10 9 13 1 13 14 9 15 14 9 11 11 2 16 3 13 9 1 10 9 2 3 13 0 1 9 0 15 2 13 1 10 9 16 13 10 9 10 0 2 0 1 16 4 13 1 9 9 15 10 0 2 15 13 9 9 1 9 2 2 13 1 9 9 15 14 15 7 9 9 15 13 14 9 9 15 2
60 10 9 10 15 13 14 13 16 9 16 13 9 11 11 2 9 15 14 9 10 9 2 1 9 9 10 9 3 2 11 11 2 11 2 3 13 3 2 7 16 9 14 9 11 11 7 14 11 11 2 9 15 14 11 2 3 13 7 15 2
15 3 9 10 9 1 2 10 9 2 13 14 10 9 13 2
37 10 9 10 0 13 9 0 14 9 9 10 9 1 9 9 10 9 10 0 13 1 9 9 11 9 13 1 9 12 9 9 10 9 1 9 11 2
9 10 9 1 9 9 2 9 13 2
29 15 13 7 13 3 16 13 16 9 10 9 13 16 13 1 9 15 10 9 1 13 14 9 15 14 12 10 9 2
9 15 13 13 15 1 9 0 3 2
22 3 13 16 9 9 10 9 3 13 15 1 9 0 13 0 7 13 1 9 0 15 2
37 3 10 9 10 0 13 1 10 9 7 1 10 9 2 1 9 2 9 1 10 9 1 10 9 7 9 0 14 9 10 9 2 1 9 9 15 2
38 10 9 10 0 13 9 10 9 16 13 10 9 10 0 2 16 1 9 15 3 13 1 9 10 9 9 16 13 13 1 9 9 9 2 9 1 9 2
8 7 3 15 9 9 1 0 2
24 1 15 2 1 9 10 13 13 9 15 10 0 14 10 9 1 10 9 10 0 14 10 9 2
23 9 15 14 9 0 13 1 9 1 9 9 0 14 10 9 1 9 1 9 9 1 9 2
55 3 16 13 3 1 9 1 9 3 2 1 9 9 9 15 2 2 13 9 9 1 9 9 9 1 9 2 16 13 9 14 9 1 9 1 12 9 0 2 16 13 1 9 9 0 16 1 15 13 9 1 9 10 9 2
33 2 1 9 10 9 13 10 9 1 9 1 9 10 9 2 2 13 10 9 7 10 9 13 3 1 9 10 9 1 9 10 9 2
18 9 4 13 9 1 10 9 1 9 10 9 10 2 12 14 10 11 2
41 12 10 9 13 3 1 10 9 1 9 0 2 10 13 11 11 2 12 9 2 13 14 11 2 13 12 2 7 11 2 12 9 2 13 1 11 2 9 12 2 2
21 11 11 4 13 14 9 15 10 12 2 3 1 15 12 9 2 7 13 1 11 2
22 10 10 9 2 11 11 11 2 11 11 2 11 11 11 2 11 11 11 2 11 11 2
5 3 2 11 11 2
30 3 13 13 1 10 9 2 16 10 9 14 11 13 10 9 10 0 3 1 10 9 10 0 7 3 7 3 1 15 2
29 12 10 9 1 9 10 9 2 10 9 7 11 2 13 1 9 11 1 9 10 9 1 10 0 7 3 13 15 2
16 11 2 16 9 15 13 11 11 2 13 1 9 14 12 9 2
39 9 0 15 13 15 1 9 10 9 1 9 0 1 10 9 10 9 9 9 7 11 9 9 2 11 9 11 7 11 11 2 10 0 16 13 14 11 2 2
27 10 9 11 2 1 9 10 9 11 2 11 2 11 2 13 3 1 10 9 10 2 12 7 3 3 13 2
27 7 10 9 1 10 9 4 13 3 1 9 10 9 1 10 9 10 0 2 1 10 9 10 0 12 2 2
22 10 9 1 11 1 10 9 10 13 3 13 3 1 9 0 7 13 3 1 9 15 2
12 12 9 13 7 10 9 3 13 3 1 11 2
16 9 10 9 13 3 12 16 10 9 14 11 13 1 9 15 2
20 1 9 11 4 13 10 9 10 0 11 11 2 16 13 1 9 9 10 9 2
12 11 13 1 10 9 10 0 1 10 9 11 2
18 13 0 1 9 14 11 13 10 9 10 0 7 13 10 9 11 11 2
22 1 9 10 9 9 0 1 9 10 9 11 11 7 11 11 2 7 10 9 3 0 2
19 9 10 9 9 9 13 1 9 9 14 11 1 13 1 10 9 10 0 2
24 7 3 1 9 15 14 11 11 13 1 10 9 1 11 11 16 3 1 15 9 1 10 9 2
24 11 9 11 2 16 13 12 2 13 3 14 11 11 16 13 1 9 15 14 10 9 11 11 2
9 9 11 9 2 3 1 10 9 2
19 3 11 9 9 9 1 9 10 9 16 13 3 1 11 1 10 9 11 2
28 1 9 9 13 3 9 9 2 16 1 15 13 10 9 10 0 14 10 9 9 10 9 2 9 10 9 2 2
21 1 11 13 3 2 12 2 11 10 0 7 10 9 11 16 13 13 1 9 9 2
23 11 9 11 2 16 13 1 10 9 10 0 9 9 2 13 1 10 9 1 10 9 11 2
11 11 11 13 14 10 9 10 0 11 11 2
35 13 10 9 9 2 3 10 9 7 10 13 16 1 15 2 16 13 1 9 7 10 9 13 7 4 13 13 9 7 3 7 1 10 9 2
20 15 13 9 1 10 9 2 7 1 15 13 9 0 7 13 13 1 10 9 2
28 3 13 3 9 15 14 9 10 9 1 9 11 11 13 1 9 9 2 16 13 1 10 9 10 0 1 11 2
35 9 15 1 9 15 14 10 1 9 10 9 16 13 1 10 9 2 16 9 15 13 1 9 9 7 9 9 2 0 3 7 3 13 3 2
29 9 15 3 3 13 9 15 1 10 9 2 7 13 7 13 14 10 9 10 0 14 9 10 9 1 10 10 9 2
15 9 9 10 9 1 9 13 7 13 14 10 9 1 11 2
24 9 15 10 0 14 11 2 16 13 13 1 9 15 9 0 2 13 1 9 14 9 9 0 2
39 3 16 0 1 1 10 9 2 9 15 14 10 9 1 11 3 13 0 3 2 7 0 3 2 1 9 15 7 3 9 15 14 11 1 10 9 10 12 2
28 7 3 16 3 0 2 9 9 10 9 1 9 3 13 3 0 2 7 1 9 13 11 14 9 15 1 11 2
17 1 9 9 10 12 13 13 16 10 9 13 1 11 11 10 0 2
17 1 9 12 13 3 1 10 9 9 10 9 7 13 9 3 0 2
67 1 13 14 9 10 9 1 10 9 2 13 14 10 9 7 13 14 10 9 1 10 9 10 0 2 15 13 9 13 2 9 2 13 9 0 1 9 10 9 2 13 7 13 10 9 1 10 9 2 13 9 0 2 13 9 9 7 13 9 9 0 1 10 9 10 0 2
38 9 10 9 10 0 7 9 10 9 10 0 3 3 13 1 9 1 16 13 1 9 10 9 2 3 13 3 9 0 2 0 14 9 15 14 11 11 2
35 1 10 9 16 13 2 1 9 0 1 12 9 9 2 13 9 11 2 11 1 9 10 9 2 7 13 1 10 9 14 10 9 10 0 2
17 10 9 2 10 9 10 0 10 0 14 9 10 9 13 9 0 2
43 1 3 13 10 9 1 9 9 10 12 13 11 11 1 9 0 2 10 9 10 0 3 16 3 13 2 7 9 10 9 13 1 12 9 9 14 10 10 9 1 9 15 2
12 3 13 10 9 2 7 3 1 9 10 9 2
52 10 9 2 11 2 13 16 10 9 10 0 13 16 9 11 11 13 0 2 7 3 0 3 2 15 13 1 13 1 9 0 16 1 15 3 13 10 9 2 7 9 10 9 2 10 9 7 10 9 10 0 2
68 1 9 15 3 13 9 2 9 10 9 13 0 1 16 13 2 10 9 13 1 9 0 1 9 9 7 1 10 9 1 10 9 1 9 10 9 2 7 10 9 10 0 13 13 9 0 1 9 7 9 1 10 9 1 9 10 9 7 9 15 2 1 9 1 9 10 9 2
24 4 13 16 10 9 10 0 10 0 13 1 9 10 9 2 15 13 1 15 9 1 10 9 2
24 7 7 1 9 15 15 3 13 13 1 10 9 16 13 10 9 10 0 1 9 9 10 9 2
22 0 3 13 14 9 10 9 16 13 1 10 9 10 0 1 9 1 9 10 9 3 2
36 9 1 15 2 1 10 9 10 0 13 1 10 9 10 0 9 9 1 9 14 12 9 2 9 16 4 13 13 15 1 10 9 1 10 9 2
21 3 9 10 9 13 3 1 9 0 1 10 9 16 13 1 10 9 1 1 12 2
117 10 9 1 10 9 13 14 10 9 1 10 9 10 0 1 9 9 1 12 7 9 10 9 10 0 1 9 0 2 1 9 2 2 1 10 9 10 0 10 9 3 15 3 16 3 13 2 7 13 1 10 9 10 0 3 1 1 10 9 1 10 9 10 0 1 10 9 2 10 9 1 9 10 9 10 0 13 1 9 7 9 2 2 7 1 9 15 13 10 9 10 0 9 1 9 9 0 1 10 9 10 0 1 9 15 1 12 7 1 12 2 3 1 11 12 2 2
16 9 15 13 0 1 12 9 2 9 10 9 7 9 10 9 2
17 10 9 7 9 1 9 10 9 1 10 9 10 0 13 1 15 2
16 9 9 0 1 9 7 9 13 9 9 10 9 1 9 0 2
26 9 9 16 13 13 1 9 13 1 9 1 9 0 3 0 2 7 4 13 3 1 9 3 2 0 2
28 13 10 9 1 9 9 9 16 13 1 10 9 10 0 1 9 0 2 3 0 2 1 9 0 0 1 0 2
35 13 10 9 16 10 9 4 13 14 10 9 10 0 1 10 9 2 16 16 15 0 13 14 10 9 10 0 1 9 2 9 7 9 9 2
28 7 13 13 3 2 13 1 9 15 10 9 14 9 10 9 10 0 1 9 9 10 9 1 10 9 10 0 2
41 10 9 1 9 9 10 9 13 3 13 1 10 9 7 3 9 1 10 9 2 7 9 1 1 9 2 10 9 14 9 0 7 9 10 9 1 10 9 14 15 2
11 0 1 15 10 9 1 10 9 10 0 2
11 10 9 13 1 9 15 9 0 1 15 2
64 1 9 16 1 15 13 3 3 12 9 0 2 7 10 4 13 12 9 0 2 13 10 9 10 0 13 1 9 15 14 9 15 10 0 2 16 13 3 12 7 12 1 10 9 10 0 1 10 9 2 12 9 1 9 7 3 2 2 7 7 13 1 15 2
23 10 9 10 3 13 13 2 16 9 10 9 13 7 13 1 9 9 0 1 9 10 9 2
49 10 9 1 9 10 9 7 1 9 0 3 2 10 9 10 0 16 13 1 9 1 10 9 14 10 9 2 10 13 13 10 9 10 0 3 1 9 10 9 14 9 10 9 1 10 9 10 0 2
19 1 11 11 15 13 14 10 9 2 1 15 15 4 13 3 14 10 9 2
14 3 13 1 10 9 10 0 9 0 2 3 0 9 2
20 12 9 13 1 12 1 12 9 15 14 9 11 1 10 9 14 9 10 9 2
53 0 9 11 2 2 11 11 2 2 13 1 9 16 10 9 2 16 15 4 13 1 9 16 1 15 10 9 13 9 0 2 3 1 9 12 2 14 10 9 2 13 9 16 4 13 9 0 1 10 10 9 2 2
45 1 9 10 9 13 1 15 12 10 9 2 10 9 10 0 11 11 2 13 14 10 9 10 0 10 15 1 0 3 2 16 13 13 14 10 9 16 15 9 0 3 1 9 15 2
35 15 13 1 15 13 14 9 15 10 0 1 10 9 14 9 0 7 14 9 0 7 3 1 10 9 14 9 11 2 7 3 14 9 3 2
13 9 11 3 13 0 2 7 15 13 14 9 15 2
34 7 16 11 13 7 13 1 10 9 2 3 1 3 2 1 9 9 7 1 9 9 10 9 2 15 4 3 1 10 9 10 0 3 2
42 9 15 1 10 9 1 11 13 1 9 15 14 9 10 9 10 0 10 0 2 16 10 9 10 0 7 10 0 10 15 4 13 13 1 10 9 16 1 9 15 13 2
22 1 12 9 15 1 10 9 13 11 10 9 10 0 3 14 11 1 10 9 10 0 2
22 9 0 13 1 9 10 9 2 13 1 9 0 0 1 9 7 13 1 15 1 9 2
13 1 11 13 13 1 15 16 15 2 9 0 2 2
7 7 11 13 3 9 0 2
16 16 16 13 9 15 1 11 2 3 13 9 15 1 9 15 2
39 1 12 15 13 1 9 9 10 9 10 0 1 10 9 2 7 3 13 3 16 13 4 13 1 10 9 13 3 14 10 9 10 0 11 11 1 11 11 2
23 11 3 13 3 9 10 9 10 0 10 0 2 7 1 10 9 15 9 10 9 10 0 2
18 3 13 9 0 3 1 10 9 11 1 9 9 0 1 10 9 11 2
7 9 15 13 3 0 3 2
24 7 1 12 13 11 13 14 9 15 2 7 14 9 15 14 9 0 0 2 1 3 2 0 2
32 15 13 2 7 2 9 1 9 0 1 9 11 2 7 13 1 15 13 1 10 9 10 0 10 0 1 10 9 2 11 11 2
13 1 11 3 13 3 9 1 10 9 7 1 11 2
30 1 9 10 9 10 0 14 15 15 13 3 14 9 15 14 9 15 2 7 14 9 15 10 0 2 0 14 9 15 2
26 15 3 13 1 11 2 1 9 9 1 10 9 2 11 11 2 2 13 9 1 11 1 9 9 15 2
44 9 9 1 2 11 2 2 11 11 2 13 1 9 1 10 9 2 1 10 9 2 0 1 9 2 15 13 1 10 9 10 0 2 1 9 0 2 2 7 0 1 9 2 2
67 1 9 11 3 2 9 1 10 9 1 10 9 1 11 2 13 10 9 2 11 11 2 1 11 2 16 9 10 9 14 11 13 1 12 9 1 10 9 9 2 16 13 9 0 1 9 15 10 0 14 10 9 10 0 2 9 0 2 9 7 9 16 9 15 11 11 2
35 1 10 9 2 1 9 9 10 9 14 11 2 13 9 15 14 11 1 10 9 10 0 2 7 3 9 15 10 3 2 0 14 9 15 2
27 11 2 7 7 13 1 12 1 9 0 1 9 10 9 14 11 11 2 3 13 1 10 9 1 9 11 2
13 15 13 16 13 13 1 11 11 7 1 11 11 2
41 15 10 0 13 10 9 10 0 10 0 2 16 13 14 9 11 1 9 15 1 12 2 16 13 14 10 9 2 9 9 2 7 13 14 11 1 2 9 0 2 2
57 11 13 2 1 15 2 1 10 9 1 2 9 14 10 9 2 2 9 1 12 9 14 9 7 9 0 1 9 10 9 10 0 2 16 13 3 9 12 9 7 9 1 10 9 10 0 1 11 2 1 13 14 15 1 9 9 2
20 15 13 9 2 0 3 1 9 15 14 9 2 1 9 10 9 14 11 11 2
30 11 3 3 13 1 10 9 13 3 1 9 15 12 9 0 7 1 9 10 9 14 15 15 13 1 15 14 9 15 2
10 16 13 10 9 13 1 11 9 13 2
18 1 15 15 3 13 2 16 2 10 9 13 1 9 1 10 9 2 2
12 1 11 15 13 14 10 9 2 9 10 15 2
18 1 11 9 2 9 1 10 9 16 13 11 13 9 14 9 2 9 2
24 0 1 9 15 13 1 11 1 9 0 14 9 9 0 1 10 9 7 1 10 9 10 0 2
27 12 10 9 10 0 3 14 10 9 13 15 16 13 1 9 14 9 14 9 2 10 9 2 9 0 2 2
29 16 0 13 13 1 9 0 1 9 2 15 13 14 15 1 9 2 13 1 9 0 2 2 7 2 9 11 2 2
17 1 9 10 9 13 3 9 1 14 15 13 1 9 1 10 15 2
22 11 2 16 13 1 10 9 1 9 14 12 9 1 9 10 9 2 13 1 9 11 2
15 9 0 1 11 13 9 0 1 10 9 7 1 10 9 2
37 3 9 13 16 9 0 1 11 10 0 2 16 9 15 10 0 13 9 10 9 10 0 2 13 14 10 9 10 0 14 15 1 9 10 3 0 2
45 11 13 1 9 0 1 9 9 2 1 9 15 13 3 4 13 14 10 9 1 10 9 10 0 1 9 7 9 0 2 13 2 7 0 7 16 3 3 13 7 13 7 13 9 2
12 1 9 9 10 9 13 10 9 2 9 13 2
45 7 3 13 2 3 10 9 10 3 2 0 1 11 13 9 0 2 7 9 15 14 10 9 10 0 2 16 15 11 11 2 13 9 1 11 1 9 1 9 9 1 9 10 9 2
29 10 9 0 3 1 10 9 9 10 9 2 11 13 1 9 10 9 2 13 15 1 9 10 9 9 14 11 11 2
51 7 10 9 11 2 7 7 13 1 9 9 3 2 10 9 11 2 13 9 10 9 3 1 3 16 13 14 10 9 2 9 1 9 15 14 11 1 9 7 9 9 1 1 10 1 9 10 9 10 0 2
37 1 9 10 9 2 9 7 9 9 2 1 9 16 13 10 9 10 0 14 10 9 2 3 4 13 1 9 14 9 2 7 16 15 0 9 3 2
39 0 9 3 13 10 4 13 1 9 9 2 13 1 9 0 7 1 10 9 1 10 15 3 16 7 13 14 11 11 13 14 9 10 9 1 9 10 9 2
22 13 16 10 9 13 1 9 15 16 13 14 10 9 11 13 9 0 1 11 1 11 2
18 7 3 2 1 9 16 1 15 13 10 9 13 3 2 0 1 9 2
26 7 9 10 9 14 9 11 2 7 3 9 15 7 9 15 2 4 3 1 9 1 10 9 10 0 2
34 3 11 13 13 9 13 1 9 9 2 3 15 3 13 13 13 1 9 15 13 9 1 9 9 2 1 13 9 9 9 0 7 0 2
38 7 3 3 10 9 11 11 2 7 13 10 9 3 11 11 2 13 16 11 13 9 16 4 13 1 9 2 7 3 13 1 15 9 15 9 1 15 2
13 7 3 3 13 1 9 10 9 1 11 10 9 2
15 7 7 2 9 10 9 1 10 9 13 1 9 3 13 2
25 11 13 11 2 7 1 13 7 11 13 3 13 13 3 13 10 9 10 0 1 9 9 10 12 2
30 13 9 16 9 1 9 16 1 15 13 9 9 1 9 13 1 14 15 2 7 13 14 10 9 1 10 9 10 0 2
8 9 15 13 2 3 1 9 2
33 10 9 11 11 2 9 10 9 10 0 16 13 1 11 2 13 16 2 10 9 16 1 9 15 4 13 14 11 1 10 9 2 2
38 7 7 15 13 9 2 1 9 16 13 1 9 0 1 2 11 11 11 2 2 3 15 13 2 13 14 9 9 10 9 1 9 0 1 10 9 2 2
24 4 16 10 9 1 9 16 0 1 0 1 10 9 10 0 13 3 1 9 11 1 9 9 2
40 7 3 15 10 9 2 7 12 1 15 2 16 11 13 3 2 0 13 14 10 9 2 16 1 9 9 15 10 0 10 9 11 13 16 15 4 13 1 15 2
74 3 15 9 16 9 10 9 11 2 7 9 0 16 15 13 3 3 2 13 9 10 9 10 0 1 9 10 9 2 7 16 3 0 1 15 9 15 13 13 1 9 12 14 10 9 2 9 7 9 2 8 1 9 14 9 2 1 10 9 2 9 11 1 11 7 9 9 10 9 1 9 15 2 2
6 7 11 13 10 0 2
45 3 3 16 13 10 9 11 2 2 15 13 16 13 9 0 1 9 1 11 2 1 9 15 14 9 10 9 1 9 15 2 7 1 9 9 1 13 9 7 9 1 10 9 2 2
21 7 3 2 9 1 10 15 0 2 7 1 0 9 13 0 16 9 13 1 9 2
29 7 16 11 13 1 10 9 1 9 9 2 16 7 13 4 13 13 3 14 10 9 10 3 2 13 1 10 9 2
13 15 9 15 14 10 9 10 0 9 2 9 15 2
33 9 15 14 11 7 10 9 13 1 9 9 1 10 9 10 9 3 13 1 9 9 2 1 9 9 2 13 14 11 1 9 15 2
52 7 16 13 1 9 15 10 0 1 10 9 16 15 4 13 3 3 7 3 13 1 11 1 11 11 7 9 15 2 4 16 10 9 13 13 1 9 15 2 7 3 7 9 10 9 13 13 13 1 12 9 2
60 7 1 9 11 4 13 1 15 1 3 13 14 10 9 1 9 15 2 7 1 9 15 14 3 9 13 1 10 9 9 2 16 1 9 9 10 9 16 13 1 9 15 13 1 9 15 10 0 14 10 9 10 9 1 9 10 9 10 12 2
32 3 9 9 2 7 3 9 0 1 10 9 2 7 1 12 10 7 10 3 9 1 9 9 2 13 4 1 9 1 10 15 2
42 1 16 9 10 9 2 1 9 10 9 11 2 3 13 1 15 14 10 9 1 10 9 2 3 15 13 1 10 9 10 0 2 2 13 9 15 14 9 15 14 11 2
20 10 15 13 1 9 16 16 3 13 13 1 12 9 9 16 13 1 9 15 2
34 1 10 9 13 9 9 14 10 9 10 0 10 0 1 11 9 9 14 9 9 10 9 1 9 16 13 1 9 15 1 9 10 9 2
25 1 9 7 9 0 13 9 10 9 1 9 15 14 9 10 9 10 0 13 14 10 9 10 0 2
18 10 9 13 13 3 13 9 14 9 1 9 2 7 13 1 9 0 2
45 9 12 10 9 16 13 1 15 14 10 9 13 2 16 10 9 1 9 9 9 0 3 10 1 3 16 13 1 15 9 10 9 10 0 16 13 1 15 9 9 0 1 9 11 2
41 7 1 9 15 13 10 9 3 13 14 9 15 1 9 15 14 10 9 2 7 13 1 9 7 1 9 10 9 14 10 9 0 10 9 16 13 1 9 9 0 2
19 3 3 13 10 9 1 9 15 14 9 10 9 10 0 2 10 9 11 2
19 1 9 15 10 12 14 10 9 13 10 9 11 1 9 15 7 1 15 2
12 9 9 15 3 13 14 9 15 1 10 9 2
20 15 13 1 9 10 9 1 9 11 2 11 2 11 7 3 4 13 13 9 2
9 2 13 1 9 15 2 2 13 2
28 2 3 13 9 10 9 14 11 11 16 10 9 13 14 10 9 1 13 14 9 15 14 10 9 10 0 2 2
7 1 15 9 13 10 9 2
25 15 13 1 9 15 14 9 9 10 9 1 10 9 10 0 7 10 9 1 9 9 0 1 9 2
34 4 3 13 1 2 9 2 16 13 1 10 9 10 0 2 10 0 2 14 11 2 16 1 15 9 9 9 15 0 1 9 10 9 2
56 4 13 1 10 9 10 0 1 10 9 2 9 9 10 9 7 9 10 9 2 16 1 2 9 9 10 9 10 0 13 9 16 13 1 9 0 13 1 9 1 9 1 9 10 9 2 16 13 14 9 15 14 9 11 2 2
18 7 4 16 10 9 13 1 9 15 9 0 1 9 10 9 10 0 2
45 9 15 13 9 0 2 1 15 1 10 15 16 13 3 1 10 9 10 0 1 10 9 10 0 2 13 9 2 16 13 9 1 9 15 7 13 1 9 15 14 9 3 2 0 2
24 9 10 9 13 14 10 9 2 1 10 9 10 0 2 14 9 10 9 1 10 9 10 15 2
53 9 9 10 9 2 11 11 2 13 1 9 11 1 9 10 9 13 1 9 10 9 16 1 11 12 13 9 11 11 9 14 9 10 9 13 1 11 9 9 2 16 13 1 10 9 10 0 10 0 1 9 11 2
15 10 9 3 13 4 3 7 13 1 15 9 10 9 9 2
25 3 2 1 13 2 13 3 11 16 13 10 9 1 10 9 16 13 11 1 9 15 1 9 11 2
22 7 7 2 10 9 14 12 13 1 9 10 9 1 10 9 16 13 13 1 10 9 2
50 7 16 11 13 3 7 3 1 9 10 9 14 11 2 15 3 13 13 16 1 13 3 7 3 9 1 9 10 11 2 15 13 14 10 9 10 0 13 16 4 13 3 14 9 15 1 15 9 15 2
43 1 9 16 13 1 9 11 13 9 11 11 16 1 15 13 11 1 9 11 7 1 10 9 1 10 9 13 9 2 16 9 12 15 15 16 13 13 14 10 9 1 15 2
28 15 13 3 14 10 9 16 13 1 9 0 0 2 16 1 15 10 9 10 0 2 0 13 0 3 1 9 2
11 1 9 15 2 9 3 13 14 10 9 2
20 13 15 2 16 16 13 10 9 13 10 9 10 0 7 13 10 9 10 0 2
88 9 15 14 9 10 9 1 9 10 9 1 9 9 10 9 2 11 13 16 10 9 13 13 3 1 10 9 13 3 1 9 9 11 14 10 9 16 13 1 15 2 2 10 9 16 13 10 9 1 9 9 10 9 7 10 9 1 11 1 9 15 10 0 4 16 15 9 0 1 15 16 10 9 13 3 3 14 9 10 9 14 15 1 10 9 10 0 2
36 4 16 10 9 13 13 16 10 9 10 0 14 11 1 10 9 10 0 1 10 9 7 1 9 15 1 15 13 7 9 16 4 13 14 15 2
28 9 0 0 0 16 13 13 1 9 9 15 13 1 15 3 2 16 1 10 9 13 16 9 13 13 1 11 2
3 3 3 2
5 9 2 15 13 2
22 9 11 10 0 13 16 9 1 10 15 14 10 9 13 1 9 0 14 9 10 9 2
57 7 16 10 10 9 2 12 9 2 13 9 0 3 1 11 7 1 10 9 2 12 9 2 2 9 15 10 0 12 9 2 0 1 10 10 9 13 16 1 11 13 14 9 15 1 11 13 1 9 2 1 13 9 1 10 9 2
8 11 11 2 9 2 11 2 2
24 11 11 13 9 1 3 9 9 2 12 9 2 7 13 14 11 11 11 1 9 1 11 12 2
39 1 10 9 1 10 9 14 11 2 16 13 1 3 1 9 12 9 1 9 2 13 3 11 11 1 12 9 7 11 11 12 2 3 1 15 9 9 2 2
8 11 11 13 12 9 1 11 2
13 11 11 13 9 0 1 11 1 11 2 12 12 2
23 11 13 3 12 9 2 7 9 10 9 13 10 9 10 0 11 11 11 2 12 9 2 2
28 11 13 9 0 1 11 1 10 11 2 12 12 2 14 11 11 13 3 10 0 1 9 10 11 1 12 9 2
31 11 13 1 11 12 12 7 11 13 1 10 9 1 11 1 9 0 1 10 11 1 11 11 12 12 2 11 12 9 2 2
20 11 11 13 1 9 15 14 11 11 12 12 2 11 11 13 12 1 11 2 2
7 11 11 13 12 1 11 2
18 12 9 0 13 3 7 3 1 10 9 10 0 14 9 11 1 9 2
32 10 9 11 9 9 13 3 1 11 1 11 11 2 1 9 9 1 9 10 9 2 12 12 1 11 1 10 9 10 0 2 2
31 10 9 9 9 2 16 13 1 10 9 10 0 1 11 11 10 0 12 12 2 13 3 14 10 9 2 3 3 1 11 2
25 9 10 9 2 10 9 9 11 2 13 14 12 9 15 1 11 11 1 11 2 1 9 10 9 2
11 3 13 10 9 10 0 7 3 10 9 2
23 9 10 9 9 11 13 1 9 2 1 9 11 2 1 11 11 1 9 10 9 10 0 2
11 1 10 9 10 0 13 10 9 12 12 2
5 11 2 11 2 2
48 9 10 9 14 10 9 10 0 13 3 1 10 9 1 10 9 2 1 10 13 11 1 9 15 10 0 11 2 16 13 12 7 13 13 1 10 9 1 9 9 15 10 0 2 0 11 11 2
24 15 13 1 9 15 1 11 9 3 1 12 9 2 1 13 14 11 11 16 13 3 9 15 2
36 11 2 2 10 9 10 0 2 1 9 9 11 2 13 1 9 10 9 1 9 9 16 13 3 1 13 10 9 2 11 11 2 3 1 9 2
12 11 13 3 12 9 3 1 2 12 9 15 2
30 1 9 10 9 14 15 13 14 15 11 1 12 9 9 2 1 9 1 10 9 10 0 7 1 9 11 1 13 9 2
26 10 9 14 11 2 1 11 11 2 13 0 7 0 3 1 7 9 15 10 0 14 9 11 10 0 2
14 9 13 1 15 9 9 12 9 2 3 2 1 9 2
21 9 15 10 0 9 13 1 9 1 10 9 10 0 1 11 11 2 16 13 12 2
20 11 2 16 13 1 2 12 9 1 9 1 10 9 10 12 2 13 14 11 2
28 11 11 10 0 2 16 13 3 14 11 11 2 13 1 9 11 14 11 9 1 9 10 9 14 15 1 11 2
25 10 9 10 9 3 2 11 11 2 11 11 11 11 2 11 11 2 11 9 11 2 9 11 11 2
53 13 9 10 9 1 10 9 11 11 1 10 13 11 11 2 12 9 16 13 3 9 1 9 11 2 11 11 13 1 9 15 12 12 1 11 1 11 7 11 13 3 12 1 10 9 1 10 9 10 0 11 2 2
22 10 9 10 0 1 9 10 9 1 9 9 13 3 1 11 2 3 13 3 10 9 2
6 10 9 13 12 9 2
20 12 1 15 13 3 2 11 11 7 11 11 2 16 13 1 9 1 12 9 2
26 1 15 13 1 9 10 9 10 0 11 11 2 16 13 1 10 9 1 10 9 1 9 1 12 9 2
6 10 9 13 11 11 2
32 15 10 9 10 0 16 1 9 15 13 9 9 0 2 8 8 8 9 10 0 2 3 16 4 16 10 9 13 3 3 0 2
5 11 2 11 2 2
30 13 9 10 9 10 0 11 11 4 13 3 1 9 12 9 2 7 3 13 13 1 9 9 1 9 1 9 1 9 2
37 10 9 10 0 7 9 9 10 9 10 0 13 3 16 15 13 3 2 12 12 9 1 9 2 7 13 3 3 2 12 9 1 9 1 9 9 2
21 11 13 3 1 9 11 2 10 9 10 0 1 2 12 9 7 9 9 9 0 2
12 12 10 9 10 13 13 1 9 9 1 9 2
24 9 10 9 1 10 9 10 0 13 9 10 9 10 3 2 0 14 11 9 9 2 11 11 2
5 9 12 7 9 2
18 13 9 9 1 11 9 9 7 13 1 15 1 10 9 9 7 9 2
23 13 12 10 13 1 9 11 16 13 1 9 11 1 2 12 2 1 9 10 9 11 11 2
27 15 13 9 0 1 11 11 1 10 9 9 11 2 1 10 9 10 0 16 13 1 9 11 1 2 12 2
26 11 13 3 2 13 3 1 10 9 2 13 1 15 9 9 13 7 12 9 16 13 13 2 7 13 2
11 15 13 13 1 15 1 9 15 1 11 2
44 1 16 11 11 0 1 10 9 2 15 13 1 9 14 9 12 2 1 10 9 10 0 12 2 2 1 10 9 7 3 1 16 1 9 9 12 13 9 0 13 14 10 9 2
19 13 14 10 9 9 9 7 1 9 15 13 1 15 9 0 3 1 11 2
30 4 9 1 10 9 10 15 1 11 2 9 10 9 1 11 12 2 2 7 7 15 13 14 10 9 10 9 14 11 2
23 10 9 11 7 11 11 13 3 7 3 1 9 0 2 10 9 10 0 1 11 12 2 2
21 15 13 1 11 1 16 13 1 15 9 16 4 13 7 10 9 3 13 1 11 2
24 15 13 16 11 9 9 4 13 1 9 10 9 1 9 11 2 10 0 16 13 0 3 2 2
20 11 0 3 2 4 13 1 10 9 7 7 1 11 9 10 9 3 3 13 2
12 9 11 13 1 10 9 14 10 9 9 9 2
10 15 0 3 7 13 1 9 10 9 2
13 3 9 9 13 12 1 12 10 0 1 10 9 2
11 12 10 9 14 15 13 9 15 10 0 2
5 11 2 11 2 2
31 9 9 11 4 13 14 10 9 10 0 1 9 9 7 9 11 2 7 10 9 1 9 1 9 9 13 3 9 10 9 2
46 2 15 0 3 1 10 9 2 13 10 9 2 11 11 2 1 13 1 10 9 10 9 10 0 1 12 10 9 10 0 2 1 16 13 9 0 2 4 13 3 1 2 12 1 11 2
30 1 10 11 10 0 13 9 11 1 9 12 1 10 9 7 13 3 12 0 2 1 9 13 9 9 9 1 10 9 2
15 10 9 3 1 10 15 13 1 11 9 9 1 9 11 2
42 9 10 9 13 1 9 10 9 9 9 13 1 9 0 2 1 9 15 14 11 11 2 1 10 9 1 10 9 9 11 2 11 1 9 11 9 9 2 16 13 3 2
47 9 10 9 11 11 13 3 1 9 9 9 9 9 11 11 16 7 10 9 13 14 9 15 13 9 0 7 13 9 9 2 15 13 1 9 0 1 9 10 9 10 0 14 9 10 9 2
40 11 13 16 9 10 9 9 9 13 1 9 0 7 13 9 9 1 10 9 14 10 9 10 9 13 9 9 7 13 9 0 1 10 9 1 9 11 2 11 2
33 9 9 10 9 7 9 10 9 9 9 2 13 16 10 9 16 13 1 15 9 0 2 7 1 9 10 9 2 13 1 9 0 2
35 9 11 11 1 11 13 13 1 9 0 2 3 1 10 9 9 10 9 2 1 9 0 16 13 1 9 14 12 9 3 2 12 12 2 2
47 9 11 1 11 3 13 3 1 9 15 2 7 1 9 15 13 1 15 9 9 2 3 16 3 9 3 1 0 13 1 15 13 1 10 9 16 13 1 1 10 9 14 10 9 10 0 2
38 9 7 2 12 9 1 10 9 13 9 11 1 11 1 9 14 12 12 3 2 7 3 9 0 14 11 11 7 11 11 13 14 10 9 1 10 9 2
20 11 1 11 13 13 9 2 7 1 9 0 13 1 9 11 13 1 10 9 2
26 1 11 13 3 10 9 11 11 2 7 7 10 9 10 12 11 13 1 10 9 7 3 13 7 9 2
18 11 13 3 1 10 9 10 0 2 12 1 12 9 14 11 1 11 2
22 11 11 2 16 13 1 10 9 1 2 12 9 2 13 13 7 7 3 13 10 9 2
5 11 11 13 3 2
15 10 0 2 3 11 11 2 13 0 1 9 15 10 0 2
21 1 9 2 3 9 11 13 1 9 9 2 16 1 9 15 13 11 7 11 11 2
8 3 13 3 16 13 9 0 2
30 9 9 10 9 14 10 9 11 1 10 9 13 10 9 1 10 9 9 15 1 9 10 9 2 14 9 9 15 0 2
20 9 2 16 13 1 15 1 9 0 1 9 15 2 13 9 9 1 11 11 2
27 9 9 10 9 11 11 11 2 16 13 1 10 9 2 13 9 7 9 1 11 11 7 13 14 9 15 2
14 9 9 13 1 9 11 1 16 11 13 1 9 0 2
13 15 3 13 3 1 9 15 7 13 1 9 13 2
21 10 9 13 1 10 9 14 11 11 7 11 11 2 16 3 13 1 9 10 9 2
14 1 15 9 0 13 1 11 9 3 0 14 9 0 2
15 10 9 13 1 9 0 1 10 9 16 13 1 11 3 2
42 3 2 10 9 10 0 13 1 10 9 10 0 10 15 13 9 9 1 14 15 2 16 13 14 10 9 10 0 3 7 13 1 15 9 1 9 7 9 9 7 9 2
27 1 10 9 16 0 1 9 15 3 10 9 10 0 2 13 1 15 14 10 9 13 1 10 9 10 0 2
23 7 13 1 15 14 9 9 10 9 7 10 9 10 0 16 0 1 11 13 9 0 0 2
21 10 9 10 0 10 15 2 13 1 9 3 0 1 9 10 9 10 0 2 0 2
27 9 14 9 2 16 11 3 13 3 13 14 15 3 1 15 13 9 13 7 15 13 3 1 9 10 9 2
2 3 2
9 3 1 15 2 15 13 3 9 2
25 13 9 16 11 13 1 9 3 0 2 14 3 1 15 1 9 15 7 3 1 15 1 9 15 2
6 7 13 3 9 0 2
24 10 9 10 15 13 13 10 16 3 9 0 1 9 0 1 11 11 7 1 10 9 1 11 2
57 7 15 13 1 9 2 16 7 15 13 1 11 7 1 10 9 1 11 2 7 7 13 1 15 9 0 3 2 16 16 1 10 9 15 13 13 9 0 2 16 13 3 13 14 10 9 1 11 7 3 13 14 10 9 1 11 2
59 15 10 9 10 0 16 11 13 1 15 2 7 15 3 13 14 10 9 10 0 7 14 13 9 1 10 9 1 11 7 10 9 10 0 4 1 9 0 13 1 9 0 2 15 4 13 14 10 9 10 0 7 13 9 14 9 14 11 2
53 10 9 10 15 13 2 16 7 3 13 1 9 16 9 9 10 9 10 0 2 9 10 9 2 13 1 10 9 2 15 13 1 15 16 3 0 0 0 2 13 13 1 10 9 10 0 1 9 10 9 1 11 2
9 15 10 9 10 0 14 10 9 2
12 15 9 15 14 10 9 16 11 13 1 15 2
50 7 13 3 1 9 2 9 15 14 10 9 13 0 2 7 4 16 9 10 9 10 0 2 16 13 14 10 9 2 13 13 14 10 9 1 9 9 9 16 13 1 10 9 10 0 3 1 10 9 2
20 4 13 1 15 16 1 11 13 9 1 10 9 10 0 16 13 1 9 15 2
21 1 12 9 1 10 9 13 10 9 16 11 13 13 10 10 9 2 7 3 13 2
20 1 10 9 13 10 9 0 2 12 12 2 2 3 1 10 9 2 12 12 2
32 9 0 1 11 1 3 2 9 9 2 2 1 9 10 9 11 9 2 7 9 1 9 0 7 3 3 0 1 9 10 9 2
22 11 13 3 12 9 2 11 12 9 7 11 12 9 2 9 12 7 2 12 9 2 2
20 9 0 1 10 15 1 12 9 2 16 4 13 14 11 2 4 13 13 0 2
27 7 3 13 1 10 9 11 11 1 10 9 10 2 12 2 7 13 13 9 1 10 9 2 12 9 2 2
27 15 3 3 13 1 10 9 1 1 10 9 2 14 15 13 14 10 9 2 13 7 13 16 16 15 13 2
20 11 11 2 12 9 2 7 11 11 2 12 9 2 13 3 3 1 10 9 2
26 11 13 14 11 11 10 0 2 13 12 9 2 13 12 9 7 14 12 10 9 13 1 11 1 9 2
25 11 13 1 9 0 2 12 1 10 9 2 7 13 10 9 16 13 1 11 14 10 9 10 0 2
20 3 11 7 11 2 16 13 12 9 1 10 9 7 13 14 11 2 13 9 2
20 11 11 3 13 12 9 0 2 7 3 13 0 7 13 10 9 1 9 0 2
46 11 13 1 9 0 7 7 13 13 1 9 1 10 9 10 2 12 2 1 11 11 2 16 1 10 9 10 0 13 1 10 9 10 2 12 14 11 7 13 14 10 9 1 9 0 2
37 3 13 10 9 1 0 0 2 0 1 11 2 7 10 3 2 9 11 2 16 13 14 11 2 3 1 11 13 1 11 14 10 9 1 10 9 2
37 1 10 9 10 2 12 3 13 12 12 1 11 1 11 13 10 9 14 11 2 7 11 13 1 9 0 12 12 7 11 13 1 9 1 14 15 2
5 11 2 11 2 2
34 10 9 10 12 14 9 11 13 3 2 1 9 1 9 11 2 1 15 13 9 11 14 11 11 12 12 1 9 9 1 2 12 9 2
24 9 13 12 12 1 9 10 9 7 13 1 10 15 1 10 9 16 13 12 12 1 9 15 2
42 1 9 0 16 13 3 1 10 9 13 11 1 9 15 1 11 11 12 12 7 13 1 10 9 10 0 1 9 10 9 2 1 12 12 1 10 9 10 0 1 11 2
25 11 1 11 13 12 12 14 11 11 11 1 9 1 13 9 2 7 10 9 13 1 9 12 12 2
26 1 9 11 13 11 1 11 14 9 11 12 12 2 7 10 9 13 1 15 1 11 12 12 7 13 2
39 11 0 0 13 10 9 9 9 1 10 9 16 3 13 1 9 0 7 7 10 9 10 0 7 10 9 10 0 2 1 10 9 2 15 13 13 1 0 2
20 10 9 2 1 9 0 1 10 9 10 0 2 3 13 9 15 1 9 9 2
46 9 15 10 0 2 11 7 11 2 13 1 9 1 1 10 9 2 14 11 13 1 9 11 2 9 2 7 15 13 13 9 3 1 11 7 1 11 10 0 16 13 15 1 9 0 2
23 9 10 9 13 3 1 9 0 14 11 7 11 2 16 13 7 13 9 9 15 1 9 2
14 11 9 9 13 9 1 16 13 1 10 9 10 9 2
28 9 10 9 11 7 11 13 14 16 13 1 15 7 13 14 9 10 9 16 13 1 15 2 3 12 9 2 2
27 10 9 13 3 1 11 2 16 3 13 13 1 0 10 9 2 7 1 13 10 9 11 16 13 9 0 2
11 10 9 13 1 9 15 1 9 10 9 2
54 9 13 9 7 1 10 9 10 2 12 13 9 10 9 1 9 12 2 12 9 1 10 9 13 1 10 9 9 12 12 2 7 14 13 9 1 10 9 13 9 0 1 11 1 9 9 7 15 13 1 12 9 9 2
20 9 10 9 1 9 9 9 1 10 9 3 13 9 7 10 9 13 1 9 2
16 1 10 9 13 1 10 9 9 12 3 2 10 9 9 9 2
14 12 9 14 15 1 12 14 9 9 13 14 10 9 2
17 9 10 9 13 3 1 9 1 11 1 10 9 1 9 10 9 2
41 9 10 9 13 3 1 9 0 3 14 12 9 1 9 2 7 7 16 1 9 0 14 10 9 13 10 9 2 7 1 9 15 14 9 13 7 13 1 9 0 2
37 3 9 10 9 7 10 9 13 3 1 11 2 1 9 0 2 1 10 9 1 9 10 9 7 10 9 10 0 1 9 9 10 9 1 11 11 2
23 9 10 9 7 10 9 13 1 10 9 10 0 1 11 11 1 9 9 10 9 1 11 2
30 9 15 13 0 2 7 13 1 10 9 16 13 7 1 10 9 16 13 1 10 9 1 11 11 9 10 9 10 9 2
12 9 10 9 13 1 1 9 1 9 1 11 2
21 9 15 13 1 10 9 10 9 2 7 16 1 9 10 9 13 9 0 14 9 2
23 9 10 9 13 3 1 11 11 2 7 3 13 9 10 9 7 13 1 9 9 10 9 2
43 10 9 10 0 13 1 1 12 9 1 9 2 1 9 16 0 1 12 9 1 9 2 7 16 1 9 1 10 9 13 1 9 9 10 9 9 14 1 12 9 1 9 2
30 10 9 1 9 10 9 1 9 9 10 9 13 1 9 15 1 9 16 13 2 1 15 11 13 14 9 15 1 11 2
39 10 9 1 9 10 9 13 3 1 9 9 1 2 9 10 9 2 7 1 9 0 1 9 10 9 10 0 2 3 1 10 9 1 10 9 11 7 11 2
25 10 9 1 9 10 9 1 10 9 10 0 13 1 10 9 1 10 9 10 0 10 0 14 11 2
15 9 10 9 13 13 3 1 10 9 10 0 14 9 11 2
39 9 10 9 13 1 9 11 1 9 1 9 9 0 10 13 1 11 2 7 7 3 13 10 9 13 1 16 1 10 9 3 13 1 9 0 16 13 13 2
15 9 10 9 13 1 12 9 1 9 1 10 9 10 0 2
7 9 10 9 13 13 3 2
65 9 10 9 13 1 9 0 1 3 9 7 7 10 9 10 0 1 10 9 14 9 15 2 7 3 13 10 9 13 9 7 9 10 9 10 0 2 7 1 9 9 1 9 9 10 9 2 13 3 9 10 9 1 3 1 12 9 1 9 1 10 9 10 0 2
21 1 9 9 10 9 13 3 9 2 1 9 0 1 10 9 10 0 14 9 11 2
6 2 9 13 1 11 2
41 9 15 14 11 11 13 1 10 9 10 0 14 10 9 10 2 12 14 9 10 9 1 10 9 12 12 2 1 9 13 9 2 16 13 1 9 0 1 10 9 2
38 1 10 9 1 11 9 9 1 9 11 2 13 1 9 10 9 16 15 1 10 9 10 0 2 7 1 11 16 13 1 10 9 2 9 1 14 15 2
17 14 10 9 13 11 11 7 2 11 11 1 9 10 9 11 11 2
5 15 4 1 9 2
22 11 9 9 13 14 9 15 10 0 2 1 13 9 3 13 1 10 9 11 12 12 2
17 9 11 13 3 12 9 7 3 1 9 15 13 9 1 9 11 2
37 11 11 1 11 13 13 1 1 10 9 1 10 9 9 10 9 2 7 10 9 13 1 10 9 12 12 7 11 13 3 1 10 9 10 2 12 2
32 10 9 9 9 13 1 15 14 10 9 10 0 1 11 1 9 9 1 9 10 9 1 11 9 9 12 12 2 1 9 2 2
12 10 9 9 3 3 13 1 9 10 9 3 2
21 11 11 13 9 9 1 11 11 12 12 2 16 13 14 9 15 1 9 10 9 2
9 11 13 1 9 10 9 10 0 2
28 2 12 9 1 9 9 10 9 14 9 10 9 1 10 9 16 13 1 9 10 9 14 15 1 11 1 11 2
19 3 13 1 10 9 9 14 12 9 9 1 9 2 12 9 2 1 9 2
36 11 9 10 11 13 3 15 1 2 12 9 7 13 1 15 9 9 1 2 12 9 1 9 1 9 2 1 9 9 1 10 9 1 11 11 2
16 11 11 2 9 10 9 10 0 2 13 1 12 9 1 9 2
54 9 11 2 16 13 1 9 15 3 1 3 1 11 9 15 2 7 16 13 3 16 13 14 15 1 0 10 9 14 9 15 2 3 13 14 2 9 2 2 7 3 2 11 2 2 1 10 9 10 0 3 14 15 2
62 15 7 3 2 1 9 16 15 13 1 9 15 10 0 2 9 1 10 9 2 4 13 2 3 1 9 2 16 1 9 10 9 13 9 15 1 9 15 2 16 13 13 1 9 15 1 9 9 10 9 10 12 14 13 1 11 7 13 1 10 9 2
36 2 11 2 13 9 0 1 9 0 2 11 11 11 2 9 7 9 2 16 13 13 14 9 9 11 2 9 16 9 9 0 3 13 1 15 2
25 1 9 15 15 4 13 9 0 2 16 13 1 15 10 10 9 16 13 15 1 3 9 0 0 2
7 7 16 15 13 7 9 2
19 2 9 2 13 9 16 13 3 2 1 3 9 0 1 10 9 10 15 2
97 4 16 13 15 0 1 9 15 14 11 11 2 0 1 9 15 2 2 16 13 3 9 0 2 13 1 9 15 1 9 15 14 9 11 1 11 2 13 14 10 9 10 0 2 10 9 11 11 9 2 12 2 2 7 3 3 15 9 3 2 16 1 11 2 16 3 1 15 13 11 0 2 9 15 14 10 9 2 11 2 13 9 2 16 9 10 9 10 15 13 9 10 9 1 10 9 2
14 10 9 10 15 13 1 10 9 3 1 9 10 9 2
76 3 13 3 7 3 7 1 9 9 10 9 7 10 9 2 16 13 1 9 16 1 15 13 10 9 10 0 1 12 9 10 9 2 16 13 14 12 10 9 16 1 15 13 11 14 10 9 10 0 16 15 13 1 9 15 2 9 1 9 9 10 9 2 9 10 9 2 9 15 7 9 10 9 1 15 2
44 10 9 10 0 14 10 9 13 1 9 1 9 2 16 1 15 13 11 3 3 14 9 15 2 10 0 7 10 0 2 7 3 14 10 10 9 16 15 13 13 1 9 15 2
44 10 9 13 1 11 11 16 0 2 1 11 16 13 1 11 14 15 2 1 9 9 0 16 1 13 14 15 1 0 1 15 13 15 1 10 9 2 16 1 10 9 13 9 2
62 14 10 9 1 9 15 14 9 2 0 2 0 2 13 1 15 10 9 11 9 2 9 10 9 10 0 2 2 10 0 2 11 11 14 10 9 10 15 2 10 4 13 14 10 9 11 2 9 2 2 16 14 15 13 11 1 9 1 9 10 9 2
7 11 13 9 0 10 9 2
46 1 13 14 10 3 0 15 4 13 10 9 9 7 3 1 9 10 9 15 13 1 0 7 0 2 1 3 16 13 1 9 9 2 9 7 1 9 16 13 1 15 9 1 9 15 2
20 9 10 9 14 9 10 9 14 11 13 2 16 9 4 1 9 7 1 9 2
45 15 9 9 0 10 9 2 9 16 13 10 9 14 9 0 16 1 9 9 15 13 14 10 9 1 10 9 1 9 15 1 9 15 14 10 10 2 4 2 7 10 10 2 13 2
42 10 9 2 16 1 15 13 10 9 10 0 1 10 12 2 13 2 3 2 7 1 1 9 10 9 13 9 7 13 1 9 7 1 9 9 7 13 1 10 9 9 2
23 11 2 13 1 15 3 2 13 1 10 9 10 0 1 9 16 13 4 13 3 1 9 2
48 3 13 15 9 0 2 7 15 13 13 1 9 16 13 1 15 10 9 13 3 1 15 9 16 4 1 9 0 2 7 16 13 1 15 3 9 1 9 9 0 2 7 2 9 1 10 13 2
42 10 9 10 0 16 13 11 11 1 1 10 15 16 11 4 13 1 15 2 13 9 1 9 15 2 9 10 9 2 9 14 15 2 9 10 9 10 0 7 10 9 2
36 3 9 15 2 16 13 14 9 10 9 1 10 0 13 9 1 9 2 1 16 15 13 1 9 2 7 2 1 9 1 9 15 14 10 9 2
95 1 11 2 2 2 16 13 1 10 9 7 1 9 0 1 9 15 2 3 3 3 16 13 11 1 11 2 7 3 3 9 9 2 2 1 9 2 9 2 16 7 9 10 9 16 13 14 9 14 13 7 13 0 2 7 2 14 13 1 15 16 15 13 9 2 14 13 1 9 9 14 9 7 13 1 15 16 10 9 13 9 16 13 1 9 1 15 7 3 15 4 13 1 15 2
7 7 2 1 9 10 9 2
30 7 1 13 1 10 9 10 15 4 11 13 14 10 9 14 15 2 10 9 0 10 9 7 10 9 14 9 10 9 2
16 3 16 15 13 1 9 15 15 13 1 15 14 11 1 9 2
56 9 15 2 7 0 3 9 2 13 14 15 10 10 9 2 7 7 15 2 16 0 1 9 15 2 13 1 9 15 1 10 9 10 0 1 9 15 14 9 15 2 7 9 15 10 0 13 9 10 9 1 11 1 10 9 2
36 13 7 16 2 11 2 13 3 9 0 2 9 9 0 9 14 9 2 10 13 15 1 9 9 7 9 7 13 15 1 9 9 15 10 0 2
24 14 9 15 14 11 2 7 1 9 15 10 0 14 11 2 13 10 9 7 15 13 13 13 2
34 7 3 9 2 9 10 9 16 13 11 13 9 0 7 7 10 9 10 0 13 9 0 2 9 0 3 1 9 15 10 0 14 11 2
25 3 16 3 2 13 3 11 9 0 1 9 10 9 2 7 15 9 0 1 9 10 9 10 0 2
25 1 9 15 13 11 9 0 1 9 14 9 10 9 10 0 2 1 1 9 10 9 11 1 11 2
21 1 9 0 1 11 2 3 3 16 13 1 11 13 16 13 1 11 14 9 15 2
15 16 11 2 1 10 10 9 2 13 9 13 1 9 15 2
67 14 11 13 1 9 15 16 13 13 2 15 13 14 10 9 7 1 16 15 2 13 1 9 0 2 2 14 10 9 2 2 15 13 16 10 9 9 0 13 7 2 10 0 16 1 15 13 16 15 15 0 13 1 1 15 16 13 4 13 14 9 10 9 10 0 2 2
10 11 13 7 9 13 1 9 9 15 2
19 7 3 16 13 11 13 13 3 9 15 14 9 15 16 13 1 9 0 2
55 11 13 1 10 9 1 9 12 9 2 9 2 9 2 9 0 2 9 0 1 9 7 0 9 2 11 9 15 2 3 16 13 7 13 1 15 1 11 9 9 1 11 2 9 12 0 7 9 0 9 7 3 12 9 2
36 10 9 13 1 9 9 1 9 0 14 10 9 1 10 9 7 1 9 15 14 9 13 1 11 3 10 9 7 10 9 10 0 2 10 0 2
62 10 0 1 10 9 13 11 2 16 16 16 15 13 1 9 15 3 15 13 9 1 11 2 7 16 9 15 13 1 9 7 15 13 13 7 13 13 2 1 9 10 9 2 2 13 1 15 11 16 3 13 7 13 1 9 15 2 9 14 9 2 2
16 3 15 13 1 1 10 9 7 13 1 9 15 14 10 9 2
13 16 16 13 9 15 10 0 14 11 2 13 11 2
45 15 3 2 11 1 9 9 7 11 10 13 2 13 1 9 10 9 16 13 1 10 9 7 13 1 11 13 14 9 15 1 16 15 13 2 13 1 15 9 1 9 10 9 2 2
10 1 9 15 14 9 13 11 1 9 2
33 15 13 1 10 9 1 9 0 2 16 15 13 1 9 9 7 9 2 13 9 1 9 9 1 9 7 13 0 1 12 10 9 2
54 0 3 13 10 9 16 13 14 10 9 16 13 1 11 2 11 10 0 1 9 10 9 16 13 1 10 9 7 10 9 11 16 13 13 14 16 13 1 9 10 9 7 1 9 15 14 9 13 14 11 1 10 9 2
83 1 9 15 13 11 1 10 9 3 3 13 11 2 7 13 9 0 2 11 13 10 9 2 11 13 9 0 2 11 13 10 9 16 13 13 3 2 16 16 13 11 2 2 11 3 13 2 15 13 3 3 2 3 13 2 1 9 10 9 2 7 3 13 2 7 9 9 15 13 1 9 15 14 9 2 1 15 16 13 1 15 2 2
27 7 16 16 16 13 11 2 2 3 3 13 9 2 7 2 1 2 9 16 15 13 13 16 3 3 15 2
12 1 3 1 3 2 16 13 2 13 9 2 2
19 7 1 2 15 15 13 2 2 15 13 3 1 9 2 15 13 0 2 2
49 2 11 2 13 9 0 1 9 2 0 1 9 7 0 1 3 1 9 2 3 3 1 9 15 10 0 2 7 3 1 13 0 1 9 0 16 13 0 7 3 1 9 11 1 9 0 9 11 2
28 1 9 0 14 11 11 7 3 3 1 15 15 9 2 0 7 13 9 0 7 1 9 15 4 3 1 9 2
14 7 7 12 9 13 1 9 10 9 1 9 14 9 2
22 10 12 2 3 3 11 13 14 11 10 9 2 7 3 14 15 15 13 1 10 9 2
41 10 9 13 1 9 11 1 10 9 16 13 11 1 9 15 14 11 2 9 16 9 13 13 1 15 2 1 16 11 3 13 13 1 10 9 7 3 4 13 13 2
37 7 11 16 13 2 13 14 10 9 1 9 14 9 7 15 10 9 16 13 13 1 15 2 1 11 2 2 15 13 13 14 9 15 14 10 9 2
26 15 13 13 1 15 10 10 9 14 13 1 9 7 13 14 10 9 16 13 1 15 1 9 15 2 2
26 7 14 3 13 1 15 2 16 7 13 1 15 2 15 13 2 2 15 13 16 13 14 9 15 2 2
45 11 9 9 10 9 2 11 9 10 9 2 11 16 10 9 14 15 1 10 9 0 7 0 7 3 2 0 2 13 7 10 9 16 13 0 1 15 16 13 1 9 15 14 11 2
32 3 10 9 14 15 1 11 1 9 10 9 13 1 15 16 15 9 0 7 1 16 4 13 2 4 13 16 13 1 10 9 2
24 10 9 10 12 16 13 3 3 1 10 9 13 10 9 3 13 11 11 14 10 9 10 15 2
18 9 15 4 13 13 2 7 7 13 3 9 16 13 1 9 10 9 2
25 9 16 10 9 1 9 15 13 13 1 15 2 3 13 0 7 3 0 2 3 7 13 13 3 2
13 3 9 2 7 1 16 1 10 15 13 13 9 2
18 9 15 14 11 2 16 13 3 2 13 1 10 9 1 9 10 9 2
15 11 11 13 14 10 9 1 11 2 1 16 13 1 15 2
46 7 16 16 13 0 7 9 15 14 11 13 0 3 1 9 15 13 15 13 13 1 10 9 14 10 9 7 13 9 1 10 9 16 10 9 10 0 13 1 9 15 1 9 1 15 2
109 1 15 4 13 14 2 11 2 3 3 7 13 14 9 15 1 9 15 14 10 9 10 0 2 10 0 2 16 1 15 15 13 3 14 10 9 2 13 13 3 14 10 9 10 9 2 7 3 14 11 2 10 9 10 9 2 10 9 0 10 9 2 9 0 7 0 16 13 16 13 9 1 9 15 2 7 16 13 1 9 10 9 13 9 2 10 9 16 13 13 9 7 13 1 9 9 15 0 10 9 9 9 1 16 13 9 7 9 2
41 13 9 1 15 2 16 10 9 1 9 2 11 2 13 1 9 15 14 11 3 1 9 9 10 9 10 12 7 1 10 9 10 0 2 1 9 10 9 1 11 2
95 7 13 3 11 14 16 13 15 1 15 9 1 1 9 15 14 9 0 2 3 2 9 0 2 7 9 1 9 9 2 3 13 16 13 1 0 13 7 13 1 15 3 1 9 0 0 14 15 2 3 12 10 9 10 0 16 13 1 9 1 10 9 2 1 2 9 10 9 2 2 9 16 1 1 10 9 10 0 14 15 2 15 9 0 7 0 2 9 1 10 9 7 10 9 2
46 1 9 15 1 9 10 9 1 9 9 9 11 11 2 13 1 15 9 10 9 2 1 10 9 10 0 7 1 9 14 9 2 14 10 9 1 10 9 16 13 4 13 14 10 9 2
21 3 16 13 3 1 11 13 16 10 9 14 9 10 9 3 13 0 2 7 3 2
53 9 3 15 16 4 13 15 2 9 9 7 9 13 1 9 1 9 15 14 9 16 13 1 9 10 9 2 3 1 9 0 2 9 16 13 1 9 9 10 9 7 7 9 2 7 1 9 15 9 1 10 9 2
8 3 13 4 13 16 15 13 2
37 9 14 9 0 1 9 13 1 9 1 9 16 1 15 13 9 9 16 13 1 10 9 2 3 1 9 9 16 13 1 10 9 10 0 2 0 2
36 16 16 13 9 10 9 1 9 0 1 10 9 10 0 2 13 9 9 1 9 10 9 0 3 7 3 7 13 10 9 1 9 0 14 9 2
36 3 2 1 9 9 10 9 2 13 10 9 4 1 9 15 7 1 9 15 2 7 10 9 7 13 1 9 10 9 10 0 1 9 13 15 2
30 3 10 9 13 1 15 9 0 7 3 3 9 0 1 9 9 16 13 1 9 10 9 9 2 10 9 7 10 9 2
17 7 13 1 15 9 2 16 16 13 1 10 9 16 13 1 9 2
32 9 1 10 15 2 16 9 15 13 1 9 15 13 14 9 15 2 13 1 9 1 16 13 1 9 9 2 9 2 7 9 2
46 9 1 10 15 4 13 1 10 13 1 9 10 9 7 10 9 1 10 9 7 15 2 4 13 2 13 9 1 9 15 14 10 9 7 1 9 0 14 15 16 13 0 1 9 15 2
24 13 3 9 13 14 9 10 9 1 9 9 0 16 4 1 9 15 13 1 9 9 1 9 2
41 1 10 9 10 0 2 3 7 10 9 10 3 0 14 10 9 1 9 10 9 2 13 1 9 14 10 9 9 9 2 7 3 9 0 2 1 9 0 7 0 2
33 9 15 2 16 13 1 9 1 10 9 2 1 9 0 10 9 2 2 3 13 14 10 9 16 13 9 13 1 15 14 9 15 2
31 10 9 1 11 13 1 9 0 7 3 0 2 16 13 1 15 9 0 7 13 9 0 1 10 9 10 0 14 10 9 2
40 10 9 13 1 10 9 10 9 7 10 9 7 1 9 9 15 7 9 15 10 0 2 13 1 10 9 10 0 14 9 15 10 0 7 10 0 14 10 9 2
33 3 16 9 15 10 0 7 10 0 13 9 1 10 9 13 1 15 9 14 9 16 13 14 9 10 9 7 7 13 1 15 9 2
19 10 9 0 16 13 9 1 9 1 10 9 13 3 3 1 9 9 15 2
27 7 16 15 16 13 3 9 13 13 1 9 7 9 2 1 9 0 7 0 2 1 9 13 1 9 13 2
29 7 13 9 0 1 9 10 9 1 10 9 2 9 15 12 13 14 9 10 9 10 0 7 14 10 9 10 0 2
38 4 13 16 9 10 9 13 9 16 13 1 9 9 15 14 10 9 0 7 9 0 3 7 7 10 9 15 13 13 14 10 9 1 2 9 9 15 2
16 10 9 13 13 14 9 15 2 3 7 10 9 13 1 15 2
18 3 1 9 7 9 13 10 9 16 13 7 10 13 1 9 10 9 2
21 4 3 13 7 13 16 9 15 14 9 3 13 2 16 1 15 10 9 3 13 2
26 1 9 13 15 10 9 2 10 9 7 10 9 2 7 10 9 13 1 9 10 9 10 0 9 15 2
46 10 9 1 9 10 9 11 11 7 9 10 9 11 11 13 3 2 1 16 11 13 13 14 9 15 14 11 11 2 1 9 9 11 2 1 9 9 11 1 9 10 9 7 10 9 2
23 11 2 16 15 9 9 10 9 2 13 1 9 11 1 9 2 1 10 9 14 9 11 2
13 14 13 11 1 9 10 9 13 9 1 10 9 2
21 3 13 9 15 14 11 1 9 2 1 10 9 2 7 11 13 13 14 9 15 2
30 1 9 15 13 14 9 15 2 11 9 2 16 7 15 13 1 10 9 2 16 9 15 13 1 2 12 1 9 15 2
32 10 9 13 14 9 15 14 11 2 7 1 1 9 15 13 2 1 9 0 2 1 11 11 2 9 11 7 9 15 14 11 2
16 11 13 7 13 1 9 2 7 13 1 11 13 9 9 2 2
7 10 9 3 13 1 11 2
50 9 1 9 11 2 16 13 3 13 11 1 11 2 13 9 0 1 9 10 9 2 16 2 13 9 1 9 10 9 16 13 1 9 0 1 9 10 9 10 0 7 1 9 10 9 2 1 9 15 2
28 15 13 16 9 15 13 3 1 9 2 7 9 15 1 11 2 7 16 9 10 9 15 13 13 13 1 15 2
17 15 13 16 1 9 13 13 9 14 9 1 10 9 1 9 11 2
27 10 9 11 13 13 3 14 9 15 2 11 11 2 1 9 9 2 11 2 2 9 1 9 11 2 11 2
17 11 2 16 13 1 9 9 9 9 11 2 13 9 9 10 9 2
18 3 13 11 14 9 9 10 9 2 11 11 2 1 9 2 11 2 2
24 3 13 11 13 14 11 11 2 9 9 10 9 7 9 1 9 11 2 1 9 9 10 9 2
34 11 13 9 14 15 13 14 11 11 2 9 15 14 11 2 1 12 9 15 9 11 7 9 10 9 1 9 10 9 10 0 1 11 2
27 13 1 11 13 14 9 9 10 9 2 11 11 2 1 9 9 2 9 2 1 11 9 2 11 16 13 2
19 9 10 9 11 11 1 10 9 13 13 1 9 13 9 1 9 10 9 2
29 9 13 1 3 13 11 1 9 9 7 9 9 0 3 13 1 15 2 7 3 3 9 16 1 9 15 4 13 2
31 1 10 9 13 9 1 9 10 9 16 13 1 9 9 1 9 15 7 1 10 9 13 1 9 9 10 9 7 10 9 2
46 10 9 3 13 1 10 9 2 7 7 2 13 3 11 2 1 16 13 1 15 16 9 11 13 12 9 9 1 9 10 9 7 10 9 2 7 16 1 15 3 13 9 1 9 15 2
26 9 10 9 13 3 1 9 10 9 13 9 1 11 1 12 10 9 10 9 2 10 9 7 10 9 2
47 7 9 10 9 7 10 9 11 11 2 16 13 9 1 9 10 9 1 11 7 10 9 10 0 2 13 4 1 9 9 1 9 15 2 7 3 11 13 13 3 3 1 9 1 10 15 2
54 1 16 13 11 1 9 16 13 1 15 13 10 9 1 11 16 9 15 1 9 10 9 2 9 11 2 3 13 1 9 9 9 10 9 1 11 7 1 9 15 13 10 9 1 9 9 1 10 9 1 9 10 9 2
44 1 10 9 2 13 3 9 1 10 9 13 14 9 10 9 11 1 9 15 11 11 2 3 16 7 1 15 13 10 9 2 3 4 13 3 7 13 10 2 11 2 7 9 2
26 1 9 9 0 2 13 3 9 9 10 9 13 14 10 9 10 0 2 11 11 2 1 9 10 9 2
52 9 11 11 2 16 13 1 10 9 2 13 3 13 1 9 1 9 9 7 9 2 1 9 9 1 10 9 1 9 15 1 9 15 14 10 9 3 11 11 2 7 10 9 13 13 14 10 9 1 10 9 2
38 9 0 13 1 9 10 9 16 11 13 1 9 1 9 9 7 9 1 16 3 13 3 1 10 9 1 9 10 11 1 9 9 15 14 9 11 11 2
26 9 11 11 13 16 11 13 4 1 9 1 9 15 10 0 2 16 1 15 13 14 11 1 10 11 2
18 11 13 3 16 1 9 10 9 13 10 9 13 1 9 9 1 15 2
29 15 13 16 9 10 9 9 11 11 13 1 9 15 14 10 9 16 3 9 15 1 9 9 7 9 13 9 0 2
40 11 13 2 9 0 2 7 2 11 2 11 2 7 11 11 2 16 13 14 9 15 1 9 10 9 2 1 13 10 9 16 13 1 9 1 9 9 7 9 2
50 11 13 16 1 9 9 16 13 1 15 3 13 10 9 11 7 11 11 1 9 10 9 2 7 7 15 13 1 9 9 7 9 2 7 2 9 15 2 13 1 10 9 10 0 9 13 14 10 9 2
12 3 2 11 13 13 2 9 1 9 10 9 2
56 10 9 13 16 9 9 10 11 9 11 13 16 15 13 13 14 9 2 13 10 9 2 1 10 9 2 7 11 4 13 15 3 3 1 9 1 9 9 7 9 2 7 2 3 3 1 13 2 9 9 0 1 9 10 9 2
35 10 9 13 1 9 1 9 1 9 10 9 13 1 9 0 3 0 16 1 15 13 9 10 9 7 10 9 2 9 10 9 7 10 9 2
44 9 10 9 13 16 9 10 9 13 14 10 9 16 15 13 1 2 9 11 2 1 9 9 10 9 1 11 7 13 15 1 9 0 0 7 1 10 9 10 0 14 10 9 2
11 1 9 11 4 13 13 9 9 10 9 2
32 1 10 9 1 9 10 9 3 13 9 1 10 9 1 10 9 16 13 1 15 2 7 1 9 13 13 14 10 9 1 9 2
71 7 1 10 9 16 13 3 1 9 9 9 10 9 7 10 9 11 11 2 9 9 9 10 9 9 11 11 2 9 10 9 10 0 7 10 9 1 10 9 2 11 11 2 7 9 9 10 9 1 10 9 2 13 9 11 16 13 1 15 9 13 14 9 9 15 1 9 12 1 9 2
43 1 10 9 13 16 10 9 1 9 10 9 13 1 9 10 9 7 10 9 9 12 9 1 9 10 9 14 11 16 13 3 1 10 9 1 9 10 9 1 9 10 9 2
21 11 13 1 10 9 2 7 1 10 9 1 9 10 9 13 16 3 13 14 15 2
33 9 10 9 10 0 1 10 9 13 1 9 10 9 1 9 10 9 7 7 1 9 10 9 1 10 9 13 1 10 9 10 0 2
34 1 10 9 1 9 10 9 13 3 7 13 1 11 13 14 10 9 1 10 9 10 0 2 2 7 15 3 4 13 1 9 15 2 2
28 10 9 1 1 10 9 10 0 1 10 9 16 1 9 9 11 7 9 10 9 13 14 10 9 7 9 15 2
22 9 3 0 15 1 9 10 9 13 3 1 10 9 1 10 9 10 0 14 10 9 2
15 9 10 9 1 10 9 13 16 3 13 9 14 9 0 2
20 9 10 9 2 1 9 10 9 2 13 2 9 0 2 2 10 12 1 15 2
28 3 14 13 1 9 9 15 10 9 1 10 9 13 10 9 10 9 1 10 9 7 13 13 2 13 10 9 2
17 7 3 13 9 10 9 13 1 9 15 9 16 13 1 10 9 2
43 1 10 9 16 13 1 9 10 1 10 9 10 9 13 2 1 10 9 2 16 1 2 9 11 13 10 9 9 1 10 9 2 7 3 15 13 9 9 12 1 10 9 2
25 1 11 9 10 9 13 1 15 9 1 9 16 15 0 1 10 9 10 0 16 13 9 10 9 2
35 2 11 9 2 9 9 10 9 1 10 9 2 13 1 9 2 2 10 9 10 9 13 1 10 9 2 16 10 9 13 9 1 10 9 2
58 1 9 15 2 10 9 13 2 1 9 0 7 3 0 2 2 13 1 10 9 2 14 10 9 9 11 7 13 9 0 14 10 9 1 9 9 1 9 0 7 9 0 0 0 14 12 10 9 16 1 15 13 9 1 10 9 2 2
38 1 16 9 10 9 14 11 13 3 1 9 9 15 2 13 9 9 10 9 1 9 10 9 13 9 0 14 12 12 9 1 9 9 9 1 10 9 2
47 13 16 10 9 13 1 10 9 10 0 1 9 9 10 9 2 7 9 1 10 9 13 2 3 1 9 9 10 9 3 13 9 14 9 9 2 7 3 10 9 16 13 1 15 3 13 2
82 9 9 9 2 9 2 11 9 2 13 1 15 16 9 10 9 13 14 10 9 16 13 3 1 9 15 1 9 2 9 2 9 10 9 2 1 9 11 1 9 2 9 2 7 15 1 9 16 10 9 1 15 13 10 9 13 9 0 7 16 10 9 1 15 13 10 9 14 10 9 16 1 15 13 10 9 13 3 1 12 9 2
15 1 9 9 2 1 9 10 9 13 1 10 9 9 0 2
37 9 15 13 3 9 9 9 2 9 2 9 16 13 1 10 9 16 13 1 9 9 9 10 9 2 13 1 10 9 1 10 9 1 9 10 9 2
32 9 10 9 13 13 14 10 9 7 3 13 1 10 9 16 13 1 15 9 0 7 13 1 15 1 9 9 0 1 10 9 2
54 9 10 9 13 1 10 9 2 16 10 9 13 1 13 1 9 7 9 0 2 16 13 1 9 16 13 1 9 0 2 16 9 10 9 14 15 1 10 9 13 1 2 9 9 2 2 2 9 10 9 2 7 3 2
42 1 9 10 9 13 3 9 10 9 1 9 15 15 7 3 1 10 9 16 13 2 1 9 15 2 3 2 1 9 9 16 13 1 9 0 16 13 1 9 10 9 2
40 1 9 15 1 10 9 13 9 2 16 9 10 9 13 13 3 9 0 2 16 9 10 9 13 14 15 1 9 2 1 13 9 1 10 9 1 9 9 9 2
33 1 9 15 2 10 9 1 9 9 9 9 2 4 13 14 10 9 1 9 0 7 1 9 10 9 13 13 1 10 9 9 0 2
46 1 12 10 9 13 9 1 13 2 16 3 4 1 15 16 1 9 10 9 3 13 3 9 1 9 2 9 7 1 9 15 16 13 1 11 2 9 2 9 7 9 0 1 10 9 2
27 15 13 2 16 10 9 13 13 1 9 15 13 1 10 9 9 9 0 7 13 1 15 1 3 9 0 2
41 9 9 10 9 2 11 9 2 13 16 10 9 15 14 9 10 9 13 13 14 10 9 1 9 14 12 2 12 12 9 2 9 10 9 1 9 10 9 0 2 2
44 3 13 2 16 1 9 0 2 1 14 11 9 2 9 2 13 10 9 1 10 9 1 9 15 13 1 9 1 9 10 9 2 12 9 1 1 10 9 7 3 12 12 9 2
15 10 9 10 0 10 0 1 11 13 9 9 1 9 11 2
28 1 9 16 13 3 1 9 10 9 1 11 13 2 16 1 10 9 10 13 13 9 1 12 1 9 10 9 2
21 10 9 13 13 1 9 11 10 0 2 7 13 1 15 9 9 7 9 9 11 2
29 1 9 15 13 10 9 1 9 9 1 9 11 1 9 11 7 13 1 9 10 9 2 9 10 9 7 9 11 2
39 9 10 9 1 9 9 11 2 11 11 2 13 1 10 9 16 13 1 9 9 16 13 1 2 9 9 9 10 9 10 0 14 11 1 11 2 11 11 2
36 11 13 1 9 10 9 10 0 2 7 12 10 9 1 10 9 11 11 1 9 9 2 9 2 11 2 9 13 1 12 9 9 1 9 11 2
45 1 10 9 2 13 12 9 1 10 12 1 10 9 16 13 1 9 9 10 9 1 9 9 2 1 9 2 1 9 9 0 7 1 9 9 0 1 11 13 11 2 11 7 11 2
32 1 10 9 10 0 13 10 10 9 1 12 1 12 2 7 3 13 9 11 9 1 9 1 9 9 10 9 10 0 14 11 2
31 10 9 10 0 1 9 7 1 9 13 1 9 15 3 2 13 1 10 9 9 1 9 9 10 9 10 0 1 10 9 2
36 9 10 9 9 10 9 1 9 10 9 2 9 7 9 10 9 13 1 9 10 9 1 9 16 13 1 12 1 9 10 9 1 9 10 9 2
106 9 10 9 10 0 1 9 10 9 10 0 1 10 9 16 13 1 9 10 9 10 0 1 9 7 1 9 7 16 13 3 9 10 9 13 9 1 9 10 9 10 0 7 9 15 2 2 9 1 10 9 2 7 2 9 1 10 9 2 2 9 9 9 9 1 9 9 2 9 9 7 9 10 9 9 9 1 10 9 2 9 2 9 0 2 2 9 9 9 9 1 10 9 1 9 0 7 9 10 9 16 13 1 9 9 2
61 11 11 2 9 9 9 0 7 0 1 9 10 9 2 13 16 9 15 2 16 13 1 10 9 16 13 1 2 12 2 13 14 10 9 10 0 14 10 9 7 13 14 9 10 9 7 10 9 1 9 10 9 1 10 16 13 1 9 9 0 2
34 11 13 2 16 9 9 0 1 10 9 13 9 9 0 1 9 0 1 9 7 9 9 0 7 0 2 9 0 2 9 13 7 3 2
15 10 9 10 0 1 10 16 13 1 9 14 9 10 9 2
21 10 9 13 1 9 14 9 10 9 2 9 10 9 2 9 10 9 7 9 9 2
47 1 2 9 9 2 1 12 10 9 10 0 13 1 10 9 10 0 1 12 12 9 1 9 0 14 10 9 2 9 14 10 9 1 10 9 2 9 9 14 10 9 1 10 9 7 3 2
23 3 13 1 10 9 16 9 15 13 7 13 1 2 9 10 9 10 0 14 9 10 9 2
36 10 9 10 0 14 9 10 9 13 1 9 0 13 9 7 13 1 9 10 9 2 7 3 13 9 1 9 9 10 9 1 10 9 1 9 2
22 10 9 1 9 13 10 3 0 1 16 9 10 9 4 13 9 0 1 9 2 9 2
16 15 13 16 13 9 0 7 16 13 9 1 9 0 7 0 2
16 3 13 9 1 9 9 9 0 1 9 10 9 1 9 0 2
32 10 9 13 1 10 9 14 9 10 9 1 9 10 9 10 0 2 7 3 10 9 13 9 1 9 2 7 1 9 7 9 2
20 7 2 9 10 9 7 10 9 13 14 9 15 1 9 10 9 1 9 15 2
35 10 9 13 3 13 10 9 16 1 15 13 9 10 9 7 10 9 2 7 3 14 9 2 10 9 16 1 9 15 13 14 10 9 15 2
13 10 9 13 13 9 7 13 9 1 9 1 9 2
19 3 1 9 15 14 10 9 4 9 10 9 7 10 9 13 1 9 9 2
15 13 1 9 15 16 10 9 13 9 1 9 9 10 9 2
23 10 9 4 13 0 7 0 7 9 15 13 9 0 7 0 1 9 14 1 12 12 9 2
47 13 14 9 15 15 1 9 10 9 11 11 2 1 9 10 9 11 11 2 1 9 10 9 11 11 2 1 9 10 9 11 11 2 11 2 7 1 10 9 10 0 1 10 9 11 11 2
32 10 9 1 9 15 14 9 1 10 15 13 9 9 0 1 10 9 2 16 13 7 10 9 13 1 2 9 9 10 9 3 2
37 10 9 10 13 14 9 10 9 1 11 13 3 9 0 1 9 9 0 2 1 9 16 13 1 10 9 1 11 7 13 1 9 10 9 10 0 2
38 10 9 13 14 10 9 13 1 10 9 3 1 9 9 1 10 9 10 0 1 10 9 1 9 1 10 9 10 0 16 13 9 10 9 7 10 9 2
63 9 1 15 2 1 2 10 9 2 13 16 1 9 9 10 9 10 0 13 9 9 10 9 2 11 11 2 1 9 10 9 2 11 11 2 13 1 15 1 10 9 1 12 1 9 10 9 13 9 1 10 9 1 1 9 1 9 1 10 9 10 0 2
38 10 9 1 10 9 13 1 9 9 0 16 13 9 10 9 1 9 9 10 9 10 0 1 10 9 10 0 2 1 9 15 10 0 14 11 1 12 2
41 9 15 3 13 1 10 9 13 14 9 9 10 9 1 11 1 1 9 9 9 3 2 0 2 7 13 14 9 15 1 9 9 0 1 10 9 10 3 2 0 2
19 1 9 10 9 13 16 9 15 13 1 9 10 9 7 10 9 1 12 2
23 3 2 1 10 9 13 14 9 10 9 1 12 2 13 9 10 9 1 9 9 10 9 2
42 1 9 9 15 13 9 1 9 10 9 1 10 9 10 0 1 9 10 9 10 0 1 9 9 2 16 1 15 13 9 1 10 9 2 1 10 9 7 1 10 9 2
20 15 2 13 1 9 10 9 10 0 2 16 1 15 13 9 3 1 10 9 2
27 9 11 13 9 16 13 1 9 9 0 7 13 9 1 10 9 1 9 9 1 9 10 9 7 10 9 2
20 3 13 11 11 2 9 10 9 1 9 9 2 16 13 1 9 1 10 9 2
42 11 13 9 2 9 1 10 9 1 15 13 11 2 1 9 0 0 16 13 1 15 2 1 9 15 2 14 10 9 16 1 2 9 15 13 10 9 1 9 9 0 2
29 1 9 15 13 1 11 9 16 13 1 9 7 13 10 9 16 13 1 9 2 7 13 13 14 15 1 10 9 2
37 3 13 16 11 13 1 10 9 1 9 9 14 9 10 9 1 9 16 1 15 15 13 9 2 1 16 10 9 13 1 9 9 9 1 15 9 2
21 10 9 3 2 9 11 11 2 1 9 1 9 10 9 10 0 14 9 10 9 2
42 1 9 15 2 10 9 7 10 9 3 3 13 14 9 10 9 16 13 1 9 15 1 10 9 2 9 10 9 10 9 1 10 9 1 12 9 1 10 9 10 0 2
32 9 0 1 10 9 14 2 9 1 10 0 2 2 13 11 2 13 10 9 16 13 1 10 9 16 13 1 10 9 10 0 2
24 1 12 9 13 16 16 10 9 13 13 9 9 1 9 0 1 15 2 16 13 1 9 13 2
38 9 10 9 13 9 9 14 12 9 1 10 10 9 1 10 9 10 0 13 3 2 16 16 13 15 9 9 11 2 11 11 2 9 0 1 10 9 2
38 3 1 9 1 16 13 9 0 2 16 1 9 15 9 9 10 9 2 7 2 9 10 9 1 10 9 2 2 13 10 9 7 13 3 14 10 9 2
25 7 15 13 10 9 10 0 1 15 2 16 1 10 9 3 3 13 16 10 9 13 1 10 0 2
19 7 4 13 12 9 9 0 1 10 9 1 10 9 10 0 2 4 13 2
19 9 1 9 9 16 13 9 10 9 7 10 9 2 3 13 1 10 11 2
19 1 9 10 9 11 2 10 9 13 9 1 9 16 0 13 1 9 15 2
42 7 1 3 16 13 10 9 2 3 1 9 13 1 16 9 10 9 7 10 9 13 1 9 1 9 10 9 16 13 1 10 9 1 9 9 16 13 1 9 10 9 2
14 7 1 16 15 13 3 2 3 4 13 14 10 9 2
23 3 13 10 9 2 1 9 3 13 1 9 9 1 9 15 2 7 13 13 1 9 0 2
11 3 13 14 10 9 10 0 14 10 9 2
35 3 9 13 9 10 9 16 13 1 10 9 16 13 1 10 9 2 9 10 1 9 2 7 10 10 9 16 1 10 9 13 1 9 15 2
18 15 9 13 1 15 16 10 9 13 13 1 10 9 1 9 10 9 2
18 7 15 3 3 13 14 10 10 9 16 13 1 10 9 1 10 9 2
20 3 13 1 10 9 16 13 1 10 9 1 9 9 7 1 9 9 9 9 2
28 7 1 10 9 2 1 10 3 16 13 1 10 9 1 9 15 1 9 12 2 3 0 16 3 13 9 0 2
47 1 13 3 9 1 10 9 10 0 16 13 1 9 10 9 1 2 9 9 9 0 2 13 1 10 0 1 3 9 1 10 9 2 3 9 1 9 10 9 7 3 9 1 9 9 0 2
18 7 3 13 9 16 10 9 13 0 3 2 16 16 13 1 3 13 2
24 7 3 1 15 2 9 9 10 9 13 14 9 10 9 1 9 13 3 9 0 1 10 9 2
19 9 13 3 1 9 0 2 7 10 9 14 11 13 16 4 13 9 15 2
15 7 3 13 3 9 1 9 12 9 1 9 2 10 9 2
38 9 9 10 9 11 11 7 9 13 1 9 15 1 9 10 9 14 10 9 10 0 2 1 16 13 1 10 9 16 13 1 9 9 0 1 9 0 2
35 1 9 10 9 10 0 14 10 9 10 0 13 10 9 9 2 9 0 2 7 1 9 15 9 11 2 11 2 11 7 9 7 11 11 2
40 1 9 0 13 1 10 9 16 9 10 9 10 0 13 1 9 15 14 9 9 11 2 16 7 13 14 9 10 9 1 9 15 14 10 9 10 0 1 9 2
21 13 16 9 3 13 1 10 9 16 15 3 13 1 9 10 9 14 9 10 9 2
18 1 10 9 16 13 13 9 9 1 9 10 9 14 10 9 0 0 2
23 1 9 10 13 9 11 11 11 1 9 10 9 14 10 9 10 0 1 9 11 14 11 2
45 9 1 10 9 13 16 3 13 9 0 1 10 9 10 0 2 14 9 11 7 9 13 14 9 15 14 9 11 11 2 11 2 16 15 9 10 9 10 12 14 10 9 10 0 2
24 9 9 1 9 9 9 14 9 0 0 13 3 1 9 10 9 2 1 9 9 1 11 2 2
17 9 11 7 9 4 13 1 9 10 9 10 0 14 9 11 11 2
14 9 0 0 1 9 9 10 9 13 1 9 10 9 2
13 9 11 7 9 13 1 10 9 1 9 9 11 2
19 10 9 1 9 9 10 9 14 10 9 10 0 13 1 9 0 14 9 2
17 15 13 1 9 0 14 9 2 16 13 1 9 10 9 10 0 2
35 1 9 15 10 0 13 10 9 10 0 1 10 9 9 0 14 9 9 1 10 9 10 0 1 10 9 1 10 9 16 1 1 12 9 2
59 9 15 13 12 1 15 16 13 1 9 0 16 13 1 9 10 1 2 9 2 10 9 10 0 1 9 0 7 0 2 16 13 1 10 9 10 0 1 9 10 9 1 9 10 9 10 0 2 7 13 1 9 10 9 14 9 10 12 2
15 10 9 10 2 0 2 14 9 2 11 13 13 9 15 2
20 9 9 15 13 1 9 10 9 1 10 9 10 0 3 2 13 1 10 9 2
31 3 13 16 10 9 16 13 3 1 10 9 10 0 13 3 3 1 9 0 7 1 9 10 9 10 0 1 9 2 11 2
62 1 12 9 0 13 10 9 2 1 10 9 10 0 10 3 2 0 16 13 1 9 10 12 1 9 9 2 11 2 1 10 9 10 0 1 10 9 10 0 3 1 11 7 1 11 2 7 1 10 9 1 10 9 10 0 2 3 1 9 10 9 2
55 10 9 13 2 1 10 9 2 3 13 1 9 0 1 0 2 7 1 15 13 9 11 11 9 0 2 7 10 9 13 13 3 16 10 9 1 9 15 13 14 9 0 2 1 7 10 9 2 7 13 13 1 9 0 2
14 7 10 9 13 7 13 13 2 13 1 9 0 0 2
22 7 7 10 9 13 13 2 1 10 9 10 0 16 15 13 2 7 13 1 9 0 2
45 9 11 11 2 11 13 16 1 9 2 11 2 1 16 13 13 1 9 7 9 2 9 10 9 10 0 7 10 9 10 0 2 10 9 10 0 3 13 13 1 9 15 7 0 2
30 9 11 11 13 16 9 11 11 2 16 13 1 9 10 9 10 0 2 13 14 10 9 1 9 1 9 0 1 0 2
55 1 10 9 10 0 1 9 10 12 7 1 10 12 16 13 13 10 9 2 16 1 9 15 10 0 2 12 1 9 10 9 14 15 2 13 9 0 1 10 9 10 0 10 0 2 7 3 1 9 10 9 1 10 9 2
33 9 11 11 13 16 10 9 13 3 9 0 7 9 0 16 13 2 1 10 9 1 9 9 2 9 1 9 1 11 7 9 0 2
35 9 11 11 13 16 1 16 10 9 10 0 13 3 1 10 9 10 0 10 0 2 10 10 9 10 0 13 0 0 1 10 9 10 9 2
44 13 1 10 9 2 16 1 10 9 16 13 14 2 10 9 10 0 2 1 9 14 9 16 13 3 3 1 13 7 13 1 15 2 13 1 9 15 9 0 14 9 7 9 2
42 1 9 2 1 9 10 12 14 10 12 10 12 2 16 13 9 0 1 9 2 7 9 2 10 9 1 11 2 13 9 9 1 9 16 13 2 3 2 14 10 9 2
92 9 10 9 10 0 1 10 9 7 1 10 9 10 0 1 9 10 12 12 13 1 9 0 14 9 9 0 1 9 7 9 2 1 2 1 9 9 11 11 2 1 10 9 1 9 2 9 2 7 1 9 9 11 11 1 10 9 10 0 16 13 1 10 9 13 9 9 0 2 9 9 15 14 9 11 1 11 1 11 2 7 9 10 9 14 11 11 1 9 2 9 2
19 1 9 10 9 13 10 9 2 3 13 14 9 2 11 1 9 10 12 2
35 9 11 9 13 16 4 13 1 9 15 10 0 7 9 15 10 0 1 9 0 14 9 10 9 10 12 7 1 10 9 16 13 1 15 2
40 9 10 9 13 1 10 9 16 9 10 9 10 0 7 10 9 10 0 13 1 10 9 3 3 0 1 16 16 10 9 10 0 13 13 1 10 9 10 0 2
57 1 10 9 16 13 3 1 9 2 10 9 10 0 1 10 9 1 9 2 9 2 13 10 9 11 11 2 1 9 9 10 9 7 10 9 14 9 11 2 14 10 9 1 9 10 9 16 13 3 1 10 9 1 9 9 12 2
19 9 10 9 3 13 1 9 10 9 1 10 9 1 9 12 1 10 9 2
36 10 9 11 13 16 7 16 13 1 10 9 9 1 10 9 10 0 2 13 10 9 1 9 15 1 1 10 9 10 0 1 9 2 10 9 2
43 1 10 9 13 9 9 9 11 16 10 9 16 13 1 9 11 2 7 9 15 13 9 10 9 2 13 1 9 9 1 10 9 7 1 9 9 1 15 13 3 1 9 2
33 10 9 13 16 10 9 13 1 9 14 9 12 1 9 15 2 11 11 2 9 9 9 1 9 10 9 2 16 16 13 10 9 2
25 11 13 1 9 16 13 1 10 9 9 1 9 0 16 13 1 9 7 9 9 9 1 9 11 2
22 1 10 9 3 13 9 10 9 2 16 13 9 1 15 13 14 9 15 1 10 9 2
48 10 9 10 0 1 9 2 9 13 3 9 1 9 14 12 12 9 16 13 9 10 9 11 1 9 10 9 11 11 2 9 9 9 1 9 2 9 2 7 1 11 11 9 9 9 1 11 2
69 1 10 9 16 13 1 9 9 13 13 9 9 10 9 2 9 11 11 2 16 12 10 9 13 1 9 10 9 9 2 1 9 2 1 9 9 9 1 9 9 10 9 2 7 10 9 16 13 1 11 13 9 10 9 16 13 1 9 9 10 9 2 7 16 13 4 13 2 2
23 9 10 9 2 13 1 10 9 2 13 10 9 1 9 14 10 9 16 13 1 10 9 2
6 3 13 9 9 13 2
45 9 0 1 11 11 2 16 13 9 12 9 14 9 0 2 0 9 1 11 9 11 7 9 9 7 9 13 1 10 9 16 13 3 9 1 9 1 11 1 9 11 9 7 9 2
24 10 9 7 9 15 11 11 13 3 1 9 2 10 9 10 0 9 1 9 14 12 12 9 2
81 9 10 9 2 9 11 11 2 13 1 9 10 9 16 13 1 9 0 7 13 1 9 15 14 9 3 2 0 1 10 9 2 16 13 1 9 15 14 10 9 7 1 9 0 14 10 9 2 9 10 9 2 2 16 1 9 0 14 9 9 0 13 13 14 9 15 7 9 15 7 13 1 9 9 2 9 2 9 7 9 2
25 9 10 9 13 10 9 2 9 0 14 9 9 0 2 9 9 0 7 9 0 1 9 10 9 2
32 1 2 15 13 9 10 9 16 13 1 9 10 9 7 13 1 15 9 0 1 13 9 0 0 2 1 9 1 10 9 2 2
48 1 9 9 10 9 2 13 1 15 9 9 10 9 16 15 4 13 9 7 7 3 1 9 1 10 9 10 0 2 9 1 9 11 11 2 16 7 3 3 3 13 10 9 9 14 10 9 2
34 1 9 10 9 2 1 9 1 10 9 14 10 9 1 10 9 10 0 2 1 15 13 10 9 9 0 14 12 9 2 13 10 9 2
6 3 3 13 9 9 2
30 12 9 16 13 1 9 10 9 12 2 12 7 12 1 9 11 1 11 2 1 11 13 3 9 14 9 1 13 9 2
18 10 9 16 13 1 9 2 9 10 9 1 11 13 1 1 12 9 2
48 9 10 9 2 9 11 11 2 13 1 9 10 9 16 9 10 9 2 10 9 2 13 1 9 9 15 1 9 11 11 2 16 1 9 13 1 2 9 13 9 7 3 9 15 13 1 13 2
16 9 10 9 2 1 9 10 9 2 13 9 9 0 7 0 2
5 3 13 9 9 2
49 9 2 10 9 10 0 1 9 2 9 13 3 9 9 0 1 15 1 9 9 13 1 9 7 9 14 9 9 1 9 9 2 11 2 1 1 9 1 10 9 16 1 10 9 1 9 10 9 2
13 10 9 1 9 12 10 9 13 1 12 1 11 2
29 1 12 10 9 10 0 14 10 9 13 12 9 1 9 7 1 9 9 1 9 2 1 9 0 14 12 12 9 2
20 9 15 13 1 2 10 9 2 1 9 10 9 1 8 8 9 1 9 11 2
52 1 12 9 1 9 10 9 2 12 12 9 2 13 1 9 10 9 10 0 2 12 9 1 9 11 2 12 9 1 9 11 2 12 9 1 9 11 2 9 9 2 0 16 13 9 1 10 9 10 0 2 2
12 10 10 9 13 1 9 10 9 7 10 9 2
34 10 9 14 9 11 13 16 3 13 9 2 9 0 1 9 10 9 1 11 2 3 13 9 0 1 10 10 9 16 13 13 1 9 2
24 1 2 9 10 9 10 0 2 13 1 10 9 13 1 9 1 1 12 9 1 9 9 15 2
32 16 16 10 9 1 10 9 3 13 1 9 9 1 10 9 2 13 9 11 13 9 0 1 10 9 16 13 1 9 1 9 2
32 10 9 10 0 13 1 12 9 1 12 10 9 10 0 14 10 9 2 1 10 9 10 0 3 2 7 13 1 12 12 9 2
35 1 10 9 10 0 1 9 13 3 16 1 12 12 9 1 9 15 13 1 9 9 9 10 9 2 7 12 12 9 1 9 9 7 9 2
34 1 9 11 7 11 13 10 9 14 9 10 9 16 13 1 11 1 3 1 12 9 1 11 7 11 2 1 9 10 9 1 10 9 2
26 1 11 2 11 3 13 10 9 0 1 12 12 9 7 13 0 1 12 9 1 10 9 10 0 3 2
14 10 9 0 13 1 12 9 7 13 1 12 12 9 2
14 1 9 11 2 13 10 9 10 0 1 12 12 9 2
16 10 9 13 1 12 12 9 2 7 10 9 1 12 12 9 2
19 1 11 7 11 13 10 9 10 0 1 12 9 1 12 10 9 16 13 2
23 9 15 13 1 9 1 10 9 1 12 9 1 16 1 10 9 1 15 9 2 13 9 2
50 1 10 9 10 0 13 10 9 1 9 7 1 10 9 1 12 12 9 1 9 1 9 2 0 1 12 9 1 10 0 10 0 1 11 7 11 1 9 14 12 9 1 9 15 1 11 7 11 3 2
39 9 9 1 9 2 7 9 7 9 2 13 1 12 12 9 1 9 1 9 1 11 7 11 7 13 0 1 12 9 1 10 9 1 12 10 9 16 13 2
16 9 9 9 13 1 12 9 7 13 1 12 12 9 1 9 2
8 9 9 9 13 1 12 9 2
27 1 11 13 9 10 9 1 12 12 9 2 12 9 9 0 2 12 9 9 9 2 7 12 9 9 0 2
41 10 9 10 0 13 1 10 9 10 0 1 12 12 9 1 9 1 9 2 0 1 12 9 1 12 10 9 16 13 1 9 1 9 14 12 9 1 11 7 11 2
17 10 9 1 9 10 9 2 10 9 7 10 9 13 1 12 9 2
16 1 15 2 13 9 1 10 9 14 9 10 9 7 10 9 2
40 1 9 10 9 13 9 14 12 9 1 10 9 10 0 2 7 7 1 10 9 10 0 13 9 14 12 9 2 7 15 13 1 12 12 9 1 9 1 9 2
20 9 16 13 9 9 1 9 10 9 2 13 1 9 1 9 9 9 10 9 2
16 9 0 15 13 1 9 10 9 10 0 1 9 15 1 9 2
37 9 10 9 13 1 10 9 16 13 9 9 10 9 2 9 0 1 9 9 9 7 10 9 1 9 10 9 9 11 9 7 9 10 9 10 0 2
41 10 9 13 16 1 9 10 9 12 7 1 9 0 2 13 9 9 2 9 9 14 9 1 9 9 0 2 1 9 1 9 15 1 2 9 10 9 10 0 2 2
88 1 9 10 9 12 2 13 9 9 1 10 9 10 0 7 9 10 9 10 0 7 1 9 15 9 10 9 3 13 1 10 9 1 9 10 9 10 0 16 13 1 9 0 2 2 13 1 9 9 0 1 10 16 13 1 10 9 1 10 9 10 0 2 7 13 2 3 2 1 9 10 9 9 13 9 1 9 9 1 10 9 10 0 1 9 10 9 2
31 10 9 13 16 10 9 3 13 14 10 9 1 9 10 9 16 13 1 9 0 2 7 13 1 15 1 9 9 10 9 2
83 9 2 9 10 9 10 0 9 2 9 2 9 2 10 9 11 11 7 11 11 2 13 16 9 10 9 13 7 7 3 1 9 16 13 1 10 9 2 7 2 1 9 15 9 3 1 10 9 16 10 9 13 13 13 1 9 10 9 12 3 1 10 9 2 7 1 15 13 4 13 10 9 10 0 7 9 15 13 15 7 13 15 2
83 1 9 9 9 10 9 1 9 9 2 9 10 9 10 0 2 2 4 9 13 9 1 9 10 9 10 0 1 9 9 10 9 2 7 7 3 2 13 1 9 15 10 0 14 10 9 2 2 7 7 10 9 16 13 1 9 10 9 12 13 13 2 1 9 15 10 0 2 14 10 13 1 10 9 7 3 13 1 9 9 10 9 2
67 3 13 9 16 9 10 9 10 0 13 12 9 1 10 9 10 0 16 13 3 1 2 9 0 2 13 9 9 10 9 15 2 16 13 16 9 10 9 14 10 9 10 0 1 9 10 9 12 13 12 9 3 2 1 13 1 9 9 15 14 10 2 9 10 0 2 2
50 3 13 9 16 10 9 1 2 9 10 9 2 14 10 9 10 0 9 2 9 2 1 9 9 14 12 9 1 10 9 10 0 1 9 0 2 13 7 9 9 2 16 3 13 1 9 9 10 9 2
30 9 9 10 9 13 1 10 9 10 0 13 1 9 0 7 0 2 1 9 9 1 9 9 15 14 1 9 10 9 2
9 13 16 10 9 13 1 11 15 2
21 13 1 15 3 2 16 1 9 9 15 1 9 10 9 2 13 13 13 1 9 2
23 8 9 10 9 2 2 13 1 9 15 14 9 9 10 9 14 10 9 10 0 1 9 2
22 11 13 16 1 15 13 3 13 2 16 15 10 9 10 0 14 15 1 9 10 9 2
32 1 10 9 13 16 9 10 9 16 13 10 9 1 10 9 1 10 9 10 0 13 9 0 1 2 1 16 10 9 13 3 2
41 1 2 9 10 9 1 15 13 11 2 7 9 10 9 2 13 11 2 2 0 11 2 7 10 9 11 2 7 13 9 1 10 9 13 13 1 15 9 0 0 2
39 8 1 9 9 10 9 16 13 3 10 9 10 0 1 9 13 9 10 9 2 16 13 9 12 1 9 10 9 2 7 13 1 9 9 1 9 9 9 2
38 1 9 10 9 2 16 13 1 10 9 10 0 2 13 10 9 13 1 12 9 2 3 16 13 1 10 9 1 10 9 7 1 9 10 9 10 0 2
28 8 2 9 9 10 9 10 0 2 13 3 1 2 9 9 11 2 9 16 13 1 9 10 9 1 10 9 2
29 9 13 16 1 10 9 1 9 10 9 7 9 10 9 7 10 9 2 13 1 9 10 9 1 10 9 1 11 2
13 13 16 10 9 13 9 0 16 13 1 9 15 2
27 3 13 11 13 14 9 10 9 16 4 13 1 2 11 11 2 2 16 13 13 14 10 9 1 10 9 2
11 9 13 16 4 13 15 1 12 1 11 2
22 8 10 9 3 13 3 1 10 9 16 13 1 9 10 9 10 0 1 9 10 9 2
38 3 13 9 2 1 9 15 2 9 2 9 13 1 9 1 10 9 10 0 16 13 1 9 2 10 9 10 0 1 11 1 10 9 16 0 12 9 2
58 1 9 15 13 9 2 16 13 1 9 0 13 1 9 10 9 2 16 1 15 13 9 1 10 9 1 9 9 15 10 0 1 10 9 10 9 7 1 7 10 9 9 0 9 7 1 9 10 9 7 7 1 9 9 15 10 0 2
12 9 9 13 16 2 10 9 0 7 0 2 2
4 10 9 13 2
61 1 9 10 9 13 3 9 10 9 9 10 9 7 10 9 3 8 8 10 9 10 0 3 13 1 9 10 9 2 7 9 10 9 7 9 10 9 10 0 13 14 10 9 1 15 2 7 9 15 14 10 9 13 3 1 9 15 14 10 13 2
44 10 9 1 10 9 1 10 9 2 13 1 9 10 9 9 1 9 10 9 10 0 1 10 9 2 2 7 1 15 13 1 15 13 9 9 1 9 10 13 2 1 9 15 2
29 11 13 16 1 9 1 9 10 9 7 1 9 10 9 10 0 1 10 9 2 4 13 9 1 9 7 1 9 2
28 1 9 9 16 13 12 9 1 9 13 12 9 2 9 2 7 1 3 16 13 12 9 1 9 13 12 9 2
31 1 15 16 13 13 7 13 16 1 9 9 9 13 9 1 9 15 10 0 2 13 11 16 4 13 9 9 1 9 9 2
30 1 2 1 10 9 2 2 9 10 9 14 9 10 9 1 9 11 2 13 16 13 10 9 10 9 1 9 10 9 2
25 2 1 10 9 2 13 14 10 9 16 13 3 1 9 9 0 1 15 13 2 9 9 10 9 2
42 13 9 1 2 1 10 9 2 2 7 7 1 9 12 2 1 10 9 16 13 15 9 0 1 10 9 13 14 9 10 9 2 1 10 9 16 3 13 9 1 9 2
27 8 8 1 9 10 9 2 10 9 1 10 9 1 9 10 9 7 9 2 13 13 1 9 15 1 11 2
16 11 13 14 9 15 1 10 9 1 12 9 2 1 13 9 2
18 11 3 3 13 3 13 2 7 13 16 13 0 7 13 16 15 9 2
40 8 2 12 2 9 9 10 9 1 9 11 2 11 2 9 2 9 2 1 9 10 9 2 13 1 9 9 10 9 14 9 11 2 9 9 1 10 9 2 2
10 11 2 0 1 2 10 9 2 2 2
50 9 11 13 16 9 10 9 10 0 16 13 1 9 15 1 11 1 9 11 7 11 13 1 9 10 9 14 9 9 0 2 0 0 2 1 9 16 13 9 0 1 11 2 16 11 13 0 1 15 2
16 3 13 9 10 9 2 11 11 2 1 9 9 15 1 11 2
49 15 10 9 10 12 2 1 10 9 10 0 14 9 0 1 11 2 16 13 16 11 0 1 9 9 0 1 11 1 11 1 9 9 16 13 9 1 12 10 9 2 7 13 9 0 1 10 9 2
52 9 10 9 13 2 1 9 9 1 9 11 2 16 13 3 9 14 9 7 9 0 1 10 9 10 0 2 7 16 2 4 13 9 15 14 9 1 9 0 1 12 10 9 2 16 13 1 9 14 9 2 2
47 3 13 10 9 2 1 9 9 1 9 0 2 16 1 11 13 1 10 9 16 11 13 9 0 14 9 1 9 11 2 7 13 2 7 15 3 7 11 13 9 1 15 7 3 7 3 2
20 2 13 1 15 9 9 1 9 16 13 2 2 13 9 0 1 9 10 9 2
32 12 10 9 16 13 1 10 9 13 1 9 15 9 0 14 9 9 1 11 1 9 10 9 10 0 2 16 13 9 9 0 2
33 1 9 1 10 15 2 7 2 13 9 1 9 0 2 0 1 13 9 16 1 15 9 10 9 14 12 10 9 13 14 15 9 2
19 11 13 2 1 10 9 2 16 11 13 9 1 9 1 11 2 7 13 2
15 9 10 9 3 13 1 10 9 16 11 13 7 11 13 2
23 9 12 16 1 15 3 13 9 0 1 9 10 9 1 12 10 9 13 10 9 10 0 2
31 12 10 9 10 0 10 13 14 11 13 10 9 1 9 1 9 10 9 10 0 16 13 1 10 13 1 11 7 1 11 2
32 9 9 10 9 14 11 2 13 3 16 11 2 13 1 9 0 1 11 1 10 10 9 2 16 3 9 10 9 1 10 9 2
16 15 13 7 13 14 9 10 2 9 10 0 2 16 11 13 2
29 9 0 0 1 11 13 13 1 10 9 2 7 13 7 9 10 9 10 0 13 3 1 9 0 1 9 10 9 2
35 9 9 15 14 10 9 11 11 2 9 10 9 14 9 10 9 16 9 15 13 2 13 3 1 9 2 10 9 1 9 11 11 7 9 2
38 9 15 16 13 1 9 9 13 1 10 9 14 9 10 9 10 11 10 0 11 2 16 15 1 9 10 9 14 9 10 9 11 16 1 9 9 0 2
42 10 9 14 9 11 11 9 7 9 2 1 15 13 9 10 9 2 13 1 9 9 12 9 1 9 11 12 2 1 9 9 10 9 2 3 13 11 14 10 9 15 2
12 1 9 15 4 13 12 9 1 9 10 9 2
28 10 9 13 1 2 9 9 11 11 1 9 9 11 7 11 2 16 15 10 9 1 9 9 10 9 14 11 2
59 12 9 13 1 9 10 9 2 9 11 2 16 12 1 9 15 13 11 11 2 16 13 9 9 9 2 9 14 9 0 2 9 11 1 9 2 9 2 16 9 15 13 1 10 9 10 9 2 0 2 10 9 11 11 2 9 11 11 2
41 10 9 10 0 16 13 1 10 9 13 12 12 9 2 7 10 9 13 14 10 9 1 9 1 9 10 9 10 0 16 13 1 9 2 10 9 10 0 1 11 2
32 10 9 13 3 1 9 0 14 12 9 2 1 16 10 9 13 1 12 12 9 2 1 1 12 9 3 1 3 16 13 3 2
12 3 1 10 9 13 10 9 1 12 12 9 2
15 1 10 9 13 9 3 13 9 2 11 1 9 10 9 2
45 9 9 10 9 10 0 13 3 14 11 11 1 9 15 1 9 10 9 7 9 10 9 10 0 14 10 9 2 7 13 9 1 9 10 9 11 11 7 1 10 9 9 10 9 2
22 1 11 13 1 9 15 10 9 10 0 1 12 9 10 9 1 9 10 9 10 0 2
25 10 9 13 1 1 9 0 0 16 13 3 1 11 1 9 9 10 9 1 9 10 9 10 0 2
57 9 10 9 13 1 10 9 1 9 15 1 10 9 2 1 10 9 1 11 1 11 2 7 15 13 1 15 1 16 13 1 9 1 11 2 16 1 15 13 1 15 1 9 11 7 1 9 13 9 10 9 14 9 9 10 9 2
35 1 10 9 13 3 9 10 9 11 11 2 9 9 9 2 11 2 1 9 10 9 1 10 9 2 7 3 13 9 15 1 9 10 9 2
37 11 15 3 13 3 1 10 9 2 1 16 3 13 13 14 15 1 9 16 13 0 2 16 16 10 9 13 1 9 14 9 10 9 14 10 9 2
25 1 2 9 9 15 14 11 7 9 15 2 9 11 7 11 2 13 13 14 10 9 16 16 13 2
15 8 8 1 10 1 10 12 9 10 9 13 1 10 9 2
13 9 1 9 10 9 10 0 3 13 1 10 9 2
39 1 2 9 9 15 14 11 11 2 9 9 9 9 10 9 2 13 13 1 9 14 10 9 13 14 11 7 9 15 7 13 10 9 2 16 16 13 11 2
6 10 9 13 9 12 2
39 10 9 13 16 13 1 9 10 9 13 14 11 1 9 15 1 9 10 9 10 0 2 1 16 9 15 13 13 3 1 10 9 1 11 1 9 10 9 2
18 12 1 9 10 9 13 1 9 15 14 11 2 12 13 7 12 13 2
33 11 11 13 3 1 13 16 10 9 7 10 9 13 0 2 7 16 15 13 13 1 9 2 10 9 1 9 13 14 9 10 9 2
38 1 10 9 2 9 0 2 13 3 11 16 11 13 9 16 13 1 15 1 9 9 1 9 10 9 2 1 9 14 9 9 16 13 14 10 9 15 2
36 11 13 16 1 10 9 13 3 9 1 9 10 9 9 10 9 2 9 9 11 2 7 13 14 10 9 1 2 9 14 9 9 10 9 2 2
31 11 13 1 9 14 11 1 13 16 15 13 0 13 1 9 9 10 9 10 0 7 16 13 1 9 0 1 9 10 9 2
19 8 8 11 13 1 9 16 9 9 10 9 7 10 9 13 1 10 9 2
37 15 13 16 10 9 13 1 2 9 9 11 7 13 1 9 16 15 15 13 2 7 13 16 11 13 1 15 1 9 16 13 0 1 9 10 12 2
16 2 13 13 13 1 10 9 16 13 1 15 9 1 9 15 2
10 15 3 4 16 11 13 1 9 15 2
32 15 16 13 1 15 1 10 9 13 14 9 15 1 9 15 2 7 11 13 10 0 16 4 13 9 1 10 9 14 9 2 2
56 9 11 11 2 9 9 9 9 2 9 1 9 9 11 2 13 3 16 1 9 15 13 9 9 0 2 16 1 15 13 9 10 9 10 0 1 9 0 16 13 1 15 9 9 7 9 0 1 2 9 9 16 13 10 9 2
17 3 9 10 9 10 0 13 9 2 16 10 9 1 15 13 0 2
40 9 9 15 13 13 16 1 9 10 9 7 9 15 13 3 9 9 1 10 9 10 0 2 1 10 9 7 1 10 9 2 7 3 3 9 9 7 9 15 2
40 1 9 10 9 13 3 9 15 14 9 10 9 10 0 2 1 2 3 9 14 9 9 14 10 9 1 10 9 2 1 10 9 16 13 1 10 9 10 0 2
50 9 9 13 1 9 10 9 7 10 9 2 11 11 2 7 1 9 9 11 2 11 11 2 1 9 9 10 9 1 10 9 1 9 10 9 2 16 13 1 9 10 9 1 9 9 14 9 10 9 2
37 3 13 9 10 9 1 9 9 10 9 7 9 10 9 13 9 0 1 10 9 1 9 9 1 9 14 12 9 1 10 10 9 1 9 10 9 2
41 9 10 1 9 10 9 1 10 9 2 13 11 1 9 9 10 9 2 9 11 11 2 7 13 1 15 16 10 9 3 13 9 1 10 9 1 13 1 9 15 2
11 11 13 16 9 1 9 12 9 0 3 2
23 11 13 1 10 9 7 13 14 11 13 1 9 15 10 0 14 10 9 2 1 9 11 2
31 9 10 9 2 10 9 11 11 7 9 9 10 9 11 11 2 13 1 10 9 11 7 13 1 15 1 9 15 14 11 2
13 11 13 1 11 7 13 1 15 13 9 1 9 2
28 15 13 16 1 9 13 1 9 7 13 4 13 1 9 15 1 9 16 13 1 9 9 15 1 9 9 9 2
13 11 13 16 10 9 13 9 1 9 15 10 0 2
25 10 9 13 3 14 10 9 1 9 9 10 9 7 1 9 15 13 9 9 10 9 7 10 9 2
38 12 1 10 9 13 13 14 9 10 9 7 10 9 13 14 9 10 9 10 1 16 13 13 14 9 10 9 2 1 0 1 10 13 1 9 10 9 2
9 9 0 13 13 14 9 10 9 2
17 9 15 13 13 1 9 9 10 9 14 10 9 1 9 1 9 2
14 9 10 9 13 3 1 9 10 9 1 9 10 9 2
11 10 10 9 13 13 3 14 9 10 9 2
19 9 11 11 2 11 13 16 1 10 9 13 9 0 1 9 9 10 9 2
17 1 10 9 13 9 10 9 1 2 9 2 9 11 2 11 2 2
17 3 13 9 15 1 2 9 9 2 14 9 10 9 7 10 9 2
13 15 13 16 9 9 10 9 13 1 9 10 9 2
36 9 11 9 13 16 13 9 0 1 9 9 10 9 2 7 7 13 1 9 16 1 15 9 10 9 1 10 9 13 1 7 1 1 10 13 2
26 11 13 10 9 10 0 16 13 14 9 10 9 1 12 1 11 12 7 1 3 1 9 14 12 9 2
10 10 9 1 15 13 9 14 10 9 2
27 10 9 1 9 10 9 1 10 9 2 11 11 2 13 16 10 10 9 1 11 13 1 9 1 10 9 2
13 9 10 9 13 7 7 10 9 1 15 13 3 2
16 1 15 2 13 10 3 9 16 9 15 13 3 1 10 9 2
27 7 2 1 9 15 10 9 13 3 1 10 9 7 3 4 10 9 13 14 9 10 9 7 9 10 9 2
15 11 13 16 9 10 9 1 11 0 1 10 9 1 11 2
20 1 9 9 9 2 15 13 1 9 10 9 2 7 3 1 9 1 9 0 2
25 9 10 9 2 11 11 2 13 16 1 11 2 11 13 9 9 14 12 9 1 10 9 10 0 2
10 11 3 13 14 10 9 1 9 15 2
21 1 11 13 1 9 9 1 9 10 9 2 16 13 14 9 15 1 11 2 11 2
20 11 13 3 16 1 3 13 9 9 14 1 12 12 16 1 9 9 10 9 2
28 7 9 10 9 13 1 9 1 9 15 10 0 2 7 16 1 9 1 9 10 9 13 9 14 12 12 16 2
9 1 10 16 13 1 9 10 9 2
11 13 1 15 9 1 10 9 7 10 9 2
32 1 10 9 10 0 13 1 10 9 7 1 10 11 9 9 16 13 13 1 10 9 13 14 10 9 10 0 1 9 10 9 2
20 10 9 13 13 7 13 1 10 9 10 0 2 1 10 16 13 1 15 2 2
35 9 15 13 3 9 10 9 2 11 11 2 1 9 9 16 13 10 9 10 0 1 9 1 9 10 9 10 0 7 9 15 1 10 9 2
35 3 13 9 10 9 2 16 1 9 12 4 9 0 1 10 9 10 0 7 1 9 10 9 14 10 9 2 1 2 9 1 10 9 2 2
40 10 9 10 0 1 9 10 9 13 1 12 12 9 2 7 13 1 3 1 12 12 2 7 1 9 11 10 9 1 9 10 9 13 10 9 13 9 1 9 2
36 1 9 15 2 13 1 10 9 10 0 9 0 2 16 13 9 14 9 11 7 9 9 1 10 9 10 0 2 7 10 9 3 3 3 0 2
43 1 9 15 1 9 10 9 13 11 9 0 1 10 9 16 13 1 16 9 10 9 13 14 10 9 2 1 16 10 9 14 9 10 9 1 9 7 9 0 13 1 9 2
41 2 13 10 9 13 1 9 1 11 9 0 14 12 9 1 9 2 14 10 9 10 0 1 9 9 1 9 10 9 13 1 12 12 9 1 9 2 2 13 11 2
33 9 9 11 2 10 9 11 11 2 13 16 9 10 9 13 3 1 9 9 7 9 14 9 10 9 2 16 16 13 1 9 0 2
20 2 1 9 7 1 9 1 9 10 9 2 10 9 3 13 2 2 13 11 2
17 2 1 9 10 9 13 9 0 1 9 10 9 1 10 9 15 2
16 7 10 9 3 13 13 1 9 12 2 13 15 9 0 2 2
19 9 10 9 2 11 11 2 13 16 3 13 1 10 9 9 14 9 9 2
48 1 9 15 2 13 1 10 9 9 0 2 7 15 3 13 14 9 10 9 1 10 9 2 1 9 9 1 9 10 9 1 10 10 9 2 9 9 10 9 1 9 7 9 1 9 10 9 2
26 9 9 10 9 2 11 11 2 13 16 9 10 9 1 9 9 10 9 13 0 2 7 16 9 0 2
44 2 10 9 13 13 2 9 10 9 0 3 7 3 0 2 7 3 13 13 1 9 15 14 9 10 9 7 10 9 2 11 11 2 1 9 10 9 7 10 9 1 15 2 2
48 3 13 9 1 9 10 9 2 9 9 10 9 11 11 2 10 9 11 11 1 9 9 2 9 2 9 9 10 9 9 11 11 2 9 9 11 11 11 2 7 9 9 10 9 9 11 11 2
34 9 9 11 13 1 10 9 10 0 1 9 1 9 9 10 9 16 13 1 9 0 2 3 16 15 4 13 1 9 0 1 10 9 2
41 14 10 9 13 10 9 1 10 9 2 1 9 16 1 10 9 10 0 13 10 9 13 14 9 10 9 10 0 14 15 1 10 9 10 0 16 13 1 10 9 2
35 10 9 13 3 1 9 10 9 16 13 1 9 12 2 1 15 4 13 14 9 10 9 14 10 9 10 0 1 10 16 13 1 9 0 2
22 1 9 15 13 16 4 16 1 10 9 10 0 13 9 0 0 1 9 9 10 9 2
18 10 9 16 13 7 10 9 13 1 9 1 9 9 10 9 2 9 2
26 3 16 13 1 10 9 13 3 10 9 1 9 2 16 9 15 13 1 3 1 9 10 9 14 15 2
28 9 0 2 16 13 1 10 9 1 9 10 9 1 9 10 9 2 13 15 1 3 1 9 0 1 10 9 2
4 9 0 3 2
13 13 1 9 0 0 2 16 13 1 9 9 9 2
28 9 10 9 11 13 9 0 14 12 9 2 11 12 9 2 11 12 9 2 11 12 9 2 7 11 12 9 2
22 3 0 7 3 9 10 9 14 10 9 10 0 2 7 11 7 11 2 13 9 0 2
22 10 9 10 0 13 12 12 9 1 9 2 9 11 2 1 9 9 11 1 10 9 2
16 1 10 9 13 12 9 0 1 9 9 10 13 1 9 9 2
27 7 13 1 15 3 9 1 12 9 16 13 1 9 1 10 9 2 9 9 7 1 10 9 1 10 15 2
27 10 9 1 15 13 1 10 9 10 0 13 1 9 15 14 9 1 9 0 2 9 2 9 9 7 9 2
38 1 9 15 13 1 9 10 9 10 0 13 9 1 10 9 2 7 13 1 9 0 14 9 1 11 7 2 9 2 1 10 9 10 0 11 7 9 2
36 9 1 9 1 9 9 11 2 16 13 9 9 1 9 2 9 9 7 9 1 10 9 2 13 1 11 10 0 2 1 9 14 12 12 9 2
26 1 10 9 9 10 11 2 10 9 10 0 7 9 9 2 16 9 15 1 10 9 13 10 0 3 2
11 1 3 13 10 9 10 0 12 9 9 2
4 2 11 2 2
39 9 9 10 9 1 9 2 9 13 3 9 9 1 2 9 7 9 0 1 11 11 7 11 11 2 9 9 10 9 7 10 9 11 9 7 9 0 9 2
10 11 7 11 13 1 9 9 1 9 2
33 1 9 10 9 2 13 10 9 13 9 1 9 12 9 16 13 1 9 9 2 16 13 14 9 15 1 9 9 1 9 9 9 2
13 3 2 3 13 10 9 10 9 1 9 10 9 2
16 11 13 1 12 9 9 1 2 9 7 1 9 14 12 9 2
15 11 13 1 12 9 9 1 2 9 7 9 14 12 9 2
7 9 11 13 1 12 9 2
14 11 7 11 13 14 9 10 9 1 9 9 9 0 2
25 9 1 15 13 1 9 9 9 1 9 9 10 9 2 11 11 2 1 9 9 7 9 1 11 2
52 1 9 2 7 9 16 13 3 1 11 13 16 1 9 9 1 11 1 9 9 10 9 10 0 14 11 2 11 2 13 16 1 10 12 1 11 1 10 12 1 11 13 1 11 9 14 12 9 9 1 11 2
12 14 10 9 13 9 9 10 9 1 10 9 2
32 9 10 9 13 1 9 10 9 2 7 7 13 14 9 10 9 1 9 0 2 1 15 4 13 1 9 10 9 2 11 11 2
32 12 9 9 1 11 13 1 9 9 14 11 1 11 2 16 13 1 9 9 9 9 10 9 7 10 9 14 11 2 11 2 2
11 10 9 13 1 9 9 11 2 11 11 2
15 1 10 9 13 9 9 11 7 3 9 9 0 1 11 2
10 9 10 9 13 1 9 10 9 11 2
31 9 9 10 9 13 1 9 15 1 10 13 2 16 1 10 9 1 11 13 12 9 2 13 10 9 1 11 12 9 11 2
28 1 9 11 2 13 1 9 10 9 1 9 10 9 14 11 2 16 13 13 7 13 14 11 1 9 9 12 2
29 2 11 2 2 9 10 9 1 9 0 2 13 14 9 15 1 9 11 1 9 9 2 7 9 14 12 12 9 2
33 1 2 10 9 2 13 16 3 1 12 10 9 10 0 14 10 9 2 1 10 9 10 0 1 9 9 7 1 11 2 13 9 2
22 10 9 13 1 9 15 14 9 10 9 11 11 16 13 1 9 11 11 9 7 9 2
14 10 9 13 1 1 9 9 1 9 11 12 9 9 2
31 10 9 2 1 9 14 1 12 9 13 1 9 15 14 9 10 9 11 11 2 10 9 14 9 1 9 7 9 9 9 2
24 9 10 9 13 13 9 9 14 1 12 9 1 9 2 7 12 9 1 9 2 3 13 9 2
22 15 13 1 9 10 9 2 16 13 1 10 9 1 9 9 0 2 1 12 12 9 2
19 10 9 13 14 10 9 1 11 11 16 13 14 10 9 1 9 14 9 2
21 3 13 11 1 2 10 9 2 16 9 10 9 13 1 12 9 1 9 10 9 2
27 15 13 13 9 9 7 13 1 9 0 1 11 11 2 16 13 1 9 10 9 13 9 9 1 10 9 2
19 9 10 9 13 1 11 13 14 9 10 9 1 12 9 2 7 11 13 2
35 1 9 0 7 9 7 9 13 3 10 9 1 9 9 1 15 13 10 9 1 11 1 12 1 11 7 13 10 9 10 0 1 10 9 2
24 1 2 10 9 2 13 16 3 12 10 9 10 0 14 10 9 1 9 1 9 9 1 9 2
40 9 9 10 9 1 9 10 9 11 11 2 11 2 13 13 14 10 9 7 13 10 9 14 9 10 9 10 0 13 1 9 12 9 1 9 11 1 9 0 2
71 9 9 11 13 1 9 15 9 1 9 9 10 9 10 0 2 11 9 2 16 1 15 15 13 16 10 9 13 9 15 1 9 11 1 9 0 2 13 9 1 9 10 9 7 9 1 10 9 14 10 9 2 2 16 15 9 1 10 9 10 0 14 10 9 2 2 1 9 10 9 2
51 10 9 13 1 9 15 13 9 1 10 9 1 9 10 9 7 3 1 9 0 14 9 15 7 3 13 1 10 9 13 1 9 1 9 15 13 1 9 9 14 10 9 7 15 1 9 0 1 9 0 2
78 9 15 14 9 10 9 1 9 9 10 9 10 0 13 1 9 1 10 9 16 9 10 9 13 1 9 10 9 11 11 7 1 9 10 9 11 11 2 1 12 9 2 16 1 15 13 16 9 1 9 10 9 16 13 1 10 9 1 9 9 2 13 1 10 9 1 9 13 2 16 16 13 1 9 2 11 2 2
11 10 9 13 3 1 12 9 1 9 11 2
24 12 9 1 10 9 13 1 11 2 9 9 14 11 9 7 12 9 1 10 9 13 10 9 2
37 9 9 10 9 10 0 13 3 1 9 2 16 10 9 3 13 14 9 15 1 9 10 9 7 7 9 15 1 9 0 14 9 13 2 0 2 2
29 1 9 15 2 9 15 14 10 9 1 10 9 1 9 0 2 13 1 10 9 2 7 7 15 13 13 1 15 2
19 9 13 16 12 9 0 2 0 7 0 2 13 1 9 9 1 10 9 2
27 9 10 9 11 11 7 9 10 9 11 11 13 13 3 1 9 0 1 9 9 9 1 10 9 10 0 2
19 10 9 10 9 3 13 2 7 15 13 16 10 13 1 10 9 10 0 2
48 10 9 13 1 10 9 13 1 9 0 1 9 10 9 3 3 1 10 9 16 13 1 15 3 2 7 7 3 1 9 0 1 15 13 9 9 2 1 9 9 9 10 9 7 9 10 9 2
23 9 10 9 1 9 0 2 11 11 2 13 3 1 11 1 9 10 9 10 0 10 0 2
28 9 15 2 11 11 2 13 9 1 9 13 14 9 10 9 1 9 0 1 9 0 2 7 3 1 9 0 2
19 3 13 9 15 14 10 9 10 0 7 11 13 9 9 2 1 15 13 2
59 1 13 1 9 10 9 1 10 9 2 13 1 10 9 10 0 3 9 9 0 2 13 11 16 10 9 13 4 13 1 9 9 16 13 1 9 0 2 3 3 16 10 9 1 9 15 13 0 1 9 10 9 10 0 7 1 9 0 2
26 16 1 9 10 9 2 13 14 9 10 9 1 9 9 2 13 9 13 14 9 10 9 16 1 15 2
17 9 15 13 12 9 1 9 1 9 9 2 1 12 9 1 3 2
6 9 0 13 12 9 2
12 1 3 13 10 9 1 9 15 1 12 9 2
19 1 9 11 13 9 10 9 10 0 7 10 9 13 14 9 9 10 9 2
26 9 10 9 13 9 0 1 9 9 1 9 11 11 1 11 9 9 10 9 10 0 3 1 9 15 2
23 1 9 9 10 9 13 3 9 12 9 9 2 7 1 15 9 1 9 9 1 9 11 2
10 10 9 13 1 3 12 12 9 9 2
18 3 13 10 9 12 9 9 0 1 11 1 9 9 10 9 10 0 2
16 1 10 9 16 13 10 9 13 10 9 10 9 1 10 9 2
26 3 13 9 11 7 11 2 9 9 1 9 10 9 7 9 0 11 2 11 2 1 9 1 9 0 2
10 11 2 0 1 2 10 9 2 2 2
26 1 10 9 10 0 3 1 11 13 3 10 9 2 0 2 10 9 2 7 1 15 13 9 10 9 2
40 10 9 2 16 13 9 11 11 7 10 13 1 9 14 12 9 2 13 1 2 9 10 9 11 10 0 2 1 10 9 16 13 1 9 15 2 11 7 11 2
33 9 10 9 14 11 11 13 3 12 9 14 9 9 3 16 13 1 3 12 9 1 10 9 14 10 9 14 11 1 12 9 3 2
15 10 9 13 9 0 1 9 10 9 7 10 9 10 0 2
14 1 10 9 13 12 9 2 7 13 1 15 12 9 2
26 10 9 11 2 16 13 1 15 9 0 3 1 11 2 13 1 9 10 9 10 0 3 1 11 11 2
27 9 10 9 1 11 13 10 0 3 16 13 1 15 1 3 2 7 15 13 1 15 3 1 12 12 9 2
36 1 13 9 1 15 2 1 9 14 9 9 1 11 7 9 9 1 9 2 13 10 9 1 1 9 9 1 11 1 9 14 1 12 12 9 2
80 10 9 11 11 1 9 2 10 9 1 10 9 1 9 2 9 13 9 9 3 13 10 9 1 9 9 1 10 9 1 9 9 12 1 9 2 9 2 1 1 10 9 16 13 1 9 15 1 10 12 1 11 2 1 15 13 9 15 14 10 9 3 14 10 9 13 14 10 9 10 0 1 9 9 9 1 10 9 9 2
23 10 9 13 3 1 16 13 1 9 10 9 13 14 10 9 1 9 2 10 9 11 11 2
32 11 11 11 13 1 12 9 9 7 9 10 9 14 9 2 9 14 10 9 10 0 16 13 1 9 2 9 1 10 9 9 2
43 11 13 1 9 15 1 9 1 10 9 2 1 9 9 12 2 1 2 9 9 10 9 9 10 9 2 1 16 13 1 15 9 9 13 1 9 0 14 3 1 12 9 2
30 1 15 2 1 9 12 2 13 11 2 1 9 11 11 2 9 1 9 2 10 9 1 10 9 1 9 1 10 9 2
54 11 13 13 15 3 1 9 9 10 9 1 9 2 7 13 1 15 9 1 9 9 15 10 4 1 10 9 2 9 9 0 1 9 10 9 2 9 9 2 9 9 0 7 3 2 1 9 0 14 1 12 12 9 2
38 10 9 13 3 13 14 9 9 1 10 9 1 9 2 9 1 9 14 12 12 9 2 1 13 16 1 11 13 1 3 13 10 9 1 9 16 13 2
24 1 9 1 9 2 10 9 13 9 11 11 16 10 9 10 0 13 13 7 13 3 9 0 2
21 3 2 13 1 9 2 7 9 10 9 13 1 10 9 3 1 1 12 12 9 2
31 3 2 1 16 13 9 2 9 0 1 9 2 10 9 10 0 1 9 2 7 3 1 9 7 1 9 2 13 9 0 2
7 9 10 9 4 13 3 2
28 1 15 2 10 9 13 9 1 10 9 9 1 10 9 7 13 13 1 11 1 9 9 1 10 9 1 15 2
9 1 2 15 13 10 9 1 9 2
52 9 10 9 1 9 11 2 11 11 2 13 1 9 1 9 10 9 7 10 9 13 1 9 10 9 1 9 13 2 16 4 13 1 15 9 2 7 1 15 13 15 1 9 13 1 9 9 0 7 9 0 2
49 11 13 16 1 9 11 13 1 9 10 9 1 11 9 1 9 9 9 0 1 10 9 2 7 14 9 10 9 13 1 9 9 13 7 0 16 13 3 1 10 9 2 7 3 1 9 10 9 2
59 1 10 9 10 0 14 9 10 9 1 9 11 16 13 3 13 16 1 10 9 10 0 13 9 1 10 9 1 9 1 9 10 9 2 3 9 1 9 3 0 2 7 1 10 9 10 0 16 13 1 13 10 9 2 10 9 13 0 2
39 1 10 9 13 16 9 9 10 9 1 9 9 11 2 13 1 10 9 10 0 9 1 9 1 9 10 9 14 9 10 9 1 9 13 9 1 9 15 2
56 9 10 9 2 11 11 2 13 16 3 12 9 2 1 15 12 9 7 12 9 0 2 13 1 10 9 10 0 1 9 0 1 9 10 9 16 13 1 9 9 1 9 11 1 9 10 9 2 7 9 10 9 7 10 9 2
16 10 9 10 0 14 9 11 1 11 13 9 9 1 9 11 2
23 1 9 16 13 3 1 9 10 9 1 11 2 13 1 10 9 1 12 1 9 10 9 2
25 10 9 13 13 1 9 11 10 0 7 13 1 15 9 9 9 11 7 1 15 9 9 7 9 2
30 1 9 10 9 13 10 9 13 9 9 1 9 11 1 9 11 7 9 1 9 10 9 2 9 10 9 7 9 11 2
5 11 2 11 2 2
37 9 9 13 1 11 2 11 10 0 7 11 2 13 3 9 0 1 10 9 16 13 1 9 11 2 16 9 15 9 13 9 1 10 9 10 0 2
29 2 10 9 13 16 13 3 9 0 2 2 13 9 10 9 14 11 2 11 11 2 1 9 15 14 12 9 13 2
39 2 4 13 9 1 10 9 2 2 13 1 16 13 1 10 9 14 9 10 12 2 8 2 16 13 1 9 10 9 14 10 9 10 3 2 13 1 12 2
72 9 10 9 10 0 2 11 11 2 13 9 0 1 10 9 16 1 9 11 1 11 2 1 13 16 15 13 9 16 13 13 13 14 2 9 11 2 1 9 11 2 1 9 15 14 9 12 9 2 16 13 1 15 9 9 1 9 9 10 9 14 9 10 9 7 10 9 1 12 1 11 2
39 10 9 10 0 14 11 2 11 11 2 13 1 15 3 9 14 12 9 2 1 9 13 14 10 9 1 9 10 9 1 9 9 16 13 14 9 10 9 2
12 11 2 11 2 0 1 2 10 9 2 2 2
39 1 11 11 2 11 16 13 1 9 1 11 11 13 3 1 10 9 9 9 1 9 1 9 12 2 9 1 9 2 9 0 7 9 3 0 14 9 9 2
35 9 1 9 12 13 10 9 10 0 3 16 1 15 4 13 9 1 9 1 9 11 2 11 2 16 13 13 1 9 14 9 9 10 9 2
27 9 10 9 13 1 9 15 14 10 9 1 9 10 13 2 11 2 1 11 2 3 15 13 1 9 15 2
25 10 9 16 1 15 13 11 2 11 2 16 13 1 9 9 7 9 9 2 13 1 9 0 0 2
20 9 15 10 0 2 11 2 13 1 9 15 0 1 9 0 0 0 7 9 2
37 9 15 14 10 9 2 11 11 2 13 3 14 10 9 16 13 13 14 10 9 1 9 11 1 12 9 2 1 16 13 9 0 0 3 13 15 2
21 10 9 2 16 3 13 4 13 1 9 15 2 13 1 9 15 1 9 9 0 2
7 15 13 16 13 14 11 2
21 1 9 9 1 9 16 1 15 13 11 2 11 2 13 10 9 13 16 13 3 2
28 1 9 9 3 13 10 9 16 13 1 10 9 2 11 11 2 16 4 16 10 9 1 10 9 3 13 3 2
40 1 9 9 11 2 11 13 9 10 9 10 0 1 9 1 10 9 7 9 10 9 2 11 2 11 2 16 13 13 7 1 10 9 13 9 3 2 0 15 2
13 1 3 3 13 10 9 1 15 13 10 9 0 2
23 12 10 9 13 16 11 11 2 11 2 9 10 9 2 13 16 9 15 13 3 1 9 2
31 10 9 1 10 9 13 16 13 16 11 2 11 13 9 9 2 7 1 9 15 13 9 0 14 9 16 13 1 9 9 2
11 10 9 13 3 0 1 9 9 1 11 2
16 1 10 9 16 13 1 9 15 3 13 9 1 9 9 9 2
38 10 9 10 0 1 9 9 10 11 2 16 1 15 13 1 2 9 10 9 11 2 11 1 11 2 13 7 7 3 13 10 9 13 3 13 14 15 2
29 1 12 1 9 15 14 11 2 11 13 10 9 9 7 1 15 9 0 1 10 9 10 0 2 0 1 9 11 2
40 10 9 16 13 0 16 13 1 9 15 2 1 9 1 10 9 1 9 11 1 11 2 11 2 13 1 2 9 10 9 2 7 13 16 15 13 9 9 0 2
33 3 13 16 10 9 13 1 9 15 1 9 11 2 11 2 16 1 15 13 1 9 9 7 9 1 9 10 9 10 0 1 11 2
32 1 9 10 9 2 11 11 2 2 9 1 10 9 13 11 2 11 4 13 1 9 9 15 10 0 1 9 10 9 1 11 2
27 10 9 13 2 1 9 9 1 9 10 9 10 0 2 16 11 2 11 13 1 9 14 13 1 10 9 2
20 9 10 9 13 16 1 10 9 16 1 10 9 13 11 2 11 12 9 9 2
10 8 13 1 1 9 2 13 1 11 2
14 3 13 1 9 2 10 9 2 9 1 9 14 11 2
33 1 10 9 13 1 9 2 10 9 2 11 2 9 10 9 2 7 13 16 9 1 9 15 13 1 9 15 1 10 9 10 0 2
22 1 9 15 2 13 14 11 1 9 0 1 10 9 2 7 13 14 15 13 1 15 2
14 11 13 13 1 9 16 13 1 9 7 1 9 15 2
17 10 16 13 4 13 13 2 2 15 13 2 7 15 10 9 2 2
31 9 9 10 9 2 1 9 9 2 10 9 11 14 11 2 13 3 1 9 2 10 9 10 0 1 9 1 9 10 9 2
34 10 9 13 1 9 2 10 9 9 9 2 9 0 2 1 15 13 9 1 9 9 14 9 1 9 16 13 1 15 1 9 10 9 2
40 10 9 2 1 9 12 2 13 16 10 1 13 10 9 1 10 9 1 9 10 9 1 9 2 13 9 10 9 4 13 1 9 9 10 9 14 9 10 9 2
27 10 9 1 10 9 1 9 10 9 13 1 12 2 7 7 3 13 9 10 9 13 1 9 9 10 9 2
44 10 9 10 0 14 9 10 9 2 11 11 2 13 16 10 9 13 4 13 1 10 13 2 7 16 9 9 10 9 13 3 1 9 2 7 9 1 9 10 9 1 10 9 2
25 1 9 1 15 13 10 9 1 9 2 7 9 1 9 10 9 2 7 1 10 9 13 9 0 2
34 10 9 1 10 9 3 13 14 10 9 2 16 13 16 9 10 9 13 13 14 9 15 1 10 9 2 7 16 13 9 1 9 0 2
24 9 10 9 13 2 1 15 2 16 10 9 1 10 9 13 4 1 15 13 3 14 9 15 2
14 10 9 1 9 2 10 9 3 13 1 9 9 15 2
33 9 9 10 9 1 11 2 11 11 2 13 1 9 0 14 9 10 9 1 10 9 2 7 1 9 9 10 9 1 9 10 9 2
24 3 2 13 11 2 4 13 3 14 10 9 1 9 10 9 2 16 3 3 13 9 10 9 2
3 2 12 2
26 9 15 2 16 13 1 10 9 1 10 9 2 10 9 2 2 13 1 2 9 9 10 9 10 0 2
40 1 10 9 10 0 10 9 3 7 3 13 2 1 16 9 15 13 1 9 9 10 9 11 14 11 2 16 13 1 10 9 1 10 9 1 9 9 10 9 2
44 9 15 2 16 4 9 3 1 9 0 2 3 3 1 9 0 2 13 13 1 10 12 1 9 15 14 9 15 10 0 2 1 10 9 1 9 10 9 1 9 9 7 9 2
19 10 9 13 13 1 10 9 13 14 9 10 9 16 15 13 13 1 15 2
33 3 1 15 10 9 13 14 9 10 9 1 9 9 14 10 9 16 13 1 9 9 7 10 13 9 0 1 15 14 9 10 9 2
27 10 9 3 4 1 10 9 13 7 1 9 15 1 9 9 3 7 9 0 16 13 3 9 9 7 9 2
18 9 9 11 14 11 13 14 9 10 9 13 1 9 1 9 10 9 2
22 11 11 2 9 10 9 2 13 1 9 1 9 9 10 9 7 3 1 9 9 9 2
18 13 1 9 15 16 15 13 14 10 9 14 10 9 1 15 15 13 2
25 1 15 2 13 9 10 9 1 13 1 9 1 10 9 1 9 9 9 10 0 16 9 15 13 2
32 3 13 10 9 1 9 1 12 10 9 10 0 16 13 1 9 0 2 9 2 1 15 12 16 13 1 15 13 1 10 9 2
29 9 1 9 15 13 3 1 9 10 9 7 0 13 9 16 0 3 1 9 9 2 1 15 13 9 7 9 9 2
43 10 9 10 0 14 9 9 10 9 10 0 1 9 11 1 11 2 13 13 1 12 9 9 1 9 15 10 0 14 12 9 15 2 1 10 9 16 13 14 9 10 9 2
34 9 10 9 13 13 9 0 2 1 1 9 9 0 10 4 1 9 15 1 9 15 1 9 15 14 10 9 7 1 9 13 9 9 2
21 9 15 3 13 1 9 15 1 10 9 10 0 10 0 14 9 10 9 10 0 2
26 9 9 9 9 13 3 9 9 1 9 13 0 9 2 1 2 9 10 9 10 0 16 0 1 11 2
27 9 10 9 10 0 13 1 9 9 10 9 1 9 9 10 9 2 16 13 9 1 9 14 12 12 9 2
16 10 9 13 16 13 1 9 9 10 13 1 10 9 10 0 2
28 9 10 9 2 11 11 2 13 14 9 15 14 10 9 10 0 1 9 10 9 1 9 10 9 7 10 9 2
18 1 9 12 9 0 1 10 9 2 11 11 2 11 11 7 9 11 2
13 11 2 1 11 2 13 1 9 9 1 9 0 2
15 1 10 9 12 13 1 9 9 10 9 1 9 9 0 2
21 9 11 1 11 13 9 9 11 7 11 9 16 13 1 9 10 9 1 9 12 2
10 15 13 14 10 9 14 15 1 9 2
22 9 15 10 0 1 11 13 1 9 15 1 9 9 9 9 11 10 0 2 11 11 2
11 15 13 1 9 10 9 0 7 0 0 2
21 1 10 9 13 16 1 10 12 1 12 10 9 10 0 13 9 0 1 11 11 2
68 9 10 9 13 1 9 9 15 14 9 15 16 13 13 9 1 10 9 2 1 9 10 9 7 10 9 1 9 15 14 9 10 9 7 10 9 1 10 9 10 9 7 10 9 13 1 9 9 9 15 1 9 12 12 9 9 1 9 0 7 9 0 1 10 9 10 9 2
28 13 16 9 10 9 14 10 9 7 9 10 9 1 9 1 9 10 9 1 9 14 1 12 12 9 2 9 2
60 9 10 9 13 1 10 9 7 1 9 10 9 13 1 9 10 9 14 15 13 15 13 1 9 14 9 0 1 9 16 13 1 15 1 2 9 9 10 9 2 7 1 9 14 9 0 16 13 12 1 10 9 16 13 1 2 9 10 9 2
37 1 9 15 1 9 10 9 13 9 10 9 2 11 11 2 16 10 9 14 9 0 14 10 9 1 10 9 13 9 0 1 10 9 1 9 15 2
37 1 10 9 13 16 1 9 15 4 9 10 9 7 10 9 13 3 1 10 10 9 7 3 13 9 0 1 9 9 2 9 1 9 1 9 15 2
30 11 1 11 2 11 1 11 7 11 2 11 2 9 11 1 9 2 10 9 13 9 1 9 7 9 1 9 10 9 2
13 1 10 9 13 9 1 9 7 1 9 14 9 2
8 11 11 13 9 14 9 11 2
15 11 2 11 2 9 11 13 9 1 9 11 9 11 11 2
30 10 9 13 16 13 14 10 9 10 0 2 16 13 11 2 11 2 11 2 1 9 1 9 1 9 10 9 14 9 2
27 10 9 1 9 10 9 13 0 1 11 2 1 11 10 0 2 1 10 9 10 0 7 1 11 2 13 2
10 11 2 0 1 2 10 9 2 2 2
71 9 11 2 9 9 12 2 16 13 1 9 11 1 9 11 1 10 9 2 13 9 1 9 0 2 15 10 9 10 0 16 13 1 9 15 16 13 13 1 10 9 10 0 2 15 10 9 10 0 1 10 9 2 7 15 10 9 10 0 3 16 13 3 2 3 1 10 9 10 0 2
21 11 13 3 1 9 12 9 9 10 9 7 10 11 7 9 10 9 7 10 9 2
38 7 12 9 1 10 9 1 15 13 1 10 9 10 12 14 10 9 2 16 13 1 9 0 3 2 13 3 1 1 9 15 14 12 10 9 3 3 2
13 13 16 11 13 1 10 9 3 1 9 10 9 2
20 15 13 0 1 10 9 10 0 3 1 9 15 1 9 10 9 7 10 9 2
35 3 1 9 15 13 7 13 16 13 1 9 9 7 9 9 9 12 9 0 1 15 13 3 10 9 10 0 7 3 1 9 1 9 11 2
28 7 1 10 9 10 0 2 3 15 13 1 10 9 1 9 15 2 7 15 13 3 1 10 9 3 13 9 2
13 2 13 13 1 10 12 1 10 9 2 2 13 2
55 10 9 10 0 14 15 2 11 11 1 10 9 10 0 2 13 13 1 9 9 9 10 9 9 1 10 9 2 1 9 9 0 2 7 1 9 16 9 10 9 10 0 13 3 2 9 1 10 9 7 13 1 9 15 2
7 9 11 13 1 12 9 2
14 13 1 15 9 0 2 7 1 9 15 9 0 0 2
32 10 9 16 15 13 1 9 10 9 9 15 2 1 9 9 2 13 1 15 9 0 0 1 7 16 15 13 13 1 10 9 2
46 9 9 10 11 10 0 1 9 2 1 9 12 10 0 1 10 9 1 9 9 1 10 9 10 0 2 1 1 9 2 13 9 0 0 1 9 0 0 1 15 13 10 9 10 0 2
6 10 9 16 13 0 2
30 10 9 1 9 7 10 9 10 0 16 13 1 15 2 13 1 9 9 2 1 9 1 9 0 1 9 7 9 0 2
13 10 9 13 13 9 2 3 4 13 0 3 3 2
19 4 13 1 9 16 9 10 9 10 9 13 0 7 1 10 9 10 0 2
26 14 3 16 13 13 9 10 9 1 9 2 11 11 2 1 2 9 9 2 7 3 2 9 0 2 2
23 3 3 15 2 9 10 9 1 9 1 2 12 13 1 9 0 1 9 12 1 12 9 2
14 9 10 9 16 13 13 3 3 1 2 12 12 9 2
12 1 2 12 12 1 10 9 1 9 10 9 2
6 10 9 13 12 9 2
5 10 9 9 0 2
8 9 12 0 2 12 12 9 2
8 12 9 1 10 9 1 9 2
11 13 16 13 9 0 1 9 12 9 3 2
13 1 10 9 10 0 3 13 9 10 9 12 9 2
8 12 1 15 13 1 9 9 2
32 1 10 9 2 13 10 9 1 9 3 9 0 2 10 9 1 9 0 2 9 9 2 9 1 9 9 2 9 9 1 9 2
11 3 13 9 9 7 9 1 10 10 9 2
5 15 13 10 9 2
5 8 8 8 13 2
10 11 2 2 15 9 14 3 16 13 2
22 1 12 15 13 3 12 9 1 10 2 12 12 2 16 3 3 13 3 9 10 9 2
9 10 9 13 1 2 12 7 12 2
14 3 15 13 1 9 1 2 12 9 1 9 9 2 2
14 11 13 1 9 14 9 0 7 13 2 2 15 13 2
13 13 13 13 1 9 0 7 3 13 3 1 15 2
8 1 15 10 9 0 3 2 2
21 13 1 10 9 1 9 9 9 9 14 12 12 9 2 1 9 16 13 12 12 2
7 13 1 15 1 12 12 2
18 13 9 13 1 9 16 10 9 13 16 3 1 15 15 3 4 13 2
11 13 16 1 10 9 13 12 8 2 8 2
16 3 2 1 3 1 9 0 2 9 10 9 13 12 12 9 2
11 13 1 2 12 9 7 13 9 10 9 2
17 8 8 8 1 9 9 1 10 9 10 9 2 3 13 1 9 2
5 15 13 9 0 2
6 10 9 4 13 3 2
10 4 13 1 9 12 16 16 15 13 2
7 3 9 9 13 9 0 2
9 1 10 9 16 0 3 4 13 2
11 1 10 9 10 15 3 9 0 3 13 2
9 3 4 13 9 7 9 1 9 2
4 13 9 9 2
6 13 9 1 10 9 2
5 10 9 3 13 2
8 15 13 1 10 9 10 0 2
4 10 9 13 2
25 13 9 1 9 16 13 4 2 7 3 13 9 2 16 15 3 13 1 9 9 9 7 9 11 2
22 10 9 2 13 10 9 1 9 1 3 2 1 10 9 7 10 10 9 13 1 9 2
22 10 9 14 9 13 1 9 10 9 16 13 2 10 13 1 10 9 7 3 10 9 2
9 10 9 13 12 1 9 9 13 2
2 8 2
5 13 1 15 9 2
5 13 1 15 9 2
7 15 13 13 9 9 0 2
7 10 9 13 13 1 9 2
6 12 13 9 0 3 2
25 15 13 9 1 10 9 1 9 0 2 3 0 9 10 9 1 15 15 13 1 10 9 10 0 2
26 10 9 13 1 2 12 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 2
14 13 3 12 12 9 1 9 10 9 2 1 9 0 2
5 3 3 13 9 2
19 10 9 13 14 10 9 10 3 2 0 1 10 9 1 10 9 10 0 2
13 13 13 1 9 1 10 9 16 13 1 9 0 2
13 13 9 7 13 9 0 0 1 10 9 10 0 2
6 10 9 1 11 0 2
12 7 13 9 1 10 9 1 10 9 1 11 2
6 13 1 15 9 9 2
18 13 9 16 13 1 15 9 9 7 13 9 1 9 1 9 10 9 2
15 3 2 4 13 1 9 9 16 13 3 7 3 13 3 2
9 1 10 9 10 0 3 13 3 2
12 8 8 8 0 2 3 1 10 9 10 0 2
22 10 9 0 7 13 9 9 2 7 1 10 15 13 9 1 10 9 10 3 2 0 2
12 11 2 2 15 3 13 16 13 1 15 9 2
17 10 9 4 13 16 15 13 1 3 2 9 2 1 3 2 9 2
8 7 13 1 9 15 13 2 2
29 9 9 15 13 1 10 9 1 9 2 1 9 2 1 9 2 1 9 2 1 9 2 1 9 7 3 1 9 2
46 1 13 9 2 15 13 1 9 1 9 0 1 11 2 2 7 13 1 9 1 11 16 1 15 12 12 9 1 2 12 10 9 16 15 13 13 1 2 12 9 7 15 1 2 12 2
4 15 9 0 2
8 9 0 4 13 1 11 2 2
6 7 10 9 13 13 2
6 13 1 9 3 0 2
8 11 13 16 2 15 3 13 2
6 13 16 13 1 11 2
12 7 3 2 4 13 1 11 7 1 9 11 2
17 3 3 1 9 11 16 13 1 15 12 9 1 9 1 9 2 2
10 10 9 1 9 0 1 15 4 13 2
4 9 2 7 2
42 15 13 14 10 9 10 0 16 13 1 11 2 1 10 9 3 13 1 9 10 9 2 7 1 15 10 9 10 3 2 13 1 10 9 10 12 1 10 9 10 0 2
15 2 3 2 4 13 10 10 9 7 13 13 9 13 2 2
26 1 11 13 1 11 14 10 9 10 0 1 9 1 9 9 2 1 16 13 12 9 1 2 12 0 2
12 15 13 1 2 12 9 14 11 11 1 11 2
12 1 10 9 13 11 12 9 1 11 12 9 2
6 10 9 13 1 11 2
28 8 1 9 9 13 1 9 9 16 13 1 9 10 9 1 9 9 2 1 16 13 12 9 1 2 12 9 2
10 15 13 14 11 11 1 11 1 9 2
11 8 13 3 1 9 9 10 9 1 11 2
9 10 12 2 11 11 7 11 11 2
8 15 13 1 9 1 12 9 2
17 8 1 9 2 11 11 12 12 2 11 9 9 9 0 12 12 2
8 10 9 11 11 11 12 12 2
27 8 13 1 11 1 10 9 10 12 1 9 11 1 11 2 16 13 1 10 9 14 11 11 12 2 12 2
18 1 9 10 9 13 11 14 11 11 12 12 2 12 12 2 12 12 2
12 11 13 14 11 1 11 12 12 2 12 12 2
19 1 10 9 1 9 13 11 7 11 11 14 11 7 11 11 12 2 12 2
38 8 9 1 11 13 1 11 9 0 1 2 12 9 1 10 9 10 0 1 9 9 1 16 13 12 9 2 10 9 10 0 2 11 11 12 9 2 2
13 11 13 14 11 11 1 9 9 1 2 12 9 2
17 8 1 9 13 1 9 11 1 9 11 11 16 13 1 9 11 2
33 10 9 13 1 9 11 12 9 1 2 12 9 2 1 13 1 2 12 9 14 11 11 1 9 9 16 13 1 10 9 16 13 2
29 11 2 11 11 2 11 2 11 2 9 2 11 2 11 2 9 2 2 11 2 11 2 9 2 2 11 2 11 2
6 10 9 2 11 11 2
30 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 2 9 2 11 11 2 11 2 11 2 11 2 11 2 2
7 10 9 2 11 11 11 2
10 13 11 11 2 12 9 2 1 11 2
37 3 2 11 9 9 13 14 9 12 12 2 7 13 14 10 9 1 0 16 13 1 9 11 1 10 9 1 11 2 15 3 13 14 3 16 13 2
8 9 15 7 13 1 9 9 2
40 15 3 13 2 1 9 11 7 9 15 2 16 3 10 9 13 1 11 11 2 1 9 9 9 7 9 15 16 13 9 1 10 9 1 9 15 13 10 9 2
20 10 9 13 1 9 14 9 10 9 16 1 15 13 11 1 9 15 10 0 2
78 9 11 2 11 2 11 2 11 7 11 16 13 14 11 10 0 2 13 9 0 1 9 10 9 7 1 9 14 11 1 10 9 10 12 13 1 9 2 12 2 2 11 13 1 9 13 1 10 9 10 0 2 13 9 1 9 10 9 7 11 13 1 3 16 13 3 7 1 10 9 1 2 12 9 13 12 12 2
44 9 1 10 9 16 13 13 10 9 1 12 9 2 9 12 1 9 15 2 14 10 13 10 0 13 11 11 16 13 1 9 1 11 11 7 13 14 9 15 10 0 14 11 2
11 1 10 9 10 2 12 12 12 1 11 2
23 11 11 13 9 0 1 9 16 13 1 9 11 7 3 13 13 3 1 9 15 14 11 2
63 9 15 14 11 10 0 1 10 9 10 12 7 1 10 9 10 12 9 15 10 0 14 11 11 1 11 13 1 9 1 9 10 9 2 16 9 11 13 13 1 9 11 7 13 1 10 9 10 2 12 1 9 12 14 11 9 1 9 11 1 10 9 2
29 10 9 13 1 13 1 9 15 2 3 11 13 1 9 10 9 7 11 11 7 11 1 9 0 13 1 9 11 2
3 11 2 2
31 3 16 13 13 14 11 11 7 14 11 11 2 13 4 13 1 10 9 10 15 1 11 1 11 2 16 13 9 1 3 2
22 11 13 1 3 1 9 0 1 12 9 7 13 1 12 12 1 10 11 10 3 13 2
21 11 13 3 3 14 9 10 2 12 2 12 9 2 7 13 10 9 14 10 11 2
19 11 11 2 12 9 2 7 11 11 2 12 9 2 3 13 14 10 0 2
39 10 9 10 0 16 3 13 1 3 13 11 2 16 13 1 10 9 11 3 16 3 13 13 1 15 1 9 10 11 2 11 3 13 1 9 15 12 12 2
28 10 9 11 11 1 12 9 7 2 12 9 7 10 9 11 2 16 13 12 9 2 13 0 1 9 10 9 2
27 9 11 16 13 12 9 13 14 9 1 9 0 1 11 11 2 12 12 2 10 9 10 0 14 10 11 2
10 11 13 9 0 1 11 11 12 12 2
9 11 11 11 13 1 11 12 12 2
11 11 11 13 13 2 3 14 11 12 12 2
8 11 13 12 9 1 10 9 2
26 11 13 14 11 12 12 2 11 13 1 11 12 12 2 11 1 11 12 12 7 11 1 11 12 12 2
34 9 10 9 16 13 9 1 9 11 2 11 11 11 11 12 12 2 11 11 11 11 12 12 2 11 11 12 12 2 11 11 12 12 2
29 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 2 11 2 11 2 11 2 2
6 10 9 2 11 11 2
29 11 2 11 2 11 2 11 2 11 2 11 11 2 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 2
6 10 9 2 11 11 2
11 13 11 11 2 12 9 2 1 9 12 2
28 11 11 13 3 9 1 10 9 10 0 2 1 16 9 12 13 14 15 1 9 10 9 2 14 13 12 12 2
22 10 9 10 0 14 9 12 13 16 15 13 9 7 13 9 2 16 16 10 9 13 2
18 10 9 16 13 14 12 10 9 11 7 11 2 13 14 9 10 9 2
25 1 10 9 13 9 9 9 9 2 11 11 2 16 13 9 1 9 15 7 13 13 13 9 9 2
4 9 3 13 2
28 9 15 14 11 11 16 13 1 10 9 1 9 2 13 14 10 9 7 15 10 9 10 12 16 15 13 9 2
16 11 11 13 13 1 9 9 15 14 9 15 1 9 10 9 2
26 9 15 0 2 3 0 2 4 1 9 1 9 7 13 1 13 16 13 1 9 3 1 10 10 9 2
11 10 9 13 0 7 4 13 14 10 9 2
38 9 12 13 3 1 10 9 10 0 2 7 1 10 9 10 12 13 9 13 1 11 13 9 2 16 11 13 1 0 7 11 13 7 13 1 9 15 2
12 10 9 10 0 13 1 10 9 10 2 12 2
48 11 11 13 9 1 9 11 2 11 13 1 11 16 13 1 10 9 10 0 14 9 10 2 12 7 11 13 14 10 9 2 13 14 10 9 7 3 3 13 9 0 1 9 10 9 10 0 2
12 12 9 1 1 3 13 11 9 1 9 15 2
35 11 13 9 1 11 16 13 15 1 9 10 12 2 1 10 9 13 13 11 7 11 2 7 11 13 7 11 13 14 10 9 1 9 11 2
13 11 11 13 13 14 10 9 7 13 14 15 3 2
25 1 10 9 10 2 12 13 11 1 1 9 10 9 2 11 13 7 13 14 10 9 1 10 9 2
10 11 2 9 2 9 10 9 2 2 2
23 11 11 13 2 16 4 13 1 9 1 10 9 16 15 13 0 1 12 9 1 12 9 2
19 1 9 10 9 16 13 3 1 11 13 11 11 14 10 9 11 12 12 2
8 14 12 10 9 13 11 11 2
16 11 11 13 9 2 12 1 11 2 9 12 1 12 9 2 2
21 10 9 1 10 9 2 11 2 12 9 2 2 13 12 12 1 9 9 14 9 2
4 11 10 0 2
13 9 0 2 11 12 11 12 2 11 12 11 12 2
25 11 1 9 11 1 9 10 9 14 15 3 1 10 9 10 0 1 11 13 9 10 9 11 11 2
16 2 11 13 16 15 4 1 9 14 9 1 13 1 9 2 2
7 11 13 12 1 12 9 2
53 9 15 14 11 13 1 9 14 9 10 9 13 14 10 9 10 0 10 0 2 16 3 13 13 1 11 1 10 9 1 11 1 11 2 7 3 13 1 9 9 0 7 3 13 9 9 15 1 9 2 12 9 2
20 11 2 12 9 2 13 1 10 9 7 13 1 10 13 1 9 15 14 11 2
26 1 12 16 13 1 15 1 12 9 2 11 7 11 2 9 9 2 11 13 1 11 7 11 1 11 2
22 10 9 10 9 10 12 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2
14 12 9 2 9 0 1 11 2 13 3 1 9 9 2
16 11 11 13 1 9 11 1 9 0 11 1 16 13 12 9 2
16 1 9 10 9 1 9 12 13 11 11 2 16 13 12 9 2
21 13 10 9 11 1 11 13 1 9 10 9 1 10 9 10 0 2 1 9 11 2
14 1 9 11 13 10 11 11 1 9 11 1 12 9 2
6 10 9 13 1 11 2
43 11 11 1 11 2 7 10 9 11 2 13 9 9 1 9 11 1 9 1 10 9 10 0 2 1 13 1 11 11 16 13 14 10 9 1 9 9 1 9 11 10 0 2
22 9 10 9 13 1 9 11 1 9 1 9 11 2 1 9 10 9 1 9 9 11 2
27 1 9 11 13 12 9 2 1 9 11 9 12 7 1 1 10 9 10 0 12 9 2 9 1 9 11 2
22 2 9 10 9 14 9 11 2 4 13 1 9 9 15 1 9 11 2 13 1 11 2
11 11 13 1 9 1 9 9 15 10 0 2
21 1 9 0 16 13 1 15 1 11 13 2 16 15 4 13 1 13 14 10 9 2
19 3 13 10 9 11 1 10 9 7 3 15 13 1 9 0 14 9 11 2
35 9 10 9 2 16 13 13 1 9 1 10 9 1 10 9 11 1 9 11 1 11 2 13 1 9 1 9 10 9 1 1 9 10 9 2
32 11 13 1 10 9 1 10 9 11 11 2 16 13 1 10 9 2 13 1 9 10 9 2 7 13 1 11 13 14 10 9 2
24 10 9 13 1 10 9 3 1 2 12 1 10 9 2 1 16 13 1 9 9 1 10 9 2
9 1 9 9 10 9 13 10 9 2
14 1 9 15 11 3 3 13 1 9 10 9 11 11 2
18 9 10 9 14 10 9 11 11 13 16 11 13 7 13 1 10 9 2
16 11 16 13 1 9 1 10 9 13 13 7 13 13 12 9 2
8 15 13 14 14 11 1 9 2
10 9 10 9 13 9 1 9 10 9 2
20 3 1 10 13 16 11 13 3 1 9 10 11 1 9 10 9 14 9 15 2
41 10 9 10 0 1 9 13 3 1 9 10 9 10 2 12 1 9 14 9 2 1 9 10 9 1 9 1 11 2 9 10 9 7 11 1 9 11 1 10 9 2
42 12 10 9 16 13 1 9 16 13 7 15 16 13 3 4 13 9 1 9 15 14 10 9 2 9 15 7 9 10 9 1 15 2 7 3 4 13 9 7 3 9 2
25 2 13 1 9 1 10 15 12 9 2 2 13 1 15 1 9 10 9 9 11 9 9 11 9 2
56 10 9 13 3 1 13 1 9 9 15 2 7 1 9 16 9 0 13 7 16 1 11 9 9 3 13 4 1 1 10 9 13 13 1 10 9 10 0 1 9 10 9 10 0 2 16 13 1 15 9 1 10 11 2 11 2
22 1 11 9 9 13 3 3 9 16 3 13 14 10 9 1 15 1 10 9 9 15 2
21 1 10 9 10 0 11 11 2 1 15 11 11 7 11 11 2 7 1 11 11 2
49 9 13 1 15 3 14 10 9 16 11 11 2 9 9 13 1 10 15 2 13 1 10 9 10 0 7 16 11 13 1 9 0 2 1 11 2 16 4 13 7 13 7 13 0 3 3 1 15 2
36 2 15 16 11 3 13 1 12 9 2 4 1 15 13 14 10 9 16 10 9 11 13 10 0 1 10 9 7 9 15 13 2 2 13 9 2
23 2 1 11 1 11 2 16 3 1 15 9 0 2 4 13 1 9 1 1 9 10 9 2
9 3 13 4 1 11 9 9 3 2
19 9 10 9 13 1 9 15 9 7 3 9 3 13 2 1 1 10 9 2
42 3 16 13 1 10 9 1 3 13 11 11 2 9 10 9 11 2 16 1 10 9 10 12 14 15 1 10 9 3 2 1 15 13 14 10 9 11 11 13 9 13 2
34 3 11 13 3 1 12 9 9 1 12 2 7 13 1 15 14 11 9 9 2 12 12 2 7 14 10 9 9 9 2 12 12 2 2
45 9 0 16 4 1 9 2 13 16 10 9 11 13 3 1 9 16 13 7 3 2 13 2 1 15 7 1 10 15 13 13 9 2 9 1 10 9 1 10 9 1 11 9 9 2
19 2 3 16 13 1 9 15 14 9 15 10 11 2 11 2 2 13 11 2
27 2 0 16 3 9 16 13 1 10 9 2 9 13 1 15 9 12 9 2 7 15 3 13 1 10 9 2
23 11 9 9 13 1 10 9 1 1 9 0 2 7 3 10 9 10 0 13 1 10 9 2
17 10 9 14 15 13 13 1 10 9 10 0 2 1 10 9 9 2
30 15 13 16 13 9 0 1 16 3 2 7 3 13 1 9 10 9 7 13 1 9 12 9 1 11 2 13 0 2 2
47 3 1 9 9 10 9 10 0 11 11 2 16 15 9 12 14 15 2 12 1 11 7 2 12 1 11 2 9 0 2 2 1 12 10 9 10 0 13 10 9 1 11 1 9 15 2 2
13 1 15 13 11 2 2 11 4 13 14 10 9 2
7 15 13 16 15 3 13 2
8 15 4 13 3 3 1 11 2
8 10 9 13 1 10 9 2 2
6 3 11 1 11 13 2
31 13 11 2 2 3 1 10 9 16 13 13 9 10 9 1 10 9 10 0 2 7 15 13 3 13 1 9 15 14 9 2
11 15 3 13 16 11 13 1 12 10 9 2
10 1 9 15 3 9 12 13 1 9 2
12 3 13 9 12 2 7 3 13 1 10 9 2
37 7 13 1 12 1 12 10 9 10 0 1 10 9 9 9 2 11 9 9 7 10 9 9 0 15 13 9 0 2 16 13 1 15 9 3 2 2
26 11 13 16 10 9 3 13 14 9 15 2 16 16 9 13 2 1 9 15 10 13 14 10 9 15 2
24 1 10 9 13 9 0 2 10 9 11 2 11 9 9 7 11 9 10 11 13 1 10 9 2
6 1 10 12 13 12 2
6 1 10 12 9 0 2
32 8 8 10 9 10 0 1 10 9 7 1 10 9 2 10 9 1 10 9 11 11 13 1 11 1 10 9 11 2 12 2 2
18 9 0 1 9 9 9 1 9 10 9 10 13 14 11 2 12 2 2
18 10 9 10 9 11 13 1 10 0 1 10 9 2 1 9 10 11 2
9 9 0 13 9 0 2 12 2 2
17 11 9 9 13 1 11 7 13 1 3 1 9 0 2 12 2 2
37 10 9 9 0 13 13 1 9 11 14 9 9 15 1 11 2 3 1 11 9 9 2 16 13 12 9 9 0 1 10 9 10 0 2 12 2 2
19 10 9 11 4 13 14 9 15 1 13 1 9 1 11 11 2 12 2 2
34 1 10 9 1 10 9 9 13 12 12 1 9 0 1 9 15 14 11 11 2 13 9 10 9 1 11 13 1 11 1 9 10 9 2
9 11 13 12 12 3 1 12 9 2
18 3 13 15 11 9 16 13 1 10 9 10 2 12 9 14 11 11 2
18 1 10 9 10 2 12 13 1 10 9 9 11 11 11 14 11 11 2
20 11 11 2 10 9 10 0 16 4 13 3 1 11 2 13 1 2 12 9 2
20 9 13 9 12 1 10 9 2 12 14 15 3 2 1 10 9 10 2 12 2
18 8 8 13 11 11 14 10 9 10 12 2 3 15 1 9 14 11 2
33 10 9 1 10 9 2 11 2 13 3 1 12 10 9 10 0 1 13 12 7 13 1 12 9 1 9 12 1 9 0 1 11 2
24 11 11 13 12 12 1 11 1 10 9 10 2 12 7 11 11 13 1 10 9 10 2 12 2
17 1 10 9 10 2 12 13 11 1 9 12 1 9 14 11 11 2
17 9 11 2 10 9 11 11 2 13 13 1 10 9 1 2 12 2
8 3 13 12 10 9 10 0 2
24 3 9 14 11 11 1 10 9 10 2 12 7 1 15 14 11 11 1 10 9 10 2 12 2
9 11 13 12 12 14 11 9 11 2
24 10 9 1 11 2 11 11 2 12 2 2 11 11 11 2 12 2 2 11 11 2 12 2 2
9 11 2 9 11 2 12 12 2 2
8 1 9 0 4 13 13 9 2
54 1 10 9 1 9 1 11 11 2 13 3 12 9 1 9 2 9 2 9 12 2 11 11 2 11 11 2 7 9 10 9 1 11 11 1 11 1 10 9 10 0 2 0 11 11 16 13 14 10 9 1 9 9 2
61 11 9 2 16 13 1 10 9 16 13 1 9 11 1 11 11 2 13 3 9 0 1 10 9 1 9 1 9 10 9 10 0 11 11 1 10 9 10 2 12 2 7 13 1 2 12 12 1 9 15 1 11 16 13 1 10 9 10 2 12 2
16 1 10 9 10 2 12 13 11 11 9 2 12 1 11 9 2
23 9 11 2 9 11 2 13 9 0 3 1 10 9 10 2 12 1 9 1 2 12 9 2
39 9 10 9 14 11 13 1 9 2 12 14 11 11 2 16 3 1 10 15 13 14 10 9 16 13 1 9 1 10 9 1 9 15 14 9 11 11 11 2
27 8 8 13 0 1 10 9 10 12 1 12 9 1 9 12 12 1 11 2 16 13 0 1 12 9 3 2
21 10 9 1 10 9 2 11 2 12 9 2 2 13 12 12 1 10 9 1 11 2
19 10 9 13 1 2 12 9 1 9 9 9 16 13 1 9 1 10 9 2
18 13 16 12 9 13 1 9 10 13 7 2 12 0 13 1 9 0 2
15 1 10 9 10 0 13 9 9 7 13 9 1 10 9 2
64 9 0 1 10 9 10 12 2 11 12 11 12 2 11 12 11 11 12 2 11 12 11 12 2 9 11 12 11 11 12 2 11 12 11 12 2 11 12 11 12 2 11 11 12 9 11 12 2 11 12 9 9 12 2 11 12 11 12 2 11 12 11 12 2
37 15 13 1 13 14 10 9 1 10 9 1 9 10 9 2 1 15 13 1 9 11 10 0 2 12 1 11 2 10 9 10 0 14 11 7 11 2
30 15 13 9 10 9 14 11 1 10 9 10 3 0 2 7 7 1 11 13 15 9 12 1 10 9 1 11 12 12 2
7 1 9 15 13 3 11 2
31 11 13 3 16 1 10 9 2 16 13 3 2 12 12 9 2 9 0 9 12 12 9 16 13 9 1 10 9 10 0 2
11 10 9 9 15 13 3 2 12 12 9 2
20 1 16 10 9 0 2 9 10 9 13 7 10 13 13 1 3 2 12 9 2
17 10 9 10 0 13 1 9 1 9 0 2 16 13 1 12 9 2
20 11 13 16 13 14 10 9 1 9 10 9 11 11 7 10 0 13 9 9 2
15 10 9 10 0 13 3 14 10 9 1 10 9 1 11 2
22 1 10 9 3 13 9 0 7 13 1 15 12 9 11 11 2 11 11 7 11 11 2
31 3 13 9 9 1 10 9 11 1 10 9 10 0 7 1 9 11 9 9 0 1 10 9 9 9 1 10 9 10 0 2
19 3 9 12 13 12 10 9 10 0 13 9 1 9 9 10 9 10 0 2
55 1 9 9 13 15 9 9 2 1 10 9 10 12 14 10 9 2 1 16 13 7 13 9 1 13 14 10 9 1 9 11 11 2 16 13 1 9 9 7 9 2 7 1 9 2 1 10 9 10 0 3 1 9 15 2
39 1 9 3 13 10 9 9 12 10 0 16 3 3 13 2 7 14 10 9 13 12 10 9 10 0 16 3 3 13 9 2 11 9 2 11 2 11 2 2
18 7 16 12 10 11 13 2 11 11 14 11 9 3 13 14 10 9 2
61 1 12 9 1 15 3 13 13 7 13 9 3 1 2 12 2 13 3 11 11 1 9 15 12 12 14 10 9 1 15 1 10 9 2 10 9 9 11 2 1 13 1 9 10 9 1 12 9 7 9 0 3 1 9 10 9 2 12 12 2 2
30 1 9 11 13 3 12 9 9 10 0 1 15 2 16 13 7 13 1 10 9 13 14 10 9 10 15 1 9 15 2
47 1 10 9 10 12 13 11 11 2 16 13 1 10 9 7 13 1 9 15 1 9 12 13 14 9 15 10 0 3 2 12 12 2 2 1 9 0 0 14 12 9 1 10 15 1 15 2
37 11 11 13 1 10 9 10 12 1 16 13 9 0 1 10 9 9 9 2 16 13 15 9 10 9 14 15 2 12 12 2 1 9 14 11 11 2
50 11 9 9 13 14 9 15 10 12 2 3 1 9 1 11 2 3 12 7 13 1 13 14 10 9 7 13 14 10 9 16 1 12 10 9 10 0 13 10 9 10 0 16 10 9 3 13 1 15 2
48 10 9 11 13 14 11 11 12 1 12 10 9 10 0 16 3 3 13 9 2 16 13 1 10 9 12 12 7 13 14 15 1 9 2 1 9 1 12 9 10 9 1 11 7 1 9 9 2
32 10 9 10 0 1 9 9 13 1 10 9 14 10 9 7 10 9 13 13 1 9 9 2 16 13 14 9 15 1 10 9 2
27 3 13 9 15 14 10 9 1 9 10 9 2 16 1 11 11 13 14 10 9 10 9 0 1 12 9 2
23 14 10 10 12 13 9 15 10 0 2 9 9 0 0 7 0 2 7 3 9 9 0 2
36 1 10 9 10 2 12 13 12 9 2 13 12 9 7 13 2 1 9 9 9 2 9 10 9 2 12 12 9 2 9 14 12 9 1 9 2
43 1 10 9 16 10 9 13 1 9 13 2 7 13 16 3 16 13 3 15 2 3 2 3 2 16 13 2 13 1 15 10 9 2 16 3 15 0 16 3 13 0 3 2
42 9 0 15 2 16 9 15 3 3 1 9 2 9 7 1 9 9 7 9 2 13 1 15 1 10 9 16 9 0 2 9 7 9 2 13 1 9 9 1 9 9 2
20 1 16 13 1 9 15 2 1 9 0 3 2 1 10 9 10 0 14 15 2
79 1 10 9 1 11 7 1 11 2 13 1 10 9 16 13 1 11 9 0 1 10 9 2 1 13 1 9 14 10 9 10 0 7 13 14 10 9 10 0 1 10 9 10 0 2 10 9 10 3 0 10 0 14 15 1 9 11 14 10 9 10 0 1 11 2 1 9 12 1 11 2 16 13 3 14 11 7 11 2
26 9 15 13 9 1 10 9 1 11 2 7 16 3 13 14 10 9 10 0 7 13 3 9 9 0 2
53 10 9 10 0 3 13 2 7 10 9 11 11 7 11 11 13 14 10 9 1 9 10 9 10 0 10 0 2 1 9 10 9 7 1 9 10 9 2 3 3 7 13 1 9 0 2 7 13 1 9 0 3 2
36 1 9 15 2 13 10 9 1 12 9 0 2 3 10 9 10 0 10 0 2 1 1 9 12 2 4 13 3 1 16 16 13 1 9 15 2
25 7 3 9 10 9 10 15 2 16 16 15 13 7 13 10 9 10 9 2 3 0 1 9 15 2
60 3 7 4 3 13 1 9 0 1 9 2 1 9 9 0 14 0 1 9 0 3 9 0 9 2 16 0 3 1 10 9 9 0 2 7 3 2 16 4 13 15 1 9 12 1 11 2 11 2 11 2 11 2 11 2 11 7 11 11 2
13 13 11 2 11 11 7 11 2 7 13 9 0 2
13 3 16 13 0 1 9 2 9 2 10 9 13 2
13 9 2 10 9 13 3 9 1 9 2 9 0 2
9 10 9 10 0 3 13 1 15 2
36 9 15 14 11 2 11 2 11 2 11 2 11 2 11 11 7 0 13 1 9 0 2 7 3 16 13 14 15 1 9 12 12 13 3 13 2
25 3 3 13 9 15 1 9 1 9 12 12 2 7 9 15 1 10 9 13 1 3 7 13 9 2
6 3 3 1 10 9 2
33 15 13 1 9 0 2 1 9 0 2 14 1 10 9 16 1 9 15 9 0 3 7 1 10 9 10 0 1 9 10 9 3 2
22 1 10 10 9 2 3 9 15 10 0 4 13 1 15 1 10 9 2 1 10 9 2
41 7 3 10 13 7 10 9 16 1 15 2 7 13 3 14 9 2 11 11 2 11 2 11 2 11 9 10 9 14 15 7 13 1 15 7 13 3 10 1 15 2
21 10 9 14 15 13 14 9 10 9 14 9 9 15 0 2 3 3 1 9 15 2
34 13 10 9 0 13 3 1 9 9 0 0 2 13 7 0 2 16 3 13 1 10 9 16 13 7 13 1 15 14 9 2 10 9 2
26 10 9 1 12 9 2 14 1 11 12 13 14 9 10 9 10 0 3 1 9 0 2 13 1 9 2
28 9 10 9 2 1 12 2 2 16 13 1 9 12 1 11 2 13 1 15 3 9 0 7 3 9 3 0 2
36 4 13 2 16 9 0 13 10 9 10 2 0 2 14 9 11 1 9 0 2 16 13 3 1 9 0 14 10 9 10 0 1 10 9 15 2
21 15 10 9 1 10 9 10 0 14 11 2 11 2 11 7 9 0 1 10 9 2
17 3 9 0 2 3 2 14 1 9 10 9 9 12 1 9 9 2
37 7 13 16 1 9 15 2 1 9 2 9 2 9 7 9 2 13 10 9 13 1 9 9 1 9 1 11 2 16 10 3 13 13 1 15 3 2
71 3 3 16 16 15 0 3 1 9 9 2 9 7 9 2 3 3 1 16 0 1 15 9 1 9 0 2 9 7 9 2 7 3 3 16 16 9 13 2 16 10 9 10 0 16 15 13 0 1 10 9 7 13 13 1 9 12 1 10 9 7 10 9 2 10 9 7 9 10 9 2
22 3 16 13 1 9 0 1 12 9 2 3 3 1 15 3 7 3 1 9 0 0 2
71 14 10 9 4 13 1 10 9 2 1 9 10 9 2 1 9 10 9 2 1 10 9 10 0 2 1 10 9 2 1 10 9 7 3 1 9 10 9 7 1 10 9 16 13 14 15 2 1 10 9 1 9 0 7 0 16 13 1 9 0 1 10 1 9 15 10 0 14 9 0 2
20 10 9 10 0 3 13 2 13 9 2 2 7 3 13 1 10 9 10 0 2
37 13 1 15 9 9 1 14 15 3 1 10 9 7 13 3 9 7 9 7 15 13 9 9 0 2 9 9 1 9 2 9 2 9 9 7 9 2
20 9 10 9 10 0 13 1 10 9 2 3 10 9 14 15 13 1 16 13 2
14 10 3 9 2 9 7 9 2 3 3 9 7 9 2
91 1 9 9 10 0 2 1 3 13 9 2 14 1 10 9 13 9 2 14 1 11 13 13 2 1 3 13 9 2 9 7 9 2 9 2 14 9 13 1 9 7 1 9 1 1 9 7 1 9 13 9 0 1 9 9 1 9 7 13 3 2 13 2 1 10 9 1 9 10 9 16 1 9 10 9 2 7 1 9 10 9 10 0 16 1 10 9 1 9 11 2
23 3 13 1 9 10 9 9 0 7 9 9 2 7 13 9 0 7 3 2 12 1 9 2
14 7 7 13 3 15 2 3 2 13 14 10 10 9 2
28 11 7 9 11 2 16 13 1 9 1 9 15 1 9 1 12 9 0 1 11 11 3 13 1 13 1 11 2
30 3 13 9 11 11 13 1 9 15 14 10 9 10 0 2 3 1 9 0 2 3 1 3 13 1 10 9 11 11 2
4 11 2 11 2
11 11 2 11 2 2 11 2 11 2 11 2
18 11 2 11 2 11 11 2 11 2 11 2 11 2 2 11 2 11 2
6 10 9 2 11 11 2
4 11 2 16 2
11 11 2 11 2 11 2 2 11 2 11 2
20 11 2 11 11 2 11 2 2 11 11 2 11 2 11 2 11 11 2 11 2
6 10 9 2 11 11 2
11 13 11 11 11 2 12 9 2 1 11 2
20 1 9 13 10 9 10 9 0 10 0 1 10 9 1 11 12 12 9 0 2
49 3 13 1 10 9 10 9 0 10 0 2 1 10 9 1 11 2 3 1 2 12 9 7 3 15 13 1 9 10 9 10 0 2 1 1 9 10 9 16 13 3 0 1 9 10 9 10 0 2
17 1 11 15 13 9 9 0 16 1 9 15 13 1 9 10 9 2
39 10 9 13 9 1 9 9 0 7 0 16 13 3 14 9 11 7 13 1 9 10 9 14 15 2 7 3 13 3 1 10 9 10 0 2 9 0 2 2
23 10 10 9 13 1 12 9 10 2 12 2 14 3 3 13 10 9 13 1 9 10 9 2
19 3 13 9 1 10 9 7 9 10 9 13 7 7 3 1 9 1 0 2
12 9 9 15 13 1 9 0 7 1 9 9 2
41 1 9 10 9 10 0 7 9 10 9 10 0 2 13 10 9 3 14 1 10 9 13 10 9 1 10 9 2 3 1 16 10 9 13 1 10 9 0 10 9 2
6 11 13 1 9 15 2
11 11 11 13 3 7 11 11 13 0 3 2
12 3 10 10 9 3 13 1 9 15 10 0 2
37 3 1 10 9 10 2 12 13 10 9 3 1 10 9 2 7 13 15 11 11 16 13 1 2 12 9 7 11 11 13 1 9 0 1 10 9 2
32 1 10 9 10 2 12 13 11 11 2 1 10 9 10 0 14 15 2 1 9 1 2 12 9 7 10 9 13 1 10 9 2
42 7 1 10 9 10 2 12 2 1 10 9 10 0 16 13 1 10 9 10 12 1 10 9 2 13 11 3 7 15 13 9 0 1 2 12 9 1 1 9 10 9 2
51 3 1 9 9 0 15 13 10 9 7 13 10 9 1 10 9 2 7 13 15 9 15 14 10 9 16 13 13 2 9 12 1 9 2 1 9 0 2 7 3 1 9 15 10 12 7 13 1 9 0 2
34 9 2 7 16 13 10 9 1 10 9 10 0 1 11 2 13 9 1 10 9 10 0 14 10 9 10 0 1 15 13 9 3 13 2
16 3 13 10 12 1 10 9 16 3 13 9 2 12 12 2 2
17 10 9 11 13 14 10 9 16 13 1 15 1 9 0 1 9 2
12 3 10 9 10 0 14 10 9 4 1 9 2
41 3 1 9 10 9 10 0 10 0 13 9 0 1 10 0 2 10 9 11 2 16 13 12 12 14 11 11 7 1 15 12 9 3 1 11 16 13 14 10 9 2
17 1 10 9 10 12 13 11 11 16 13 14 10 9 11 12 12 2
19 11 11 13 13 9 3 12 12 1 11 11 7 13 1 10 9 10 12 2
19 11 11 13 12 12 14 11 11 7 13 1 10 9 10 12 1 10 12 2
17 10 9 11 13 1 9 9 12 12 1 16 13 12 12 1 11 2
10 3 11 7 11 13 1 9 12 12 2
12 9 9 7 9 10 9 13 1 9 12 12 2
25 12 9 2 16 13 1 10 9 1 11 13 1 9 0 1 9 0 1 10 9 15 1 10 9 2
19 10 9 13 1 10 9 10 0 14 10 9 7 10 9 10 0 14 11 2
7 13 9 2 9 7 9 2
13 9 10 9 13 1 9 7 13 9 0 7 0 2
9 1 9 10 9 10 0 13 9 2
10 13 11 11 2 12 9 2 1 11 2
22 11 11 11 1 9 10 9 3 13 13 9 15 1 13 1 11 11 1 9 10 9 2
42 10 9 16 13 1 9 0 13 1 9 15 1 9 1 10 9 10 0 2 7 10 0 2 16 13 14 10 9 10 12 1 9 2 13 13 7 13 13 1 9 0 2
24 10 9 10 0 1 9 15 13 14 11 11 11 9 1 10 9 2 1 13 3 1 10 9 2
13 13 11 11 2 11 2 12 9 2 1 9 11 2
19 11 8 8 1 9 9 12 0 13 10 9 11 1 9 10 9 3 3 2
20 1 10 9 10 2 12 13 11 11 14 11 1 9 1 9 1 2 12 9 2
28 1 10 9 10 2 12 13 14 9 15 10 2 12 3 2 1 10 9 10 0 2 1 9 11 1 10 9 2
22 12 9 3 3 13 11 14 11 1 10 9 7 11 11 13 14 10 9 1 9 12 2
14 11 11 13 9 9 15 1 9 12 9 1 10 9 2
10 13 11 11 2 12 9 2 1 11 2
19 11 8 8 9 1 9 0 14 11 2 1 9 0 14 11 16 13 9 2
32 1 9 11 2 16 13 13 2 13 11 11 9 12 3 2 1 13 1 9 15 9 14 12 9 1 9 16 13 4 1 15 2
10 13 11 11 2 12 9 2 1 11 2
21 11 8 8 0 0 3 7 1 10 9 9 1 9 10 9 16 13 1 12 9 2
11 10 9 13 9 9 1 11 1 10 9 2
24 16 13 13 2 16 10 9 11 13 13 9 13 13 9 14 9 1 9 11 11 7 11 11 2
16 1 12 9 13 10 9 12 9 16 13 3 0 1 9 15 2
10 13 11 11 2 12 9 2 1 11 2
8 11 8 8 0 7 0 9 2
39 9 10 9 13 0 3 1 9 16 13 1 1 10 9 10 0 14 11 11 2 10 9 10 0 7 10 0 14 9 9 2 1 15 13 15 9 12 3 2
11 13 11 11 2 12 9 2 1 11 11 2
25 11 3 10 0 16 13 12 12 1 9 10 9 10 0 13 9 1 16 13 1 10 9 10 9 2
21 1 10 9 10 12 13 11 14 9 15 7 10 9 16 13 13 3 9 14 9 2
10 9 1 10 9 13 13 14 10 9 2
11 13 11 11 11 2 12 9 2 1 11 2
10 11 1 12 9 0 3 13 1 11 2
14 9 15 14 11 11 1 11 11 13 1 9 10 9 2
9 15 13 12 9 7 13 12 12 2
10 13 11 11 2 12 9 2 1 11 2
45 10 9 10 0 1 9 2 11 9 9 2 13 3 1 10 9 10 12 1 9 11 1 10 9 2 1 16 13 1 11 2 11 2 14 11 12 12 2 12 2 12 2 12 2 2
12 10 13 2 11 11 2 11 11 7 11 11 2
28 11 2 16 13 3 1 10 9 10 0 1 9 9 12 12 2 13 1 10 9 10 12 1 9 11 10 0 2
29 1 10 9 1 9 13 9 13 10 9 9 9 2 1 16 13 1 10 9 12 12 1 10 9 10 0 11 11 2
22 10 9 10 0 1 12 10 9 2 16 13 3 15 1 11 2 13 10 9 12 12 2
38 9 11 1 9 2 9 10 9 9 11 2 13 12 12 2 12 2 12 2 12 2 1 10 9 10 0 1 9 11 1 10 9 1 11 11 1 11 2
10 9 10 9 13 3 15 3 1 11 2
30 13 10 9 9 11 13 9 9 10 9 10 0 2 1 16 13 3 1 10 9 1 9 11 12 12 1 9 11 11 2
18 3 1 10 9 10 0 16 13 1 11 13 10 9 10 0 12 12 2
18 1 10 9 10 12 1 9 13 10 9 1 9 10 9 7 1 9 2
12 10 9 1 10 9 1 9 9 2 9 13 2
20 9 0 13 1 9 10 9 2 9 9 13 1 9 9 1 9 7 9 9 2
22 3 16 13 16 10 9 16 13 1 10 9 13 1 10 9 13 2 7 3 13 9 2
18 3 9 10 9 13 1 1 15 1 9 10 9 7 7 13 1 9 2
23 3 3 3 15 13 9 7 9 2 1 15 9 16 1 15 15 13 1 13 9 0 0 2
21 3 15 16 9 16 1 15 13 9 0 2 9 9 13 3 3 0 14 10 9 2
21 9 9 3 0 4 13 9 0 2 14 15 13 1 10 9 7 3 1 9 9 2
16 3 9 13 1 9 9 7 1 9 9 1 10 9 13 9 2
10 3 13 9 1 9 3 7 1 9 2
36 1 10 9 10 0 2 1 12 7 1 12 1 11 13 9 14 10 9 10 0 1 9 0 1 9 9 2 1 9 12 7 9 1 10 9 2
29 1 9 14 9 0 3 2 1 10 9 10 0 7 10 0 14 9 0 2 13 13 16 3 13 13 9 7 9 2
2 3 2
22 7 10 9 1 9 10 9 1 15 9 2 9 11 2 2 13 1 9 9 9 3 2
36 9 2 9 9 11 13 9 1 15 1 9 1 9 11 2 1 13 9 0 2 2 1 9 0 1 9 1 3 10 9 16 13 1 10 9 2
22 10 9 10 0 1 10 9 3 13 1 9 10 9 10 0 7 13 14 15 1 0 2
15 7 2 10 9 10 0 1 10 9 13 9 9 10 9 2
22 1 9 15 1 10 9 1 9 13 10 9 1 10 9 16 10 9 13 9 1 9 2
16 1 10 9 3 13 1 15 16 3 13 9 3 7 1 9 2
21 1 9 10 3 0 3 2 7 0 3 14 15 13 1 15 2 13 1 15 3 2
29 1 10 9 13 3 3 9 1 9 0 16 13 1 9 10 9 2 7 15 13 3 1 10 9 1 9 10 9 2
9 1 0 1 15 15 13 1 9 2
9 9 1 9 0 13 1 10 9 2
21 14 15 13 1 9 16 13 1 9 1 9 0 2 10 9 1 15 7 0 3 2
26 7 10 9 10 0 2 3 13 14 15 1 10 9 10 12 7 15 4 13 3 7 3 3 7 3 2
20 1 9 9 13 9 0 13 14 10 9 1 9 9 2 7 3 13 16 13 2
35 1 1 9 13 11 1 10 9 10 0 14 9 2 16 2 1 3 4 13 9 7 13 1 15 1 10 9 2 2 7 2 1 9 9 2
22 10 9 2 16 13 3 2 13 14 10 10 9 1 9 9 0 16 13 1 10 9 2
16 14 13 1 9 15 14 10 9 2 13 16 10 9 13 0 2
24 3 9 12 3 13 1 10 9 1 9 15 2 7 1 10 0 3 13 1 10 9 10 0 2
17 1 9 15 13 10 9 3 3 2 7 9 3 13 13 9 9 2
19 1 9 0 14 15 2 13 9 9 16 10 13 13 3 2 1 9 9 2
18 1 9 15 13 10 13 1 9 2 9 1 9 9 2 9 1 9 2
18 1 9 1 10 9 13 9 14 9 3 1 2 9 9 1 9 0 2
14 1 9 11 7 1 9 0 10 9 13 12 9 3 2
23 7 16 1 11 13 1 9 0 3 9 16 1 12 9 2 7 1 9 0 1 9 9 2
8 1 9 10 9 13 9 3 2
26 1 9 0 2 1 15 2 13 1 9 10 9 9 0 7 7 3 7 1 9 16 0 1 12 9 2
20 13 9 16 9 0 15 2 1 9 9 2 9 3 0 2 13 1 10 9 2
15 9 10 9 1 9 10 9 3 13 2 9 7 9 2 2
38 7 3 2 16 9 10 9 13 9 2 10 16 13 1 9 9 9 1 9 10 9 1 10 0 1 10 9 2 9 9 2 10 9 2 13 1 15 2
39 9 10 9 13 1 11 11 9 1 9 7 9 2 7 15 13 1 9 9 2 2 14 13 13 14 10 9 10 15 1 9 0 2 7 13 1 15 9 2
14 15 1 15 9 2 13 1 10 9 1 11 1 12 2
49 13 9 9 12 2 7 1 16 13 3 0 13 1 10 9 7 10 10 9 2 10 9 1 10 9 10 0 7 10 9 10 0 16 15 13 13 14 15 1 12 1 15 2 13 1 15 1 3 2
28 10 9 14 10 9 13 1 15 9 0 13 1 9 2 16 3 15 3 3 9 7 3 9 1 10 9 2 2
27 9 10 9 2 15 13 14 15 2 13 9 0 0 7 0 2 16 13 1 10 9 14 9 15 13 9 2
35 9 10 9 13 1 15 9 0 2 13 9 1 9 2 7 9 15 13 2 2 7 3 15 3 13 13 1 9 7 9 16 3 3 13 2
14 13 2 9 2 9 7 9 2 13 2 13 2 13 2
23 15 13 9 9 7 9 2 13 1 9 9 7 9 2 9 9 1 10 9 9 7 9 2
17 4 13 16 15 10 9 10 0 16 13 1 10 9 10 15 2 2
15 3 3 3 4 11 13 1 9 7 9 16 3 3 13 2
13 2 13 1 10 9 2 1 15 9 9 1 9 2
20 13 1 15 16 9 10 9 10 15 0 3 1 10 9 16 1 15 13 15 2
35 15 13 9 16 7 9 2 1 15 2 3 10 9 16 13 3 13 9 2 9 2 16 3 13 9 1 9 3 1 10 9 16 15 9 2
5 15 3 3 0 2
12 2 9 0 0 14 15 13 10 9 10 0 2
26 15 3 13 14 15 2 7 3 4 13 16 15 13 16 15 0 2 16 13 1 10 9 3 3 3 2
15 9 1 9 15 15 10 9 16 13 1 12 11 2 11 2
20 1 9 16 13 1 15 15 13 2 15 3 9 2 7 3 4 13 14 15 2
12 15 13 16 10 15 3 3 0 1 9 15 2
40 13 1 15 16 7 13 14 10 9 14 9 1 9 15 1 9 1 10 9 14 9 0 2 13 16 9 15 14 10 9 1 9 10 9 13 3 3 0 2 2
18 14 10 9 15 13 11 13 1 10 9 7 1 10 9 1 10 9 2
20 11 2 10 9 10 0 2 13 1 11 2 9 0 2 1 9 3 3 0 2
29 1 9 15 13 9 0 1 10 9 1 9 7 9 2 13 11 1 9 7 13 14 9 10 9 16 13 9 0 2
25 10 12 13 1 9 0 1 9 2 7 1 16 13 10 9 2 13 7 13 10 9 1 10 12 2
17 11 2 9 9 0 2 13 0 7 0 2 9 9 7 9 13 2
20 15 3 4 13 1 11 16 10 9 13 1 15 1 2 9 1 10 9 2 2
20 10 9 10 0 13 1 15 2 9 2 2 9 0 7 15 13 13 1 11 2
36 11 0 2 0 9 2 0 2 7 4 13 10 9 1 13 14 9 15 2 3 7 10 9 13 1 9 1 10 13 14 15 2 1 15 11 2
25 1 10 9 13 3 9 9 1 9 9 7 1 9 16 13 1 9 15 9 0 1 9 10 9 2
12 11 13 14 15 3 1 11 7 3 1 11 2
21 2 1 11 13 3 14 9 10 9 2 16 13 7 15 3 13 14 15 1 15 2
24 13 1 15 9 1 9 2 7 1 15 15 13 13 2 13 7 13 1 12 9 1 9 12 2
18 11 2 1 10 0 14 15 2 13 9 1 10 9 14 11 1 13 2
18 1 9 15 15 13 3 9 0 14 15 2 3 15 13 1 10 9 2
29 3 15 13 14 9 15 1 10 9 2 10 9 7 10 9 14 10 0 2 7 10 9 10 15 13 3 13 2 2
7 14 10 9 13 11 11 2
23 13 1 15 11 11 2 11 11 2 11 2 11 11 2 11 11 2 11 11 7 11 11 2
22 10 9 13 1 9 10 9 2 7 11 13 16 9 10 9 13 2 10 10 9 2 2
36 15 13 16 1 10 9 10 0 16 13 1 10 9 2 13 1 9 10 9 7 10 9 14 9 0 2 1 16 13 14 9 15 1 9 13 2
51 9 0 1 16 13 11 11 1 11 2 1 10 9 10 12 1 9 15 2 13 10 9 1 9 15 14 9 10 9 10 12 1 10 9 2 9 11 2 2 16 14 15 15 13 1 9 15 1 10 9 2
18 9 12 10 9 10 0 13 3 2 7 1 1 9 13 3 12 9 2
13 10 9 13 13 1 9 10 9 1 9 9 11 2
16 1 1 9 13 11 1 2 9 10 9 13 9 0 1 9 2
13 3 10 9 1 15 13 1 13 9 10 9 3 2
23 11 13 16 9 15 1 9 10 9 3 13 0 3 2 7 4 13 16 3 15 10 9 2
9 1 11 13 9 0 1 9 9 2
35 1 10 9 13 12 9 2 2 10 9 13 14 14 15 2 2 10 0 2 12 2 7 2 13 14 10 9 2 2 10 9 2 12 2 2
43 16 16 11 13 3 2 3 1 9 0 1 2 11 2 7 3 1 9 15 1 9 15 14 11 11 1 9 11 2 13 1 15 13 12 1 12 9 10 9 1 9 0 2
18 15 13 1 9 15 2 11 2 13 9 15 1 9 10 9 10 0 2
26 10 9 7 9 15 13 1 15 9 14 10 9 2 14 10 12 13 7 13 1 9 15 14 10 9 2
12 10 9 13 14 9 15 14 9 0 0 3 2
45 10 9 2 11 11 2 9 9 1 9 0 2 10 9 2 11 11 2 9 2 10 9 2 11 11 2 9 2 9 7 10 9 2 11 11 2 13 14 9 15 1 9 10 13 2
12 10 9 13 1 10 9 7 1 9 10 9 2
32 11 13 1 10 9 16 15 13 0 1 10 9 10 0 14 10 9 2 7 10 9 3 13 1 9 15 7 1 9 9 15 2
27 11 13 1 15 16 10 9 16 13 1 10 9 10 0 1 3 3 13 1 9 0 1 2 9 10 9 2
12 1 9 15 2 3 16 15 3 13 9 15 2
20 1 9 10 9 7 9 10 9 2 15 13 2 3 13 10 9 13 9 0 2
26 2 9 1 11 9 16 13 3 13 3 9 0 14 10 9 10 0 2 15 12 10 9 16 13 3 2
18 13 3 3 12 9 16 15 0 3 2 7 7 10 9 13 13 2 2
25 11 13 1 9 0 2 2 9 14 9 3 13 3 9 10 9 14 9 9 1 11 2 7 2 2
23 11 13 16 1 9 10 9 3 13 9 1 9 15 2 16 13 1 9 0 2 11 2 2
13 10 9 10 0 13 1 10 9 7 1 10 9 2
10 15 13 16 15 13 9 0 7 0 2
11 1 10 9 15 13 1 9 14 9 13 2
48 11 2 11 11 2 11 11 2 11 11 7 11 11 2 7 1 9 15 9 14 9 0 2 1 9 9 1 12 9 2 13 1 10 9 16 13 14 10 9 2 10 9 10 0 10 0 2 2
23 10 9 13 1 9 9 11 1 9 7 1 9 7 1 9 10 11 10 0 2 9 9 2
9 1 9 15 13 1 3 12 9 2
20 9 7 1 15 9 2 9 9 7 9 10 9 13 9 16 13 1 10 9 2
31 2 10 9 13 13 9 0 14 10 9 10 0 1 10 9 1 15 13 10 9 2 2 13 11 11 2 1 9 10 9 2
15 10 9 13 13 1 10 9 2 7 9 9 1 9 0 2
16 2 1 9 9 0 2 15 13 3 9 0 2 2 13 11 2
20 1 10 9 1 10 9 13 10 9 1 12 1 9 1 9 10 9 16 13 2
15 1 10 9 13 1 10 9 10 0 1 12 1 12 9 2
6 3 3 13 12 9 2
46 10 9 13 1 9 1 10 9 1 10 9 2 1 9 1 9 10 9 2 1 9 0 7 3 2 2 7 15 3 9 10 9 2 13 9 2 7 16 9 13 1 9 1 15 2 2
20 9 0 2 7 9 1 9 2 13 1 9 9 0 7 13 1 9 9 9 2
10 10 9 13 1 9 11 1 10 12 2
37 2 2 1 2 9 9 14 11 11 2 13 11 11 14 2 15 13 1 15 1 9 1 9 2 2 10 9 16 13 1 9 15 10 0 14 11 2
26 10 9 13 1 10 9 1 9 15 7 15 13 1 15 1 9 13 7 1 9 11 11 14 11 11 2
44 15 9 15 14 9 2 11 11 2 2 9 9 9 2 16 13 14 9 15 2 11 2 11 11 2 2 7 4 2 7 3 13 2 2 1 10 3 13 10 2 3 3 2 2
43 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 2 11 11 2 11 11 7 13 0 2 13 14 9 15 14 11 3 1 10 9 2
28 10 9 10 9 2 0 2 1 9 10 9 2 13 9 0 2 2 13 14 15 3 1 9 0 14 9 15 2
65 11 13 9 0 16 2 13 10 10 9 9 0 2 2 3 0 1 9 9 15 2 11 11 2 2 13 1 9 15 14 9 15 11 2 11 2 13 14 15 14 9 15 1 9 10 9 2 13 14 9 7 13 16 13 1 9 15 10 9 16 1 15 15 13 2
9 10 9 13 9 10 9 10 15 2
25 11 2 9 11 10 0 7 10 0 2 11 11 2 2 13 1 10 9 1 9 9 15 1 9 2
26 10 9 13 1 10 9 1 10 9 10 0 7 10 9 2 16 1 9 13 7 15 13 9 10 9 2
49 7 15 3 9 2 7 15 13 3 1 11 9 11 2 11 11 2 2 11 13 1 9 15 7 1 15 10 9 10 9 2 10 9 7 10 9 2 16 9 13 1 15 14 13 10 9 10 0 2
11 3 9 13 2 16 15 13 3 1 9 2
16 10 9 16 13 1 10 9 7 10 9 14 11 0 3 3 2
81 10 9 13 1 9 10 9 10 0 1 9 1 9 2 9 10 9 10 0 13 9 0 2 7 3 13 10 9 1 9 2 16 11 7 10 9 13 14 10 9 14 15 2 1 9 7 9 2 1 10 9 14 10 9 2 13 1 15 11 11 2 1 9 9 0 2 7 13 1 11 11 14 2 9 9 10 9 14 15 2 2
21 1 10 9 3 2 1 10 9 7 1 9 10 9 2 13 9 9 1 9 0 2
49 9 10 9 2 11 2 13 1 10 9 2 1 9 10 9 10 0 1 9 15 2 12 2 1 9 12 1 10 9 2 2 1 11 2 3 15 13 1 9 15 9 9 1 9 9 15 12 9 2
19 1 15 13 2 1 9 9 16 13 2 1 9 9 9 7 1 9 15 2
47 2 9 1 9 0 2 13 1 9 9 2 9 2 1 10 12 7 1 10 12 1 11 1 10 9 2 1 10 12 1 11 1 9 12 7 1 10 12 1 11 1 9 12 1 10 9 2
46 9 9 16 1 15 9 16 13 1 13 0 3 2 2 13 9 1 9 9 0 1 10 9 2 16 9 10 9 0 2 10 9 14 15 13 1 9 1 10 9 16 13 2 11 2 2
28 1 10 9 13 2 1 10 9 2 16 2 9 10 9 10 0 14 9 9 9 13 14 10 9 1 0 2 2
53 3 13 10 9 1 10 9 16 13 14 10 9 16 13 1 9 15 2 13 10 10 9 2 1 9 0 2 2 9 9 9 2 2 2 16 10 9 10 0 1 10 9 10 0 13 10 9 16 13 1 11 12 2
13 1 10 9 13 9 16 13 14 9 9 10 9 2
36 10 9 2 16 1 13 0 13 13 1 9 9 10 9 7 9 15 10 0 2 13 1 10 9 13 9 0 2 7 3 13 1 15 9 0 2
19 3 2 15 13 2 3 10 13 3 1 9 9 2 7 1 9 9 0 2
24 3 2 2 9 10 9 10 0 2 9 15 16 1 15 13 9 3 1 4 13 14 9 15 2
18 3 2 10 9 2 15 13 1 15 2 1 9 15 2 13 12 9 2
17 1 9 15 1 15 15 13 2 2 3 3 9 7 3 10 9 2
11 3 10 9 13 9 14 10 13 10 0 2
18 13 7 13 9 1 9 9 0 7 13 10 9 16 13 0 1 15 2
7 3 2 9 2 9 2 2
32 3 13 14 15 13 3 13 14 10 9 10 0 15 1 9 10 9 2 16 13 3 1 10 9 10 0 2 9 9 9 2 2
75 13 16 9 10 9 13 1 10 9 1 10 9 2 10 9 2 1 9 9 0 1 9 9 0 2 13 14 10 9 2 9 2 2 3 1 10 15 2 9 2 2 2 7 3 13 13 14 10 9 2 9 2 1 9 0 2 9 0 13 14 2 9 2 2 9 10 9 13 1 2 9 2 7 3 2
27 1 3 13 10 2 9 2 2 7 2 3 13 10 2 9 16 13 1 13 0 3 2 1 9 10 9 2
25 1 9 10 9 13 1 9 13 2 7 3 13 3 9 13 12 2 10 10 9 13 1 9 12 2
103 1 9 2 7 1 9 0 4 10 13 13 1 10 9 1 9 2 16 10 9 13 1 15 12 9 1 10 9 7 10 9 16 13 1 10 9 2 9 2 15 4 13 1 9 1 9 3 1 9 12 2 7 1 10 9 10 0 13 10 13 9 0 1 9 14 9 0 2 7 3 9 9 2 16 16 13 10 13 1 9 2 1 16 13 1 10 9 12 9 13 1 9 9 13 1 9 12 1 9 3 1 9 2
62 3 3 2 13 2 3 1 9 1 10 9 16 13 1 9 9 0 1 9 9 10 9 2 1 15 2 10 9 10 0 13 13 1 9 10 9 2 16 7 13 13 14 2 10 9 16 13 1 13 0 3 2 2 13 1 10 9 1 9 1 9 2
27 1 10 9 14 10 9 10 0 13 13 1 9 11 2 16 13 1 1 12 9 7 13 1 9 14 9 2
3 9 0 2
51 10 0 13 2 16 15 9 0 2 1 15 1 9 0 2 13 1 10 13 9 0 2 9 16 1 15 9 9 2 7 1 16 13 1 10 9 16 13 1 13 0 3 2 2 7 9 9 1 9 12 2
8 9 15 3 13 1 10 9 2
15 10 9 13 1 9 15 2 3 13 1 10 9 16 13 2
31 13 14 15 7 13 4 3 1 9 10 9 2 1 9 10 9 7 2 3 2 1 9 9 9 10 9 10 0 14 15 2
40 10 10 9 16 13 3 1 10 13 10 0 2 13 14 15 1 9 2 13 7 13 2 7 7 3 2 9 2 1 9 9 9 13 9 16 4 1 9 0 2
75 10 9 1 9 7 1 9 13 1 3 1 3 2 1 9 9 15 1 13 7 9 2 14 10 9 2 9 0 9 2 2 7 13 3 16 10 9 2 10 9 2 1 9 15 13 2 1 9 10 9 2 1 12 9 1 12 9 2 7 3 1 10 9 10 0 2 7 7 9 1 9 13 9 0 2
10 4 13 14 10 9 1 9 3 0 2
15 1 10 9 2 10 9 13 3 3 1 9 9 10 9 2
35 13 14 9 10 9 10 0 2 11 12 2 11 12 2 2 10 9 10 0 13 1 12 9 2 9 10 9 1 9 13 1 12 9 3 2
24 13 16 13 1 15 9 2 13 4 1 9 0 7 3 13 13 9 0 10 9 0 1 15 2
20 15 13 2 16 10 9 1 9 0 1 9 15 3 7 10 9 16 13 9 2
18 7 15 2 9 9 1 9 14 12 9 1 11 12 13 9 0 0 2
50 7 13 9 10 9 13 14 10 9 3 1 10 9 10 0 9 1 9 13 9 0 3 2 3 3 16 10 9 4 1 9 1 10 9 2 10 9 0 7 9 10 9 2 10 9 7 10 9 0 2
44 9 11 1 9 9 2 2 11 2 2 3 3 13 14 10 9 2 7 1 15 13 1 15 1 15 3 2 3 13 1 9 16 13 9 13 12 9 1 10 9 2 1 12 2
27 13 1 15 9 14 9 15 1 9 9 1 10 9 2 16 13 9 2 9 1 9 1 9 12 9 2 2
26 9 16 13 1 9 15 1 10 9 2 13 12 9 2 12 1 9 10 9 7 12 3 1 10 9 2
8 3 13 1 10 9 10 15 2
50 1 9 0 13 1 9 2 11 2 13 14 9 10 9 1 9 12 9 2 16 10 9 13 1 9 10 9 2 7 7 13 2 16 7 10 9 3 13 14 9 10 13 16 13 3 14 9 10 9 2
27 1 9 15 13 2 16 9 2 11 2 4 13 14 10 9 1 9 3 7 1 15 4 13 1 9 15 2
25 2 3 3 2 2 13 10 9 10 0 11 11 11 2 2 15 9 16 15 13 1 9 0 3 2
13 7 1 10 9 15 4 13 3 2 3 3 3 2
16 3 3 13 1 9 0 1 9 15 2 3 3 13 13 2 2
34 11 11 13 1 3 16 13 1 9 1 12 10 9 16 1 15 13 14 9 15 10 0 7 0 10 9 2 1 9 15 13 1 9 2
33 15 13 16 15 13 2 7 3 1 15 15 2 13 9 0 2 1 16 10 9 13 1 9 15 14 11 11 2 9 0 2 0 2
38 9 10 9 14 11 11 13 2 1 9 15 2 1 9 10 9 14 15 1 10 9 14 11 7 9 15 16 10 9 4 13 7 13 1 9 9 0 2
49 7 1 9 15 1 10 11 10 0 16 1 9 15 1 10 11 10 0 14 15 13 10 9 10 0 2 10 0 7 9 10 9 10 0 16 2 9 15 3 13 0 2 1 9 15 1 10 9 2
10 3 3 15 13 1 9 15 10 0 2
60 10 9 10 0 7 10 0 1 10 9 2 1 9 10 9 10 0 2 2 16 13 15 3 1 9 10 9 1 10 9 2 11 2 11 11 11 2 2 13 16 13 1 9 1 12 1 10 9 14 9 15 2 1 9 10 9 14 9 9 2
31 1 10 9 15 13 16 9 15 10 0 3 13 3 14 9 15 1 9 15 10 0 1 9 15 10 0 14 9 10 9 2
24 10 9 9 11 2 9 9 9 2 13 9 1 10 9 2 1 13 9 0 13 7 0 3 2
57 9 15 13 1 9 10 9 7 9 10 9 14 9 10 9 16 15 13 1 9 15 10 0 11 11 2 1 9 15 1 9 0 7 1 9 15 1 9 9 0 2 1 10 9 10 0 7 10 0 16 15 13 1 9 9 9 2
20 10 9 16 12 1 15 13 1 10 9 13 14 9 15 10 0 14 9 11 2
33 10 9 13 14 9 15 1 9 15 2 7 11 11 2 16 15 3 13 1 15 12 9 2 13 1 10 10 9 9 7 9 0 2
37 15 1 16 9 15 14 9 11 1 9 15 10 0 2 9 13 2 13 1 9 11 0 15 2 7 11 11 13 16 13 1 15 9 1 14 15 2
44 2 10 9 13 1 9 16 13 1 10 9 1 13 1 9 0 0 2 1 13 13 9 0 7 3 0 2 2 13 11 11 9 10 12 14 13 3 1 3 1 11 2 11 2
28 2 15 13 16 1 10 15 13 10 9 2 15 13 1 10 9 14 15 9 2 9 16 1 15 15 13 2 2
22 1 13 14 9 15 10 0 1 9 13 10 9 2 2 9 13 9 1 9 10 9 2
7 15 9 13 14 9 15 2
8 1 9 13 10 9 1 9 2
13 7 10 9 13 9 0 12 9 15 13 1 9 2
18 7 15 13 9 14 9 10 9 13 9 2 9 2 9 7 9 2 2
20 16 13 3 13 1 9 0 13 11 11 16 15 13 16 10 9 13 1 15 2
29 2 10 9 1 15 13 0 1 0 1 9 10 9 14 15 15 2 9 16 13 1 10 9 14 15 2 2 13 2
7 7 13 3 9 0 3 2
15 10 9 13 1 10 9 2 15 9 10 9 14 10 9 2
16 11 11 13 16 1 9 10 9 9 15 13 9 1 10 9 2
15 2 15 13 0 1 9 15 14 10 9 2 2 15 13 2
36 2 7 10 9 13 16 3 3 9 0 7 0 0 7 3 15 9 7 9 0 15 16 1 15 15 13 2 13 1 10 9 7 13 14 15 2
21 13 1 10 9 9 0 1 14 15 2 16 16 15 13 16 10 9 13 1 15 2
8 15 9 1 9 10 9 2 2
31 9 15 9 13 1 10 9 1 9 9 9 2 1 10 9 13 9 15 1 9 15 10 3 2 0 7 10 0 2 0 2
27 1 16 13 1 10 3 13 7 13 1 9 15 10 0 2 13 11 11 1 9 10 9 16 13 14 15 2
20 2 9 12 2 16 13 14 9 15 2 13 1 9 15 10 9 13 1 9 2
21 15 13 9 9 7 0 2 7 3 13 13 3 13 10 9 16 1 15 13 2 2
29 1 12 9 15 1 9 2 16 1 15 13 3 1 12 9 13 11 11 15 3 13 1 9 9 1 16 13 3 2
57 1 9 15 1 9 1 2 9 1 9 2 7 2 9 15 10 0 14 11 11 2 2 16 1 15 10 9 13 11 1 9 15 7 9 15 2 10 9 1 2 1 9 10 9 10 0 2 13 3 0 7 0 2 13 7 0 2
17 2 9 1 9 9 13 9 3 0 1 15 2 2 13 10 9 2
5 2 15 0 3 2
7 7 3 13 1 10 9 2
12 1 9 9 10 9 14 15 0 7 3 13 2
20 7 9 15 1 9 7 9 13 9 13 7 0 2 9 16 13 9 7 9 2
17 10 9 3 13 9 0 1 13 1 10 9 14 9 7 9 9 2
7 13 14 15 9 0 2 2
7 10 9 13 10 9 0 2
9 11 11 13 1 9 1 13 9 2
18 2 10 9 13 14 15 13 2 2 15 13 2 2 3 9 13 9 2
12 15 9 7 13 1 15 3 3 1 9 2 2
18 9 16 9 15 3 3 9 10 9 7 3 9 1 10 9 9 15 2
27 1 9 9 9 15 13 2 7 7 3 1 10 9 10 0 1 10 9 16 13 1 15 1 3 9 15 2
9 9 10 9 10 0 13 13 15 2
16 9 10 9 14 10 9 1 11 13 1 9 0 1 10 9 2
43 3 1 16 2 10 9 10 0 2 0 12 9 2 4 9 10 9 2 1 2 9 9 12 1 9 10 9 10 0 2 13 9 1 14 15 1 9 1 10 9 10 0 2
39 7 7 10 9 13 1 9 0 2 7 7 9 15 13 13 14 15 7 3 3 1 10 9 14 15 2 4 3 13 14 9 15 14 9 10 9 14 15 2
26 10 9 10 0 13 1 2 9 15 10 0 14 10 9 10 0 2 2 13 9 1 9 9 1 11 2
20 1 9 14 13 9 13 15 9 0 0 1 9 9 2 11 2 11 2 11 2
21 9 7 9 2 9 9 2 9 9 7 9 0 13 9 9 15 14 9 0 0 2
14 10 9 13 13 9 2 13 10 9 10 0 11 11 2
7 9 9 13 1 9 0 2
14 1 1 15 2 2 10 9 13 13 1 10 9 2 2
12 15 13 3 0 1 9 13 7 1 9 13 2
17 10 9 1 10 9 10 0 7 10 9 13 9 0 1 10 9 2
71 10 9 3 13 1 2 9 0 2 14 9 15 2 13 10 9 10 0 1 9 2 9 1 11 2 11 11 2 10 9 13 2 4 1 15 13 7 15 4 13 9 2 2 13 1 10 9 7 13 14 9 15 1 2 9 9 16 13 0 7 9 9 2 2 9 16 13 4 1 9 2
27 3 10 10 9 1 9 9 2 9 16 13 1 10 9 1 9 0 1 11 13 1 9 9 2 13 11 2
18 9 7 9 0 16 13 1 9 0 13 3 12 1 9 14 9 0 2
13 15 13 14 9 15 7 13 9 2 9 13 13 2
17 10 9 4 13 3 1 9 0 2 16 9 0 13 1 9 0 2
15 16 13 1 9 10 9 4 9 13 0 3 1 9 15 2
26 9 9 12 13 1 10 9 3 13 9 15 9 10 12 1 9 0 7 13 13 14 15 1 9 9 2
13 10 9 13 13 9 9 7 9 13 14 15 9 2
45 9 9 1 9 16 1 9 15 9 0 3 2 9 1 9 15 2 15 7 9 1 9 10 9 1 9 0 13 9 0 13 14 9 15 1 9 3 3 1 15 16 13 1 15 2
22 10 9 10 0 11 11 2 11 13 16 9 13 13 1 9 15 14 10 9 1 9 2
34 11 2 11 2 9 9 9 7 9 1 9 9 16 4 13 2 13 1 9 15 14 9 2 16 9 15 9 10 12 13 1 10 9 2
31 1 9 3 13 10 9 16 1 9 12 13 10 9 14 9 9 10 9 14 15 2 16 16 10 9 13 13 3 9 12 2
13 10 9 13 9 9 16 10 9 13 1 10 9 2
8 10 9 13 1 9 10 9 2
12 10 9 13 14 10 9 9 3 1 10 15 2
13 3 13 10 9 1 9 7 13 1 9 10 9 2
18 3 0 9 13 13 9 1 9 10 9 13 1 9 16 13 1 9 2
14 15 13 14 10 9 10 0 1 11 1 13 14 15 2
41 1 11 11 2 12 2 2 9 9 9 2 9 2 13 10 9 1 12 9 15 2 11 9 10 12 7 11 9 10 12 2 16 16 13 13 14 15 1 9 9 2
27 12 9 1 1 3 13 9 15 2 11 11 2 1 9 16 1 15 13 10 9 2 13 14 15 1 9 2
17 1 9 9 0 13 10 9 9 7 9 9 7 13 1 10 9 2
16 15 13 13 14 9 15 1 9 1 11 1 13 14 15 3 2
41 1 9 11 2 11 11 2 11 13 11 2 13 1 10 9 16 13 3 1 10 9 10 0 7 13 1 9 10 9 2 2 13 14 15 2 9 13 14 15 2 2
13 10 9 7 10 9 13 7 10 9 13 9 9 2
25 9 9 9 1 9 16 13 1 9 0 1 11 2 13 1 9 9 0 0 14 9 1 9 15 2
22 3 12 2 1 3 13 14 9 10 9 14 10 9 2 13 10 9 9 0 7 0 2
16 13 9 0 0 1 10 9 2 7 9 0 4 13 9 0 2
23 3 12 9 7 9 0 1 9 12 2 12 13 1 3 12 1 9 10 9 11 1 11 2
8 3 9 2 10 9 13 13 2
12 10 9 2 13 9 2 2 13 9 10 9 2
13 9 1 9 7 3 2 9 13 13 14 14 15 2
24 1 9 0 1 9 2 9 0 13 9 3 7 3 2 16 16 4 13 11 11 2 9 12 2
29 1 9 10 9 10 0 13 10 9 1 9 3 3 1 15 1 9 2 2 15 13 14 15 3 16 3 13 2 2
30 16 9 9 2 10 9 10 0 11 1 11 13 1 11 13 1 9 9 15 13 13 1 9 2 9 0 0 1 11 2
16 3 3 13 1 15 9 1 10 9 7 13 9 1 9 9 2
21 11 13 1 10 9 1 9 9 7 1 9 0 7 13 9 1 9 7 1 9 2
29 3 2 9 14 10 9 10 0 1 11 1 9 0 13 1 9 0 10 9 1 9 9 2 7 3 1 9 9 2
26 1 9 12 13 9 15 14 11 1 9 2 10 9 2 16 3 13 13 3 1 9 15 1 9 0 2
13 15 13 7 15 3 9 1 9 9 9 7 9 2
13 7 13 1 15 9 2 13 2 13 1 15 9 2
5 7 9 10 9 2
23 2 9 2 9 2 2 13 11 2 2 15 13 1 15 1 10 9 7 13 1 15 2 2
19 3 4 16 10 9 13 1 9 2 9 0 7 13 3 2 13 10 9 2
10 2 10 3 13 13 13 9 9 2 2
6 9 15 13 13 9 2
24 9 0 13 3 9 13 7 13 1 9 15 14 10 9 2 7 9 15 10 13 13 14 15 2
24 9 1 15 2 1 9 10 9 13 10 9 1 9 1 9 10 9 10 12 1 9 10 9 2
13 1 11 13 9 10 9 1 9 9 1 10 9 2
18 13 9 9 7 10 9 13 13 1 9 15 16 1 10 9 13 9 2
15 1 12 9 13 10 9 10 0 16 13 3 1 9 0 2
25 3 4 13 1 9 10 9 14 9 10 9 2 16 3 13 13 1 15 10 2 3 1 9 0 2
33 9 9 10 12 2 13 1 10 9 2 9 9 0 0 7 3 0 2 13 10 9 10 0 1 9 15 16 13 1 15 9 9 2
21 1 10 9 15 13 13 10 9 1 16 4 13 1 15 3 3 9 1 14 15 2
14 3 3 13 9 15 2 1 9 11 2 13 1 11 2
22 11 9 10 12 7 11 9 10 12 13 3 15 13 1 10 9 7 13 9 1 15 2
10 2 3 3 2 3 2 2 13 11 2
11 11 11 13 16 16 13 3 15 9 15 2
37 9 0 2 9 1 11 2 11 11 2 13 16 1 10 9 14 9 13 1 11 2 2 9 1 9 7 9 2 2 13 16 15 2 1 9 2 2
12 3 4 16 9 16 13 9 13 1 15 9 2
31 10 9 13 1 10 9 2 9 2 11 2 2 16 0 1 9 10 11 2 2 1 9 9 10 9 16 13 1 10 9 2
18 3 13 1 15 16 13 1 9 9 2 7 16 10 9 13 1 9 2
23 16 16 13 9 0 7 10 9 3 13 2 13 1 10 9 1 9 10 9 1 10 9 2
31 1 9 15 14 9 10 9 1 9 9 2 9 11 11 2 13 9 10 11 16 13 14 10 10 9 10 0 1 9 0 2
46 9 10 9 7 9 10 11 2 11 11 2 13 1 9 1 9 15 16 3 13 9 1 10 9 7 3 13 1 10 9 10 9 10 9 0 7 1 15 13 10 9 2 1 9 2 2
21 10 9 11 13 14 9 15 1 9 1 9 0 2 16 1 9 15 3 15 13 2
24 13 1 9 1 9 2 11 2 2 16 13 7 15 1 11 2 1 9 9 11 1 10 11 2
22 1 10 9 13 1 11 2 2 9 0 1 9 15 2 7 3 2 9 2 12 9 2
18 1 9 0 13 1 11 2 2 9 0 0 2 1 9 9 10 9 2
23 1 12 10 9 10 9 1 11 13 2 2 0 1 9 0 9 2 9 9 12 9 2 2
24 13 10 13 2 7 10 9 0 1 9 0 9 2 3 4 16 15 13 9 3 0 14 9 2
35 9 9 10 9 1 9 10 9 2 11 11 2 16 13 14 10 9 2 13 16 1 9 15 2 10 9 13 1 9 1 10 9 10 0 2
24 13 2 16 7 1 10 9 10 0 2 3 10 9 10 0 13 13 14 9 10 9 1 9 2
17 13 10 9 2 3 10 9 10 0 14 9 7 13 1 9 0 2
51 11 13 2 16 1 9 10 9 13 14 10 9 7 13 1 15 14 10 9 2 1 9 0 13 1 9 9 12 9 9 2 7 7 1 9 0 1 12 9 9 2 2 7 3 13 1 10 9 10 0 2
21 11 13 2 16 1 7 16 10 9 13 1 10 9 2 13 1 15 3 1 13 2
8 9 2 4 13 14 10 9 2
5 1 2 10 9 2
23 10 9 13 1 10 9 10 0 7 13 14 1 10 9 14 9 10 9 7 9 10 9 2
16 9 12 13 1 10 9 14 10 9 2 7 0 1 10 9 2
26 10 9 13 1 10 9 10 0 14 9 10 9 7 10 9 7 13 3 1 9 10 9 14 9 11 2
14 10 9 13 9 1 11 7 9 0 1 9 7 9 2
12 9 0 0 3 13 3 2 7 13 12 9 2
27 1 13 1 9 10 9 2 13 10 9 14 9 10 9 14 10 9 2 7 13 14 9 15 1 10 9 2
15 9 1 9 1 10 15 13 1 12 9 2 13 9 2 2
30 9 16 13 1 9 0 4 13 1 10 9 1 9 0 7 13 1 12 9 10 9 1 10 9 7 1 9 10 9 2
53 9 1 10 9 10 0 1 9 9 2 16 13 16 10 3 16 13 1 15 9 7 9 9 13 13 9 1 9 10 9 9 15 2 13 9 11 2 16 15 9 9 0 2 16 1 9 9 0 4 13 9 9 2
32 11 11 2 16 9 9 15 13 1 9 12 7 3 2 13 1 9 10 9 10 0 2 16 13 1 9 14 10 9 10 0 2
36 15 13 9 1 9 9 7 1 9 1 9 1 11 11 7 11 11 2 16 13 1 9 15 13 1 9 14 3 9 7 7 13 1 15 9 2
25 11 13 14 10 9 7 13 14 15 9 1 9 2 3 1 15 7 1 2 15 1 9 7 9 2
22 1 9 13 9 10 9 1 15 7 15 13 13 9 1 9 2 9 7 1 9 0 2
34 1 9 2 3 13 13 1 9 10 9 1 10 9 1 10 9 16 13 1 9 9 0 1 9 2 10 9 11 11 1 9 2 12 2
12 15 13 3 9 7 13 1 15 1 9 0 2
30 11 13 2 16 13 1 15 9 7 9 1 16 13 1 9 0 2 16 16 13 10 9 1 9 7 3 13 1 9 2
32 9 15 13 1 10 9 0 2 14 1 9 15 10 9 16 10 9 10 0 13 15 16 13 1 10 9 7 1 9 10 9 2
22 9 0 2 9 0 7 9 2 4 13 1 9 1 9 10 9 7 1 9 10 9 2
17 3 13 11 11 3 2 3 1 9 0 2 1 9 7 9 9 2
22 15 3 13 1 9 15 1 9 1 9 16 13 1 9 9 0 9 2 9 7 3 2
40 2 1 10 9 10 0 2 2 13 11 2 2 9 10 9 13 9 14 9 10 9 7 4 13 1 10 12 2 16 16 3 4 13 1 9 0 7 9 9 2
33 1 10 9 10 0 2 1 15 2 9 10 9 13 1 10 9 10 0 7 9 9 13 1 10 9 10 0 7 3 10 0 2 2
31 1 9 1 10 9 13 9 0 1 9 1 9 0 2 13 11 2 16 16 15 4 9 1 10 9 2 3 9 0 0 2
15 16 13 2 13 9 16 9 15 13 7 13 14 10 9 2
19 7 16 10 9 4 13 1 9 0 2 9 10 9 4 9 0 7 0 2
9 4 13 15 1 9 9 9 0 2
37 16 13 9 9 2 1 10 9 10 0 3 7 1 1 10 0 2 13 16 10 9 13 13 1 9 13 7 10 9 13 1 9 7 3 0 3 2
19 1 9 15 1 9 2 10 9 7 9 10 9 13 9 1 9 10 9 2
25 10 9 2 13 11 2 4 13 0 1 10 9 7 1 9 15 7 3 3 1 10 9 10 0 2
14 2 9 1 9 9 13 9 14 10 9 7 10 9 2
27 7 9 13 9 9 3 1 9 9 0 2 15 4 13 14 10 9 10 10 9 1 13 14 3 16 13 2
33 9 16 13 3 9 0 13 1 10 9 13 1 15 14 10 9 10 0 1 9 0 1 10 9 2 7 3 13 3 9 1 9 2
24 15 13 14 10 9 13 14 9 15 16 16 13 1 10 9 2 14 13 1 15 9 0 2 2
34 10 9 10 0 1 9 10 9 13 9 9 16 13 1 10 9 10 0 1 10 9 2 16 1 15 9 0 1 9 10 9 10 0 2
36 2 9 10 9 13 0 7 0 2 2 13 11 2 2 7 4 13 2 16 16 9 0 4 13 9 7 1 9 0 1 9 9 10 9 2 2
34 10 9 2 2 13 1 9 15 1 9 12 2 1 9 12 7 12 2 14 15 13 1 15 9 0 16 13 1 3 3 1 12 9 2
17 13 2 16 3 10 3 16 13 1 9 15 3 13 1 9 15 2
38 11 2 16 13 9 9 9 2 13 1 9 15 1 9 0 2 3 1 9 0 2 1 9 15 7 1 9 15 14 13 1 10 9 7 9 1 12 2
35 9 1 10 9 15 13 1 9 15 14 0 2 9 13 7 13 1 2 9 9 9 16 13 1 15 2 7 9 2 3 2 3 13 3 2
18 1 9 0 13 11 9 0 14 9 1 9 15 14 10 9 11 11 2
27 10 9 13 13 1 9 15 9 7 9 14 9 7 15 13 13 14 10 2 9 2 1 9 15 10 0 2
41 1 9 0 2 16 13 1 12 1 9 11 1 9 10 12 14 10 12 10 0 2 13 10 9 1 9 1 12 1 9 15 14 11 7 1 3 13 1 9 0 2
47 11 11 10 9 2 9 2 10 9 1 10 9 2 2 13 1 10 9 2 7 1 9 10 9 13 1 9 15 2 16 13 1 10 9 2 2 15 10 9 3 0 14 15 2 9 2 2
35 10 9 3 13 14 9 9 15 2 13 9 0 1 9 15 2 7 13 2 2 13 1 15 3 9 12 0 1 15 2 7 15 15 2 2
18 11 10 9 13 1 9 1 16 13 9 10 9 16 13 14 10 9 2
29 2 4 13 15 2 9 2 2 15 13 1 9 2 2 1 9 2 14 15 13 1 15 13 1 9 15 3 2 2
50 1 10 9 2 9 10 9 2 2 1 11 11 10 9 2 13 10 9 11 2 9 16 9 15 13 13 1 15 9 2 3 1 9 15 2 2 9 1 10 9 2 16 13 1 9 9 0 7 0 2
44 10 9 2 1 9 15 10 0 2 13 3 2 16 3 4 13 1 11 14 10 10 9 16 13 1 15 2 7 3 13 1 15 16 10 10 9 16 13 1 9 15 3 13 2
35 1 9 13 10 9 9 12 1 9 9 15 14 11 1 9 10 9 10 0 10 0 2 12 1 10 12 2 12 1 10 12 7 3 3 2
27 11 13 14 9 10 9 7 13 1 10 9 16 13 1 9 15 9 10 9 16 13 3 3 1 10 9 2
20 15 13 1 15 9 0 7 13 1 9 15 14 9 0 2 3 1 9 15 2
33 11 13 14 9 15 1 10 9 10 0 16 1 2 11 2 2 1 9 12 2 7 2 9 11 7 9 11 2 2 1 9 12 2
44 11 2 16 13 9 3 2 13 1 10 9 7 1 10 9 10 0 10 13 1 15 2 7 9 15 16 15 13 14 10 9 15 7 13 14 9 10 9 10 0 7 10 0 2
33 9 15 0 1 9 15 14 10 9 1 10 9 10 9 2 1 1 12 7 12 9 16 1 15 15 9 2 9 1 10 9 0 2
21 3 1 9 15 13 1 15 9 15 14 9 10 9 2 16 13 13 1 9 11 2
11 10 9 13 1 10 9 7 4 13 13 2
23 1 11 13 2 16 13 13 14 9 15 1 9 7 1 15 13 13 1 9 15 9 0 2
4 2 9 2 2
5 2 3 10 9 2
4 2 9 2 2
5 2 9 15 2 2
27 3 13 10 9 14 9 15 7 13 13 1 15 1 9 2 7 3 13 1 10 9 9 0 14 9 13 2
16 1 9 0 1 12 9 13 11 7 10 9 1 9 9 0 2
19 9 10 9 3 13 2 7 10 9 10 13 13 9 13 3 1 15 9 2
105 1 10 9 1 10 9 13 3 9 1 10 9 10 15 2 16 9 15 1 11 13 9 1 12 2 16 15 13 13 3 1 10 9 14 10 9 10 0 1 11 2 10 3 16 13 1 15 9 1 9 15 7 0 1 10 9 10 0 2 13 16 13 3 9 0 1 10 13 1 10 9 1 10 9 16 4 13 1 10 9 2 7 10 9 15 2 3 2 4 13 0 2 7 3 3 1 10 9 14 11 11 1 9 9 2
8 9 9 1 10 9 9 15 2
24 1 9 10 9 1 10 9 2 7 9 9 0 13 1 9 9 10 9 1 10 9 10 0 2
56 11 11 2 9 9 10 9 1 11 2 13 1 10 9 7 13 9 1 2 11 2 1 11 2 9 10 9 1 11 7 1 11 2 9 10 9 10 0 1 11 2 9 10 9 9 9 1 9 2 10 11 7 3 13 0 2
36 1 9 15 14 9 11 1 11 13 9 1 9 12 1 9 3 2 0 1 9 2 9 1 9 2 2 16 13 1 11 16 1 11 3 9 2
15 10 9 1 9 2 13 11 2 13 13 3 1 9 0 2
12 13 1 15 12 9 0 0 2 0 7 0 2
14 10 9 10 0 13 1 10 9 1 9 0 7 0 2
22 9 0 13 14 10 9 7 13 14 15 2 7 4 13 9 16 13 0 1 10 9 2
34 9 0 2 1 0 2 0 7 0 2 13 1 9 14 0 2 1 9 0 2 1 0 7 0 2 16 13 1 9 9 2 1 0 2
25 10 9 10 0 13 1 10 9 16 1 9 15 13 0 3 2 1 16 9 0 13 14 10 9 2
13 10 10 9 15 13 1 9 1 9 9 10 9 2
17 1 9 9 9 9 1 9 9 2 7 2 13 11 1 9 0 2
17 4 1 15 13 7 10 9 1 10 9 13 1 9 0 7 0 2
33 3 13 14 9 10 9 1 9 13 7 1 9 16 13 14 10 9 10 3 0 1 12 9 9 1 15 9 9 2 2 15 13 2
10 10 9 10 12 13 10 9 10 0 2
10 10 9 13 1 10 9 7 13 9 2
22 9 0 2 1 9 2 13 9 2 9 0 13 9 9 9 7 9 0 13 9 9 2
13 11 13 13 1 9 10 9 1 10 9 10 0 2
12 9 0 1 9 13 1 9 9 1 9 0 2
33 1 9 10 13 11 1 11 13 11 9 0 2 16 13 1 12 9 9 10 13 2 1 9 14 0 1 0 9 7 1 0 0 2
19 2 10 9 10 0 1 0 1 0 13 1 9 9 1 10 9 10 0 2
29 1 15 2 10 9 10 0 13 9 0 2 7 1 9 10 9 16 13 14 9 15 1 10 9 1 9 13 2 2
15 3 10 9 10 0 13 14 11 1 9 15 1 9 0 2
28 15 13 15 10 9 10 0 7 10 0 14 10 9 2 15 9 10 9 2 15 9 13 9 10 9 7 3 2
31 9 15 13 1 9 9 3 1 9 9 0 2 16 13 1 9 0 7 0 13 1 15 14 10 9 7 13 14 10 9 2
33 1 10 9 1 9 9 11 2 7 2 13 11 1 9 10 0 14 10 9 7 9 10 9 7 10 9 13 1 9 0 2 0 2
26 1 9 10 9 13 11 9 2 9 14 10 9 2 13 1 9 15 7 13 9 1 10 9 10 0 2
20 1 9 10 9 7 9 10 9 1 9 1 10 10 9 2 13 9 10 9 2
20 11 13 1 10 9 7 13 13 9 1 9 9 10 9 7 10 9 10 0 2
41 2 3 13 2 2 13 11 2 2 16 1 10 9 16 13 7 9 15 13 13 9 10 9 14 10 9 2 7 1 9 1 15 13 3 9 15 7 9 15 2 2
45 9 15 13 13 1 9 14 9 10 9 1 10 9 10 0 2 7 13 14 9 11 1 9 2 9 1 9 0 2 16 13 14 10 9 7 13 1 10 9 16 13 1 10 9 2
21 0 13 1 9 10 9 9 9 2 16 13 1 9 9 2 9 2 9 9 0 2
37 15 9 16 13 1 9 10 9 1 10 9 16 1 15 13 1 9 15 2 16 16 13 1 9 9 1 10 9 2 1 10 9 7 1 10 9 2
48 14 9 9 13 1 9 10 12 11 11 2 9 15 14 9 11 7 11 11 2 16 13 1 9 10 12 14 10 12 10 0 14 9 10 9 7 14 9 15 1 10 9 16 13 1 10 9 2
34 9 11 7 11 11 13 14 10 9 1 9 10 9 7 10 9 10 0 1 10 9 10 0 2 7 13 14 9 9 10 9 7 11 2
37 1 9 15 13 10 9 9 9 2 16 1 15 13 9 14 9 7 9 2 16 13 1 9 10 9 7 1 10 9 1 10 9 16 1 9 15 2
21 10 9 10 0 2 16 9 15 12 9 2 13 1 9 9 2 13 1 9 13 2
29 10 9 13 1 9 1 9 2 7 1 10 12 1 15 13 9 16 13 9 0 2 9 7 9 1 9 10 9 2
20 1 9 9 9 16 13 1 10 9 13 10 9 1 9 10 9 1 10 9 2
27 3 13 1 10 9 10 9 1 9 10 9 2 10 9 7 10 9 1 9 10 9 2 9 1 10 9 2
29 9 11 2 7 2 13 1 10 9 1 9 14 9 9 7 9 2 13 1 9 9 0 7 13 1 9 10 9 2
35 9 10 9 13 14 9 15 14 9 10 9 2 16 13 1 9 9 15 1 9 9 10 9 2 7 1 10 9 13 9 1 9 10 9 2
13 10 9 10 0 13 1 12 1 12 9 10 12 2
11 10 9 13 1 9 13 1 9 1 9 2
53 3 13 1 9 11 1 9 9 10 9 7 10 9 2 16 1 15 13 9 11 7 1 9 15 9 9 2 9 2 2 13 1 9 9 16 13 1 10 9 7 1 10 9 7 13 14 9 10 9 1 9 11 2
9 10 9 13 1 9 9 10 9 2
11 13 9 16 13 9 0 1 9 9 0 2
45 1 16 1 9 11 13 1 12 10 9 1 12 10 9 2 7 1 9 10 9 13 1 9 1 9 2 1 9 11 9 15 13 1 9 9 10 11 2 16 14 15 13 9 11 2
44 14 10 9 13 1 10 9 16 13 1 9 10 9 1 9 12 10 9 2 7 9 15 3 13 3 1 9 10 9 2 3 15 13 1 9 10 9 2 9 2 7 10 9 2
54 3 16 13 1 9 15 14 10 9 2 4 1 15 13 9 15 3 1 9 15 2 1 10 13 2 2 16 13 9 1 10 9 2 9 15 13 1 15 2 7 7 13 1 15 9 9 13 1 15 1 9 0 2 2
11 1 10 9 13 9 0 1 12 10 9 2
35 1 10 9 4 13 1 9 10 9 2 1 15 13 14 10 9 2 7 3 13 2 7 13 10 9 2 13 10 9 2 13 10 9 2 2
30 1 9 15 9 10 9 1 9 15 2 7 1 12 9 10 9 4 13 14 10 9 10 0 1 10 9 1 9 9 2
14 10 9 13 1 10 9 1 9 15 14 9 10 9 2
9 10 9 13 1 9 1 9 0 2
9 1 9 13 9 9 7 9 9 2
21 9 9 1 10 9 7 1 9 10 9 13 12 9 1 9 2 12 9 1 9 2
14 9 10 9 1 10 9 10 0 13 9 2 12 9 2
9 10 9 0 1 9 7 1 9 2
21 1 9 9 13 10 9 1 9 12 2 1 9 7 7 1 9 9 1 12 2 2
12 4 13 14 10 9 3 9 1 9 10 9 2
24 1 9 9 1 9 9 9 13 7 9 0 4 13 1 9 12 2 7 1 11 12 11 12 2
12 10 9 11 4 3 13 1 9 9 1 9 2
43 10 9 13 14 9 15 1 10 9 13 1 10 9 2 14 13 16 2 1 9 0 4 13 1 9 7 9 0 2 2 7 2 1 9 0 2 10 9 13 14 10 9 2
15 11 13 3 14 9 15 1 10 9 2 7 3 14 15 2
10 1 3 10 12 13 1 15 9 0 2
21 1 10 9 16 11 13 16 4 9 0 2 15 13 1 9 15 12 12 9 9 2
45 11 1 9 13 13 9 15 13 9 9 0 2 1 12 9 0 2 1 9 0 2 1 9 11 2 1 9 9 7 3 15 3 14 13 1 9 9 0 1 10 9 7 1 9 2
33 1 9 2 3 10 9 13 9 1 9 9 15 14 9 16 13 1 9 13 1 9 9 2 14 3 15 13 1 2 9 9 0 2
15 15 7 16 13 16 14 10 9 1 9 9 15 4 13 2
37 9 15 14 9 0 9 1 9 13 1 9 9 13 13 1 9 15 1 9 15 2 7 2 14 9 0 1 9 9 1 16 13 1 15 9 0 2
21 9 11 13 13 1 9 0 1 1 13 9 15 2 7 13 14 15 1 9 0 2
9 9 15 14 10 9 15 13 13 2
8 13 1 15 9 9 7 9 2
30 7 1 10 9 9 9 15 13 13 3 9 1 9 10 9 10 0 14 15 2 7 9 15 13 9 9 15 10 0 2
15 9 10 9 13 3 14 9 15 7 13 1 15 9 0 2
39 11 2 1 3 16 13 1 9 9 1 11 16 13 9 1 9 7 9 2 1 11 7 1 10 9 2 1 9 15 13 14 10 9 10 0 14 9 15 2
15 10 9 0 13 14 9 15 16 13 1 10 9 10 0 2
20 1 9 9 14 9 2 13 1 15 1 9 10 9 10 0 10 0 2 0 2
34 15 4 13 2 16 10 9 10 0 16 13 1 15 13 3 1 15 2 10 9 1 9 2 7 13 1 15 14 10 9 1 9 0 2
15 4 13 1 9 15 16 13 3 1 9 0 1 10 9 2
48 9 9 1 9 1 9 15 14 9 11 11 2 9 9 9 2 2 2 10 9 2 12 2 13 13 9 16 13 1 9 10 9 7 1 10 9 16 13 1 15 1 10 9 10 0 10 0 2
54 4 13 16 10 9 10 0 16 13 4 13 14 10 9 10 9 2 13 9 0 1 9 2 13 1 2 9 13 2 2 16 15 2 3 2 10 9 10 0 14 9 0 1 9 2 9 0 0 1 9 10 9 2 2
34 10 9 14 2 9 13 2 13 1 10 9 9 1 9 1 11 1 2 2 9 1 9 2 2 9 11 11 2 7 9 15 10 0 2
28 1 9 10 9 10 0 1 10 9 13 14 15 9 11 11 7 11 11 2 10 0 1 9 10 9 1 11 2
21 1 9 15 1 9 10 9 10 0 1 9 1 9 12 13 14 15 9 11 11 2
50 1 9 15 1 9 2 10 9 1 9 10 9 13 1 9 10 9 1 11 2 7 13 1 9 9 11 11 1 9 15 14 10 9 1 9 10 9 2 3 1 9 11 11 1 9 10 9 1 11 2
15 1 10 9 10 0 10 15 13 13 9 9 13 7 0 2
14 9 15 10 0 14 9 10 9 1 11 13 1 9 2
23 15 16 13 3 1 9 0 7 3 1 9 0 1 13 1 9 14 10 9 10 0 13 2
22 1 1 15 15 13 16 9 10 9 13 13 14 10 9 10 0 7 13 14 10 9 2
51 9 10 9 13 13 14 11 1 9 12 7 9 10 9 13 1 9 10 9 1 9 10 0 7 10 0 2 1 1 9 0 1 9 14 9 9 2 1 15 13 10 9 14 9 9 15 1 9 10 9 2
19 9 13 16 1 9 12 13 10 9 13 2 7 16 15 13 4 13 9 2
36 10 9 2 10 9 2 9 7 9 13 13 1 9 15 10 0 10 0 2 1 9 0 2 7 13 1 15 1 9 15 10 0 1 10 9 2
22 16 1 9 4 13 1 14 15 2 4 13 9 13 7 0 2 7 4 3 13 13 2
16 10 9 13 13 1 11 11 7 13 1 15 9 13 14 11 2
2 3 2
2 11 2
2 3 2
2 11 2
2 3 2
8 13 13 1 11 9 13 9 2
14 6 3 13 14 10 9 14 11 11 2 11 7 3 2
31 10 9 13 13 1 10 9 1 11 2 13 1 15 2 13 2 13 1 14 15 7 13 13 14 10 9 7 3 13 9 2
26 13 1 10 9 9 13 1 11 7 10 11 2 7 3 13 1 15 9 13 1 3 9 3 3 13 2
32 16 3 10 9 10 0 1 9 2 9 3 13 2 9 3 4 13 7 10 9 3 13 14 10 9 7 13 14 10 9 13 2
24 7 3 13 10 9 13 3 1 10 9 16 13 1 15 13 1 10 9 2 13 9 15 13 2
22 9 2 9 2 9 11 11 13 3 16 13 16 13 1 9 10 9 10 0 1 11 2
6 1 11 11 4 13 2
12 1 9 15 2 13 4 13 14 9 9 15 2
21 11 11 13 9 0 2 7 3 1 9 15 11 11 13 7 4 13 1 9 15 2
4 2 11 2 2
44 9 10 9 10 0 1 9 2 9 13 9 1 2 9 7 10 9 1 10 9 10 0 7 10 0 2 14 9 0 1 11 7 9 15 1 11 2 7 3 13 1 9 15 2
46 10 9 2 11 11 9 12 2 1 9 2 10 11 13 1 9 9 1 9 15 7 1 9 15 14 11 9 1 9 2 9 2 16 13 14 15 13 1 9 15 2 3 15 9 11 2
16 11 13 1 9 16 10 9 10 0 1 15 13 12 9 9 2
41 1 9 10 9 13 2 16 10 9 13 9 2 9 0 1 16 9 15 10 0 13 1 9 15 1 10 9 7 9 9 12 9 15 7 9 15 13 1 9 15 2
18 10 9 13 1 10 9 1 9 1 11 2 9 7 9 1 12 9 2
26 7 1 10 9 10 0 16 13 1 15 10 9 10 0 3 4 13 13 14 15 1 9 11 7 11 2
12 1 15 13 14 15 1 9 0 1 9 9 2
53 10 9 11 11 13 1 9 10 9 2 16 10 9 10 0 16 10 9 13 1 15 9 15 1 15 9 1 1 9 15 10 0 2 7 1 9 3 10 9 10 0 1 15 1 9 15 13 1 15 1 9 0 2
27 10 9 13 13 1 9 15 7 13 1 15 9 14 9 7 9 9 1 10 9 7 12 9 1 2 9 2
26 11 1 9 9 10 9 10 0 13 3 1 10 12 10 12 1 10 9 7 13 1 15 9 0 0 2
14 3 15 9 2 9 0 1 9 9 10 9 10 0 2
39 1 9 9 13 1 9 0 9 2 9 2 0 1 9 9 2 12 14 11 2 1 16 11 13 3 13 14 9 9 10 9 10 15 16 13 1 9 15 2
21 15 9 0 16 9 10 9 10 0 13 1 10 9 10 0 1 10 9 10 0 2
21 1 3 9 10 9 13 1 10 9 12 9 1 10 9 1 9 10 9 10 0 2
33 10 9 13 1 10 9 1 9 14 9 10 9 7 14 9 7 9 0 2 16 10 9 10 0 13 7 13 14 9 15 14 11 2
30 9 11 13 13 1 9 15 1 10 9 16 13 2 1 13 14 10 9 10 0 7 14 9 15 10 0 14 10 9 2
18 10 9 13 9 9 2 0 1 10 9 7 1 9 14 9 7 9 2
17 1 9 11 16 1 11 13 9 10 12 9 7 16 10 9 0 2
20 3 13 10 9 14 10 9 2 9 15 1 10 9 2 1 9 9 2 9 2
23 1 11 13 1 9 9 12 1 10 9 2 7 10 9 1 10 9 9 15 0 3 10 2
10 10 9 10 0 13 13 1 9 12 2
45 9 0 13 1 15 1 10 9 1 9 10 9 7 10 9 7 1 10 9 10 0 10 0 2 16 13 1 10 9 12 12 14 9 1 9 10 9 7 1 10 9 10 9 0 2
18 1 10 9 3 3 9 10 9 7 13 1 15 16 13 1 9 15 2
17 1 12 1 11 13 1 11 16 1 11 9 0 3 1 9 15 2
22 9 0 3 1 10 15 13 1 9 9 1 11 9 9 12 2 16 13 1 10 9 2
18 15 13 14 9 15 14 9 16 13 1 9 10 9 10 1 9 15 2
14 10 9 13 1 9 0 9 12 16 13 1 10 9 2
23 1 10 9 10 15 13 9 2 16 9 1 9 15 13 3 7 3 1 10 9 10 15 2
21 3 10 9 10 0 10 0 2 16 13 1 9 9 0 2 13 3 1 10 9 2
16 10 9 16 13 1 10 9 13 3 1 10 9 14 10 9 2
56 13 1 15 13 3 1 9 9 9 2 1 2 9 2 1 16 9 10 9 0 7 10 9 0 2 0 13 9 2 9 13 1 9 0 2 7 13 16 13 13 1 10 9 1 10 9 2 16 13 1 15 10 9 10 0 2
18 3 16 0 1 9 10 9 2 7 1 9 15 2 0 1 10 9 2
33 11 2 10 0 2 2 16 13 1 9 1 9 9 10 9 10 0 2 9 10 9 10 0 2 13 1 9 0 1 9 9 9 2
25 9 9 10 9 1 10 9 13 1 9 15 16 1 9 11 3 13 12 12 9 16 13 1 9 2
30 7 2 13 10 9 1 10 12 1 11 13 1 9 0 14 10 10 9 7 9 9 10 9 1 10 9 1 9 0 2
23 9 13 1 10 9 2 10 0 2 1 9 14 9 1 12 9 2 3 7 1 9 15 2
6 3 9 10 9 13 2
50 10 9 13 13 14 9 15 14 9 10 9 13 9 0 1 10 9 16 13 1 10 9 2 1 9 16 10 9 13 1 15 9 1 10 9 10 0 7 10 0 7 1 9 9 0 0 1 9 9 2
16 1 10 12 1 11 13 9 9 1 9 9 10 9 10 0 2
31 9 9 15 13 13 1 9 15 14 9 9 10 9 16 13 9 10 9 2 16 10 9 1 13 2 9 15 14 11 13 2
31 9 10 9 2 16 13 1 9 0 0 2 13 13 14 9 9 10 9 2 1 9 1 12 9 3 1 9 10 9 2 2
29 1 10 9 13 9 3 1 9 1 9 0 1 10 9 2 16 13 1 9 0 1 10 9 10 0 1 11 3 2
34 9 15 13 1 9 15 14 11 1 12 9 0 2 9 2 9 7 9 2 7 1 9 15 14 3 9 1 10 9 10 0 10 0 2
29 1 9 15 13 13 1 9 10 9 16 0 3 2 7 3 9 10 9 16 13 1 10 9 3 9 1 14 15 2
23 3 9 15 0 1 10 9 10 0 7 10 0 14 11 2 7 15 13 1 9 10 9 2
27 11 10 0 13 3 1 9 15 2 7 16 9 1 9 15 13 1 9 15 7 0 1 10 9 10 0 2
39 9 0 13 3 1 12 12 14 9 2 16 13 1 10 9 1 9 10 9 14 11 12 2 16 1 15 9 13 3 2 13 12 7 13 12 9 2 9 2
20 9 13 3 3 1 11 7 1 11 2 7 3 3 1 9 11 7 1 11 2
15 3 9 0 13 14 9 15 7 13 9 0 1 10 9 2
19 1 10 10 9 3 13 10 10 9 2 7 12 12 9 13 3 1 9 2
12 1 15 2 13 3 9 7 3 10 9 9 2
16 1 10 9 11 2 7 2 13 1 9 1 12 9 1 9 2
17 3 16 13 1 10 9 13 9 10 9 16 13 1 9 10 9 2
33 9 0 1 10 9 16 13 1 9 15 13 1 10 9 16 13 1 9 10 9 3 2 10 3 2 0 11 9 2 9 10 9 2
21 3 13 14 10 9 1 10 9 1 13 14 9 9 10 9 1 9 9 10 9 2
64 4 13 16 10 9 10 15 13 1 9 11 9 13 1 9 10 9 12 12 9 1 9 9 2 9 1 9 9 10 9 1 9 0 0 1 9 9 2 16 13 1 9 10 9 10 3 2 0 7 1 9 10 9 10 0 14 10 9 9 0 1 10 9 2
27 11 9 2 12 9 9 9 15 7 3 9 9 2 13 1 9 10 9 10 0 14 12 10 9 10 15 2
76 7 13 1 9 2 10 9 1 9 10 9 2 3 15 3 16 9 15 13 7 9 15 1 10 9 10 0 13 1 10 9 2 7 16 15 13 13 1 9 0 14 9 15 10 0 2 11 2 9 10 9 10 0 2 10 9 1 9 15 1 11 2 16 9 15 13 1 7 1 1 9 15 1 10 9 2
26 1 2 9 9 10 9 13 3 9 7 9 9 10 9 1 10 9 2 1 13 14 10 9 10 0 2
18 9 10 9 13 7 4 16 9 10 9 13 13 14 9 9 10 9 2
28 1 15 2 10 9 10 0 13 1 15 9 7 3 13 11 10 0 1 9 1 9 0 1 10 9 10 0 2
42 1 10 9 16 1 15 13 1 9 1 9 10 9 7 1 9 10 9 2 13 9 1 10 9 10 0 11 16 1 11 2 9 0 1 10 9 1 11 1 10 9 2
26 11 14 9 10 12 2 13 7 13 7 13 9 9 0 2 1 9 7 1 9 1 9 11 14 3 2
14 7 3 1 9 15 13 9 9 9 2 12 14 11 2
10 11 2 0 1 2 10 9 2 2 2
43 9 0 16 13 14 9 9 15 14 10 9 10 0 10 0 9 11 11 11 2 13 9 0 14 9 0 1 10 9 10 0 14 15 2 7 3 1 9 10 9 14 15 2
65 9 10 9 16 13 1 9 9 11 2 9 11 11 1 9 11 1 11 2 16 13 3 1 9 10 9 1 9 15 14 11 2 13 3 1 9 0 16 3 13 9 1 10 15 14 9 1 9 15 14 10 9 10 0 10 0 2 1 9 16 13 9 1 9 2
29 9 11 2 16 13 1 11 14 9 10 9 14 15 1 9 12 2 13 3 16 15 13 1 9 1 9 10 9 2
34 1 15 2 4 13 16 10 9 13 13 14 10 9 14 11 2 16 16 11 7 10 9 14 15 1 9 10 9 13 3 1 10 9 2
33 11 11 11 2 9 9 16 13 14 10 9 1 9 9 14 0 1 11 1 9 10 12 7 10 12 2 13 1 9 12 1 9 2
60 10 9 10 0 2 16 13 3 1 10 9 2 11 11 11 2 3 2 13 1 9 16 9 0 13 13 9 16 13 1 9 11 2 1 16 10 9 1 9 15 13 9 9 1 9 9 9 15 14 11 1 9 9 10 9 10 0 14 15 2
24 10 9 13 1 9 9 1 10 9 1 9 10 9 10 0 7 10 0 1 10 9 16 13 2
56 9 0 2 16 13 1 9 9 10 9 2 13 16 13 13 1 9 10 9 10 0 14 9 10 2 9 2 10 0 2 10 2 9 2 9 2 2 2 16 4 13 3 1 11 2 7 3 1 9 9 0 1 9 10 9 2
11 10 9 4 13 9 0 0 1 9 11 2
43 8 8 8 16 13 14 9 15 14 9 11 11 11 1 9 14 9 0 2 13 16 11 13 1 9 0 1 9 0 3 3 1 9 0 7 3 13 14 15 1 9 15 2
38 10 9 13 13 3 9 10 9 10 0 1 9 11 2 7 13 1 10 9 16 13 1 9 15 10 9 3 2 16 11 13 9 14 9 7 9 0 2
20 9 10 9 14 11 13 9 1 9 10 9 1 9 15 14 12 9 9 0 2
65 10 2 11 11 11 2 13 1 9 15 3 2 16 1 10 9 14 11 13 9 0 14 9 1 9 7 1 9 0 14 9 0 2 11 11 2 16 13 1 9 0 2 1 9 15 14 10 9 16 13 14 11 1 9 15 2 9 0 1 9 10 9 14 11 2
49 10 9 13 16 11 3 13 14 9 15 14 11 1 10 9 10 0 14 15 2 7 13 1 15 9 3 3 1 9 10 9 14 15 2 7 16 13 1 9 0 1 9 0 1 10 9 14 11 2
19 12 10 9 10 0 14 9 9 11 2 1 12 9 0 2 13 3 3 2
41 10 2 11 2 13 1 10 9 14 15 3 2 16 9 1 9 10 9 1 9 11 13 13 3 9 2 16 13 16 9 0 1 9 15 14 11 13 1 9 0 2
38 1 10 9 16 13 13 9 0 14 9 9 0 2 11 11 2 16 13 16 11 11 11 13 9 9 1 9 1 10 9 2 9 10 9 1 9 15 2
20 1 10 9 13 16 0 3 9 1 9 9 2 11 2 1 9 2 11 2 2
19 10 9 13 1 13 16 2 3 13 1 15 9 7 3 1 9 0 2 2
27 1 9 15 13 3 3 2 16 1 10 9 14 11 2 16 13 1 11 1 9 11 2 3 13 9 11 2
16 10 9 14 9 11 0 7 0 7 13 0 1 15 14 11 2
30 10 9 14 15 13 3 3 1 9 0 1 9 11 2 7 3 1 9 16 13 1 10 9 2 7 9 10 9 3 2
30 0 10 9 2 16 9 11 7 9 11 15 1 9 9 11 2 16 15 10 9 10 0 1 10 9 1 9 10 9 2
12 7 1 15 13 10 9 16 1 12 10 9 2
13 11 7 11 0 1 9 0 7 13 1 9 0 2
17 13 13 16 1 9 9 11 13 9 10 9 9 11 12 2 11 2
24 13 9 10 14 9 11 7 13 16 1 9 10 9 13 1 9 9 10 9 3 2 1 9 2
52 1 9 10 9 16 13 1 10 9 13 10 9 10 0 14 11 9 9 2 11 11 11 9 3 0 15 9 1 9 0 1 9 10 9 2 7 13 3 9 0 2 7 1 12 1 10 15 1 9 15 13 2
14 1 9 3 13 9 0 1 11 1 9 11 1 11 2
14 1 10 9 13 3 9 9 9 7 9 9 1 9 2
8 1 10 9 13 16 15 13 2
47 7 16 13 13 14 10 9 1 9 2 13 1 10 9 1 9 10 9 7 13 7 4 13 1 15 1 9 11 9 7 9 9 0 2 13 1 15 9 7 10 9 0 1 9 15 2 2
37 1 9 11 1 10 9 13 9 0 1 10 9 7 13 12 9 2 16 1 10 12 1 15 12 9 9 2 9 2 9 7 3 2 0 7 0 2
13 13 13 14 9 10 9 2 7 9 10 11 13 2
9 9 15 14 9 10 9 13 11 2
14 3 13 9 0 14 9 1 9 9 11 1 9 9 2
10 10 9 13 1 15 0 1 10 0 2
11 13 1 10 9 10 0 2 0 11 11 2
42 1 9 2 15 13 1 15 2 1 11 2 13 1 15 16 13 14 10 9 10 9 7 13 16 13 9 1 10 9 15 2 7 16 15 0 1 10 0 7 13 3 2
15 15 13 13 1 15 1 9 0 9 0 1 9 9 0 2
33 10 9 16 13 1 11 13 1 9 9 2 16 3 1 3 2 13 9 1 9 9 8 2 15 13 14 15 1 9 7 1 9 2
8 9 0 1 9 1 12 9 2
31 11 11 13 1 10 9 7 10 9 1 9 15 14 11 2 16 10 9 14 15 13 0 7 0 7 9 9 13 1 15 2
25 9 11 2 16 9 7 9 13 14 9 15 10 0 2 13 9 3 2 3 1 9 7 1 9 2
22 3 7 1 10 9 10 0 3 9 13 1 9 15 14 11 2 7 7 13 1 15 2
23 15 13 9 0 2 16 13 1 9 14 9 1 9 0 2 7 10 9 13 1 10 9 2
5 15 13 1 9 2
12 15 13 16 13 12 9 2 7 14 10 9 2
7 7 16 10 9 13 0 2
40 7 15 13 7 13 14 9 11 11 7 13 1 15 9 2 7 13 1 9 0 14 11 2 11 2 16 13 13 14 10 9 7 4 16 13 1 15 9 0 2
19 9 10 9 13 1 9 9 7 9 1 9 3 2 9 7 1 9 9 2
15 15 13 1 9 13 14 10 0 7 13 9 1 10 11 2
27 1 10 9 16 13 13 11 11 14 9 9 11 2 16 13 9 1 10 9 1 9 0 1 9 1 9 2
8 7 15 13 1 9 9 0 2
7 7 3 3 1 9 15 2
18 3 9 0 1 9 16 13 1 9 0 13 13 1 9 7 1 9 2
12 15 13 1 10 9 2 2 1 11 3 13 2
6 7 13 13 1 9 2
5 15 13 9 2 2
7 9 2 9 13 1 11 2
29 9 0 13 1 10 9 2 16 3 13 1 15 9 2 7 3 15 13 1 10 9 2 7 16 10 9 3 13 2
22 7 3 1 15 11 11 2 7 1 10 9 16 13 13 1 10 9 16 1 1 15 2
17 13 14 10 9 10 0 10 9 1 11 11 2 9 9 10 9 2
16 9 16 13 0 7 0 9 2 9 0 1 9 1 9 2 2
7 7 11 13 3 0 3 2
36 11 11 7 11 9 2 1 9 1 9 15 10 0 14 11 11 2 13 1 1 9 2 7 13 9 0 1 9 15 14 3 16 13 1 9 2
47 13 11 16 13 1 9 10 9 9 0 2 7 13 14 10 9 3 13 2 1 9 15 14 3 16 13 1 12 12 9 1 10 9 2 7 10 9 3 13 9 10 9 10 0 14 15 2
19 11 11 2 1 9 0 2 13 4 7 13 7 13 1 9 1 10 15 2
50 11 13 1 9 10 9 2 0 7 0 2 12 12 9 2 9 1 10 9 2 2 13 11 11 1 10 9 1 9 10 9 2 1 10 9 1 10 9 10 0 1 9 11 10 0 1 11 2 11 2
26 10 9 10 0 2 10 9 14 9 2 11 2 1 9 9 2 7 7 15 13 10 9 10 13 3 2
18 2 9 2 11 2 13 3 2 13 14 2 9 2 11 13 3 2 2
50 10 9 10 0 14 11 1 11 2 9 14 11 11 2 9 7 9 11 2 11 2 9 7 1 9 11 2 11 2 9 7 11 2 11 2 11 2 13 1 9 12 9 2 16 10 9 9 7 9 2
19 3 2 9 9 13 1 10 9 2 7 1 9 15 15 13 1 9 0 2
32 10 9 1 9 0 13 1 0 2 1 1 9 0 7 0 2 0 1 9 2 2 7 4 9 3 1 9 0 2 0 3 2
8 1 11 13 3 11 2 11 2
14 9 10 9 14 11 13 1 12 2 1 9 11 11 2
9 11 2 11 13 12 9 1 15 2
69 10 9 13 3 2 1 10 9 2 14 9 11 2 11 2 11 2 14 2 11 11 2 2 9 9 16 13 1 9 2 2 9 9 9 2 9 2 9 9 2 7 1 12 3 14 2 11 9 2 2 9 10 9 2 16 13 3 9 0 14 12 9 2 1 9 14 12 9 2
27 1 1 10 9 16 13 1 9 11 2 12 9 2 2 13 16 13 1 9 11 2 11 2 11 3 13 2
18 7 13 16 12 10 9 13 13 3 1 9 2 10 9 14 10 9 2
9 7 1 10 9 13 10 9 13 2
9 10 9 10 0 14 11 13 3 2
7 13 9 0 2 13 3 2
31 9 13 16 11 11 2 10 9 10 0 14 11 2 11 2 11 2 13 3 1 9 0 7 9 15 13 1 9 10 9 2
8 1 11 13 14 9 2 11 2
41 9 10 9 14 11 2 11 2 11 2 16 13 1 10 9 1 12 3 1 10 9 10 0 1 10 9 14 11 1 11 2 3 13 9 14 9 2 1 9 0 2
66 4 13 1 9 10 9 14 9 10 9 10 0 7 1 9 1 9 10 9 14 2 11 11 2 2 4 13 9 16 13 3 2 9 1 3 2 9 2 7 13 14 11 11 13 14 10 9 1 9 2 13 1 10 9 14 9 7 13 1 9 2 9 1 10 9 2
42 1 9 0 2 1 9 10 9 2 13 1 11 2 11 12 9 2 9 2 7 10 9 10 0 13 1 10 9 14 11 7 14 11 2 11 2 11 1 12 1 9 2
16 1 1 10 9 10 0 10 15 13 1 11 3 9 11 11 2
23 15 13 3 9 7 1 15 12 9 9 7 12 9 14 9 1 9 16 13 1 10 9 2
31 1 11 13 9 1 15 2 1 12 13 14 9 9 15 1 11 1 10 9 7 13 14 10 9 1 9 9 0 7 0 2
13 15 13 3 1 12 12 9 1 10 9 10 0 2
20 10 9 2 16 13 1 12 9 1 9 2 13 1 11 1 9 1 10 9 2
25 9 2 9 7 9 9 0 13 9 9 2 7 10 9 13 16 13 1 15 9 16 13 9 9 2
11 10 9 15 9 2 7 0 7 0 3 2
39 1 10 9 10 0 16 13 14 10 9 13 1 9 10 9 3 11 2 16 13 14 10 9 1 9 0 1 10 9 10 0 2 16 13 3 1 10 9 2
13 9 9 15 14 9 2 11 13 16 13 13 15 2
23 9 15 2 10 9 2 7 10 10 9 10 9 2 0 7 13 2 13 1 15 1 9 2
13 10 9 13 3 15 3 1 10 9 1 9 11 2
15 9 13 1 9 0 2 0 3 7 1 10 15 13 13 2
13 1 10 9 13 10 9 13 14 9 15 10 0 2
25 10 9 13 1 10 9 7 1 10 9 13 1 15 9 2 11 1 9 1 9 0 1 9 15 2
26 1 10 9 15 9 16 13 3 1 9 15 2 7 10 9 10 0 13 16 13 9 0 1 9 15 2
16 1 3 13 1 9 1 9 9 1 9 10 9 14 11 11 2
18 1 9 9 0 13 13 2 9 2 1 9 15 14 9 0 2 0 2
52 13 1 10 9 14 9 0 1 10 9 3 9 0 2 15 13 14 10 9 1 12 9 2 9 9 7 9 2 16 7 13 1 15 9 13 1 10 15 13 13 13 1 10 9 1 9 16 13 1 15 9 2
18 7 3 3 15 2 7 16 1 10 9 10 0 13 3 9 13 9 2
39 9 15 13 1 9 0 9 0 7 13 14 9 10 9 2 7 3 3 9 14 9 9 1 9 15 10 0 9 2 9 2 9 2 9 2 9 7 3 2
20 13 1 11 9 1 10 3 16 13 1 11 2 11 2 11 2 7 7 3 2
24 12 9 0 1 9 13 11 1 9 1 11 2 9 16 13 1 15 14 11 2 11 2 11 2
36 1 11 9 9 12 9 1 9 9 9 2 7 15 13 14 15 1 10 9 16 13 3 1 9 9 2 1 9 0 2 7 13 9 14 3 2
40 13 1 10 9 9 9 2 7 1 15 2 13 10 13 2 13 10 9 1 10 9 2 1 9 0 2 7 10 9 13 14 15 1 9 15 7 1 9 15 2
15 9 11 1 9 2 10 9 16 1 11 3 13 3 0 2
40 1 2 11 11 2 7 10 9 16 13 1 9 1 10 9 14 11 2 11 2 11 2 13 1 11 14 11 11 2 2 13 10 9 7 14 2 9 9 2 2
9 9 0 7 3 2 0 3 3 2
40 1 16 11 11 13 14 10 9 1 9 10 9 14 2 9 10 9 2 2 15 13 9 0 1 10 9 7 13 14 15 1 9 16 1 15 13 9 14 9 2
35 1 9 7 1 9 0 1 9 10 9 2 3 15 13 14 10 9 13 14 9 10 9 2 1 1 9 10 9 10 0 16 1 10 9 2
14 13 14 9 10 9 7 13 14 15 1 1 9 0 2
16 12 10 9 13 14 9 10 9 1 10 9 2 1 9 15 2
27 1 9 10 9 13 1 9 7 13 1 1 10 9 1 9 10 9 2 12 1 9 11 2 16 13 3 2
29 10 9 13 3 13 14 9 10 9 2 12 9 1 10 12 9 2 2 16 13 13 14 10 9 7 14 10 9 2
16 10 9 16 13 1 9 10 9 13 9 0 1 9 10 9 2
34 1 9 10 9 10 9 4 13 7 10 2 9 2 13 2 2 9 2 3 2 15 13 2 13 3 14 2 1 9 1 10 9 2 2
18 13 3 9 16 1 15 13 9 2 9 1 10 9 7 1 10 9 2
28 3 1 11 7 3 1 11 2 11 2 11 10 9 9 0 1 10 9 7 13 1 10 9 1 9 9 0 2
11 7 1 12 10 9 13 9 1 10 9 2
20 10 9 13 1 9 14 9 9 0 2 7 7 9 10 9 13 1 9 9 2
8 10 9 13 1 9 0 3 2
70 9 11 1 10 9 14 10 9 2 1 2 11 11 2 2 13 9 16 13 1 11 11 2 16 13 1 15 9 9 1 2 11 2 2 2 9 2 7 3 2 9 1 10 9 14 2 9 2 15 13 2 2 1 11 11 2 1 9 15 14 11 11 2 7 2 9 10 9 2 2
54 4 13 1 9 15 10 0 14 11 11 2 16 13 0 3 1 9 9 10 9 1 9 10 9 14 11 2 11 2 11 2 7 4 3 13 14 10 9 14 9 10 9 1 10 9 2 7 13 1 11 9 3 0 2
17 12 9 9 0 13 1 10 9 1 12 2 11 11 7 9 11 2
33 10 9 16 9 15 2 11 2 11 2 13 14 10 9 1 9 1 9 9 15 14 9 13 1 11 7 11 2 9 11 7 0 2
15 10 9 10 0 7 10 0 13 9 13 1 9 7 9 2
25 4 13 7 15 9 16 13 1 9 9 2 7 9 9 16 13 14 10 9 10 0 1 9 9 2
22 3 7 3 2 15 9 1 9 10 9 10 0 14 10 13 1 11 2 11 2 11 2
22 9 8 14 10 13 1 10 9 4 13 1 9 0 3 7 9 7 9 1 9 0 2
15 10 9 1 12 10 9 7 13 1 9 0 14 10 9 2
24 1 11 2 11 2 11 13 1 11 14 10 10 12 2 1 11 1 9 10 12 7 10 12 2
16 1 12 10 9 13 9 11 2 7 10 9 7 10 0 0 2
22 1 11 13 11 11 2 9 0 2 13 1 10 9 7 10 9 0 1 13 2 0 2
20 9 10 9 0 2 7 1 10 9 13 9 14 11 2 11 7 11 2 11 2
20 1 12 10 9 10 9 13 9 9 7 9 2 10 12 9 9 1 14 15 2
34 1 11 2 11 2 11 13 14 2 9 11 9 2 2 16 1 15 13 14 10 9 2 11 2 2 10 9 10 0 1 9 10 9 2
27 15 13 1 10 13 16 13 1 2 11 2 7 3 13 3 2 7 13 9 1 3 16 13 14 10 9 2
27 1 15 2 10 2 11 9 9 2 1 11 2 10 0 3 1 10 9 2 0 1 9 9 7 13 0 2
6 3 13 1 9 9 2
17 3 9 9 0 2 0 2 1 11 2 13 1 10 9 10 9 2
16 3 13 3 9 0 1 9 15 1 9 15 7 1 9 15 2
5 3 9 13 3 2
14 10 9 10 0 14 11 1 9 15 13 9 9 0 2
22 9 14 12 9 2 9 13 1 9 0 2 7 10 9 13 14 9 10 9 1 9 2
19 1 10 16 13 1 9 10 9 7 10 9 2 13 1 11 10 3 13 2
21 1 11 2 11 2 11 13 12 1 10 9 1 9 2 1 9 0 7 1 9 2
23 15 10 9 10 0 13 1 12 10 9 1 9 13 14 10 10 9 10 0 1 10 9 2
27 1 11 9 13 14 10 9 1 10 9 10 0 2 1 16 10 9 13 0 1 1 11 2 11 2 11 2
28 9 13 1 10 9 7 4 13 15 13 1 10 9 10 0 2 13 1 10 9 10 0 2 7 10 9 13 2
15 13 9 16 10 10 9 3 0 3 1 10 9 10 0 2
27 9 0 2 16 13 1 9 9 12 1 12 9 2 3 13 9 15 7 9 15 1 9 9 14 10 9 2
28 3 7 13 16 10 9 10 0 14 11 2 11 2 11 13 1 10 9 1 9 15 2 15 3 13 13 9 2
9 1 12 13 3 12 9 9 0 2
48 2 9 10 9 2 2 16 13 1 10 9 14 11 11 2 13 1 9 9 2 13 1 15 9 2 9 2 9 9 7 9 2 9 3 9 0 2 7 9 1 9 9 10 12 7 10 12 2
36 10 9 10 0 2 16 13 1 9 12 9 2 13 3 7 15 10 2 11 1 11 2 9 9 2 1 9 7 1 9 2 9 0 7 9 2
32 1 9 10 9 14 11 2 11 9 0 2 7 13 1 10 9 10 0 10 0 16 3 13 1 9 15 2 15 13 0 3 2
27 11 13 4 13 1 9 9 10 9 16 1 11 2 11 2 9 0 1 9 10 9 1 10 9 10 0 2
27 1 11 3 13 3 12 9 9 2 2 9 10 9 2 2 12 9 2 7 2 11 2 2 12 9 2 2
16 1 9 11 13 9 12 2 9 10 9 2 2 12 9 2 2
26 1 9 10 9 10 15 4 13 3 1 10 9 14 11 2 11 1 9 0 0 7 1 9 2 9 2
32 1 12 13 13 1 11 2 11 3 12 9 9 2 1 12 9 2 2 9 1 9 9 2 9 9 2 9 7 3 9 9 2
24 10 9 1 11 13 1 10 9 14 11 7 1 12 9 10 9 7 10 9 16 1 10 9 2
10 11 2 0 1 2 10 9 2 2 2
38 1 10 9 10 0 13 9 0 16 13 13 14 11 11 1 10 9 1 11 11 2 1 10 9 10 0 1 10 9 2 16 13 1 10 12 1 11 2
46 9 16 13 1 11 13 16 15 13 1 9 10 9 2 11 11 2 14 9 15 1 9 14 2 9 9 2 2 9 16 13 1 15 1 13 1 3 13 14 10 9 7 10 9 13 2
24 10 9 10 0 13 15 13 1 9 13 1 10 9 1 9 10 9 1 10 9 1 12 9 2
39 1 11 2 9 0 16 1 15 9 0 0 2 13 9 15 14 10 9 1 12 9 1 10 9 1 9 12 2 16 10 9 13 1 9 15 1 10 9 2
15 10 9 13 1 9 12 1 10 9 7 10 9 10 0 2
36 1 10 9 11 2 16 13 3 7 3 9 14 10 9 2 13 10 9 14 10 9 14 15 1 9 10 9 2 14 15 13 3 1 12 9 2
36 13 16 9 10 9 1 9 10 9 0 1 15 16 1 10 9 10 0 2 16 1 15 13 1 9 2 9 3 9 1 12 10 9 10 0 2
36 9 9 10 9 13 9 14 10 9 10 0 1 9 1 10 9 10 0 2 1 9 1 10 9 2 1 9 10 9 7 1 9 9 10 9 2
16 1 15 13 3 9 2 9 0 2 16 13 0 1 9 9 2
26 1 9 10 9 10 0 13 9 2 7 9 15 14 9 10 9 1 9 9 0 1 10 9 10 0 2
15 1 9 15 13 1 9 15 9 9 10 9 13 11 11 2
27 13 14 9 2 10 9 1 9 10 9 1 9 2 10 9 7 13 1 9 1 9 2 11 2 1 11 2
15 1 10 9 15 13 9 3 0 2 13 1 9 9 0 2
20 10 9 0 9 9 7 13 1 9 0 2 16 13 1 10 9 1 9 0 2
20 11 13 14 10 9 1 9 11 7 13 14 10 10 9 10 0 1 9 12 2
17 14 10 9 13 11 1 9 9 2 7 13 9 1 9 9 0 2
23 3 13 11 14 9 9 15 1 9 1 9 9 2 2 9 2 13 1 9 9 7 9 2
28 10 9 13 1 9 2 9 2 9 2 9 7 3 9 0 16 13 14 15 2 7 9 15 13 9 14 11 2
18 15 13 1 2 9 9 10 9 2 1 9 16 11 15 13 7 13 2
18 4 13 14 10 9 1 10 9 1 9 9 1 9 2 9 1 12 2
12 11 11 13 7 13 9 9 0 1 9 0 2
19 10 9 16 15 13 1 15 13 9 1 11 2 16 13 2 9 10 9 2
29 1 13 14 10 9 2 16 0 9 1 9 0 2 13 14 15 11 1 9 9 7 13 14 15 1 9 9 9 2
33 1 1 3 15 13 14 10 9 1 9 10 2 9 2 9 2 9 2 9 2 9 2 9 9 2 9 9 2 9 0 7 3 2
29 1 10 9 2 10 3 16 1 9 15 13 9 10 9 2 16 4 3 1 9 1 10 9 2 2 3 13 9 2
16 10 9 13 1 9 15 3 9 2 1 9 1 9 10 9 2
31 10 9 2 1 9 12 9 7 1 12 9 2 13 1 12 9 1 10 9 10 0 7 1 12 9 1 10 9 10 0 2
4 9 2 12 2
9 11 11 13 9 0 1 9 9 2
18 1 9 11 0 15 13 1 15 11 2 11 2 11 0 1 9 0 2
34 9 10 9 2 9 2 11 13 1 10 10 9 7 1 10 10 9 2 7 1 15 9 0 14 9 2 9 2 9 7 9 0 0 2
39 1 9 0 14 10 9 10 0 9 2 9 2 9 0 1 9 13 7 3 2 13 11 14 9 10 11 2 11 2 11 7 13 14 15 1 9 10 11 2
16 1 9 10 9 15 13 9 1 9 9 1 13 14 10 9 2
17 4 13 14 10 9 1 9 9 0 3 1 9 16 10 9 13 2
11 9 10 9 12 9 2 0 1 9 15 2
4 9 2 12 2
11 11 2 11 2 11 13 9 1 9 13 2
12 15 13 3 1 9 2 9 7 9 0 3 2
18 10 9 16 13 1 9 10 9 13 1 10 9 10 0 14 10 9 2
19 11 13 14 9 10 9 2 13 14 15 2 7 1 9 10 9 3 13 2
18 15 13 3 1 9 9 2 16 14 15 15 13 1 9 14 9 9 2
12 1 10 9 13 11 9 16 13 1 9 0 2
63 10 9 2 11 2 11 2 1 9 9 7 0 2 11 2 9 0 16 1 9 15 4 13 1 15 9 2 7 9 2 11 2 2 16 1 9 15 13 1 12 9 2 0 1 10 9 10 0 2 1 10 9 10 12 9 0 7 1 10 9 0 0 2
10 1 9 15 13 11 3 9 7 9 2
15 10 9 2 9 12 9 2 9 12 9 7 9 12 9 2
4 9 2 12 2
10 16 13 7 13 1 12 12 9 3 2
28 3 13 9 9 9 11 11 11 2 11 1 9 9 1 10 9 10 0 10 0 1 9 10 9 14 10 9 2
19 9 10 9 10 0 1 11 9 0 7 9 3 3 13 1 12 12 9 2
27 11 2 11 13 16 10 9 1 10 9 10 0 13 0 1 9 14 12 12 9 2 16 13 1 10 9 2
36 10 9 1 10 9 13 3 1 1 9 10 9 1 2 9 9 10 9 2 16 13 12 12 9 1 10 9 2 7 10 9 10 0 10 0 2
30 9 10 9 1 10 9 10 0 13 1 10 9 1 9 10 9 7 10 9 16 1 9 0 13 1 15 9 0 3 2
50 11 2 11 2 16 13 3 1 13 9 10 9 7 10 9 1 9 10 9 2 13 16 9 10 9 1 10 9 10 0 16 15 3 13 7 13 12 9 1 9 10 9 13 1 10 9 12 12 9 2
15 15 13 16 13 1 10 9 9 0 1 9 9 9 15 2
20 1 9 10 9 1 9 12 13 16 1 9 10 9 13 9 14 12 12 9 2
21 11 2 11 13 16 9 15 0 7 9 15 13 1 10 9 10 0 16 13 3 2
25 1 10 9 10 0 3 13 9 0 1 2 9 9 15 7 15 13 1 10 9 10 0 10 0 2
28 10 9 1 11 13 7 10 9 10 0 7 10 9 16 13 3 3 13 9 0 1 9 10 9 7 10 9 2
17 10 9 10 13 14 9 11 1 9 12 13 1 3 12 12 9 2
36 9 9 10 9 13 16 15 9 1 9 0 3 1 10 9 10 0 10 0 2 7 15 9 14 9 0 0 7 9 9 1 10 9 10 0 2
43 1 15 2 10 9 1 10 9 13 3 1 10 9 16 13 1 10 9 7 10 9 13 1 10 9 13 14 10 9 16 13 1 10 9 1 9 1 9 15 1 9 11 2
26 3 16 1 9 15 9 9 2 13 7 13 2 13 9 9 2 9 10 9 1 9 13 10 0 3 2
13 1 15 2 10 9 1 9 9 13 10 0 3 2
21 15 13 1 9 9 9 16 13 10 9 1 9 10 9 1 10 9 1 10 9 2
43 3 9 10 9 1 10 12 9 2 9 9 9 9 14 9 9 2 2 9 12 9 9 2 9 2 1 12 9 9 2 1 9 2 12 9 9 12 9 9 1 9 12 2
37 12 11 16 13 13 9 9 0 13 9 1 9 9 10 9 1 9 15 16 13 10 9 2 9 9 1 12 1 12 9 2 0 1 9 10 9 2
8 9 0 1 12 1 12 9 2
7 9 1 12 1 12 9 2
14 9 9 0 1 12 1 12 9 2 0 1 10 9 2
8 13 9 1 12 1 12 9 2
52 9 10 9 1 9 10 9 13 2 16 1 9 1 10 9 16 13 2 10 9 10 9 13 1 9 0 1 9 9 10 9 2 7 16 3 13 3 2 1 15 2 1 9 0 13 9 9 14 1 12 9 2
11 13 9 16 4 13 9 9 1 10 9 2
13 10 9 1 9 0 3 2 0 3 7 0 3 2
33 10 9 1 9 0 3 2 7 16 15 13 14 10 9 1 10 9 7 13 9 0 2 2 2 1 15 10 9 4 13 9 0 2
35 9 9 2 1 9 2 4 3 15 2 3 2 13 0 2 16 16 15 13 14 9 10 9 7 13 14 10 9 2 7 7 0 9 9 2
14 16 13 1 9 7 1 9 2 4 3 13 9 9 2
22 3 4 1 10 9 13 1 9 9 7 9 1 10 9 2 7 3 3 1 9 9 2
32 9 10 9 16 13 3 1 9 9 13 9 0 2 16 13 13 14 10 9 7 16 13 9 9 3 7 10 9 13 1 15 2
22 2 11 13 3 0 1 9 10 9 2 15 13 13 14 15 1 9 9 3 2 0 2
16 7 13 1 9 9 10 9 10 0 7 1 9 9 9 9 2
12 15 13 2 16 10 9 16 13 1 15 13 2
19 11 13 3 10 9 14 15 2 16 16 10 11 16 1 9 15 3 0 2
62 15 13 1 15 10 3 3 2 2 3 13 1 9 2 7 1 10 9 10 0 2 10 9 11 2 1 9 15 2 11 11 0 2 9 9 10 9 14 9 9 10 9 2 16 13 3 1 9 9 1 9 10 11 2 1 9 10 9 1 9 9 2
34 11 13 1 9 9 1 9 10 9 16 13 1 11 2 9 9 3 1 16 13 1 11 1 10 9 10 0 14 9 9 9 10 9 2
42 9 0 13 14 11 11 1 9 15 10 0 2 1 15 9 7 9 3 2 9 11 2 9 9 2 9 12 10 9 10 3 2 0 14 9 9 9 7 9 10 9 2
31 1 10 9 10 0 13 1 15 9 10 9 2 11 11 2 16 13 1 9 15 10 0 14 11 11 7 9 15 10 0 2
22 3 1 10 15 13 9 15 14 11 1 9 0 14 9 11 2 9 1 11 2 11 2
17 0 1 9 9 9 10 9 13 10 9 1 9 10 9 16 13 2
13 2 11 2 13 15 1 15 0 2 0 7 13 2
12 3 10 9 13 14 9 15 1 9 3 9 2
31 10 9 13 1 15 2 3 1 3 16 1 9 9 13 1 9 10 9 2 3 1 9 15 10 0 1 9 9 10 9 2
47 3 15 13 1 15 13 9 0 1 10 9 1 10 9 16 13 13 10 9 9 12 2 2 13 1 9 13 9 9 9 10 9 2 11 11 2 1 10 9 2 1 9 1 9 10 9 2
9 2 9 9 9 10 9 13 9 2
16 13 14 9 15 14 12 1 9 10 9 2 9 9 7 9 2
8 9 9 1 9 15 10 0 2
6 13 13 1 10 9 2
5 14 16 13 13 2
10 9 15 7 9 15 13 1 15 3 2
26 13 1 9 7 13 9 9 7 15 13 13 7 13 1 9 2 2 13 9 9 10 9 2 11 11 2
22 9 10 9 2 13 7 13 2 2 13 13 14 15 2 13 14 15 7 13 14 15 2
9 11 13 9 0 2 0 7 0 2
26 1 9 9 15 10 0 2 13 1 15 3 9 7 3 9 7 15 13 1 15 3 1 9 15 2 2
22 2 13 1 9 15 9 3 2 0 1 9 10 9 1 9 16 3 13 1 9 15 2
28 10 9 1 10 9 0 3 7 7 1 10 9 2 16 13 9 0 7 9 0 1 9 15 2 2 13 11 2
19 9 10 9 16 13 1 9 10 9 14 9 10 9 13 13 14 9 15 2
81 10 9 7 9 10 9 13 1 9 0 0 7 0 2 13 2 2 7 3 10 9 13 13 1 10 9 3 13 1 1 10 9 2 1 10 13 9 10 9 7 10 9 1 10 9 16 10 9 4 13 2 15 9 10 9 16 13 1 15 2 1 10 9 14 9 10 9 1 9 10 9 13 7 15 9 10 9 14 10 9 2
41 16 2 1 9 2 9 13 1 10 9 16 9 0 0 3 1 15 16 0 9 9 0 2 4 1 10 9 13 7 15 0 3 1 10 9 2 7 1 10 9 2
15 1 10 12 1 10 9 16 0 1 10 9 9 7 9 2
14 16 16 10 9 0 3 1 9 2 3 13 9 15 2
38 7 13 9 16 13 13 1 9 15 14 10 9 10 0 2 1 16 4 13 1 12 10 9 2 3 9 0 1 10 9 2 7 3 0 1 10 9 2
26 10 9 10 15 0 1 10 9 10 0 2 7 1 1 10 9 10 0 4 3 16 13 1 10 9 2
17 4 13 1 10 9 16 1 9 10 9 1 15 16 1 10 9 2
34 7 1 10 9 10 0 2 1 9 15 10 0 14 10 9 10 9 0 9 2 3 16 13 3 9 2 13 9 2 7 9 13 9 2
23 10 9 10 0 4 13 9 2 7 0 1 9 1 9 0 7 13 11 2 11 2 11 2
12 9 16 13 13 13 2 3 4 9 7 9 2
35 11 11 11 2 9 9 9 7 9 15 1 10 9 1 9 1 9 10 9 2 13 16 1 15 13 9 2 1 9 16 15 1 9 0 2
24 1 9 15 2 10 9 10 0 2 16 13 1 9 10 9 2 13 1 9 1 10 0 3 2
15 16 1 0 2 3 15 4 13 9 2 7 16 13 13 2
20 7 15 13 2 16 1 10 9 13 3 10 9 9 16 0 1 9 0 3 2
9 1 3 13 9 0 1 9 0 2
9 10 9 0 1 9 2 9 2 2
12 9 9 10 9 13 9 9 14 9 10 9 2
19 10 9 0 1 9 10 9 7 9 15 2 16 9 15 1 11 10 0 2
24 15 9 0 2 3 1 10 9 1 9 10 9 2 7 7 13 14 15 1 9 1 9 0 2
17 10 9 13 15 1 15 2 7 10 9 13 1 9 9 7 9 2
13 10 10 9 1 10 9 13 1 10 9 10 0 2
20 10 9 16 13 1 10 9 13 9 1 9 2 16 13 14 15 1 9 9 2
20 10 9 0 1 9 9 9 2 3 9 0 7 9 9 16 3 13 1 9 2
33 1 9 9 13 9 10 9 13 1 10 9 10 0 14 10 9 16 13 1 15 3 2 9 2 9 2 9 0 7 1 0 2 2
16 14 10 9 13 3 1 9 0 7 1 3 16 13 13 9 2
21 9 10 9 13 9 14 9 10 9 1 15 13 2 9 10 9 7 9 10 9 2
39 10 9 13 4 13 14 9 10 9 16 1 1 10 9 2 7 3 3 13 1 15 7 13 1 9 10 9 2 7 13 9 1 10 9 7 1 10 9 2
57 9 1 9 0 13 1 10 9 1 9 1 9 2 7 16 15 9 2 0 2 2 15 0 7 13 13 1 9 0 1 9 10 9 2 10 9 2 1 3 10 9 10 0 2 13 9 2 0 2 2 16 4 13 9 0 2 2
21 10 9 3 0 3 1 9 2 7 10 9 4 13 1 9 0 3 14 10 9 2
14 1 15 9 15 0 1 9 0 1 15 14 10 9 2
18 9 10 9 1 12 10 9 4 13 1 12 9 1 10 9 10 0 2
19 10 9 13 9 0 3 7 0 3 1 9 2 9 7 10 9 10 9 2
46 9 1 9 15 4 13 1 10 9 2 16 16 10 9 13 1 9 2 9 1 9 9 2 9 0 7 0 3 1 10 11 7 9 15 2 16 13 1 15 1 9 9 14 10 9 2
16 10 9 10 0 2 1 9 9 10 9 2 13 1 10 9 2
53 9 13 2 1 1 9 7 1 9 2 3 1 9 2 9 14 9 1 9 0 2 2 1 2 9 0 2 16 13 1 9 14 9 0 7 9 1 9 2 2 1 9 9 0 2 7 3 0 3 1 9 9 2
14 11 11 13 2 16 9 9 4 16 13 0 7 0 2
28 0 2 16 16 15 13 7 13 9 0 1 9 10 9 2 0 2 16 16 3 15 13 3 9 1 10 9 2
65 1 9 10 9 2 3 9 10 9 10 0 1 9 2 9 12 9 9 12 9 9 12 9 12 9 9 12 9 2 1 12 9 9 2 9 12 9 2 1 12 9 9 2 2 9 2 1 2 9 9 2 9 10 9 10 0 1 9 0 13 12 9 12 9 2
20 16 16 10 9 10 0 0 3 2 3 9 15 1 9 2 3 2 0 3 2
36 2 1 10 9 13 16 10 9 2 10 9 7 10 9 13 9 10 9 10 0 3 2 7 1 9 15 13 1 15 9 1 10 9 10 0 2
19 1 10 9 4 13 2 16 9 15 16 15 13 9 0 2 3 1 9 2
29 13 9 9 16 13 9 1 9 2 9 14 9 1 9 0 1 9 9 2 1 15 9 16 0 1 15 10 9 2
20 10 2 9 2 13 1 12 9 9 0 2 16 10 9 1 15 1 12 9 2
20 9 9 10 9 13 2 16 9 15 13 13 9 2 16 16 4 13 1 9 2
28 15 16 16 10 9 10 0 13 1 15 1 9 9 0 2 7 3 1 9 10 9 13 1 9 9 10 9 2
27 1 9 0 2 9 10 9 13 16 3 4 13 3 9 13 1 10 9 2 9 0 1 10 9 10 0 2
25 11 11 13 2 16 10 9 10 0 16 13 1 9 10 9 13 9 14 9 3 0 14 10 9 2
26 1 9 15 2 9 0 3 2 1 9 0 7 1 9 9 0 14 10 9 2 13 9 1 10 9 2
12 10 2 13 9 15 2 13 10 9 10 0 2
22 9 15 13 1 9 0 14 9 0 2 9 1 9 7 9 3 14 10 9 1 9 2
26 9 10 9 13 1 9 10 9 10 13 7 1 9 10 9 2 7 2 9 10 9 7 9 10 9 2
28 13 10 9 16 10 9 13 1 9 2 0 10 1 9 2 3 15 13 9 7 13 2 7 7 15 4 13 2
29 9 10 9 0 3 3 1 10 9 10 0 7 1 10 9 2 7 15 13 13 1 10 9 10 0 1 16 13 2
26 10 2 1 10 9 2 13 9 2 0 2 7 0 1 10 9 9 16 13 1 10 9 1 9 15 2
21 11 11 13 2 16 1 9 0 2 13 1 9 0 2 3 1 9 15 10 0 2
46 9 15 10 0 14 10 2 1 9 10 9 2 13 1 15 2 16 13 1 9 15 1 9 9 16 3 4 13 15 8 2 1 9 0 7 0 2 9 9 0 2 9 2 7 3 2
14 9 9 10 9 14 15 1 9 1 15 14 9 9 2
31 1 10 9 10 0 10 9 13 3 3 12 7 3 1 15 14 9 1 9 9 2 1 9 0 3 7 9 9 0 3 2
21 10 13 13 1 10 9 7 1 9 10 9 15 13 1 2 9 10 9 10 0 2
25 10 9 0 3 13 1 10 9 7 13 9 9 0 2 1 16 13 16 1 10 9 13 9 0 2
24 3 2 13 10 1 9 10 9 1 9 10 9 7 10 9 1 9 3 13 9 1 10 15 2
55 10 9 10 0 13 9 0 3 2 7 1 9 10 9 13 10 9 10 0 2 10 9 13 9 0 12 9 12 9 9 1 9 10 9 2 1 10 9 4 13 1 9 1 9 10 9 2 7 4 13 1 9 1 9 2
32 8 13 1 10 9 2 9 1 9 15 2 3 10 9 2 2 9 1 9 15 2 11 2 11 2 11 9 2 9 7 9 2
16 9 15 14 9 13 3 12 1 9 10 9 2 13 11 11 2
39 9 13 9 0 3 2 7 9 10 9 16 15 13 13 3 1 9 15 2 7 3 1 9 10 9 14 10 9 10 0 1 9 2 9 2 9 7 3 2
34 9 15 14 10 9 10 0 13 1 12 1 12 9 1 9 2 9 10 9 10 0 3 2 16 13 11 2 13 1 12 9 1 9 2
18 11 2 9 0 16 13 1 9 13 2 0 1 12 9 1 10 11 2
19 9 11 2 11 2 16 13 7 15 1 9 0 2 0 3 3 1 11 2
9 9 15 4 13 1 9 0 0 2
42 10 9 4 13 7 13 9 0 1 9 0 3 2 7 14 10 9 10 0 2 16 13 9 0 16 13 9 1 9 2 9 7 3 7 13 9 16 4 13 14 15 2
34 11 11 2 9 9 11 2 13 16 4 13 3 9 0 2 16 13 1 9 1 9 7 9 2 1 9 10 9 16 13 1 10 9 2
11 13 9 16 13 9 0 15 1 9 15 2
50 1 15 15 13 1 3 16 13 9 9 1 9 0 14 9 2 3 13 1 9 0 15 7 13 16 3 10 9 2 10 9 7 10 10 9 10 0 2 16 13 1 9 1 9 7 9 2 13 9 2
21 9 2 1 10 9 0 9 9 0 9 16 13 14 10 9 10 0 2 11 2 2
45 9 15 13 13 7 1 10 9 10 0 14 9 1 9 9 2 9 7 9 2 7 3 10 16 15 1 9 1 9 2 7 4 13 1 13 1 9 15 10 0 2 13 11 11 2
33 7 16 1 10 9 13 12 9 2 0 16 1 9 10 9 2 1 3 1 9 10 9 2 13 9 0 1 9 10 9 16 13 2
60 1 9 2 10 9 1 9 9 1 9 10 9 13 3 1 9 15 2 16 16 9 15 13 13 1 9 9 2 16 16 13 1 10 9 2 10 9 1 10 9 1 10 9 4 9 9 7 9 2 7 1 9 9 9 2 0 7 9 2 2
15 1 10 9 10 0 13 14 9 10 9 7 9 2 9 2
18 1 9 11 2 9 9 10 9 13 12 10 9 1 9 9 10 9 2
24 1 3 13 1 15 3 9 11 2 11 7 11 2 7 1 9 9 0 13 9 11 7 11 2
20 7 1 10 9 2 9 15 13 1 9 10 9 7 1 9 15 1 9 9 2
25 10 9 13 4 13 9 15 1 9 10 9 2 7 1 9 10 9 13 16 13 3 3 14 15 2
13 3 9 0 16 13 1 10 9 13 9 10 9 2
52 13 14 9 10 9 14 15 1 9 7 14 9 2 16 13 1 9 2 10 9 1 10 9 13 12 12 9 1 9 7 9 0 2 1 9 0 2 7 3 12 12 9 9 2 1 9 1 9 14 12 9 2
33 9 10 9 13 3 14 9 10 9 1 10 9 2 9 1 9 2 1 13 2 1 9 0 2 1 9 2 1 9 7 1 9 2
55 9 2 9 11 2 2 1 9 9 2 9 2 16 13 1 9 9 1 9 7 9 2 13 3 1 9 0 2 9 9 10 9 10 0 1 2 9 9 10 9 3 2 1 12 9 1 9 15 14 9 0 1 15 9 2
32 7 16 10 9 15 16 13 1 10 9 14 9 15 2 7 15 3 10 0 3 1 9 2 13 1 9 15 1 13 9 0 2
48 10 9 10 0 0 1 2 1 9 0 2 7 1 9 9 2 14 9 10 2 13 10 9 1 10 9 0 2 1 10 10 9 16 13 1 10 9 2 7 9 9 4 13 1 12 9 3 2
20 10 9 13 14 9 9 10 9 1 9 2 7 4 13 2 1 9 0 2 2
14 9 10 2 1 9 10 9 13 1 10 9 16 13 2
29 15 9 8 8 1 11 2 11 2 11 2 1 10 9 16 1 15 10 9 13 1 9 9 2 9 7 9 0 2
20 10 9 3 13 1 9 1 9 0 2 9 12 9 2 9 1 12 9 2 2
27 10 9 13 9 2 1 9 1 13 2 9 12 9 9 12 9 9 12 9 9 12 9 1 9 9 0 2
45 12 9 9 12 9 9 12 9 1 9 0 9 9 15 14 9 9 12 9 2 1 12 9 2 1 9 13 1 2 12 9 2 1 10 9 16 13 1 9 9 0 7 9 0 2
4 2 11 2 2
35 1 9 10 9 10 0 1 9 2 9 13 1 9 11 9 9 1 11 11 2 9 12 1 11 2 16 13 1 2 9 1 10 9 2 2
23 9 10 9 2 16 13 1 9 12 9 2 13 1 11 12 9 14 9 9 1 9 0 2
43 10 9 2 9 11 11 2 13 16 1 1 9 7 9 13 11 9 0 14 9 9 1 9 9 2 1 16 15 13 1 9 7 13 1 15 1 9 10 9 7 9 15 2
32 1 9 1 10 9 2 13 1 9 10 9 2 7 13 11 1 9 1 13 14 9 10 9 7 1 13 1 10 9 1 9 2
14 9 9 10 9 14 11 13 1 3 1 12 12 9 2
36 1 9 16 13 1 2 9 9 10 9 15 13 1 10 9 1 9 2 1 15 13 1 9 9 10 9 10 9 2 7 13 3 1 9 0 2
49 1 9 10 9 13 3 2 16 1 9 10 9 1 9 11 1 9 2 9 2 13 10 9 1 9 10 9 2 16 9 15 10 0 0 1 10 9 2 7 13 13 14 15 1 9 9 10 9 2
46 8 8 8 10 9 10 0 1 11 13 10 9 1 10 9 1 10 9 16 9 10 9 13 1 9 15 2 7 3 13 11 1 10 9 9 1 9 14 10 9 7 13 1 10 9 2
24 3 1 9 11 1 9 2 9 13 10 9 2 1 13 1 12 9 2 9 9 14 10 9 2
48 1 9 9 10 9 1 9 9 1 9 2 9 13 11 2 1 13 1 12 9 1 9 10 9 2 3 9 14 12 9 1 12 1 9 10 9 2 16 13 1 10 9 14 10 9 16 13 2
44 1 9 10 9 1 10 9 10 0 1 11 2 13 1 10 9 12 10 9 16 13 1 10 9 1 9 10 9 3 13 1 10 9 14 10 9 2 7 16 13 1 9 9 2
11 15 13 1 11 1 9 13 1 15 13 2
16 1 9 13 11 9 12 1 10 9 7 10 9 13 13 3 2
27 1 9 10 9 1 9 9 10 9 1 11 2 13 9 10 9 1 10 9 10 0 1 15 13 10 9 2
19 10 9 13 1 15 14 10 9 7 13 1 15 13 1 10 9 10 12 2
15 10 9 13 1 9 15 7 13 16 16 11 13 1 15 2
25 1 9 10 9 1 9 9 0 2 0 1 9 11 1 11 2 13 1 10 9 9 14 10 9 2
22 11 13 1 15 13 3 1 9 10 9 7 13 1 15 2 2 15 13 1 15 2 2
36 7 13 14 9 9 15 2 13 11 9 12 16 13 1 9 9 1 10 9 2 16 9 15 13 1 10 9 7 13 14 10 13 1 10 9 2
27 1 9 1 9 10 9 1 9 2 9 1 11 2 13 12 10 9 13 1 9 10 9 13 1 10 9 2
17 11 13 1 15 7 13 1 15 1 9 15 13 1 9 10 9 2
24 10 9 13 7 3 1 16 10 9 13 1 9 15 2 13 10 9 7 13 1 9 10 9 2
38 11 3 13 1 9 14 12 9 1 9 9 9 10 9 1 9 2 9 2 7 13 1 10 9 9 16 0 1 12 1 9 10 9 16 13 12 9 2
33 8 8 8 13 1 9 10 9 13 14 10 9 1 9 14 12 9 1 9 10 9 2 9 15 7 10 9 10 0 14 10 9 2
37 15 13 16 10 9 10 0 1 10 9 1 10 12 1 12 10 9 13 12 9 2 7 1 15 4 9 14 12 9 2 16 13 1 9 10 9 2
25 10 9 13 16 11 13 1 10 9 1 10 9 16 13 1 15 7 7 3 13 16 10 9 13 2
17 10 9 13 3 1 9 10 9 13 14 11 11 1 9 10 9 2
40 15 13 16 1 9 10 9 16 13 2 1 9 0 7 1 9 0 2 15 13 3 16 15 13 9 1 10 9 2 7 16 0 9 16 13 1 9 10 9 2
8 10 9 1 10 9 13 3 2
50 9 10 9 7 10 9 11 11 13 1 9 10 9 1 9 11 13 1 9 10 9 2 1 9 9 10 9 2 16 3 13 1 10 9 2 13 9 1 9 9 2 16 1 15 13 11 1 9 9 2
13 1 3 13 9 1 9 9 1 9 1 11 3 2
41 1 9 10 9 13 16 9 15 14 11 13 13 3 14 9 9 10 9 1 10 9 2 16 9 15 13 3 1 12 9 1 9 10 9 2 1 12 1 9 11 2
26 1 9 10 9 13 3 16 9 15 1 13 1 10 9 10 0 16 13 13 9 0 1 9 10 9 2
32 9 10 9 13 14 9 15 1 9 10 9 1 10 0 1 12 9 7 13 0 1 9 11 16 13 3 7 1 9 10 9 2
32 3 13 1 9 10 9 16 12 10 9 10 0 1 10 9 3 13 9 9 7 15 4 13 1 10 9 1 10 9 10 0 2
10 11 2 0 1 2 10 9 2 2 2
33 9 0 3 13 1 9 11 1 9 10 12 2 3 1 9 9 10 11 2 11 2 9 2 7 13 9 0 1 9 3 2 0 2
14 15 13 1 9 16 13 1 11 7 1 9 0 0 2
15 10 9 15 13 3 1 9 10 9 1 11 7 1 11 2
15 9 10 9 13 13 1 9 1 9 14 9 0 1 11 2
16 15 13 1 13 1 9 10 1 10 9 10 0 14 9 11 2
12 1 1 9 13 9 10 9 14 15 1 11 2
28 1 10 9 13 1 11 14 10 9 14 10 9 1 10 3 2 9 16 13 1 12 14 9 10 9 1 11 2
7 1 9 15 13 12 9 2
27 10 3 2 9 13 3 1 9 13 1 9 2 7 9 1 11 2 1 16 3 13 9 1 9 10 9 2
27 1 9 1 11 1 10 9 13 9 15 14 10 9 11 11 2 16 13 9 9 10 9 1 9 10 12 2
19 2 9 11 2 2 16 16 13 9 10 9 1 11 2 13 1 9 15 2
23 10 9 13 3 1 11 2 1 9 10 12 2 1 9 13 1 10 9 10 0 14 11 2
18 3 1 11 13 9 14 10 9 15 13 3 1 12 7 13 1 12 2
21 1 11 3 13 9 14 10 9 2 1 9 9 2 7 13 1 9 15 9 0 2
20 9 15 13 13 9 1 9 9 2 9 7 9 0 2 1 9 14 9 0 2
28 1 11 13 9 16 13 9 1 9 1 10 9 10 0 1 9 3 2 0 0 1 9 2 11 10 0 2 2
33 9 0 1 11 13 1 10 9 2 16 10 9 13 1 16 10 10 9 13 0 2 7 10 9 10 0 13 13 9 16 9 15 2
21 9 10 9 10 0 11 13 16 9 10 9 13 1 9 15 14 10 9 10 0 2
31 9 15 13 1 9 7 1 9 1 2 9 0 2 7 2 9 0 2 2 3 3 1 9 11 7 3 1 9 10 9 2
10 13 13 13 1 10 9 7 3 4 2
15 9 3 0 1 10 9 3 4 13 1 10 9 10 0 2
12 13 9 2 15 13 3 3 1 9 2 9 2
17 7 15 13 14 9 9 10 9 2 9 3 2 0 15 12 9 2
20 7 7 9 0 13 13 15 1 2 9 9 15 1 9 9 10 9 10 0 2
23 1 9 10 9 13 9 14 9 1 0 7 0 10 0 13 7 10 0 13 1 9 9 2
32 15 16 13 13 2 0 2 7 7 3 3 2 1 9 9 1 9 2 9 2 15 13 13 15 1 9 0 14 9 2 9 2
37 9 15 3 13 7 13 1 10 9 10 3 2 13 14 10 9 2 16 4 1 9 15 13 9 2 13 2 13 9 2 1 13 9 7 13 9 2
41 3 9 9 0 2 9 13 9 0 1 10 9 14 10 9 10 0 14 3 7 1 9 10 9 14 10 9 10 0 14 3 2 1 13 13 10 12 1 10 9 2
39 7 1 10 9 16 13 1 9 15 2 1 9 0 7 1 9 0 1 10 9 2 4 13 3 12 9 13 1 9 10 9 2 16 3 13 9 10 9 2
52 3 13 9 2 9 0 2 9 0 1 10 9 13 1 10 9 2 16 3 2 13 2 10 9 0 1 9 10 9 2 13 10 3 2 9 2 10 9 14 9 11 13 2 7 10 9 13 9 0 1 11 2
31 7 10 9 10 0 2 10 0 7 10 0 13 1 9 0 3 2 1 10 16 13 2 7 2 1 9 9 2 10 9 2
19 10 9 10 0 13 1 9 3 13 1 9 10 9 10 0 7 10 0 2
11 7 1 9 9 2 3 9 13 14 15 2
42 15 16 13 13 1 10 9 1 1 9 10 9 13 9 1 10 9 10 0 1 10 10 9 2 1 9 0 14 9 7 9 2 3 3 16 13 1 2 9 0 2 2
23 10 9 10 0 11 3 13 3 16 3 16 3 13 13 1 10 9 13 13 14 15 3 2
32 9 15 14 9 0 13 9 1 10 9 2 7 9 15 10 0 1 9 10 9 2 16 16 15 2 4 13 3 9 1 9 2
43 9 10 9 10 0 2 3 7 13 9 15 13 1 9 0 9 2 9 0 2 13 15 3 1 10 9 10 0 13 1 9 11 2 1 15 9 14 9 7 14 9 9 2
39 3 2 4 13 16 9 10 0 1 9 10 9 10 0 2 0 13 1 9 9 15 14 9 10 9 2 16 13 15 9 9 14 9 2 9 0 1 9 2
23 10 10 9 10 0 13 1 9 10 9 1 9 9 2 7 3 1 9 15 13 10 9 2
42 0 10 9 2 9 9 9 0 2 13 9 0 7 13 14 9 15 1 10 9 10 0 14 10 9 2 1 15 13 15 16 13 9 7 9 1 10 9 7 3 3 2
36 7 3 13 16 10 9 1 10 9 13 1 10 10 9 10 15 2 16 16 13 1 9 9 10 12 7 10 12 2 9 0 2 3 9 9 2
28 15 13 1 15 14 10 15 16 3 13 3 2 16 3 13 2 7 1 10 9 10 15 10 9 13 1 9 2
30 7 3 10 0 14 9 9 10 12 13 1 9 10 9 10 0 7 3 13 1 9 15 1 9 7 1 3 9 9 2
30 7 7 2 1 2 9 2 15 2 9 10 9 13 9 9 2 9 10 9 10 0 2 15 3 9 14 9 10 9 2
22 1 9 15 14 10 9 13 1 15 1 2 9 9 15 7 15 13 14 9 9 15 2
28 10 9 1 9 10 9 10 0 14 9 10 9 1 2 9 9 14 9 0 2 13 1 15 16 9 3 13 2
16 9 9 10 9 16 1 15 13 9 9 3 13 1 9 7 2
83 4 13 1 12 9 1 10 9 16 13 1 10 9 15 12 9 2 11 2 9 9 16 1 9 15 13 9 1 10 9 10 0 1 9 10 9 13 14 15 1 9 2 13 3 14 9 15 10 3 2 0 2 0 7 13 1 9 15 1 3 1 2 9 9 0 2 16 13 9 3 2 0 7 9 9 0 1 9 10 9 1 15 2
30 11 2 13 9 0 2 1 10 9 7 1 10 9 2 1 13 1 9 0 9 0 2 1 10 9 10 0 2 0 2
28 9 15 13 1 9 9 10 9 16 1 9 15 13 3 3 1 9 10 9 1 10 9 10 0 14 10 9 2
9 1 10 9 13 9 1 9 15 2
41 4 13 15 13 7 7 3 1 10 9 2 16 13 1 10 9 2 9 9 2 2 1 10 9 10 0 14 9 0 2 1 11 1 10 9 7 11 1 10 9 2
48 4 3 13 1 9 14 9 2 9 2 16 13 13 1 10 9 14 9 10 9 2 1 13 9 0 1 10 9 7 1 10 9 2 7 3 13 14 9 15 1 9 1 9 10 9 10 0 2
18 12 10 9 14 10 9 7 14 9 10 9 4 1 9 0 7 0 2
48 7 3 4 13 1 15 16 3 13 9 0 2 9 13 2 2 16 15 3 4 13 1 10 9 10 0 3 1 15 16 13 1 9 10 9 10 0 2 16 13 0 10 9 7 10 9 0 2
19 8 8 9 10 9 10 0 13 1 10 9 1 16 13 16 13 1 9 2
10 1 10 9 13 9 9 7 9 9 2
24 9 10 9 2 11 2 11 2 13 1 9 15 14 9 10 9 2 7 16 13 14 9 15 2
63 10 9 11 9 13 2 2 3 3 13 10 9 10 0 14 13 1 9 10 9 14 15 1 10 9 10 0 1 9 10 9 12 9 1 9 15 1 9 10 9 2 16 9 15 13 1 9 1 9 7 9 15 13 1 9 9 15 7 1 9 9 0 2
34 7 13 3 10 9 2 3 13 10 9 7 9 10 9 3 1 9 9 15 14 9 9 7 9 9 2 1 16 13 14 9 10 9 2
19 2 9 10 9 13 16 9 10 9 2 16 13 1 12 9 2 13 0 2
15 13 3 9 16 9 15 3 13 0 1 9 9 10 9 2
35 9 1 15 2 9 10 9 16 9 15 13 1 9 15 3 2 0 7 10 10 9 16 13 7 10 9 16 13 13 1 9 1 10 9 2
31 2 13 10 9 2 7 2 16 10 9 13 1 9 10 9 13 9 15 1 3 16 13 7 13 16 9 13 15 13 13 2
14 15 13 16 9 10 9 10 0 13 0 7 3 0 2
32 13 13 9 14 9 2 7 7 13 9 16 14 15 13 10 9 1 9 15 7 1 9 2 16 13 1 15 9 7 9 0 2
14 7 7 15 13 14 10 9 7 13 14 9 10 9 2
28 2 15 13 13 15 15 16 13 14 9 10 9 10 0 2 16 1 12 9 13 16 15 13 4 1 9 15 2
26 3 15 16 13 14 10 9 1 10 9 10 0 13 3 15 16 13 14 10 9 1 10 9 10 0 2
48 2 0 1 10 13 10 9 2 3 10 10 9 7 10 9 2 1 10 9 10 0 2 13 1 9 12 9 1 10 9 16 4 13 1 9 1 9 0 3 7 15 4 13 1 9 10 9 2
15 7 13 10 9 15 16 13 2 3 13 9 15 0 2 2
32 11 11 1 2 9 10 12 14 11 2 2 15 11 3 2 7 10 9 16 13 13 14 15 1 3 13 9 9 13 7 13 2
56 1 1 10 9 10 0 13 13 16 1 10 9 10 0 13 10 9 1 9 1 9 11 10 0 2 16 13 13 1 12 9 1 10 9 10 0 7 1 9 10 9 11 2 7 1 9 15 14 11 2 1 9 15 7 0 2
47 10 15 1 9 15 14 1 12 9 9 0 7 1 9 14 11 13 1 10 0 2 7 3 15 2 3 1 11 2 16 14 15 13 3 1 3 2 13 1 10 9 12 7 3 2 2 2
13 7 9 15 13 0 3 1 1 10 9 10 0 2
39 1 9 15 13 7 13 10 9 2 12 9 11 2 11 7 11 13 13 9 0 0 3 2 0 2 16 9 15 16 13 13 1 9 15 14 9 10 9 2
65 11 11 2 10 9 10 9 2 0 3 2 13 1 9 1 11 11 1 11 2 7 13 13 1 9 15 16 3 1 9 15 13 14 9 15 1 9 9 10 9 3 2 7 3 1 9 9 10 9 10 0 3 2 7 9 10 9 10 0 3 2 1 9 9 2
23 3 11 2 9 9 11 3 2 13 1 9 1 11 1 9 13 14 10 9 1 9 9 2
31 3 13 14 2 9 10 9 2 14 10 9 1 9 9 11 1 12 9 1 9 10 9 10 12 7 1 9 10 9 15 2
32 9 0 0 13 1 10 9 10 0 1 11 2 7 1 9 15 2 9 0 1 9 0 2 1 9 9 2 10 9 10 0 2
22 3 1 11 13 9 1 9 15 10 0 14 11 2 7 1 9 15 9 9 3 0 2
12 11 13 2 13 7 13 7 15 9 1 11 2
37 3 3 13 16 11 13 1 10 9 10 0 10 0 1 11 12 9 0 2 16 13 1 11 10 0 7 13 2 3 1 9 9 9 1 11 2 2
24 11 11 13 3 13 16 10 9 13 2 1 9 15 10 0 7 10 0 14 11 1 11 2 2
41 3 9 10 9 14 9 15 2 13 13 14 9 10 9 2 1 9 15 14 9 0 7 0 9 2 14 11 7 11 2 16 1 11 2 1 9 0 1 10 9 2
108 1 9 1 9 10 9 14 15 9 3 13 11 11 13 2 1 9 10 9 14 11 2 9 15 7 9 15 2 2 1 9 10 9 14 15 1 9 9 2 1 9 10 9 14 11 2 9 15 7 9 15 2 2 16 2 11 13 10 9 10 12 14 11 7 1 10 15 15 13 3 2 7 16 16 13 10 9 16 13 1 15 13 1 9 15 7 13 1 15 2 3 3 13 9 9 10 9 10 0 7 10 10 9 14 10 9 2 2
49 13 2 16 11 13 1 10 9 7 1 10 9 14 10 9 16 13 1 9 10 9 1 15 13 11 1 9 14 11 2 1 9 1 10 9 10 0 2 7 1 9 10 9 14 9 11 10 0 2
7 7 3 3 13 10 9 2
49 13 2 7 3 13 9 1 15 16 11 13 16 13 2 1 1 12 9 2 1 9 1 11 1 9 15 13 1 9 15 10 0 14 11 2 16 13 13 9 13 14 10 9 1 10 9 10 0 2
25 9 15 14 11 1 11 13 1 9 0 2 3 1 9 10 9 7 3 1 9 9 2 10 9 2
46 11 13 1 9 0 1 9 2 1 10 9 10 0 10 0 16 13 1 15 9 10 9 7 9 2 10 9 1 9 2 16 3 13 1 9 1 10 9 1 9 16 13 14 10 9 2
22 1 15 4 13 2 3 2 13 10 9 10 0 10 0 16 13 12 10 9 1 11 2
75 4 13 13 0 1 15 9 2 16 1 9 10 9 4 11 13 14 9 15 10 0 1 9 9 15 7 1 10 9 1 10 9 10 0 16 13 1 9 15 1 9 10 9 7 3 15 2 9 10 9 7 9 2 10 9 13 2 3 1 9 15 14 10 9 2 13 9 0 1 12 12 9 1 11 2
84 11 4 13 1 9 9 15 2 7 9 9 15 15 2 7 7 3 1 12 1 10 9 10 0 2 7 0 3 1 9 15 2 1 9 0 1 15 2 9 14 3 1 9 10 9 10 0 2 16 14 9 15 13 13 10 9 1 10 9 9 15 2 9 14 3 1 9 10 9 14 11 2 1 9 9 10 9 16 13 1 9 9 15 2
35 4 13 16 9 9 15 10 0 14 11 2 1 9 10 9 1 9 7 1 9 2 13 0 1 15 9 7 15 13 4 13 1 9 15 2
38 3 4 13 3 9 15 3 13 14 15 9 0 12 2 1 3 13 1 11 11 10 10 9 10 0 10 0 16 13 1 15 3 1 9 15 1 11 2
45 11 11 2 7 13 1 9 10 9 16 13 1 10 9 2 13 13 1 9 11 13 9 1 10 9 10 0 1 9 10 9 2 1 15 9 9 2 9 9 7 13 9 2 2 2
37 7 3 13 9 11 11 3 2 4 10 9 16 13 3 1 9 13 9 0 12 9 2 1 9 7 1 9 2 1 10 9 10 3 10 3 0 2
20 4 1 9 10 9 10 0 13 1 10 9 10 3 10 3 0 13 1 15 2
44 1 10 9 7 1 10 9 10 0 1 10 9 13 9 1 9 15 14 9 11 11 2 11 2 1 9 9 2 1 9 9 9 9 9 10 9 1 9 11 11 1 9 11 2
15 9 15 13 1 11 1 10 9 16 13 1 9 9 11 2
41 9 0 1 10 9 2 7 1 9 15 9 1 10 9 2 13 16 4 13 1 9 0 15 14 9 9 9 10 9 2 3 9 16 11 13 14 9 9 10 9 2
23 3 9 10 9 7 10 9 11 11 2 16 11 13 1 9 15 2 3 13 1 10 9 2
24 1 15 2 1 9 1 11 2 13 11 1 11 16 13 9 13 1 15 9 1 9 10 9 2
18 3 13 1 10 9 16 3 4 13 1 11 12 9 1 9 10 9 2
22 3 13 1 9 15 10 9 11 9 2 1 9 9 9 10 9 2 7 9 11 11 2
35 1 9 10 9 10 0 13 1 15 1 9 9 11 11 11 1 11 2 7 1 9 10 9 16 13 1 11 3 9 11 13 1 10 9 2
21 9 0 1 10 9 13 16 2 10 10 9 13 0 7 3 13 1 10 9 2 2
34 9 1 10 9 13 3 16 3 4 16 11 13 1 9 9 2 1 13 9 0 1 9 10 9 9 11 11 2 16 13 1 9 0 2
30 1 11 13 9 9 9 10 9 7 10 9 2 7 7 2 3 13 10 9 12 9 14 9 9 10 9 1 9 11 2
23 9 2 9 11 13 1 9 16 2 9 10 9 1 10 9 7 1 9 10 9 13 3 2
38 13 9 1 15 2 7 1 15 13 9 16 10 9 3 13 1 9 9 9 9 10 9 2 1 9 16 9 10 9 13 1 9 0 1 10 9 2 2
10 9 7 13 13 9 13 1 10 9 2
22 11 11 2 12 2 2 9 0 2 13 1 9 1 9 11 2 13 3 1 9 15 2
19 15 13 1 9 15 1 10 9 1 9 0 1 10 9 11 2 1 11 2
6 15 13 1 9 15 2
35 11 11 2 12 2 2 13 13 14 9 15 1 9 9 1 9 11 2 1 3 13 10 9 10 0 1 9 15 2 11 2 9 10 12 2
13 10 12 13 13 14 9 15 14 11 1 9 0 2
7 10 9 13 14 15 3 2
11 1 11 13 16 10 9 13 1 10 9 2
21 2 13 2 2 13 1 9 13 1 9 15 2 2 13 13 1 15 9 9 2 2
22 1 9 7 9 13 10 9 13 1 10 9 2 1 15 9 2 10 9 13 0 3 2
5 9 15 13 13 2
23 11 13 1 9 15 1 9 11 2 3 13 14 15 13 1 10 9 7 13 1 9 15 2
22 1 2 9 9 10 9 2 15 13 9 9 9 0 1 9 15 7 13 1 10 9 2
23 2 15 13 14 9 9 15 2 13 1 9 1 9 15 11 1 10 9 2 7 3 13 2
43 9 10 9 1 11 13 3 1 10 9 16 11 3 4 13 13 1 9 15 2 7 9 1 10 9 13 10 9 2 11 11 2 1 9 16 13 14 9 15 1 10 9 2
21 12 12 9 1 11 2 1 15 1 1 12 12 9 7 9 2 13 1 9 11 2
16 3 3 0 13 9 15 14 9 15 7 13 1 9 10 9 2
43 9 15 14 10 9 2 16 9 15 10 0 2 16 13 2 7 9 10 9 10 0 14 15 13 14 9 15 14 10 9 7 14 9 2 13 9 16 13 9 0 7 9 2
21 9 7 13 13 2 15 13 1 9 10 9 2 3 15 14 10 9 7 10 0 2
15 1 10 9 15 9 1 9 7 9 0 2 3 7 3 2
17 1 12 9 9 15 15 13 3 12 1 9 10 9 1 10 9 2
17 3 9 0 7 9 9 13 3 13 9 1 10 13 1 9 0 2
46 9 1 9 9 10 9 1 9 0 0 4 3 13 14 10 9 1 10 9 1 9 11 2 13 14 10 9 10 0 2 16 3 3 13 1 15 3 9 0 2 1 9 9 9 12 2
10 7 9 7 9 3 13 1 9 0 2
16 7 3 0 2 16 13 9 10 9 13 9 1 9 10 9 2
29 3 2 9 0 0 1 9 11 3 13 1 3 15 1 9 9 0 0 2 7 13 1 15 1 9 15 1 3 2
32 9 0 13 14 10 9 7 13 2 1 10 9 2 1 10 9 1 9 10 9 2 7 9 11 13 13 9 0 1 10 9 2
48 7 3 9 0 16 13 13 0 2 13 3 1 13 10 9 1 10 16 13 1 9 7 9 2 3 1 16 9 13 13 1 10 9 1 9 15 7 0 7 13 13 13 1 9 15 10 0 2
28 9 16 13 1 9 7 9 1 9 1 10 9 13 1 9 9 1 9 7 1 13 9 1 9 15 14 9 2
19 10 9 13 13 13 1 9 9 0 7 1 9 9 16 13 0 1 15 2
23 9 0 9 12 2 7 2 13 13 12 9 1 16 10 9 1 11 13 13 1 15 9 2
18 9 12 13 1 9 2 9 2 2 9 9 1 9 7 9 1 9 2
15 3 13 1 9 15 9 0 7 3 13 9 1 9 15 2
24 9 15 14 10 9 13 1 9 15 9 7 13 13 14 15 13 1 9 15 2 16 13 13 2
23 1 10 9 10 0 2 9 13 9 14 9 1 9 15 2 2 13 9 10 9 11 11 2
28 1 9 10 9 13 10 9 14 10 9 2 1 10 9 13 14 10 9 2 9 0 7 0 13 9 9 9 2
50 1 2 9 10 9 2 3 2 0 10 9 7 10 9 1 11 1 3 9 10 12 2 16 13 10 9 11 11 11 2 11 2 10 9 10 0 2 9 11 10 0 2 13 1 9 9 1 9 15 2
36 9 13 13 1 12 12 9 1 10 9 7 12 9 1 10 9 2 7 10 9 0 13 13 13 15 16 15 13 13 1 9 14 9 9 15 2
9 7 9 1 9 2 10 9 0 2
30 13 3 13 10 9 13 2 9 10 9 2 7 2 10 9 13 10 9 2 10 9 13 9 7 9 13 1 9 2 2
18 3 3 9 13 3 3 10 9 10 12 2 3 10 0 2 14 11 2
13 1 15 2 10 9 15 13 0 9 3 7 3 2
27 7 16 10 9 13 1 3 1 9 2 7 3 16 10 13 1 9 0 2 13 15 3 0 3 0 3 2
47 3 2 10 9 13 1 9 15 9 2 16 1 9 1 9 15 13 1 9 0 1 9 10 9 2 2 13 10 9 11 11 1 9 15 2 9 1 9 10 9 2 2 11 2 12 2 2
23 1 2 9 10 9 4 9 13 9 2 13 1 9 15 7 13 1 9 15 1 9 15 2
28 15 13 4 1 9 15 2 7 2 1 9 3 13 4 13 13 1 10 9 1 10 9 0 2 2 13 11 2
20 15 13 1 10 12 10 12 2 7 10 9 13 3 1 9 10 9 10 0 2
21 3 1 10 9 10 0 9 15 14 10 9 13 0 3 7 1 10 9 10 0 2
12 15 2 3 1 9 10 9 10 0 10 3 2
26 9 13 3 7 13 1 9 15 3 0 3 2 1 9 1 10 15 2 1 10 9 4 3 3 3 2
54 15 13 1 9 9 10 9 2 15 9 9 0 2 10 9 1 15 13 7 13 2 13 1 9 9 1 9 16 13 0 9 2 1 10 9 0 2 7 10 9 3 13 14 9 15 1 10 9 2 10 9 10 0 2
41 1 9 9 7 9 9 1 9 2 13 9 15 1 10 9 16 13 1 11 1 9 13 7 13 1 15 2 1 1 9 9 10 9 15 13 1 9 13 7 0 2
15 1 10 9 10 9 2 0 16 15 13 4 13 10 9 2
7 10 9 13 3 9 9 2
6 15 13 1 9 9 2
9 10 9 10 0 13 4 13 3 2
6 9 15 13 9 15 2
11 15 3 13 4 13 9 1 9 0 15 2
15 2 3 16 13 3 13 3 9 0 2 2 13 9 0 2
25 1 10 4 10 9 13 9 13 10 9 11 1 9 15 0 10 9 2 12 9 0 14 11 2 2
25 10 9 13 3 2 1 9 15 14 11 10 0 1 11 2 13 14 15 11 9 15 1 9 15 2
7 12 9 13 10 9 15 2
11 7 13 1 9 1 9 11 4 1 15 2
17 2 3 2 9 15 14 10 9 13 3 1 9 2 2 13 11 2
15 1 10 9 2 1 10 9 2 13 10 9 14 10 9 2
45 9 15 14 11 13 1 9 14 9 0 2 7 13 1 15 9 0 2 15 13 3 1 9 0 16 13 0 1 9 15 9 0 7 13 3 1 10 9 2 1 11 1 10 9 2
37 9 7 9 0 1 11 13 1 9 9 9 2 9 2 9 7 9 0 2 9 2 9 7 9 2 9 1 10 9 14 10 9 7 3 10 9 2
15 7 9 13 1 10 9 1 9 2 13 3 9 7 9 2
13 3 13 9 1 9 10 9 2 1 9 10 9 2
19 7 16 2 1 9 2 13 9 3 2 13 3 9 9 1 9 10 9 2
23 9 9 0 7 0 13 9 15 1 11 2 1 11 7 1 11 2 1 12 1 12 9 2
19 7 10 9 13 13 9 9 0 2 7 4 13 14 10 9 1 10 9 2
5 3 13 9 0 2
4 10 9 13 2
21 3 0 10 9 13 4 13 7 3 3 13 2 16 16 13 1 15 1 9 0 2
8 13 9 1 11 16 13 9 2
19 15 13 9 9 16 13 16 9 0 1 10 9 13 10 9 1 9 15 2
13 4 3 1 10 9 13 7 15 13 1 10 9 2
11 9 13 14 10 9 2 7 10 9 13 2
26 3 2 10 10 9 16 4 13 1 9 9 9 15 13 7 13 2 7 14 10 10 9 3 13 9 2
15 1 9 0 13 10 9 1 10 9 1 12 1 12 9 2
23 1 11 13 9 0 1 9 0 2 16 4 13 1 10 9 14 10 9 13 1 9 11 2
17 1 9 1 10 15 2 10 9 4 13 1 9 1 12 12 9 2
24 9 10 9 1 9 11 0 1 9 0 16 10 9 1 10 9 13 1 15 10 9 10 0 2
7 7 3 3 3 15 0 2
16 9 9 12 13 9 0 1 9 15 16 13 1 9 1 11 2
16 2 13 3 13 14 15 2 2 13 3 3 1 9 10 9 2
8 9 13 3 3 1 9 9 2
14 1 10 9 16 13 13 12 9 10 13 1 9 9 2
41 11 11 2 12 2 13 14 9 15 3 2 11 11 2 12 2 2 13 14 15 7 13 14 15 2 7 13 14 9 15 10 0 2 11 9 10 12 2 1 11 2
18 9 0 3 1 10 15 13 10 9 10 0 11 11 1 9 9 15 2
15 15 13 1 9 0 13 1 9 15 10 0 3 14 11 2
32 9 12 13 1 15 11 2 13 1 15 16 15 2 9 2 16 2 0 1 9 2 2 13 1 15 7 13 14 15 12 9 2
9 10 9 13 16 3 1 9 13 2
27 9 9 10 9 1 9 1 10 9 2 11 11 2 13 13 14 9 15 1 10 9 13 1 9 1 11 2
21 10 9 13 1 16 9 9 10 9 14 11 13 12 9 0 7 13 9 7 9 2
29 9 10 9 1 9 1 10 9 13 9 9 10 9 2 1 16 13 10 9 1 9 13 1 9 16 13 1 11 2
31 1 10 9 2 16 13 1 9 1 9 10 9 2 13 16 10 16 13 13 1 9 1 11 4 16 13 3 14 9 15 2
26 10 9 13 1 12 9 9 16 13 9 1 11 2 7 13 1 9 10 9 1 9 10 9 1 11 2
30 10 9 13 13 1 10 3 16 13 1 9 1 11 14 9 10 9 7 13 1 9 15 14 10 9 7 13 1 11 2
12 3 13 9 1 10 10 9 16 13 1 11 2
30 9 11 13 1 10 9 10 0 14 9 15 1 10 9 10 0 10 0 2 3 1 9 9 9 10 9 1 9 11 2
18 13 16 9 9 15 13 16 13 14 9 11 16 13 1 11 1 9 2
16 9 15 13 14 10 9 1 9 9 9 1 9 1 9 11 2
19 1 13 1 15 13 10 9 13 14 10 9 1 9 16 13 1 9 9 2
36 15 13 14 9 10 9 1 9 10 9 1 11 1 11 7 1 11 2 7 3 3 13 4 13 1 3 1 9 1 9 2 1 1 10 9 2
8 3 13 10 9 1 10 9 2
24 9 9 13 16 7 13 3 10 9 13 14 10 9 3 13 1 11 2 3 13 13 1 15 2
89 2 13 10 9 13 1 9 0 13 14 9 15 1 9 16 1 15 13 1 15 9 0 2 2 13 10 9 2 2 7 16 16 9 10 9 10 0 13 9 1 9 10 9 1 9 0 13 1 9 1 10 9 16 13 1 0 1 15 2 3 9 1 10 9 10 0 1 11 16 13 1 15 13 1 9 1 9 1 9 16 1 15 13 9 1 9 0 2 2
40 13 1 9 10 9 2 11 2 11 2 11 2 11 7 0 2 13 1 9 10 9 10 0 14 15 2 3 9 1 9 0 1 9 9 10 9 7 9 9 2
22 1 9 15 13 1 9 10 9 14 11 2 16 15 1 10 9 16 13 1 9 15 2
20 1 9 1 15 13 16 10 9 0 1 9 9 11 16 4 13 1 9 0 2
23 3 16 13 13 1 9 12 14 10 10 9 7 3 10 1 15 2 4 13 1 9 3 2
12 1 9 9 12 3 3 13 13 14 10 9 2
19 10 9 2 1 9 9 2 11 2 2 13 1 9 14 12 9 12 9 2
24 1 9 10 9 13 3 9 14 9 1 9 0 1 9 9 2 7 3 9 11 1 9 0 2
60 3 4 13 3 2 1 10 9 2 9 9 1 9 1 12 9 2 9 9 1 9 1 12 9 2 9 0 3 2 1 9 9 1 9 2 1 12 9 2 7 9 9 0 2 0 2 1 9 0 2 1 12 2 1 12 9 1 10 9 2
18 3 13 9 2 9 2 1 10 9 1 12 9 2 1 9 0 3 2
27 9 9 7 9 9 13 10 0 3 1 9 15 2 13 11 11 2 16 13 14 10 9 1 11 1 11 2
18 9 1 9 13 14 9 10 9 10 0 7 10 0 1 9 12 9 2
13 10 9 2 13 1 12 9 7 1 1 12 9 2
9 10 9 1 12 7 1 1 12 2
22 9 9 13 1 1 9 12 7 9 9 1 1 9 12 2 7 3 1 10 10 9 2
27 9 9 1 9 9 11 2 1 9 0 0 2 13 12 9 1 12 9 1 10 9 2 7 10 9 0 2
20 9 9 14 2 11 2 3 13 1 9 0 2 12 9 1 12 1 10 9 2
54 1 10 9 13 10 9 11 0 0 2 1 1 12 9 2 1 12 9 2 2 11 1 9 7 1 9 11 2 11 13 12 9 2 9 9 0 1 9 7 3 9 0 14 9 2 9 1 9 9 13 1 12 9 2
37 3 4 13 3 14 11 2 11 2 9 16 9 0 13 1 15 1 7 10 9 10 0 2 9 0 2 2 1 12 9 2 2 1 12 9 2 2
18 3 9 9 13 2 1 9 12 9 2 10 9 0 1 10 9 2 2
25 1 9 10 9 4 13 14 2 11 2 2 16 1 2 11 2 13 9 1 10 9 1 10 9 2
6 9 11 13 12 9 2
60 9 9 1 9 11 2 1 9 0 2 13 12 1 12 9 2 1 9 9 10 9 13 12 9 2 9 9 1 9 9 15 13 12 9 2 9 0 2 1 12 2 1 10 9 13 9 9 2 11 2 9 2 12 2 1 12 1 12 9 2
22 13 3 9 9 11 1 9 2 11 2 7 2 11 2 2 9 9 11 13 12 9 2
14 2 11 2 3 13 7 13 9 2 11 2 1 11 2
22 9 1 3 1 9 0 13 3 12 9 1 12 9 2 9 1 3 16 13 9 0 2
10 9 11 0 13 12 9 7 12 9 2
24 1 10 9 10 0 13 3 9 9 2 9 0 1 9 0 16 13 13 1 10 9 10 0 2
16 10 9 3 13 1 10 9 7 13 1 9 13 14 10 9 2
36 9 9 13 12 7 1 9 10 9 3 0 2 9 9 1 9 2 9 9 1 9 16 13 1 0 2 13 12 9 1 12 9 1 9 0 2
26 3 13 2 11 2 1 9 1 9 2 11 2 10 0 16 13 14 10 9 13 9 15 1 10 9 2
33 13 1 11 1 9 0 1 9 3 0 1 9 0 9 10 9 9 2 7 4 13 16 1 10 9 13 3 15 1 9 10 9 2
56 4 13 1 2 11 2 1 15 16 10 9 14 9 10 9 16 4 13 2 1 9 10 9 2 1 10 9 2 0 1 15 1 9 9 16 13 1 10 9 3 1 10 9 2 3 16 3 10 9 0 9 15 1 10 9 2
52 9 10 9 13 1 9 2 9 2 1 9 10 11 12 2 1 9 2 11 2 1 9 10 9 2 9 11 2 1 11 2 1 11 2 1 9 11 12 2 1 11 2 1 9 11 7 1 9 10 9 12 2
6 2 11 2 11 2 2
13 11 9 11 13 3 13 14 9 15 1 9 0 2
24 9 10 9 10 0 13 1 9 10 9 16 13 3 9 1 9 9 13 0 7 9 0 0 2
24 2 9 10 9 13 1 16 13 10 9 10 0 2 2 13 10 9 1 9 10 9 10 0 2
15 11 13 1 3 1 9 0 1 3 13 10 9 1 12 2
15 10 9 1 9 13 14 10 9 1 9 0 1 10 9 2
31 1 11 13 16 12 9 13 3 14 15 13 1 9 1 9 1 9 10 9 1 7 10 9 16 13 10 9 1 9 15 2
23 9 10 9 13 16 15 13 9 1 9 1 10 9 10 0 16 13 13 9 1 9 11 2
15 1 10 9 13 1 9 0 7 0 2 7 1 15 13 2
10 10 9 10 0 13 14 15 1 0 2
8 3 13 3 9 1 10 9 2
24 9 15 13 14 15 1 9 0 0 7 13 1 15 9 13 1 10 9 1 10 9 10 0 2
10 9 10 9 1 10 9 13 0 3 2
12 3 13 16 0 13 13 9 1 9 10 9 2
13 3 3 3 13 9 1 10 9 7 13 1 15 2
14 3 2 1 10 9 10 0 13 9 0 1 9 0 2
27 7 13 9 15 1 9 0 10 3 2 1 9 9 9 2 13 9 16 9 10 9 3 3 13 3 0 2
39 9 10 9 7 10 9 3 13 3 3 1 9 1 9 15 2 3 1 9 10 9 2 1 10 11 2 2 7 3 13 14 9 15 14 10 9 10 0 2
2 3 2
7 3 1 9 15 13 9 2
9 9 10 9 13 1 9 10 9 2
14 13 10 9 16 13 1 9 15 2 3 1 9 9 2
19 1 10 9 16 13 1 9 9 13 10 1 15 9 2 7 10 13 13 2
11 7 1 9 3 13 13 1 15 9 0 2
10 1 10 9 9 13 9 9 7 9 2
9 15 9 14 9 15 7 3 3 2
27 1 10 9 13 9 0 2 11 2 9 2 16 1 9 15 13 9 1 10 9 2 7 3 9 14 15 2
21 1 9 1 10 15 2 16 1 15 12 12 9 2 13 16 13 9 1 9 9 2
30 3 13 13 14 10 9 2 7 13 10 9 1 15 16 10 11 13 16 13 1 9 9 7 13 14 15 1 9 9 2
2 3 2
12 10 9 10 9 10 0 13 9 1 10 9 2
33 13 9 9 7 9 2 16 1 15 9 3 11 11 2 7 15 13 1 10 9 14 9 10 9 2 10 9 10 0 10 0 2 2
5 10 9 13 0 2
18 15 13 13 1 9 10 9 10 0 2 7 3 15 9 1 10 9 2
22 13 9 16 15 13 1 9 15 9 0 2 9 2 3 9 2 7 9 9 7 11 2
26 10 9 13 1 9 9 16 10 9 3 3 13 13 2 7 1 9 15 9 10 9 1 10 9 13 2
19 1 9 9 2 1 9 10 9 13 11 0 11 0 16 13 1 15 9 2
18 7 1 3 3 13 14 15 2 7 7 13 1 9 1 9 3 0 2
18 13 13 1 9 15 2 7 15 13 1 9 15 1 9 1 14 15 2
24 1 9 10 9 10 0 10 9 1 10 11 13 3 9 0 3 7 1 10 11 1 10 9 2
15 13 13 3 16 4 13 14 10 11 13 14 9 9 15 2
10 3 2 10 9 1 9 10 9 0 2
7 10 9 13 0 7 0 2
12 1 10 9 7 10 9 9 9 2 15 0 2
8 7 15 13 1 9 10 9 2
14 0 9 9 1 9 9 9 10 9 7 10 9 3 2
19 10 9 10 0 3 1 9 15 13 11 11 2 9 15 14 11 11 2 2
7 10 3 13 15 10 9 2
5 16 13 9 0 2
6 3 3 13 9 0 2
5 3 13 9 0 2
14 7 10 9 1 9 11 13 2 3 2 1 10 9 2
21 1 1 9 2 9 10 9 10 0 1 10 9 13 14 9 9 15 14 10 9 2
18 1 9 0 2 1 15 2 15 13 3 1 9 3 1 3 2 3 2
19 16 16 10 9 10 0 13 2 4 13 9 0 3 1 10 9 10 0 2
14 9 3 13 1 10 9 13 4 13 10 9 10 0 2
21 1 11 13 3 9 0 0 3 2 16 16 10 9 1 10 9 10 0 3 13 2
7 13 1 15 3 9 0 2
27 7 1 9 15 2 13 10 9 1 15 16 9 15 13 1 9 1 10 9 10 0 2 7 1 9 0 2
23 0 16 3 11 11 13 9 16 9 15 13 1 9 15 2 7 15 13 3 1 9 0 2
17 15 13 1 9 0 7 0 1 10 9 2 9 2 11 2 11 2
15 3 15 13 1 9 1 9 0 1 10 9 1 11 11 2
6 1 15 13 14 15 2
28 7 1 7 9 15 10 0 14 10 11 2 11 2 9 2 15 3 13 3 13 16 9 1 10 15 3 0 2
9 3 1 15 16 3 13 0 3 2
16 1 12 2 16 13 1 10 9 2 13 1 15 1 9 0 2
8 3 3 13 14 15 1 9 2
25 3 2 3 1 15 12 9 2 13 9 11 1 10 9 1 9 16 13 9 0 0 14 10 9 2
14 7 1 9 14 9 2 13 10 9 1 9 0 0 2
13 1 12 9 9 10 9 13 12 9 7 9 9 2
13 1 3 3 13 7 7 9 12 1 10 9 15 2
12 10 9 7 9 3 13 14 10 9 1 15 2
17 13 9 16 10 13 1 9 10 9 13 13 14 10 9 10 0 2
59 10 9 13 1 15 14 9 10 9 10 0 2 7 7 10 9 11 11 13 16 9 1 10 9 10 0 2 1 2 10 9 1 9 0 2 2 0 1 10 9 15 16 16 15 4 2 13 1 10 9 14 9 10 9 7 10 9 2 2
24 12 12 9 9 10 9 13 2 1 9 9 1 10 9 2 13 1 10 9 1 9 10 9 2
26 14 10 9 13 2 10 9 10 0 10 0 14 11 2 9 9 16 13 14 9 10 9 1 10 9 2
44 1 16 1 10 9 3 13 9 1 9 9 1 9 9 10 9 2 13 9 16 15 13 2 7 7 1 10 9 10 0 1 12 13 10 9 9 7 9 9 1 13 9 0 2
13 1 10 15 13 16 10 9 3 13 9 1 11 2
35 1 12 9 13 10 9 11 10 9 10 0 16 13 1 10 9 1 3 10 9 10 0 2 16 13 1 12 1 9 9 10 9 10 0 2
17 9 15 14 11 13 13 1 9 7 1 9 15 13 12 9 9 2
50 10 9 11 2 1 9 9 2 13 4 13 9 0 2 7 9 9 15 10 0 2 0 16 9 10 9 3 2 11 11 11 2 13 1 10 9 2 13 1 3 13 1 16 11 13 1 9 9 0 2
11 11 15 13 1 9 9 10 9 10 0 2
66 9 11 11 11 2 16 1 9 15 2 1 9 9 10 12 2 13 1 10 13 9 0 7 12 9 1 9 9 0 1 10 9 10 0 2 13 10 9 10 13 1 1 1 9 2 16 9 10 9 10 0 13 16 10 9 13 1 9 10 9 3 13 1 10 9 2
43 1 10 9 13 3 12 10 9 10 13 9 9 11 9 3 2 11 11 2 1 2 9 10 9 10 0 2 10 0 2 7 11 11 11 1 2 9 10 9 10 0 2 2
44 12 10 9 13 1 9 9 0 1 13 14 11 1 10 9 10 0 2 7 0 1 10 9 7 9 11 2 16 13 9 1 10 13 1 2 9 10 0 14 10 9 11 2 2
38 13 16 10 12 4 13 15 1 15 9 0 2 1 1 9 2 7 9 1 15 3 13 13 1 3 1 12 9 1 10 9 1 10 9 10 0 3 2
24 9 12 2 1 1 12 9 2 13 11 2 11 2 11 7 12 9 1 10 9 14 9 11 2
104 11 11 2 9 9 9 9 14 12 9 1 11 2 13 3 1 9 15 14 9 1 9 2 13 0 1 9 10 9 2 9 15 11 2 1 9 9 0 2 13 1 11 1 9 2 9 1 9 9 1 10 11 2 7 3 15 13 9 13 3 1 10 9 10 3 0 14 15 2 9 15 11 9 10 12 13 3 1 11 2 7 1 9 10 9 13 3 9 9 2 2 1 16 3 13 1 9 1 10 9 10 0 2 2
14 9 9 11 13 13 1 9 14 9 10 9 10 0 2
34 1 11 15 13 1 10 12 1 11 2 7 1 9 10 9 3 13 1 9 9 15 14 9 15 14 11 1 9 10 9 1 9 9 2
8 9 3 3 13 1 10 9 2
27 1 15 13 1 12 1 1 12 10 9 16 13 14 9 10 9 10 0 1 11 1 9 10 9 10 0 2
49 1 10 9 16 13 3 1 3 1 10 9 11 2 11 1 9 2 10 13 10 9 0 1 10 12 10 12 2 2 13 10 9 1 9 11 11 14 9 15 14 10 9 1 9 15 14 10 9 2
20 2 3 16 13 14 10 9 1 10 9 13 10 9 10 0 16 13 1 15 2
19 10 9 4 13 1 9 10 9 9 0 7 0 2 1 3 9 0 2 2
30 10 10 9 1 10 9 2 9 10 9 10 0 2 3 13 3 14 10 9 1 9 0 1 9 9 15 7 9 15 2
38 1 9 0 13 10 9 10 0 1 12 9 15 10 11 2 10 9 10 0 7 10 9 10 0 1 10 9 10 0 14 2 9 0 1 10 9 2 2
32 10 13 1 9 9 2 0 2 16 1 9 15 13 10 9 1 10 9 2 13 1 10 9 7 13 1 15 14 10 10 9 2
32 10 9 10 0 2 12 9 1 9 1 9 9 12 9 2 13 1 9 10 9 14 10 9 7 13 1 15 9 1 10 9 2
13 10 9 4 13 1 10 9 9 9 12 1 9 2
18 10 9 9 0 2 1 9 14 12 9 1 9 2 13 1 10 9 2
20 9 1 9 13 1 10 9 9 0 14 9 2 16 13 1 9 7 1 0 2
9 7 9 9 0 15 13 9 0 2
27 9 10 9 14 10 9 2 16 13 1 9 0 7 0 0 2 13 3 9 12 16 13 14 9 10 9 2
20 9 15 10 0 14 9 10 9 1 10 9 10 2 0 2 3 13 7 15 2
15 7 16 10 9 7 1 15 9 10 9 13 14 14 15 2
22 10 9 10 0 13 2 7 12 9 13 3 14 9 15 10 0 1 10 9 10 0 2
24 9 13 13 3 10 1 15 7 3 13 1 10 9 1 1 10 9 10 0 16 13 1 9 2
18 1 10 9 10 15 16 1 10 9 1 11 1 10 9 9 9 0 2
14 10 9 1 11 13 1 15 9 9 0 1 10 9 2
52 9 0 9 9 0 7 3 2 0 0 13 14 10 9 16 13 1 10 9 1 10 9 1 9 1 2 9 0 1 10 9 2 1 2 9 9 1 9 9 2 16 13 9 1 10 10 9 14 10 9 2 2
27 13 16 13 16 10 9 1 11 13 10 9 16 13 1 10 9 2 11 2 2 9 2 9 2 9 2 2
31 11 9 2 9 9 9 7 12 10 9 14 9 2 9 0 1 10 9 2 2 13 2 2 10 9 13 16 9 15 9 2
12 13 1 15 3 12 9 13 16 15 3 15 2
14 3 1 9 0 15 13 16 15 1 10 15 3 2 2
22 9 0 1 9 11 13 14 10 9 1 9 2 9 16 13 1 9 2 9 7 9 2
17 14 11 11 2 9 0 1 11 2 13 1 9 15 1 9 11 2
27 1 12 9 13 1 11 11 10 9 7 9 15 10 9 7 13 13 1 9 2 9 2 3 1 9 0 2
9 1 10 9 10 0 3 13 9 2
25 1 10 9 7 1 10 9 10 0 2 16 15 13 1 9 11 1 9 2 3 13 14 10 9 2
12 1 9 13 1 9 10 9 7 13 9 9 2
5 10 9 13 9 2
23 2 3 13 9 1 10 9 2 2 13 11 2 12 2 2 2 7 10 9 13 0 3 2
6 13 16 15 1 9 2
12 1 9 0 1 10 9 2 0 2 3 0 2
4 13 7 13 2
7 3 13 14 15 10 9 2
16 10 3 16 13 1 10 9 1 11 7 3 13 2 0 3 2
6 3 13 16 15 9 2
12 3 15 13 16 15 0 2 7 15 0 2 2
23 1 7 10 9 10 0 10 15 2 3 13 1 9 15 16 1 9 15 13 1 10 9 2
10 15 9 9 0 7 13 13 1 3 2
33 11 11 2 10 9 14 9 11 2 13 1 9 2 2 7 13 9 10 9 11 13 1 10 9 2 13 13 9 1 16 3 13 2
14 10 9 13 1 15 7 9 10 9 13 1 15 2 2
28 3 9 9 11 2 16 13 1 1 9 1 10 9 11 16 1 9 11 2 13 16 10 9 13 9 1 15 2
45 10 9 2 11 2 9 9 0 9 2 10 9 2 11 2 13 9 2 10 9 2 11 2 12 2 2 13 13 9 9 1 10 9 2 7 7 13 9 0 1 10 9 10 0 2
30 3 1 9 9 15 13 1 10 9 10 0 2 11 2 9 0 2 16 13 1 9 0 3 14 10 9 1 10 9 2
24 13 16 9 13 9 16 0 13 1 15 2 16 1 9 13 9 0 2 13 3 2 13 9 2
20 1 9 7 9 1 11 9 9 11 3 13 16 10 9 3 13 1 10 9 2
15 3 10 9 13 9 2 7 15 3 1 15 2 15 13 2
28 2 10 9 1 10 9 13 16 13 9 2 2 13 11 2 1 15 4 13 3 14 10 9 2 1 10 9 2
21 15 13 16 10 9 16 3 13 9 1 10 9 1 11 2 13 13 1 10 9 2
19 14 13 1 15 10 9 2 7 3 13 9 2 15 13 1 10 9 2 2
25 10 9 11 2 2 1 10 9 3 13 10 13 9 2 10 13 9 2 3 13 9 1 10 9 2
10 3 15 0 2 7 15 3 10 9 2
15 15 13 16 10 9 16 13 1 10 9 3 13 13 3 2
14 15 13 14 10 9 7 15 13 9 0 1 10 9 2
5 3 15 3 2 2
17 7 11 11 13 2 2 15 0 3 7 13 1 15 1 9 2 2
18 0 1 10 9 10 0 13 13 1 9 15 13 1 15 9 1 9 2
20 9 13 1 15 14 9 10 9 1 10 9 10 0 2 14 10 9 10 0 2
23 9 10 11 2 11 11 2 13 3 16 4 13 9 0 14 9 1 9 15 14 10 9 2
16 3 4 16 9 13 1 10 9 1 16 15 13 1 9 11 2
23 3 13 16 15 13 1 10 9 7 13 14 15 1 10 9 2 1 16 13 2 15 13 2
14 7 13 9 16 4 13 9 0 1 10 9 1 9 2
8 1 9 10 9 13 10 9 2
15 10 9 13 9 7 13 1 11 9 1 10 9 10 0 2
20 3 10 9 13 1 10 9 3 1 3 16 15 13 1 10 9 9 0 0 2
25 9 0 14 10 9 1 9 13 16 12 9 12 9 1 10 9 4 13 9 14 9 1 10 9 2
19 1 2 7 9 15 3 10 9 13 3 1 13 14 9 15 14 10 9 2
27 4 13 16 15 13 1 10 9 1 9 7 1 9 2 1 9 15 14 12 9 9 2 1 15 9 9 2
13 11 11 13 16 10 9 13 13 1 9 9 15 2
28 15 13 15 1 9 9 2 7 1 15 16 9 10 9 13 1 10 9 1 9 9 7 1 9 1 9 9 2
23 10 9 13 16 3 13 1 10 9 16 13 7 13 2 7 3 15 3 13 14 15 2 2
14 11 13 3 3 1 10 9 10 0 14 9 10 9 2
8 3 16 13 3 13 1 10 2
5 10 9 13 13 2
19 1 10 9 10 15 15 13 14 10 9 14 10 9 1 10 9 10 0 2
30 3 10 9 13 3 13 3 9 0 2 7 10 9 10 0 13 1 10 9 14 10 9 13 4 1 9 1 9 15 2
12 1 15 4 16 15 13 3 10 15 13 2 2
4 2 11 2 2
22 9 13 14 9 11 7 9 0 1 9 13 1 9 7 1 9 9 10 9 1 11 2
40 1 9 10 9 13 12 9 10 9 2 9 1 12 2 16 9 15 13 1 9 2 1 9 16 13 9 14 9 11 7 9 0 1 10 9 1 9 1 11 2
20 12 10 9 13 3 1 10 12 1 11 2 7 3 13 9 9 1 10 9 2
45 1 9 7 13 1 9 10 9 9 9 10 9 14 9 11 2 16 1 10 12 1 11 3 13 12 9 1 9 9 2 9 16 12 10 9 13 1 9 15 9 0 1 12 9 2
18 1 9 15 13 10 9 16 10 9 13 1 15 9 9 7 9 0 2
26 10 9 13 3 16 10 12 13 13 1 15 9 0 7 13 1 15 1 1 9 1 10 9 9 11 2
10 1 9 13 1 10 9 9 9 0 2
13 1 9 10 9 13 16 1 10 9 13 9 0 2
26 9 10 9 13 16 12 1 10 9 13 1 10 9 7 13 9 13 1 15 9 9 1 9 9 15 2
36 10 9 11 11 13 1 9 15 16 13 9 0 1 10 9 16 13 9 10 9 14 10 9 2 16 13 1 9 16 13 1 9 1 9 9 2
22 1 9 15 2 1 10 9 13 16 10 9 13 7 13 1 9 15 7 1 9 15 2
35 2 13 16 3 1 9 1 9 10 9 16 13 1 9 9 10 9 2 3 0 13 1 9 9 16 3 1 9 9 2 2 13 10 9 2
30 15 13 13 14 9 15 14 12 1 10 9 1 12 7 12 9 7 7 10 9 10 12 13 1 9 14 12 12 9 2
14 16 10 9 13 3 1 10 9 2 4 13 9 9 2
9 9 16 13 9 3 1 9 0 2
9 3 9 0 2 7 3 3 0 2
25 12 9 7 3 13 1 15 1 9 10 9 16 13 2 12 9 3 2 12 9 14 9 9 0 2
59 7 1 10 15 2 3 9 0 3 1 10 9 9 15 16 13 7 13 3 13 9 7 9 1 15 9 0 16 13 9 9 2 1 3 13 11 2 11 2 11 10 0 1 11 16 15 13 13 14 15 9 2 10 9 1 9 10 9 2
34 8 2 8 7 12 7 9 9 2 7 3 3 13 16 9 0 15 13 1 9 7 13 13 1 9 0 9 0 14 9 13 7 13 2
6 3 16 3 13 9 2
12 3 13 3 7 3 9 0 9 14 9 13 2
15 9 15 1 9 15 3 9 9 0 16 3 13 1 15 2
25 2 9 9 12 1 9 15 14 9 2 11 10 9 2 0 13 1 9 2 9 16 1 10 15 2
6 9 3 13 1 15 2
33 9 13 16 1 9 9 15 15 3 13 9 16 3 13 9 1 10 9 2 7 1 9 9 15 13 13 9 15 1 9 0 2 2
22 3 7 13 9 9 13 3 2 7 3 2 3 0 1 10 9 7 13 1 10 11 2
5 7 13 7 13 2
1 2
4 9 9 0 2
1 2
3 3 3 2
33 7 3 2 1 3 13 3 16 13 1 10 9 2 13 9 16 1 15 3 13 10 9 1 9 15 9 0 13 14 9 10 9 2
15 11 2 11 2 9 2 9 2 7 3 9 10 9 0 2
25 7 1 10 9 14 9 0 2 7 1 9 2 9 1 10 9 10 0 14 9 10 9 10 0 2
2 3 2
11 10 9 13 1 10 9 10 0 10 15 2
16 13 9 16 13 3 15 9 0 14 10 9 1 9 10 9 2
15 16 7 2 7 7 1 9 9 3 4 3 13 3 13 2
15 10 9 15 13 3 9 0 0 7 0 2 9 13 9 2
16 3 2 4 13 9 1 9 7 13 2 3 13 3 7 3 2
19 1 9 9 15 13 16 0 7 13 13 9 2 7 13 7 13 13 9 2
17 3 1 15 13 16 0 13 3 9 2 7 13 7 13 13 9 2
4 7 9 3 2
7 3 13 9 2 13 0 2
3 13 13 2
9 13 9 2 9 2 9 2 9 2
4 7 3 3 2
31 16 7 10 9 10 0 16 13 1 9 10 9 3 13 13 1 15 3 14 10 9 10 0 1 9 1 9 15 10 0 2
8 3 3 13 2 1 10 9 2
23 7 7 3 13 1 10 9 2 3 9 15 10 0 14 10 9 1 10 9 13 9 0 2
13 9 3 13 16 10 11 13 1 15 14 10 9 2
14 1 9 15 13 1 9 15 9 7 9 1 10 9 2
6 0 2 0 7 0 2
32 9 7 9 9 13 13 9 13 7 9 0 7 0 1 9 10 9 1 10 9 1 9 15 2 1 10 9 10 0 10 15 2
50 15 13 1 15 9 1 9 15 14 10 9 2 9 1 9 15 1 9 15 10 0 2 9 1 9 15 1 15 16 13 1 9 2 10 9 7 13 1 15 2 7 3 3 7 3 9 0 7 0 2
17 9 0 7 0 9 0 1 9 0 7 13 1 9 15 16 13 2
28 7 3 1 15 13 1 15 16 15 3 3 13 1 9 0 9 2 7 13 1 15 14 10 9 3 1 9 2
24 3 10 9 16 13 1 10 9 10 11 2 11 2 0 10 15 16 10 9 13 1 15 3 2
36 2 13 16 1 9 0 2 3 1 16 13 9 15 14 3 9 0 2 4 3 13 14 9 9 15 10 0 14 10 9 2 0 2 15 2 2
2 2 2
39 10 9 10 3 2 13 13 2 1 10 10 9 2 3 15 2 7 9 0 13 16 10 9 13 2 7 10 9 10 0 10 15 13 16 15 3 3 13 2
8 15 3 3 3 13 14 15 2
6 3 3 9 2 9 2
8 3 13 1 15 1 10 9 2
5 4 13 14 15 2
56 9 10 9 10 0 11 11 2 9 15 10 0 14 9 9 2 13 13 1 10 9 10 0 14 10 9 1 12 10 9 10 0 14 12 2 1 9 15 10 0 14 9 10 9 1 9 11 1 10 9 10 9 11 1 11 2
17 9 10 9 13 13 9 9 16 13 1 10 9 10 0 1 15 2
29 11 13 13 1 10 9 1 9 16 10 9 0 3 7 13 13 14 10 9 16 13 1 15 16 13 14 10 9 2
6 15 13 13 2 13 2
30 15 13 1 10 9 1 10 9 2 1 15 13 9 12 12 9 2 7 13 1 10 9 9 10 9 13 1 9 15 2
19 11 13 13 1 15 3 13 14 10 9 10 0 14 10 9 1 10 9 2
18 9 9 2 16 13 13 1 9 15 1 9 10 9 2 13 1 9 2
31 1 9 15 14 9 2 1 9 13 2 13 1 9 10 9 10 0 7 1 9 15 10 0 1 9 9 10 9 9 15 2
29 1 2 9 9 9 15 14 9 1 11 12 4 11 2 1 9 11 2 13 12 12 9 1 12 9 1 9 9 2
33 12 9 1 9 15 13 1 13 2 7 3 12 12 1 9 3 2 0 1 9 2 14 10 0 16 1 15 1 10 12 1 11 2
35 1 9 9 7 9 15 14 11 1 3 2 9 10 9 16 13 1 15 14 13 14 10 9 2 13 9 16 15 13 13 14 9 10 9 2
40 9 10 9 14 9 13 1 9 15 10 0 14 11 11 2 9 7 9 9 10 9 10 0 14 9 11 10 0 2 1 9 9 7 9 14 9 10 9 9 2
26 11 2 16 9 9 15 10 0 13 1 11 2 13 14 9 15 1 9 3 1 9 15 1 9 11 2
46 1 9 13 16 1 10 9 10 0 13 11 14 9 10 9 16 1 9 15 1 9 2 16 13 3 1 9 10 9 16 13 1 10 9 10 0 1 9 10 9 1 10 9 1 11 2
39 11 15 13 16 13 9 9 9 2 11 11 2 13 3 1 10 9 10 0 10 0 14 10 9 2 3 9 10 9 2 10 9 2 10 9 7 10 9 2
31 1 15 13 11 1 9 15 13 3 9 0 2 16 13 0 1 9 9 10 9 1 10 9 1 9 2 7 1 9 15 2
11 1 3 13 14 9 15 11 11 2 11 2
32 1 9 13 16 11 2 11 2 16 15 9 1 9 10 9 14 9 2 13 13 9 1 9 10 9 1 10 9 14 10 9 2
21 1 9 11 12 9 12 9 7 12 9 16 13 1 10 9 10 0 1 10 9 2
17 1 0 1 10 9 2 13 10 9 1 15 9 1 9 9 13 2
16 9 10 9 1 10 9 13 1 9 2 9 14 12 9 0 2
18 9 10 9 7 10 10 9 10 0 13 13 1 9 11 15 9 0 2
14 10 10 9 13 1 9 10 9 7 10 9 9 0 2
35 1 10 9 2 1 10 9 7 1 10 0 2 16 13 13 1 9 10 9 2 13 3 4 13 2 7 0 9 16 13 13 1 9 0 2
32 2 10 9 10 0 2 3 14 10 0 2 9 12 9 1 9 1 11 2 13 9 1 10 9 10 0 1 10 12 1 11 2
45 3 2 1 9 10 0 2 13 10 9 10 0 9 12 14 9 10 9 1 2 11 2 2 13 16 9 15 13 1 9 11 7 13 13 1 10 9 10 0 1 12 12 10 0 2
36 1 9 1 9 12 12 9 2 12 12 9 1 9 10 9 10 0 2 13 10 9 10 0 13 9 14 9 2 16 13 14 9 15 10 0 2
39 2 15 13 13 1 9 10 9 16 9 1 9 10 9 2 7 1 9 9 10 11 9 2 1 11 2 2 13 11 11 2 9 15 14 10 9 10 0 2
11 1 10 9 13 4 3 13 14 10 9 2
18 1 9 10 9 13 9 12 9 2 13 11 2 10 0 16 1 15 2
12 1 10 9 13 9 0 16 13 2 0 2 2
21 15 13 1 10 15 1 9 15 3 2 1 9 16 13 13 9 0 15 7 0 2
15 7 3 2 16 13 9 15 14 11 2 13 9 0 3 2
27 10 9 10 0 15 13 9 9 2 0 2 7 11 13 9 1 9 13 14 9 0 1 10 9 10 0 2
16 9 0 13 9 12 2 9 13 1 9 13 9 0 7 3 2
30 9 11 2 11 11 2 13 16 15 13 1 10 9 1 9 0 7 13 9 0 0 7 0 1 9 10 9 10 0 2
24 7 10 9 4 13 0 1 9 12 9 1 9 0 2 1 1 10 9 7 1 1 10 9 2
32 16 16 13 9 0 1 10 9 10 3 0 2 11 2 2 2 3 16 11 13 1 11 2 10 9 10 0 13 1 11 2 2
11 10 9 1 11 1 10 0 13 0 9 2
34 9 10 9 14 11 13 1 10 12 10 12 1 10 9 10 0 3 7 9 15 14 11 9 7 10 9 10 0 2 10 0 14 15 2
43 1 9 10 9 1 11 13 10 10 9 2 1 9 1 11 1 1 10 9 10 0 2 2 0 2 2 7 1 9 9 0 2 2 1 9 10 9 13 3 9 0 2 2
13 10 10 9 1 11 13 0 9 14 12 9 9 2
11 9 10 9 13 1 11 10 0 1 12 2
20 1 10 12 1 11 3 13 10 0 9 15 1 9 0 14 12 9 1 11 2
13 9 13 9 1 10 9 7 9 13 2 11 0 2
25 2 10 9 14 15 3 3 13 9 0 2 2 13 10 9 11 11 2 2 10 9 13 0 2 2
30 10 9 0 10 9 14 10 9 10 0 2 10 0 13 15 3 1 9 10 11 10 0 2 16 13 9 2 1 11 2
19 7 1 9 10 9 13 9 7 9 1 9 9 0 1 10 12 10 12 2
24 2 10 9 14 15 3 0 3 2 7 10 9 14 15 0 3 2 2 13 10 9 11 11 2
20 9 10 9 10 0 13 3 13 14 10 9 10 0 1 2 9 9 10 9 2
8 7 13 16 10 9 13 0 2
35 9 0 13 3 13 9 2 9 0 3 1 10 9 10 0 2 13 9 0 1 10 9 7 13 14 9 11 1 9 11 1 9 10 9 2
47 15 13 13 14 12 10 0 16 13 1 9 1 10 9 1 11 2 1 11 2 1 9 11 7 1 11 2 3 13 3 1 12 12 0 2 2 1 13 14 9 15 14 10 9 10 0 2
38 2 15 4 13 10 9 1 10 9 1 10 9 2 2 13 11 11 1 9 10 9 10 0 2 11 2 2 16 13 16 2 4 3 16 9 13 2 2
21 9 13 1 9 9 2 7 3 9 13 1 9 9 0 3 7 1 9 0 3 2
34 1 9 9 9 0 2 9 1 9 0 13 1 10 9 16 13 9 14 12 12 9 2 12 12 9 2 2 16 14 9 3 13 11 2
14 11 13 1 9 1 12 12 9 1 9 9 10 9 2
23 2 1 12 9 3 13 1 9 2 2 13 11 11 2 9 9 9 9 10 9 10 0 2
19 2 15 13 13 14 9 15 1 2 9 9 9 0 3 1 9 15 2 2
47 9 15 13 0 2 11 13 9 10 9 10 12 1 9 15 1 9 10 9 7 13 1 15 9 9 0 2 1 9 10 9 14 11 2 16 13 12 9 1 9 10 9 14 9 10 9 2
25 10 9 10 0 13 13 14 11 13 1 9 15 14 10 9 1 9 10 9 1 9 1 9 9 2
10 9 0 15 13 1 9 1 9 9 2
25 9 0 2 0 7 9 1 12 2 13 16 1 10 9 10 0 3 13 10 9 1 9 9 0 2
13 15 13 16 1 9 10 9 13 7 9 0 12 2
12 2 9 13 1 10 9 7 13 1 9 0 2
24 7 10 12 13 13 3 13 15 2 2 13 11 11 2 9 10 9 10 0 2 11 11 2 2
8 2 10 12 3 13 1 15 2
7 13 1 15 10 9 2 2
20 9 0 13 16 1 15 13 1 9 1 11 1 16 4 13 13 14 10 9 2
9 7 0 13 16 15 3 10 9 2
30 9 13 9 9 0 3 7 9 9 0 0 3 2 7 7 10 9 3 3 13 14 10 9 1 9 10 9 10 0 2
25 2 15 13 13 9 1 10 9 1 13 1 9 2 2 13 11 11 2 9 9 0 0 1 11 2
16 10 9 15 9 10 9 16 13 10 0 1 11 13 3 0 2
22 11 0 13 1 9 0 0 1 11 2 1 3 1 9 0 1 11 2 7 13 13 2
14 13 9 1 15 16 9 3 15 3 4 1 10 9 2
18 2 15 9 0 3 2 2 13 11 11 2 9 1 10 9 10 0 2
20 2 15 10 3 4 1 16 9 13 13 13 1 10 9 7 13 1 15 2 2
13 9 9 0 13 16 9 3 13 1 15 3 9 2
26 2 15 13 14 10 9 14 15 2 2 13 11 11 2 9 9 9 9 10 9 1 10 9 10 0 2
16 2 7 15 3 13 3 13 1 15 14 10 9 14 15 2 2
15 9 3 13 1 9 9 16 13 1 9 0 16 13 9 2
24 10 9 1 11 13 1 9 9 1 9 0 16 13 14 10 9 1 9 0 12 1 10 9 2
19 2 3 9 13 1 10 9 14 15 1 9 1 10 9 0 1 10 9 2
11 2 13 11 11 2 9 9 0 1 11 2
10 2 13 10 9 13 1 15 9 2 2
13 9 15 14 11 13 3 1 9 0 1 11 11 2
16 13 16 9 0 13 16 15 13 1 9 15 14 9 10 9 2
22 16 13 1 11 1 11 2 13 11 2 2 15 13 1 15 13 10 16 15 4 2 2
9 9 0 0 13 9 15 1 0 2
11 2 11 13 3 9 2 2 13 11 11 2
15 2 15 13 1 15 3 15 9 7 1 3 15 13 2 2
36 10 3 11 13 1 11 1 9 0 3 1 11 2 7 10 9 13 16 13 1 9 0 3 1 9 15 14 15 7 9 15 4 13 9 0 2
25 2 1 12 9 13 11 9 16 9 15 13 9 2 2 13 9 10 9 14 9 11 2 11 11 2
10 2 10 9 13 7 13 13 1 9 2
23 10 9 13 1 15 9 4 9 13 2 2 7 1 15 9 13 10 9 3 14 9 11 2
21 13 1 15 9 1 16 9 0 15 13 13 2 7 3 3 15 13 1 9 0 2
20 7 2 16 16 15 9 0 3 2 4 1 9 0 13 1 9 15 10 0 2
31 10 9 2 16 13 1 9 2 13 12 9 16 13 9 1 9 0 12 2 7 15 13 13 1 15 1 10 9 10 9 2
32 10 9 13 1 12 9 7 12 9 2 9 0 7 0 7 9 9 9 2 9 16 13 9 1 10 9 10 0 14 10 9 2
20 10 9 0 1 11 2 7 16 10 9 13 13 1 15 11 2 9 15 3 2
17 15 13 1 10 9 1 9 9 1 9 11 2 3 1 9 11 2
38 1 16 11 3 13 16 15 0 9 0 2 13 11 1 10 9 14 11 16 1 15 13 9 15 1 10 9 2 11 1 16 13 1 9 15 10 0 2
26 10 9 10 12 1 9 9 15 13 11 2 9 15 14 11 2 16 3 13 9 1 11 1 9 15 2
2 0 2
4 3 10 3 2
10 7 3 3 3 1 9 15 14 9 2
13 4 13 1 10 9 7 11 7 11 13 13 3 2
14 7 13 1 10 9 9 0 16 13 1 9 0 15 2
32 10 9 0 1 9 0 14 9 7 9 16 13 9 14 9 1 9 12 2 13 1 15 7 13 1 15 3 1 9 0 0 2
40 9 9 7 9 15 13 3 1 9 0 14 9 7 9 2 7 7 15 4 13 1 10 9 16 1 10 9 10 15 3 13 1 11 2 11 7 9 0 0 2
38 3 16 13 14 10 9 13 10 9 16 1 9 15 10 3 2 0 15 2 1 10 15 2 9 0 2 7 10 9 10 0 13 1 15 1 9 0 2
44 3 16 10 9 13 9 2 16 3 11 11 3 13 13 13 0 1 15 2 10 9 10 0 13 1 15 9 14 9 7 9 16 13 14 15 1 0 3 1 3 16 15 3 2
30 10 9 0 3 1 9 10 9 2 11 9 11 2 16 13 14 11 2 7 11 11 2 16 13 14 9 15 14 11 2
24 11 13 9 14 9 0 0 7 0 2 1 10 15 16 13 1 10 9 11 11 7 11 11 2
23 14 10 9 13 11 11 2 9 15 14 10 9 10 0 11 11 2 16 13 1 9 0 2
33 15 9 15 10 0 1 9 2 7 13 9 0 1 10 9 16 15 13 13 14 10 9 14 15 1 9 0 7 0 1 9 15 2
29 13 1 10 9 9 14 9 7 9 2 7 2 15 13 9 0 3 2 7 15 13 13 1 15 7 1 9 15 2
35 9 11 13 1 9 11 1 10 9 1 9 9 11 2 11 2 12 9 3 1 9 10 9 1 9 11 2 1 9 9 1 9 10 11 2
38 9 11 13 1 9 1 9 15 1 16 13 1 9 0 7 1 9 14 9 1 9 10 11 16 13 3 3 1 10 9 16 1 9 1 9 10 9 2
11 10 9 13 9 9 2 9 7 9 11 2
21 15 13 1 10 9 11 2 11 7 11 9 2 11 9 2 12 9 3 1 11 2
25 1 9 10 9 13 7 13 10 9 16 13 14 10 9 1 9 1 9 1 9 11 7 1 11 2
26 9 11 13 1 9 9 0 3 2 1 9 9 0 7 1 9 14 12 9 3 0 1 9 10 9 2
32 9 0 13 16 10 9 1 10 9 13 1 9 9 1 9 0 3 1 11 2 9 10 9 7 9 1 9 9 1 9 12 2
34 8 8 8 13 16 9 11 13 10 10 9 7 13 9 9 16 13 14 9 11 1 9 9 7 9 1 11 7 9 1 9 10 9 2
30 10 9 13 16 10 9 13 9 1 9 11 1 10 9 13 1 9 0 0 1 9 14 9 1 9 1 9 10 9 2
34 9 11 13 1 9 10 9 16 9 10 9 10 0 11 13 1 11 1 9 11 1 13 1 9 10 9 10 0 11 13 1 9 11 2
26 9 10 9 11 11 13 1 9 11 1 9 10 9 1 11 7 13 14 10 9 10 0 1 9 9 2
20 9 10 9 13 9 1 10 9 2 1 15 3 1 9 9 10 9 11 11 2
46 1 9 10 9 16 13 13 9 0 0 1 9 10 9 16 10 9 10 0 11 2 16 1 9 1 9 10 9 2 13 9 0 7 4 16 10 9 1 15 13 1 9 9 9 11 2
25 10 9 1 11 13 16 9 11 10 3 2 0 13 13 9 14 9 0 1 10 9 1 9 11 2
31 3 9 11 11 2 9 9 2 13 16 1 10 9 10 0 10 3 13 9 0 15 13 1 10 9 14 9 0 1 11 2
33 9 11 13 16 1 10 16 13 1 15 2 13 9 1 11 1 9 10 9 7 15 13 4 13 9 0 1 10 15 1 9 11 2
40 9 0 1 11 13 14 10 9 16 13 1 11 2 7 1 9 16 13 1 10 9 1 9 16 13 10 9 1 9 11 2 13 16 10 9 13 1 9 0 2
45 10 10 9 1 10 9 13 2 16 9 13 12 10 9 16 1 15 13 14 15 10 9 10 0 1 9 2 10 9 1 9 9 0 2 7 9 15 10 0 13 9 0 7 0 2
21 14 13 1 9 2 9 2 4 13 1 15 2 3 10 2 13 7 13 1 9 2
42 3 2 4 3 13 1 10 9 16 4 1 9 13 13 9 7 13 9 1 10 9 10 0 2 7 3 15 1 10 9 16 13 3 1 9 10 9 1 9 2 9 2
15 1 15 0 16 4 13 9 0 14 10 9 16 13 13 2
9 10 9 13 13 1 10 9 2 2
57 9 16 13 13 14 15 1 9 0 2 4 16 3 13 3 2 16 15 13 9 9 1 10 10 13 1 10 9 2 1 10 9 2 1 10 13 2 1 9 2 10 9 10 0 2 2 7 3 3 7 3 2 1 10 9 15 2
33 9 15 14 10 9 11 11 2 12 1 12 9 16 13 1 10 9 10 0 1 10 9 2 13 9 1 9 16 13 13 14 15 2
30 9 15 1 10 9 14 11 13 13 2 9 15 13 0 7 0 2 9 2 7 9 10 9 14 15 13 0 7 0 2
34 3 4 13 9 1 10 9 1 10 9 15 2 7 9 0 4 13 14 9 10 9 14 15 7 13 2 3 3 2 14 9 10 9 2
10 9 0 13 3 1 9 11 7 11 2
18 11 13 14 15 1 9 15 14 9 9 7 9 16 3 13 1 15 2
14 3 1 10 9 14 11 13 9 10 9 1 9 9 2
17 9 9 10 9 11 11 13 1 10 9 9 0 14 9 2 9 2
16 9 15 0 7 0 2 13 14 10 9 7 13 14 10 9 2
28 15 13 13 9 14 9 7 9 2 7 16 10 11 14 15 0 10 2 3 16 15 13 1 15 10 9 0 2
97 10 13 3 3 1 10 9 1 10 9 10 0 14 10 9 2 3 13 3 9 15 14 10 11 2 1 10 9 1 2 9 11 2 2 7 3 1 10 9 1 2 9 10 9 2 14 11 2 10 11 7 10 11 13 1 10 11 1 10 9 2 2 13 16 1 11 13 10 9 10 0 14 9 10 9 7 9 10 9 2 7 10 9 10 0 10 0 14 1 15 13 9 1 9 0 0 2
33 1 9 15 13 3 9 0 0 7 0 2 7 3 3 13 3 10 9 1 9 10 9 7 1 9 10 9 10 0 14 10 9 2
45 3 9 12 10 9 1 2 11 11 2 14 11 16 13 2 1 9 2 9 9 1 10 9 13 0 3 1 9 10 9 14 11 7 14 10 9 10 0 7 1 9 0 2 0 2
19 3 16 9 15 14 10 9 10 0 2 11 11 2 13 0 7 3 0 2
13 3 1 9 9 10 9 1 9 10 9 10 0 2
36 10 9 16 13 14 9 15 14 10 9 10 0 7 10 9 10 0 10 0 1 9 16 13 1 2 11 2 1 11 4 13 1 9 10 9 2
40 1 9 2 9 11 2 2 7 2 16 13 1 9 9 14 10 9 16 1 10 9 2 9 10 9 10 0 13 0 3 2 1 9 11 11 1 2 11 2 2
30 1 11 12 13 9 7 9 9 12 9 1 9 12 12 9 2 1 9 9 14 12 12 9 12 9 1 9 10 9 2
21 9 1 15 15 13 12 9 1 9 12 12 9 12 9 1 9 10 9 10 0 2
23 1 11 3 15 13 12 9 1 9 0 14 12 12 9 12 9 1 9 10 9 9 15 2
31 1 11 13 12 10 9 16 13 9 1 9 0 2 3 2 14 12 12 9 1 12 9 1 9 9 11 14 2 11 2 2
13 10 9 13 9 9 1 9 0 7 1 9 0 2
41 9 9 1 12 10 9 10 0 13 10 9 10 0 14 9 9 0 1 10 9 10 0 7 13 13 9 9 0 1 11 2 1 9 10 11 7 1 9 9 11 2
31 11 13 1 9 10 9 10 0 3 1 9 10 9 10 0 2 7 1 9 9 15 13 13 9 0 1 10 9 10 0 2
18 1 3 13 10 9 2 16 9 15 14 9 10 9 10 9 3 13 2
13 9 0 1 15 13 1 10 12 1 11 1 11 2
17 1 15 9 13 11 11 9 0 14 9 0 1 10 12 10 12 2
30 15 13 10 9 10 0 1 9 15 16 13 0 1 10 9 2 7 3 13 3 1 9 1 10 9 1 9 0 0 2
13 15 13 9 15 14 9 16 13 11 1 9 0 2
51 11 2 9 15 14 9 9 0 2 16 13 12 10 9 1 9 15 1 11 2 13 1 9 9 15 13 1 9 10 9 14 9 9 0 7 13 1 9 9 10 9 7 10 9 14 9 11 1 9 11 2
14 3 15 12 1 12 2 12 9 16 13 1 9 15 2
16 15 3 13 1 9 10 9 1 9 0 1 10 12 10 12 2
28 9 15 2 11 11 2 13 14 15 1 9 10 12 1 13 1 12 10 9 10 0 1 9 0 9 9 15 2
25 14 13 9 1 14 15 1 12 2 13 10 9 13 9 0 1 9 0 7 9 0 0 1 12 2
22 15 13 9 9 1 9 0 0 2 13 1 12 2 7 13 13 14 10 9 1 11 2
22 10 1 9 12 9 0 13 1 11 12 14 9 2 11 2 1 9 0 14 9 9 2
9 10 9 1 11 13 9 10 9 2
29 10 9 2 16 13 1 9 1 10 9 14 11 1 11 2 3 13 4 13 1 9 3 0 2 7 13 4 13 2
27 1 15 10 9 3 13 4 13 14 9 15 10 0 3 1 9 0 0 2 16 1 9 9 15 13 0 2
7 7 10 9 13 9 0 2
21 1 12 10 9 16 13 1 9 13 12 2 1 12 12 9 2 12 12 9 2 2
13 9 10 9 1 10 9 13 12 1 12 12 9 2
23 16 16 13 11 2 10 9 1 9 0 16 1 15 9 0 13 1 9 10 12 10 0 2
24 1 9 10 12 10 0 13 10 9 9 2 7 9 10 9 10 0 13 0 1 9 1 15 2
37 10 9 1 9 14 9 1 9 0 13 16 13 14 10 9 14 10 9 2 10 9 7 10 9 10 0 14 10 12 10 12 1 10 9 10 0 2
35 7 13 10 9 1 11 2 1 9 0 2 9 1 10 16 13 1 9 16 13 10 9 1 9 9 0 1 10 12 10 12 7 10 12 2
17 9 10 9 13 1 9 1 9 16 13 1 10 9 10 0 3 2
40 9 14 9 11 1 11 11 2 16 10 9 14 15 13 14 9 15 1 9 10 9 10 0 2 13 1 12 12 9 1 1 10 9 10 0 14 12 12 9 2
16 9 0 13 3 1 2 11 14 11 2 1 11 2 1 12 2
25 9 15 2 16 13 13 0 3 1 9 0 2 13 1 12 12 9 12 9 1 10 9 10 0 2
23 1 10 9 16 13 13 10 9 1 11 2 11 14 9 15 13 7 13 9 1 9 9 2
54 1 9 0 14 2 11 2 1 10 12 1 11 13 11 2 10 9 10 13 1 9 14 9 0 0 1 11 2 12 9 9 16 0 3 3 12 1 10 9 10 0 1 9 1 9 1 10 12 10 12 7 10 12 2
34 10 9 13 3 13 1 9 10 9 10 0 1 10 9 10 0 2 16 16 13 1 15 10 9 1 9 10 12 1 9 9 10 12 2
45 1 9 12 15 13 14 10 9 10 0 3 2 7 1 9 0 13 13 1 10 9 10 0 14 9 0 2 16 9 0 14 9 9 0 1 9 15 4 1 9 9 1 10 9 2
36 7 4 13 2 16 9 0 0 16 15 2 7 2 3 0 2 7 9 9 15 14 9 0 1 11 2 9 2 11 7 11 3 13 1 9 2
30 1 10 9 10 0 3 13 11 13 1 9 16 13 1 10 9 7 1 15 2 7 16 9 9 15 3 4 1 9 2
31 1 9 9 9 9 15 13 10 9 13 13 9 9 9 0 2 13 9 14 15 16 13 1 0 3 2 7 3 13 9 2
29 1 9 11 9 1 2 11 2 2 9 9 0 13 1 11 1 9 0 7 1 9 0 1 16 16 13 1 3 2
29 9 10 9 7 10 9 2 11 11 2 13 13 1 9 9 10 9 1 10 9 10 0 2 3 10 9 10 0 2
18 11 13 14 10 9 1 9 16 13 1 9 10 9 1 9 9 11 2
40 1 9 10 9 2 10 9 16 13 1 9 0 1 9 9 15 1 9 10 9 1 10 9 13 3 3 1 9 9 9 0 2 7 3 1 9 14 9 0 2
43 11 13 3 16 15 13 1 9 9 9 0 2 16 13 1 9 9 1 10 9 16 10 9 13 9 0 14 10 9 2 7 13 9 16 3 13 1 10 9 1 9 15 2
31 15 9 13 1 10 9 1 9 2 16 1 15 13 10 9 10 0 1 0 7 13 3 14 10 9 10 0 14 10 9 2
26 9 13 9 10 9 1 10 3 16 13 1 9 14 9 10 9 13 1 9 9 10 9 7 10 9 2
47 3 2 14 13 9 11 1 9 9 0 1 9 10 9 2 1 9 0 1 9 10 9 7 9 15 10 0 1 9 9 10 9 2 13 1 10 9 7 9 15 13 14 10 9 10 0 2
76 1 9 0 16 1 15 13 9 15 14 9 10 9 2 11 11 2 7 3 9 10 9 2 11 9 2 3 13 9 2 7 14 13 10 9 16 13 13 9 0 2 3 13 1 15 9 9 11 7 9 15 9 0 13 9 2 16 10 12 13 13 15 15 9 0 2 9 1 9 9 15 7 1 9 15 2
41 7 9 10 9 1 9 10 9 2 13 9 16 9 9 11 2 7 9 10 9 10 0 14 9 10 9 2 3 13 13 1 9 16 1 10 15 1 9 10 9 2
42 1 9 10 9 13 16 13 2 16 9 9 15 14 9 11 13 1 9 2 7 16 1 10 9 9 15 13 3 1 9 9 9 9 7 9 2 9 16 3 3 13 2
50 11 2 1 15 2 13 16 13 1 9 9 1 10 15 3 1 13 9 16 13 1 15 15 9 3 2 15 13 7 7 13 13 9 0 0 2 7 15 12 10 9 16 1 15 4 13 14 9 15 2
74 10 9 1 9 9 0 1 10 9 1 9 10 9 2 9 9 11 7 9 9 1 9 15 2 9 15 10 0 14 9 10 9 10 0 2 9 11 11 2 7 3 9 15 10 0 1 9 14 9 9 9 9 2 9 11 9 2 10 15 13 1 10 9 10 0 1 9 9 0 9 1 10 9 2
25 1 9 9 0 2 1 12 9 0 1 9 9 2 9 7 3 13 1 10 9 7 1 10 9 2
16 9 10 9 13 1 10 9 10 0 1 9 0 9 9 0 2
18 9 13 3 1 9 10 9 7 13 1 9 0 1 9 1 10 9 2
32 3 3 13 1 10 9 2 16 16 3 13 3 3 9 15 1 10 9 2 16 13 1 9 9 1 9 10 9 14 10 9 2
9 10 9 10 15 9 13 13 9 2
14 15 13 13 16 10 9 16 13 1 15 0 7 0 2
17 9 9 0 1 9 1 10 15 3 13 1 10 9 15 9 0 2
25 7 13 9 16 10 9 7 10 9 13 2 1 9 7 9 7 7 9 9 14 9 7 9 9 2
19 10 9 1 10 9 13 3 9 0 7 9 14 9 13 9 15 14 0 2
30 3 9 10 9 7 3 10 9 0 1 10 9 10 3 2 0 10 15 7 13 16 3 1 1 9 13 1 10 9 2
47 9 10 9 10 0 1 10 9 13 1 10 9 1 9 9 9 11 10 0 2 9 0 2 0 7 0 3 2 16 10 9 1 15 0 7 16 13 9 9 1 10 9 7 1 10 9 2
85 13 1 9 1 9 15 9 9 10 9 2 9 11 11 2 9 9 10 9 10 0 2 9 11 11 2 9 9 10 9 2 9 11 11 2 9 9 9 9 2 9 2 9 11 11 2 7 9 9 10 9 1 9 14 10 9 2 9 11 11 9 2 16 1 1 1 9 13 1 9 9 10 9 7 16 13 1 15 9 0 0 1 10 9 2
47 3 1 10 9 10 15 16 3 13 1 10 9 2 0 9 15 13 1 12 10 9 10 0 10 0 2 1 9 10 9 10 0 2 9 9 10 9 2 7 9 10 9 14 9 10 9 2
45 1 9 15 13 1 9 10 9 1 10 9 10 0 14 10 9 1 9 9 15 14 9 11 10 0 2 3 1 9 10 9 10 0 7 3 1 9 9 9 10 9 7 10 9 2
15 1 10 9 10 13 2 9 11 13 1 9 11 10 0 2
18 10 9 14 10 9 13 1 9 10 9 10 0 2 1 9 10 9 2
10 4 16 13 1 10 9 3 9 11 2
59 10 9 9 13 1 9 0 2 3 15 1 10 9 10 0 7 9 10 9 2 1 9 9 0 2 3 1 9 9 2 9 2 2 13 9 10 9 10 0 3 2 1 10 9 0 2 7 1 15 9 0 7 9 0 2 10 9 2 2
79 1 9 10 9 13 14 10 9 13 10 9 2 16 9 10 9 1 11 7 9 10 9 7 9 15 2 3 1 9 3 2 0 2 13 9 16 13 9 14 9 0 7 0 14 9 7 9 10 9 1 10 9 2 1 9 15 14 9 0 7 0 1 9 9 2 16 3 1 9 15 13 13 10 9 15 1 9 11 2
25 1 3 13 11 0 1 10 9 10 0 2 16 13 1 11 1 10 9 7 1 11 1 10 9 2
29 1 9 10 9 10 0 10 0 2 10 9 10 0 13 1 9 10 9 3 2 7 9 15 13 1 9 2 12 2
32 1 10 9 7 7 1 9 10 9 13 13 16 13 2 16 9 9 11 1 10 9 10 0 2 13 7 1 9 9 0 3 2
49 13 16 1 10 9 16 13 2 16 1 15 13 10 9 1 9 10 9 1 9 9 11 2 1 9 9 15 14 10 9 11 2 16 13 1 9 0 2 3 10 9 9 3 13 13 1 10 9 2
34 13 16 13 1 10 9 10 0 2 3 1 13 16 10 9 13 9 1 9 9 10 9 7 3 3 1 13 9 9 0 1 10 9 2
49 16 13 14 9 10 9 10 0 13 2 16 7 3 13 3 10 12 9 0 1 10 9 7 3 9 0 14 9 7 9 2 1 9 11 1 9 9 2 3 13 10 9 1 9 10 9 10 0 2
11 15 9 0 13 10 9 9 9 7 9 2
20 10 9 13 9 1 10 15 1 10 9 2 7 10 9 3 13 1 10 9 2
27 3 2 1 10 9 1 9 10 9 10 0 2 13 9 10 9 16 13 1 11 12 9 0 1 9 9 2
15 7 7 2 9 15 14 15 1 15 13 1 15 10 9 2
41 1 9 9 10 9 10 0 2 11 11 2 13 9 11 2 1 3 9 10 9 2 1 9 0 1 12 9 2 16 13 1 9 9 1 10 10 9 1 10 9 2
10 9 9 15 13 2 1 9 3 2 2
29 9 1 9 12 9 1 10 9 14 9 11 2 1 9 9 10 9 10 0 1 10 9 2 13 3 9 0 3 2
27 15 7 3 2 9 10 9 13 9 16 9 1 10 9 10 9 13 1 15 2 7 1 9 0 14 9 2
24 9 9 10 9 10 0 1 9 15 2 15 13 2 13 1 9 10 9 1 10 9 10 9 2
32 10 9 9 13 2 16 7 3 13 9 0 2 13 9 14 9 10 9 2 16 13 1 10 9 1 9 11 2 1 9 11 2
31 10 9 13 2 16 13 1 15 9 13 15 1 9 15 7 16 10 9 13 1 9 10 9 7 3 1 9 9 10 9 2
26 1 10 9 2 1 9 9 2 1 9 9 10 0 1 10 9 2 4 9 15 14 10 9 13 9 2
24 10 9 13 2 16 1 9 9 11 1 9 10 9 1 11 2 3 3 13 10 9 9 9 2
52 9 11 3 13 2 3 2 13 1 9 10 9 9 0 14 9 9 2 16 13 1 10 9 13 14 9 15 10 0 1 10 9 2 1 0 1 10 9 16 13 1 9 15 1 9 10 9 1 9 10 9 2
19 1 9 15 13 9 11 1 10 9 10 0 15 9 0 1 9 10 9 2
25 13 1 9 9 0 2 16 13 3 1 9 1 9 0 2 1 9 7 1 9 1 9 10 9 2
43 3 13 1 9 9 7 9 0 1 10 9 7 3 1 9 1 10 9 10 0 14 15 7 1 10 9 1 15 2 7 1 9 0 2 0 7 0 14 10 9 10 0 2
38 9 0 4 13 1 9 0 14 9 10 9 2 13 1 10 9 7 13 1 10 9 16 13 9 0 1 9 15 7 3 13 1 15 13 9 0 3 2
62 3 1 11 12 13 9 9 10 9 2 11 11 2 9 2 16 13 1 9 1 9 9 10 9 7 9 9 7 9 0 2 7 1 15 13 1 9 1 9 15 14 9 10 9 1 2 9 9 0 16 13 1 9 10 9 7 9 9 10 9 2 2
52 1 9 16 9 15 2 2 9 10 9 9 10 9 2 10 9 7 10 9 2 2 13 10 9 2 1 10 9 2 3 14 10 9 16 1 9 15 13 9 11 13 14 9 10 9 10 0 1 9 10 9 2
34 2 4 13 16 10 9 14 9 9 0 16 13 1 15 2 4 13 1 9 9 1 9 3 1 9 0 0 2 2 13 1 10 9 2
41 1 10 9 14 9 10 9 13 10 9 14 9 10 9 14 10 9 7 9 9 10 9 1 9 9 7 9 9 0 14 9 9 2 9 15 7 9 1 9 15 2
18 10 9 13 3 14 10 9 14 9 9 7 9 9 1 9 10 9 2
64 15 13 1 9 16 13 1 9 10 9 7 1 9 10 9 1 9 9 15 10 0 2 2 9 10 9 2 1 9 9 0 7 9 14 9 10 9 2 4 13 9 15 1 10 9 14 12 9 0 2 9 7 9 2 9 9 2 9 0 7 9 0 0 2
66 1 9 9 15 1 10 9 13 7 13 1 10 9 10 0 3 12 9 0 2 16 13 12 1 10 9 2 1 10 9 10 0 2 11 2 9 7 9 1 9 9 2 11 2 9 7 9 1 9 10 9 7 9 9 13 2 11 2 9 9 9 7 9 9 0 2
11 9 0 3 1 9 9 9 13 10 9 2
18 1 9 0 2 9 15 14 10 9 13 1 9 0 14 9 10 9 2
14 2 9 0 13 9 0 0 7 13 1 9 10 9 2
19 9 0 1 10 9 4 13 1 12 9 2 0 2 0 2 13 7 0 2
39 1 10 9 10 15 2 16 13 9 9 10 9 1 9 2 13 3 1 9 1 9 7 9 1 10 16 13 1 9 10 9 1 10 9 1 9 10 9 2
64 1 9 10 9 13 9 2 16 9 9 0 13 9 2 3 13 9 0 7 13 2 3 3 1 9 9 0 1 10 9 14 9 10 9 16 13 2 7 13 13 1 10 9 10 0 2 1 10 9 1 9 14 9 10 9 1 9 15 10 0 14 10 9 2
12 9 9 0 1 9 10 9 4 13 9 15 2
25 3 3 16 9 11 13 1 9 10 9 9 13 1 9 0 0 2 9 16 3 13 0 1 3 2
26 1 9 15 13 9 10 9 1 9 0 2 3 1 9 9 15 2 1 9 1 9 10 9 10 15 2
20 1 9 10 9 10 13 2 13 10 9 10 0 14 10 9 12 2 12 9 2
44 9 12 2 1 9 3 2 9 2 13 9 9 0 1 9 10 9 2 10 9 7 10 9 2 7 9 0 2 1 9 9 2 9 2 13 9 9 7 9 1 9 10 9 2
19 1 9 15 3 9 10 9 13 13 1 10 9 14 15 1 9 10 9 2
46 1 10 9 10 0 3 13 9 10 9 1 12 9 9 0 7 0 3 1 9 9 9 2 1 9 9 10 9 14 9 10 9 2 1 10 9 13 14 9 10 9 10 0 14 15 2
18 1 10 9 2 3 2 13 1 9 2 0 2 1 1 9 10 9 2
24 1 9 10 9 13 16 10 9 10 0 16 13 1 10 9 3 13 1 10 9 1 10 9 2
32 1 10 9 2 1 16 13 10 9 10 0 3 3 13 1 9 10 9 9 1 9 1 10 9 7 1 10 9 14 10 9 2
35 10 9 16 13 9 9 1 10 9 1 9 9 10 9 2 1 9 9 0 7 3 9 9 1 9 10 9 10 0 2 3 3 13 0 2
36 9 1 9 10 9 10 0 2 13 9 9 10 9 10 0 9 16 13 14 10 9 10 0 2 1 9 15 2 1 9 15 1 9 10 9 2
66 1 10 9 13 1 10 9 9 10 9 11 11 2 7 9 15 11 11 2 16 2 9 2 10 9 13 1 12 1 12 9 2 10 9 13 1 1 12 9 1 10 9 16 1 15 13 10 9 1 9 15 2 7 16 10 9 10 0 14 10 9 13 1 12 9 2
61 4 13 1 9 10 9 10 15 2 16 7 9 15 10 0 13 13 9 1 10 9 7 13 1 15 1 10 9 2 7 3 1 10 9 16 4 13 1 10 9 10 0 1 9 10 9 1 9 9 2 16 1 9 15 13 10 9 1 9 11 2
21 7 9 10 9 14 10 9 13 13 7 13 13 1 10 9 10 0 14 10 9 2
22 9 10 9 1 11 13 1 9 9 2 16 9 7 13 1 15 1 15 9 0 0 2
35 10 9 15 13 1 9 0 2 16 1 15 13 9 11 1 9 10 9 1 10 9 14 10 9 10 0 1 9 1 10 9 14 10 9 2
31 9 1 9 15 13 15 1 3 2 1 9 2 9 2 10 9 10 0 2 14 9 10 9 7 9 9 10 13 10 0 2
30 7 1 9 10 9 13 10 9 1 9 15 7 11 11 2 11 11 7 11 11 10 0 2 3 13 14 9 10 9 2
66 3 15 3 16 10 9 10 0 14 9 10 9 1 9 9 15 1 9 9 14 10 9 13 1 10 9 1 9 15 15 13 0 1 9 9 0 0 7 16 10 9 10 13 1 15 1 9 9 15 0 1 10 9 0 16 13 1 13 9 9 0 2 7 12 9 2
14 15 9 3 0 1 10 9 0 0 7 3 2 0 2
26 16 16 9 9 10 9 13 1 9 10 9 10 0 2 15 13 3 3 1 9 9 10 9 10 0 2
42 3 15 9 13 9 9 16 9 15 13 1 9 9 0 1 12 9 2 0 1 12 9 2 13 9 14 12 9 2 16 0 3 15 1 12 9 7 13 1 10 9 2
63 1 9 11 2 9 15 2 3 10 12 4 13 9 9 2 10 3 16 13 13 9 16 13 14 9 10 9 2 9 16 13 7 13 1 15 14 10 9 1 10 9 2 7 10 9 15 2 9 16 3 10 9 9 10 9 13 1 15 1 10 9 2 2
40 10 9 10 0 14 9 9 9 13 13 1 9 11 2 11 7 9 15 2 13 14 9 10 9 1 9 0 1 9 0 14 9 10 9 1 9 9 0 0 2
45 7 13 10 9 10 13 1 9 9 10 9 7 13 1 10 9 10 0 9 2 4 16 9 10 9 13 13 7 13 9 0 16 13 14 10 9 1 9 16 13 1 9 10 9 2
20 15 2 1 13 14 9 10 9 1 12 9 7 13 14 9 15 1 12 9 2
24 9 9 0 1 10 15 13 9 0 0 14 10 9 10 0 1 10 9 1 10 9 10 13 2
57 1 1 9 13 9 10 9 10 0 9 0 2 16 1 15 7 9 13 1 9 10 9 7 13 9 15 9 2 13 9 16 13 3 1 10 15 1 9 1 9 9 10 9 2 7 1 10 9 1 10 9 2 0 1 10 9 2
39 1 9 9 16 13 1 9 14 12 9 1 12 2 13 16 10 9 10 0 13 7 10 9 13 7 7 13 1 10 9 2 1 1 9 7 1 1 9 2
12 10 9 13 14 10 9 10 0 2 9 2 2
27 7 9 10 9 2 11 11 2 13 14 10 9 10 15 2 7 13 16 3 1 9 15 10 9 1 15 2
33 11 13 16 1 9 9 10 12 13 9 10 9 14 9 15 2 7 10 9 13 1 9 9 0 1 10 9 7 1 9 10 9 2
17 1 10 9 10 15 2 13 3 10 9 14 9 7 9 1 9 2
45 13 10 9 16 13 1 15 1 9 10 9 1 9 16 13 1 9 15 1 10 9 2 7 16 13 14 10 9 2 7 13 0 16 15 13 3 1 9 15 14 10 9 10 0 2
46 10 9 13 2 3 0 2 0 2 10 9 13 1 10 9 1 9 15 1 9 10 9 7 13 1 9 10 9 2 7 7 10 9 16 1 15 13 4 13 13 7 13 1 9 0 2
42 9 10 9 13 1 9 15 14 10 9 16 1 15 3 9 4 13 9 1 9 15 14 10 9 1 9 15 1 10 9 2 7 15 13 14 9 15 1 9 10 9 2
50 1 13 14 9 10 9 1 10 9 2 13 10 11 14 9 12 2 11 2 1 9 10 9 2 7 13 16 2 9 1 9 16 13 9 1 9 1 9 10 9 13 0 1 10 9 1 9 0 2 2
27 7 3 2 7 2 13 9 16 13 1 9 10 9 1 9 10 9 1 9 16 10 9 4 13 1 15 2
41 7 9 15 14 10 9 13 1 10 9 2 7 1 15 10 9 16 10 9 16 13 14 10 9 2 13 9 1 10 9 7 13 1 10 9 9 13 14 15 2 2
72 9 10 9 13 16 9 10 9 4 13 14 10 9 16 13 1 9 1 9 15 3 7 9 15 2 13 9 2 1 16 16 15 13 13 7 1 16 3 4 13 15 1 9 10 9 2 2 7 3 16 10 9 13 16 2 9 0 13 13 7 13 14 13 10 9 1 13 14 10 9 2 2
24 9 12 2 11 2 13 9 0 1 9 0 14 9 9 10 9 1 10 9 1 9 10 9 2
29 1 10 15 1 15 13 1 9 10 9 10 0 9 9 16 13 14 9 15 14 9 2 16 13 1 3 0 9 2
24 3 2 7 2 13 16 9 9 16 10 9 13 1 10 9 2 1 15 1 10 9 1 9 2
41 1 1 3 2 13 16 3 1 9 9 16 13 9 1 9 15 1 9 2 7 13 9 16 10 9 13 1 9 10 9 7 1 9 15 2 2 9 11 2 2 2
21 10 9 15 13 2 3 2 9 3 0 1 9 10 9 10 0 1 9 10 9 2
27 10 9 13 1 9 9 0 13 1 9 12 2 11 2 7 13 9 1 9 16 13 1 15 1 10 9 2
18 1 9 15 14 11 11 2 7 2 13 9 2 10 9 10 13 2 2
23 12 10 9 2 16 13 1 9 10 9 10 0 2 13 1 9 10 9 9 1 10 9 2
30 9 9 10 9 13 9 10 9 16 2 9 13 2 13 1 2 9 2 2 7 7 9 15 1 10 9 4 13 0 2
15 10 9 10 0 14 9 12 2 11 2 13 1 12 9 2
18 1 9 9 2 16 7 15 13 1 10 9 2 13 2 9 9 2 2
49 9 16 13 13 14 9 15 1 9 10 9 13 1 3 16 2 13 9 2 2 7 7 13 9 15 1 10 9 0 1 10 9 3 7 13 10 9 16 9 0 13 14 15 13 1 9 10 9 2
44 9 15 13 3 1 2 9 2 2 3 1 10 16 13 1 10 9 10 0 1 9 10 9 2 7 3 13 1 10 9 10 0 9 0 13 14 10 9 16 4 13 9 9 2
25 3 13 16 13 9 0 1 9 15 2 7 0 16 9 10 9 3 13 9 1 10 9 16 13 2
19 3 2 13 1 10 9 16 13 1 9 15 14 2 9 9 2 16 9 2
9 13 15 2 15 13 14 10 9 2
16 3 9 10 9 2 16 10 9 10 0 2 0 13 10 13 2
31 9 15 14 9 12 2 11 2 13 16 10 9 13 13 1 9 13 2 1 9 10 9 10 0 1 10 9 1 9 0 2
36 7 7 7 13 9 1 9 0 1 9 1 10 9 2 7 1 1 3 13 1 10 9 2 13 3 1 10 9 10 9 13 14 15 9 0 2
24 10 9 16 1 15 13 9 10 9 3 13 2 9 1 10 9 2 1 9 15 14 10 9 2
14 7 3 2 10 9 16 9 13 1 9 9 3 13 2
36 0 16 10 9 1 10 9 13 9 0 2 7 13 1 15 1 13 1 9 10 9 16 9 0 3 1 9 10 9 4 13 1 9 1 9 2
13 9 10 9 13 1 9 1 9 15 2 9 2 2
43 15 13 16 3 15 9 14 9 16 13 1 9 10 9 2 13 9 9 16 13 9 10 9 1 9 10 9 2 7 1 15 13 13 1 10 9 16 13 2 9 9 2 2
47 13 1 15 16 7 9 13 2 13 7 1 0 2 7 3 4 13 15 2 13 9 15 1 10 9 0 3 7 13 10 9 16 9 15 13 2 1 9 2 7 2 13 13 9 9 2 2
13 9 15 0 1 9 2 9 0 2 10 0 3 2
38 1 15 13 16 7 3 13 10 9 15 14 9 15 1 10 9 2 13 9 15 4 1 9 1 9 0 1 16 4 10 9 13 14 15 1 9 15 2
29 1 10 11 3 13 9 9 1 9 10 9 10 0 2 16 13 9 11 11 7 16 9 15 9 2 9 11 2 2
16 3 16 0 13 16 10 9 3 3 13 14 10 9 10 0 2
32 7 10 9 16 3 10 9 10 0 7 3 15 16 13 2 13 1 9 15 14 9 2 3 13 14 10 9 16 10 9 0 2
25 9 13 10 0 13 14 10 9 1 9 9 10 9 1 10 9 1 10 9 1 9 0 1 9 2
31 1 3 13 3 16 13 1 9 2 1 9 7 1 9 2 10 1 10 9 10 0 1 9 10 9 10 0 14 10 9 2
37 1 9 10 9 13 16 1 1 3 13 1 9 15 2 16 13 13 1 9 15 2 10 1 9 10 9 10 0 16 13 1 9 15 14 10 9 2
21 1 9 9 10 9 2 11 11 2 13 1 9 14 12 9 7 3 1 10 9 2
27 9 15 14 9 13 10 0 13 1 9 10 9 13 1 15 9 16 13 14 15 1 12 10 9 10 0 2
24 12 10 9 1 9 16 13 3 13 1 15 9 0 1 9 15 14 15 16 13 1 10 9 2
23 3 1 12 9 3 12 1 10 10 13 1 9 11 1 10 9 10 0 13 1 9 15 2
28 1 2 9 13 16 4 13 9 13 9 2 9 2 7 13 1 9 0 7 13 14 10 9 10 0 10 0 2
38 0 1 15 2 13 1 9 0 1 9 0 1 10 9 10 0 2 16 13 2 1 10 9 2 9 9 0 1 10 9 7 1 10 9 9 9 9 2
36 16 16 15 2 4 13 3 14 10 9 16 13 1 9 15 2 1 2 1 13 14 9 15 1 10 9 10 0 2 2 10 9 13 0 2 2
62 1 3 16 13 9 1 9 1 10 9 1 9 2 15 4 13 16 13 1 9 9 1 9 9 9 0 0 3 2 10 10 9 13 9 9 12 2 9 10 9 0 1 10 9 10 0 14 10 9 2 10 9 13 9 2 9 2 7 9 9 0 2
23 10 9 0 13 16 13 1 15 9 1 9 9 16 0 1 9 9 1 9 0 2 0 2
16 3 2 7 3 2 13 10 9 16 13 1 10 9 9 0 2
20 16 16 13 1 15 9 0 2 3 2 2 7 3 15 4 3 13 9 0 2
6 15 9 0 1 11 2
28 7 2 7 15 13 9 1 9 9 1 10 9 1 9 0 15 13 9 0 16 13 1 15 9 0 7 0 2
21 7 15 13 15 1 9 9 0 1 15 9 2 13 1 15 3 9 7 3 9 2
37 10 9 10 0 13 16 10 9 1 9 1 10 9 13 9 7 4 1 9 7 1 9 9 2 7 9 10 9 14 10 9 13 1 9 10 9 2
23 1 9 10 9 10 0 13 9 0 1 10 15 2 3 1 10 9 2 3 1 10 9 2
7 9 0 15 13 3 0 2
28 10 9 10 0 16 13 2 9 9 11 2 1 9 1 9 10 9 10 10 9 10 0 2 13 13 9 15 2
27 10 9 10 3 2 0 13 13 9 1 10 9 2 13 13 13 9 0 7 15 0 3 7 4 1 9 2
10 2 10 9 13 1 10 0 3 2 2
21 9 15 13 1 15 16 9 10 9 1 10 9 0 3 7 1 10 9 10 0 2
30 1 10 9 1 9 9 10 9 0 3 1 12 9 1 9 1 10 9 2 9 9 15 13 9 9 7 9 9 2 2
12 3 2 13 10 9 16 13 9 1 10 15 2
15 3 3 13 10 9 3 1 9 0 1 9 9 7 9 2
42 10 9 1 10 9 4 13 0 7 0 3 1 10 9 1 10 9 2 7 15 4 13 1 10 9 10 9 1 10 9 2 1 9 9 1 10 9 1 15 15 13 2
38 7 10 9 13 16 9 10 9 10 0 10 0 1 9 13 10 9 1 10 9 0 3 3 1 9 10 9 10 0 7 1 15 16 13 1 10 9 2
34 1 9 10 9 4 13 14 10 9 1 10 9 16 13 1 10 9 10 0 2 7 1 9 10 9 16 13 1 10 9 1 10 9 2
17 12 13 13 9 0 1 9 16 13 2 9 12 2 1 9 9 2
30 10 9 13 0 2 12 9 1 9 10 9 1 10 9 13 9 9 0 1 9 0 2 7 9 0 13 9 0 0 2
22 1 10 10 9 13 2 3 2 9 9 0 7 0 1 10 9 1 10 9 10 0 2
19 10 9 13 9 2 7 3 9 13 9 15 1 10 9 7 1 10 9 2
26 13 14 10 9 15 3 3 0 10 9 1 9 16 13 1 15 2 7 9 0 1 9 1 9 15 2
30 1 9 0 1 10 9 10 0 2 9 10 9 1 9 13 9 0 0 7 13 3 7 10 9 1 10 9 10 0 2
20 15 16 16 9 10 9 10 0 1 10 9 13 0 3 2 7 16 3 0 2
40 1 9 1 9 14 10 9 1 9 2 9 10 9 1 9 9 10 9 13 7 2 11 2 12 9 2 11 2 11 2 12 9 2 7 11 2 11 12 9 2
33 9 9 11 2 11 1 10 9 10 0 2 2 1 10 0 3 2 2 13 7 1 9 10 0 7 10 0 1 10 9 10 0 2
64 3 16 13 1 9 15 16 9 15 1 9 2 9 15 1 9 7 1 10 9 10 0 7 9 15 1 10 9 9 15 2 13 3 13 9 3 0 1 9 0 7 13 1 12 9 9 11 11 2 13 14 9 15 16 13 1 15 13 9 15 1 9 0 2
71 1 13 1 10 9 1 9 7 15 13 16 10 9 0 3 1 10 9 10 0 15 4 13 9 12 2 3 16 13 1 9 15 14 9 15 13 9 1 9 15 7 1 9 15 13 9 16 13 1 15 9 7 13 1 15 9 3 1 9 0 2 3 1 9 0 7 3 1 9 0 2
38 9 10 9 2 11 11 2 13 13 3 1 9 10 9 14 9 3 2 9 15 14 10 9 1 9 10 9 2 1 9 9 0 14 9 9 10 9 2
32 10 9 3 13 0 10 3 13 9 10 9 7 10 9 2 11 11 2 1 9 15 13 1 10 9 16 9 10 9 3 13 2
63 1 9 15 10 13 14 10 9 1 9 10 9 2 13 9 10 9 1 9 10 9 13 2 1 1 11 2 14 10 9 14 9 10 9 1 10 10 9 2 7 9 9 1 9 10 9 1 11 2 16 13 1 9 1 10 9 1 2 9 9 10 9 2
41 9 9 10 9 2 1 15 10 9 1 9 10 9 3 13 14 9 10 9 1 10 9 2 13 1 3 2 9 15 14 10 9 13 9 14 9 9 1 10 9 2
31 7 9 9 1 10 9 2 3 10 9 4 13 1 10 9 9 13 10 9 2 16 13 1 3 1 12 12 9 1 9 2
27 3 2 9 10 9 1 10 9 1 9 10 9 13 3 14 9 15 14 10 10 9 16 13 1 9 15 2
64 3 3 13 9 2 1 9 10 9 11 2 11 7 11 2 16 9 15 14 10 9 1 9 10 9 13 9 16 13 14 10 9 1 9 9 1 10 9 13 0 2 7 16 3 3 15 13 13 10 9 16 13 1 15 1 13 1 9 15 14 9 10 9 2
6 7 0 3 9 11 2
29 15 13 1 9 0 1 9 10 9 10 0 3 2 7 9 15 1 9 1 10 9 1 10 9 13 0 1 3 2
7 15 13 1 15 9 2 2
21 9 15 13 10 9 11 11 1 9 1 9 1 9 9 10 9 1 11 7 11 2
52 3 2 3 4 13 13 1 9 0 3 2 7 9 10 9 2 16 1 15 9 12 10 9 13 12 1 9 9 1 9 1 9 0 2 13 13 14 1 15 2 16 11 7 11 3 2 13 1 15 9 2 2
59 10 9 2 16 1 2 9 15 13 9 15 2 13 1 10 9 16 1 15 10 9 1 9 10 9 1 9 10 9 13 14 9 15 3 1 10 9 10 9 2 0 2 9 14 9 15 13 4 13 14 9 10 9 16 13 1 10 9 2
46 9 10 9 1 11 7 9 9 0 14 10 9 10 0 1 11 13 9 0 1 11 7 11 2 7 1 10 0 16 13 9 0 1 10 9 10 0 2 16 9 15 2 9 0 2 2
54 11 13 2 1 2 9 9 10 9 2 1 9 0 2 7 9 15 14 10 9 10 0 1 11 13 9 16 4 1 15 13 1 15 2 11 11 4 13 13 14 15 2 7 10 9 10 0 13 1 10 9 10 0 2
45 7 3 13 1 9 15 16 3 13 14 15 3 1 9 15 2 1 9 13 2 1 9 9 1 10 15 2 13 14 10 9 16 13 3 14 11 2 11 7 11 1 9 10 9 2
18 16 16 11 13 1 13 2 15 13 13 1 10 9 13 1 9 15 2
18 11 4 13 0 1 9 9 9 15 1 2 9 9 10 9 10 0 2
18 9 10 9 1 11 13 2 16 9 0 1 11 3 13 1 9 0 2
45 15 9 13 2 16 15 13 1 15 1 9 2 13 0 3 2 7 10 9 10 0 13 13 14 11 1 10 16 13 1 9 15 14 10 9 10 0 2 1 11 7 1 11 15 2
57 7 10 9 2 9 0 2 13 9 9 3 14 11 13 4 3 13 1 9 0 1 10 9 10 0 2 3 4 11 13 2 16 10 9 13 1 15 2 1 9 9 7 1 9 9 2 14 9 10 9 1 9 10 9 10 0 2
10 0 13 2 16 9 15 3 3 13 2
23 10 9 1 11 13 1 10 9 14 10 9 13 14 10 9 2 16 13 1 15 1 3 2
22 10 9 10 0 13 3 13 14 9 9 10 9 1 9 10 9 16 15 13 1 11 2
28 10 9 0 13 9 15 7 7 13 1 15 2 3 13 14 11 1 10 9 14 11 2 16 15 3 13 9 2
18 11 13 13 1 9 15 2 7 15 13 9 15 15 1 10 10 9 2
27 1 15 2 15 13 3 13 1 9 10 9 7 15 13 1 9 1 11 3 1 9 1 10 9 14 15 2
61 7 15 4 1 9 0 2 7 7 10 9 10 0 10 0 1 9 11 4 13 14 11 2 3 15 0 13 1 15 14 10 9 16 13 1 9 10 9 10 0 7 13 1 9 15 14 9 10 9 1 9 16 13 1 15 7 3 7 1 11 2
35 10 9 10 0 14 9 10 9 13 1 9 0 1 9 1 9 1 9 10 9 1 9 10 9 2 1 10 9 1 9 10 9 1 9 2
12 10 9 13 9 2 9 7 9 1 10 9 2
23 10 9 13 1 9 0 14 9 9 10 9 2 16 13 1 9 10 9 1 9 2 9 2
22 12 1 9 10 9 13 13 1 9 1 9 1 10 9 2 7 13 3 13 14 15 2
29 1 9 2 9 10 9 2 11 11 2 13 13 9 9 13 1 10 9 1 9 9 10 9 1 10 9 10 0 2
15 10 9 7 13 1 9 9 9 1 9 9 1 10 9 2
54 8 8 8 16 13 9 10 9 1 9 9 15 14 9 0 1 9 10 9 1 10 9 1 9 10 9 2 13 3 1 9 1 9 9 10 9 7 10 9 2 9 10 9 2 9 9 10 9 7 10 9 10 0 2
42 1 2 9 10 9 16 13 9 10 9 2 11 11 2 13 1 9 1 9 1 12 9 1 12 9 1 10 9 10 0 14 9 10 9 16 13 9 1 9 1 9 2
7 10 9 13 1 12 9 2
31 1 9 10 9 13 10 9 9 1 9 7 1 9 1 10 9 10 0 2 16 13 1 9 9 0 7 1 9 9 0 2
26 10 9 13 1 9 15 9 9 1 9 14 3 12 9 1 9 15 10 0 1 12 10 9 10 0 2
40 1 9 10 9 2 10 9 16 13 9 10 9 1 9 10 9 4 2 1 9 15 2 13 1 15 12 9 1 9 10 9 2 9 10 9 7 9 10 9 2
16 1 15 2 13 16 10 9 13 1 10 9 13 0 3 12 2
37 9 7 9 9 2 11 2 13 1 1 12 9 2 13 15 16 13 2 13 14 10 9 2 7 16 3 13 1 10 9 16 13 1 15 9 9 2
35 1 9 2 12 7 1 11 2 10 9 14 10 9 2 16 1 3 13 1 9 1 10 9 7 1 9 9 1 10 9 15 13 12 3 2
31 3 15 13 2 7 15 2 16 1 9 15 14 11 13 12 12 9 2 13 13 12 12 7 13 16 13 1 12 12 2 2
18 3 9 10 9 10 0 2 1 9 2 11 2 7 1 9 10 9 2
21 13 9 16 10 9 2 9 13 1 9 10 9 1 16 13 2 3 1 9 0 2
16 4 16 7 10 9 15 13 13 1 10 9 10 0 10 0 2
14 3 3 13 10 9 1 16 13 9 15 1 10 11 2
18 7 13 16 3 4 13 14 9 15 16 1 10 9 1 9 9 15 2
18 3 13 15 10 9 10 0 1 9 15 1 11 1 10 9 10 0 2
25 12 10 9 16 13 1 1 12 9 3 13 9 14 9 7 3 3 10 9 16 13 1 9 9 2
45 1 16 9 9 10 9 10 0 13 16 3 13 14 9 15 10 0 1 9 9 7 9 2 13 15 9 2 16 9 10 9 10 0 16 1 15 3 13 1 15 16 1 9 11 2
26 13 16 9 0 14 10 9 13 15 9 3 2 10 13 3 1 9 10 13 10 0 1 10 9 9 2
40 9 10 9 16 13 1 9 2 10 9 10 15 2 13 0 1 10 9 16 13 1 10 9 2 1 1 9 0 3 14 10 9 2 16 13 13 1 9 15 2
23 4 13 16 3 9 1 9 9 10 9 2 10 9 13 9 11 2 7 9 15 10 0 2
22 9 15 13 9 11 2 7 10 9 13 1 9 2 1 9 2 1 9 7 1 11 2
13 1 9 2 2 10 9 10 0 2 1 10 9 2
28 3 10 9 10 15 13 1 13 1 9 10 9 16 1 11 0 7 0 7 16 1 9 15 16 13 1 9 2
18 15 3 9 3 2 7 3 3 9 4 13 2 7 3 13 1 15 2
38 0 1 15 2 1 11 7 1 2 11 2 13 9 0 1 9 0 14 10 9 2 1 9 9 15 15 13 9 1 9 1 9 2 9 2 7 9 2
26 3 1 15 2 4 13 14 11 1 9 15 10 0 2 7 3 13 1 10 9 7 9 15 13 15 2
24 1 9 15 14 9 15 13 3 3 7 9 0 9 0 7 3 0 2 7 1 10 15 9 2
29 3 1 10 9 10 0 7 10 0 16 1 10 9 13 9 0 13 14 9 15 14 15 16 13 13 14 9 15 2
19 1 3 9 15 10 0 14 11 1 9 9 1 10 9 10 0 14 15 2
46 13 9 7 9 3 1 10 15 16 13 1 2 9 9 15 10 0 16 10 10 9 1 15 2 16 13 1 9 1 10 9 1 9 2 11 2 2 13 1 10 10 13 1 10 9 2
19 3 11 13 14 10 9 16 1 10 9 7 9 7 7 13 1 15 3 2
33 10 9 10 0 13 9 14 10 9 10 0 10 0 3 2 16 13 14 10 9 1 9 10 9 7 13 1 9 9 9 0 0 2
27 12 9 9 15 14 10 9 13 1 9 0 14 10 9 9 2 16 10 9 1 10 9 13 3 2 0 2
29 1 9 1 10 9 13 10 9 13 7 16 9 9 1 10 9 13 9 1 10 9 10 0 7 1 9 10 9 2
49 13 15 3 13 16 1 9 9 15 14 10 9 13 9 0 2 16 13 9 2 9 14 9 15 1 10 9 2 9 15 14 10 9 10 0 9 15 9 9 2 0 1 10 9 2 1 10 9 2
35 1 9 9 15 1 10 9 2 14 10 9 10 15 3 2 4 13 1 10 9 0 2 16 9 13 9 2 9 2 9 15 14 9 11 2
34 7 7 9 10 9 13 9 13 2 10 9 10 0 1 10 9 10 0 10 15 13 9 10 9 7 9 15 1 9 9 7 1 9 2
10 15 10 9 14 9 10 9 10 0 2
41 10 3 10 9 1 10 9 7 10 9 1 1 10 9 3 13 1 9 0 1 9 10 9 10 0 2 10 10 13 1 10 9 10 0 1 10 9 13 7 13 2
11 10 15 13 10 9 7 3 2 11 2 2
13 11 3 13 7 13 14 10 9 10 0 10 15 2
7 11 2 11 7 11 2 2
22 9 14 9 9 13 7 13 1 11 1 9 9 10 9 16 13 1 9 1 9 9 2
42 12 9 0 13 1 11 1 9 11 2 3 13 10 9 1 11 2 1 9 10 9 10 0 7 9 10 9 1 9 9 3 0 7 1 9 0 1 10 9 16 13 2
39 9 9 13 3 1 11 2 9 0 1 9 11 2 7 1 10 9 10 0 13 9 1 9 0 2 1 9 12 9 1 9 10 9 1 10 9 10 0 2
18 9 10 9 13 1 10 9 16 13 1 11 1 9 10 9 10 0 2
32 12 9 9 0 13 14 9 9 10 9 10 0 1 9 1 9 16 13 13 1 10 9 1 9 9 10 9 10 0 10 0 2
47 9 13 16 7 16 3 13 1 10 9 12 9 14 9 1 9 10 9 2 3 15 4 13 1 9 9 0 2 16 13 1 9 1 9 9 10 9 14 10 9 7 10 9 1 9 0 2
36 9 10 9 2 9 9 2 16 13 3 9 14 9 9 0 16 3 13 1 15 12 9 2 13 14 9 10 9 7 13 16 13 1 15 9 2
27 1 9 11 16 13 13 10 12 9 1 9 9 15 14 9 11 3 11 2 16 13 1 10 9 1 12 2
24 15 13 1 9 15 1 9 10 9 1 11 2 3 13 10 9 3 0 1 10 9 10 0 2
50 10 9 1 10 9 1 11 13 9 1 9 10 9 1 10 9 1 9 10 9 2 7 13 9 0 1 2 9 12 9 7 1 15 9 1 9 9 1 10 9 7 11 4 13 9 7 13 1 9 2
14 1 9 10 9 13 3 10 9 10 0 14 10 9 2
22 10 9 13 1 9 10 9 1 10 9 7 1 9 10 9 16 13 1 9 10 9 2
28 1 9 10 9 7 10 9 0 2 10 9 13 3 1 10 11 9 0 1 10 9 10 0 1 9 10 9 2
34 1 9 0 15 13 3 1 3 13 11 11 1 9 11 11 13 14 11 7 11 11 13 14 9 10 9 10 3 2 0 1 10 9 2
7 3 11 11 13 1 11 2
7 3 13 1 9 15 13 2
8 10 9 1 12 13 9 0 2
26 11 11 7 11 11 7 11 11 7 11 11 1 9 10 9 10 0 1 9 9 1 10 9 1 11 2
36 15 13 1 9 10 9 1 12 10 9 7 15 1 10 9 14 10 9 2 7 9 2 10 9 1 10 9 1 10 9 10 0 1 9 0 2
61 3 13 1 10 9 9 11 11 2 16 7 9 15 13 14 9 10 9 7 10 9 2 3 9 0 14 10 9 10 0 2 7 1 9 2 3 9 0 14 11 1 10 9 2 7 9 3 2 7 3 9 1 10 9 2 7 1 9 0 3 2
5 11 11 13 13 2
8 15 1 9 1 9 7 9 2
26 7 13 15 9 13 1 9 10 9 1 9 7 9 3 1 11 2 3 1 9 9 10 9 10 0 2
46 3 13 1 9 15 1 2 9 10 10 9 7 9 1 10 9 16 13 1 10 9 2 16 13 1 11 13 14 10 9 1 9 10 11 2 1 16 13 14 9 15 1 15 1 15 2
8 3 13 9 15 1 10 9 2
6 3 1 10 9 13 2
15 11 11 13 13 1 15 3 9 13 1 2 11 11 2 2
39 15 13 1 15 9 2 9 2 16 1 9 11 3 4 10 11 13 14 9 15 10 0 2 7 3 13 1 10 9 9 0 16 13 1 9 14 10 9 2
35 9 9 10 9 1 9 10 9 2 13 11 1 9 2 3 1 9 11 11 2 3 13 14 11 1 10 9 1 9 7 9 16 13 3 2
8 7 3 15 13 13 3 3 2
13 3 13 1 10 11 14 11 1 10 9 10 9 2
12 3 13 7 13 14 9 15 1 9 10 9 2
25 1 1 15 16 7 1 10 9 1 10 9 1 9 2 11 3 13 3 9 9 10 9 13 9 2
11 9 15 14 9 11 13 14 9 10 9 2
22 3 9 15 7 11 1 9 9 10 9 13 13 2 16 10 9 1 10 9 13 9 2
28 3 9 11 2 16 9 10 9 10 0 1 9 10 9 3 13 14 11 1 9 1 10 13 3 2 13 0 2
11 3 16 13 13 13 13 1 9 7 9 2
14 11 7 11 13 3 1 16 9 11 7 11 13 0 2
11 15 13 1 10 9 10 0 14 10 9 2
51 1 16 15 13 13 1 10 9 13 14 9 15 1 15 2 13 9 0 7 13 1 10 9 7 1 10 9 7 1 9 2 9 3 0 7 13 9 0 1 9 9 7 9 0 1 11 1 9 10 9 2
21 1 9 1 9 15 3 4 3 13 9 1 9 2 10 9 14 10 9 10 0 2
35 15 13 1 9 9 0 7 0 1 14 15 2 16 13 3 7 13 1 15 9 2 16 13 1 9 10 9 10 0 14 11 1 9 0 2
17 9 11 7 0 3 1 9 15 10 0 13 9 9 1 10 9 2
15 3 13 3 9 1 10 9 3 1 11 2 11 7 11 2
11 1 10 9 3 1 11 2 11 7 11 2
66 13 9 1 9 11 1 9 10 11 2 10 9 7 9 8 8 1 9 9 9 0 2 1 9 3 2 0 1 10 9 16 13 9 15 1 10 9 2 7 1 9 0 14 10 9 2 16 3 13 3 9 9 7 3 2 7 1 3 15 0 1 10 9 10 0 2
45 7 9 8 8 10 0 1 9 1 11 2 16 15 13 7 0 10 3 3 13 1 15 13 9 9 1 9 9 15 8 8 8 2 13 1 9 3 9 7 9 1 10 9 9 2
7 15 3 0 1 9 11 2
15 3 16 3 13 1 9 11 1 11 3 13 7 3 13 2
18 9 10 9 13 1 9 10 9 7 13 16 3 13 1 15 9 0 2
8 11 3 13 1 15 1 11 2
30 1 9 7 9 13 1 9 2 10 9 10 0 14 10 9 7 1 2 12 9 1 11 14 10 9 4 13 9 0 2
62 1 9 1 9 8 8 10 0 1 11 7 9 10 9 2 13 9 15 14 10 11 11 11 1 11 13 3 1 10 9 2 16 13 1 9 15 9 0 1 11 2 1 15 16 10 9 13 13 14 11 1 9 15 10 0 7 10 0 1 10 9 2
26 9 13 13 2 16 1 3 13 10 9 1 10 9 2 13 10 9 10 0 1 13 1 11 9 0 2
31 16 13 14 11 1 9 2 10 9 10 0 2 16 15 13 2 13 1 10 9 16 3 3 10 9 13 1 15 9 0 2
42 1 9 0 2 13 9 16 1 15 11 13 1 13 9 1 10 9 10 0 3 1 10 9 10 0 1 10 9 10 0 1 15 13 1 15 9 0 1 9 9 0 2
41 1 15 2 1 9 0 2 7 1 15 1 10 15 16 1 1 10 9 13 1 9 2 13 10 9 3 9 0 1 10 9 10 0 7 9 9 0 0 1 9 2
42 1 11 13 16 13 3 2 16 3 9 10 9 13 14 9 15 14 11 1 9 0 7 9 15 2 16 1 11 13 10 9 9 0 7 7 3 1 10 9 10 0 2
31 1 9 15 14 3 9 0 0 7 9 0 2 1 9 14 9 0 0 2 13 9 10 9 8 8 8 1 12 10 9 2
56 9 11 11 2 1 10 9 1 9 0 1 9 11 2 13 16 11 4 13 15 13 1 3 16 13 1 9 15 14 9 10 9 1 10 9 2 1 13 1 10 9 14 11 2 7 1 3 16 13 1 9 9 9 0 0 2
42 9 15 14 10 9 16 13 1 10 9 10 0 13 1 9 1 15 16 11 13 13 1 9 0 3 2 16 16 3 13 9 10 9 2 1 10 9 0 1 9 15 2
19 7 9 15 14 9 0 12 3 1 9 11 13 9 0 0 1 9 0 2
22 9 15 14 11 2 3 7 3 13 1 15 2 4 13 1 9 9 0 1 10 9 2
49 1 9 1 10 15 2 1 9 15 14 9 0 1 11 1 11 2 4 10 9 10 0 13 9 2 16 13 1 9 9 15 1 0 7 13 1 10 9 16 3 15 13 14 9 15 14 10 9 2
53 9 0 1 9 10 9 13 1 9 10 9 2 16 13 10 9 13 1 8 8 1 9 3 2 1 10 9 10 0 10 0 2 1 10 16 13 8 8 8 10 0 14 12 10 9 2 10 13 1 9 14 9 2
13 1 9 10 9 10 0 2 13 2 13 10 9 2
28 10 9 13 8 8 8 8 1 10 15 0 9 14 9 3 0 1 10 9 2 16 3 13 9 13 9 3 2
33 9 0 0 13 3 9 0 1 10 9 2 16 13 1 9 0 0 2 16 1 15 13 12 9 9 0 2 0 2 0 7 0 2
50 9 9 3 14 9 1 10 15 1 10 9 10 0 10 0 1 10 9 4 13 1 9 2 16 1 9 15 13 9 9 10 9 11 2 7 10 9 10 0 16 13 1 11 1 15 2 1 9 9 2
36 9 15 14 9 9 10 9 10 0 1 11 12 9 1 16 13 2 13 13 9 1 10 9 10 0 16 13 1 9 9 10 9 1 10 9 2
17 7 2 3 10 13 3 1 9 3 14 10 9 10 0 10 0 2
26 13 9 0 1 9 9 1 12 10 9 1 9 9 15 10 0 14 11 1 14 9 0 1 10 9 2
40 1 12 10 9 2 1 11 7 1 11 2 13 10 9 2 16 3 7 13 11 1 13 3 14 9 11 2 3 13 9 0 1 16 11 13 13 15 1 15 2
50 10 9 10 0 10 13 7 10 9 1 9 9 15 10 0 14 11 11 13 1 9 10 9 10 0 3 16 13 4 1 15 13 1 9 0 1 9 9 10 9 1 15 7 1 9 10 9 10 0 2
14 3 13 3 1 9 9 0 9 9 10 9 1 11 2
7 1 11 9 0 13 15 2
38 9 15 14 9 10 9 1 11 13 1 9 10 9 1 11 14 10 9 16 13 1 9 10 9 1 12 10 9 2 16 4 13 1 9 1 15 9 2
23 3 1 9 15 14 11 4 9 2 16 9 15 9 7 9 1 9 10 9 10 3 0 2
30 4 13 16 9 1 9 1 15 13 3 2 1 9 9 15 1 11 14 9 9 10 9 2 1 9 10 9 11 11 2
40 10 9 13 3 1 11 14 1 9 10 9 3 9 9 7 9 2 7 13 9 16 9 15 13 13 14 10 9 10 0 3 1 10 10 0 1 9 10 9 2
24 10 9 1 10 9 13 1 9 15 3 9 15 14 9 9 1 9 9 1 10 9 10 0 2
27 10 9 13 1 9 1 12 9 10 9 10 0 1 9 9 2 16 13 1 9 9 10 9 14 10 9 2
23 1 10 9 10 0 13 9 14 9 9 1 11 2 16 13 9 16 13 1 12 12 9 2
30 10 9 10 12 13 8 8 8 10 0 2 14 9 10 9 2 11 11 2 13 9 14 12 12 11 0 1 10 9 2
40 11 2 16 9 10 9 14 15 13 1 9 9 1 9 0 2 2 9 2 2 2 13 1 9 10 9 2 1 9 16 9 10 9 14 15 13 1 9 0 2
39 12 9 15 3 13 13 7 13 9 9 9 13 2 9 9 2 2 7 3 13 14 9 10 9 2 1 9 13 14 9 9 15 14 9 0 1 10 9 2
23 1 9 8 8 14 9 9 9 3 13 16 10 9 13 13 1 9 9 9 1 9 0 2
28 1 9 9 9 13 16 10 9 16 4 13 1 9 9 15 14 9 9 1 9 9 1 9 13 1 10 9 2
26 10 9 16 3 13 13 1 9 10 9 1 10 9 10 12 14 12 2 16 13 1 10 9 10 0 2
28 13 16 1 9 9 13 9 3 1 12 8 8 10 0 14 12 2 7 3 1 10 9 10 12 14 10 9 2
24 10 9 1 8 8 2 11 11 2 13 8 8 8 10 0 9 1 12 10 9 1 9 9 2
16 1 10 9 1 8 8 3 13 14 15 1 9 9 9 0 2
20 3 3 13 3 3 1 9 0 1 10 16 13 1 9 9 9 1 9 9 2
25 9 0 13 14 9 9 9 9 1 9 12 10 9 2 1 13 14 9 10 9 7 9 1 15 2
21 3 13 9 9 1 9 1 9 9 9 9 1 9 9 1 9 0 1 9 15 2
9 13 3 14 10 9 13 1 9 2
25 1 9 10 9 10 0 13 11 1 9 14 2 11 2 1 10 11 7 13 14 15 2 3 13 2
12 15 13 16 15 13 13 3 9 1 10 9 2
15 13 1 15 14 10 9 2 10 9 3 13 2 13 11 2
15 13 1 15 14 10 9 2 10 9 3 13 2 13 11 2
14 1 10 9 13 3 1 10 9 16 11 13 1 15 2
18 14 15 13 9 2 13 9 11 1 9 10 9 7 3 10 9 13 2
32 1 11 3 13 16 13 1 2 8 8 13 14 10 9 1 9 0 14 9 10 9 1 9 16 13 1 15 9 1 10 9 2
32 10 9 1 9 1 10 15 13 0 2 16 13 1 9 10 9 7 1 3 16 13 1 9 10 9 14 9 0 1 10 9 2
48 1 10 9 10 15 13 11 1 9 11 10 0 2 1 9 0 2 1 9 15 14 9 11 1 9 2 9 2 14 13 1 3 10 9 1 9 9 10 9 1 9 10 9 1 9 10 9 2
41 1 9 11 13 14 9 15 2 13 1 9 15 11 9 16 13 1 15 9 1 10 9 2 1 15 11 13 1 9 7 13 1 10 9 10 0 13 14 10 9 2
28 2 7 13 3 13 14 10 9 2 2 13 11 1 2 10 9 2 2 2 4 13 9 0 7 3 0 2 2
28 11 2 10 9 16 1 10 9 1 11 7 9 11 2 13 1 10 9 10 0 1 9 16 13 1 10 9 2
26 15 13 1 15 1 9 15 1 10 11 7 1 9 2 11 2 1 11 2 3 13 10 9 10 0 2
27 1 9 9 15 10 0 13 9 0 2 13 9 15 2 16 11 13 13 3 7 13 1 9 1 9 15 2
44 12 1 15 2 7 2 13 3 13 1 9 0 13 9 1 9 11 2 1 16 13 16 15 13 9 9 1 10 9 7 13 1 15 13 3 1 10 9 1 9 9 10 9 2
19 11 13 1 9 15 2 16 13 9 0 3 1 9 15 13 1 10 9 2
37 1 9 1 10 15 2 15 13 2 9 2 7 15 3 13 2 11 2 2 2 13 1 10 9 12 10 9 2 9 10 0 16 9 1 10 9 2
27 8 8 1 15 3 9 0 2 13 9 9 1 9 10 9 2 16 13 13 9 1 4 3 14 10 9 2
14 14 13 1 15 2 13 1 15 2 3 3 1 15 2
21 13 9 16 13 14 9 15 7 3 3 1 15 13 9 7 3 1 15 13 9 2
29 11 13 13 1 10 9 16 13 3 1 9 11 10 0 2 7 13 2 1 9 15 13 1 10 9 1 11 1 2
29 15 1 10 9 16 13 9 1 9 9 15 10 12 2 7 10 9 16 11 3 13 14 11 1 10 9 10 0 2
30 2 13 4 13 1 15 2 2 13 11 2 2 7 3 1 15 13 1 12 2 14 15 4 13 1 10 9 14 15 2
21 9 15 10 0 7 10 0 1 11 13 13 1 9 10 9 16 15 13 1 15 2
14 15 13 1 11 3 3 0 7 10 9 14 15 0 2
19 3 10 9 13 16 13 1 15 9 2 7 3 15 16 13 13 15 2 2
6 11 2 11 11 2 2
31 10 9 1 11 13 1 9 11 1 9 0 1 11 2 16 13 1 10 9 9 0 9 2 0 7 13 14 9 10 9 2
52 2 9 15 13 1 10 9 10 0 3 14 10 9 10 0 7 14 9 10 9 2 2 13 10 9 1 9 16 13 12 9 3 1 10 9 10 0 7 16 13 1 10 10 9 10 9 16 13 12 12 9 2
11 10 9 10 0 13 1 10 9 10 0 2
30 10 9 2 16 1 9 0 13 14 10 9 2 7 13 2 1 10 9 10 0 2 13 14 9 14 9 1 10 9 2
32 2 1 9 10 9 13 10 9 14 9 9 0 2 10 9 13 7 10 9 13 14 10 9 2 2 13 1 10 9 10 0 2
41 8 8 8 11 13 13 14 10 9 10 0 1 9 0 1 10 9 1 9 11 2 16 13 1 9 9 10 9 1 15 13 10 9 7 1 9 15 13 9 0 2
22 9 9 1 10 9 10 0 13 14 10 9 2 13 1 10 9 7 13 1 15 2 2
14 1 9 10 9 10 0 13 10 9 1 1 10 9 2
34 10 9 11 2 16 9 13 1 10 9 14 15 1 11 2 3 13 1 10 9 1 15 13 10 9 14 10 9 1 10 9 10 0 2
15 3 9 10 9 11 2 9 12 2 3 13 1 10 9 2
43 10 9 10 0 14 9 9 9 9 13 1 10 9 14 9 10 9 1 12 1 9 9 0 2 10 13 16 13 14 9 10 9 10 0 14 10 9 1 1 9 7 9 2
61 10 9 13 9 13 1 10 9 14 11 9 2 11 2 9 9 10 9 2 16 13 1 9 10 9 1 10 9 2 7 3 14 12 10 13 11 11 7 9 11 2 1 9 16 13 1 9 2 11 1 15 16 13 1 15 3 13 14 10 9 2
36 1 9 11 1 9 7 9 13 9 9 0 12 9 9 2 1 15 9 2 11 2 16 16 13 9 9 1 9 9 9 1 10 9 10 0 2
15 1 15 13 9 10 9 13 9 2 7 10 9 13 13 2
19 13 10 9 7 10 9 3 13 9 1 10 9 7 13 13 14 10 9 2
9 3 13 2 9 2 1 10 9 2
42 9 10 9 14 10 9 2 16 13 14 10 9 2 13 16 10 9 13 7 9 0 2 16 13 14 9 10 9 1 9 10 9 1 9 10 9 1 10 9 10 0 2
8 9 10 9 13 1 10 9 2
14 12 10 9 13 1 10 9 1 9 10 9 10 0 2
31 3 4 13 3 1 11 9 9 10 9 9 11 2 9 11 2 1 13 1 9 0 1 9 10 9 10 0 9 10 9 2
15 10 9 10 0 13 16 9 10 9 4 1 15 12 9 2
26 1 9 11 2 1 16 10 9 15 13 14 10 9 13 1 10 9 2 15 13 1 9 11 1 11 2
41 10 9 13 14 9 10 9 1 11 1 9 10 9 2 1 13 9 15 14 9 0 9 9 9 10 9 2 11 11 11 2 13 1 9 15 9 13 14 10 9 2
20 9 9 9 0 13 13 1 1 10 9 1 9 14 9 9 1 9 10 11 2
36 7 1 10 9 1 9 12 3 13 10 9 14 9 11 1 9 15 2 13 14 10 9 1 11 7 3 15 13 13 3 14 9 9 1 11 2
27 10 9 13 1 15 16 13 1 15 3 9 9 11 7 3 13 9 1 9 15 1 9 10 9 10 12 2
20 9 10 9 13 13 1 9 9 2 9 11 11 2 1 13 1 9 10 9 2
17 1 10 9 1 9 9 1 9 2 9 13 10 9 13 9 9 2
19 1 10 9 1 10 9 13 9 3 13 9 1 10 9 1 1 9 0 2
64 1 9 9 10 9 7 10 9 1 9 9 2 9 11 11 7 1 9 10 9 16 3 13 9 1 9 10 9 1 9 9 2 10 3 3 13 1 10 11 9 1 9 9 2 13 10 9 16 3 3 13 13 1 9 10 9 1 1 9 14 10 10 9 2
13 13 16 9 10 9 13 0 1 9 15 14 9 2
31 10 9 13 1 9 2 1 10 9 2 14 10 10 9 16 13 1 10 9 3 2 1 9 10 9 2 1 9 9 0 2
20 10 9 3 4 3 1 9 10 9 2 11 11 2 13 1 9 9 10 9 2
68 9 10 9 7 10 9 14 10 11 1 9 9 11 11 13 9 1 9 9 2 16 4 13 1 10 9 13 1 9 10 9 2 7 9 1 9 10 9 1 9 1 9 10 9 3 13 9 1 10 9 11 2 13 1 9 15 9 10 9 1 9 12 7 12 1 10 9 2
16 9 13 1 9 0 7 9 16 13 1 9 14 12 12 9 2
36 9 10 9 13 1 9 10 9 13 3 2 9 1 9 9 2 1 13 9 9 7 13 14 10 9 1 16 13 1 9 10 9 10 0 3 2
28 9 9 10 9 9 11 11 2 11 2 11 2 13 9 0 1 9 10 9 1 9 3 9 9 1 9 9 2
30 9 11 13 16 9 10 9 14 10 9 13 1 10 9 2 13 9 14 9 9 10 9 1 10 9 7 1 9 15 2
46 1 9 10 9 16 13 1 9 15 13 9 10 9 9 9 16 13 1 9 1 13 1 9 10 9 7 10 9 13 9 16 13 1 9 9 10 9 16 13 14 9 9 1 9 0 2
28 9 9 10 9 7 10 9 2 9 11 11 13 1 9 2 2 9 9 9 13 9 1 9 1 9 10 9 2
32 7 1 16 10 9 3 13 1 9 15 16 1 10 9 13 14 10 9 10 0 1 9 9 2 3 4 13 14 10 9 2 2
36 9 11 13 8 8 8 8 10 0 13 1 9 10 9 13 13 9 1 10 9 1 9 9 0 1 9 12 12 1 9 9 2 9 11 2 2
28 15 1 16 13 16 1 12 9 14 9 3 13 10 9 1 9 15 13 1 9 1 9 10 9 1 10 9 2
30 9 10 9 13 13 10 9 10 0 10 0 1 9 9 9 11 7 13 1 10 9 1 9 1 9 9 1 10 9 2
98 7 1 16 13 16 10 9 13 13 1 9 9 12 9 1 9 10 9 1 9 9 14 12 9 1 12 9 1 9 15 2 7 3 13 13 1 9 9 9 7 10 9 14 10 9 1 10 9 10 9 1 10 9 2 1 10 9 1 9 9 9 9 10 13 10 0 1 15 10 0 1 9 13 10 0 2 2 13 13 14 10 9 7 13 1 9 1 13 9 0 1 9 10 9 1 10 9 2
61 1 9 1 9 16 13 1 9 10 9 9 10 9 10 0 1 10 9 10 0 2 9 11 11 2 13 16 10 9 10 0 14 9 13 0 1 9 10 9 1 9 11 12 13 12 9 2 9 15 14 9 9 12 9 2 14 9 0 12 9 2
5 9 15 13 9 2
12 7 9 15 13 13 14 10 9 1 9 9 2
22 10 9 13 16 9 15 14 9 9 15 13 1 12 1 9 0 1 12 1 9 0 2
36 1 13 1 15 13 10 9 13 14 10 9 1 9 9 9 2 9 16 4 13 14 9 15 1 9 0 16 13 1 12 1 12 9 1 9 2
37 9 10 9 2 1 9 9 11 2 13 13 14 9 15 14 9 2 9 7 9 2 10 13 1 12 9 1 9 10 9 1 12 9 1 12 9 2
58 9 15 14 9 1 9 9 11 13 12 9 1 9 7 10 9 13 13 1 12 9 2 13 9 2 2 9 0 14 10 9 13 13 14 9 10 9 1 12 9 1 12 9 1 9 2 7 14 10 9 1 12 1 12 9 1 9 2
30 1 15 13 10 9 13 1 12 9 14 9 15 14 9 13 16 9 15 10 0 3 13 12 9 7 13 1 12 9 2
4 9 13 9 2
53 9 11 13 16 2 10 9 10 0 13 13 1 9 9 0 1 9 15 1 12 9 1 10 9 13 3 1 10 9 10 0 7 7 3 1 12 9 13 1 9 15 16 16 10 9 13 15 2 13 1 9 2 2
15 3 0 9 0 16 13 4 13 1 9 1 10 15 0 2
23 10 9 1 9 15 13 13 1 9 1 9 7 13 14 11 1 9 1 2 10 0 2 2
24 10 9 1 9 10 9 11 11 13 1 9 1 9 2 16 13 1 9 9 7 1 9 0 2
11 1 15 13 10 9 2 11 11 11 2 2
62 1 10 9 2 16 13 1 9 16 13 9 16 13 14 10 9 2 13 16 9 9 15 13 16 11 2 11 11 13 1 9 0 7 1 9 0 13 9 1 9 2 11 2 2 16 10 9 1 15 13 3 1 11 1 9 1 13 16 13 1 9 2
16 9 0 13 14 10 9 2 9 10 9 14 9 10 12 2 2
24 3 13 9 16 12 1 10 9 1 10 9 13 1 9 9 7 13 9 0 7 9 1 9 2
11 10 9 13 16 1 9 10 9 13 3 2
55 1 9 16 13 3 1 9 2 9 0 1 11 2 13 12 9 1 9 10 9 1 9 14 9 11 2 16 12 9 1 10 13 16 13 9 2 9 9 15 15 1 9 9 0 1 9 9 7 9 7 1 9 11 0 2
17 7 9 15 2 13 9 13 1 9 15 7 13 14 9 10 9 2
32 9 0 1 10 9 10 0 1 9 13 1 10 9 16 1 10 9 13 9 16 10 9 3 13 1 9 9 7 1 9 0 2
44 8 8 8 2 11 11 11 2 13 3 16 1 11 12 13 1 11 9 9 2 7 1 9 1 9 0 16 13 1 9 0 1 9 15 2 13 1 9 1 9 9 10 0 2
15 1 10 9 16 13 13 11 9 14 12 9 1 9 15 2
16 15 13 9 14 9 9 1 10 9 16 0 1 9 11 11 2
15 9 10 9 11 11 13 14 11 1 9 0 2 0 3 2
23 2 15 3 13 1 9 2 13 13 9 1 9 7 1 10 9 13 13 1 9 10 9 2
10 3 13 1 10 9 1 9 0 2 2
20 11 13 16 11 13 1 9 9 7 13 3 1 10 9 1 10 9 10 9 2
14 16 13 9 15 14 11 1 10 9 2 13 11 13 2
20 1 9 15 14 11 13 9 14 9 9 7 9 16 13 1 9 9 2 0 2
34 9 10 9 13 9 16 11 2 16 13 9 9 1 9 11 16 1 11 2 13 13 9 1 11 11 7 13 16 13 13 14 9 15 2
25 9 1 9 11 11 13 16 13 13 14 10 9 10 0 14 10 9 16 1 15 13 11 1 11 2
11 15 13 14 10 9 10 0 1 10 9 2
25 10 9 16 13 3 1 9 9 10 11 1 11 2 13 1 10 9 7 1 9 9 1 10 9 2
22 12 1 10 9 13 3 1 10 9 10 0 1 9 0 9 12 9 16 13 1 9 2
19 9 15 13 1 9 9 2 16 13 9 9 10 9 1 1 10 9 3 2
23 1 15 2 13 10 9 10 0 3 3 1 9 10 9 10 0 10 0 16 13 1 11 2
31 10 9 13 3 9 10 9 2 7 10 9 13 1 10 9 7 13 1 10 9 10 0 16 13 1 10 9 1 11 3 2
19 1 9 10 9 2 13 1 10 9 9 9 2 16 13 9 11 2 11 2
29 1 3 13 10 9 1 10 9 14 9 9 10 9 1 9 1 9 9 2 16 10 9 16 13 1 9 0 3 2
19 3 2 4 9 11 13 1 9 10 9 12 9 0 1 9 15 14 9 2
15 1 3 2 13 10 9 13 1 9 9 9 1 10 9 2
36 15 2 7 10 9 10 0 1 10 9 16 13 9 1 9 10 9 7 9 15 2 10 13 1 10 9 1 10 9 2 1 10 9 10 0 2
10 11 2 0 1 2 10 9 2 2 2
47 9 11 2 11 2 11 7 11 13 1 9 11 1 10 9 16 13 1 10 9 10 0 2 7 11 13 1 10 9 9 1 9 10 9 1 9 12 2 16 13 14 10 9 1 9 0 2
18 9 11 2 16 13 1 15 2 13 16 3 13 9 11 1 9 15 2
9 11 3 3 13 1 9 10 9 2
66 10 9 2 11 11 2 13 3 2 16 9 11 13 13 14 9 15 1 9 10 9 10 3 2 0 3 1 9 11 2 7 3 15 13 13 3 14 10 9 2 16 16 15 13 2 16 9 10 9 1 10 9 1 9 15 4 13 14 9 10 9 10 3 2 0 2
5 11 2 9 2 2
27 12 10 9 1 9 9 10 9 10 0 13 9 13 1 9 9 0 2 16 13 1 11 7 1 9 0 2
10 3 13 10 9 2 11 2 1 11 2
51 9 10 9 1 11 13 2 16 9 10 9 7 10 9 14 9 9 15 13 1 9 0 7 16 9 10 9 7 10 9 16 1 15 13 9 2 13 1 9 0 7 15 13 1 9 10 9 1 10 9 2
63 9 0 0 13 16 10 9 16 13 3 1 9 15 14 9 9 10 9 13 3 13 9 15 14 9 2 10 9 2 1 9 3 0 2 3 16 16 10 9 13 16 10 9 14 10 9 1 9 15 14 9 10 9 3 13 1 9 14 9 12 9 0 2
52 2 13 1 9 10 9 2 16 9 0 13 13 1 9 9 15 14 10 9 2 16 16 13 1 9 15 13 13 1 9 0 1 9 7 1 9 0 1 11 2 11 7 11 3 13 9 10 9 14 10 9 2
25 1 13 1 15 13 9 9 1 13 1 9 10 9 1 9 0 7 0 0 2 2 13 10 9 2
42 9 0 1 11 2 9 11 11 2 13 16 13 9 0 16 4 13 14 9 15 14 9 0 1 10 9 2 7 3 13 3 14 10 9 10 0 7 13 14 10 13 2
70 11 2 16 15 9 7 9 1 9 1 9 11 7 3 9 10 9 1 9 0 14 10 9 7 10 9 1 10 9 1 9 14 10 9 2 13 16 1 9 10 9 16 13 1 9 10 9 2 13 16 15 13 9 0 1 9 7 1 9 9 1 0 0 3 7 1 10 9 9 2
32 1 16 13 1 10 9 1 12 13 11 9 9 1 9 1 9 11 16 1 11 7 13 1 10 9 10 0 1 9 9 3 2
75 7 1 9 10 9 10 0 10 0 2 16 1 15 13 9 1 12 1 10 9 10 0 1 9 15 2 9 13 14 10 9 7 10 9 10 0 2 9 9 15 10 0 2 7 9 10 9 7 9 15 2 13 11 13 9 1 9 15 1 10 9 10 0 2 7 13 14 10 9 10 9 1 9 0 2
46 9 10 9 13 3 1 9 0 1 2 11 11 2 1 9 7 2 12 2 10 0 2 7 13 1 9 0 3 1 9 2 11 7 3 1 9 9 2 7 1 9 14 9 10 9 2
75 11 13 1 2 10 9 2 16 13 1 9 0 15 1 2 1 13 1 10 9 1 10 9 2 16 15 4 1 9 1 10 9 10 0 14 9 15 2 7 7 7 3 2 4 13 9 1 9 0 16 13 1 3 3 1 10 9 2 10 9 7 9 0 3 13 4 13 1 15 9 7 13 9 15 2
18 11 13 3 16 9 0 0 4 13 1 9 9 10 9 1 9 11 2
22 13 16 11 13 14 9 15 10 3 2 0 14 10 9 3 2 1 9 1 9 0 2
71 1 9 9 2 9 3 0 2 1 9 10 2 9 9 2 10 0 2 15 13 3 16 9 0 14 10 9 13 9 2 9 2 14 9 9 16 13 1 9 1 11 9 2 7 13 1 12 9 14 10 9 1 12 9 2 1 16 3 9 0 3 3 13 1 10 9 1 9 9 15 2
69 9 1 9 2 0 2 2 7 2 9 16 10 9 10 0 14 15 13 1 9 2 16 9 0 13 1 15 2 13 16 1 16 10 10 9 16 13 1 15 9 0 13 1 9 2 15 16 13 1 15 10 9 16 1 10 9 13 2 7 1 9 3 13 1 15 9 9 15 2
13 3 13 9 10 9 1 9 10 9 7 10 9 2
26 7 15 2 11 13 16 3 13 3 3 14 9 9 10 9 14 9 10 9 1 9 9 7 9 0 2
51 4 13 16 10 9 13 0 1 9 1 9 9 1 10 9 10 0 2 3 7 10 9 13 1 9 0 14 9 13 2 9 0 4 13 3 9 2 7 3 13 9 13 9 0 1 9 10 9 10 0 2
5 11 2 9 2 2
39 10 9 10 0 1 9 10 9 1 10 9 13 9 9 3 2 0 2 16 13 1 9 0 1 9 11 1 11 7 1 1 3 3 1 10 9 10 0 2
44 10 9 10 0 2 11 9 16 13 1 15 13 16 10 9 10 0 14 10 9 10 0 2 16 1 9 15 13 11 9 1 10 9 2 13 2 9 0 1 11 1 9 0 2
17 9 9 3 2 0 1 9 1 9 15 10 0 14 11 1 11 2
44 7 12 10 9 10 13 7 10 9 10 3 2 0 10 0 3 13 1 9 13 9 2 13 10 9 1 9 3 2 0 0 2 16 9 9 15 7 9 15 13 0 7 0 2
18 9 1 9 13 10 9 1 11 1 9 0 7 13 10 9 1 15 2
14 9 0 2 0 2 0 3 13 9 0 15 1 11 2
26 10 9 10 3 2 0 13 14 9 15 7 13 3 1 9 10 9 10 0 2 3 10 9 10 0 2
45 9 10 9 16 13 9 1 9 10 9 14 11 11 2 13 1 10 9 10 0 14 10 9 13 1 11 13 1 10 9 10 0 16 1 15 13 1 9 1 9 1 9 10 9 2
41 1 9 10 9 13 9 1 9 9 10 9 16 11 13 1 15 2 11 2 11 1 9 11 7 10 9 1 9 10 9 10 0 2 7 9 1 9 9 10 9 2
32 10 9 10 3 2 0 13 1 10 9 10 0 10 9 0 2 1 9 13 9 1 9 14 11 7 1 9 16 13 1 15 2
13 10 9 13 2 7 16 3 13 9 1 10 15 2
24 2 3 13 1 11 14 10 9 16 3 13 1 15 9 2 2 13 9 16 13 1 10 9 2
32 1 10 9 8 14 9 10 9 13 16 11 2 10 9 7 9 3 13 13 1 11 1 1 10 9 16 13 1 15 1 3 2
38 1 10 9 13 10 9 13 9 0 1 9 1 9 15 14 11 2 7 10 13 16 1 15 13 10 9 13 14 15 2 1 16 13 1 15 10 9 2
15 3 13 9 0 1 9 10 9 2 16 3 13 9 0 2
25 7 15 0 3 9 16 11 2 16 13 1 3 9 1 9 9 10 9 14 11 2 13 13 15 2
11 3 3 4 13 13 14 9 15 14 11 2
32 1 9 11 15 13 16 10 9 10 3 2 0 13 9 1 9 15 2 7 13 16 1 9 0 3 10 9 4 13 9 15 2
9 9 1 10 9 13 14 9 15 2
43 9 13 1 10 9 1 9 10 9 2 3 1 10 9 10 0 2 1 9 15 14 9 10 9 13 14 9 10 9 1 9 10 9 10 0 7 1 9 9 14 9 9 2
25 9 10 9 13 1 9 10 9 1 9 14 9 1 9 11 7 11 2 16 13 1 12 12 9 2
28 9 10 9 13 13 1 9 10 9 1 12 1 11 2 7 13 13 9 14 12 9 1 9 1 9 10 9 2
32 9 10 9 11 11 13 1 9 16 13 13 1 9 10 9 1 9 10 9 7 13 1 15 9 1 9 10 9 2 7 3 2
27 9 9 13 3 16 10 9 13 9 1 9 10 9 1 9 10 9 1 10 9 10 0 7 1 9 9 2
18 1 9 15 2 1 9 9 13 16 1 15 3 1 9 15 13 9 2
31 15 13 14 9 10 9 1 9 9 12 12 9 1 9 1 9 1 9 12 7 1 9 1 9 9 16 10 9 13 3 2
37 9 1 9 13 14 9 10 9 16 2 13 14 10 9 1 9 9 2 2 16 3 2 9 10 9 9 15 1 9 10 9 13 14 9 10 9 2
26 9 10 9 1 9 9 14 9 13 3 1 10 9 2 1 1 10 9 16 13 1 10 9 10 0 2
21 10 9 2 16 13 1 9 0 3 1 10 9 2 13 1 9 1 9 10 9 2
37 9 9 10 9 14 10 11 2 9 11 11 2 11 2 2 13 9 0 1 9 10 9 1 9 10 11 1 9 9 14 9 9 1 9 10 9 2
44 9 11 13 14 9 10 9 16 13 14 9 9 1 9 9 1 9 9 10 9 2 7 15 1 10 9 14 9 10 9 13 1 10 9 14 9 10 9 1 9 1 9 15 2
33 9 11 13 16 9 9 10 9 2 3 4 13 14 10 9 1 9 9 3 1 10 9 10 0 2 7 3 1 9 9 9 0 2
53 9 9 10 9 2 9 11 11 11 2 11 2 2 13 1 9 7 9 0 1 9 9 10 9 11 0 2 7 13 13 1 9 9 14 9 9 15 14 10 9 2 1 9 9 9 10 9 1 10 9 10 0 2
48 11 13 16 2 1 10 9 15 1 9 10 9 14 9 10 9 2 16 1 9 13 14 10 9 10 13 2 4 13 14 9 10 9 7 13 9 1 10 9 2 1 2 9 9 10 9 2 2
64 15 13 16 1 9 15 13 1 9 0 14 9 10 9 1 9 1 10 9 16 1 15 13 10 10 9 16 1 9 15 13 9 1 10 9 10 0 14 9 2 7 13 1 2 9 15 14 9 15 10 0 14 10 9 2 7 9 9 15 1 9 10 9 2
10 11 2 0 1 2 10 9 2 2 2
29 9 11 2 11 11 2 13 3 1 11 9 9 9 2 16 1 9 15 13 9 3 2 9 1 9 15 1 11 2
39 10 9 13 14 10 9 1 12 10 9 1 9 0 14 9 2 7 15 13 1 9 9 1 9 0 2 16 13 14 9 15 14 11 7 11 1 9 0 2
31 10 9 2 1 9 14 12 9 2 13 9 16 9 0 14 11 7 11 13 3 0 1 13 14 10 9 14 12 10 9 2
22 3 7 2 13 9 10 9 3 9 12 1 9 2 7 9 10 9 3 9 1 9 2
30 1 9 10 9 13 11 7 11 1 9 9 0 1 9 10 9 2 10 9 2 9 10 9 2 9 10 9 7 3 2
21 11 13 9 13 1 9 11 9 0 7 0 0 2 16 9 15 10 0 3 13 2
34 1 9 1 15 13 11 1 9 0 13 14 9 10 9 10 0 1 9 2 11 7 13 9 0 1 12 12 10 9 16 13 1 11 2
17 10 9 10 0 1 10 9 10 15 3 13 1 1 12 12 11 2
36 9 15 14 11 1 11 13 1 9 0 3 2 7 13 1 15 9 0 1 10 9 1 15 16 10 9 10 0 13 1 9 0 1 9 11 2
40 9 1 15 13 3 16 9 10 9 2 11 11 2 13 1 9 15 10 0 2 11 2 11 11 2 1 9 1 10 9 11 2 1 9 9 2 11 3 2 2
20 11 13 9 9 15 14 11 2 7 3 15 13 13 1 15 9 1 9 0 2
18 11 1 9 15 13 14 11 1 9 15 1 11 2 9 1 9 11 2
26 1 9 0 1 10 9 11 13 11 1 10 9 2 7 12 13 1 15 1 9 2 11 2 11 2 2
27 1 11 13 10 9 10 0 1 13 14 11 1 10 9 10 0 1 9 1 9 15 14 10 9 10 0 2
23 1 9 10 9 13 11 2 16 9 1 9 15 13 9 0 7 13 2 16 13 9 0 2
20 15 13 2 16 11 13 9 9 16 13 9 0 1 3 16 13 1 15 9 2
34 11 1 9 15 13 2 16 9 15 13 1 11 1 9 9 3 2 7 13 1 9 9 15 1 16 3 15 13 1 9 15 14 11 2
10 11 11 2 0 1 2 10 9 2 2
46 11 11 2 9 2 9 10 9 2 14 9 10 9 11 11 11 2 13 1 9 15 1 10 9 12 12 9 3 1 9 10 9 1 15 13 3 3 13 3 10 2 11 11 11 2 2
18 1 10 9 12 12 13 11 9 10 12 9 9 0 9 12 12 9 2
28 15 13 12 12 9 1 9 12 2 7 13 1 15 1 9 16 9 15 10 0 13 10 0 3 1 9 11 2
42 3 13 10 2 11 2 2 16 1 9 14 12 9 14 15 13 11 1 11 2 9 9 15 7 9 15 10 13 2 13 16 9 10 9 13 1 15 3 12 9 3 2
34 1 9 9 9 7 9 1 15 13 10 9 2 13 9 1 10 9 10 0 14 11 9 9 12 7 3 12 9 1 10 9 10 0 2
24 9 9 9 0 1 10 9 13 1 10 9 16 9 10 9 14 11 1 10 9 13 12 9 2
20 9 14 10 3 2 9 13 14 9 10 9 1 2 13 7 13 9 0 2 2
13 9 9 15 14 11 4 13 3 2 3 3 3 2
29 1 10 13 2 15 13 1 12 9 9 14 9 1 9 14 9 16 13 1 9 15 2 7 13 1 12 12 9 2
30 1 10 9 10 0 8 8 10 9 13 2 3 13 2 11 11 2 1 9 11 2 1 1 9 16 13 1 10 9 2
32 11 16 13 1 3 9 10 9 10 12 1 10 9 2 13 9 7 9 1 11 2 1 10 9 10 0 7 1 11 10 0 2
18 2 10 9 13 1 10 9 9 10 9 2 2 13 2 11 11 2 2
23 9 10 9 10 9 13 1 12 12 9 1 12 1 12 12 1 12 2 13 1 10 9 2
25 9 1 9 9 13 12 12 11 2 12 12 9 2 1 12 12 11 2 12 12 9 2 1 12 2
25 9 9 1 9 10 9 13 1 12 12 11 2 12 12 9 2 1 12 12 2 12 12 9 2 2
31 10 9 1 9 10 9 10 0 13 1 12 12 11 2 12 12 9 2 1 9 1 12 12 2 12 12 9 2 1 12 2
53 10 9 13 1 9 16 1 15 13 16 2 10 9 10 0 1 11 7 9 9 9 0 0 1 11 9 15 16 9 10 9 13 1 10 9 3 1 9 0 16 13 1 10 9 7 13 1 9 1 10 9 2 2
20 2 9 11 7 11 1 9 15 13 1 10 9 10 0 2 2 13 10 9 2
28 11 11 13 3 1 9 9 16 13 1 9 9 2 9 7 9 1 9 0 7 9 0 2 0 2 7 0 2
19 10 9 13 1 2 9 10 9 11 11 1 9 10 9 1 11 2 11 2
49 11 2 9 9 12 2 13 1 15 14 11 11 11 16 13 14 9 9 10 9 1 16 10 9 10 0 10 0 2 13 9 10 9 2 7 10 9 13 9 1 9 3 2 9 10 9 16 13 2
26 2 15 13 16 10 9 10 0 13 9 1 9 9 9 15 12 2 2 13 10 9 1 9 10 9 2
12 8 8 14 11 13 10 0 3 1 9 11 2
31 9 15 14 11 11 11 13 12 9 3 1 12 9 1 9 10 9 7 13 1 9 10 9 14 11 11 7 9 10 9 2
13 11 15 13 13 9 7 13 1 10 9 14 11 2
15 11 13 16 13 1 15 9 1 10 9 1 9 10 9 2
23 11 13 16 9 15 10 0 13 13 9 1 10 9 1 10 9 7 13 10 9 0 0 2
11 9 11 13 1 11 12 9 1 10 9 2
29 12 10 9 13 16 1 9 4 11 13 14 10 9 14 10 9 10 0 10 0 2 16 9 13 13 1 15 3 2
37 10 9 11 13 16 15 13 0 1 10 9 13 1 9 9 0 14 9 9 10 9 2 1 11 13 1 9 9 7 9 9 1 9 9 7 0 2
36 7 7 7 11 11 13 10 9 10 0 10 0 16 13 4 13 1 15 14 10 9 3 2 3 13 1 10 9 7 13 14 10 9 1 15 2
38 9 0 1 11 2 11 13 16 9 11 13 9 9 1 10 9 10 0 16 13 1 16 13 10 9 1 10 9 1 10 9 1 9 10 9 1 11 2
20 8 8 14 11 13 14 9 15 10 0 1 9 15 2 1 15 13 9 0 2
30 9 9 9 2 9 9 0 7 9 9 13 14 9 15 14 11 1 9 16 13 1 9 15 1 9 3 1 9 15 2
31 10 9 10 0 16 13 13 1 15 9 1 9 0 7 13 13 1 15 1 13 1 9 15 2 9 0 0 14 9 9 2
14 10 9 13 14 15 7 13 14 15 1 9 10 9 2
17 10 9 1 9 10 9 13 1 10 9 14 9 9 1 9 11 2
5 2 15 3 0 2
8 3 13 1 9 1 10 15 2
9 3 15 13 14 10 9 10 0 2
11 15 3 4 3 2 2 13 12 1 15 2
26 0 13 14 11 1 2 9 0 14 15 13 10 9 10 0 3 1 10 9 14 10 9 10 0 2 2
32 1 9 9 10 9 1 9 9 7 0 16 13 1 11 1 9 15 13 11 1 9 0 3 16 3 13 16 13 1 15 9 2
48 10 9 10 0 2 9 1 10 9 11 13 1 9 14 9 7 9 9 1 9 10 9 10 0 13 14 9 10 9 1 9 0 1 10 9 10 0 1 10 9 1 12 9 1 3 12 9 2
22 9 9 9 7 9 1 10 9 10 0 13 1 9 15 7 13 13 15 1 10 9 2
13 1 1 15 13 12 10 9 1 11 7 1 11 2
23 1 9 10 9 1 12 9 15 16 1 9 11 13 12 9 9 1 9 10 9 10 0 2
8 9 0 0 13 1 9 11 2
19 1 1 10 15 13 11 1 9 0 0 16 13 1 3 9 11 1 11 2
23 10 9 13 1 9 0 1 9 10 9 7 10 9 7 9 16 13 1 9 3 2 0 2
4 2 11 2 2
24 9 0 2 12 1 9 15 2 13 1 9 11 1 9 11 1 9 10 9 1 9 2 9 2
14 10 9 13 1 9 10 9 12 9 1 9 10 9 2
18 9 0 13 14 10 9 10 0 14 10 9 7 10 9 13 1 15 2
10 1 9 11 13 9 1 9 10 9 2
21 1 9 11 13 9 9 2 7 1 9 11 1 10 9 13 1 10 9 9 13 2
18 1 12 10 9 10 0 13 9 9 14 13 10 9 16 13 1 9 2
17 7 15 13 9 7 13 9 0 9 12 1 10 9 1 10 9 2
31 10 9 13 1 12 9 1 9 7 13 3 1 15 9 2 16 16 10 9 1 9 11 7 1 9 11 13 1 9 15 2
29 1 9 11 13 1 10 9 9 2 1 9 9 1 9 9 2 7 13 1 9 10 9 2 13 10 9 10 0 2
15 9 9 11 13 16 13 13 1 3 3 12 1 10 9 2
20 2 1 16 15 13 1 10 9 10 12 2 15 4 13 3 9 2 2 13 2
9 11 2 9 2 9 2 9 2 2
21 12 9 0 16 13 3 9 14 9 10 9 10 0 13 1 9 10 9 10 0 2
27 12 10 9 7 9 9 15 14 10 9 16 13 1 9 15 1 11 1 11 13 1 16 9 1 15 13 2
27 11 11 2 9 0 14 9 9 11 2 13 1 1 9 10 9 16 15 13 1 9 0 7 13 9 9 2
23 1 11 13 9 1 9 1 9 2 9 10 9 7 10 9 2 16 3 13 13 1 3 2
26 1 10 9 13 16 10 9 13 13 1 10 9 13 2 1 9 10 9 10 0 1 9 7 9 9 2
20 13 1 15 10 9 13 1 10 9 7 1 10 9 2 2 13 1 10 9 2
31 12 10 9 13 1 10 9 1 9 9 15 10 13 7 13 2 2 7 13 14 9 15 13 15 1 9 1 9 11 2 2
31 10 9 13 1 9 11 13 14 10 10 9 10 0 2 13 9 1 10 9 10 0 7 13 14 10 9 1 9 0 13 2
34 3 13 10 9 16 11 13 14 10 10 9 1 11 1 16 10 9 13 1 9 0 7 9 9 0 16 13 1 11 13 9 14 9 2
23 1 11 16 13 13 12 9 9 0 16 13 1 9 9 7 13 14 10 9 13 1 11 2
8 15 13 7 3 13 1 11 2
16 9 9 10 9 7 10 9 13 3 14 9 15 14 12 15 2
28 10 9 1 11 7 1 1 15 13 1 10 9 10 0 16 13 14 10 9 1 9 1 9 9 0 1 9 2
32 1 11 13 1 11 9 1 10 9 10 0 7 10 9 10 0 13 1 3 13 14 10 9 1 10 9 16 13 1 9 13 2
8 9 10 9 0 13 1 9 2
4 2 11 2 2
22 1 9 9 16 13 1 9 11 1 10 9 1 9 9 2 10 0 11 13 9 9 2
18 9 1 9 12 13 7 12 9 13 2 1 15 3 12 1 9 0 2
27 10 9 13 9 1 11 2 16 13 1 11 1 12 9 7 13 1 9 11 11 2 16 0 1 9 11 2
11 3 13 1 12 9 1 10 9 1 11 2
40 1 1 9 12 13 12 10 9 2 16 0 1 9 9 1 11 2 1 9 9 2 11 11 2 13 10 9 7 13 1 13 10 9 2 14 15 1 9 15 2
29 1 10 9 13 1 15 9 12 9 2 9 7 9 2 9 2 16 9 15 13 1 10 9 7 13 1 10 9 2
23 10 9 10 12 13 9 3 7 1 10 16 13 2 1 9 1 15 2 9 12 13 3 2
23 12 1 10 9 13 1 9 10 13 11 9 10 9 7 12 1 15 1 11 9 2 9 2
25 12 9 13 3 1 9 10 13 7 12 3 13 1 9 10 13 11 9 2 9 7 11 10 9 2
5 9 15 13 3 2
30 9 12 13 7 12 13 3 1 9 9 0 16 13 1 9 11 1 10 9 1 9 11 9 2 9 1 9 10 9 2
15 10 9 7 10 9 13 1 9 9 1 9 11 9 9 2
36 11 11 2 9 12 2 1 9 9 2 13 1 11 2 16 9 11 1 15 13 1 9 1 9 15 2 13 1 9 9 2 1 9 9 9 2
29 10 9 2 11 9 11 1 9 11 2 7 9 0 11 11 2 9 12 2 13 3 7 13 1 9 11 1 11 2
22 10 9 13 9 16 10 9 2 16 1 9 15 9 9 10 9 3 2 13 1 9 2
9 10 9 13 1 9 12 1 9 2
30 12 9 13 1 9 9 1 9 11 1 9 2 14 9 0 13 9 9 1 9 11 7 13 1 9 16 13 1 15 2
13 9 12 13 1 9 0 7 10 9 1 9 0 2
17 10 9 13 1 9 10 13 11 7 9 11 2 11 2 1 11 2
21 9 9 12 1 11 2 13 3 1 9 11 1 9 2 1 9 9 1 10 9 2
28 10 9 13 14 10 9 1 9 0 9 12 1 9 9 10 9 2 16 3 1 9 9 7 1 9 9 13 2
15 9 0 13 1 9 12 1 9 2 9 2 13 1 9 2
24 9 9 0 14 9 9 0 13 14 15 1 9 0 1 10 9 10 0 11 1 9 2 9 2
15 1 10 9 2 16 13 1 9 15 2 3 13 9 9 2
43 9 10 9 14 9 9 11 2 16 1 9 9 10 9 2 13 13 14 9 15 14 11 11 1 9 15 1 9 10 9 2 16 13 1 9 15 1 9 0 14 12 9 2
35 1 2 3 13 10 9 13 9 14 10 9 10 0 14 9 10 9 14 10 9 2 7 13 1 9 15 1 9 15 14 11 1 9 15 2
43 11 2 16 13 1 9 9 10 9 10 0 9 1 13 1 9 15 10 0 14 9 10 9 1 10 9 10 0 14 9 11 2 3 13 1 10 9 16 13 1 9 11 2
41 1 15 13 1 9 9 10 9 9 1 15 2 16 1 15 15 4 13 1 9 1 9 1 9 12 9 2 1 9 16 13 9 0 16 13 14 10 9 1 15 2
25 9 9 10 9 13 4 13 14 9 15 1 9 1 9 2 7 13 9 2 12 14 9 10 9 2
30 9 9 10 9 14 9 9 11 11 9 2 13 1 11 2 1 15 13 1 15 9 0 16 15 13 13 1 10 9 2
14 9 10 9 13 1 9 15 14 11 9 1 10 9 2
22 11 3 3 13 1 9 10 9 1 9 11 11 2 1 15 13 1 13 1 9 15 2
16 1 1 3 13 16 10 9 13 14 9 15 1 13 1 15 2
28 1 9 11 13 16 9 10 9 3 13 14 10 10 9 16 13 1 15 2 16 16 9 1 10 15 3 13 2
20 10 9 13 9 13 1 15 16 1 9 10 9 13 9 16 4 13 9 15 2
44 8 8 10 9 13 9 9 10 9 14 9 11 2 1 9 15 11 11 2 10 9 9 11 11 2 7 9 9 9 11 2 16 15 9 2 9 14 10 9 2 9 11 11 2
21 9 10 9 7 9 9 2 11 13 3 1 9 10 9 1 3 1 12 12 9 2
15 1 9 15 14 11 3 13 9 0 1 10 9 16 13 2
9 9 9 13 1 16 13 9 15 2
30 13 9 9 1 9 0 3 2 7 13 9 1 9 12 9 2 16 3 13 3 1 9 10 9 2 7 13 1 9 2
16 1 9 9 10 9 3 13 9 0 1 9 10 9 14 11 2
12 3 13 13 1 15 14 10 10 9 10 0 2
30 1 9 10 9 13 1 9 10 9 9 13 14 10 9 7 7 13 3 9 9 1 10 9 10 0 14 9 10 9 2
33 1 10 9 10 0 13 9 10 9 13 14 10 9 7 13 1 15 14 10 9 13 9 0 2 1 9 13 14 11 1 9 15 2
21 3 13 10 9 10 0 13 14 9 10 9 1 9 12 7 14 9 9 10 9 2
24 11 11 13 1 9 2 2 13 1 9 16 13 3 7 15 13 1 15 13 1 9 1 9 2
17 10 9 14 15 13 9 9 0 16 13 14 10 10 9 1 15 2
8 1 1 15 15 3 13 13 2
8 15 3 13 1 9 10 9 2
7 15 3 0 1 9 15 2
15 13 1 10 10 9 2 13 9 0 1 13 9 0 2 2
3 3 4 2
26 1 10 9 13 9 16 1 9 10 9 14 10 9 13 3 16 9 3 13 1 10 9 1 9 11 2
19 1 3 13 10 9 16 3 1 9 7 1 9 0 4 13 1 9 9 2
10 4 16 13 9 13 9 9 0 3 2
17 9 10 9 10 0 2 13 13 1 10 9 1 9 3 2 9 2
19 10 9 1 9 9 16 13 1 9 2 4 13 9 16 13 0 1 9 2
18 9 12 2 4 3 16 9 13 1 10 9 3 1 9 7 1 9 2
29 1 2 3 4 13 7 15 13 16 3 13 1 10 9 9 7 9 14 9 7 9 0 14 10 9 15 1 15 2
18 10 9 10 0 14 9 1 9 13 9 0 1 9 9 1 10 15 2
29 1 2 9 10 9 10 0 2 0 1 10 9 16 7 15 13 1 15 1 9 2 15 4 13 1 15 1 9 2
38 13 9 16 1 10 9 16 13 1 9 10 9 10 9 13 9 1 10 10 9 10 0 16 13 1 2 9 10 9 10 0 14 9 0 9 9 0 2
22 0 16 15 9 3 1 9 16 3 13 1 10 9 2 1 10 9 10 0 10 0 2
31 15 13 3 9 14 9 0 16 13 1 10 9 10 0 7 4 13 7 3 3 13 14 15 7 13 1 13 14 9 15 2
2 3 2
19 10 9 10 0 10 15 2 13 0 9 7 9 1 9 15 14 10 9 2
39 15 3 13 9 9 0 14 9 0 2 1 13 14 9 15 10 0 14 10 9 7 13 9 9 10 9 1 9 16 13 9 1 15 1 10 9 10 0 2
46 15 13 16 3 16 13 1 10 9 10 15 2 13 1 10 10 9 16 13 1 15 7 9 1 15 16 13 9 1 15 3 1 11 2 13 13 1 9 15 7 1 10 9 14 15 2
33 1 9 1 10 9 0 9 14 9 2 9 7 9 2 16 4 1 13 10 9 13 7 13 14 10 9 10 0 16 13 1 15 2
10 11 2 0 1 2 10 9 2 2 2
50 10 9 10 0 11 11 2 16 13 1 10 9 16 13 14 9 15 1 16 13 14 9 9 15 14 9 15 1 10 9 10 0 2 13 3 1 10 9 10 0 1 9 9 15 11 2 1 9 11 2
33 15 13 14 9 15 1 9 2 9 1 9 9 10 9 10 0 2 9 11 2 2 16 15 7 9 15 9 1 15 15 12 9 2
40 15 13 2 16 15 13 16 13 1 9 10 9 14 15 13 1 10 9 10 15 2 13 1 2 9 15 7 13 2 2 7 13 2 9 0 2 1 10 9 2
28 10 9 16 13 14 11 2 11 11 13 3 2 16 3 15 13 9 1 9 1 11 7 1 9 0 1 15 2
35 15 13 2 16 1 10 9 1 10 9 13 2 9 15 2 2 16 7 3 15 2 9 0 7 0 13 13 15 14 15 1 9 0 2 2
37 11 2 9 9 12 1 9 10 9 2 9 10 9 10 0 2 13 1 9 11 16 13 14 11 11 2 1 10 9 10 0 10 0 3 1 11 2
51 9 11 13 10 9 10 0 3 14 10 9 1 10 9 1 11 2 7 15 13 1 2 9 1 9 0 1 9 15 10 0 14 2 11 11 11 2 2 7 1 9 10 9 0 2 10 9 2 11 2 2
33 10 9 10 0 14 9 10 9 13 1 9 9 14 9 11 1 9 9 15 14 11 1 10 9 10 0 7 1 10 9 10 0 2
37 9 0 1 11 13 2 16 10 9 10 15 2 1 9 10 9 10 0 14 11 7 16 3 1 9 15 2 13 1 10 9 10 0 1 9 15 2
14 15 13 1 15 9 0 1 9 15 7 1 1 15 2
31 1 9 10 11 10 0 1 11 2 16 11 13 12 1 9 15 2 13 1 9 11 10 9 10 0 9 0 1 10 9 2
42 9 1 10 9 10 0 14 11 13 1 9 1 9 9 15 14 11 2 7 13 1 9 7 9 13 1 11 9 1 11 2 3 1 16 13 1 9 2 1 9 11 2
42 9 9 10 9 14 11 2 10 9 10 0 11 11 2 13 1 9 0 1 11 2 16 2 11 13 9 10 2 3 0 2 16 10 9 0 0 13 1 15 3 2 2
7 11 3 3 13 1 11 2
39 10 9 1 9 15 2 16 13 1 10 9 1 12 9 0 2 13 3 1 9 11 1 11 11 2 1 9 10 9 10 0 14 10 9 10 0 1 11 2
22 11 13 9 9 15 14 11 1 11 2 1 9 10 9 10 0 1 10 9 1 12 2
26 10 9 13 14 11 2 16 15 3 3 13 1 9 15 14 11 1 11 7 1 11 9 16 11 13 2
60 1 9 0 1 11 1 9 15 13 11 1 9 9 0 1 11 2 16 15 9 0 14 11 2 7 13 1 10 9 1 10 9 10 0 2 7 2 15 13 16 15 13 14 10 9 14 9 0 2 9 11 2 16 15 4 13 14 11 2 2
40 11 13 2 2 1 15 9 2 1 9 11 2 4 9 13 0 1 9 0 7 15 3 13 0 1 9 10 9 1 11 2 16 14 15 15 13 1 9 0 2
32 15 13 2 16 13 10 9 2 7 9 2 7 10 9 2 7 15 13 16 1 9 15 14 9 13 9 15 14 9 1 9 2
14 7 15 13 3 1 10 9 10 0 7 1 11 2 2
34 1 9 10 9 13 10 9 10 0 2 16 15 13 16 2 1 9 15 14 9 13 9 15 14 9 2 7 15 13 16 15 13 13 2
33 2 10 9 10 0 2 2 13 11 2 2 13 4 13 2 16 7 3 15 13 9 0 7 0 13 15 14 15 1 9 0 2 2
35 3 13 11 2 9 15 10 3 2 0 11 2 7 9 9 10 9 14 15 11 11 2 1 9 9 11 1 9 10 11 10 0 14 11 2
45 9 9 10 11 2 11 11 2 13 2 16 1 10 9 1 9 15 14 11 13 13 2 3 2 9 14 9 10 9 2 16 13 14 15 10 2 3 0 1 9 2 2 1 11 2
41 9 9 11 2 2 11 11 2 2 13 1 9 15 10 0 9 3 2 0 1 11 2 16 13 2 2 15 13 1 13 14 11 11 2 7 13 13 1 9 11 2
7 15 4 13 9 0 2 2
34 9 11 11 2 11 2 13 9 0 1 9 10 9 2 1 9 1 9 10 9 7 10 9 13 14 9 10 9 1 9 15 10 0 2
35 9 11 13 16 3 4 16 9 9 15 16 13 1 9 9 15 2 9 1 9 2 13 13 9 2 1 3 2 9 9 1 2 11 2 2
25 1 9 15 2 10 9 9 2 9 13 1 3 12 1 9 15 2 12 1 15 1 9 9 12 2
18 9 15 13 13 1 12 9 1 9 14 12 12 9 1 2 11 2 2
40 11 11 13 1 9 11 2 13 9 1 13 1 10 9 10 0 13 14 10 9 7 13 16 16 13 1 9 0 16 13 1 9 9 11 3 1 9 15 2 2
29 9 10 9 11 11 7 9 10 9 11 11 13 13 9 1 10 9 16 13 10 12 1 9 1 9 9 9 9 2
15 3 13 9 10 9 13 14 10 9 16 13 14 11 11 2
18 11 13 1 9 14 11 11 2 3 9 9 9 10 9 7 10 9 2
14 11 13 13 1 9 14 9 9 10 9 2 11 11 2
35 7 9 15 14 11 1 9 15 14 11 2 13 16 10 12 1 10 9 13 1 10 9 14 9 15 2 7 9 10 9 13 1 10 12 2
34 9 11 13 12 9 2 1 15 12 9 9 10 9 2 9 10 9 11 11 2 9 10 9 11 11 2 7 9 9 10 9 11 9 2
35 1 9 10 9 12 9 1 10 9 2 9 16 13 1 10 9 7 10 0 1 9 10 9 11 11 2 7 9 10 9 10 0 11 9 2
21 3 13 1 10 9 1 9 10 9 11 11 11 2 7 9 15 14 11 11 11 2
23 1 2 9 9 11 13 1 10 9 11 11 2 3 10 9 1 9 10 9 1 10 9 2
27 9 11 2 11 11 2 13 3 16 9 10 9 13 9 2 16 1 15 13 9 10 9 14 12 10 9 2
10 11 7 11 13 13 3 1 10 9 2
21 11 13 16 15 13 16 10 9 13 1 2 9 9 10 9 10 0 14 10 9 2
23 9 9 2 3 13 1 9 1 9 10 9 2 11 11 2 13 14 9 11 1 9 0 2
38 1 9 15 13 9 2 3 16 11 13 1 9 9 9 16 16 13 1 10 9 2 7 13 1 9 10 9 13 14 10 9 1 9 10 9 10 0 2
24 1 9 15 1 11 13 9 2 3 16 3 13 9 0 1 9 15 7 9 15 14 9 11 2
18 9 15 13 1 9 1 9 13 1 9 7 1 9 13 1 9 0 2
61 1 9 15 2 1 9 11 1 9 9 2 13 9 2 3 1 10 9 1 9 9 2 16 13 9 0 1 2 9 9 16 13 1 9 15 1 9 9 16 4 13 1 9 15 14 9 7 1 9 15 2 7 1 9 1 9 9 1 15 2 2
38 9 15 14 10 9 11 11 2 16 13 3 1 10 9 1 9 10 9 1 11 1 9 9 0 1 11 2 13 13 3 7 15 3 13 1 9 9 2
20 11 13 3 1 12 9 1 9 11 9 2 9 7 3 13 1 9 10 9 2
23 1 9 10 9 3 13 11 7 9 15 14 9 10 9 2 16 16 13 10 9 13 3 2
18 10 13 9 11 11 11 9 12 1 11 2 13 1 9 15 7 13 2
43 11 2 9 11 7 9 1 9 9 14 10 9 2 13 1 11 1 9 9 10 9 16 13 1 10 9 1 3 10 9 1 9 10 9 2 1 10 9 7 1 9 11 2
30 3 1 1 9 12 1 10 9 2 13 11 1 12 1 9 15 1 9 10 9 1 9 10 9 2 1 9 9 0 2
19 3 13 1 9 9 1 9 10 9 12 9 0 2 14 9 0 1 9 15
25 9 15 1 10 9 9 13 1 15 2 13 14 15 1 10 9 7 13 14 10 9 1 9 15 2
25 2 15 13 1 9 11 2 2 13 3 9 2 2 13 14 15 1 10 9 7 13 14 10 9 2
10 10 9 13 7 13 13 14 10 9 2
5 9 13 3 2 2
36 12 10 9 10 0 16 13 1 10 9 13 1 10 13 1 9 9 10 9 10 0 7 13 1 9 1 3 9 2 11 2 16 1 9 15 2
9 10 13 13 1 9 0 7 13 2
16 1 9 15 13 16 15 9 11 16 13 1 9 11 2 11 2
18 1 9 13 13 9 1 11 7 3 1 10 9 13 1 9 1 11 2
31 15 13 1 9 9 1 9 10 9 2 13 9 0 7 3 13 3 1 9 9 10 9 2 13 1 9 10 9 7 13 2
24 16 13 12 10 9 1 9 10 9 13 10 13 14 10 9 1 9 15 7 13 14 11 11 2
15 1 9 0 13 1 10 9 9 9 0 7 9 14 9 2
18 15 13 9 0 1 11 11 2 16 13 9 0 7 13 14 9 15 2
14 11 13 1 11 9 2 9 14 15 1 9 7 13 2
31 1 9 0 1 9 9 15 13 3 1 9 10 9 2 3 13 9 1 9 10 9 7 9 10 9 16 13 1 10 9 2
25 9 15 14 10 13 16 13 1 10 9 13 0 2 7 3 15 13 1 11 9 9 3 13 9 2
33 10 9 7 9 15 3 13 9 9 7 3 1 10 9 13 9 10 9 9 9 11 11 1 10 9 1 10 9 13 1 9 15 2
11 1 10 13 3 13 9 0 2 7 0 2
32 15 13 3 1 9 10 11 2 16 13 13 3 13 1 9 0 2 7 13 1 9 9 7 3 3 13 10 9 1 9 15 2
11 11 13 16 13 4 13 9 1 10 15 2
14 15 13 14 10 9 14 10 9 16 13 1 10 9 2
14 2 7 3 3 13 13 7 13 14 10 13 2 13 2
33 11 13 13 3 1 11 7 10 10 9 3 13 9 9 2 7 16 13 16 13 9 16 10 9 13 13 3 7 15 13 13 9 2
38 10 9 13 16 10 9 13 1 9 15 14 10 9 16 1 11 1 9 11 2 1 13 9 16 13 9 15 1 11 1 10 9 10 0 7 1 9 2
15 1 10 9 13 10 9 7 10 10 9 13 14 10 9 2
15 15 10 9 10 12 14 9 9 1 15 9 1 12 9 2
20 10 9 1 9 10 9 1 10 9 13 9 13 9 0 1 9 0 1 9 2
21 12 1 15 13 2 10 9 2 2 9 16 13 14 9 10 9 10 0 14 15 2
36 9 10 2 11 2 13 1 9 10 9 1 9 9 1 10 9 2 11 2 7 1 9 10 9 1 9 0 1 10 9 1 10 9 10 0 2
51 10 9 16 13 14 9 10 9 13 16 9 0 16 13 1 9 15 1 12 9 2 4 13 1 15 9 0 0 1 10 9 10 9 7 13 1 10 9 10 0 7 10 9 14 9 10 9 1 10 9 2
39 11 13 1 9 10 9 1 10 9 2 1 16 13 1 12 9 2 9 0 1 10 9 10 0 2 7 9 0 14 9 9 10 9 1 10 9 1 15 2
21 1 9 10 9 13 9 11 2 10 9 1 9 0 2 9 10 9 7 9 13 2
22 12 10 9 16 13 13 1 10 9 12 9 1 9 2 9 2 9 2 7 9 0 2
37 10 9 16 13 1 10 9 13 9 9 0 7 0 2 7 9 15 0 2 16 13 1 9 0 1 9 15 2 7 13 9 0 1 9 10 9 2
36 1 9 9 10 9 1 9 0 1 10 9 1 9 0 2 10 9 16 13 13 1 9 0 1 15 13 9 0 1 9 9 9 1 10 9 2
24 10 13 9 11 11 13 3 13 1 9 15 7 1 9 10 9 16 13 1 15 1 12 9 2
30 10 9 13 1 9 10 9 10 0 14 9 10 9 1 9 9 0 7 13 1 9 9 1 9 7 1 9 1 9 2
31 1 10 9 10 0 13 9 7 9 1 10 10 9 1 9 15 7 13 9 16 13 9 13 1 10 9 16 13 1 15 2
22 9 11 9 16 13 7 13 1 9 9 1 9 7 1 9 1 9 9 2 3 13 2
25 9 0 9 0 11 11 2 16 13 7 13 1 9 9 1 9 7 1 9 1 9 9 3 13 2
49 10 13 10 0 3 10 9 9 9 11 11 16 13 7 13 1 9 9 1 9 7 1 9 1 9 9 2 13 3 16 10 9 14 10 9 14 15 13 3 13 1 9 10 9 7 9 10 9 2
34 1 9 15 1 9 0 15 13 1 9 2 7 1 10 9 7 9 10 9 2 10 9 13 3 13 1 9 10 9 10 0 1 9 2
17 1 15 2 13 3 11 16 3 1 10 9 13 10 9 10 0 2
48 9 0 9 11 11 2 10 0 16 13 1 9 9 14 9 1 10 9 7 9 1 9 9 2 13 13 1 9 9 9 15 9 10 9 11 11 2 7 1 9 15 3 13 10 9 10 0 2
30 7 3 13 9 11 9 1 9 10 9 10 0 1 9 2 15 13 1 9 10 9 10 3 0 3 16 13 1 9 2
35 3 10 9 10 0 13 3 13 1 8 10 9 2 7 1 9 16 15 1 10 9 16 13 13 9 2 13 3 10 9 10 0 9 0 2
55 7 1 9 9 11 11 10 9 1 9 11 11 13 1 9 15 1 9 10 9 7 9 10 9 2 7 10 9 1 16 13 10 9 2 13 14 10 9 1 16 13 1 15 16 1 11 13 1 9 15 7 15 13 9 2
11 7 3 9 15 14 9 9 11 11 13 2
57 1 10 9 10 0 13 1 10 9 10 0 14 9 10 9 1 10 10 13 1 10 9 10 0 16 9 15 13 1 9 11 11 1 10 9 10 0 2 16 13 3 14 10 9 7 13 1 10 9 14 9 11 3 9 11 11 2
35 1 10 16 13 1 9 11 11 7 1 3 9 11 11 2 10 9 10 0 10 0 3 13 7 13 1 9 10 9 1 10 9 14 15 2
30 9 10 9 1 9 0 1 10 9 10 0 11 2 9 11 11 2 13 1 9 9 11 7 11 11 0 1 9 12 2
15 10 9 1 9 12 12 9 0 13 1 9 9 9 0 2
21 9 11 13 9 12 1 9 9 10 9 10 0 14 9 10 9 2 9 11 11 2
24 10 9 13 1 15 1 9 9 15 7 9 15 10 0 7 10 0 1 9 10 9 10 0 2
47 9 11 13 16 10 9 13 1 10 9 1 9 9 0 16 13 1 9 9 1 9 7 9 9 2 7 1 9 1 9 9 2 1 1 9 10 9 1 9 1 9 9 7 9 9 0 2
13 15 10 9 10 12 16 10 9 13 1 9 9 2
47 1 10 9 13 14 10 9 9 11 11 1 10 9 10 0 2 11 2 2 13 11 11 2 1 9 10 9 1 9 10 9 1 9 11 11 7 9 11 11 1 9 10 13 11 1 11 2
10 11 2 0 1 2 10 9 2 2 2
63 9 9 1 11 13 16 10 9 11 13 14 10 9 10 0 1 9 10 9 14 11 1 11 1 9 10 9 2 1 16 10 9 10 0 1 11 13 2 7 1 9 10 9 10 0 2 16 1 15 13 9 0 1 9 9 9 1 9 11 7 9 11 2
48 9 10 9 2 16 13 3 1 9 1 10 9 10 0 1 9 10 9 2 13 16 4 13 16 11 13 13 9 0 1 9 10 9 10 0 10 0 1 11 2 16 13 3 3 1 9 11 2
46 1 11 1 11 3 13 9 9 3 0 1 9 7 1 9 11 13 9 10 9 2 16 1 9 15 13 12 12 7 3 12 14 9 1 9 10 9 1 9 11 2 1 9 10 9 2
61 10 9 14 9 1 9 9 1 11 2 3 2 13 16 9 0 14 9 11 13 1 1 9 11 2 11 14 10 9 10 0 2 3 16 0 9 0 1 10 9 1 10 0 10 0 16 1 9 9 0 1 9 11 1 9 9 15 14 10 9 2
14 11 13 3 13 9 1 9 10 9 14 11 1 11 2
30 9 10 9 14 11 2 11 11 2 13 3 16 10 9 13 13 13 14 10 9 16 13 1 10 9 1 9 14 9 2
30 9 15 13 9 1 9 10 9 2 16 13 1 1 9 16 1 9 15 13 14 10 9 16 13 1 11 1 9 0 2
25 9 0 13 16 9 10 9 13 13 14 10 9 10 0 1 11 7 13 16 9 0 4 13 3 2
36 9 0 4 16 10 9 0 3 2 7 13 9 0 10 2 3 1 10 9 2 3 13 9 13 1 10 9 1 13 14 15 16 1 10 9 2
48 9 9 16 13 1 10 9 10 0 1 9 10 9 2 13 16 9 10 9 13 1 9 9 0 1 10 9 13 1 10 9 13 14 10 9 1 11 2 1 16 11 11 2 13 1 9 2 2
56 2 10 9 13 13 1 11 9 0 2 16 3 2 4 13 1 15 2 16 15 0 2 2 13 3 9 10 9 2 11 11 2 1 9 15 1 11 1 9 9 9 1 11 2 11 2 11 2 11 2 11 2 11 7 11 2
26 1 9 15 2 13 14 9 9 10 9 15 1 9 1 9 1 11 2 7 10 9 10 0 3 13 2
21 1 9 9 15 13 11 3 1 9 10 9 14 11 2 1 9 16 13 1 11 2
48 11 13 3 16 10 9 16 13 14 9 10 9 10 9 2 0 1 10 9 13 0 2 7 16 9 10 9 10 0 13 1 10 9 10 9 13 1 13 1 10 9 10 0 13 14 9 15 2
10 11 13 3 1 9 11 2 11 11 2
17 12 10 9 13 16 10 9 1 11 0 7 0 7 7 13 3 2
32 10 12 1 15 3 13 14 10 9 10 0 1 13 14 11 13 1 11 2 7 11 13 16 13 3 1 9 14 9 11 0 2
27 9 15 14 11 1 11 13 10 0 3 2 16 16 9 0 13 16 3 15 0 7 9 0 13 1 9 2
12 11 13 9 15 10 0 14 11 1 9 15 2
35 1 9 15 1 11 13 11 1 9 10 9 2 11 11 2 16 9 10 9 14 10 11 13 3 13 9 1 9 1 13 14 11 1 11 2
32 9 10 9 2 11 11 2 4 16 10 9 16 3 13 1 2 9 10 9 4 9 1 11 2 7 13 13 9 0 1 15 2
18 11 13 1 11 16 11 7 11 3 13 9 1 9 9 1 10 15 2
31 9 0 13 2 1 9 9 0 1 9 14 9 10 9 2 16 11 13 1 9 15 14 10 9 13 0 1 9 1 11 2
32 9 1 11 13 16 1 10 9 10 0 13 10 9 13 14 10 9 1 11 11 1 10 9 10 0 7 1 10 9 10 0 2
64 1 10 9 10 0 2 13 10 9 1 10 9 10 9 1 10 9 10 3 2 0 2 13 9 0 7 13 9 0 1 10 11 2 1 13 1 9 10 9 16 13 9 1 9 1 11 2 1 9 10 9 2 16 11 13 3 1 9 9 15 1 10 11 2
33 1 10 9 10 0 2 13 9 0 0 1 9 2 10 9 2 9 2 1 13 1 9 9 14 12 9 1 9 10 9 10 0 2
36 1 9 10 9 10 0 2 13 9 15 10 0 14 10 9 10 9 2 0 1 9 10 9 10 0 7 13 3 9 15 10 0 7 10 0 2
53 1 9 9 13 11 2 16 10 9 13 2 1 10 9 2 12 13 9 2 9 9 2 3 1 12 9 7 9 7 12 9 1 9 9 2 12 2 11 2 12 2 16 13 1 9 10 9 10 0 10 0 3 2
13 10 9 13 3 12 9 9 16 13 3 1 11 2
39 9 10 9 13 1 9 10 9 10 0 7 13 15 10 9 10 0 10 0 10 0 3 1 9 0 1 3 11 2 9 11 1 11 13 1 12 1 12 2
31 9 0 1 10 9 1 12 10 9 13 9 0 1 15 16 11 3 13 1 15 1 13 1 9 9 10 9 1 10 9 2
33 1 10 9 13 3 9 9 10 9 11 11 2 9 9 15 14 11 2 16 15 10 9 10 0 3 1 9 10 9 14 10 9 2
36 1 10 9 10 0 13 13 1 11 9 0 14 0 2 16 13 1 9 1 10 9 2 1 10 9 3 2 0 0 16 13 13 1 9 0 2
75 9 9 2 9 16 13 1 9 16 13 1 9 16 13 1 10 9 1 9 10 9 10 0 2 1 9 10 9 1 9 10 9 10 0 2 2 13 16 12 9 1 10 13 10 0 13 1 9 10 9 10 0 1 10 9 7 3 12 9 14 9 10 9 13 16 15 13 1 9 10 9 10 0 3 2
33 9 10 9 14 11 7 14 11 2 9 11 11 11 2 9 7 11 11 2 11 2 13 3 1 10 9 11 1 9 10 9 11 2
41 15 13 1 10 9 3 13 1 9 0 0 1 11 7 3 13 1 9 9 16 13 11 13 1 9 10 9 14 10 11 2 16 1 15 13 3 9 0 1 11 2
14 11 13 12 12 9 0 1 11 1 10 9 10 0 2
14 1 9 13 1 11 12 9 0 7 12 12 9 0 2
28 9 0 0 13 1 9 11 2 16 11 3 13 9 9 1 9 10 9 14 10 11 1 9 1 9 1 11 2
18 11 13 3 16 3 13 13 1 9 11 16 13 9 1 9 1 11 2
10 9 10 9 11 11 13 3 1 11 2
19 15 10 9 10 0 14 9 14 9 16 13 1 9 0 1 9 10 9 2
15 11 13 16 10 9 11 1 9 0 13 13 1 9 13 2
25 1 9 9 15 1 9 15 10 0 13 11 16 1 11 7 1 11 9 0 1 9 1 10 9 2
32 1 9 9 1 11 13 9 11 2 11 11 2 16 13 3 16 13 16 4 13 13 9 1 10 9 10 3 2 0 1 11 2
26 15 13 16 4 13 14 10 10 9 10 0 7 10 0 1 13 14 10 9 1 10 9 1 9 9 2
29 9 1 9 15 14 10 9 10 9 2 0 2 11 11 2 1 9 1 11 2 13 3 9 9 1 9 10 9 2
19 11 13 1 15 1 11 12 9 2 9 1 11 2 1 15 1 12 9 2
24 10 9 10 0 1 11 13 1 11 1 10 9 2 1 16 1 10 9 10 0 13 1 15 2
39 10 9 1 9 10 9 11 1 10 9 13 1 9 10 9 16 13 1 11 2 7 9 15 14 9 9 2 10 9 13 1 9 9 15 16 13 1 11 2
29 10 9 10 0 1 11 2 11 11 11 2 11 2 13 1 9 11 16 9 0 1 9 11 13 14 10 10 9 2
20 10 9 13 14 9 15 10 9 1 9 10 9 11 1 9 9 1 10 9 2
55 1 9 1 9 0 0 13 11 2 2 15 13 14 10 9 14 15 1 3 9 7 10 9 13 14 10 9 14 10 10 9 7 10 10 9 2 1 16 15 13 13 9 9 1 11 1 9 0 0 2 1 9 0 2 2
14 1 9 10 9 13 1 9 10 9 1 9 10 9 2
31 9 10 9 13 1 10 9 9 14 1 12 9 14 9 1 10 9 2 16 3 13 13 1 11 3 1 10 9 10 0 2
6 15 13 9 9 0 2
20 9 1 9 10 9 13 16 10 9 13 13 9 15 14 9 9 0 1 11 2
23 3 1 11 13 1 9 10 9 2 13 9 0 0 7 13 9 15 1 11 14 9 0 2
28 9 0 13 1 12 9 9 7 1 12 9 1 9 1 9 1 9 9 2 16 13 1 9 10 9 1 11 2
23 9 0 13 16 3 13 9 1 9 9 10 9 1 9 1 9 9 2 3 1 9 0 2
38 1 9 10 13 11 13 9 9 12 2 11 11 2 11 2 1 9 10 9 11 2 16 13 1 9 1 2 9 9 9 2 1 16 13 1 9 9 2
34 3 13 9 2 9 1 10 9 14 11 11 2 9 12 2 1 9 10 9 11 2 1 11 13 1 10 9 11 11 11 2 9 12 2
21 9 9 1 11 13 1 11 9 2 11 2 9 12 2 1 9 10 9 10 0 2
4 15 13 3 2
23 1 9 11 13 1 9 11 11 11 2 9 12 2 15 13 3 7 13 1 9 10 13 2
14 1 11 13 12 9 1 9 1 9 9 1 9 9 2
22 9 9 9 11 2 9 2 9 11 11 2 13 16 10 9 13 14 10 10 9 15 2
13 1 9 15 2 13 2 13 1 9 1 9 0 2
25 7 7 9 0 13 16 10 10 9 13 1 9 9 9 2 1 16 1 9 1 10 0 9 0 2
11 8 8 8 8 13 1 9 11 9 0 2
14 9 0 13 1 12 9 16 13 1 9 1 10 9 2
8 9 11 13 16 3 13 9 2
13 3 13 10 9 1 10 9 10 9 1 10 9 2
13 9 0 13 16 7 13 9 2 13 10 9 3 2
15 8 8 8 10 9 13 1 9 0 14 9 1 10 9 2
17 1 9 11 13 9 0 1 9 10 9 10 12 1 9 10 9 2
12 10 9 10 9 10 0 13 13 1 9 0 2
34 9 0 13 16 1 9 1 9 10 9 1 10 9 13 9 11 2 9 12 2 9 9 10 9 9 9 11 2 1 9 1 9 15 2
43 1 10 11 14 11 13 3 9 14 9 10 9 10 0 1 9 11 1 9 9 1 9 9 2 10 9 10 0 2 1 11 7 1 9 15 14 9 10 9 2 11 11 2
28 1 10 9 13 9 1 9 10 9 2 7 9 11 13 9 9 1 9 0 16 1 10 9 1 13 13 9 2
11 13 1 9 9 16 13 9 15 14 9 2
42 1 9 10 9 13 11 9 1 10 9 11 2 11 1 9 11 2 1 16 9 9 13 13 14 13 10 9 2 9 11 2 9 12 2 16 13 1 9 9 1 11 2
5 10 13 3 13 2
34 7 12 9 2 7 13 14 9 10 9 2 1 13 14 10 9 10 0 1 9 10 9 1 9 12 2 16 13 1 10 9 1 9 2
29 1 9 0 1 11 13 10 9 1 9 9 10 9 1 10 9 2 3 9 10 9 2 1 9 9 9 10 9 2
35 3 13 10 9 16 3 13 4 13 1 9 9 0 1 10 9 16 13 1 9 10 9 2 16 16 13 10 9 10 0 14 9 10 9 2
33 1 10 9 1 10 9 1 9 10 9 13 3 11 11 2 9 15 10 0 14 9 10 9 2 1 10 9 1 9 9 10 9 2
30 1 9 11 13 3 9 9 11 11 11 16 3 13 9 1 9 9 10 9 1 10 9 2 1 13 14 9 10 9 2
39 4 13 16 1 1 9 2 16 13 10 9 1 10 9 10 0 1 9 10 9 7 9 11 2 13 9 9 0 1 12 10 9 1 9 10 9 10 0 2
41 1 9 11 13 16 4 13 9 10 3 0 1 9 15 14 9 0 2 16 13 9 0 1 10 9 2 7 7 1 10 9 13 1 9 10 9 1 1 9 0 2
25 1 10 9 13 13 1 9 0 1 9 9 10 9 1 9 0 2 7 10 9 0 3 3 13 2
31 9 1 10 9 13 16 13 10 9 1 9 15 13 14 9 9 10 9 2 7 13 16 9 15 4 13 1 9 10 9 2
18 8 8 1 11 13 10 9 1 10 9 1 9 12 1 9 9 0 2
29 7 2 7 10 9 3 13 13 14 9 10 9 16 13 1 10 9 2 15 13 13 1 9 10 9 1 9 0 2
19 15 1 10 3 2 9 1 9 15 14 10 9 13 14 10 9 10 0 2
38 1 15 0 3 2 9 1 9 10 9 10 0 2 16 16 3 13 3 10 9 13 1 10 9 10 0 2 7 10 9 13 1 12 12 1 12 12 2
9 9 12 13 1 3 12 12 9 2
49 9 9 10 9 3 3 13 2 16 9 10 9 13 1 9 10 9 16 15 13 12 12 9 1 9 15 1 10 9 10 0 2 1 9 9 9 10 9 7 9 0 1 9 9 10 9 3 9 2
35 3 1 10 9 10 0 1 10 11 13 3 9 0 1 9 10 9 13 1 9 10 9 10 0 7 13 1 10 9 10 9 13 9 9 2
15 10 9 13 1 9 1 9 10 9 10 0 1 9 7 2
45 1 9 9 13 9 10 9 1 9 0 1 10 9 1 10 9 10 0 7 13 1 9 0 3 1 10 9 1 10 9 10 0 2 16 9 15 13 3 1 9 10 9 10 0 2
19 10 9 13 13 1 9 1 9 10 9 11 13 14 9 10 9 1 11 2
33 9 13 16 10 9 10 0 13 1 9 14 9 0 7 10 9 10 0 13 1 15 16 9 15 13 7 13 1 10 9 10 0 2
30 10 9 1 9 10 9 11 13 1 9 10 9 1 11 13 1 9 9 1 9 9 9 10 9 10 0 1 9 11 2
34 1 9 9 15 2 16 13 1 9 7 2 13 9 10 9 10 0 1 12 9 3 1 1 9 14 12 9 16 13 1 9 10 9 2
51 3 1 15 2 10 9 13 16 1 9 10 9 1 9 10 9 7 10 9 2 13 9 15 1 9 0 1 10 9 1 9 11 7 13 16 13 1 15 1 13 1 10 9 10 0 1 10 9 1 11 2
27 8 8 8 13 7 13 1 9 7 1 10 9 1 10 9 7 10 9 10 0 1 9 10 9 1 11 2
43 10 9 13 16 9 10 9 14 9 12 10 9 10 13 10 13 13 1 9 13 1 9 10 9 1 9 10 9 13 1 9 15 10 0 14 10 11 1 10 9 10 0 2
20 10 11 13 7 13 1 9 14 12 9 1 9 14 12 9 1 9 10 9 2
23 9 9 15 14 10 9 10 0 14 11 13 14 9 10 9 1 9 9 9 2 3 13 2
44 9 9 11 11 9 9 9 1 10 9 10 0 1 11 7 11 13 1 9 15 9 1 9 10 9 2 7 1 15 13 1 9 10 9 1 9 9 1 9 9 1 10 9 2
18 14 10 9 1 9 10 9 13 9 10 9 1 10 9 2 11 11 2
29 11 13 16 10 9 9 13 4 13 13 12 9 9 1 10 9 2 10 9 1 10 9 7 10 9 1 9 11 2
14 9 10 9 10 0 3 13 9 9 1 9 9 15 2
38 1 9 15 2 10 9 1 9 10 9 1 10 9 1 9 10 9 10 0 13 3 13 1 9 2 7 9 9 10 9 10 0 3 13 14 10 9 2
33 9 10 9 13 3 12 1 9 10 9 1 9 14 9 9 1 10 9 2 1 9 16 13 1 0 2 1 9 10 9 10 0 2
28 10 9 13 13 3 14 9 10 9 16 13 1 9 10 9 1 10 9 1 10 9 10 0 1 9 10 9 2
46 9 13 10 0 13 1 9 1 12 1 9 10 9 10 0 2 1 9 0 1 9 10 9 2 13 1 9 9 9 9 1 9 13 2 11 2 1 11 2 1 15 14 9 11 11 2
13 11 13 1 9 1 9 9 2 1 9 10 9 2
59 1 15 13 3 9 7 9 10 9 10 0 14 10 9 2 9 11 11 2 1 9 1 9 15 14 9 9 11 2 11 11 2 16 9 9 11 13 9 1 10 9 2 7 16 9 15 14 9 9 9 1 2 11 2 13 1 9 15 2
17 11 13 1 9 9 13 14 9 10 9 1 9 14 9 7 9 2
33 1 9 11 13 9 1 9 13 10 0 16 13 1 15 3 9 9 14 12 12 9 2 7 1 9 13 1 15 13 1 9 0 2
27 1 9 3 13 11 16 1 9 15 13 13 1 9 0 1 2 9 11 2 2 7 13 14 9 10 9 2
19 1 9 7 9 1 10 9 15 13 9 9 16 4 13 1 9 1 12 2
30 9 9 13 1 9 11 16 13 4 13 9 0 1 0 2 7 16 10 9 13 1 10 9 10 0 1 9 10 13 2
26 1 9 10 9 2 13 9 11 1 15 9 13 1 9 10 13 11 1 9 1 10 9 10 0 11 2
16 9 11 13 16 10 9 13 1 9 1 9 10 9 14 15 2
39 1 9 9 9 10 9 14 10 9 2 9 11 11 2 2 1 10 10 9 1 9 15 14 11 2 13 13 9 16 9 1 12 10 9 13 9 9 2 2
30 11 7 13 9 15 1 9 9 10 9 2 7 13 16 2 10 13 1 9 0 14 9 9 7 9 1 9 0 2 2
32 9 9 13 1 11 7 10 9 11 11 13 16 9 13 10 0 13 14 9 11 16 16 13 9 0 7 1 9 0 1 15 2
30 1 9 15 13 3 9 11 1 9 9 16 13 1 9 9 2 1 9 9 9 1 9 10 13 10 0 11 1 11 2
46 1 15 1 9 2 13 10 9 2 15 3 13 13 1 9 9 0 1 10 9 1 9 0 1 11 1 9 10 13 11 2 1 7 16 13 1 10 9 3 12 9 1 9 13 0 2
27 9 11 13 16 9 9 13 4 13 14 9 11 9 1 10 9 7 13 13 1 10 9 10 0 10 0 2
42 9 11 13 13 1 9 10 9 2 7 1 9 16 13 3 1 2 11 2 15 13 2 2 10 9 15 13 16 13 1 15 1 9 14 12 9 13 3 1 9 11 2
13 13 16 15 13 1 10 9 10 0 7 9 9 2
22 13 16 10 9 10 0 14 10 9 1 9 10 13 11 13 1 9 15 7 7 13 2
24 13 3 16 10 9 0 13 1 9 7 1 9 16 13 1 15 9 8 8 8 10 13 11 2
14 10 9 16 13 13 0 1 9 7 0 1 10 13 2
6 7 10 9 3 13 2
23 13 1 15 9 14 9 3 13 3 1 15 2 7 15 13 3 13 1 15 3 9 2 2
45 9 0 1 9 7 9 1 9 0 14 12 12 9 2 16 13 1 9 0 7 0 2 13 1 9 10 9 14 10 9 10 3 2 0 1 9 11 2 11 16 13 3 1 11 2
16 10 9 13 1 9 9 2 9 2 9 2 9 7 9 9 2
26 14 11 13 1 10 9 9 9 10 9 7 10 9 7 10 9 10 0 14 9 10 9 7 10 9 2
18 14 11 13 9 9 10 9 2 10 9 2 7 9 10 9 10 0 2
28 11 11 2 9 9 10 9 2 13 16 9 15 13 9 1 9 1 15 13 9 9 0 0 2 1 9 0 2
25 1 9 12 2 13 10 9 10 13 1 9 1 9 10 9 1 10 9 10 0 1 1 12 9 2
15 10 9 10 3 2 0 1 9 7 9 13 1 9 12 2
36 1 9 15 2 13 11 7 11 10 12 12 12 9 1 10 9 2 14 10 9 1 10 9 13 1 9 9 0 1 9 10 9 7 10 9 2
14 1 9 10 9 2 13 9 10 9 1 12 12 9 2
24 9 12 2 1 1 12 9 2 13 11 2 11 2 11 7 12 9 1 10 9 14 9 11 2
102 11 11 2 9 9 9 9 14 12 9 1 11 2 13 3 1 9 15 14 9 1 9 2 13 0 1 9 10 9 2 9 15 11 2 9 9 0 2 13 1 11 1 9 2 9 1 9 9 1 11 2 7 3 15 13 9 13 3 1 10 9 10 3 0 14 15 2 9 15 11 9 10 12 13 3 1 11 2 7 1 9 10 9 13 3 9 9 2 2 1 16 3 13 1 9 1 10 9 10 0 2 2
14 9 9 11 13 13 1 9 14 9 10 9 10 0 2
33 1 11 15 13 1 12 1 11 2 7 1 9 10 9 3 13 1 9 9 15 14 9 15 14 11 1 9 10 9 1 9 9 2
8 9 3 3 13 1 10 9 2
27 1 15 13 1 12 1 1 12 10 9 16 13 14 9 10 9 10 0 1 11 1 9 10 9 10 0 2
23 9 0 1 10 9 2 16 15 9 0 1 10 9 2 16 13 3 13 1 9 10 9 2
47 1 9 16 13 3 1 3 1 9 11 2 11 1 9 2 10 13 10 9 0 1 10 12 10 12 2 2 13 10 9 1 9 11 11 14 9 15 14 10 9 1 9 15 14 10 9 2
23 2 3 16 13 1 10 9 14 10 9 1 10 9 13 10 9 10 0 16 13 1 15 2
21 3 3 4 10 9 13 1 9 10 9 9 0 7 0 2 1 3 9 0 2 2
15 9 11 13 10 0 16 13 1 9 10 9 1 10 9 2
33 10 10 9 1 10 9 2 9 10 9 10 0 2 3 13 3 14 10 9 1 9 0 1 9 9 15 7 9 15 14 10 9 2
38 1 9 0 13 10 9 10 0 1 12 9 15 10 9 2 10 9 10 0 7 10 9 10 0 1 10 9 10 0 14 2 9 0 1 10 9 2 2
30 10 13 1 9 9 2 0 2 16 1 9 15 13 10 9 1 9 2 13 1 9 7 13 1 15 14 10 10 9 2
32 10 9 10 0 2 12 9 1 9 1 9 9 12 9 2 13 1 9 10 9 14 10 9 7 13 1 15 9 1 10 9 2
13 10 9 4 13 1 10 9 9 9 12 1 9 2
18 10 9 9 0 2 1 9 14 12 9 1 9 2 13 1 10 9 2
20 9 1 9 13 1 10 9 9 0 14 9 2 16 13 1 9 7 1 0 2
9 7 9 9 0 15 13 9 0 2
27 9 10 9 14 10 9 2 16 13 1 9 0 7 0 0 2 13 3 9 12 16 13 14 9 10 9 2
20 9 15 10 0 14 9 10 9 1 10 9 10 2 0 2 3 13 7 15 2
25 7 16 10 9 7 1 15 9 10 9 13 14 14 15 7 13 9 3 1 2 9 10 9 2 2
22 10 9 10 0 13 2 7 12 9 13 3 14 9 15 10 0 1 10 9 10 0 2
25 9 13 13 3 10 1 15 7 3 13 1 10 9 1 1 10 9 10 0 16 13 1 10 9 2
16 10 9 10 15 16 1 10 9 1 11 1 10 9 13 0 2
12 10 9 13 1 15 9 9 0 1 10 9 2
57 9 0 9 9 0 7 3 2 0 0 13 14 10 9 16 13 1 10 9 1 10 9 1 9 1 2 9 0 1 10 9 2 1 2 9 9 1 9 9 2 16 13 9 1 10 9 10 9 2 2 7 16 10 9 0 3 2
28 13 3 16 13 16 10 9 1 11 13 10 9 16 13 1 10 9 2 11 2 2 9 2 9 2 9 2 2
18 9 15 1 10 9 0 7 0 9 0 2 16 13 14 9 10 9 2
31 11 9 2 9 9 9 7 12 10 9 14 9 2 9 0 1 10 9 2 2 13 2 2 10 9 13 16 9 15 9 2
12 13 1 15 3 12 9 13 16 15 3 3 2
12 3 1 9 0 15 13 16 15 3 9 2 2
13 9 2 1 9 9 2 13 3 9 13 1 9 2
15 3 1 3 13 9 9 9 1 11 1 9 1 10 9 2
15 3 1 11 13 14 15 2 3 13 14 10 9 11 2 2
24 7 3 13 9 0 1 9 11 14 10 9 1 9 2 9 16 13 1 9 2 9 7 9 2
17 14 11 11 2 9 0 1 11 2 13 1 9 15 1 9 11 2
27 1 12 9 13 1 11 11 10 9 7 9 15 10 9 7 13 13 1 9 2 9 2 3 1 9 0 2
9 1 10 9 10 0 3 13 9 2
14 1 10 9 7 1 10 9 10 0 10 9 13 13 2
13 1 9 15 13 1 9 10 9 7 13 9 9 2
5 10 9 13 9 2
23 2 3 13 9 1 10 9 2 2 13 11 2 12 2 2 2 7 10 9 13 0 3 2
6 13 16 15 1 9 2
12 3 9 0 1 10 9 2 0 2 3 0 2
4 13 7 13 2
7 3 13 14 15 10 9 2
16 10 3 16 13 1 10 9 1 11 7 3 13 2 0 3 2
6 3 13 16 15 9 2
12 3 15 13 16 15 0 2 7 15 0 2 2
23 1 7 10 9 10 0 10 15 2 3 13 1 9 15 16 1 9 15 13 1 10 9 2
9 15 9 9 0 7 13 13 3 2
33 11 11 2 10 9 14 9 11 2 13 1 9 2 2 7 13 9 10 9 11 13 1 10 9 2 13 13 9 1 16 3 13 2
14 10 9 13 1 15 7 9 10 9 13 1 15 2 2
28 3 9 9 11 2 16 13 1 1 9 1 10 9 11 16 1 9 11 2 13 16 10 9 13 9 1 15 2
45 10 9 2 11 2 9 9 0 9 2 10 9 2 11 2 13 9 2 10 9 2 11 2 12 2 2 13 13 9 9 1 10 9 2 7 7 13 9 0 1 10 9 10 0 2
30 13 1 9 9 15 13 1 10 9 10 0 2 11 2 9 0 2 16 13 1 9 0 3 14 10 9 1 10 9 2
24 13 16 9 13 9 16 0 13 1 15 2 16 1 9 13 9 0 2 13 3 2 13 9 2
20 1 9 7 9 1 11 9 9 11 3 13 16 10 9 3 13 1 10 9 2
15 3 10 9 13 9 2 7 15 3 1 15 2 15 13 2
27 2 10 9 1 9 13 16 13 9 2 2 13 11 2 1 15 4 13 3 14 10 9 2 1 10 9 2
20 15 13 16 10 9 16 3 13 9 1 10 9 1 11 2 13 13 1 9 2
19 14 13 1 15 10 9 2 7 3 13 9 2 15 13 1 10 9 2 2
26 10 9 11 13 2 2 1 10 9 3 13 10 13 9 2 10 13 9 2 3 13 9 1 10 9 2
10 3 15 0 2 7 15 3 10 9 2
15 15 13 16 10 9 16 13 1 10 9 3 13 13 3 2
14 15 13 14 10 9 7 15 13 9 0 1 10 9 2
5 3 15 3 2 2
29 11 11 2 9 10 9 2 13 9 1 10 9 14 9 10 9 2 2 15 0 3 7 13 1 15 1 9 2 2
18 0 1 10 9 10 0 13 13 1 9 15 13 1 15 9 1 9 2
37 9 13 1 15 14 9 10 9 1 10 9 10 0 2 14 9 10 9 10 0 16 13 1 15 2 1 1 9 2 7 1 1 9 7 13 9 2
23 13 9 11 2 11 11 2 13 3 16 4 13 9 0 14 9 1 9 15 14 10 9 2
16 3 4 16 9 13 1 10 9 16 16 15 13 1 9 11 2
23 3 4 16 15 13 1 10 9 7 13 1 10 9 14 15 2 1 16 13 2 15 13 2
15 7 13 9 16 4 13 9 0 1 10 9 1 9 2 2
8 1 9 10 9 13 10 9 2
15 10 9 13 9 7 13 1 11 9 1 10 9 10 0 2
20 3 10 9 13 1 10 9 3 1 3 16 15 13 1 10 9 9 0 0 2
25 9 0 14 10 9 1 9 13 16 12 9 12 9 1 10 9 4 13 9 14 9 1 10 9 2
19 1 2 7 9 15 3 10 9 13 3 1 13 14 9 15 14 10 9 2
27 4 13 16 15 13 1 10 9 1 9 7 1 9 2 1 9 15 14 12 9 9 2 1 15 9 9 2
13 11 11 13 16 10 9 13 13 1 9 9 15 2
28 15 13 15 1 9 9 2 7 1 15 16 9 10 9 13 1 10 9 1 9 9 7 1 9 1 9 9 2
26 2 10 9 13 16 3 13 1 10 9 16 13 7 13 2 7 1 10 9 15 3 13 14 15 2 2
14 11 13 3 3 1 10 9 10 0 14 9 10 9 2
13 2 3 16 13 3 13 1 3 2 2 15 13 2
6 2 10 9 13 13 2
13 1 9 15 4 13 1 9 13 9 0 1 9 2
21 3 10 9 13 3 13 1 15 3 9 0 2 7 4 1 15 13 1 9 15 2
20 10 9 10 0 13 13 1 10 9 14 10 9 13 4 1 9 1 9 15 2
12 1 15 4 16 15 13 3 10 15 13 2 2
27 2 13 9 0 1 15 1 10 9 0 2 2 13 11 9 2 9 1 9 9 11 1 10 9 10 0 2
14 2 1 9 15 14 9 2 15 13 14 15 3 2 2
17 9 15 15 13 14 9 10 9 16 13 14 10 9 1 10 9 2
17 0 9 16 9 10 9 13 1 10 9 2 3 3 1 10 13 2
34 7 2 7 2 13 13 1 9 10 9 2 16 13 13 10 9 7 9 1 10 9 1 9 9 2 1 9 1 9 9 1 10 9 2
32 9 15 14 9 10 9 10 0 2 11 11 2 13 9 1 9 16 13 1 15 9 2 15 9 9 2 13 9 1 9 0 2
26 3 2 1 9 1 9 9 2 1 9 9 1 9 10 9 2 13 10 9 10 0 1 9 10 9 2
38 1 9 1 9 15 2 4 13 1 9 14 9 10 9 14 9 11 2 2 7 1 11 1 11 13 10 9 16 13 1 15 9 2 15 9 13 2 2
7 11 2 9 2 11 2 2
6 11 11 13 13 9 2
7 11 1 9 7 1 9 2
43 9 1 3 13 9 10 11 9 16 3 13 3 13 15 2 9 12 9 1 10 9 10 0 1 11 11 2 16 13 9 1 10 9 16 13 2 11 11 11 12 12 2 2
25 11 13 1 10 9 12 12 7 13 9 0 14 11 11 1 9 9 2 1 9 2 1 2 12 2
14 3 1 10 9 10 12 13 10 11 9 2 12 9 2
15 1 9 11 2 11 11 2 13 15 10 9 10 2 12 2
27 12 9 13 3 1 2 12 9 1 11 2 16 10 9 10 0 14 10 9 13 11 11 11 2 12 9 2
16 1 11 2 11 12 2 11 11 11 1 9 15 10 0 12 2
14 11 11 2 12 9 2 13 9 12 9 1 10 9 2
14 15 13 10 9 10 0 1 10 9 16 11 11 13 2
14 11 11 13 12 9 1 10 9 7 11 12 1 11 2
42 11 11 13 1 11 12 12 2 11 1 11 11 14 10 11 12 12 2 11 13 14 10 11 1 11 11 12 12 7 11 11 1 11 2 9 11 2 14 11 12 12 2
18 9 0 2 11 11 12 12 2 11 11 12 12 2 11 11 12 12 2
31 9 2 9 13 9 1 9 9 7 1 9 0 2 1 12 9 1 9 11 3 2 1 9 9 10 9 13 3 9 0 2
44 10 9 13 1 9 9 2 1 9 7 1 9 0 1 13 3 1 2 12 9 2 13 1 15 13 9 2 16 13 1 11 1 10 9 11 2 13 9 10 9 2 11 11 2
12 1 9 11 1 10 9 13 12 9 9 0 2
21 15 13 9 9 1 9 0 1 16 13 9 1 9 2 1 9 9 9 1 11 2
4 12 9 13 2
35 1 12 9 9 16 13 15 2 13 2 0 2 13 1 11 1 11 9 1 9 9 9 12 16 13 1 9 1 10 9 1 10 9 11 2
16 12 9 13 14 10 9 16 13 1 12 9 1 1 9 11 2
12 10 9 13 2 16 10 9 13 1 9 9 2
28 12 9 9 14 9 10 9 0 7 15 3 13 14 10 9 11 11 2 1 10 9 1 11 1 3 9 11 2
34 10 9 16 13 1 11 3 2 12 2 13 10 9 14 9 11 1 9 15 2 1 10 9 10 13 12 12 1 9 10 9 1 11 2
27 1 10 9 16 13 3 1 10 9 1 9 9 1 11 12 9 2 13 9 0 11 11 1 11 9 9 2
47 12 10 9 13 1 10 9 10 0 2 10 9 11 11 2 11 11 2 16 13 1 9 9 0 2 10 9 10 0 11 11 1 10 9 9 11 7 10 9 11 11 11 1 10 9 11 2
6 2 10 9 13 0 2
33 15 13 13 3 1 10 9 16 13 2 7 13 1 9 10 9 7 10 12 1 10 12 3 13 14 10 9 2 2 13 11 11 2
19 3 3 13 3 9 12 1 10 9 10 13 1 10 9 16 13 1 11 2
17 10 9 11 13 1 9 0 1 10 0 16 13 13 3 1 11 2
41 2 15 3 3 0 1 9 10 9 2 7 13 1 15 9 0 7 15 13 13 2 16 10 9 0 13 14 15 1 10 9 2 1 10 9 1 9 10 9 2 2
23 15 13 14 15 12 12 1 10 9 16 13 1 10 9 2 7 10 9 14 15 13 9 2
13 13 3 13 1 10 9 14 15 2 2 13 11 2
6 9 11 2 9 2 2
25 1 9 0 16 13 1 11 7 1 10 9 10 0 13 1 9 15 12 9 0 1 9 1 11 2
45 9 15 10 0 7 9 15 10 0 13 1 10 9 10 0 16 13 1 15 1 10 9 10 0 1 10 9 10 0 2 7 3 1 10 9 16 15 3 0 3 1 9 9 0 2
22 1 15 2 7 4 13 13 9 1 9 3 2 13 10 9 15 3 3 1 11 9 2
24 13 1 15 13 13 1 9 11 1 9 10 9 7 13 1 9 15 1 9 10 9 14 15 2
14 2 15 13 16 13 10 9 10 0 16 13 1 11 2
35 15 9 15 4 13 7 13 1 11 7 1 9 15 2 2 13 9 11 11 11 2 11 2 9 10 9 10 0 16 13 1 9 10 9 2
32 1 9 10 9 10 0 13 1 10 9 12 9 1 9 9 2 7 13 1 9 9 1 2 2 11 2 11 2 10 9 2 2
10 9 13 9 0 1 9 9 10 9 2
13 2 13 10 9 13 1 9 15 7 13 1 11 2
15 13 10 9 13 1 10 9 2 2 13 1 12 10 9 2
24 10 9 10 0 14 10 9 3 13 12 9 2 7 3 3 12 1 15 13 9 1 10 9 2
26 9 11 2 11 13 16 15 13 13 1 9 0 7 1 9 3 3 7 13 16 13 3 9 1 9 2
25 1 11 13 9 16 9 10 9 13 13 9 1 10 9 1 9 16 15 13 14 10 9 1 15 2
14 3 3 13 3 13 10 9 1 9 10 9 7 13 2
25 1 10 9 13 16 15 13 9 1 10 9 10 0 10 0 16 13 1 11 7 10 13 12 9 2
27 9 9 11 13 1 10 9 10 0 3 16 13 1 3 12 9 1 9 9 7 9 1 9 9 13 9 2
17 10 9 10 0 1 15 13 9 13 11 2 16 1 10 9 9 2
23 3 13 12 9 1 13 1 10 12 16 3 13 8 1 9 9 10 9 1 9 9 11 2
15 1 9 0 2 10 9 11 16 1 11 2 13 12 9 2
24 3 13 9 1 11 2 9 2 11 2 9 2 11 2 11 2 11 2 11 7 9 2 11 2
18 10 9 13 3 9 1 12 9 1 9 2 9 15 1 9 10 9 2
34 9 10 9 2 11 11 2 13 16 10 9 10 0 13 1 9 2 11 2 9 2 9 2 11 2 1 11 2 11 7 9 2 12 2
30 1 13 9 13 14 15 10 9 1 9 9 9 9 1 10 9 10 9 2 7 1 9 16 15 3 13 1 12 9 2
15 3 13 9 9 11 12 9 1 9 0 1 9 2 11 2
13 9 10 9 1 9 7 9 2 1 9 12 9 2
20 10 9 13 1 9 9 12 12 12 9 2 7 1 9 10 9 12 12 9 2
25 1 11 13 10 9 1 3 12 1 9 10 9 1 9 1 9 9 1 9 10 9 14 10 9 2
24 15 13 12 9 1 9 16 1 12 9 1 9 2 7 13 1 12 1 12 12 9 1 9 2
22 1 11 13 10 9 9 14 12 9 2 1 9 12 9 2 1 9 9 1 10 9 2
29 9 11 9 2 16 9 15 13 1 10 9 10 9 2 0 2 13 1 10 9 7 13 1 10 9 12 12 9 2
23 11 2 16 1 9 15 13 10 9 11 11 2 13 1 11 1 9 0 2 3 1 9 2
24 1 10 9 10 0 13 9 13 9 7 9 16 13 1 9 9 0 1 9 0 2 0 3 2
35 1 10 9 13 9 13 7 13 9 9 0 2 7 3 16 3 13 1 3 10 9 14 9 1 9 0 2 16 13 3 3 1 9 0 2
28 9 1 9 10 9 13 2 1 9 11 9 2 9 1 9 12 9 1 9 10 9 14 11 1 9 2 11 2
24 10 9 13 13 1 9 10 9 12 9 1 9 9 0 3 2 16 16 10 9 13 9 0 2
32 1 3 13 10 9 1 9 1 9 2 9 2 3 13 1 12 9 1 9 2 7 1 15 13 9 0 1 9 9 10 9 2
28 9 0 2 9 9 13 9 9 12 9 1 9 14 12 9 1 1 12 9 1 9 9 11 1 9 2 9 2
18 10 9 16 13 13 9 0 2 16 13 1 9 14 12 9 1 9 2
17 9 0 13 1 10 9 10 0 1 9 10 9 1 9 2 9 2
9 9 10 9 13 1 1 12 9 2
52 3 10 9 1 10 9 1 10 9 2 9 9 12 9 1 9 11 1 11 2 9 15 13 1 1 12 9 12 12 9 2 13 1 9 15 14 9 3 1 16 9 15 13 1 12 12 9 9 14 12 9 2
31 9 1 9 10 9 1 11 2 16 9 15 13 12 12 9 2 13 3 1 12 12 9 2 7 3 3 13 1 15 9 2
28 9 9 1 9 16 13 1 0 2 16 9 15 13 1 1 12 9 12 12 9 2 13 3 1 12 12 9 2
20 9 9 10 9 13 10 1 9 11 1 9 10 9 1 11 1 12 12 9 2
11 10 9 13 1 9 0 0 14 12 9 2
28 15 13 0 1 9 11 2 16 12 1 9 15 2 11 11 2 13 14 9 15 2 12 9 2 1 10 9 2
15 9 10 9 13 14 9 10 9 1 9 9 14 12 9 2
31 1 9 10 9 11 2 16 13 14 10 12 10 9 1 10 9 2 13 9 1 9 7 9 2 1 9 1 12 9 0 2
48 1 1 9 13 9 10 9 9 9 0 2 1 9 15 13 1 9 10 9 10 0 11 2 11 2 11 14 9 15 1 9 9 2 11 9 11 1 9 2 9 2 3 3 1 12 12 9 2
17 10 9 10 0 1 9 1 9 15 13 1 3 12 9 1 9 2
33 10 9 2 16 13 1 9 14 12 9 1 9 0 1 10 9 7 3 12 9 1 9 9 0 2 13 1 9 10 9 11 9 2
22 11 9 13 13 9 9 9 1 9 12 12 9 2 0 1 9 10 9 1 10 9 2
21 8 1 9 9 10 9 1 9 2 9 9 2 1 11 9 2 13 13 14 15 2
30 13 1 9 0 2 16 13 12 9 9 1 3 1 9 0 0 16 13 9 2 14 1 9 15 9 0 1 9 9 2
28 1 9 11 11 1 11 9 13 16 13 1 9 15 12 9 0 1 9 1 9 2 16 9 15 13 7 13 2
19 1 10 9 13 3 12 12 9 2 1 12 12 1 9 16 13 10 9 2
18 11 11 2 9 15 14 11 2 13 14 10 9 13 9 1 10 9 2
12 15 7 13 12 12 9 1 9 2 7 13 2
12 3 13 10 9 0 1 9 0 1 11 9 2
33 9 13 16 1 10 9 1 10 9 2 13 9 9 12 9 2 12 9 2 1 9 2 11 11 2 1 11 9 1 12 12 9 2
22 9 0 14 12 9 2 12 9 2 1 9 2 9 9 2 2 13 1 12 12 9 2
48 8 9 10 9 11 11 13 13 9 1 10 9 2 1 9 13 1 15 14 10 9 1 9 11 12 1 9 2 9 2 16 13 1 10 9 10 0 14 9 10 9 11 2 7 13 7 9 2
32 9 10 9 13 13 9 9 14 1 12 9 1 9 2 3 13 9 2 1 10 9 16 9 15 12 9 7 12 9 1 9 2
19 1 16 3 13 13 1 9 13 1 9 10 9 1 9 1 9 9 15 2
39 11 2 9 15 14 9 1 9 7 9 9 9 2 10 13 1 15 16 9 15 14 9 11 13 2 4 13 14 9 10 9 7 13 1 12 9 1 9 2
21 15 13 1 10 9 14 11 11 2 1 9 11 2 13 1 9 9 14 12 9 2
5 11 2 11 2 2
22 11 13 12 12 14 11 7 13 1 10 9 10 0 1 10 9 10 0 1 12 9 2
46 1 11 12 9 2 14 13 1 15 1 9 9 3 2 11 16 13 1 10 9 12 12 14 11 7 11 16 13 3 15 1 12 9 1 9 9 1 12 1 11 10 0 1 10 9 2
33 1 9 10 9 3 13 12 9 2 16 10 10 9 16 13 14 11 1 9 11 2 13 1 9 15 1 10 9 10 3 2 0 2
50 10 9 10 0 14 11 1 11 2 13 0 1 10 9 10 0 11 11 2 16 3 3 13 14 11 1 10 9 2 1 9 15 14 10 9 1 11 2 7 3 13 14 15 13 14 10 9 10 12 2
16 11 11 13 14 9 10 9 14 11 1 10 9 10 2 12 2
9 3 1 10 9 13 11 12 12 2
28 10 9 14 11 16 13 1 9 9 2 13 12 9 1 2 15 7 10 2 12 13 1 9 12 14 11 11 2
34 10 9 14 11 13 3 1 9 11 11 16 13 1 10 9 10 0 1 10 9 10 2 12 7 13 3 14 10 9 1 9 10 9 2
31 1 11 2 16 1 9 13 14 10 9 1 10 9 2 1 10 9 10 0 1 12 9 2 13 15 9 12 1 12 9 2
28 1 9 11 16 13 13 12 12 14 11 11 10 0 7 13 1 9 10 9 1 10 9 10 0 1 13 9 2
45 9 11 11 2 16 13 1 9 9 9 10 9 14 11 10 0 2 13 1 11 12 12 1 9 0 1 12 10 9 2 1 9 14 11 11 11 2 12 2 7 11 2 12 2 2
41 10 9 14 11 10 9 10 12 14 11 1 9 10 13 1 11 13 1 9 1 9 12 1 10 9 10 2 12 1 9 11 11 2 10 9 10 0 1 10 9 2
11 15 13 9 15 10 12 3 1 10 9 2
37 11 2 16 13 1 9 10 9 1 10 9 10 0 2 13 1 9 1 10 9 10 2 12 2 1 16 10 0 14 11 11 11 13 9 2 12 2
18 10 9 10 3 2 0 11 11 13 9 1 9 11 12 12 1 11 2
24 14 10 9 10 0 1 11 2 16 13 1 10 9 10 12 1 9 11 2 13 11 7 11 2
4 11 2 11 2
27 11 2 16 13 14 11 9 1 9 11 2 13 14 11 12 12 1 9 14 11 7 11 1 2 12 9 2
5 11 13 1 11 2
21 10 9 14 11 13 1 9 15 1 9 11 16 13 1 9 10 9 1 11 11 2
56 11 2 16 13 14 10 9 11 7 14 11 11 2 9 15 13 1 9 0 2 2 3 13 13 14 10 9 10 0 14 11 7 13 3 1 9 2 9 16 13 14 15 1 9 12 2 1 10 9 10 12 1 12 9 3 2
40 9 0 2 11 12 2 11 15 2 11 2 11 12 2 11 12 11 12 2 9 2 9 15 2 2 11 12 2 11 2 11 2 11 12 2 11 2 11 2 2
22 10 9 11 13 3 1 10 9 10 0 1 16 13 9 12 12 1 11 16 13 0 2
22 11 13 14 9 15 1 11 14 10 13 1 9 10 9 2 11 2 12 12 1 11 2
25 10 9 1 11 2 11 2 12 2 2 11 2 12 2 2 11 2 12 2 2 11 2 12 2 2
8 1 11 2 11 2 12 2 2
45 9 0 1 9 10 9 2 11 12 11 12 2 11 12 11 12 2 11 11 12 11 12 2 11 12 11 12 2 11 12 11 11 11 12 2 9 12 11 12 2 11 12 11 12 2
23 11 13 1 10 9 10 12 1 16 13 3 1 10 9 1 9 9 14 11 9 12 12 2
23 10 9 1 11 2 11 11 2 12 2 2 11 11 2 12 2 2 11 11 2 12 2 2
19 1 9 2 11 11 2 12 1 2 12 9 2 2 11 11 2 12 2 2
38 11 11 11 11 2 14 15 13 10 9 11 11 2 13 1 10 9 10 0 2 1 9 9 12 12 1 11 1 9 14 11 1 10 9 10 2 12 2
33 1 11 12 9 1 12 9 2 7 15 13 1 9 9 14 10 9 11 11 16 13 1 9 15 7 13 3 1 9 12 1 11 2
26 9 0 2 11 11 12 11 12 2 11 11 12 11 12 2 11 12 11 12 2 11 11 12 11 12 2
52 9 12 2 11 12 11 12 2 11 12 11 12 2 11 11 12 11 12 2 11 12 11 12 2 11 12 9 11 12 2 11 12 11 12 2 11 12 11 12 2 11 11 11 12 2 11 11 11 12 11 12 2
16 10 9 2 11 12 2 11 11 12 2 11 12 2 11 12 2
40 9 12 2 11 11 12 11 12 2 11 11 12 11 12 2 11 11 12 11 11 12 2 11 11 12 11 12 2 11 11 12 11 12 2 11 11 12 11 12 2
14 10 9 2 11 12 2 11 11 12 2 11 11 12 2
22 11 2 1 15 13 11 11 2 13 3 12 12 1 10 9 1 11 11 16 13 0 2
7 11 13 12 12 14 11 2
43 9 0 2 9 11 12 11 11 12 2 11 11 12 11 11 12 2 11 12 11 12 2 11 12 11 12 2 11 12 11 11 12 2 11 12 11 12 2 11 12 11 12 2
20 10 9 2 9 12 2 2 11 12 2 11 12 2 11 12 2 11 11 12 2
50 9 12 2 11 12 11 12 2 11 12 11 12 2 1 9 15 12 11 12 2 11 12 9 12 2 9 12 11 12 2 11 12 11 12 2 11 12 11 12 2 11 12 11 12 2 11 12 11 12 2
21 10 9 2 11 12 2 11 12 2 11 12 2 9 12 2 11 12 2 11 12 2
8 11 13 1 9 11 10 0 2
16 15 9 12 16 13 9 9 13 14 11 1 9 1 9 0 2
40 1 9 12 13 11 11 2 3 9 10 9 2 11 2 7 11 2 16 9 15 0 2 13 3 1 11 11 7 13 1 15 1 15 9 1 9 11 1 9 2
22 1 15 13 1 11 11 1 10 11 7 13 13 1 11 1 11 1 9 11 11 7 11
16 11 13 9 0 3 16 4 13 13 1 11 1 1 10 9 2
18 15 13 14 11 3 13 14 11 11 2 9 11 11 11 2 16 13 2
29 1 9 10 9 1 15 11 2 13 1 15 1 10 9 2 13 3 1 11 1 9 15 14 9 9 0 1 9 2
18 12 1 11 13 10 9 10 0 1 9 9 0 10 9 7 1 11 2
20 10 3 2 13 9 0 3 1 10 9 2 9 9 13 9 0 14 9 0 2
14 1 10 9 13 1 10 9 1 9 0 1 15 9 2
17 10 9 2 14 15 2 2 16 13 1 11 2 13 2 11 2 2
10 9 9 0 13 9 1 10 9 11 2
10 13 1 11 7 2 13 2 14 11 2
9 3 1 11 13 7 13 1 11 2
22 16 10 9 9 9 13 1 9 10 13 12 9 9 0 7 11 11 15 1 15 11 2
8 1 10 9 10 0 9 9 2
14 14 15 13 9 1 10 15 1 10 9 15 3 13 2
7 15 3 13 1 15 9 2
6 15 3 13 14 15 2
40 13 14 15 2 16 13 14 11 11 1 9 1 10 9 2 16 9 15 13 1 9 0 1 10 9 2 7 1 10 10 9 15 13 1 10 9 14 9 15 2
25 13 14 15 2 16 15 13 14 11 11 13 1 10 9 2 13 9 2 7 3 13 1 10 9 2
13 15 2 1 9 2 3 10 9 7 3 9 9 2
19 7 3 1 10 9 10 12 9 9 16 13 1 10 9 11 12 1 11 2
34 11 11 13 1 11 1 9 9 2 11 11 13 1 11 2 11 11 13 1 11 9 2 7 3 12 9 9 16 13 1 3 16 13 2
6 3 3 12 1 11 2
8 0 16 9 13 14 11 11 2
10 3 16 15 2 1 9 15 2 13 2
3 9 0 2
2 9 2
10 9 12 7 13 1 10 9 10 9 2
30 13 7 13 7 13 3 7 3 2 3 7 3 7 3 2 0 7 0 7 0 1 1 10 9 10 3 13 10 15 2
11 11 16 3 13 2 11 16 9 3 13 2
19 13 9 1 10 9 2 11 13 11 7 10 9 10 15 3 3 15 9 2
6 9 13 3 9 15 2
33 3 16 4 13 13 9 9 0 2 13 3 1 9 3 2 0 2 1 9 13 9 7 0 14 11 11 16 13 1 9 12 12 2
16 11 11 13 0 7 13 14 12 1 11 1 10 9 10 0 2
43 1 11 13 9 1 9 15 2 12 9 13 3 2 11 12 2 11 12 2 11 12 2 11 12 2 7 10 9 11 13 3 14 9 15 7 13 12 9 2 12 9 2 2
6 11 13 13 9 0 2
20 9 15 10 0 2 9 0 0 7 9 0 3 14 9 10 9 11 7 11 2
9 11 13 1 10 9 1 9 0 2
14 10 9 13 1 9 15 14 11 1 10 9 10 12 2
11 9 15 14 11 13 14 11 1 9 9 2
44 12 9 0 14 11 1 9 2 1 9 9 0 14 11 7 11 2 7 9 0 14 11 2 12 9 1 10 9 10 12 2 13 14 10 9 10 0 16 13 1 1 10 9 2
34 1 10 9 10 0 2 14 10 9 3 13 4 1 9 2 13 11 1 9 0 1 9 15 14 11 2 16 13 9 1 9 10 9 2
26 11 13 13 1 13 14 9 10 9 1 10 9 10 0 16 13 1 15 1 10 9 16 13 1 11 2
25 1 9 13 10 9 1 9 9 13 14 9 10 9 10 0 14 10 9 7 13 1 9 9 0 2
14 1 9 10 9 3 13 10 9 9 7 1 9 15 2
37 1 9 15 14 11 11 2 13 9 0 1 10 9 7 13 14 10 9 2 12 2 9 12 2 2 12 2 9 12 2 2 12 2 9 12 2 2
29 1 9 3 13 9 1 10 9 10 0 10 0 14 11 2 16 13 12 9 7 13 14 9 9 15 1 9 0 2
13 11 7 11 16 13 1 15 2 13 1 12 9 2
11 7 15 3 3 4 13 13 14 10 9 2
