241 11
21 13 10 9 7 10 9 15 2 10 15 13 1 0 9 10 9 2 14 13 3 2
15 3 13 12 9 1 9 1 14 13 0 10 9 10 9 2
23 13 7 10 9 15 10 9 13 10 0 9 10 0 9 1 10 9 10 9 10 9 15 2
23 1 9 15 2 13 14 13 10 0 9 10 9 2 1 15 13 14 13 7 9 1 9 2
26 10 9 10 0 9 0 10 9 2 3 13 10 0 9 10 0 2 13 10 9 13 0 9 10 9 2
22 1 9 10 9 2 10 9 13 0 7 0 10 15 3 3 1 15 2 1 9 9 2
15 13 1 10 9 0 9 1 10 0 9 7 10 9 9 2
28 10 9 10 9 1 9 13 7 2 10 0 9 13 9 12 1 9 15 13 9 2 1 9 1 10 12 2 2
28 1 3 10 9 9 9 13 1 0 9 15 13 14 13 1 9 1 9 14 13 0 14 13 9 1 0 9 2
20 10 9 9 2 0 1 10 0 9 10 9 2 13 0 9 1 9 10 9 2
32 10 9 10 9 2 10 9 7 10 0 9 13 14 13 3 1 15 15 9 1 10 9 7 10 9 10 9 7 10 9 15 2
34 10 9 1 0 9 2 7 0 9 13 14 13 0 2 15 9 13 14 13 0 9 1 9 7 14 15 13 1 10 0 7 0 9 2
38 0 9 13 7 2 10 0 9 15 13 10 9 10 9 10 9 9 13 7 13 13 0 9 7 13 10 9 7 10 9 9 14 13 3 10 9 2 2
8 10 9 9 13 10 9 15 2
15 13 1 10 9 10 0 9 14 13 10 9 0 9 2 2
37 10 9 9 13 1 2 2 7 10 12 15 13 10 0 9 7 10 12 13 1 10 9 10 9 7 13 1 12 9 9 2 7 1 9 13 0 2
33 9 10 9 2 9 7 10 9 9 9 13 7 10 12 10 9 13 7 10 9 1 9 14 13 10 0 9 7 10 9 0 9 2
11 12 9 3 2 10 9 13 10 9 13 2
4 13 0 9 2
17 1 9 10 9 13 1 10 9 2 9 3 13 2 10 9 9 2
34 1 9 10 9 13 1 9 1 9 10 12 0 0 2 1 10 9 10 12 15 13 13 1 9 1 9 9 15 13 1 10 9 9 2
31 10 9 9 13 10 0 15 1 10 9 2 7 13 7 10 9 14 13 10 0 14 13 10 9 15 7 14 13 10 9 2
37 10 0 9 13 10 0 9 2 15 13 10 0 9 1 9 10 9 2 7 15 13 0 1 0 2 1 10 0 7 0 9 7 3 1 10 9 2
33 3 3 10 0 10 9 14 13 0 2 10 2 13 0 1 10 9 10 9 9 7 10 9 10 9 3 1 9 7 10 9 0 2
15 2 7 9 13 0 9 1 10 9 10 9 9 1 9 2
39 10 9 10 9 13 1 9 10 0 9 10 9 1 9 2 10 15 13 10 9 2 13 0 9 1 0 9 1 10 9 2 7 3 13 0 9 7 9 2
26 10 9 13 3 10 9 14 13 0 9 1 0 9 7 13 0 9 7 9 7 10 9 13 10 9 2
52 1 9 10 9 13 10 9 10 0 2 10 0 9 10 9 1 10 0 9 2 10 9 10 9 13 7 13 1 9 10 9 10 0 9 7 10 0 9 10 9 13 10 12 9 7 13 0 0 7 0 9 2
11 13 10 12 12 10 9 9 1 0 9 2
24 10 9 14 13 10 3 9 10 9 15 1 9 2 15 7 15 15 15 13 10 9 1 9 2
36 10 9 9 2 13 0 13 9 15 13 9 13 1 9 7 10 9 9 13 3 1 0 9 10 0 9 2 7 1 0 9 10 9 10 9 2
27 10 0 9 1 10 0 9 9 1 9 10 9 12 13 3 10 9 2 10 9 2 1 9 10 9 15 2
1 9
9 13 3 9 7 13 3 1 0 2
21 10 0 9 10 2 14 13 1 10 9 9 7 1 10 9 9 2 9 7 9 2
52 10 0 9 13 1 10 9 15 2 10 9 1 9 2 13 10 9 15 13 3 3 1 10 0 9 10 9 10 0 9 15 13 1 3 7 14 13 14 13 7 1 9 2 9 2 13 9 10 0 15 9 2
9 9 2 9 3 1 10 0 9 2
28 10 0 13 7 2 1 12 9 13 10 12 9 1 10 9 10 9 10 0 9 2 7 3 13 10 12 9 2
50 3 3 2 0 9 13 10 9 1 0 9 2 1 10 15 7 14 13 10 9 0 0 9 7 10 0 0 1 10 9 7 13 10 0 1 9 9 10 0 0 9 10 15 13 1 0 9 7 9 2
6 7 13 9 14 13 2
36 10 0 9 10 9 13 1 12 9 2 13 10 9 10 0 0 9 1 9 10 9 2 7 7 9 15 13 0 9 1 9 7 1 0 9 2
33 10 9 2 13 1 10 9 10 0 9 2 2 10 9 2 10 9 7 10 9 13 10 0 9 10 9 7 13 10 9 15 13 2
20 10 9 13 1 0 3 10 0 9 1 0 9 9 2 15 13 13 10 9 2
25 7 14 13 0 0 9 9 2 10 9 14 13 1 9 10 9 9 1 9 3 1 10 0 9 2
7 3 10 0 9 13 0 2
31 3 2 13 1 10 9 2 3 1 9 12 9 2 3 10 9 2 7 3 1 0 9 2 7 14 14 13 3 10 9 2
34 3 3 13 2 10 0 9 13 3 7 9 10 9 7 13 14 15 13 3 1 10 0 9 10 9 2 3 1 9 15 13 13 3 2
18 1 9 2 3 10 0 0 9 14 13 13 1 9 2 13 3 9 2
29 10 9 9 13 3 10 9 10 1 9 9 7 13 10 9 3 10 9 3 7 10 9 1 0 10 9 10 9 2
16 3 2 1 10 9 2 13 9 15 14 13 3 10 0 9 2
15 13 15 3 12 9 1 14 13 9 7 14 3 14 13 2
1 9
15 13 7 10 9 9 13 10 0 9 10 9 1 9 12 2
18 12 1 10 9 10 9 13 14 13 10 9 10 14 13 0 1 9 2
4 2 2 1 2
40 1 10 9 15 13 3 0 14 13 15 10 9 2 3 7 10 9 10 9 15 14 13 0 1 15 10 9 1 10 0 9 9 2 9 7 10 9 0 9 2
39 14 13 3 10 9 2 3 1 10 15 14 13 1 9 10 9 7 13 13 3 3 10 9 10 0 9 13 1 9 9 10 9 0 9 10 9 10 9 2
25 7 2 10 0 9 13 9 1 0 9 0 0 9 14 13 9 1 9 2 1 0 9 7 9 2
28 10 0 9 2 13 10 0 9 2 1 9 10 9 2 10 15 13 1 10 9 10 9 14 13 3 1 9 2
16 10 9 9 10 9 13 0 2 7 10 9 10 9 13 0 2
10 10 0 9 14 13 1 12 9 2 2
20 13 14 13 7 2 3 1 10 0 15 9 2 10 9 10 9 13 3 3 2
5 1 9 10 9 2
33 3 13 10 0 0 9 2 10 9 9 2 9 7 9 15 13 1 9 10 9 2 13 1 10 9 9 2 9 9 7 0 9 2
25 1 10 9 10 9 10 9 2 10 9 13 10 0 15 9 2 13 10 9 7 13 10 9 9 2
37 7 13 3 14 13 10 9 1 0 9 7 1 0 9 2 14 13 14 13 10 9 9 1 0 9 15 14 13 10 9 14 13 7 14 13 3 2
17 3 0 9 13 10 9 15 13 1 0 9 1 10 0 0 9 2
42 10 9 10 9 13 0 2 7 13 7 9 1 10 9 10 9 2 7 7 1 10 9 2 10 9 2 10 9 2 10 9 2 10 9 2 10 9 7 10 9 9 2
11 3 13 10 9 7 10 9 9 1 9 2
14 15 15 13 1 9 3 13 15 9 9 14 15 13 2
5 15 13 13 3 2
17 10 9 3 1 9 13 14 13 7 14 13 0 7 10 9 15 2
18 3 12 9 13 1 10 9 1 9 2 13 10 9 3 1 9 9 2
19 1 15 14 13 1 9 10 9 15 13 10 2 9 1 9 10 9 2 2
48 10 9 9 10 2 2 9 9 2 13 1 9 2 9 2 10 0 9 2 3 1 9 15 10 9 15 13 10 9 1 9 7 9 2 10 15 7 14 13 13 0 9 7 15 0 9 9 2
34 10 9 15 13 13 10 9 9 2 9 7 9 15 13 14 13 7 14 13 10 9 10 9 9 2 1 7 14 13 10 15 13 3 2
19 10 9 15 10 9 2 10 15 13 1 9 10 12 2 13 3 0 9 2
9 7 2 10 9 13 14 13 3 2
14 13 7 0 10 9 1 14 13 9 1 15 13 0 2
32 0 13 7 10 0 9 9 2 1 15 13 9 1 9 1 9 7 10 9 7 10 9 10 9 9 2 10 15 13 3 9 2
33 3 13 10 0 10 9 1 10 9 15 13 10 2 9 9 2 13 14 13 7 10 0 10 2 9 9 13 14 13 3 0 9 2
16 13 9 12 9 7 13 1 10 0 9 7 0 0 9 15 2
14 10 9 13 13 1 9 7 14 13 10 9 10 9 2
37 1 10 9 15 10 9 10 9 2 9 9 2 13 9 1 10 9 10 9 9 7 2 14 13 0 10 0 9 3 1 10 0 9 10 9 2 2
27 1 10 0 9 7 10 9 13 0 9 1 10 9 7 10 0 9 10 9 2 1 0 9 7 0 9 2
18 2 10 9 15 13 7 10 9 10 0 9 1 10 9 14 13 0 2
25 1 9 10 0 9 2 1 3 2 13 13 10 9 10 0 9 10 9 2 10 9 10 0 9 2
11 1 10 9 2 10 9 13 14 13 3 2
30 12 13 10 3 9 10 9 2 9 9 2 7 10 0 0 1 10 0 0 9 1 9 2 10 9 9 2 13 12 2
20 10 9 13 1 10 9 9 15 13 13 7 13 2 3 1 10 9 10 9 2
8 10 9 10 9 13 9 1 9
17 13 14 13 3 9 9 10 9 10 15 10 0 13 13 1 9 2
14 10 0 9 1 9 9 13 14 13 10 9 10 9 2
20 10 9 10 9 13 13 10 9 10 0 0 9 1 9 3 3 1 10 9 2
24 7 13 9 7 15 14 13 3 2 13 10 1 9 9 7 7 13 9 9 15 13 10 9 2
10 13 0 9 1 10 9 10 9 15 2
26 3 2 10 9 13 10 9 1 9 12 2 1 10 9 10 0 9 1 9 10 12 10 9 9 12 2
27 1 15 13 0 15 10 9 1 9 2 15 13 1 9 9 10 0 9 2 14 13 9 1 15 10 9 2
17 13 2 9 9 2 7 10 9 13 14 13 3 0 10 0 9 2
27 13 10 9 2 7 10 9 13 14 13 10 0 9 9 7 14 13 1 15 1 14 13 10 0 0 9 2
38 10 9 1 15 13 10 9 15 13 7 15 10 9 10 9 13 14 13 3 2 13 10 9 9 9 14 3 1 15 1 9 2 7 7 1 3 9 2
23 10 9 9 10 9 2 9 9 9 2 13 7 2 10 9 15 14 14 13 1 9 2 2
24 13 10 0 9 2 1 10 9 10 9 2 15 13 9 9 7 13 10 9 1 10 9 9 2
20 9 10 0 9 10 9 7 10 9 9 13 2 1 9 9 9 14 13 13 2
34 7 14 13 10 9 1 10 15 10 9 9 13 0 7 0 2 10 9 15 13 0 1 10 0 0 9 1 9 1 10 9 10 9 2
34 10 9 15 13 3 1 2 7 10 0 9 2 3 1 9 1 9 7 13 12 9 1 10 9 10 9 10 0 9 2 9 9 9 2
8 10 9 13 10 9 1 9 12
11 12 9 13 3 1 10 9 9 10 9 2
13 13 1 10 0 9 2 7 7 13 10 9 9 2
20 13 10 9 10 0 9 9 12 2 3 13 0 0 9 2 1 9 12 9 2
1 9
16 13 7 13 14 13 10 9 15 3 7 14 15 13 0 9 2
31 3 2 10 9 9 13 3 1 10 9 9 10 9 2 9 9 2 3 7 1 10 9 9 10 0 9 2 9 9 9 2
26 7 15 2 3 13 10 2 9 2 13 9 9 0 15 0 9 2 1 10 15 7 10 0 10 9 2
27 3 3 10 9 13 9 10 9 9 2 13 3 10 9 9 1 10 9 1 9 3 1 10 9 10 9 2
17 1 15 2 13 15 14 13 3 1 10 9 7 1 9 1 10 9
26 1 10 9 2 10 9 13 1 2 2 3 13 1 9 10 9 2 7 10 12 13 1 9 1 9 2
16 10 0 9 10 15 10 0 9 0 9 10 9 13 14 13 2
35 10 9 0 9 14 13 9 10 12 9 2 7 13 9 15 13 1 15 9 7 10 9 13 7 15 14 13 1 9 14 13 10 0 9 2
17 10 0 10 9 13 9 12 9 7 13 10 9 9 9 12 9 2
28 10 9 1 10 0 0 9 2 1 10 9 10 0 10 9 2 1 10 9 2 9 2 13 1 12 9 9 2
5 13 1 0 9 2
23 13 14 13 14 13 7 10 9 9 14 13 14 13 1 9 10 9 15 1 10 9 9 2
48 10 9 10 0 9 1 10 9 9 1 9 7 10 0 9 1 10 9 10 9 10 9 2 13 10 9 10 9 10 9 14 13 1 9 15 7 3 10 9 1 10 9 10 9 1 10 9 2
25 7 2 10 9 2 3 10 9 2 13 9 10 0 7 10 0 9 2 7 10 2 13 15 9 2
14 1 9 15 10 9 7 10 9 13 14 13 0 9 2
31 9 9 2 10 9 9 3 1 10 9 9 9 13 14 13 0 10 9 15 13 1 9 9 3 10 0 9 10 0 9 2
35 1 12 9 10 15 13 9 1 9 10 9 9 0 9 7 9 10 9 2 13 0 9 1 9 14 13 3 10 0 9 1 10 0 9 2
45 3 1 10 0 0 9 1 10 0 9 2 2 0 1 12 9 9 13 9 1 12 9 2 9 10 0 9 2 7 0 0 13 3 10 9 9 1 0 9 7 10 0 9 2 2
39 3 13 14 13 9 7 14 13 7 15 15 13 0 1 9 2 9 2 9 7 1 9 1 9 10 9 7 10 0 10 9 13 14 13 1 10 0 9 2
24 3 1 9 10 9 9 2 10 9 13 12 9 9 2 7 10 9 15 14 13 10 0 9 2
64 10 9 13 3 10 9 15 13 10 0 9 1 9 10 9 1 9 15 13 1 9 10 0 9 3 1 10 0 7 10 0 9 7 1 15 15 13 10 0 2 0 7 0 9 2 7 13 10 9 15 14 13 10 9 3 10 0 3 7 10 12 15 9 2
31 13 0 9 1 10 2 2 1 15 0 9 13 2 7 10 9 13 3 1 9 10 9 13 7 10 9 7 10 9 2 2
24 13 7 13 1 3 10 9 14 13 10 9 15 7 2 7 13 3 2 14 13 10 0 9 2
18 10 9 10 9 9 13 3 9 14 13 9 10 9 10 9 9 9 2
16 10 0 9 0 9 13 1 0 9 2 13 10 0 9 9 2
29 3 2 7 13 10 9 10 9 10 9 7 10 9 2 14 13 3 9 2 7 10 9 13 3 9 1 15 9 2
17 14 13 1 15 9 10 9 7 10 9 1 10 9 13 1 9 2
13 14 13 14 13 0 15 9 1 10 9 10 9 2
16 13 9 9 10 12 9 2 10 9 13 14 13 10 9 15 2
10 10 0 9 10 9 13 3 1 9 2
18 3 2 7 2 14 13 3 14 13 2 7 7 14 13 7 14 13 2
47 3 15 2 10 9 13 15 0 9 2 0 0 9 2 10 14 9 3 7 12 9 10 0 9 2 9 15 15 13 1 9 15 13 9 10 0 9 2 15 13 12 1 10 9 10 9 2
20 13 14 13 10 9 14 13 1 10 9 7 10 9 10 9 7 14 13 9 2
30 10 9 15 9 14 13 0 2 7 3 13 3 3 10 9 1 10 12 9 2 10 15 13 14 13 3 1 0 9 2
35 1 15 10 9 14 13 10 9 15 13 0 9 1 0 9 3 9 10 0 9 15 13 13 1 9 10 9 0 9 1 0 10 0 9 2
26 3 1 9 2 10 0 9 13 7 13 2 3 0 2 9 1 10 9 10 9 1 10 9 1 2 2
38 10 9 14 13 14 13 12 0 9 2 12 15 14 13 1 9 9 3 3 1 9 15 2 7 12 15 15 14 13 1 9 9 7 15 13 0 9 2
17 3 2 9 9 2 14 13 1 9 3 1 10 9 7 10 9 2
19 10 9 13 13 3 7 2 2 3 13 10 9 2 13 0 10 9 2 2
32 3 1 9 2 1 9 10 15 1 12 9 3 10 12 9 13 14 13 9 1 9 15 2 9 0 1 15 15 13 10 2 2
18 13 14 13 1 10 9 2 10 2 13 9 9 1 9 1 9 9 2
32 3 2 10 0 9 13 1 9 10 0 9 7 13 14 13 10 9 15 1 9 7 10 9 10 9 7 1 9 1 10 9 2
4 10 9 9 2
21 9 9 2 13 10 0 9 15 1 9 15 7 10 2 13 14 13 10 9 15 2
23 13 3 10 9 14 13 12 9 10 9 10 9 15 7 10 0 15 13 0 10 12 9 2
18 9 9 2 14 13 7 15 14 15 13 1 10 9 15 3 12 9 2
56 3 2 13 10 9 10 0 9 15 14 13 15 9 1 9 15 1 14 13 15 10 9 7 14 13 14 13 3 7 10 9 9 13 1 9 10 0 9 1 10 9 15 13 1 9 10 9 2 14 13 9 1 15 10 9 2
26 9 10 9 10 9 9 13 7 2 10 9 10 9 10 9 9 13 7 13 10 9 7 14 13 3 2
36 15 14 13 2 7 3 13 10 9 2 7 13 7 1 10 0 9 2 7 13 1 9 15 0 9 3 1 10 9 10 9 7 10 0 9 2
33 10 9 10 9 13 7 2 10 0 9 10 9 13 13 10 0 9 2 7 3 10 12 10 9 9 12 9 13 1 15 10 9 2
10 15 10 9 13 14 13 14 13 0 2
3 2 9 2
23 3 1 10 9 10 9 13 1 9 10 9 9 2 10 15 7 13 10 9 15 1 9 2
48 3 10 9 10 9 3 7 10 9 1 9 15 13 9 3 1 15 7 10 9 13 14 13 0 9 1 10 9 10 0 9 10 9 10 0 9 7 10 9 15 14 13 1 9 1 15 9 2
40 1 15 10 9 13 3 0 7 13 7 13 10 0 9 1 9 2 7 1 0 9 10 9 9 1 10 0 0 9 14 13 15 10 0 9 9 15 13 3 2
42 7 2 15 9 3 10 9 2 10 9 2 10 2 7 3 10 9 13 1 10 9 2 7 15 13 10 0 9 7 2 14 13 1 0 9 9 1 10 9 15 2 2
38 13 0 1 10 9 9 7 10 9 9 7 1 10 0 9 10 9 7 10 9 10 0 0 9 13 14 13 9 1 9 7 1 10 3 0 0 9 2
3 15 13 2
53 7 2 13 7 3 1 10 9 9 13 10 0 9 7 1 0 9 10 0 9 1 15 15 0 1 15 13 14 13 7 13 0 1 10 0 9 10 0 9 3 13 10 9 10 9 10 9 10 9 1 15 13 2
40 13 15 14 13 1 9 3 9 2 7 13 7 10 9 13 14 13 10 9 2 12 7 13 10 9 2 12 2 12 2 12 2 12 2 12 2 12 7 12 2
10 9 15 13 10 9 14 13 10 0 9
10 9 2 9 0 9 1 10 9 9 2
42 1 9 2 3 1 10 9 10 9 2 10 9 13 10 9 10 9 12 2 10 15 2 13 10 0 7 0 9 10 9 2 15 13 2 15 13 7 15 13 1 9 2
33 3 2 14 13 14 13 1 9 10 0 9 7 10 0 9 2 7 7 1 9 10 9 1 0 9 2 1 10 12 2 12 9 2
39 1 14 13 10 9 1 10 9 0 9 10 9 1 10 9 2 10 9 15 14 13 14 13 10 9 15 1 10 9 15 2 7 3 3 1 10 9 15 2
6 1 15 15 13 7 2
28 10 9 9 13 13 1 0 9 1 9 15 2 10 12 2 1 9 1 0 9 2 1 10 15 13 12 9 2
22 1 9 13 10 0 9 2 10 0 10 9 7 1 9 13 10 9 10 9 10 9 2
16 10 0 9 13 1 9 10 9 7 10 9 3 13 0 9 2
6 3 13 10 12 9 2
15 9 10 9 9 1 9 9 7 9 1 0 9 10 0 2
42 1 15 3 1 15 9 2 13 10 0 9 12 9 2 9 10 9 9 12 1 9 10 12 2 9 2 10 15 13 13 7 15 9 13 10 9 10 9 9 2 9 2
7 10 12 9 13 3 0 2
21 10 9 13 9 1 0 9 10 2 1 9 2 7 10 9 2 0 3 2 13 2
21 3 2 1 9 14 13 9 1 10 7 10 9 9 14 13 1 9 15 1 9 2
14 0 1 12 9 13 13 9 2 13 10 9 0 9 2
6 14 13 10 0 9 2
28 10 9 15 13 3 10 2 9 13 3 10 0 2 3 3 7 0 2 9 10 9 15 13 1 9 10 9 2
11 10 9 9 13 1 10 9 9 1 9 12
33 15 9 2 3 0 7 7 13 2 13 9 3 7 13 1 0 9 10 9 15 2 7 3 1 10 0 9 1 0 10 9 9 2
24 10 9 13 14 13 15 9 10 9 3 2 7 10 0 0 9 14 14 13 0 10 0 9 2
14 2 10 9 9 13 3 0 2 2 13 9 10 9 2
9 9 2 1 10 0 9 1 10 9
33 10 1 9 9 13 3 1 9 9 2 1 1 9 9 10 9 2 10 15 7 15 13 1 9 9 7 1 15 13 1 0 9 2
12 13 1 0 10 0 9 10 9 10 0 9 2
19 7 13 14 13 10 9 15 3 0 9 2 3 13 14 13 1 0 9 2
13 3 2 7 2 13 10 0 7 1 10 0 9 2
33 3 1 9 10 9 2 13 10 0 0 9 1 10 12 9 15 13 10 9 15 2 10 9 2 10 9 2 10 9 7 10 9 2
38 9 13 13 1 0 9 3 1 0 9 1 10 0 9 9 9 2 9 2 2 1 0 0 9 1 12 9 15 13 1 9 2 10 9 7 15 9 2
4 10 9 9 2
20 0 1 10 9 13 9 3 2 0 15 2 2 7 2 9 1 10 9 2 2
18 1 10 9 15 2 10 9 13 14 13 1 9 15 10 9 10 9 2
11 10 9 13 3 9 1 10 9 0 9 2
55 13 14 13 7 1 15 9 10 9 13 3 0 7 7 10 9 10 12 9 13 1 10 9 15 10 9 15 13 1 0 9 9 2 13 3 1 9 15 9 9 10 9 14 13 15 3 0 0 9 1 10 0 0 9 2
14 7 2 10 9 15 14 13 14 13 10 9 15 9 2
27 1 10 0 2 2 9 15 10 0 9 13 10 9 2 10 9 3 10 9 7 10 0 9 9 2 9 2
17 10 0 9 2 7 2 13 7 2 15 9 14 13 1 9 2 2
32 10 0 9 15 1 10 9 9 1 10 9 9 13 13 10 2 2 10 15 13 7 2 10 0 9 13 14 13 0 9 2 2
38 9 9 2 15 13 3 0 1 10 7 13 1 10 9 14 13 1 0 9 2 1 9 15 2 9 1 10 0 1 9 9 3 1 10 9 10 9 2
20 12 3 9 2 15 13 1 9 2 10 9 9 9 2 13 0 10 0 9 2
36 10 0 9 13 14 13 1 9 1 10 9 10 0 9 15 13 13 10 9 10 9 7 13 3 14 13 1 0 9 14 13 10 9 10 9 2
17 10 9 13 3 1 9 7 10 0 9 1 10 9 13 3 0 2
22 1 9 1 2 9 9 2 10 9 13 3 9 1 0 9 3 1 10 9 15 13 2
29 13 7 14 13 9 7 7 10 0 10 9 10 9 13 13 7 10 9 10 9 14 14 13 13 3 1 10 9 2
14 10 9 13 10 9 10 9 1 12 9 1 1 12 2
24 3 1 9 2 13 3 1 15 2 13 10 9 2 10 9 0 0 9 2 0 9 7 9 2
12 10 9 10 0 9 13 3 14 13 14 13 2
21 1 10 0 9 13 10 12 0 9 10 0 9 1 14 13 1 9 1 0 9 2
20 10 0 9 13 10 3 0 9 2 13 7 13 13 3 7 13 14 13 3 2
21 12 9 13 14 13 1 9 10 9 2 1 9 2 7 10 9 13 9 1 9 2
38 10 9 15 14 14 13 2 3 7 7 13 1 9 9 1 15 9 2 14 13 10 9 7 10 9 10 9 2 10 15 13 10 0 9 0 0 9 2
8 10 9 13 9 9 15 1 2
25 2 3 1 10 9 15 2 10 2 14 13 10 0 9 1 9 10 9 2 2 13 10 9 9 2
39 0 15 13 14 13 10 0 9 1 10 9 2 1 9 10 9 2 10 9 15 13 3 0 1 9 1 10 9 10 13 1 10 9 9 7 1 10 9 2
27 10 0 9 9 2 9 9 2 13 7 10 0 9 1 9 10 9 13 3 2 13 3 2 10 0 9 2
8 10 15 9 14 13 3 0 2
8 1 15 13 14 13 10 12 2
32 3 13 14 13 10 9 7 14 13 10 9 15 9 10 9 15 2 10 3 0 9 2 3 14 13 3 10 9 15 14 13 2
15 10 9 10 0 9 13 3 10 0 9 10 9 10 9 2
31 1 15 13 3 2 13 0 10 0 9 15 13 1 9 9 10 9 9 9 2 9 0 7 12 1 10 0 9 10 9 2
22 10 9 13 0 1 2 3 10 9 7 10 9 7 1 9 1 9 7 3 1 9 2
26 10 9 15 13 7 10 9 2 10 15 13 10 9 14 2 14 13 9 15 14 13 9 1 9 2 2
25 10 9 10 0 9 2 9 9 2 1 12 9 13 0 9 1 9 2 7 13 1 9 10 9 2
25 1 14 13 2 14 13 10 0 7 0 9 1 9 3 14 13 10 9 10 9 1 10 0 9 2
21 7 10 9 10 0 9 10 9 13 0 2 10 9 1 10 9 10 9 13 0 2
25 3 14 13 9 7 10 9 13 1 15 9 14 13 9 9 10 9 2 7 13 14 15 13 15 2
12 10 9 15 14 13 3 13 9 15 10 9 2
42 3 2 1 9 9 9 0 9 14 13 10 9 10 15 14 13 14 13 10 0 7 3 2 3 1 9 10 0 9 2 10 9 10 9 13 14 13 1 9 10 9 2
5 14 13 15 9 2
25 10 9 13 9 7 9 1 14 13 1 12 10 9 2 1 10 9 14 13 9 1 9 12 9 2
