559 17
23 11 9 9 13 9 1 9 0 1 9 2 9 2 9 2 7 9 0 15 13 9 9 2
35 11 11 13 1 9 0 2 3 0 1 9 11 11 2 0 1 9 11 11 2 0 1 11 11 11 2 7 0 3 1 9 11 11 11 2
51 9 10 3 13 1 10 9 9 15 2 1 2 11 11 11 7 11 11 11 2 2 9 11 11 1 15 3 13 1 9 2 3 13 9 1 11 7 9 9 11 2 7 7 9 9 9 7 11 9 9 2
14 16 11 13 9 3 9 15 13 1 9 7 9 14 2
8 11 11 11 13 9 9 12 2
18 12 9 13 1 9 12 9 2 12 9 1 11 7 10 9 1 11 2
21 11 11 9 11 13 1 13 9 9 2 9 9 2 7 9 9 1 9 9 9 2
35 9 9 3 0 1 11 1 3 7 9 9 9 12 2 12 7 12 1 9 9 0 2 1 9 13 0 1 13 9 9 13 1 9 12 2
14 11 9 10 11 11 1 9 11 11 1 9 15 0 2
39 9 10 3 13 9 2 9 1 11 11 12 9 11 2 11 9 11 11 9 12 2 11 2 12 2 11 13 9 11 11 1 9 9 13 9 11 7 11 2
28 9 2 9 0 3 13 3 3 1 13 10 9 15 3 13 1 9 9 0 1 9 9 9 7 9 9 9 2
22 11 13 1 9 9 10 9 15 13 1 9 9 2 16 1 9 9 14 13 1 10 2
9 16 3 1 9 9 11 7 11 2
22 9 9 13 1 11 11 11 2 15 13 1 11 11 1 9 12 1 11 9 2 11 2
24 11 13 10 9 9 1 10 9 0 9 7 9 0 9 15 13 9 7 9 10 14 13 3 2
16 3 11 11 1 9 13 9 11 15 3 0 1 12 9 9 2
14 11 3 13 1 11 2 7 15 13 3 13 1 11 2
16 11 9 11 13 0 1 9 9 11 11 1 9 12 2 12 2
17 9 1 11 11 11 3 13 15 13 9 7 9 15 10 2 10 2
25 11 0 7 9 2 11 3 13 7 13 9 9 15 1 9 2 9 9 11 1 9 7 9 0 2
38 9 0 1 9 9 9 13 9 9 2 9 2 9 2 11 2 11 2 11 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 2
14 11 11 1 11 2 2 9 0 3 15 13 1 11 2
33 11 2 9 10 13 1 9 12 12 9 7 10 9 11 13 9 1 9 15 13 16 10 9 14 3 13 9 9 0 1 9 11 2
20 9 10 3 13 1 9 15 13 11 11 11 15 13 1 11 1 12 11 12 2
13 7 9 0 13 11 11 2 13 10 9 13 11 2
29 3 9 13 1 9 2 15 3 13 1 2 9 2 16 1 10 9 15 3 13 12 1 9 15 3 13 9 0 2
6 11 3 13 9 9 2
13 11 13 9 11 1 9 9 7 9 15 13 9 2
3 1 9 2
43 1 13 9 2 9 9 3 13 9 9 9 15 0 2 3 9 9 9 15 13 9 2 9 7 9 15 3 1 1 9 1 0 1 9 9 7 9 2 9 2 7 9 2
4 3 13 11 2
8 9 15 0 13 13 0 9 2
7 3 10 9 13 9 0 2
34 11 11 5 9 9 13 10 9 9 1 9 9 2 9 15 13 1 9 9 2 9 15 13 1 9 9 7 12 1 12 9 11 11 2
22 1 11 12 2 7 9 9 1 11 2 11 7 11 11 9 10 13 9 13 11 11 2
16 10 2 10 0 9 13 10 9 2 9 9 15 0 7 0 2
77 11 11 0 1 11 2 11 11 2 16 14 0 16 10 9 11 0 10 3 13 9 2 1 1 11 2 11 2 11 11 2 11 11 2 11 11 2 11 2 11 11 2 11 2 11 11 2 11 11 2 11 2 11 2 11 2 11 11 2 11 2 11 11 11 2 11 2 11 2 11 11 2 11 2 11 11 2
41 11 11 7 11 11 2 12 5 12 2 12 11 12 2 2 13 2 11 2 1 9 13 9 11 15 13 1 11 11 2 13 9 11 1 12 11 1 12 11 12 2
11 3 1 11 11 15 3 0 13 1 11 2
16 7 16 15 3 14 13 1 9 2 3 15 13 1 1 9 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
7 11 11 12 2 12 12 2
11 1 13 2 9 10 3 13 1 11 11 2
66 1 9 12 2 11 11 11 11 11 11 2 11 2 2 1 9 15 13 1 11 11 11 11 11 11 2 11 2 1 12 1 9 12 2 13 9 1 9 9 9 1 9 1 9 0 2 16 1 9 10 3 13 16 9 9 1 9 14 3 0 1 13 1 0 9 2
25 9 2 9 11 13 16 11 3 0 2 0 9 3 13 9 2 11 7 11 2 11 1 12 9 2
6 9 3 15 13 9 2
29 9 10 13 1 9 15 14 13 1 9 9 11 1 11 11 7 13 1 9 11 11 7 9 9 9 2 13 2 2
43 11 11 2 11 2 13 1 11 2 10 9 9 9 9 9 15 13 9 13 1 11 11 10 13 1 9 2 9 9 0 15 2 1 1 9 9 11 2 11 2 7 11 2
11 11 11 15 13 9 11 11 13 1 9 2
19 9 9 11 2 11 13 9 2 1 9 9 15 3 10 2 10 12 9 2
18 9 10 13 9 1 9 15 2 3 13 9 1 13 9 1 9 9 2
27 11 2 15 13 10 9 3 13 1 10 9 9 2 13 11 16 13 9 11 11 7 13 1 9 11 11 2
33 16 2 1 9 2 9 10 13 1 11 11 7 11 11 11 1 9 12 11 12 1 9 11 11 11 11 11 11 2 12 2 12 2
24 13 13 14 13 1 9 7 9 15 13 1 9 9 3 13 1 9 7 9 1 9 0 10 2
11 1 9 15 14 11 11 11 11 3 13 2
27 10 9 3 0 13 16 15 13 9 10 13 9 9 9 7 9 9 2 11 11 0 2 12 2 12 2 2
43 16 3 10 9 1 11 11 1 9 11 2 9 15 3 3 13 1 9 11 9 9 2 2 9 1 11 1 9 0 1 9 11 1 3 1 12 9 3 13 1 9 9 2
18 15 13 16 1 10 3 13 0 1 11 11 7 13 9 1 11 11 2
47 15 13 1 13 10 9 9 0 15 3 15 13 2 7 13 9 2 9 1 9 11 11 1 10 1 9 9 0 2 7 16 15 13 9 0 1 13 9 2 9 11 11 0 1 11 11 2
140 1 9 2 9 9 9 2 9 1 1 9 9 11 11 7 11 11 11 11 11 10 3 0 13 9 9 1 9 9 15 1 11 12 13 10 9 9 11 11 11 2 11 2 1 9 2 9 7 9 9 0 1 10 9 11 7 11 11 9 9 12 1 13 9 9 15 13 9 13 11 11 15 13 7 13 11 2 1 0 9 12 2 9 9 9 11 11 1 13 11 11 10 1 9 9 9 9 12 11 11 2 11 11 2 9 9 9 11 11 2 9 11 11 2 11 11 7 10 9 0 13 11 11 7 11 11 11 2 11 11 11 11 2 3 15 13 1 11 11 2
32 9 0 1 9 10 13 9 2 1 9 0 12 5 1 9 2 1 9 3 12 5 2 11 11 13 1 10 9 1 9 10 2
16 11 3 13 1 11 7 13 10 9 2 16 11 2 11 2 2
25 10 9 1 11 11 13 1 3 13 10 9 3 2 2 11 0 11 13 9 13 15 13 1 9 2
19 16 15 13 1 9 10 2 15 14 3 13 9 2 9 16 13 9 11 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
23 9 11 13 16 9 9 15 3 0 2 16 16 15 13 1 9 16 11 3 13 13 11 2
13 11 13 9 10 7 13 2 16 9 15 3 13 2
29 3 2 11 11 11 2 11 2 13 1 0 1 9 9 11 11 11 12 1 9 0 1 13 11 11 15 13 9 2
29 11 11 11 3 13 16 15 13 9 9 15 0 1 9 13 2 7 9 11 3 13 1 9 12 2 9 2 11 2
150 11 12 2 11 11 11 2 0 9 9 0 15 13 1 9 12 11 2 11 10 13 7 13 1 9 2 9 11 9 12 11 2 11 11 11 11 2 9 9 9 0 15 13 1 9 12 11 2 11 10 13 7 13 9 12 11 2 9 11 11 11 2 9 9 9 0 2 0 1 11 2 3 13 1 9 12 11 2 11 10 13 7 13 12 11 12 2 11 11 11 2 9 9 9 0 15 13 1 9 12 12 2 11 10 13 7 13 1 9 2 9 11 9 12 11 2 11 11 11 11 11 2 9 9 9 0 15 13 1 9 12 11 2 11 10 13 1 9 9 2 9 11 7 13 1 0 1 9 12 2
22 9 2 9 9 15 13 1 9 2 13 9 15 0 1 9 15 0 7 13 9 0 2
21 16 11 13 0 1 11 2 15 3 13 16 15 13 9 15 0 2 0 7 0 2
28 10 9 9 11 1 9 11 11 7 11 13 1 9 11 1 13 9 1 9 0 11 2 11 11 2 7 11 2
8 15 13 1 9 11 11 11 2
5 9 5 9 9 2
21 9 9 13 1 9 0 7 16 9 9 10 13 15 0 2 7 1 9 0 9 2
8 11 13 13 12 9 2 7 2
63 11 2 11 2 11 2 2 2 13 9 9 9 11 1 9 1 9 11 11 11 2 11 11 2 11 11 11 2 11 11 11 7 11 11 11 2 2 13 1 11 2 3 13 11 1 12 9 2 11 11 12 9 2 11 11 12 9 7 9 11 12 9 2
14 16 15 13 1 15 2 2 10 10 9 15 13 9 2
10 11 11 3 13 1 9 11 11 11 2
20 9 10 13 1 11 11 15 13 12 5 1 11 11 2 9 9 11 11 11 2
25 9 15 11 13 1 13 9 3 3 2 16 15 14 13 16 9 3 13 1 9 9 7 9 9 2
21 2 2 9 13 2 7 11 13 11 1 13 2 7 13 9 1 11 1 13 9 2
28 16 9 10 13 1 9 9 9 2 11 13 9 3 1 13 9 11 11 2 11 10 15 13 13 9 13 9 2
25 9 9 13 9 0 0 7 0 2 0 0 2 16 9 9 2 11 2 11 2 2 13 0 0 2
12 10 13 1 9 9 15 3 14 3 13 9 2
27 11 13 1 10 9 2 3 1 1 9 11 11 2 11 11 2 11 11 2 11 2 11 2 11 7 11 2
18 1 11 2 11 13 11 2 15 9 13 1 9 10 10 9 1 11 2
13 11 11 3 3 13 1 9 0 13 9 9 11 2
39 9 10 13 1 9 2 9 15 13 9 2 9 9 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 7 3 3 3 2
17 9 2 9 11 13 1 13 15 0 2 13 9 2 9 15 13 2
9 11 11 13 1 9 1 10 9 2
12 11 11 12 12 12 12 12 2 12 12 12 2
13 9 10 13 11 11 1 11 11 15 3 0 9 2
11 11 13 9 1 11 11 11 11 2 11 2
10 9 10 13 1 12 9 1 12 9 2
26 10 9 15 3 13 1 3 3 1 9 2 7 14 3 13 1 9 11 2 9 10 3 13 11 11 2
18 15 3 13 9 0 1 11 11 1 11 7 11 1 11 11 2 11 2
17 11 13 9 1 11 11 2 11 11 7 11 2 11 11 2 11 2
13 1 9 9 11 2 11 11 13 1 11 11 11 2
12 16 12 9 2 15 13 13 9 15 7 13 2
7 9 7 9 9 2 2 2
23 3 16 2 9 9 9 3 3 13 2 1 9 2 9 2 9 2 9 2 7 13 9 2
15 9 9 11 11 13 9 11 3 13 7 13 9 11 11 2
28 9 9 11 13 11 2 2 2 7 11 11 2 2 11 11 2 11 2 2 2 2 15 3 3 13 3 11 2
26 11 11 11 11 11 11 11 11 11 13 10 9 1 11 15 3 13 9 9 11 1 11 2 11 2 2
40 1 9 9 11 11 2 14 13 11 2 9 2 11 11 7 11 11 13 10 10 9 1 11 11 2 7 13 9 9 9 11 2 11 11 11 2 11 2 11 2
20 1 12 9 13 2 9 11 1 11 11 13 0 16 3 13 2 13 9 2 2
19 9 10 3 13 9 9 9 1 13 1 9 9 1 9 11 1 11 11 2
110 9 13 11 2 11 11 11 11 2 0 1 9 11 11 7 9 0 1 9 0 2 11 11 2 11 13 1 11 9 9 2 9 1 9 9 13 1 9 15 13 1 9 9 2 9 15 13 1 9 9 11 12 1 10 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 9 2 2 11 11 2 11 2 9 2 11 2 11 2 11 2 11 2 2 11 2 11 2 11 2 2 11 11 2 11 2 7 11 2 11 2 11 2 11 2 2
45 9 10 13 11 11 2 15 13 9 11 2 13 10 10 9 9 15 0 1 9 11 11 12 2 11 11 12 13 11 11 1 9 15 3 13 7 3 13 2 16 10 9 9 0 2
17 11 11 13 9 9 1 11 2 2 7 10 10 9 0 1 11 2
11 9 9 9 9 10 13 7 9 9 0 2
25 10 9 9 9 9 1 3 13 13 9 9 9 2 10 9 15 3 13 1 10 9 9 9 9 2
28 11 11 2 13 12 11 12 1 11 2 11 11 2 13 12 11 12 1 11 2 2 13 10 9 0 9 11 2
21 10 9 13 1 12 9 3 0 2 0 0 2 0 2 0 2 9 2 7 0 2
15 1 9 9 9 1 9 11 11 2 9 9 11 3 13 2
12 9 10 13 9 15 13 2 11 11 11 2 2
35 12 9 1 9 12 2 15 13 1 10 9 2 7 1 9 2 9 2 9 15 13 2 1 9 2 13 1 11 11 2 13 1 9 12 2
18 11 9 2 9 0 7 9 2 13 1 9 1 9 12 1 12 9 2
28 1 9 11 1 9 11 1 9 11 2 11 15 0 2 11 3 13 9 1 9 11 15 3 13 1 9 0 2
9 1 9 3 13 7 9 11 11 2
16 7 16 16 9 3 13 2 12 9 0 7 9 1 11 13 2
12 3 9 10 13 9 2 15 14 13 1 9 2
24 1 10 9 15 0 2 1 9 12 5 9 3 13 2 9 14 13 3 3 13 9 9 9 2
13 1 9 10 2 15 13 11 11 11 1 9 12 2
74 11 2 12 11 12 2 11 11 12 2 12 11 11 13 1 11 5 11 11 2 0 9 12 13 9 2 11 11 2 2 9 11 11 7 10 9 0 11 11 2 7 9 1 9 11 7 9 11 11 13 1 11 2 9 13 1 9 11 11 11 2 11 2 11 11 15 13 9 11 1 10 9 0 2
9 3 3 9 11 16 13 9 10 2
60 10 9 2 9 11 9 10 13 11 11 2 15 3 13 9 9 1 2 11 11 2 2 15 13 1 13 9 2 9 15 13 1 9 10 2 13 9 9 15 3 13 9 9 9 10 2 7 13 9 1 10 9 9 9 15 0 2 9 2 2
9 1 12 9 9 13 9 3 13 2
28 9 2 9 0 2 2 11 11 2 7 2 11 11 11 2 13 1 9 12 9 9 11 16 13 1 9 12 2
16 9 11 3 13 0 16 13 1 9 11 2 16 3 13 2 2
9 11 11 11 13 1 12 9 9 2
12 0 0 9 9 0 1 11 2 11 7 11 2
6 9 2 3 9 11 2
9 11 11 9 9 1 11 11 0 2
18 11 13 9 15 13 1 11 11 2 11 11 11 2 11 11 2 11 2
11 11 11 13 11 11 11 13 9 12 11 2
11 9 0 9 13 1 11 2 15 13 9 2
11 1 9 12 11 13 9 11 1 9 12 2
6 2 3 13 14 3 2
13 11 13 9 1 11 11 2 11 2 11 2 11 2
14 16 11 13 1 9 0 2 11 2 11 13 3 11 2
28 11 13 11 11 1 11 1 9 12 2 1 9 13 9 9 9 9 2 15 13 9 1 1 11 13 13 11 2
19 16 2 13 16 9 9 9 13 1 13 9 2 11 2 8 2 5 12 2
8 0 9 9 9 11 7 11 2
9 11 11 2 11 13 9 12 9 2
44 1 11 11 2 11 13 13 11 11 1 11 1 9 1 11 2 13 2 12 2 7 11 2 13 2 12 2 1 13 1 9 9 9 2 3 9 11 1 11 11 1 11 11 2
26 16 16 15 13 13 11 3 2 3 2 3 11 2 11 11 2 15 13 9 11 13 1 13 3 9 2
17 9 9 2 12 12 9 11 2 12 12 9 11 2 12 9 12 2
10 3 11 11 11 0 1 11 11 11 2
22 11 11 13 9 11 1 10 11 13 11 11 1 12 1 9 9 11 2 9 9 2 2
57 9 10 15 13 0 9 1 2 3 9 10 13 9 15 13 7 13 9 9 16 1 12 9 14 13 9 15 13 2 16 11 13 9 1 11 11 2 10 9 0 15 3 13 9 2 7 1 11 11 2 11 13 9 14 3 13 2
33 1 11 11 11 11 2 9 9 10 9 13 12 12 2 7 1 9 10 2 12 2 12 9 13 9 16 12 2 12 9 13 9 2
16 1 9 9 11 2 9 9 13 1 9 9 0 1 9 0 2
49 1 11 2 11 2 11 11 2 7 11 2 3 13 1 10 9 1 13 9 1 9 3 2 9 11 2 9 11 2 11 11 2 7 11 2 9 11 2 11 11 2 1 13 9 9 15 15 13 2
11 15 13 1 11 11 2 11 2 11 11 2
10 11 13 9 1 9 7 9 9 9 2
22 16 13 7 13 1 9 10 11 2 7 13 9 9 2 15 13 1 9 2 2 9 2
13 1 9 11 2 11 13 10 10 9 9 9 9 2
36 11 13 9 1 9 1 11 11 1 9 1 9 1 1 9 11 12 2 2 14 15 13 2 16 15 15 13 9 1 9 13 15 0 7 0 2
24 9 10 13 1 9 12 2 12 1 9 0 1 9 11 2 11 2 11 2 7 9 2 9 2
11 3 0 2 10 9 13 1 0 13 0 2
13 1 9 11 12 2 13 10 9 0 1 11 11 2
29 9 0 1 11 2 13 9 7 2 9 3 13 9 2 7 9 2 9 2 7 9 13 10 9 13 9 7 9 2
13 1 10 3 2 9 11 11 13 1 9 9 0 2
35 1 9 12 2 12 2 2 9 11 13 1 9 9 16 13 9 9 7 3 13 11 2 15 9 3 3 13 1 9 9 2 1 11 11 2
21 9 9 13 9 11 1 10 9 9 13 1 9 11 2 9 11 2 7 9 0 2
16 9 13 9 9 1 9 11 11 1 13 9 9 1 9 10 2
14 11 13 12 1 12 9 7 9 15 13 1 9 11 2
19 16 13 9 9 9 2 9 0 2 1 11 11 2 3 9 10 14 13 2
25 15 13 1 9 1 9 2 7 1 9 1 11 11 1 12 15 13 11 11 11 7 13 1 9 2
21 11 11 2 2 13 10 9 9 9 13 9 15 13 1 9 11 1 9 9 9 2
25 11 11 3 13 16 2 1 9 0 3 13 1 9 2 9 0 2 3 9 7 9 2 2 2 2
12 1 3 2 9 13 9 9 2 13 3 9 2
21 9 9 0 13 3 13 1 9 15 13 1 9 9 12 2 12 7 12 2 12 2
41 1 9 0 2 13 9 13 9 0 2 1 11 7 11 11 11 7 11 11 11 11 2 7 9 9 0 2 1 12 11 2 11 11 11 11 11 11 7 11 11 2
26 11 13 16 9 11 1 11 11 13 1 13 9 9 9 2 11 11 2 13 1 11 1 11 12 2 2
9 1 9 10 9 9 13 9 9 2
14 1 9 15 13 13 11 11 11 15 13 1 11 11 2
35 11 11 11 13 2 9 11 1 9 11 2 11 11 1 11 11 7 11 11 13 9 9 1 9 11 2 11 11 7 9 11 1 9 11 2
20 11 11 13 9 12 9 1 9 11 11 2 11 11 2 11 11 11 2 11 2
11 9 9 1 9 10 13 11 2 11 11 2
30 9 10 13 16 1 13 9 9 3 3 13 9 9 2 1 9 10 16 13 13 1 9 9 3 13 1 9 15 0 2
72 9 10 13 1 9 11 11 1 11 11 2 1 9 1 12 2 9 10 13 13 12 9 2 11 11 2 11 11 2 7 11 11 2 11 11 2 15 13 1 9 1 11 11 7 9 11 2 9 9 0 11 2 15 13 1 11 2 11 11 2 10 9 2 15 13 1 9 11 2 9 11 2
15 14 2 15 13 3 14 2 2 13 2 15 13 3 14 2
8 9 10 13 9 1 12 9 2
8 11 9 10 13 1 9 12 2
17 13 9 9 12 2 9 11 1 13 3 13 3 0 1 13 9 2
11 11 11 13 10 9 1 9 9 11 11 2
48 13 11 1 11 10 2 2 16 3 9 2 3 9 13 9 10 2 15 14 3 13 2 14 3 13 7 14 3 13 2 14 3 13 9 7 13 9 2 16 14 3 13 15 1 9 7 9 2
69 1 12 9 7 12 9 2 9 9 1 3 13 1 9 9 11 2 7 3 3 15 13 1 9 11 1 9 10 2 15 3 9 3 3 13 1 9 0 2 1 9 9 1 2 12 11 2 11 3 13 9 9 11 1 9 9 11 1 11 2 9 2 9 12 2 12 9 2 2
13 11 11 9 1 2 11 11 15 13 1 11 2 2
21 11 13 9 9 15 13 16 9 9 9 2 9 10 13 1 9 0 7 9 9 2
12 11 13 9 15 13 1 9 11 11 2 11 2
9 1 12 9 3 13 13 0 11 2
33 11 13 9 0 1 3 13 1 1 12 9 0 2 9 11 7 9 11 5 11 1 13 9 1 12 9 9 9 9 12 9 10 2
8 9 9 10 0 1 9 11 2
34 11 1 9 9 7 9 13 9 0 1 11 15 13 1 9 1 0 12 11 2 11 13 9 0 1 12 9 9 3 0 1 11 11 2
18 9 9 0 1 9 10 13 9 2 9 2 9 2 9 2 9 9 2
20 9 9 9 10 13 1 10 9 11 2 11 11 2 15 3 13 9 9 10 2
16 11 13 10 9 1 11 11 2 11 11 2 11 11 2 11 2
41 1 9 10 9 15 13 2 11 2 13 1 9 9 9 9 9 2 11 11 2 2 9 10 13 13 12 9 9 13 1 9 9 1 10 9 9 11 2 9 2 2
46 1 9 11 11 2 1 9 9 3 13 16 9 9 2 9 9 11 13 9 9 0 7 9 2 9 2 9 7 9 0 1 9 2 9 9 0 2 7 9 2 9 0 1 9 9 2
35 10 9 16 9 0 13 9 1 13 0 7 0 1 9 2 1 9 15 7 9 15 2 1 10 10 9 0 1 9 9 2 9 7 9 2
3 2 9 2
20 11 3 3 13 9 1 0 16 15 13 1 9 2 9 9 2 7 9 9 2
35 1 11 3 13 10 9 15 0 7 3 13 2 1 0 11 11 11 2 11 2 11 11 11 2 11 11 7 3 13 9 9 1 11 0 2
42 1 13 1 9 1 10 2 1 9 13 1 13 2 16 9 13 15 3 3 13 9 13 15 3 13 9 7 13 9 9 9 2 1 2 1 7 9 2 1 2 9 2
19 16 9 9 9 0 1 9 0 1 0 13 9 9 9 2 12 11 11 2
19 9 11 13 1 11 16 1 9 10 2 11 11 3 13 1 9 9 11 2
22 9 9 0 15 13 1 11 13 9 0 2 9 2 9 2 0 2 7 9 9 0 2
32 11 9 0 2 11 11 2 3 0 1 9 7 15 0 13 9 9 9 9 2 11 2 11 11 2 7 11 2 11 11 2 2
11 11 13 9 15 13 1 11 11 2 11 2
9 3 11 14 3 13 1 11 10 2
11 9 12 1 13 9 1 9 9 5 9 2
12 9 11 12 13 2 11 11 2 11 11 2 2
27 11 9 0 11 2 11 11 11 11 11 2 3 13 1 11 2 13 10 9 9 0 1 9 11 11 0 2
23 11 10 13 1 9 11 11 10 3 13 1 11 11 2 11 11 7 9 2 9 11 0 2
61 9 15 3 13 1 11 7 9 2 9 13 9 11 15 3 13 0 9 2 9 12 9 1 12 9 2 1 9 0 1 2 15 13 1 9 13 9 2 2 7 2 1 9 15 13 9 0 2 2 2 1 10 10 2 15 13 9 0 15 0 2
34 16 9 13 11 1 9 1 9 11 12 2 9 10 13 2 13 10 9 0 2 2 16 13 9 2 9 3 15 13 1 9 12 9 2
33 11 11 13 1 9 15 3 0 16 10 15 13 1 1 3 15 13 9 1 9 9 9 7 1 9 1 0 2 0 7 1 9 2
14 15 3 13 1 11 11 1 11 2 11 2 7 11 2
13 16 9 10 13 1 0 15 2 14 15 13 9 2
13 3 0 9 13 9 7 7 3 13 9 7 9 2
8 0 9 1 9 9 11 11 2
49 11 9 1 11 11 13 9 9 2 9 3 2 9 13 7 13 1 9 9 9 2 9 9 7 11 13 1 9 9 9 9 2 16 15 0 3 13 1 9 9 2 9 0 13 1 9 9 0 2
24 11 1 9 9 1 9 11 11 7 9 2 13 10 10 9 1 11 7 9 15 14 13 9 2
18 11 13 2 16 15 14 3 13 9 10 2 3 9 2 11 2 13 2
7 10 13 9 9 0 11 2
9 9 9 9 11 13 9 15 0 2
32 11 13 0 16 14 13 0 2 0 16 10 9 9 9 11 11 1 11 11 3 13 1 11 11 15 13 9 1 9 13 11 2
24 11 12 13 1 13 9 9 1 11 11 2 13 9 9 1 9 11 2 12 9 1 1 9 2
6 9 15 3 13 0 2
11 11 9 13 9 0 1 9 15 13 0 2
15 9 13 1 9 12 5 12 2 11 12 5 12 2 11 2
5 5 15 3 10 2
18 9 9 13 13 11 11 11 9 13 10 9 15 9 13 1 11 11 2
37 10 13 9 2 11 11 2 11 2 11 11 2 1 3 11 2 11 11 2 11 2 11 2 7 11 9 0 2 7 10 9 13 9 9 9 11 2
14 15 3 13 1 11 11 16 11 11 13 1 9 12 2
12 11 13 9 1 11 11 7 3 13 9 0 2
12 10 10 1 15 13 1 11 2 9 15 0 2
38 1 9 9 9 9 2 9 9 0 1 9 15 13 13 3 13 2 1 15 13 9 13 9 9 7 9 9 9 1 9 9 2 9 2 7 10 9 2
21 16 9 11 3 3 13 9 9 11 2 15 9 13 0 11 14 13 9 9 0 2
7 13 15 1 9 7 9 2
12 11 9 13 3 1 0 1 11 11 11 11 2
11 11 14 13 2 16 11 10 9 7 3 2
16 3 1 13 9 15 12 9 3 13 3 9 9 13 1 9 2
11 11 13 9 9 11 11 2 11 11 11 2
40 9 10 3 13 1 2 9 0 1 9 9 15 13 1 11 1 9 9 12 11 12 7 12 11 12 2 7 3 13 1 9 9 9 1 12 9 1 9 12 2
14 9 0 13 1 9 9 2 16 9 9 13 1 9 2
20 1 10 9 9 0 2 11 13 9 1 9 2 2 9 15 13 9 9 9 2
76 1 9 9 9 11 11 11 9 2 12 5 9 5 9 5 12 5 12 9 12 9 12 2 13 9 9 9 2 1 9 11 2 11 2 11 11 7 13 1 9 2 11 11 2 9 2 11 11 11 2 9 2 2 9 2 11 2 11 11 2 9 2 11 2 9 2 11 7 11 11 2 11 2 9 2 2
21 11 11 11 11 11 13 11 11 0 15 13 1 11 2 11 11 11 2 12 11 2
22 11 11 13 10 10 9 15 13 1 9 11 11 2 11 11 11 2 11 11 2 11 2
14 11 11 11 13 9 15 13 1 9 11 11 2 11 2
16 9 3 13 9 9 16 13 11 2 9 9 2 1 9 12 2
14 15 13 9 3 2 3 13 9 0 7 0 1 9 2
25 3 3 0 16 9 10 3 13 9 11 15 13 2 16 9 10 11 13 1 9 11 11 15 13 2
7 9 13 0 7 0 0 2
9 11 11 3 13 3 7 1 0 2
4 9 9 13 2
26 9 10 3 9 10 9 9 0 1 2 9 9 2 9 0 1 9 11 11 2 7 9 0 11 11 2
60 13 9 9 9 10 15 13 1 11 11 15 0 2 13 9 1 13 11 11 2 1 9 9 1 9 2 15 13 9 1 11 2 11 2 9 9 11 2 11 2 1 9 1 13 11 11 2 15 13 9 9 1 0 7 13 9 2 9 0 2
29 1 9 11 2 1 9 12 2 12 2 11 13 9 1 13 9 1 9 11 11 11 2 11 1 9 1 9 11 2
71 11 11 11 13 1 9 12 11 1 9 12 11 12 1 11 11 11 2 12 9 3 13 1 11 1 9 0 13 11 11 11 2 9 0 0 15 13 1 9 10 2 11 2 13 1 12 9 2 9 16 13 9 9 1 9 12 2 12 2 9 9 2 1 9 11 2 12 2 11 12 2
12 15 15 13 15 1 9 11 15 3 0 10 2
16 15 9 10 11 11 11 13 2 14 1 15 13 3 9 2 2
9 1 9 12 2 11 3 13 9 2
25 9 9 7 9 1 9 11 13 9 11 1 9 0 1 9 15 13 13 2 7 3 1 9 9 2
31 16 15 3 15 13 1 9 0 1 1 9 13 3 2 16 16 13 1 9 9 15 0 1 9 2 0 7 0 2 0 2
16 15 13 9 12 7 13 2 11 2 2 16 15 13 1 11 2
15 11 9 13 9 9 15 13 1 11 11 2 11 2 11 2
19 11 9 3 13 1 10 9 7 9 1 11 1 9 1 9 0 7 9 2
13 11 13 1 9 9 1 11 1 11 2 11 2 2
22 11 11 13 10 9 9 0 2 1 9 1 12 9 2 11 2 9 0 7 9 0 2
14 1 12 9 1 12 2 12 9 0 13 1 9 0 2
8 10 13 9 15 0 13 9 2
24 11 5 9 2 15 13 1 9 0 13 9 0 15 3 0 2 3 9 0 15 13 2 13 2
13 11 11 3 13 9 9 10 9 15 13 9 10 2
12 11 11 3 13 13 9 9 1 1 9 11 2
23 10 9 1 11 11 7 11 11 15 13 13 9 7 3 3 3 9 9 9 1 13 9 2
23 11 9 10 13 1 13 9 2 9 11 2 11 11 11 15 3 13 13 11 13 11 11 2
8 11 10 13 9 0 1 11 2
24 9 10 13 1 13 12 9 9 11 2 9 2 9 7 9 2 1 9 9 9 9 1 11 2
20 1 9 11 13 1 10 9 9 11 15 0 13 9 2 9 7 9 1 13 2
12 7 3 13 11 11 7 11 11 7 11 11 2
10 9 13 11 15 13 1 9 2 11 2
9 11 10 3 13 1 11 7 11 2
7 1 9 15 13 13 9 2
8 11 11 13 10 9 1 11 2
9 9 11 11 11 13 1 2 11 0
23 9 11 13 1 9 12 7 12 3 13 1 11 11 1 13 9 11 12 15 13 9 9 2
11 16 9 0 13 12 9 9 0 15 13 2
14 11 13 9 1 11 11 2 11 11 2 11 2 11 2
7 1 9 9 13 10 9 2
11 9 13 2 15 13 1 9 7 1 9 2
46 11 11 11 11 11 11 13 11 11 11 15 13 9 12 1 11 2 11 13 3 3 13 1 9 9 12 2 12 2 16 13 1 11 11 7 11 11 13 1 11 1 11 2 11 11 2
10 9 2 9 9 10 14 13 1 0 2
26 10 9 13 9 11 13 3 1 11 2 16 15 0 3 13 1 11 2 9 11 3 13 1 11 2 2
40 9 15 13 9 1 9 11 2 11 11 11 10 3 13 1 12 9 2 13 1 12 9 7 12 9 2 9 9 9 0 1 9 1 3 3 3 13 1 15 2
21 9 13 1 9 12 2 15 13 9 3 13 1 1 9 11 7 13 13 12 5 2
30 16 9 10 7 9 9 1 11 11 2 11 13 9 9 13 11 2 7 16 11 11 3 13 9 0 1 9 2 9 2
19 2 15 13 15 15 15 13 13 1 9 10 2 7 10 14 9 15 13 2
12 9 10 13 1 11 11 7 13 1 9 0 2
20 11 11 13 9 1 11 11 11 2 11 11 2 11 11 11 2 11 2 11 2
48 9 0 13 1 13 9 9 1 9 9 1 9 9 9 2 9 9 9 2 9 9 7 9 9 2 9 0 1 13 9 13 9 15 3 0 2 0 7 9 2 15 13 9 0 7 11 11 2
16 13 9 9 1 13 11 1 11 1 9 9 15 3 13 9 2
50 11 13 9 1 11 15 13 1 11 12 1 9 11 2 11 2 2 11 2 9 2 2 11 2 9 2 2 11 2 11 2 2 11 2 11 2 2 7 11 2 9 2 2 9 9 10 13 9 9 2
24 11 11 2 2 13 10 9 9 9 13 9 15 13 1 9 11 11 11 3 13 1 9 9 2
57 1 9 11 2 9 10 13 1 9 11 15 16 15 3 13 1 9 1 9 11 12 1 9 15 1 11 2 11 11 2 7 11 11 11 2 1 9 12 11 9 10 13 1 9 11 7 9 9 16 15 3 13 9 1 11 11 2
68 11 11 12 5 12 13 12 9 0 9 9 15 13 2 3 2 3 2 11 9 12 5 12 3 0 13 9 9 9 1 1 2 9 9 11 9 12 9 12 3 3 13 2 11 9 12 5 12 2 7 3 11 11 11 5 11 2 14 13 9 3 1 9 7 9 9 9 2
86 1 9 0 2 9 0 1 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 13 1 9 0 2 16 11 11 13 9 12 2 12 11 11 1 9 12 2 12 2 12 2 12 7 9 1 11 11 2 11 11 13 9 1 11 2 11 11 1 9 12 2 12 2 12 2 12 2 12 2 12 2
14 9 10 13 9 12 7 13 9 1 11 11 11 12 2
26 7 16 9 11 13 9 11 2 11 13 10 9 0 15 13 1 11 11 1 13 9 0 1 9 9 2
12 1 9 13 3 9 2 9 0 7 9 9 2
21 11 1 1 13 9 9 1 9 2 3 1 13 9 9 1 9 13 9 9 13 2
20 11 9 2 9 2 9 2 11 2 2 11 11 2 13 9 7 9 15 0 2
43 9 9 13 15 13 3 13 9 11 1 9 11 2 7 13 11 11 1 9 2 11 15 3 2 3 0 7 3 13 1 9 0 16 14 13 9 11 11 7 9 9 9 2
20 1 9 12 2 1 9 9 11 1 11 11 2 9 11 11 3 13 12 9 2
11 16 16 9 13 11 2 15 3 13 3 2
7 9 15 15 13 1 11 2
19 11 13 10 10 9 1 9 9 9 2 9 11 2 11 11 11 2 11 2
7 2 3 15 13 9 11 2
28 2 12 12 11 12 12 2 11 2 16 15 13 7 13 1 9 9 7 9 2 9 3 13 9 15 13 0 2
27 11 3 13 13 0 1 9 9 7 9 2 9 0 15 0 1 9 2 7 13 1 9 9 1 9 9 2
38 11 2 11 2 9 2 11 2 11 2 13 10 9 15 13 10 9 1 9 13 2 13 2 9 9 7 3 13 1 9 1 13 9 9 15 3 13 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
24 9 10 3 13 1 11 7 11 2 16 3 15 10 13 11 7 11 1 13 11 2 11 2 2
12 9 11 3 13 12 2 12 9 7 9 0 2
11 11 9 15 13 9 2 9 9 13 9 2
43 0 1 11 1 9 1 11 9 9 9 1 11 11 11 11 13 1 9 12 9 9 2 13 1 11 11 1 11 12 2 10 9 13 11 11 11 11 1 13 9 13 13 2
6 11 11 13 9 0 2
21 11 11 13 9 9 9 1 9 11 11 2 9 11 11 2 11 11 11 2 11 2
43 9 12 9 2 12 2 10 9 1 11 11 13 1 9 12 9 2 9 11 11 13 9 9 1 12 9 9 2 1 9 12 9 7 12 9 2 1 9 1 11 11 11 2
33 1 9 12 2 10 9 9 9 9 11 3 13 9 1 0 7 3 13 9 9 10 15 9 3 3 13 1 9 9 15 13 0 2
14 16 10 2 11 11 11 11 3 13 9 1 9 10 2
9 1 9 2 15 13 9 11 11 2
14 7 11 13 2 2 13 9 0 9 2 11 1 11 2
23 9 9 0 2 11 11 11 2 11 2 2 13 10 10 9 9 15 3 13 1 11 11 2
8 11 1 13 9 1 1 9 2
41 1 9 15 13 2 11 11 11 1 11 12 2 12 2 15 13 9 11 12 15 13 9 11 2 9 2 1 9 9 2 11 11 13 9 1 9 11 1 9 12 2
28 9 15 13 1 11 14 9 0 9 2 1 9 9 9 1 9 9 2 9 0 7 9 2 15 0 2 0 2
18 11 13 10 10 9 1 11 11 11 2 11 11 2 11 11 2 11 2
14 1 9 9 0 2 9 1 9 9 13 1 13 9 2
16 10 11 7 11 13 1 15 12 9 1 13 11 1 9 10 2
15 11 11 13 9 1 9 11 2 11 2 11 11 2 11 2
16 9 13 9 1 11 11 2 11 2 9 0 1 9 2 11 2
16 1 12 1 12 15 13 1 13 9 13 9 15 13 1 12 2
42 9 0 11 1 11 11 1 11 11 13 1 9 0 1 10 9 9 2 3 13 9 9 1 11 11 1 9 12 11 12 15 15 11 11 13 9 9 1 11 1 11 2
10 1 9 9 11 13 7 13 1 11 2
41 15 13 16 13 10 9 1 9 11 2 11 2 1 9 12 11 12 1 11 2 11 2 11 7 13 1 11 11 1 11 2 11 2 15 13 1 0 1 9 12 2
18 1 9 0 2 11 13 13 9 3 3 0 1 9 1 11 11 11 2
13 9 10 13 1 9 9 11 2 9 11 11 11 2
19 3 2 0 9 3 13 1 0 9 7 13 0 7 1 9 15 3 0 2
7 11 9 9 13 11 11 2
17 11 9 10 3 13 9 9 2 9 9 2 7 11 2 11 11 2
9 11 13 1 9 9 11 2 11 2
13 3 2 1 13 9 2 9 13 13 1 9 10 2
16 9 9 7 11 11 13 10 10 9 15 13 1 9 9 13 2
18 11 13 10 9 9 1 9 11 2 11 11 2 11 11 11 2 11 2
19 15 13 3 13 1 9 11 15 3 13 1 9 1 9 15 13 9 9 2
6 9 9 9 1 11 2
25 11 11 13 1 9 9 9 2 11 2 9 1 11 11 11 2 11 11 2 11 11 2 11 11 2
17 9 9 3 0 2 16 13 2 10 9 3 9 2 9 13 9 2
17 9 0 1 9 1 9 15 13 1 9 0 7 0 1 9 11 2
12 11 11 3 13 9 2 9 2 7 9 9 2
5 9 9 10 10 2
9 9 15 13 13 9 1 9 0 2
14 11 11 13 10 9 1 11 11 11 2 11 2 11 2
18 9 10 13 9 9 7 9 15 13 9 12 7 13 0 1 9 12 2
17 9 0 11 13 1 12 2 12 2 7 13 9 3 1 12 9 2
49 9 2 9 0 15 13 1 13 11 11 7 11 11 7 9 2 9 9 2 15 15 13 1 11 11 2 11 2 11 11 11 2 13 1 9 0 2 0 9 9 2 1 12 5 1 9 11 11 2
47 11 13 1 9 9 14 13 11 11 12 7 11 11 12 2 10 9 13 9 15 0 2 15 13 14 13 9 15 3 0 2 9 10 3 13 9 9 15 13 9 3 13 1 9 1 9 2
10 9 10 11 13 11 11 1 9 12 2
19 1 10 9 11 1 11 15 13 9 2 11 2 13 1 9 11 11 11 2
14 10 9 13 1 13 9 10 9 15 13 13 9 0 2
19 9 9 10 13 12 9 3 11 11 11 2 11 11 11 7 11 11 11 2
17 11 1 9 9 14 3 13 9 2 16 9 0 14 3 13 9 2
13 9 0 13 10 0 9 15 1 9 2 9 15 2
26 11 11 9 11 11 1 3 1 12 9 7 3 3 13 9 9 1 11 11 11 11 1 15 11 12 2
36 11 2 11 12 2 12 2 12 2 12 2 13 16 9 2 9 10 13 1 9 11 11 1 11 2 1 15 13 1 9 9 2 15 0 2 2
12 9 10 13 9 9 13 9 0 11 11 12 2
27 11 9 9 10 13 13 7 3 13 9 9 7 9 1 9 13 9 9 1 9 9 9 1 9 9 9 2
18 9 3 13 9 16 11 14 3 3 13 1 10 10 9 1 13 9 2
28 9 15 13 1 11 11 13 1 9 9 1 9 9 1 13 15 15 15 13 1 9 9 11 15 0 1 9 2
17 3 1 3 2 15 3 3 13 9 0 1 15 13 11 1 10 2
23 11 11 11 2 2 13 10 9 9 9 13 11 15 13 1 9 11 11 1 9 9 9 2
23 3 10 2 1 9 12 11 11 2 0 1 13 9 15 0 7 13 9 2 9 15 0 2
17 9 9 9 13 9 16 9 7 9 7 9 13 9 2 9 0 2
46 9 9 15 13 1 9 10 1 0 2 9 9 2 9 9 2 9 2 9 2 3 11 2 11 11 11 2 2 2 9 10 13 9 9 0 1 9 10 16 9 15 13 13 9 0 2
36 9 9 9 9 3 3 1 9 12 11 12 1 8 13 9 2 11 2 11 11 11 11 11 2 2 13 0 1 11 2 11 11 2 11 2 2
5 15 13 1 9 2
10 12 12 9 9 2 9 9 2 9 2
10 11 13 1 11 2 9 0 11 9 2
20 11 2 2 13 10 9 0 2 9 9 2 1 9 11 2 9 9 11 11 2
42 11 11 3 13 10 9 0 1 9 1 9 9 1 9 11 11 2 11 11 11 2 11 11 11 2 7 3 13 11 11 11 1 0 1 11 11 11 11 2 11 2 2
30 1 9 9 12 9 2 9 9 10 3 13 9 1 12 9 1 9 9 2 9 0 2 7 9 15 13 1 10 11 2
7 9 10 13 9 9 12 2
9 3 11 13 3 0 1 9 11 2
45 9 9 15 3 3 13 1 0 2 11 2 11 11 2 2 11 2 11 2 11 2 11 2 11 2 11 11 11 11 7 11 2 11 11 2 7 13 9 1 13 9 2 11 2 2
30 3 13 1 1 9 2 9 11 11 15 13 1 9 2 13 10 9 0 15 13 1 9 1 10 9 2 10 9 0 2
26 1 1 9 10 2 9 13 10 9 1 13 10 9 15 3 13 1 9 9 7 1 13 9 1 9 2
37 16 13 15 1 9 9 2 16 9 13 2 3 13 9 2 9 7 9 2 9 10 1 9 9 11 2 15 13 9 9 9 9 10 2 7 13 2
16 16 3 13 2 7 11 14 3 13 11 11 3 13 13 9 2
4 3 15 13 2
26 1 9 15 12 2 13 9 10 9 2 2 3 3 15 13 2 15 13 9 2 3 9 14 13 9 2
17 3 11 3 13 0 9 1 9 9 14 15 13 13 13 1 9 2
36 16 11 9 11 13 9 2 9 11 3 13 9 2 9 13 9 9 1 9 9 15 0 2 9 13 1 9 9 2 16 9 13 1 9 9 2
41 1 9 13 9 2 11 11 2 15 13 9 1 9 11 11 2 7 1 9 13 9 11 11 2 7 11 11 11 2 15 13 9 2 9 0 1 9 9 10 9 2
16 9 3 13 0 1 9 9 7 13 2 13 13 9 9 9 2
9 9 3 13 10 9 9 9 0 2
88 1 9 0 1 9 0 9 15 13 9 9 1 9 11 13 9 9 3 0 1 9 11 13 9 2 9 2 9 2 9 2 9 2 9 2 7 9 2 7 9 3 13 9 2 16 10 9 13 9 9 0 1 9 15 3 13 1 9 2 9 2 9 2 9 2 7 3 0 9 9 9 3 13 9 1 9 7 13 1 9 9 9 16 9 15 13 0 2
42 11 11 11 11 13 10 9 9 9 0 15 13 1 9 9 1 10 9 2 1 3 1 12 9 13 1 11 11 2 11 15 13 1 0 1 9 9 2 13 7 13 2
23 1 9 12 9 9 13 9 9 9 1 9 9 12 1 12 9 1 12 9 1 9 12 2
15 11 11 13 9 1 11 12 15 13 1 11 7 13 11 2
26 9 10 13 9 12 1 9 11 7 9 1 9 1 9 9 10 9 7 9 15 13 9 11 2 11 2
28 9 11 11 2 1 9 1 11 11 2 13 0 1 9 9 9 0 11 15 15 13 7 9 0 15 15 13 2
20 1 11 11 2 10 9 11 11 0 10 13 1 11 5 11 7 11 11 11 2
47 1 9 10 11 11 9 9 9 0 7 2 9 9 2 2 10 11 11 1 9 0 1 11 3 13 9 9 11 10 16 9 3 0 2 3 12 2 12 5 1 9 9 15 13 1 9 2
4 15 13 11 2
19 1 9 10 11 11 13 9 9 11 11 11 2 7 13 9 13 11 11 2
43 11 11 2 11 11 11 2 9 13 7 15 13 1 11 2 13 11 2 9 11 11 2 16 15 13 9 1 11 11 2 9 9 0 2 16 13 9 1 10 9 7 9 2
25 15 13 9 9 1 11 11 11 1 9 11 11 1 9 12 11 12 1 9 1 11 11 11 11 2
39 1 9 11 2 9 9 16 9 2 9 2 2 3 13 1 9 2 9 1 11 1 11 1 13 10 9 2 1 9 11 2 9 11 2 7 0 2 0 2
28 9 9 9 13 1 9 9 1 9 7 9 15 13 2 16 9 9 0 0 7 0 1 9 0 13 3 0 2
16 11 11 16 13 13 1 11 11 11 2 11 11 2 11 11 2
16 11 1 9 12 1 11 13 3 1 9 11 13 1 9 12 2
13 11 11 13 2 2 16 15 14 13 9 2 2 2
13 9 11 11 13 10 10 9 1 11 11 2 11 2
11 11 11 2 2 13 10 9 7 9 11 2
19 11 11 13 9 12 12 2 12 9 2 7 9 12 5 2 12 9 2 2
49 11 13 3 2 1 9 11 0 2 1 9 13 1 0 2 9 9 2 9 13 7 9 2 9 15 0 13 1 11 11 2 9 9 11 15 13 2 9 9 1 13 7 9 2 1 9 9 9 2
21 11 11 3 13 1 0 7 1 0 1 13 9 9 9 15 3 13 1 1 9 2
32 11 2 9 9 7 9 0 3 13 0 2 16 9 9 2 9 9 2 9 9 2 9 0 2 11 2 11 11 2 7 9 2
19 11 11 13 9 0 15 13 1 9 11 11 7 11 11 11 1 11 11 2
12 9 9 10 13 1 12 9 2 9 7 11 2
16 1 9 12 2 9 10 13 9 1 12 9 7 12 9 9 2
32 9 1 9 10 13 11 1 13 10 9 13 2 1 2 11 11 2 2 2 11 11 2 2 2 11 11 2 7 2 11 2 2
29 11 11 11 2 2 2 2 2 2 13 10 9 0 1 11 11 2 15 13 10 10 9 11 2 12 11 2 0 2
48 11 0 2 11 11 13 9 15 13 11 11 13 3 0 1 9 2 9 15 13 2 1 9 9 9 0 2 11 11 7 9 9 1 9 1 9 9 11 2 7 1 10 9 2 1 9 9 2
14 9 9 3 0 1 9 9 9 9 7 9 9 9 2
33 10 9 13 13 9 0 1 11 1 9 12 7 12 13 1 10 9 1 11 11 11 1 11 12 2 11 11 11 2 2 12 2 2
37 10 9 0 3 13 9 7 13 1 9 13 9 9 0 10 2 13 16 10 9 3 3 13 1 9 9 0 1 12 9 7 13 1 9 10 9 2
42 11 15 13 3 13 16 9 10 13 1 9 9 9 9 9 9 11 9 9 11 12 13 1 11 11 11 2 15 13 1 9 2 9 9 2 2 11 2 11 11 2 2
24 11 0 11 10 13 9 13 9 9 15 3 0 1 9 9 2 9 9 9 10 2 13 0 2
13 15 13 13 1 9 0 2 11 1 12 11 12 2
5 7 15 15 13 2
26 1 9 12 2 11 2 11 2 13 9 15 13 2 11 2 1 9 9 2 11 2 11 2 11 2 2
16 11 11 11 11 11 2 11 11 2 13 9 0 12 1 11 2
21 11 13 16 11 13 9 0 1 13 9 9 7 13 10 15 13 1 9 15 0 2
35 1 11 7 11 15 13 9 0 16 9 9 2 9 15 0 10 13 1 0 1 9 0 1 9 0 2 13 1 9 0 1 10 9 9 2
8 11 3 3 13 1 9 11 2
6 15 13 1 9 9 2
15 11 2 11 3 13 9 10 13 9 9 1 11 2 11 2
3 13 9 2
25 15 13 9 13 1 9 9 9 7 9 0 0 1 10 9 3 3 3 13 9 9 15 3 13 2
24 1 16 10 2 9 13 11 1 13 9 0 2 16 3 13 1 9 13 0 1 9 9 11 2
11 11 9 2 13 10 9 1 11 11 11 2
38 3 1 9 2 9 9 11 2 1 9 15 13 3 13 1 9 9 1 11 11 1 9 10 9 12 5 1 1 9 11 9 9 1 11 11 13 12 2
9 1 10 11 13 1 11 11 11 2
51 9 2 9 1 11 11 15 13 11 13 1 11 11 1 12 11 13 11 11 11 2 11 11 11 2 3 13 1 9 9 9 9 9 11 1 12 11 2 9 9 1 9 11 11 13 1 11 1 12 11 2
11 9 1 9 10 3 13 9 9 7 9 2
17 11 11 13 9 11 7 9 9 3 13 1 9 9 9 11 0 2
38 11 11 11 2 12 2 13 10 9 9 9 0 9 9 9 11 11 11 9 11 2 11 10 13 15 12 1 0 16 9 9 10 13 9 9 11 11 2
10 7 2 3 11 3 13 15 3 3 2
17 11 13 10 10 9 1 11 11 2 11 11 2 11 11 2 11 2
7 9 12 5 1 9 9 2
10 11 9 10 13 1 11 11 11 11 2
29 1 0 9 2 11 13 9 9 0 15 3 13 2 13 2 7 13 9 9 9 0 7 1 0 13 1 9 9 2
40 3 3 9 15 13 11 2 16 11 13 3 13 9 1 9 2 16 9 3 13 16 11 13 3 11 3 3 13 11 2 10 9 13 9 2 11 7 11 13 2
14 9 0 15 13 9 0 1 9 10 13 11 11 11 2
12 11 11 13 9 15 13 1 9 1 12 9 2
21 11 13 9 1 9 1 12 9 9 9 9 12 12 9 10 9 1 9 13 9 2
16 15 0 11 9 0 3 13 9 11 2 15 13 9 9 0 2
57 1 12 11 12 2 16 13 1 9 9 13 11 11 2 9 13 10 9 1 9 0 1 9 13 11 1 9 12 9 11 11 11 2 11 10 13 9 13 1 9 0 12 2 12 7 13 11 1 9 9 1 9 0 12 2 12 2
12 11 13 9 1 9 11 11 2 15 13 9 2
29 16 0 2 3 13 3 16 11 13 9 11 11 12 15 13 1 9 0 2 9 0 13 11 11 1 9 12 2 2
26 16 9 9 10 3 13 10 9 1 11 11 2 10 9 3 3 13 1 0 1 9 0 10 3 13 2
41 16 11 11 13 16 9 13 14 13 9 9 1 13 9 11 2 16 1 9 12 3 10 9 1 13 1 9 2 9 13 11 11 11 11 2 11 2 9 1 11 2
34 11 2 7 3 13 9 2 7 11 2 13 9 1 9 11 11 15 13 9 1 9 9 9 2 15 3 13 3 1 9 12 1 12 2
5 9 1 9 15 2
30 0 1 11 1 9 1 11 9 9 9 1 11 11 11 11 13 1 9 12 9 9 2 13 1 11 11 1 11 12 2
11 11 13 9 9 13 1 12 2 12 9 2
26 10 9 0 13 9 1 13 9 13 7 9 2 13 9 2 2 16 10 14 13 9 9 1 9 10 2
14 1 12 15 13 13 1 11 11 1 13 11 11 9 2
31 9 11 2 7 11 2 13 13 1 9 11 2 9 15 13 1 9 11 0 1 9 11 15 13 1 9 9 9 11 11 2
20 15 13 9 9 9 11 11 2 13 1 11 11 15 13 9 1 9 11 11 2
18 9 15 0 16 9 15 13 13 9 0 2 16 13 9 1 9 10 2
20 10 9 0 13 0 1 9 1 9 7 9 2 9 13 1 9 2 9 0 2
19 1 9 9 13 9 2 9 15 0 7 0 2 7 9 11 1 11 13 2
25 7 10 13 3 1 9 9 13 1 13 11 1 13 1 11 11 2 10 9 13 1 11 2 11 2
13 9 9 15 13 9 13 9 9 16 9 13 0 2
9 9 12 9 15 13 9 1 9 2
35 1 9 9 1 9 9 2 9 2 9 15 9 1 11 11 13 13 12 9 9 2 9 10 13 9 9 2 9 0 7 9 1 10 9 2
34 1 9 9 11 2 9 1 11 3 12 9 12 2 11 7 12 9 12 2 11 2 12 9 13 1 9 9 0 7 9 2 9 9 2
32 1 9 9 9 7 9 9 2 14 13 0 10 13 9 15 3 0 7 1 9 0 3 2 13 7 13 15 1 9 10 9 2
31 1 0 9 12 2 12 2 11 3 13 13 11 15 13 1 9 11 2 1 9 12 2 11 11 13 1 9 2 9 11 2
8 11 7 11 3 3 13 11 2
13 11 9 1 11 13 12 2 9 9 7 9 9 2
26 16 9 3 13 11 2 3 13 1 5 9 2 5 9 2 5 9 2 5 12 2 7 3 0 3 2
16 11 10 13 9 9 0 15 3 0 16 9 3 13 1 0 2
49 9 12 9 0 3 13 2 16 11 11 15 13 12 9 7 11 11 15 13 9 2 16 3 13 1 12 9 9 7 10 9 9 0 2 13 11 2 11 11 1 10 9 9 15 13 1 9 11 2
23 3 9 0 13 9 0 13 9 0 2 9 13 9 0 1 9 9 15 13 9 9 0 2
11 11 11 13 9 1 9 13 10 9 0 2
17 9 13 10 9 9 1 9 11 11 2 11 11 2 11 11 11 2
29 9 0 15 13 3 13 9 2 9 15 14 3 13 0 1 11 2 11 2 1 9 11 2 11 7 9 0 0 2
27 11 11 11 11 11 11 11 3 13 9 0 9 9 9 2 11 2 1 13 9 9 1 9 10 2 10 2
16 11 11 13 9 9 9 9 0 15 13 1 9 9 9 0 2
24 13 10 10 9 15 3 13 7 10 0 3 13 9 9 9 2 1 9 13 1 13 9 10 2
30 11 9 3 13 1 11 11 7 9 3 13 1 11 11 2 1 1 11 2 12 2 11 2 12 3 3 13 1 11 2
11 11 11 2 2 13 10 9 9 1 11 2
7 3 11 3 13 1 9 2
14 9 13 9 9 2 9 2 7 9 0 2 9 2 2
21 9 3 0 2 13 1 12 9 15 3 0 2 3 12 9 2 9 2 1 9 2
15 11 11 2 11 2 13 9 9 9 15 13 1 11 11 2
46 3 13 13 9 11 11 2 16 9 9 13 9 1 9 12 11 12 2 9 10 14 13 9 16 9 10 13 9 15 0 2 7 13 2 9 0 2 15 13 1 11 11 7 11 11 2
9 9 15 3 13 1 11 7 11 2
6 11 11 13 1 11 2
18 1 9 3 2 9 7 9 9 13 1 11 2 7 11 13 9 9 2
4 3 15 13 2
4 9 13 9 2
14 16 13 11 1 15 2 2 14 11 15 13 9 9 2
22 11 9 3 13 1 12 9 7 13 1 9 0 12 2 7 3 13 10 9 13 0 2
11 11 11 11 13 9 9 9 11 9 12 2
23 3 15 13 9 10 11 2 16 1 9 13 2 9 10 13 1 9 0 7 9 2 9 2
16 11 2 11 3 13 1 9 7 9 0 3 0 1 9 0 2
17 9 10 13 9 9 10 0 1 13 7 13 1 10 9 15 13 2
19 11 11 2 9 10 2 10 1 9 11 2 13 10 9 1 9 1 11 2
54 7 9 10 13 11 11 11 11 11 2 11 11 11 15 0 13 1 10 9 7 9 2 2 9 9 10 3 13 13 1 9 12 1 11 11 11 11 11 11 11 11 2 11 11 11 2 7 15 0 13 11 11 11 2
26 9 9 2 9 2 7 9 13 9 1 12 9 2 15 13 1 13 9 9 9 12 7 9 9 11 2
44 11 11 11 11 3 13 9 2 11 2 1 11 11 11 11 11 11 11 11 2 16 13 1 9 9 11 11 11 9 2 12 5 11 2 11 5 11 2 12 5 12 5 12 2
26 9 10 3 13 1 9 11 11 2 13 1 9 12 11 12 1 11 9 11 2 12 5 12 5 12 2
13 9 10 12 9 15 13 1 13 11 1 9 11 2
30 10 9 11 11 2 1 12 5 1 9 3 2 9 2 13 1 11 2 16 9 11 11 10 0 13 1 9 0 11 2
30 11 13 13 9 1 9 2 9 9 1 11 11 2 9 9 15 13 1 11 11 2 11 2 11 11 9 7 11 11 2
10 11 11 11 11 11 13 9 9 12 2
5 15 13 1 9 2
9 11 0 13 1 11 11 11 11 2
29 11 15 13 1 11 11 12 11 2 11 11 12 11 13 9 0 15 13 0 7 3 13 7 9 9 9 9 9 2
15 1 9 12 2 11 11 11 13 2 15 3 13 11 11 2
18 16 3 13 9 0 1 13 1 9 11 2 15 11 11 13 9 10 2
15 16 11 14 13 1 9 9 11 2 11 13 11 1 9 2
53 11 13 1 13 9 15 0 2 16 11 13 0 1 9 1 10 9 3 2 7 16 11 13 9 12 5 12 1 9 12 7 13 0 1 9 9 1 11 11 2 1 9 1 9 10 2 15 13 1 11 11 11 2
12 11 2 11 11 13 9 1 11 11 11 11 2
11 14 13 9 9 2 2 3 15 13 15 2
20 9 10 1 9 13 1 9 9 2 7 9 9 9 9 15 13 10 9 9 2
19 1 9 14 0 2 15 3 13 1 9 0 7 13 0 1 10 9 0 2
9 11 11 13 1 9 12 11 12 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
8 1 9 10 3 11 11 13 2
27 11 13 1 9 9 9 11 11 11 11 11 1 9 12 7 13 9 1 9 2 9 9 1 9 9 9 2
28 11 10 13 1 11 11 7 11 11 1 9 2 11 11 1 9 2 11 11 1 9 2 7 11 11 1 9 2
20 1 9 12 2 9 1 9 9 2 11 13 11 15 13 9 9 2 11 12 2
29 1 9 1 11 11 2 11 11 13 7 13 1 9 11 2 15 13 1 0 11 2 15 3 0 13 1 11 11 2
27 9 1 9 9 10 3 11 11 13 3 13 7 9 9 10 13 9 9 9 2 11 11 11 2 11 2 2
42 11 11 2 11 2 7 2 11 11 2 11 2 9 12 9 11 2 2 13 9 0 1 9 11 10 9 15 13 1 9 12 9 11 7 11 12 2 12 1 9 11 2
18 11 11 13 10 9 1 9 11 11 2 11 11 2 11 11 2 11 2
40 10 13 7 3 13 11 2 11 2 11 11 2 11 3 13 7 13 11 15 3 13 11 11 11 11 1 11 1 9 7 9 1 11 11 11 11 1 11 11 2
