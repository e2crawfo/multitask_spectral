8907 11
11 1 9 2 13 2 14 15 13 0 9 2
9 0 9 2 13 2 15 4 13 2
8 1 9 2 15 6 13 15 2
6 3 2 15 13 9 2
13 15 2 13 15 2 6 13 14 15 13 1 15 2
9 3 2 0 6 4 13 1 9 2
9 9 15 2 6 2 13 0 0 2
8 10 9 1 9 6 13 11 2
6 14 6 4 13 0 2
5 14 13 14 13 2
5 14 15 13 3 2
6 14 15 13 14 3 2
6 14 14 15 13 3 2
5 13 14 14 13 2
5 13 14 14 13 2
5 13 14 14 13 2
13 15 6 4 14 13 10 15 13 1 15 1 9 2
13 15 6 4 14 13 10 15 13 1 15 1 9 2
6 13 14 14 15 13 2
11 7 15 1 9 6 2 6 2 6 2 2
4 15 2 6 2
6 7 13 0 1 9 2
9 11 11 6 15 13 1 9 15 2
4 13 15 9 2
8 3 11 13 1 9 15 11 2
8 0 9 15 13 12 0 9 2
11 15 13 1 9 7 15 13 0 0 9 2
8 1 9 15 4 13 0 9 2
10 1 10 9 11 13 1 0 9 3 2
6 9 1 15 13 3 2
9 1 9 15 13 9 1 0 9 2
14 3 15 13 10 9 3 2 15 4 13 14 13 3 2
7 13 15 9 1 9 11 2
6 9 15 13 0 9 2
5 9 15 13 3 2
9 9 15 4 13 1 9 1 9 2
12 10 9 2 3 1 11 2 1 9 13 11 2
15 1 9 1 9 2 1 0 9 2 15 13 0 9 9 2
11 1 1 10 9 2 9 15 13 1 9 2
13 11 11 2 1 0 15 9 2 2 13 14 13 2
12 13 3 1 9 2 9 3 4 13 1 9 2
7 3 13 9 1 9 15 2
6 3 15 9 13 9 2
8 3 0 9 13 0 15 9 2
7 0 9 13 3 7 3 2
10 3 3 15 13 1 9 1 0 9 2
8 3 9 11 15 13 3 3 2
7 9 3 3 15 4 13 2
7 3 15 13 1 9 9 2
9 15 3 6 15 13 1 0 9 2
13 15 3 13 1 10 9 2 7 3 13 14 13 2
5 11 15 13 3 2
6 11 15 13 3 3 2
8 15 13 0 2 14 13 3 2
5 15 15 13 3 2
6 3 13 2 3 13 2
11 9 1 3 1 15 15 4 13 1 9 2
5 1 9 13 9 2
4 11 13 3 2
9 1 0 9 1 9 15 13 9 2
9 1 0 9 1 9 15 13 9 2
8 13 4 15 1 10 0 9 2
7 1 0 9 13 0 9 2
7 3 15 13 0 0 9 2
8 1 10 9 15 13 0 9 2
7 1 9 15 15 13 9 2
6 0 9 3 15 13 2
9 3 7 11 7 11 13 1 9 2
10 15 3 13 1 9 7 13 1 9 2
6 9 15 13 1 3 2
7 1 9 15 13 0 9 2
6 13 9 15 1 9 2
6 3 13 1 9 15 2
6 3 13 1 9 15 2
6 11 3 13 9 15 2
7 9 15 3 15 13 9 2
7 1 9 3 13 10 9 2
5 3 13 1 15 2
5 9 13 1 9 2
7 11 13 1 9 1 9 2
6 15 15 13 3 3 2
7 9 15 15 13 1 9 2
15 9 9 9 15 4 13 1 9 1 0 9 1 0 9 2
5 11 13 1 9 2
5 1 9 13 15 2
16 13 15 1 9 15 2 13 15 2 6 13 1 9 7 9 2
10 12 9 13 0 11 1 0 15 9 2
6 9 15 13 1 9 2
6 9 15 13 1 9 2
5 13 1 0 9 2
6 11 15 13 1 9 2
5 9 13 1 9 2
6 14 15 13 1 9 2
12 3 6 15 13 1 15 2 3 13 1 9 2
6 6 2 13 2 9 2
7 1 9 13 9 7 9 2
7 15 13 15 9 7 9 2
4 13 9 9 2
4 0 15 13 2
9 9 11 11 4 13 1 0 9 2
13 13 7 12 2 11 2 11 7 9 1 9 15 2
7 13 7 15 1 9 11 2
19 3 9 2 3 7 0 9 1 0 9 13 1 9 7 9 1 0 9 2
4 15 15 13 2
4 15 15 13 2
6 12 13 9 1 9 2
8 6 13 2 9 15 2 14 2
9 9 15 13 1 15 7 15 13 2
8 0 3 2 14 13 0 9 2
6 15 1 11 13 3 2
9 10 9 2 10 9 6 15 13 2
8 7 9 2 6 2 6 13 2
5 15 3 9 13 2
5 9 2 13 3 2
6 3 9 7 9 13 2
5 12 11 6 13 2
12 11 2 11 7 15 14 13 1 9 1 9 2
12 1 9 1 9 1 9 15 13 9 1 9 2
11 0 9 1 9 13 1 12 9 1 9 2
10 9 6 13 15 1 9 1 9 15 2
6 0 1 0 6 13 2
6 0 13 2 13 3 2
5 0 6 14 13 2
8 0 3 13 2 9 15 13 2
8 9 13 1 9 1 0 9 2
7 10 9 1 9 15 13 2
6 15 13 9 1 9 2
11 15 13 0 0 9 2 15 4 15 13 2
7 14 13 15 2 0 9 2
10 15 13 10 9 9 2 0 9 13 2
6 9 11 13 0 9 2
10 9 11 15 13 1 9 1 0 9 2
10 9 9 13 9 1 9 7 13 3 2
6 9 11 13 14 13 2
8 9 11 15 13 9 1 9 2
7 9 11 13 0 15 9 2
13 15 14 4 15 13 2 13 14 15 13 15 15 2
10 16 13 9 2 15 4 13 3 9 2
8 15 15 13 1 0 0 9 2
3 14 13 2
8 11 13 3 0 1 9 15 2
6 0 2 14 4 13 2
10 13 10 9 2 1 14 13 9 15 2
10 7 13 15 9 0 2 0 7 0 2
9 0 9 14 4 13 1 0 9 2
11 3 4 13 1 9 7 9 1 0 9 2
9 9 13 9 1 9 7 15 13 2
10 0 7 0 0 9 4 13 0 9 2
14 10 9 14 14 15 4 13 1 9 3 1 9 15 2
8 9 4 13 1 9 7 9 2
12 13 15 15 2 16 3 13 3 1 0 9 2
8 15 13 9 1 3 0 9 2
14 7 1 9 6 13 1 9 2 7 15 13 1 9 2
6 9 13 0 15 9 2
12 9 13 2 15 15 13 2 7 7 15 13 2
6 0 12 9 13 0 2
12 7 15 14 15 13 3 7 3 14 13 0 2
6 11 11 13 9 15 2
5 15 15 13 9 2
8 0 13 2 7 9 6 13 2
5 3 9 13 15 2
14 13 9 7 13 9 0 2 13 15 2 13 0 9 2
5 11 13 9 9 2
7 15 15 13 1 10 9 2
6 15 13 14 15 13 2
13 9 13 2 13 1 9 7 13 3 1 0 9 2
15 3 15 6 13 15 2 7 15 13 3 7 13 0 9 2
19 10 9 4 13 2 4 13 2 13 15 4 2 7 1 9 13 15 0 2
7 13 15 9 1 0 9 2
11 13 15 11 2 3 4 13 1 0 9 2
10 15 13 3 3 7 0 1 0 9 2
10 11 9 2 3 11 9 15 15 13 2
8 11 13 1 0 9 1 9 2
12 15 6 13 9 1 10 9 2 7 13 9 2
21 1 9 15 13 0 9 2 9 2 0 9 2 7 1 15 9 1 9 13 11 2
13 3 1 9 3 13 9 2 7 3 13 0 9 2
16 7 9 15 13 1 9 2 7 1 9 15 13 9 7 9 2
16 9 15 2 0 7 0 2 13 9 2 7 9 15 13 0 2
14 1 12 9 1 15 13 11 2 7 15 6 15 13 2
12 6 13 1 9 2 7 13 14 13 9 3 2
20 10 9 0 9 3 13 0 1 0 9 2 7 3 6 4 15 13 1 9 2
10 13 15 4 2 7 9 15 15 13 2
12 13 9 2 0 10 2 7 15 6 15 13 2
17 14 15 13 14 2 14 15 13 14 2 7 14 15 13 0 9 2
10 7 15 13 2 7 3 6 15 13 2
18 7 10 9 13 3 0 1 0 9 2 7 14 13 3 3 1 9 2
15 7 13 14 13 9 15 2 7 14 15 13 1 0 9 2
7 6 13 14 13 14 13 2
8 6 4 13 14 13 14 13 2
9 0 9 4 13 14 13 1 11 2
11 1 12 9 13 14 13 14 13 0 9 2
8 9 13 14 13 0 7 0 2
7 15 13 14 13 1 15 2
12 15 15 13 14 15 13 3 2 16 15 13 2
8 1 9 13 2 16 4 13 2
6 13 2 16 13 3 2
5 13 10 15 13 2
19 10 0 9 15 13 1 9 1 0 9 7 15 13 14 13 1 9 15 2
10 13 14 15 13 3 3 14 15 13 2
15 7 14 13 14 15 13 1 15 0 2 0 15 9 9 2
7 13 15 14 15 13 3 2
10 6 13 14 15 4 13 9 1 9 2
7 6 13 14 4 13 15 2
8 6 13 14 15 13 14 15 2
9 6 13 14 3 14 13 1 15 2
9 6 13 3 14 15 13 1 9 2
9 6 13 14 15 13 14 4 13 2
9 6 13 14 4 15 13 1 15 2
8 3 4 13 14 15 13 9 2
9 13 15 3 14 13 1 10 9 2
5 13 15 15 13 2
8 13 15 14 13 0 7 0 2
6 13 3 14 13 3 2
10 13 2 16 1 10 9 13 3 0 2
9 13 15 14 6 13 14 13 9 2
6 13 15 15 4 13 2
11 3 1 9 1 0 9 13 14 13 9 2
10 0 9 4 15 13 14 13 1 9 2
8 15 13 2 16 4 13 9 2
7 16 15 13 2 13 3 2
9 14 15 13 2 16 13 10 9 2
15 15 13 2 16 3 14 13 2 1 16 4 13 1 9 2
10 1 14 13 15 2 14 13 14 15 2
10 1 14 15 13 2 15 13 9 15 2
22 9 1 0 9 13 0 2 1 3 15 13 2 16 0 0 9 13 9 14 13 0 2
12 13 3 14 13 1 15 2 1 3 13 9 2
9 13 15 1 9 3 15 13 9 2
6 13 15 3 13 9 2
14 3 15 13 3 2 15 3 6 4 13 3 10 9 2
7 3 13 2 9 6 13 2
13 7 3 3 6 13 14 15 13 2 3 4 13 2
9 15 13 14 15 13 2 3 13 2
7 13 2 3 4 15 13 2
8 9 13 2 3 14 15 13 2
13 6 15 13 2 14 15 13 2 1 15 14 13 2
13 3 2 15 13 14 13 1 9 2 3 13 3 2
9 9 2 3 15 13 2 4 13 2
8 3 7 14 13 2 3 13 2
11 1 14 13 3 0 2 13 14 13 9 2
14 1 16 15 13 9 2 15 0 9 6 13 14 13 2
9 6 13 0 2 7 6 15 13 2
10 13 4 4 14 13 2 3 4 13 2
19 1 9 13 0 0 9 2 3 9 13 0 2 0 2 0 2 1 0 2
7 13 4 2 3 15 13 2
12 13 15 3 2 7 13 14 13 0 15 9 2
7 9 14 13 14 15 13 2
8 16 15 13 2 14 15 13 2
6 16 13 2 13 3 2
6 16 13 2 13 3 2
10 16 15 13 3 2 13 14 15 13 2
10 16 15 13 9 2 4 13 1 9 2
9 16 6 13 9 2 6 13 9 2
6 16 14 13 2 13 2
11 13 1 12 7 16 6 13 2 15 13 2
9 1 9 16 13 2 14 15 13 2
9 14 13 9 2 15 4 15 13 2
8 9 14 13 2 14 15 13 2
11 3 14 15 13 2 6 13 15 9 3 2
10 13 15 14 13 2 1 14 15 13 2
7 7 15 13 14 15 13 2
7 7 15 13 14 15 13 2
5 13 14 15 13 2
8 3 9 15 13 9 14 13 2
6 13 15 14 13 9 2
7 13 3 2 3 0 13 2
13 13 3 2 3 13 9 2 16 15 6 15 13 2
16 6 13 14 13 9 1 9 2 3 13 0 1 15 1 15 2
12 15 13 3 2 3 9 15 13 0 1 9 2
16 3 3 13 3 0 2 15 15 13 1 0 9 1 9 15 2
5 13 15 14 13 2
11 14 13 2 16 14 15 13 1 0 9 2
19 7 10 9 13 14 13 2 16 9 15 13 7 9 15 13 1 9 15 2
6 4 13 2 16 13 2
13 4 15 13 1 12 9 1 9 2 3 13 9 2
9 14 13 2 16 6 4 13 9 2
9 14 13 2 16 6 4 13 9 2
9 16 13 9 2 13 14 15 13 2
9 16 13 9 2 13 14 15 13 2
12 16 14 13 2 16 13 2 13 15 1 9 2
11 16 15 13 3 1 9 2 9 13 9 2
9 7 13 12 9 2 3 13 3 2
18 3 15 13 1 9 1 9 7 16 15 13 2 3 15 13 1 15 2
9 13 15 2 1 3 14 15 13 2
9 16 13 9 15 2 14 15 13 2
16 16 15 13 0 9 1 11 2 9 13 2 16 15 13 0 2
18 9 15 13 1 0 9 7 13 1 0 9 2 3 4 15 13 3 2
14 3 3 14 13 1 9 2 15 3 15 13 7 13 2
7 3 13 2 15 13 3 2
7 3 13 2 15 13 3 2
15 13 0 9 1 10 9 1 9 2 16 0 15 13 3 2
10 7 3 13 9 15 2 15 15 13 2
16 7 9 15 13 3 3 2 3 13 12 9 1 9 1 9 2
10 3 15 13 2 6 13 3 1 9 2
11 13 2 7 1 14 15 13 2 15 13 2
15 3 14 15 13 2 9 2 13 15 9 2 16 15 13 2
12 1 14 13 1 0 9 2 0 13 2 13 2
12 15 13 0 15 9 2 3 15 13 1 9 2
11 12 9 13 3 2 3 1 11 13 9 2
12 13 14 13 12 9 2 16 13 9 1 9 2
16 3 15 13 7 13 1 9 15 2 3 15 15 13 1 9 2
8 16 13 2 13 15 1 9 2
11 16 9 13 2 3 15 15 13 1 9 2
11 16 15 13 9 1 9 2 3 9 13 2
7 15 13 9 3 14 13 2
15 13 15 9 2 10 13 14 15 13 3 1 10 0 9 2
9 10 2 15 13 2 4 13 3 2
11 14 9 15 13 1 9 3 14 4 13 2
21 3 14 9 15 13 1 9 1 10 9 2 1 10 11 15 13 1 9 1 9 2
15 13 2 9 2 9 2 14 13 9 2 15 14 15 13 2
15 13 2 9 2 9 2 14 13 9 2 15 14 15 13 2
9 10 9 13 3 2 15 13 3 2
11 3 9 2 15 4 13 2 13 0 9 2
14 7 7 1 0 9 13 9 2 3 9 13 7 13 2
14 7 1 15 7 9 2 3 13 9 2 13 0 9 2
30 1 9 1 9 13 2 16 0 9 1 10 9 1 0 9 13 9 1 9 0 9 2 10 9 15 13 1 0 9 2
11 3 7 13 10 2 15 4 13 1 9 2
8 3 14 13 15 14 15 13 2
12 3 13 2 3 0 9 4 13 1 0 9 2
6 15 13 2 3 13 2
10 9 13 2 3 6 15 13 1 15 2
7 6 13 3 14 15 13 2
12 7 13 2 16 11 3 4 13 1 9 3 2
11 9 13 2 16 13 3 2 16 13 9 2
12 3 3 13 2 16 15 15 4 13 1 15 2
8 3 13 2 16 4 13 9 2
13 3 6 13 15 2 15 14 13 14 13 10 9 2
15 9 1 9 7 9 13 2 15 13 9 1 10 0 9 2
11 0 9 1 15 13 10 9 14 15 13 2
10 14 9 15 13 2 16 9 6 13 2
16 1 0 9 9 14 15 13 1 15 7 14 15 13 1 9 2
17 12 9 13 3 0 9 2 7 9 4 13 2 7 9 4 13 2
10 11 13 2 7 13 1 11 1 9 2
9 13 9 2 7 15 13 1 9 2
20 15 13 9 7 3 3 3 7 1 9 13 1 9 1 9 7 13 1 9 2
8 7 15 13 2 7 15 13 2
9 14 13 2 7 10 13 14 13 2
7 13 0 9 1 0 9 2
6 9 13 1 0 9 2
9 13 1 0 9 2 1 0 9 2
7 1 0 0 9 13 9 2
10 10 0 9 1 9 11 15 13 9 2
12 10 0 7 0 9 13 1 0 9 1 9 2
10 3 1 9 2 0 9 13 0 9 2
10 1 0 2 0 9 15 13 1 9 2
12 15 13 0 2 0 9 1 11 1 0 9 2
10 9 13 1 0 1 9 9 1 11 2
11 0 7 0 9 13 1 0 1 9 9 2
6 13 14 3 14 13 2
16 0 9 4 13 14 13 9 7 13 0 9 1 0 0 9 2
6 13 16 13 0 9 2
6 9 13 14 13 9 2
5 9 13 14 13 2
6 9 13 14 13 3 2
15 10 0 9 4 13 14 13 10 9 1 0 7 0 9 2
5 13 14 15 13 2
13 13 15 2 9 2 13 2 7 1 0 9 13 2
6 11 13 14 13 3 2
12 14 15 15 13 11 14 13 7 1 1 9 2
12 11 13 14 15 13 7 13 3 14 13 0 2
9 7 9 13 14 15 13 1 9 2
9 9 7 9 6 13 14 15 13 2
13 3 13 14 13 9 2 3 13 9 7 9 13 2
7 0 9 15 13 14 13 2
8 9 13 2 6 13 14 13 2
7 3 11 13 14 15 13 2
6 9 13 14 15 13 2
6 11 15 13 14 13 2
7 6 13 14 15 13 14 2
6 9 13 14 15 13 2
9 1 15 6 13 7 9 14 13 2
10 9 13 14 15 13 1 9 3 3 2
15 0 15 3 9 13 14 15 13 7 14 15 13 1 9 2
9 13 14 13 2 6 13 0 15 2
4 13 13 9 2
10 15 6 13 14 13 1 9 1 9 2
15 15 6 13 14 13 9 15 2 1 14 6 13 9 15 2
6 15 13 14 13 9 2
12 14 13 14 13 10 9 2 13 15 13 3 2
8 7 14 15 13 9 7 0 2
10 7 10 0 2 0 9 9 15 13 2
5 13 0 7 0 2
7 11 15 13 3 9 3 2
11 1 0 3 9 9 15 13 0 7 0 2
18 9 9 11 2 15 13 1 0 9 1 10 0 9 7 1 0 9 2
14 7 3 15 15 13 1 12 1 0 9 1 9 15 2
9 7 3 15 13 14 15 13 0 2
5 11 13 1 0 2
9 9 3 15 15 13 0 7 0 2
7 9 15 13 0 1 9 2
7 11 15 13 1 9 15 2
13 13 15 2 13 15 1 0 2 16 15 6 13 2
7 9 15 13 0 7 0 2
6 9 15 13 10 9 2
8 11 13 0 9 1 9 11 2
6 9 15 15 13 0 2
21 1 9 7 1 9 15 15 13 0 9 1 9 7 3 2 7 3 1 0 9 2
9 13 14 15 13 0 1 0 9 2
10 13 15 9 15 2 9 15 13 0 2
6 9 1 11 13 0 2
3 13 9 2
15 15 15 13 1 0 9 2 1 0 9 2 1 0 9 2
9 10 9 15 15 13 0 1 9 2
16 15 13 2 16 10 11 3 0 13 2 3 13 15 7 9 2
14 15 13 0 7 0 2 1 15 9 1 9 13 0 2
9 15 13 0 1 0 9 1 11 2
6 15 13 7 3 9 2
7 15 13 9 1 0 9 2
10 15 13 0 2 6 13 3 1 9 2
9 1 9 15 15 13 9 1 15 2
10 13 3 0 9 14 13 1 0 9 2
8 13 15 9 9 1 10 9 2
13 11 13 9 15 7 13 3 2 16 6 13 3 2
3 10 9 2
3 10 9 2
6 13 15 9 1 9 2
5 13 9 1 9 2
6 9 15 13 10 9 2
6 13 15 9 1 15 2
21 0 15 9 13 2 1 9 0 2 2 0 9 9 13 2 2 1 10 9 0 2
9 15 13 1 9 1 10 0 9 2
8 13 14 15 13 9 1 9 2
7 13 15 9 1 0 9 2
7 15 6 13 9 1 9 2
8 9 0 2 3 0 13 15 2
7 1 10 9 13 0 9 2
6 1 10 9 13 9 2
2 14 2
3 13 15 2
7 7 3 14 13 2 13 2
3 13 15 2
5 0 9 2 14 2
5 3 0 13 9 2
6 13 1 0 0 9 2
6 1 10 9 9 13 2
3 13 9 2
10 16 13 12 9 2 6 15 13 3 2
10 16 13 14 13 2 13 15 14 13 2
7 3 13 2 3 6 13 2
9 13 0 9 2 13 15 2 13 2
9 13 15 3 1 9 1 0 9 2
6 1 9 13 10 9 2
9 9 13 9 2 9 2 9 13 2
8 9 2 9 2 9 7 9 2
8 7 15 13 2 7 15 13 2
6 9 6 13 3 3 2
5 15 15 6 13 2
10 9 3 6 4 15 13 1 0 9 2
18 14 7 14 15 13 14 15 13 1 11 2 3 15 13 14 13 3 2
7 15 6 4 13 1 15 2
7 3 1 9 15 13 9 2
9 1 10 9 15 15 6 15 13 2
16 15 13 9 2 15 13 9 2 15 13 10 0 9 1 9 2
5 15 3 9 13 2
8 7 12 4 13 2 13 9 2
7 14 13 15 2 0 9 2
5 1 9 13 9 2
10 1 9 13 14 15 13 1 10 9 2
18 3 1 0 12 9 1 9 15 15 15 13 14 13 1 0 15 9 2
18 3 1 0 12 9 1 9 15 15 15 13 14 13 1 0 15 9 2
17 1 15 13 7 9 2 7 10 0 9 2 15 3 6 13 13 2
5 9 13 14 13 2
3 13 9 2
6 15 6 13 15 13 2
8 9 6 13 15 14 15 13 2
6 15 13 14 13 9 2
12 13 14 15 9 1 9 2 13 15 13 3 2
8 6 13 14 13 14 13 3 2
11 3 15 13 10 9 0 2 0 2 0 2
19 2 3 13 2 13 15 2 2 16 13 14 13 1 9 9 15 1 15 2
15 1 9 13 10 9 2 6 15 13 7 9 2 7 9 2
7 9 15 13 1 12 9 2
10 9 13 14 13 0 2 0 2 0 2
8 3 15 13 15 2 13 9 2
6 10 13 1 10 9 2
6 3 15 13 1 15 2
5 9 13 1 15 2
5 9 13 1 15 2
14 15 3 13 9 2 3 13 3 3 14 13 1 15 2
17 3 2 13 15 1 10 9 2 15 13 3 0 1 9 1 9 2
6 9 13 3 3 3 2
6 9 13 3 3 3 2
13 15 14 13 2 7 13 2 16 9 15 13 3 2
9 9 3 3 13 14 13 3 3 2
12 13 2 16 3 13 3 7 6 13 14 13 2
16 13 15 10 14 14 9 11 2 13 14 13 2 13 9 9 2
11 15 13 9 1 12 15 9 2 13 9 2
10 15 15 13 2 15 15 13 1 9 2
9 12 0 9 15 13 9 10 9 2
5 15 15 13 9 2
8 11 3 15 13 9 1 9 2
9 1 12 9 15 13 3 1 15 2
10 3 7 3 13 9 7 9 1 11 2
15 1 0 0 9 15 3 14 4 13 14 13 0 0 9 2
8 1 10 9 15 13 9 9 2
6 1 9 13 0 9 2
6 9 15 13 1 9 2
6 3 13 3 0 9 2
6 9 13 1 12 9 2
17 16 3 9 3 13 0 9 7 0 9 2 9 3 13 0 9 2
14 1 7 1 3 9 2 6 13 14 13 3 0 9 2
9 3 3 15 13 9 1 10 9 2
9 3 9 15 15 13 1 10 9 2
6 15 15 13 3 3 2
5 15 15 13 3 2
6 13 0 2 0 9 2
9 15 13 1 12 9 7 12 9 2
16 1 0 9 7 9 2 1 0 9 7 0 9 13 0 9 2
21 9 11 15 13 7 16 13 0 2 3 0 9 2 13 15 7 15 13 1 9 2
7 13 0 9 1 0 9 2
7 9 11 13 7 15 13 2
6 10 9 13 1 9 2
17 15 9 2 1 0 15 9 2 13 15 3 9 13 14 13 9 2
10 10 9 7 10 9 13 1 9 15 2
9 1 10 9 11 6 13 0 9 2
9 10 9 2 10 9 6 15 13 2
12 13 9 2 13 9 7 0 9 9 13 9 2
7 0 9 9 13 1 11 2
5 13 9 0 9 2
13 15 13 1 9 1 9 2 1 0 9 1 9 2
10 3 4 13 3 15 13 0 15 9 2
18 9 15 13 3 1 9 1 15 7 3 3 15 13 9 14 15 13 2
19 7 9 0 1 9 0 2 7 9 2 6 13 9 1 15 14 13 9 2
7 10 9 13 9 1 15 2
13 1 9 1 15 7 1 0 9 3 13 9 9 2
21 1 0 15 0 9 3 13 9 1 9 2 3 15 13 14 13 0 0 9 3 2
14 3 15 13 10 9 3 2 15 4 13 14 13 3 2
18 9 15 13 14 13 2 7 10 3 15 13 7 15 13 14 15 13 2
15 1 9 3 15 13 9 2 10 0 9 15 13 1 9 2
8 0 9 3 13 1 9 9 2
25 7 3 4 13 7 1 9 2 7 1 9 2 14 13 2 3 13 2 1 10 0 9 7 9 2
15 15 6 13 14 15 13 1 10 9 2 1 10 0 9 2
14 1 10 0 0 9 11 6 13 7 9 2 7 9 2
7 7 0 4 13 9 11 2
13 3 15 13 0 7 15 15 13 2 16 13 3 2
6 13 12 14 15 13 2
9 13 15 3 1 0 7 0 9 2
8 9 2 0 2 13 1 9 2
17 10 9 2 0 1 0 9 7 0 9 2 13 3 0 7 0 2
11 9 2 0 7 0 2 13 3 1 15 2
16 9 15 13 3 0 7 13 9 1 9 15 2 0 7 0 2
15 9 2 0 1 0 9 1 12 15 9 2 13 1 9 2
4 9 15 13 2
11 15 13 10 9 1 9 2 3 7 9 2
20 3 2 3 3 2 1 3 1 12 9 2 9 1 9 11 4 13 10 9 2
15 1 0 9 13 0 0 9 2 9 13 2 13 15 9 2
7 15 13 9 7 9 13 2
16 9 15 13 3 7 1 9 2 9 15 13 1 10 0 9 2
20 11 13 3 2 13 9 2 13 9 2 13 15 2 13 0 9 2 13 9 2
13 3 15 9 13 9 2 7 9 15 3 9 13 2
14 9 13 9 15 2 7 13 1 9 7 13 1 9 2
19 7 15 13 1 9 7 9 2 7 15 13 7 15 13 1 9 1 9 2
9 13 9 2 7 15 13 1 9 2
10 9 13 9 2 7 9 6 15 13 2
14 3 3 13 1 0 9 2 7 1 9 9 15 13 2
13 14 13 15 9 2 7 14 13 1 9 1 9 2
10 15 6 13 9 2 3 13 0 9 2
25 15 15 13 1 9 2 13 9 2 13 15 1 9 2 7 6 13 14 13 1 0 9 1 9 2
7 15 13 2 9 6 13 2
10 15 13 1 9 1 9 2 6 13 2
14 3 13 14 15 13 2 16 9 13 7 15 13 3 2
15 15 13 0 15 9 2 10 9 3 6 15 13 1 9 2
8 7 12 13 9 14 13 9 2
9 13 1 9 14 6 4 13 9 2
10 3 15 15 13 9 14 13 9 15 2
9 6 15 13 3 3 15 13 3 2
12 15 6 13 14 0 9 13 3 0 1 15 2
12 9 2 1 14 13 2 11 15 13 1 9 2
12 9 2 1 14 13 2 11 15 13 1 9 2
14 3 2 16 15 13 1 9 9 2 13 14 13 9 2
12 9 13 3 0 2 16 9 15 13 1 9 2
15 13 1 9 9 2 3 16 0 9 13 14 13 1 9 2
20 15 13 1 15 7 13 9 2 16 14 15 13 15 13 9 16 14 15 13 2
12 16 6 4 15 13 2 13 14 15 13 9 2
11 14 6 4 13 15 2 16 9 15 13 2
9 14 15 13 2 16 14 13 9 2
17 7 9 14 13 2 13 15 1 9 2 13 9 15 7 15 13 2
19 3 13 14 13 14 9 1 15 2 1 16 9 3 15 13 1 9 15 2
19 15 6 13 14 13 0 9 1 9 2 1 16 4 13 1 9 1 9 2
7 9 15 13 14 13 3 2
13 1 9 15 13 11 3 13 9 1 9 1 9 2
10 15 15 13 2 16 15 6 4 13 2
42 13 9 2 15 13 2 13 9 2 15 13 2 13 11 2 15 13 3 1 9 2 13 9 2 15 13 2 7 13 2 16 13 0 1 10 9 2 16 3 13 9 2
25 15 15 13 1 0 9 1 9 2 3 9 13 9 1 9 2 7 3 13 0 9 7 0 9 2
6 2 13 14 15 13 2
10 11 13 14 15 13 2 16 15 13 2
4 11 15 13 2
4 2 13 15 2
6 13 14 9 1 11 2
4 2 13 15 2
7 9 13 2 16 13 0 2
3 3 13 2
4 2 3 13 2
6 6 15 15 13 3 2
5 13 9 1 15 2
5 13 9 1 15 2
6 6 13 15 14 13 2
7 6 13 14 6 4 13 2
10 13 15 15 2 16 15 13 10 9 2
7 15 4 13 10 10 9 2
6 9 9 13 12 9 2
8 3 13 14 15 13 14 13 2
5 13 15 7 15 2
7 15 6 13 3 1 15 2
6 13 15 10 0 9 2
6 10 0 9 15 13 2
8 13 14 6 4 15 15 13 2
8 13 14 6 15 15 4 13 2
8 13 14 6 4 15 15 13 2
7 13 14 4 15 15 13 2
7 13 14 4 15 15 13 2
7 13 14 15 15 4 13 2
7 13 14 4 15 15 13 2
5 13 14 13 15 2
6 13 2 16 13 15 2
5 9 15 13 0 2
5 13 15 14 13 2
5 15 13 14 13 2
5 15 13 14 13 2
5 15 13 14 13 2
5 15 13 14 13 2
5 13 15 14 13 2
6 15 6 13 14 13 2
6 14 4 15 15 13 2
12 14 4 15 15 13 2 13 13 13 14 13 2
6 15 10 13 3 3 2
5 9 3 13 3 2
9 10 10 9 1 10 9 15 13 2
7 9 13 1 15 1 15 2
9 13 15 15 2 16 13 10 9 2
5 13 15 1 9 2
3 13 14 2
3 2 13 2
6 3 13 15 14 13 2
6 6 13 15 14 13 2
5 13 15 14 13 2
8 13 14 13 14 13 14 13 2
5 13 15 14 13 2
6 6 13 15 14 13 2
5 13 15 14 13 2
8 13 15 14 15 13 14 13 2
5 13 14 13 9 2
5 3 13 14 13 2
7 3 13 2 16 4 13 2
9 9 2 15 13 15 2 4 13 2
10 15 13 15 2 3 9 15 15 13 2
10 15 13 15 2 3 9 15 15 13 2
9 15 13 9 2 1 15 13 15 2
7 13 9 14 13 1 9 2
8 13 15 9 2 3 13 15 2
5 14 13 1 15 2
6 14 15 13 3 13 2
10 15 13 3 3 2 3 15 13 3 2
7 13 1 0 3 4 13 2
6 13 2 3 15 13 2
7 13 1 9 14 13 15 2
5 13 14 15 13 2
7 9 4 13 1 9 15 2
7 9 4 13 1 9 15 2
7 9 4 13 1 9 15 2
11 15 13 2 16 9 1 15 14 13 0 2
5 15 15 13 9 2
5 15 15 13 9 2
6 15 15 13 1 9 2
6 15 15 13 1 9 2
6 15 9 14 13 3 2
8 3 1 9 2 15 15 13 2
9 3 1 9 2 15 14 13 3 2
5 9 15 15 13 2
5 9 15 15 13 2
8 15 15 13 2 14 6 13 2
8 1 12 9 14 11 14 13 2
6 13 9 15 14 11 2
6 13 14 15 15 4 2
14 15 13 9 2 15 15 13 2 16 4 13 1 15 2
8 15 13 9 2 15 15 13 2
6 13 15 9 14 13 2
7 15 13 2 16 4 13 2
12 15 13 9 2 15 15 15 13 14 4 13 2
7 15 15 13 14 4 13 2
10 11 15 13 2 16 11 15 4 13 2
9 15 15 13 2 1 14 15 13 2
7 6 13 2 1 14 13 2
5 10 9 15 13 2
5 15 15 13 3 2
7 13 15 14 15 13 3 2
6 0 1 15 9 13 2
7 13 1 15 7 1 15 2
10 15 13 0 9 2 7 15 15 13 2
8 15 13 12 0 9 0 9 2
9 13 15 9 0 2 0 7 0 2
6 9 9 13 1 9 2
6 9 9 13 1 9 2
7 9 1 9 13 1 9 2
5 15 9 14 13 2
6 9 9 13 1 9 2
6 15 13 12 0 9 2
10 12 9 15 13 1 10 1 10 9 2
5 3 9 13 3 2
6 15 15 13 3 3 2
6 10 15 13 3 3 2
6 13 14 9 1 3 2
5 13 14 9 3 2
7 13 14 9 1 10 9 2
6 13 9 1 9 3 2
8 9 1 9 1 11 13 0 2
8 9 1 9 1 11 13 0 2
8 9 1 15 14 13 0 3 2
8 9 1 15 14 13 0 3 2
8 9 1 15 14 13 0 3 2
5 15 13 15 14 2
6 15 13 0 9 9 2
7 15 13 0 9 1 9 2
6 15 13 3 3 13 2
6 15 13 3 1 9 2
7 15 4 13 1 1 9 2
7 15 15 13 1 0 9 2
6 15 15 13 1 0 2
6 10 9 6 13 0 2
5 10 9 4 13 2
7 10 9 4 13 1 9 2
5 15 13 9 3 2
6 15 13 1 15 3 2
6 9 13 9 1 15 2
5 15 13 0 3 2
5 15 13 3 3 2
5 15 4 13 3 2
7 15 13 0 1 15 3 2
5 9 13 1 9 2
5 13 15 1 9 2
6 13 1 15 1 9 2
5 13 12 9 0 2
6 13 15 1 10 9 2
6 13 15 1 10 9 2
3 2 13 2
5 10 9 13 3 2
4 10 9 13 2
4 2 13 15 2
6 15 13 0 1 15 2
6 15 13 0 1 9 2
6 15 13 0 1 15 2
6 14 15 13 1 15 2
5 0 9 15 13 2
5 0 9 15 13 2
7 9 13 1 9 7 9 2
9 11 13 2 16 15 15 4 13 2
9 11 13 2 16 15 15 4 13 2
5 9 15 14 13 2
8 13 15 2 16 11 14 13 2
8 15 13 10 9 1 15 14 2
8 15 13 10 9 1 15 14 2
11 1 9 1 9 9 15 15 13 3 3 2
11 1 9 15 9 1 9 15 13 3 3 2
11 1 9 15 9 1 9 15 13 3 3 2
5 9 15 13 3 2
6 9 15 14 13 3 2
5 9 15 15 13 2
13 15 13 2 16 11 14 13 7 14 13 1 15 2
14 15 13 2 16 15 6 13 14 11 14 13 14 13 2
7 14 4 13 2 13 3 2
9 0 13 2 16 15 6 13 3 2
7 14 15 13 3 13 3 2
8 16 15 13 3 2 13 3 2
9 13 15 15 2 16 15 13 3 2
8 13 15 9 2 16 4 13 2
10 13 15 15 3 2 16 15 13 3 2
9 16 4 13 2 15 13 1 15 2
6 13 15 15 14 13 2
6 9 15 13 14 13 2
7 10 9 13 2 14 13 2
6 15 13 2 4 13 2
7 15 13 2 13 14 13 2
9 10 9 13 2 13 14 13 15 2
9 1 10 4 15 13 2 4 13 2
6 14 13 2 13 3 2
6 6 13 14 4 13 2
8 15 13 2 16 13 14 13 2
6 14 15 13 14 13 2
6 13 15 14 15 13 2
5 15 13 14 13 2
7 15 16 4 13 15 13 2
6 13 15 14 15 13 2
6 15 13 14 13 3 2
6 15 13 14 13 3 2
6 6 13 14 4 13 2
5 13 15 14 13 2
7 13 15 3 13 1 15 2
7 13 15 14 13 1 15 2
8 13 15 2 16 13 1 15 2
8 13 9 2 16 9 4 13 2
7 13 15 14 13 1 15 2
6 13 14 13 1 15 2
7 13 15 14 13 1 9 2
6 13 9 14 13 9 2
6 3 14 13 10 9 2
9 3 14 13 10 9 14 15 13 2
9 3 14 13 14 15 13 10 9 2
5 13 15 14 13 2
7 11 15 13 14 15 13 2
7 11 15 13 14 15 13 2
9 3 14 13 10 9 14 15 13 2
8 13 15 15 14 15 13 15 2
5 13 15 14 13 2
6 13 15 14 13 9 2
6 13 15 14 15 13 2
6 13 15 2 16 13 2
5 13 15 1 9 2
10 15 13 2 16 15 4 15 13 15 2
7 14 15 13 14 15 13 2
7 13 15 14 15 13 15 2
6 13 2 16 4 13 2
6 13 14 15 13 9 2
8 13 15 1 9 2 16 13 2
6 15 13 3 4 13 2
7 13 1 10 2 16 13 2
8 13 15 3 14 13 1 3 2
5 13 2 15 13 2
6 15 13 2 15 13 2
15 1 15 13 14 9 1 10 9 2 15 14 13 9 15 2
9 15 2 15 13 9 15 2 13 2
10 9 2 15 3 4 13 2 4 13 2
17 15 13 3 9 2 16 15 13 9 1 3 0 1 9 15 9 2
13 9 2 3 14 13 15 2 6 15 13 1 9 2
13 1 10 9 13 10 9 2 3 9 15 15 13 2
10 13 15 9 2 16 15 6 13 3 2
10 10 2 16 4 15 13 2 13 9 2
10 9 2 16 4 13 2 4 13 3 2
10 13 9 14 13 2 10 9 13 3 2
8 15 13 10 2 15 15 13 2
13 15 13 1 9 1 9 2 10 9 15 13 0 2
8 13 9 2 10 6 4 13 2
8 13 9 2 10 9 6 13 2
10 9 2 10 9 13 15 2 13 0 2
12 15 13 15 1 9 2 3 9 15 15 13 2
12 15 13 15 1 9 2 3 9 15 15 13 2
8 15 13 9 2 3 13 15 2
11 9 2 15 3 15 4 13 9 2 13 2
9 13 9 2 15 14 13 1 9 2
8 13 9 2 15 14 15 13 2
10 9 2 15 15 4 13 9 2 13 2
6 15 13 14 15 13 2
11 9 2 15 14 13 15 2 6 15 13 2
9 14 13 9 2 15 14 15 13 2
12 1 10 9 13 9 2 15 14 13 1 9 2
9 13 15 9 2 15 4 13 15 2
6 3 13 14 15 13 2
6 3 13 14 15 13 2
10 15 14 15 13 9 2 3 14 13 2
7 9 15 14 13 13 0 2
5 13 10 14 13 2
6 13 15 15 14 13 2
6 13 15 15 14 13 2
5 13 10 14 13 2
6 13 15 14 15 13 2
11 14 13 1 15 2 3 16 15 13 15 2
8 6 13 0 2 1 14 13 2
10 14 13 1 15 2 16 15 13 15 2
10 14 13 1 15 2 16 15 13 15 2
10 14 13 1 15 2 3 15 13 15 2
10 14 13 1 15 2 3 15 13 15 2
8 14 15 13 2 1 1 13 2
8 14 15 13 2 1 14 13 2
8 15 13 3 14 6 15 13 2
7 15 13 2 1 16 13 2
7 14 15 13 2 3 13 2
10 15 13 3 2 1 14 6 15 13 2
10 13 15 1 15 3 2 3 15 13 2
7 4 15 13 2 16 13 2
10 15 14 15 13 2 7 14 6 13 2
10 15 15 13 2 15 7 14 15 13 2
8 15 13 2 1 14 15 13 2
9 15 15 13 3 3 15 13 9 2
10 15 13 3 2 3 16 14 15 13 2
7 13 2 1 14 15 13 2
10 15 13 3 3 2 16 15 15 13 2
9 14 15 13 2 3 7 14 13 2
6 13 14 13 1 15 2
6 16 6 13 2 13 2
8 15 13 3 2 16 13 15 2
5 16 13 2 13 2
7 14 13 2 3 15 13 2
8 6 15 13 2 3 4 13 2
6 13 2 16 15 13 2
6 13 2 3 15 13 2
9 15 13 2 3 15 7 14 13 2
7 13 2 1 15 14 13 2
9 15 13 2 3 16 6 15 13 2
7 13 14 13 15 1 9 2
10 15 15 13 14 15 13 14 13 9 2
8 15 15 13 2 1 14 13 2
9 15 13 2 1 14 15 13 9 2
7 13 14 13 14 13 9 2
8 15 13 9 15 14 13 9 2
6 13 14 15 13 15 2
9 15 13 9 15 1 14 13 9 2
8 1 14 15 13 2 13 15 2
13 14 13 3 2 1 14 13 9 1 1 12 9 2
10 15 13 3 9 2 3 15 13 9 2
12 14 15 13 1 15 2 15 7 14 13 15 2
7 15 13 2 1 16 13 2
9 14 13 2 15 7 14 13 15 2
9 15 15 13 2 3 14 15 13 2
10 15 13 3 9 2 3 15 13 9 2
12 15 14 15 13 2 10 9 7 14 15 13 2
12 15 14 15 13 2 10 7 9 14 15 13 2
6 3 15 13 2 13 2
6 3 15 13 2 13 2
6 3 13 2 15 13 2
6 3 13 2 15 13 2
5 15 13 7 13 2
9 9 2 16 15 13 2 15 13 2
8 9 2 16 13 2 15 13 2
8 9 2 16 13 2 15 13 2
9 16 15 13 2 15 13 14 13 2
6 3 15 13 1 15 2
6 9 15 13 1 15 2
7 3 4 13 9 1 9 2
5 13 14 15 15 2
4 13 14 9 2
4 2 13 4 2
8 13 15 14 15 15 13 9 2
5 10 9 15 13 2
7 13 15 14 15 13 9 2
8 10 9 15 13 14 15 13 2
7 6 13 14 6 4 13 2
5 3 15 13 3 2
10 13 14 4 13 2 1 14 15 13 2
6 6 15 13 1 9 2
6 15 3 15 15 13 2
5 13 15 15 9 2
8 15 3 15 13 3 13 0 2
7 1 9 6 15 13 9 2
5 13 15 15 15 2
6 1 9 6 15 13 2
9 16 15 14 13 3 2 13 3 2
7 13 15 2 16 14 13 2
5 13 14 15 13 2
6 13 15 15 14 13 2
5 13 15 0 9 2
6 13 15 15 0 9 2
6 3 15 13 0 9 2
7 13 15 14 15 13 3 2
7 15 13 14 15 13 3 2
6 3 13 14 15 13 2
6 13 15 14 13 3 2
9 9 1 15 14 6 15 15 13 2
7 13 14 11 13 14 4 2
5 3 4 13 11 2
7 2 11 14 3 4 13 2
8 13 14 4 9 15 11 3 2
7 9 14 1 9 4 13 2
6 9 1 9 14 13 2
5 6 4 15 13 2
5 9 15 14 13 2
5 9 14 15 13 2
5 15 13 3 14 2
6 6 9 14 13 15 2
6 9 14 6 13 15 2
5 6 15 14 13 2
5 6 13 14 15 2
7 15 6 13 3 1 15 2
5 15 13 1 15 2
5 15 15 14 13 2
6 15 13 14 15 13 2
9 15 13 2 16 11 13 14 13 2
8 15 13 2 16 15 4 13 2
7 15 16 4 13 15 13 2
6 15 3 13 14 13 2
6 15 3 13 14 13 2
5 15 15 14 13 2
7 15 13 2 16 15 13 2
5 15 10 9 13 2
6 11 13 14 4 13 2
7 15 15 13 14 4 13 2
7 11 13 2 16 13 3 2
7 13 2 16 15 13 0 2
5 15 13 13 0 2
7 15 13 2 16 13 0 2
10 15 13 2 7 4 3 13 1 9 2
9 15 13 2 7 9 15 13 3 2
8 9 13 2 16 9 4 13 2
8 9 13 2 16 4 13 9 2
7 9 13 2 16 4 13 2
7 13 2 16 9 4 13 2
9 13 15 2 16 9 14 13 0 2
6 11 13 3 14 13 2
9 15 13 15 2 7 6 13 10 2
10 9 2 16 14 13 0 2 15 13 2
6 11 13 3 14 13 2
6 11 4 13 14 13 2
6 9 15 13 9 15 2
7 1 11 0 0 9 13 2
6 13 15 0 0 9 2
5 15 15 13 9 2
5 15 15 13 9 2
8 16 13 0 2 15 13 9 2
12 13 15 0 15 9 2 7 15 6 15 13 2
8 15 15 13 9 1 9 15 2
6 13 15 10 15 9 2
9 15 15 13 9 15 1 9 15 2
5 13 15 9 15 2
5 13 15 9 15 2
5 13 15 9 15 2
6 15 4 15 15 13 2
5 15 15 6 13 2
9 15 13 1 12 9 9 10 9 2
8 9 15 15 4 13 10 9 2
6 15 15 15 4 13 2
5 15 15 6 13 2
6 15 15 15 4 13 2
9 1 12 9 9 15 13 10 9 2
5 15 13 10 9 2
5 2 15 13 15 2
7 13 15 3 9 1 9 2
6 13 15 9 1 9 2
5 9 3 4 13 2
6 13 15 14 15 13 2
8 11 13 9 1 14 15 13 2
6 11 13 9 14 13 2
6 11 13 14 13 9 2
5 9 15 13 9 2
4 6 13 15 2
12 7 9 2 7 9 2 14 7 9 6 13 2
18 3 13 9 7 13 9 2 7 15 13 1 9 7 15 13 14 13 2
7 15 13 1 9 7 9 2
8 9 15 1 9 3 4 13 2
37 3 1 11 13 0 9 1 9 1 9 1 9 1 9 1 9 1 0 11 2 0 1 0 9 1 9 1 9 2 9 2 0 9 7 0 9 2
18 12 9 13 1 15 1 9 7 15 13 1 9 15 7 3 0 9 2
12 13 3 1 15 2 9 2 9 1 9 11 2
20 16 13 14 13 9 1 0 11 2 13 13 13 14 13 0 1 9 7 9 2
10 0 15 9 1 9 15 13 3 3 2
48 1 9 7 9 1 9 9 1 9 1 0 9 1 11 2 0 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 0 9 7 11 13 0 9 1 0 9 7 13 9 7 9 2
11 9 11 4 13 7 9 0 9 1 11 2
11 3 9 11 13 14 13 9 15 1 11 2
11 3 9 11 13 14 13 9 15 1 11 2
19 7 14 15 13 2 7 14 15 13 1 0 9 2 16 15 13 3 9 2
9 15 13 0 9 1 9 1 11 2
15 7 16 9 13 0 9 7 9 2 9 15 13 0 9 2
8 10 9 3 13 0 1 9 2
12 3 7 9 1 9 1 9 15 13 3 0 2
11 3 2 15 6 13 0 7 6 13 9 2
4 13 0 9 2
7 9 13 3 0 7 0 2
4 0 13 15 2
14 1 10 9 4 13 9 1 9 1 0 9 1 9 2
7 14 15 13 15 14 13 2
11 7 10 9 6 13 7 0 2 7 0 2
7 15 6 13 10 0 9 2
22 10 9 1 11 13 0 9 7 0 9 1 10 9 2 1 12 1 9 1 0 9 2
33 0 9 2 15 6 4 13 14 13 9 1 9 1 9 1 0 9 2 0 1 0 0 7 0 9 1 11 2 9 1 0 9 2
23 15 13 0 15 9 7 13 0 0 9 2 15 13 0 9 1 9 15 2 13 15 3 2
8 12 9 4 13 1 9 15 2
21 15 13 7 9 15 2 15 15 13 14 13 1 9 15 2 7 9 3 15 13 2
11 0 15 13 14 13 0 9 1 9 15 2
31 1 10 9 0 0 9 4 13 3 0 9 1 9 1 0 1 15 0 9 1 9 1 9 7 9 1 0 9 1 11 2
28 9 15 9 11 2 13 3 1 9 1 11 2 13 15 2 1 0 9 2 1 9 1 9 2 13 7 13 2
16 13 3 1 0 9 2 3 3 15 4 3 13 1 9 15 2
16 1 1 13 3 0 2 0 7 0 0 9 2 9 13 3 2
23 6 3 13 9 1 9 1 9 1 12 9 2 7 13 9 1 9 1 3 0 0 9 2
15 13 15 9 2 13 9 2 13 15 9 2 13 0 9 2
11 7 15 6 15 13 14 13 14 15 13 2
10 13 15 2 16 13 14 13 1 11 2
11 13 4 9 9 1 12 9 14 13 0 2
14 0 9 14 15 13 1 11 1 0 9 1 10 9 2
10 13 0 9 2 7 13 12 0 9 2
12 15 6 13 0 2 7 7 15 6 13 9 2
12 15 6 13 0 2 7 7 15 6 13 9 2
15 10 9 3 13 3 0 9 7 10 0 9 13 9 15 2
13 13 14 3 3 11 14 4 13 1 10 0 9 2
10 13 15 3 1 0 0 7 0 9 2
30 1 9 1 0 9 1 0 9 1 0 15 9 2 9 13 9 1 9 1 0 1 9 9 1 9 1 9 1 9 2
15 1 9 13 3 1 0 9 7 9 1 0 9 15 13 2
14 1 16 4 13 2 9 1 0 11 3 6 4 13 2
13 3 9 14 13 1 0 9 1 9 2 13 11 2
22 11 13 9 1 9 2 1 15 9 1 0 9 15 13 2 1 14 13 0 15 9 2
22 0 11 4 13 1 9 2 1 15 13 0 9 1 9 1 9 1 9 1 0 9 2
15 0 1 9 15 2 11 3 13 9 7 15 13 1 15 2
16 13 9 1 0 9 1 11 7 1 0 9 1 0 9 11 2
20 11 13 11 2 15 4 13 1 0 9 1 9 15 2 7 15 13 1 9 2
13 15 13 3 1 15 7 3 15 13 1 15 14 2
7 1 9 1 9 13 9 2
5 9 13 1 9 2
11 13 14 15 10 0 0 9 13 1 9 2
11 13 14 15 10 0 0 9 13 1 9 2
13 3 3 13 9 2 7 0 9 6 15 13 0 2
21 7 15 6 13 2 16 10 0 9 7 0 9 1 9 1 0 9 13 0 9 2
15 0 9 6 13 7 15 13 1 9 2 14 13 9 15 2
17 13 15 14 6 15 13 1 9 15 2 7 15 7 13 10 9 2
6 6 13 7 6 13 2
23 13 1 9 2 13 15 1 9 1 9 1 11 7 1 0 1 0 9 9 13 1 9 2
22 15 13 3 3 2 3 2 3 3 15 4 13 7 15 13 1 9 2 9 13 3 2
23 10 1 0 9 1 0 9 13 0 1 0 9 2 15 13 14 13 9 1 9 1 9 2
26 1 15 2 3 2 13 9 1 0 9 2 1 15 0 0 9 14 15 13 1 0 2 3 0 9 2
13 6 15 13 7 0 9 1 9 2 7 0 9 2
11 11 11 4 13 3 3 7 13 0 9 2
12 1 9 7 1 12 9 1 9 13 0 9 2
21 3 13 3 14 15 13 1 9 10 4 13 0 7 4 13 1 9 1 0 9 2
18 9 2 15 13 9 1 10 9 2 13 9 1 9 15 1 1 9 2
5 9 13 0 9 2
13 9 2 9 2 9 2 0 9 2 9 2 9 2
14 1 9 1 9 12 9 13 0 9 1 0 7 0 2
20 9 1 11 7 11 13 9 1 9 1 0 9 14 15 13 1 9 1 11 2
14 6 13 9 1 9 7 9 2 15 14 13 10 9 2
17 13 15 3 1 0 9 2 3 14 15 13 10 0 9 1 9 2
10 7 3 3 6 15 13 7 1 15 2
20 1 9 2 15 13 2 0 0 9 13 11 14 13 11 1 9 1 0 9 2
18 13 15 0 0 9 1 9 0 9 1 9 7 9 1 3 0 9 2
3 9 13 2
11 13 9 14 15 13 1 9 0 10 9 2
17 9 1 0 9 1 9 1 0 15 9 1 9 11 13 3 0 2
9 13 9 15 7 3 13 1 11 2
16 15 3 13 14 13 10 0 0 9 1 11 1 9 1 11 2
18 0 9 13 2 16 1 10 9 6 13 0 9 1 9 1 9 11 2
15 3 13 2 16 11 4 13 6 3 9 1 0 15 9 2
11 1 9 1 0 9 4 13 9 1 11 2
15 6 2 7 1 9 1 11 3 15 13 1 9 1 9 2
19 1 9 15 13 9 1 9 1 9 1 0 9 7 9 1 0 15 9 2
16 2 9 1 9 13 14 9 1 11 7 0 11 7 0 9 2
11 11 13 2 7 9 1 15 3 13 9 2
17 9 13 3 2 16 3 3 9 3 13 9 1 11 1 0 9 2
7 15 3 15 13 1 9 2
11 15 13 9 15 2 15 15 3 14 13 2
13 15 6 13 14 6 15 13 1 3 0 15 9 2
19 1 9 1 0 9 1 9 1 0 9 1 9 4 13 9 1 9 11 2
16 7 0 9 1 11 13 2 16 9 1 0 9 6 13 0 2
15 9 1 0 9 13 0 1 9 7 9 0 9 1 9 2
13 3 0 0 9 14 13 3 1 9 1 0 9 2
14 13 14 15 0 9 7 14 13 14 0 9 1 9 2
9 14 3 13 9 1 11 1 11 2
30 1 0 9 0 9 1 0 9 4 13 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
14 2 1 9 4 13 9 1 9 1 9 1 11 11 2
8 11 6 13 14 13 9 15 2
9 11 15 15 13 1 0 15 9 2
16 15 3 4 3 13 1 9 1 9 1 11 2 11 2 11 2
12 0 9 1 0 9 13 1 9 1 0 9 2
9 3 14 13 14 13 9 1 11 2
14 15 4 13 14 13 0 0 9 1 0 9 1 11 2
8 11 13 9 7 13 1 15 2
8 11 13 9 7 13 1 15 2
5 12 9 15 13 2
12 1 0 9 13 7 9 1 0 9 11 11 2
12 11 11 13 9 1 0 9 1 9 1 11 2
11 2 7 1 10 9 11 3 15 13 15 2
8 10 9 11 6 13 14 13 2
13 13 9 1 9 11 11 1 0 9 1 0 9 2
12 1 0 9 4 13 7 0 9 1 9 11 2
14 3 3 15 14 13 9 1 9 7 1 12 15 9 2
4 1 10 9 2
33 7 14 13 12 9 7 2 14 13 1 0 9 2 7 14 13 10 14 14 9 2 10 9 13 9 11 2 13 9 2 13 9 2
6 14 14 15 13 0 2
35 1 0 4 13 9 1 9 1 9 1 9 1 9 1 9 2 9 7 9 1 9 7 9 1 0 9 14 13 9 1 9 1 10 9 2
11 13 14 10 9 7 3 15 13 10 9 2
18 1 9 1 9 7 0 9 13 10 9 2 1 15 15 13 0 9 2
5 9 1 9 13 2
9 9 1 9 13 0 7 3 0 2
6 3 13 9 1 9 2
10 13 15 1 9 7 15 13 3 3 2
9 6 2 3 13 9 2 0 9 2
7 7 3 13 7 3 9 2
17 7 10 2 15 15 13 1 9 2 13 14 13 9 1 10 9 2
11 7 15 13 3 1 0 9 1 10 9 2
23 1 9 1 9 15 4 13 0 0 0 9 1 9 1 9 1 0 9 14 13 3 9 2
19 3 14 13 9 1 0 9 1 9 2 15 3 13 14 13 2 13 9 2
12 9 1 0 9 1 0 9 14 13 0 9 2
24 15 13 0 1 9 2 7 1 9 15 4 13 3 1 9 2 15 4 13 2 0 7 0 2
16 9 3 14 4 13 7 1 10 0 9 2 15 3 15 13 2
42 3 1 0 9 1 9 1 0 9 2 1 9 1 9 1 9 1 9 7 9 1 0 9 7 1 10 9 13 7 13 14 15 13 9 2 9 7 9 1 10 9 2
11 1 15 4 13 9 1 9 1 0 9 2
45 0 4 13 1 9 1 0 9 1 0 9 1 9 1 9 7 9 15 1 9 1 9 1 0 9 2 9 1 10 9 1 9 1 0 9 1 9 7 9 1 9 1 0 9 2
18 0 9 1 9 1 9 1 9 13 9 9 2 9 2 9 2 9 2
19 13 15 0 9 2 0 9 2 1 10 0 9 2 9 1 9 1 9 2
9 3 13 2 16 9 6 13 0 2
26 13 15 4 1 9 7 9 15 9 11 7 6 3 15 6 13 2 7 4 13 7 14 15 6 13 2
27 1 10 9 0 9 14 13 9 1 9 1 9 7 0 9 3 1 0 1 10 0 9 9 1 0 9 2
27 1 9 9 1 12 9 13 9 1 9 1 11 7 13 9 1 10 9 14 13 1 9 7 9 1 9 2
18 3 15 13 1 9 1 9 15 2 3 9 15 13 2 16 13 0 2
13 3 1 9 9 15 13 1 0 1 9 1 9 2
17 1 9 13 0 0 9 2 1 15 15 13 9 1 0 0 9 2
12 1 9 9 13 2 3 14 13 3 12 9 2
16 9 1 9 13 0 2 15 13 7 15 13 1 9 1 9 2
47 9 1 9 14 15 13 1 9 9 7 9 1 0 9 7 9 2 9 1 9 7 9 1 0 9 7 9 2 7 9 14 4 13 1 9 9 7 9 1 0 9 7 9 1 0 9 2
6 13 15 3 7 3 2
23 1 15 9 1 10 0 9 1 9 13 3 12 14 15 13 9 2 1 14 13 1 9 2
11 6 13 14 2 1 10 9 13 3 9 2
12 16 15 13 2 13 2 13 7 15 15 13 2
14 3 0 2 15 0 9 13 1 9 2 13 14 13 2
20 1 9 1 9 1 0 9 1 9 1 9 2 1 0 9 4 13 0 9 2
17 16 13 2 13 2 16 15 13 2 7 13 9 2 13 7 13 2
12 2 3 13 9 1 9 1 9 1 0 9 2
22 3 14 13 2 16 1 9 1 9 1 9 14 15 13 9 1 9 1 9 1 9 2
6 13 9 1 10 9 2
17 16 13 0 9 1 9 1 0 9 2 9 1 10 9 13 0 2
13 3 16 9 1 9 1 9 13 9 1 10 9 2
22 1 9 1 10 9 0 9 1 9 1 9 14 13 9 1 9 1 9 1 10 9 2
16 0 7 0 13 9 1 9 7 9 1 0 9 1 10 9 2
30 9 1 0 9 1 0 9 13 1 0 0 9 2 13 7 13 9 1 9 2 9 1 9 7 9 1 0 0 9 2
19 15 13 3 9 1 9 1 9 7 0 9 1 0 0 9 1 10 9 2
12 14 13 14 10 9 9 3 1 0 15 9 2
5 15 6 13 9 2
24 3 15 13 2 1 0 9 2 1 0 9 9 1 0 9 2 1 14 13 9 2 13 9 2
10 15 15 13 1 10 7 14 13 9 2
11 3 9 7 9 6 15 13 9 14 13 2
3 13 9 2
22 7 3 13 9 14 13 2 16 0 9 7 0 1 0 9 13 14 13 3 1 9 2
21 9 13 3 3 14 13 9 1 0 9 2 13 14 13 1 0 0 7 0 9 2
15 15 13 0 9 1 9 1 9 1 9 2 13 0 9 2
8 1 9 14 13 9 1 9 2
12 1 9 4 13 2 16 3 9 13 14 13 2
9 3 0 9 14 13 9 1 9 2
21 1 9 4 13 15 2 7 1 9 15 3 13 1 15 2 3 1 9 1 9 2
15 15 13 2 16 15 4 13 0 9 1 9 1 10 9 2
42 1 9 1 0 9 15 13 9 7 9 1 0 9 2 13 15 9 1 9 1 9 2 13 15 9 1 9 7 15 13 9 1 0 0 9 1 9 1 9 1 9 2
13 9 13 2 16 15 14 13 0 9 1 10 9 2
4 15 4 13 2
14 13 4 10 0 9 2 13 4 0 9 1 10 9 2
36 7 15 3 15 15 13 2 13 3 9 1 0 15 9 7 13 10 2 15 1 0 15 9 13 14 15 13 1 9 2 16 3 13 1 9 2
20 1 9 1 0 9 0 7 0 9 1 9 14 13 9 1 9 1 0 9 2
37 2 0 0 9 2 3 1 9 1 0 9 7 9 2 3 7 1 0 9 2 1 15 1 9 1 0 0 9 2 0 9 4 13 10 0 9 2
22 13 15 14 13 9 1 9 1 9 1 0 9 2 16 15 14 15 13 1 0 9 2
14 15 14 13 3 9 7 9 1 0 9 1 10 9 2
7 13 15 7 13 1 9 2
17 1 15 9 1 9 1 0 13 7 15 3 15 13 1 9 15 2
20 11 2 0 1 9 7 9 1 9 2 15 13 3 1 9 7 13 9 15 2
17 13 9 1 9 1 15 14 13 7 6 13 10 9 1 10 9 2
43 9 1 9 1 10 9 14 15 13 1 9 1 9 7 9 1 9 7 10 0 9 2 3 7 1 9 1 0 9 1 9 1 9 1 9 1 9 7 1 9 1 9 2
2 9 2
3 13 3 2
22 13 2 13 2 13 15 9 2 13 9 7 9 13 3 0 2 7 6 13 3 9 2
26 7 0 1 15 9 7 9 15 13 2 16 9 7 9 13 3 2 3 9 1 9 2 9 7 9 2
35 13 4 0 9 1 9 1 9 1 9 1 0 9 2 1 9 1 0 9 1 9 7 9 1 0 9 7 0 9 1 9 1 0 9 2
13 9 13 3 3 2 7 1 9 15 13 1 9 2
28 3 15 13 0 0 9 2 13 15 7 3 3 3 1 9 2 3 3 13 3 9 2 1 14 13 1 15 2
18 0 9 13 14 4 13 1 9 3 3 9 13 9 1 9 1 9 2
12 1 10 9 14 13 0 9 1 10 0 9 2
26 0 9 2 0 1 9 1 0 9 2 15 13 1 9 1 0 9 2 15 13 0 9 1 0 9 2
13 3 13 9 2 7 6 15 15 13 1 0 9 2
27 7 3 15 15 13 1 9 1 10 0 9 2 3 14 15 13 2 16 1 10 9 1 0 9 13 9 2
16 0 9 1 9 13 9 1 0 9 2 16 13 9 0 9 2
17 3 15 14 13 9 1 9 2 15 13 14 13 9 1 0 9 2
8 9 13 14 13 1 0 9 2
26 3 3 2 16 13 9 10 0 9 14 15 13 6 1 9 1 0 9 2 7 1 9 1 0 9 2
23 3 3 0 0 9 13 9 1 0 9 2 9 1 0 7 0 9 1 10 9 1 9 2
5 3 15 13 15 2
21 1 9 13 9 2 15 13 1 0 9 2 7 15 13 3 0 2 13 1 9 2
12 7 16 13 9 1 9 2 15 13 7 13 2
11 1 14 13 9 2 13 7 13 1 9 2
46 1 9 9 1 0 9 13 9 2 16 9 1 0 9 1 0 9 1 9 1 0 9 14 13 0 9 1 0 1 10 9 9 7 0 9 1 9 1 0 15 9 1 9 1 11 2
17 3 3 0 9 13 1 9 1 0 9 2 15 4 13 0 9 2
29 9 3 15 13 1 15 1 9 2 1 15 1 1 9 1 9 1 9 15 13 7 1 0 9 7 0 0 9 2
11 1 9 1 9 15 15 13 1 1 9 2
24 14 13 12 9 1 12 9 1 9 1 9 2 1 15 4 13 1 9 1 0 7 0 9 2
24 14 13 12 9 1 12 9 1 9 1 9 2 1 15 4 13 1 9 1 0 7 0 9 2
28 2 0 9 1 9 1 9 15 13 3 1 9 1 0 9 7 9 1 9 1 9 1 0 9 1 0 9 2
12 0 9 13 1 9 1 9 1 9 1 9 2
11 0 9 1 9 4 13 1 9 1 9 2
9 0 4 13 7 13 14 4 13 2
18 2 15 13 3 2 15 13 1 11 7 3 13 0 9 1 10 9 2
20 1 0 9 3 13 9 1 9 1 0 9 1 9 7 9 1 9 1 9 2
33 1 0 9 13 3 2 16 9 1 11 2 0 0 9 1 0 9 1 0 11 2 13 14 13 0 9 1 9 7 9 1 11 2
22 9 1 11 13 9 2 16 3 4 13 9 1 0 9 1 0 9 1 11 1 11 2
12 3 0 0 9 1 11 15 13 1 3 0 2
23 3 13 0 9 1 0 9 1 0 2 0 7 0 2 15 14 6 13 1 9 1 9 2
4 3 0 13 2
29 10 0 9 15 13 1 9 1 10 9 9 2 15 3 13 0 6 3 1 11 7 11 2 7 4 13 0 9 2
22 3 13 2 16 4 13 1 11 2 13 14 14 13 1 9 2 10 4 13 1 15 2
13 9 1 9 1 0 9 2 9 1 9 1 11 2
11 15 13 9 1 0 9 2 9 7 9 2
5 1 0 7 0 2
2 9 2
17 1 10 9 15 13 7 13 1 9 2 1 15 13 9 1 11 2
14 3 13 14 4 13 1 14 15 13 0 9 1 11 2
14 1 10 9 1 9 1 11 4 13 9 1 9 9 2
19 3 0 13 9 1 9 1 0 9 1 11 1 9 1 0 9 1 11 2
24 1 0 0 9 9 1 0 9 11 11 13 9 1 9 1 9 1 9 1 0 9 1 11 2
7 1 10 9 15 15 13 2
12 15 13 9 15 1 0 9 2 3 15 13 2
5 3 3 2 3 2
30 9 7 9 1 9 2 15 15 13 1 9 1 0 9 2 9 1 9 7 0 9 2 9 1 0 9 1 0 9 2
7 13 0 1 11 0 9 2
24 10 10 9 13 1 0 9 1 9 7 0 9 2 15 15 13 3 1 0 9 7 0 9 2
7 7 12 0 9 1 9 2
11 15 4 13 3 0 9 1 0 0 9 2
11 0 7 0 13 9 1 0 9 7 9 2
8 3 13 3 0 9 1 11 2
9 1 0 9 1 11 13 0 9 2
8 0 15 9 13 1 9 0 2
9 1 0 9 9 13 9 11 11 2
10 1 10 9 1 9 13 3 0 9 2
9 1 0 0 9 14 15 13 9 2
4 13 12 9 2
8 13 11 1 0 9 1 9 2
10 3 13 0 9 1 11 1 0 9 2
7 13 15 2 13 2 9 2
5 0 9 1 9 2
15 14 13 14 13 12 9 2 7 15 3 13 1 0 9 2
16 7 13 14 9 1 9 1 9 9 1 9 2 3 15 13 2
16 2 13 9 1 9 7 9 1 9 1 9 1 9 1 9 2
18 10 0 9 13 14 13 9 1 0 9 3 2 1 10 10 0 9 2
2 13 2
6 2 9 3 15 13 2
5 9 3 15 13 2
4 9 13 0 2
6 7 0 9 15 13 2
7 7 14 13 14 15 13 2
23 14 3 6 15 15 13 14 13 9 15 1 9 2 16 15 13 9 7 13 9 1 9 2
19 3 3 13 9 1 10 9 1 10 0 11 7 0 9 1 9 1 15 2
12 10 9 2 10 9 6 13 14 4 13 3 2
8 7 10 9 6 13 1 3 2
4 15 13 0 2
20 15 13 9 1 0 9 1 9 2 9 15 13 1 15 3 16 13 1 9 2
19 9 15 15 13 7 3 13 14 13 2 16 13 3 3 14 13 3 0 2
26 0 15 13 2 7 1 16 15 13 2 13 0 7 15 13 3 1 15 2 16 9 13 1 0 9 2
17 2 3 13 9 1 0 9 14 4 13 1 0 15 1 0 9 2
7 15 14 13 10 0 9 2
29 7 13 15 14 15 13 2 16 15 3 6 15 13 2 15 13 2 16 15 13 3 0 1 9 1 0 15 9 2
16 7 15 14 13 1 10 9 1 10 0 9 1 9 1 9 2
42 1 9 7 9 1 0 9 1 9 7 9 1 9 1 9 7 0 9 6 13 0 0 15 7 0 9 1 0 9 3 1 9 1 9 2 3 7 1 0 0 9 2
22 6 13 1 9 7 9 2 16 1 0 9 1 9 15 13 9 1 0 9 1 9 2
22 7 0 0 9 2 15 13 9 1 0 9 2 10 13 0 0 9 1 9 7 9 2
23 1 11 3 3 15 13 10 9 1 9 1 10 0 9 2 9 1 0 9 1 0 9 2
16 15 13 9 2 15 14 13 9 1 9 2 15 11 14 13 2
36 0 0 9 13 14 13 10 9 2 16 13 9 1 0 9 1 9 2 9 7 9 1 9 2 1 9 1 9 1 0 0 9 1 0 9 2
5 3 14 15 13 2
29 1 9 1 10 2 15 15 13 1 9 1 9 1 9 7 9 1 9 2 15 4 13 14 15 13 1 12 9 2
22 7 3 15 13 1 9 0 9 1 0 9 7 10 9 15 13 1 10 7 0 9 2
12 0 9 1 9 1 9 7 0 9 14 13 2
8 15 13 9 1 9 11 11 2
11 1 10 9 14 15 13 3 1 0 9 2
9 1 15 9 13 14 15 13 3 2
5 1 9 1 9 2
21 6 13 15 13 2 14 13 12 9 7 1 10 9 14 13 2 13 9 1 9 2
26 13 9 2 16 9 1 11 13 3 1 9 1 0 9 7 13 3 0 9 1 9 1 0 15 9 2
24 15 13 0 7 0 0 9 2 0 9 1 9 1 9 2 0 9 7 0 9 1 0 9 2
27 10 9 13 2 16 0 9 13 10 0 9 1 3 0 9 7 15 13 14 13 7 13 9 15 1 9 2
13 1 10 9 15 13 0 7 0 9 1 0 9 2
14 0 9 13 14 15 13 9 2 1 15 13 0 9 2
6 12 9 3 15 13 2
9 6 13 9 1 0 9 1 9 2
39 15 15 13 3 2 3 1 10 0 9 2 0 15 13 1 9 2 7 1 0 9 15 13 9 15 3 1 9 7 3 15 15 13 2 9 15 4 13 2
20 13 15 0 0 9 1 9 1 0 9 14 13 3 14 13 0 9 1 15 2
8 13 14 13 3 9 1 9 2
10 3 3 13 14 15 13 9 1 9 2
23 15 2 13 2 14 13 0 9 2 7 14 13 14 15 13 1 0 9 2 0 15 9 2
19 9 13 3 7 15 13 2 16 1 3 9 13 1 0 9 1 10 9 2
10 7 13 3 3 0 13 1 9 15 2
17 1 11 3 13 2 16 0 15 9 15 13 3 2 3 7 3 2
22 9 3 13 2 16 1 10 9 13 9 2 7 15 3 15 13 1 9 1 0 9 2
12 9 13 0 9 1 9 1 9 1 0 9 2
21 3 13 2 16 1 15 15 13 0 9 2 1 14 13 10 0 9 1 0 9 2
40 0 9 2 0 1 0 9 1 0 0 9 2 13 9 1 0 9 1 0 9 1 9 1 0 9 1 0 9 7 1 0 9 1 9 1 9 1 0 11 2
30 7 1 9 1 9 1 0 9 7 9 1 0 9 15 13 14 13 1 0 9 2 3 1 15 15 13 1 0 9 2
22 0 9 1 9 1 0 0 9 1 9 1 9 13 1 9 1 9 15 1 0 9 2
10 15 13 9 2 16 15 13 0 9 2
12 2 13 2 16 1 10 9 15 13 0 9 2
15 3 13 9 2 13 4 15 1 15 7 6 13 1 15 2
21 9 13 14 13 0 9 2 1 14 15 13 9 1 9 2 15 9 3 4 13 2
17 0 9 15 13 7 1 3 0 9 3 1 9 3 7 1 9 2
8 2 6 2 9 2 10 9 2
3 13 4 2
4 13 12 9 2
4 15 6 13 2
7 2 3 13 14 13 9 2
9 2 13 14 15 2 2 13 15 2
9 2 13 14 15 2 2 13 15 2
8 2 1 15 13 2 13 15 2
3 3 3 2
7 13 15 3 2 9 9 2
7 13 15 2 0 9 9 2
7 2 3 4 13 10 9 2
7 3 6 13 1 9 3 2
8 13 9 2 13 9 7 13 2
8 3 2 3 3 14 14 13 2
7 14 13 14 9 1 9 2
7 15 3 13 14 15 13 2
7 13 14 3 14 13 9 2
5 15 13 13 13 2
8 13 11 2 13 15 1 9 2
9 2 13 14 15 13 2 13 15 2
8 2 10 13 1 9 1 9 2
7 9 6 13 14 13 15 2
7 13 15 1 9 1 9 2
8 15 6 13 2 7 13 9 2
7 15 6 15 13 1 15 2
7 0 15 9 6 13 9 2
4 3 13 9 2
7 7 15 13 1 9 15 2
7 13 9 1 10 12 9 2
8 14 2 15 6 13 14 13 2
7 12 9 1 9 1 9 2
7 11 15 13 10 0 9 2
8 2 10 9 4 13 1 9 2
8 2 9 1 0 9 3 13 2
8 2 3 14 15 13 0 9 2
7 15 13 9 1 0 9 2
7 15 13 1 9 1 9 2
7 1 10 9 13 14 15 2
7 13 14 9 1 0 9 2
7 13 14 9 1 0 9 2
7 9 3 13 1 9 15 2
6 13 2 15 6 13 2
3 13 9 2
7 9 11 15 13 1 9 2
7 13 14 15 1 10 9 2
8 13 2 16 3 13 1 9 2
7 13 12 7 0 0 9 2
7 0 1 0 9 6 13 2
7 10 9 1 9 1 9 2
7 3 9 13 1 0 9 2
7 9 3 15 13 1 9 2
8 7 9 15 13 7 6 13 2
8 9 3 6 13 9 1 9 2
8 11 3 15 13 1 9 15 2
8 15 6 13 9 1 0 9 2
8 15 13 14 13 9 1 15 2
6 13 2 16 13 0 2
4 3 13 15 2
7 13 14 15 1 12 9 2
2 13 2
8 15 6 13 7 10 15 9 2
8 15 14 13 9 1 9 15 2
10 15 2 6 2 15 13 7 1 9 2
8 9 15 13 1 9 1 9 2
8 1 10 9 3 9 13 9 2
8 13 15 7 13 3 1 9 2
8 1 9 13 1 9 1 9 2
8 7 3 12 9 13 1 15 2
9 9 13 3 0 2 3 13 15 2
9 2 14 13 14 3 9 14 13 2
9 2 3 14 13 9 1 0 9 2
9 2 10 9 14 4 13 1 9 2
9 2 3 9 14 15 13 1 9 2
10 2 0 9 2 15 13 9 1 9 2
9 3 2 7 14 13 9 1 9 2
3 13 9 2
8 10 10 9 13 0 1 9 2
8 9 1 0 15 1 9 13 2
8 9 1 0 9 1 0 9 2
8 1 10 9 13 14 13 9 2
8 9 1 9 7 9 1 9 2
8 9 3 15 13 1 9 15 2
7 13 14 15 1 10 9 2
2 13 2
3 13 15 2
9 2 15 13 3 0 9 1 9 2
9 2 3 13 9 1 9 1 9 2
9 2 13 7 0 9 1 0 9 2
9 2 13 14 0 9 1 9 15 2
5 15 13 0 9 2
4 3 13 9 2
8 0 9 14 14 13 0 9 2
9 7 1 3 0 9 2 3 3 2
9 13 2 13 9 1 9 11 11 2
9 2 3 3 13 9 1 10 9 2
9 2 9 1 9 1 0 0 9 2
3 13 9 2
6 11 15 13 1 9 2
9 14 13 14 3 9 1 0 9 2
9 3 0 13 7 13 0 1 9 2
9 7 4 13 1 15 14 13 9 2
9 7 15 3 13 9 1 9 15 2
9 14 13 14 9 7 9 1 9 2
9 9 15 13 14 13 7 1 9 2
9 3 15 13 15 1 0 15 9 2
9 7 1 10 6 13 0 15 9 2
9 1 9 1 9 1 9 1 9 2
10 15 15 13 3 2 3 15 15 13 2
5 9 13 1 9 2
5 13 14 13 9 2
8 15 13 14 13 15 1 9 2
2 13 2
9 3 3 13 9 15 1 10 9 2
9 7 15 13 1 0 14 15 13 2
5 6 1 10 9 2
9 3 15 13 9 7 9 1 9 2
9 14 3 1 9 13 9 1 9 2
4 14 2 3 2
7 9 13 9 14 15 13 2
10 6 2 3 13 0 7 0 0 9 2
3 9 13 2
8 13 9 14 13 2 3 13 2
5 9 15 13 3 2
13 2 15 4 13 3 10 9 2 3 16 3 13 2
9 9 13 1 0 9 1 0 9 2
9 15 6 13 9 1 9 1 9 2
9 13 14 15 9 14 13 1 9 2
9 15 13 0 9 1 9 1 9 2
9 10 9 13 9 1 0 1 9 2
7 13 14 15 1 10 9 2
3 6 13 2
9 15 13 14 10 9 1 0 9 2
9 10 9 12 9 4 13 3 3 2
9 1 9 1 9 15 13 14 9 2
9 1 9 10 13 14 14 15 13 2
9 9 15 13 1 9 1 12 9 2
9 9 13 1 0 9 1 0 9 2
11 3 13 2 11 13 14 15 13 1 9 2
10 10 9 15 13 3 7 13 1 15 2
11 6 15 13 7 0 9 2 13 15 11 2
11 10 15 13 2 16 14 6 15 13 9 2
4 3 13 9 2
7 13 14 14 13 0 9 2
10 7 3 10 9 13 1 9 1 9 2
10 1 9 7 1 12 3 15 6 13 2
10 15 3 13 1 9 7 9 1 9 2
11 2 3 13 14 13 9 1 15 1 9 2
12 9 2 0 1 12 9 2 13 10 0 9 2
10 11 15 13 7 13 9 15 1 9 2
10 15 13 9 1 9 7 13 10 9 2
10 1 12 9 15 13 1 9 1 9 2
11 13 9 2 15 6 15 13 10 9 3 2
11 10 6 13 9 2 15 13 14 15 13 2
11 13 15 2 13 0 9 7 3 15 13 2
11 2 1 9 1 9 1 9 1 0 9 2
10 10 9 3 13 1 9 1 10 9 2
12 2 13 10 9 2 0 9 4 13 1 9 2
11 2 13 14 10 9 9 1 0 0 9 2
11 9 1 9 2 9 7 9 1 0 9 2
10 0 0 9 4 13 1 0 15 9 2
10 3 13 0 9 1 0 9 1 9 2
10 3 13 0 9 1 9 1 0 9 2
10 3 13 9 1 0 0 9 1 9 2
11 2 10 9 4 13 0 9 1 0 9 2
4 2 15 6 2
8 10 0 9 13 1 10 9 2
10 3 2 1 15 13 9 1 0 9 2
2 13 2
11 2 13 14 10 9 1 0 0 0 9 2
13 0 9 9 2 0 9 9 2 9 9 2 9 2
13 15 3 13 9 2 16 15 13 2 7 6 13 2
12 10 0 9 13 14 13 7 9 2 7 9 2
4 15 13 3 2
4 15 13 3 2
12 13 15 15 2 16 9 15 13 0 7 0 2
9 1 9 1 9 15 13 0 9 2
3 13 9 2
11 9 15 13 7 13 3 1 9 1 9 2
11 7 15 13 15 7 6 15 15 13 9 2
12 15 13 9 2 0 7 0 9 1 0 9 2
11 13 3 15 7 1 12 9 3 15 13 2
11 1 15 6 15 13 14 13 0 9 3 2
12 10 9 13 1 9 2 15 13 1 0 9 2
11 3 13 9 1 9 1 0 9 1 9 2
11 10 9 14 15 13 14 7 1 0 9 2
11 9 1 9 7 9 1 0 9 7 9 2
15 16 13 2 13 2 13 15 2 13 7 9 2 7 9 2
11 10 9 1 9 1 9 1 9 1 9 2
11 9 1 0 9 7 0 9 1 0 9 2
12 6 13 3 14 13 2 16 9 13 9 3 2
11 13 14 15 1 9 14 4 13 0 9 2
11 9 15 13 1 9 1 9 1 0 9 2
12 15 6 13 3 15 4 13 9 7 15 13 2
6 15 13 9 1 9 2
14 9 1 9 4 13 1 9 2 9 2 9 7 9 2
12 3 14 13 9 1 9 1 9 7 0 9 2
2 2 13
10 2 7 1 15 6 13 14 13 9 2
15 2 9 13 2 16 15 13 3 3 15 13 2 13 15 2
12 13 15 1 9 7 15 13 9 1 10 9 2
5 12 13 0 9 2
8 3 0 9 13 14 15 13 2
12 13 15 1 9 7 13 14 13 3 1 0 2
12 13 14 15 1 10 9 1 9 1 10 9 2
15 13 15 2 9 9 2 1 12 9 3 2 15 15 13 2
13 16 13 1 9 7 9 2 9 14 13 3 0 2
12 7 14 13 14 3 7 9 9 1 0 9 2
9 2 9 13 0 9 14 4 13 2
13 15 13 9 2 7 3 9 13 14 13 10 9 2
14 13 15 2 16 13 3 3 2 3 6 4 13 9 2
13 13 15 9 2 7 7 15 6 13 1 0 9 2
12 10 9 15 13 1 9 1 9 1 10 9 2
12 0 9 12 13 3 14 13 1 9 1 9 2
12 9 1 0 15 9 3 13 0 9 1 9 2
12 1 9 1 9 7 9 3 0 9 15 13 2
12 1 0 9 15 13 9 7 1 0 0 9 2
12 9 1 9 1 9 1 0 9 1 0 9 2
14 2 13 14 3 0 9 1 0 9 2 9 7 9 2
13 16 15 4 13 3 2 13 3 0 9 1 15 2
13 1 9 1 9 10 9 13 0 7 15 13 9 2
18 2 13 14 9 2 15 15 13 14 13 2 1 14 6 13 1 9 2
13 0 9 1 9 1 0 9 14 13 1 9 11 2
13 1 9 3 13 9 3 14 13 0 9 1 9 2
13 0 9 4 13 1 9 7 9 15 13 14 13 2
13 9 13 9 1 0 9 1 9 1 9 1 9 2
7 3 9 2 1 10 9 2
5 15 6 13 9 2
14 15 15 13 1 9 2 3 15 3 15 13 14 13 2
13 1 0 9 9 14 13 14 9 1 10 0 9 2
13 3 3 13 9 7 9 1 9 1 10 0 9 2
13 1 9 1 0 9 13 14 15 9 7 1 9 2
13 9 13 3 1 9 7 13 1 0 9 1 9 2
13 3 1 15 0 9 13 14 13 1 9 1 9 2
16 14 10 0 9 13 2 13 2 9 2 7 15 13 0 9 2
15 9 9 2 13 9 7 14 13 2 16 9 13 10 9 2
14 2 13 14 9 9 1 9 1 9 1 0 1 9 2
8 13 14 15 15 1 0 9 2
14 13 14 2 16 0 9 13 0 1 9 1 0 9 2
2 3 2
12 1 9 14 4 13 0 9 1 9 1 11 2
13 9 13 1 0 9 1 9 1 0 9 1 9 2
13 9 1 0 7 0 9 15 13 1 0 0 9 2
14 1 0 9 14 15 13 9 1 9 2 13 3 9 2
13 13 15 1 10 3 10 9 1 0 9 1 9 2
13 1 9 1 0 9 14 13 1 9 1 0 9 2
13 7 9 13 1 0 9 2 3 13 1 0 9 2
14 11 9 13 0 9 1 0 9 2 16 15 13 9 2
13 9 1 0 9 13 9 7 9 1 0 0 9 2
15 15 13 2 16 10 9 13 0 9 2 15 13 0 9 2
16 13 15 15 2 16 6 15 13 2 3 3 3 13 9 15 2
8 13 15 7 1 3 15 13 2
9 3 13 14 15 13 7 3 13 2
7 15 13 14 2 3 13 2
5 6 13 1 9 2
15 1 3 0 9 1 0 9 13 2 16 15 15 13 0 2
14 9 1 9 1 9 13 14 15 13 3 1 12 9 2
14 13 0 15 9 2 1 14 13 10 3 0 15 9 2
4 13 15 3 2
15 3 15 13 2 16 13 10 9 7 15 6 15 13 0 2
14 3 15 13 9 7 9 1 9 1 9 1 0 9 2
12 13 9 1 9 2 3 3 9 15 13 9 2
4 13 15 15 2
6 9 13 1 0 9 2
9 15 14 13 3 0 9 1 9 2
14 0 0 9 1 0 0 9 13 0 9 1 0 9 2
15 2 1 3 9 4 13 9 1 9 1 0 15 0 9 2
14 9 1 9 1 9 1 0 9 15 13 1 0 9 2
2 13 2
14 1 10 9 14 13 7 1 0 9 1 0 0 9 2
7 1 9 15 13 0 9 2
8 15 4 13 9 1 0 9 2
15 2 1 9 1 0 9 3 0 9 13 7 10 0 9 2
14 15 14 15 13 1 10 3 0 9 14 13 9 15 2
17 9 0 4 13 9 1 9 2 9 2 9 2 9 7 0 9 2
15 2 10 9 4 13 9 1 9 1 0 9 1 0 9 2
17 2 13 14 4 9 2 3 10 3 0 1 9 9 13 1 9 2
18 9 13 14 15 13 7 13 2 1 14 15 13 9 1 9 1 9 2
9 3 0 14 13 3 9 1 9 2
7 13 14 15 1 0 9 2
2 3 2
15 9 1 9 13 14 4 13 1 9 1 0 9 1 9 2
15 1 10 9 15 13 1 0 9 7 9 1 0 0 9 2
2 15 2
15 14 13 14 3 0 9 7 9 1 10 9 7 0 9 2
17 2 13 14 2 16 14 15 13 7 9 1 10 9 1 0 9 2
16 2 9 9 2 10 13 1 9 1 9 9 14 13 12 9 2
16 9 1 9 1 9 2 9 1 9 1 0 9 1 0 9 2
16 9 13 2 16 9 1 9 13 1 0 9 1 9 1 9 2
10 9 1 0 0 9 6 13 0 9 2
6 15 0 15 13 15 2
18 3 13 2 9 7 9 2 16 13 9 2 0 6 13 0 15 9 2
16 3 13 1 9 1 9 1 9 1 9 2 0 1 0 9 2
15 1 10 0 9 15 14 13 0 1 9 15 1 0 9 2
8 14 15 13 1 10 13 9 2
16 10 9 1 0 9 13 14 13 1 0 9 2 0 14 13 2
9 3 15 13 3 1 9 1 9 2
12 3 13 2 13 0 9 1 9 1 0 9 2
6 1 3 15 13 9 2
18 12 9 7 9 2 0 1 9 1 9 1 0 9 2 13 3 9 2
18 2 13 9 1 9 15 2 7 3 3 13 14 15 13 1 0 9 2
12 2 15 13 7 1 10 3 0 0 0 9 2
4 15 13 9 2
14 13 9 14 13 3 3 2 9 4 13 9 1 9 2
14 14 15 3 14 13 7 9 1 10 9 15 13 11 2
10 3 0 3 6 13 3 3 14 13 2
18 1 11 13 3 2 16 13 9 1 9 1 0 0 9 1 9 15 2
30 11 15 13 3 2 13 1 9 1 9 1 9 2 1 15 4 13 3 2 13 10 9 7 1 9 15 13 0 9 2
6 1 9 15 13 9 2
8 9 15 13 1 1 0 9 2
6 13 1 9 1 9 2
14 2 1 10 9 3 14 4 13 0 9 1 0 9 2
22 13 15 14 2 16 1 10 3 0 9 10 9 14 13 9 1 0 0 9 1 9 2
16 4 13 1 9 3 3 14 13 9 1 9 15 1 10 9 2
11 7 3 13 2 16 10 9 6 13 0 2
11 0 9 9 2 0 9 7 9 0 9 2
25 13 4 7 9 1 9 2 9 2 9 7 9 2 15 15 13 1 9 1 9 1 0 0 11 2
25 13 4 9 1 10 9 1 0 0 9 1 0 9 1 9 1 9 1 9 7 1 0 0 9 2
38 7 0 0 9 15 13 1 9 2 15 13 14 13 0 0 9 1 0 9 1 0 9 1 0 9 11 7 9 1 9 1 0 9 1 9 1 11 2
30 15 13 3 1 9 1 0 11 2 3 1 15 15 13 1 10 0 9 7 13 9 2 15 15 13 14 13 1 15 2
17 1 9 1 0 0 9 1 15 15 13 9 2 9 7 0 9 2
26 1 9 1 0 0 9 15 4 13 1 9 1 11 2 7 0 9 1 9 1 9 13 3 0 9 2
16 11 3 13 1 9 1 9 11 14 4 13 1 0 0 9 2
17 13 4 9 9 1 9 1 0 11 14 13 9 1 0 0 11 2
40 0 13 9 2 16 1 9 1 0 9 1 11 1 0 9 1 11 9 1 0 9 14 13 0 9 1 0 9 1 0 0 9 2 15 13 1 9 1 9 2
6 13 9 1 0 9 2
14 1 9 0 13 9 7 9 2 7 3 15 9 13 2
6 0 9 13 0 9 2
10 7 2 11 13 10 9 1 10 9 2
22 6 2 10 9 1 9 3 4 13 2 7 14 9 2 0 1 0 9 2 13 9 2
8 13 1 9 2 7 15 13 2
14 3 15 13 0 9 14 13 9 2 3 13 0 9 2
9 13 9 2 1 15 4 13 9 2
9 1 9 3 14 13 1 12 11 2
8 13 14 3 7 9 1 9 2
6 3 15 6 15 13 2
24 3 4 13 9 2 16 9 1 10 9 15 13 1 9 1 0 9 1 9 7 0 0 9 2
22 9 1 9 3 15 13 2 9 15 13 3 3 7 9 15 13 1 9 7 0 9 2
15 2 9 3 4 13 13 10 9 1 9 1 9 1 9 2
15 3 15 13 15 9 7 1 10 3 1 9 13 0 9 2
32 12 9 13 9 1 9 1 9 1 0 11 7 13 9 2 16 13 0 0 9 1 9 15 1 0 9 1 0 9 1 9 2
21 9 1 0 9 1 9 1 9 1 10 1 9 1 9 1 0 9 14 4 13 2
30 1 10 9 9 13 1 9 14 13 9 1 0 9 1 9 0 1 9 7 9 1 9 2 1 0 9 1 0 9 2
24 14 3 9 13 14 13 9 14 1 9 15 2 7 15 13 2 16 13 3 14 15 13 9 2
26 2 1 9 1 9 1 9 1 9 2 9 13 9 1 0 9 1 9 2 16 15 13 1 10 9 2
9 7 13 2 16 6 15 13 0 2
23 1 10 9 9 13 14 15 13 1 9 1 0 7 0 0 9 7 9 2 13 11 11 2
27 7 9 15 13 9 7 9 15 13 9 7 7 9 1 9 2 7 9 1 9 1 9 13 14 15 13 2
23 1 9 10 9 9 15 13 1 0 9 1 11 2 1 14 13 0 9 1 9 1 9 2
38 1 9 1 9 11 1 11 4 13 9 1 0 9 7 9 1 9 1 9 1 12 0 9 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
14 13 15 1 0 9 14 15 13 11 2 11 7 11 2
13 11 3 13 9 1 9 1 9 1 9 1 11 2
10 13 11 1 9 7 6 15 13 3 2
10 15 15 13 2 16 14 13 1 15 2
6 13 15 4 1 11 2
6 1 0 11 13 0 2
9 3 13 14 13 3 13 10 9 2
13 7 16 1 9 1 9 1 15 3 13 10 9 2
4 13 15 9 2
9 9 1 11 15 13 1 10 9 2
24 14 13 2 16 10 9 13 0 0 9 7 13 9 1 9 1 0 9 1 9 1 12 9 2
25 3 12 1 0 9 1 9 1 0 9 13 9 1 9 1 9 9 1 9 7 9 1 0 9 2
30 1 0 9 1 10 9 3 13 14 15 13 9 1 0 9 7 3 13 9 1 9 1 9 1 9 1 9 1 9 2
24 11 4 13 0 9 2 0 15 1 9 1 9 2 9 1 9 2 9 1 9 7 1 9 2
16 15 13 3 0 15 9 1 9 15 2 3 3 15 4 13 2
21 15 13 0 15 1 9 9 2 3 2 1 10 9 13 7 1 9 1 9 15 2
22 13 1 9 1 14 13 1 11 2 0 9 14 13 1 9 2 0 1 0 0 9 2
16 3 16 10 9 15 4 13 7 3 3 13 2 1 1 9 2
6 13 1 9 1 9 2
12 3 13 1 11 2 4 13 3 9 1 9 2
14 1 10 9 1 11 13 1 9 0 9 1 0 9 2
15 6 15 14 13 9 1 9 14 13 1 9 1 0 9 2
22 10 9 15 13 1 0 9 1 9 1 9 1 9 1 0 9 1 9 1 0 9 2
28 3 9 13 9 1 0 1 9 11 9 1 9 1 9 1 9 1 0 9 2 15 14 4 13 1 0 9 2
14 0 9 7 0 9 1 10 9 13 9 1 9 15 2
7 15 15 13 1 11 3 2
19 7 9 15 13 9 1 9 1 10 9 2 3 4 13 3 9 1 9 2
10 11 3 13 9 7 13 1 0 9 2
6 7 3 9 3 13 2
14 9 15 13 3 1 9 2 15 3 13 1 9 15 2
11 9 15 4 13 1 0 9 1 10 9 2
28 9 1 0 9 11 11 15 13 3 1 11 11 2 9 1 9 1 0 0 2 0 7 0 9 1 0 9 2
5 7 11 13 0 2
18 0 9 3 15 15 13 2 13 15 1 10 9 2 7 13 1 9 2
12 0 0 9 13 0 9 1 11 1 0 9 2
16 13 9 1 0 9 1 11 7 1 0 9 1 0 9 11 2
16 1 0 9 13 2 16 11 13 9 1 0 9 1 0 9 2
5 3 13 10 9 2
16 11 15 6 13 2 13 9 1 9 7 13 14 13 9 15 2
17 2 14 13 14 0 9 1 0 9 1 9 1 9 7 0 9 2
16 15 3 15 13 1 9 3 3 0 7 1 0 9 1 15 2
17 3 3 15 13 1 9 7 9 1 0 9 2 15 13 1 9 2
7 14 6 13 3 1 9 2
10 0 9 1 9 13 7 10 0 9 2
5 13 15 0 9 2
6 14 13 7 0 9 2
6 13 14 15 13 9 2
21 14 2 15 13 2 9 7 9 2 0 9 1 9 2 15 13 15 7 0 9 2
18 15 13 14 13 3 0 2 16 15 13 9 14 13 9 15 1 9 2
18 15 14 13 9 1 9 1 9 7 0 9 7 1 9 1 0 9 2
23 9 2 1 15 3 15 13 0 0 9 2 6 13 14 15 13 1 0 9 1 1 0 2
15 10 9 1 9 15 13 1 9 2 1 14 13 9 15 2
6 0 15 13 1 9 2
21 0 0 9 2 15 13 3 0 1 9 1 9 2 13 0 9 1 9 1 9 2
15 9 2 15 13 7 1 9 1 10 0 7 0 0 9 2
22 3 14 13 2 16 1 15 15 13 7 1 10 9 2 15 13 9 1 0 0 9 2
10 13 15 2 16 15 6 13 0 9 2
8 0 13 9 7 1 0 9 2
5 13 7 0 9 2
22 7 3 3 6 13 14 15 13 3 9 2 3 15 15 13 9 2 15 4 13 9 2
25 0 9 1 9 14 15 13 1 0 9 2 1 14 13 14 13 9 1 0 9 2 13 3 9 2
7 1 15 13 10 0 9 2
19 2 1 9 1 9 13 9 1 0 9 1 9 1 9 1 9 1 9 2
2 13 2
14 3 1 9 13 9 15 2 7 13 3 14 15 13 2
24 13 15 0 2 13 15 1 3 2 13 1 10 9 2 7 13 9 7 15 13 3 1 15 2
23 9 2 9 1 9 2 10 9 7 9 1 9 1 9 15 13 1 9 1 9 1 9 2
7 7 15 13 14 13 9 2
14 1 9 1 9 15 13 2 16 10 9 13 1 9 2
23 13 4 9 1 9 1 0 9 7 0 9 1 9 1 0 9 2 9 7 9 1 9 2
13 13 14 2 16 1 9 13 9 1 9 15 3 2
10 1 3 12 9 13 7 9 1 9 2
14 10 1 9 15 13 2 15 13 1 9 14 15 13 2
24 1 9 1 9 12 9 3 15 13 1 9 1 9 1 9 2 3 7 1 9 1 0 9 2
23 13 14 3 0 15 9 1 9 1 9 1 9 7 0 9 7 3 3 13 3 1 15 2
14 9 2 13 3 10 9 2 16 15 13 9 14 13 2
23 1 10 9 4 13 9 1 9 1 9 1 0 9 7 0 9 1 9 1 9 7 9 2
23 9 13 0 9 9 14 13 0 0 9 1 0 9 7 1 0 9 1 9 1 0 9 2
9 13 15 3 1 9 1 0 9 2
25 1 10 9 12 13 1 0 9 1 9 2 13 15 1 12 9 7 15 13 1 12 1 0 9 2
14 13 15 1 10 9 2 13 2 9 15 15 13 3 2
8 0 9 13 0 1 0 9 2
18 3 13 0 9 2 15 14 13 9 1 9 1 9 7 9 1 9 2
14 9 7 9 1 9 1 9 13 9 1 0 0 9 2
19 3 1 9 2 15 13 9 9 2 13 13 1 0 9 1 0 15 9 2
25 1 9 1 0 9 1 9 1 9 1 9 1 9 15 13 0 9 1 9 7 9 1 0 9 2
4 9 13 0 2
23 9 1 9 13 14 13 9 1 9 15 2 7 15 1 10 9 14 13 9 15 1 9 2
26 9 1 10 9 13 0 1 0 9 1 9 1 9 2 7 1 0 9 10 9 13 9 1 10 9 2
18 13 2 16 3 13 10 9 2 15 4 13 14 13 0 9 1 9 2
18 13 2 16 3 13 10 9 2 15 4 13 14 13 0 9 1 9 2
16 9 13 1 9 1 9 1 0 9 7 0 9 1 0 9 2
18 14 15 13 2 0 9 2 1 0 9 14 15 13 1 9 1 9 2
17 1 0 9 2 9 13 1 0 9 1 9 7 9 1 0 9 2
18 0 3 13 14 2 16 9 1 9 7 9 1 9 7 9 4 13 2
4 11 15 13 2
16 6 13 15 2 13 15 9 2 16 3 3 13 10 10 9 2
18 2 3 9 1 9 1 0 9 14 15 13 1 9 15 1 0 9 2
15 2 12 1 9 2 15 13 2 13 0 9 1 0 9 2
6 3 14 15 13 15 2
18 1 10 9 2 15 13 9 1 0 9 1 9 1 9 1 0 9 2
17 3 7 3 14 4 13 9 1 9 1 9 7 9 1 0 9 2
18 15 4 13 1 3 0 0 9 2 1 9 1 9 1 9 1 9 2
18 13 15 1 10 9 1 10 0 1 15 9 2 15 13 3 1 9 2
18 1 15 3 13 0 9 2 9 1 0 9 7 9 1 9 1 9 2
8 0 0 9 13 9 7 9 2
20 9 11 2 3 15 13 9 7 3 9 15 15 13 9 2 13 14 15 13 2
5 15 6 13 15 2
19 3 2 9 1 9 1 0 9 1 9 1 9 7 1 9 1 10 9 2
18 1 9 1 9 15 9 1 9 15 13 1 9 1 0 9 7 9 2
6 3 13 10 10 9 2
23 2 6 15 13 9 2 7 15 13 9 1 9 2 3 16 6 1 10 9 13 0 9 2
18 9 7 9 1 10 0 9 13 0 9 1 0 9 7 1 0 9 2
20 0 0 9 1 0 2 0 7 0 9 13 9 7 9 1 0 9 1 9 2
18 9 1 0 9 7 0 9 13 9 1 9 1 9 1 12 0 9 2
7 13 4 0 9 1 9 2
12 9 6 4 13 1 0 9 7 13 1 9 2
20 9 1 0 0 9 2 0 1 0 0 9 2 13 14 4 13 1 0 9 2
19 1 10 9 4 13 0 9 7 13 14 4 0 9 1 0 9 1 9 2
19 0 9 13 9 1 0 0 9 7 1 9 1 0 9 1 9 15 3 2
7 9 6 13 7 14 13 2
13 13 15 3 1 15 7 9 13 9 3 1 9 2
21 2 9 1 0 9 13 7 0 9 1 0 9 2 15 4 13 1 9 0 9 2
19 13 14 4 13 9 7 9 1 0 9 1 0 9 1 9 1 0 9 2
22 9 13 0 9 2 0 1 0 9 2 0 1 9 1 9 7 0 1 10 9 9 2
15 1 9 4 13 9 1 0 9 1 0 9 1 0 9 2
9 0 9 13 0 9 1 0 9 2
14 13 3 9 1 9 13 3 1 0 9 1 0 3 2
19 13 2 13 2 13 2 13 1 0 9 7 16 15 6 13 2 6 13 2
7 3 13 14 15 13 9 2
8 1 15 13 1 9 9 15 2
19 7 13 14 7 15 13 1 0 9 2 13 3 0 9 7 13 9 3 2
14 9 15 13 14 13 10 15 13 2 3 9 13 11 2
29 9 1 9 1 9 11 1 9 1 10 0 9 2 3 1 0 9 2 1 15 1 3 9 13 15 14 4 13 2
40 16 0 0 7 0 0 9 15 13 10 0 0 9 1 11 1 0 2 0 7 0 9 1 0 0 9 2 14 15 6 13 9 1 9 7 9 1 0 9 2
26 0 9 2 0 1 0 9 7 9 1 9 2 15 15 13 1 0 9 2 6 15 13 1 0 11 2
18 0 9 1 0 9 0 1 9 9 2 9 7 9 13 9 1 9 2
17 0 9 9 2 0 9 7 9 0 9 2 0 9 7 9 9 2
24 13 2 16 15 4 3 13 14 13 7 10 9 1 0 9 1 9 1 11 1 9 1 9 2
24 13 2 16 15 4 3 13 14 13 7 10 9 1 0 9 1 9 1 11 1 9 1 9 2
38 3 1 15 15 13 3 2 13 3 2 3 15 13 3 1 9 2 6 3 14 13 9 2 7 14 13 0 9 2 9 2 0 1 3 0 0 9 2
13 2 0 13 2 16 0 9 4 13 1 0 9 2
26 1 9 2 16 15 13 3 9 1 9 1 9 7 10 9 2 13 9 15 1 0 9 1 0 9 2
14 15 15 13 9 2 13 9 7 13 2 3 15 13 2
5 11 13 1 15 2
14 12 15 13 9 14 13 7 11 3 13 9 1 9 2
26 3 0 0 9 2 0 1 0 9 1 9 2 13 1 0 9 1 0 0 0 9 3 1 12 9 2
14 9 13 3 3 7 11 13 0 15 9 14 1 9 2
24 14 10 0 9 13 9 1 0 9 2 7 9 15 13 3 0 2 16 15 13 14 15 13 2
23 9 3 13 11 14 15 13 9 1 0 9 2 7 9 3 15 13 14 15 13 1 9 2
10 9 1 9 13 1 9 1 12 9 2
18 1 9 1 10 9 12 0 9 14 13 9 1 11 1 9 1 9 2
19 13 9 14 15 13 0 9 1 9 2 3 7 0 7 0 14 13 15 2
10 0 9 13 14 15 13 9 2 9 2
41 9 7 9 1 0 9 1 9 13 14 15 13 3 7 10 0 9 2 7 0 9 2 3 0 9 6 13 9 2 7 12 1 9 1 9 1 0 9 1 9 2
9 15 13 0 9 1 0 0 9 2
18 15 13 9 1 0 14 13 1 9 1 0 9 7 0 9 1 9 2
5 7 15 15 13 2
26 16 15 13 9 1 0 0 9 2 6 15 13 14 6 14 13 1 0 0 1 9 15 1 9 9 2
4 14 13 3 2
6 3 15 3 4 13 2
11 9 2 2 13 9 15 0 9 1 9 2
24 10 9 1 9 11 2 13 15 3 7 15 13 2 2 10 9 1 9 4 13 14 15 13 2
14 14 13 3 14 15 13 2 7 14 13 10 0 9 2
8 6 10 0 9 13 10 9 2
10 14 13 1 9 15 1 9 1 11 2
55 9 1 10 9 2 15 13 2 13 16 3 3 2 3 3 13 0 0 0 9 1 9 1 10 9 7 9 1 9 1 0 9 1 0 0 0 9 2 3 3 9 9 1 9 1 0 9 13 14 13 1 9 1 11 2
17 16 15 13 1 0 9 2 3 13 16 10 9 14 13 14 13 2
3 0 9 2
34 15 13 2 0 13 2 11 9 2 14 13 2 13 14 13 0 9 1 9 2 7 1 10 11 13 15 14 15 13 7 9 15 13 2
21 7 13 14 9 2 14 15 6 13 2 7 13 15 9 7 13 1 0 9 14 2
12 0 9 1 0 9 13 1 9 1 0 9 2
8 15 13 0 9 1 0 9 2
20 16 15 6 15 13 1 10 9 1 0 9 2 15 6 13 14 13 0 9 2
9 0 9 13 0 9 1 0 9 2
19 3 15 1 9 1 0 9 2 15 6 4 13 14 13 0 1 15 9 2
28 13 14 13 0 0 9 1 9 7 1 9 1 0 9 7 9 14 15 13 9 7 9 2 1 15 15 13 2
19 10 3 13 2 3 1 9 2 16 13 0 1 10 9 1 9 1 11 2
22 1 9 1 9 1 0 0 9 9 1 0 9 13 2 16 9 1 0 9 4 13 2
16 13 14 2 16 9 1 11 13 2 3 13 14 13 0 9 2
21 7 16 14 15 13 9 15 2 13 15 1 9 15 7 15 13 1 9 1 9 2
8 13 9 7 13 3 1 9 2
18 13 9 2 3 15 13 2 7 6 15 13 2 9 14 13 1 15 2
37 1 0 9 1 0 9 2 3 12 1 9 13 0 9 2 0 10 9 13 3 0 9 1 9 1 9 2 1 14 6 15 13 9 1 0 9 2
19 13 15 2 13 15 2 0 13 7 13 2 7 0 15 13 7 13 9 2
10 14 15 13 9 1 10 2 15 13 2
24 15 1 0 4 13 1 10 10 9 14 13 14 15 13 3 13 10 0 9 2 0 15 9 2
21 7 16 15 13 2 16 14 13 0 9 1 10 9 2 15 13 14 13 0 9 2
3 2 3 2
9 15 6 3 13 14 13 0 9 2
22 7 16 15 13 14 13 10 9 1 9 1 0 9 2 13 3 14 15 15 13 9 2
12 10 9 4 13 3 1 9 9 1 0 9 2
12 9 1 9 2 9 7 9 13 6 12 9 2
10 13 13 15 14 13 0 9 1 9 2
4 2 3 13 2
20 9 13 9 1 0 9 1 9 15 2 3 7 1 9 1 0 0 0 9 2
18 11 6 4 13 15 7 3 15 13 1 9 1 10 9 1 0 9 2
17 16 4 15 13 10 9 2 3 13 14 13 3 1 0 9 9 2
6 13 15 3 1 15 2
12 11 4 13 1 9 1 9 1 0 15 9 2
14 9 1 9 1 9 1 0 0 11 15 13 3 3 2
19 9 1 0 7 0 9 13 1 0 9 1 0 9 7 0 9 1 9 2
35 1 9 4 13 9 1 9 1 9 1 9 7 10 9 1 9 1 9 7 4 13 9 1 11 7 11 14 15 13 1 9 1 0 9 2
4 11 13 9 2
22 3 7 6 13 3 15 4 13 1 11 2 7 16 13 9 15 2 15 13 1 9 2
9 11 13 1 9 1 0 0 9 2
15 7 2 1 9 1 0 2 1 0 9 1 9 1 9 2
18 3 9 1 0 9 1 9 1 9 4 13 2 16 9 3 13 9 2
40 9 13 3 1 9 2 13 11 9 15 2 9 15 13 9 7 16 13 1 9 2 13 7 9 2 7 9 2 13 1 13 7 1 0 3 9 13 12 9 2
13 9 15 13 2 9 13 2 9 3 13 10 9 2
12 11 13 9 15 1 0 9 2 13 7 9 2
13 10 9 3 15 13 2 9 15 13 1 0 9 2
12 11 15 13 1 15 2 3 13 9 2 13 2
8 0 9 13 0 9 1 11 2
13 15 13 9 1 11 2 3 3 15 13 14 13 2
13 15 13 9 1 11 2 3 3 15 13 14 13 2
40 9 3 4 13 10 0 9 2 16 3 15 13 1 10 1 3 0 0 9 2 1 15 15 6 4 13 9 14 14 15 13 2 1 14 13 1 0 0 9 2
6 11 15 13 1 9 2
20 9 1 0 0 9 1 9 11 15 13 1 0 9 7 0 0 9 1 9 2
17 0 9 1 0 9 1 9 1 9 7 9 13 9 1 0 9 2
14 1 15 4 13 10 0 9 2 0 2 0 2 0 2
17 1 1 11 15 13 1 15 2 11 3 15 13 1 10 15 9 2
9 13 15 10 0 9 1 0 9 2
6 9 13 9 1 9 2
5 13 15 0 9 2
7 13 2 16 13 1 9 2
17 13 3 9 7 9 1 9 2 16 9 15 13 2 7 0 13 2
16 1 0 9 9 1 9 1 9 7 9 1 11 13 3 0 2
11 15 15 13 0 9 1 0 9 7 9 2
11 3 1 9 10 9 15 4 13 0 9 2
7 9 1 11 6 13 0 2
8 14 1 9 13 9 1 11 2
24 1 9 11 4 13 9 1 0 0 9 7 1 9 1 0 9 2 15 4 13 3 0 9 2
20 15 15 13 9 14 13 2 13 15 12 9 2 0 1 9 15 1 0 9 2
17 13 12 9 2 3 15 4 13 1 0 9 7 3 6 13 0 2
3 0 9 2
5 13 15 1 15 2
2 13 2
17 7 14 1 9 2 15 14 13 9 1 0 9 7 14 13 9 2
22 15 13 3 0 2 3 0 9 13 1 0 9 7 3 15 13 1 9 1 0 9 2
8 1 3 3 9 13 3 0 2
13 13 15 1 9 7 1 10 9 1 10 0 9 2
23 14 3 3 15 4 13 10 0 9 1 0 9 2 15 14 13 14 15 13 1 0 9 2
24 3 13 14 13 3 0 1 9 15 1 9 1 0 9 2 3 16 13 1 9 1 0 9 2
29 13 2 16 13 14 13 0 2 3 0 2 3 0 9 2 7 9 13 7 14 13 14 13 0 9 1 10 9 2
14 9 6 13 1 10 9 1 9 2 15 3 13 3 2
15 13 15 2 16 13 3 14 15 13 9 2 15 13 0 2
15 7 3 1 15 1 9 2 15 13 2 15 13 1 15 2
17 15 13 3 3 14 13 1 9 2 7 13 0 9 14 13 9 2
4 13 1 15 2
8 13 15 2 16 15 13 9 2
4 13 0 11 2
7 15 13 0 9 1 11 2
12 2 1 9 1 9 1 9 3 13 0 9 2
3 13 9 2
6 1 9 13 14 13 2
23 12 1 9 2 1 15 0 9 1 9 3 13 14 13 1 9 1 9 2 3 13 9 2
14 1 9 1 9 9 15 15 13 7 15 13 1 9 2
10 13 0 9 2 0 9 2 0 9 2
14 7 3 9 15 13 14 13 3 1 0 9 1 9 2
17 0 2 6 13 2 16 3 13 10 9 1 0 9 7 0 9 2
14 9 1 9 13 7 9 9 1 9 1 9 1 9 2
11 15 13 14 13 7 9 1 9 1 9 2
11 3 3 6 13 14 4 13 7 10 9 2
29 2 9 1 9 13 1 10 9 2 9 13 14 13 9 2 15 14 13 9 7 14 15 13 2 3 10 15 13 2
12 14 3 13 9 1 9 2 15 13 3 9 2
20 1 9 1 9 1 11 3 2 1 15 4 13 2 16 4 13 9 1 9 2
17 15 15 13 9 14 15 13 9 2 3 3 13 9 1 0 9 2
15 1 3 1 9 13 9 1 0 9 2 15 13 1 9 2
17 1 9 13 0 9 7 15 13 14 13 1 12 1 9 1 9 2
7 12 9 15 13 10 9 2
12 7 13 14 2 3 3 13 14 13 1 15 2
22 9 15 13 2 16 14 15 13 1 15 1 0 9 2 3 6 13 14 13 0 9 2
35 11 11 13 1 0 9 2 16 15 13 2 3 13 3 2 13 0 15 9 7 13 2 16 9 15 3 6 15 13 1 9 1 0 9 2
18 3 15 13 9 7 13 3 2 16 15 13 3 1 9 2 16 13 2
23 11 11 6 13 14 15 13 1 9 14 6 13 9 14 15 13 7 14 15 13 1 9 2
19 3 15 15 13 1 10 9 2 13 11 11 7 13 14 15 13 1 9 2
11 13 14 13 3 0 1 9 1 0 9 2
2 6 2
5 15 14 15 13 2
19 7 2 3 0 2 0 9 13 14 13 9 0 9 2 0 1 0 9 2
13 1 9 1 0 9 0 0 9 13 0 1 9 2
9 1 9 13 9 1 9 7 9 2
5 2 13 1 11 2
6 1 9 3 13 3 2
15 0 9 13 0 1 9 1 0 9 7 15 3 15 13 2
5 9 15 3 13 2
8 4 13 11 2 15 13 9 2
8 7 13 13 13 15 14 2 2
9 1 9 1 9 13 15 0 9 2
7 3 6 13 14 15 13 2
10 1 9 9 13 0 9 1 0 9 2
18 9 2 1 15 15 13 2 1 14 15 13 1 10 9 2 13 0 2
12 9 1 9 13 9 1 0 7 9 1 0 2
24 11 13 1 9 2 14 15 6 13 2 16 11 3 3 15 13 2 16 15 4 13 1 15 2
6 2 13 1 12 9 2
5 13 14 15 13 2
8 15 13 1 15 1 0 9 2
7 9 3 4 13 1 11 2
8 7 0 1 0 9 3 13 2
10 0 9 1 0 9 13 0 1 9 2
15 1 9 1 11 1 0 9 11 15 13 1 3 0 9 2
6 3 15 13 0 9 2
10 3 15 13 3 1 9 1 9 11 2
4 13 0 9 2
11 11 15 13 3 1 9 3 1 0 9 2
3 13 11 2
20 0 9 1 11 2 7 7 1 11 13 3 13 9 1 0 0 9 1 9 2
19 7 0 0 9 14 4 14 13 1 11 2 3 4 13 1 9 1 9 2
25 1 9 9 1 0 9 15 13 9 1 9 1 9 2 9 1 9 1 9 2 0 9 7 9 2
17 7 16 15 13 9 2 13 15 9 1 9 7 15 13 1 9 2
17 1 9 7 12 13 2 3 13 1 10 3 9 14 13 1 9 2
19 7 15 13 2 1 14 13 9 14 13 0 2 7 13 3 14 4 13 2
5 0 9 13 14 2
18 13 15 3 3 2 16 10 0 9 1 15 15 13 7 3 15 13 2
19 13 3 14 15 13 2 16 7 9 6 4 13 2 7 14 3 15 13 2
23 9 9 13 15 2 7 13 9 2 16 16 14 15 13 14 6 15 13 3 7 9 15 2
7 13 15 9 7 15 13 2
12 13 9 11 2 13 3 7 13 1 0 9 2
8 15 13 0 7 15 13 0 2
6 13 2 16 13 3 2
24 7 9 13 1 9 2 7 3 13 10 9 2 1 0 9 13 9 2 7 6 13 3 9 2
6 14 14 3 13 9 2
17 16 3 15 13 15 1 3 0 9 1 9 2 15 3 13 3 2
24 16 15 13 2 13 15 1 3 9 2 7 13 2 13 15 1 9 7 9 15 13 1 9 2
23 13 15 2 13 1 9 7 3 16 13 9 2 10 0 9 1 0 9 15 13 1 9 2
9 10 9 4 13 1 9 1 15 2
23 1 9 1 9 1 11 7 0 9 1 11 2 0 13 14 15 13 7 1 0 0 9 2
24 2 10 14 15 13 1 9 1 9 1 10 10 9 2 15 15 13 1 0 1 0 0 9 2
11 9 15 13 2 1 15 14 4 15 13 2
16 7 7 0 9 15 13 2 3 16 15 3 13 1 0 9 2
26 14 14 4 15 13 2 3 13 9 2 14 15 13 9 1 9 7 13 14 13 2 16 6 13 9 2
25 13 2 16 3 1 10 9 6 13 14 4 13 7 0 9 2 6 13 14 4 13 7 0 9 2
14 11 15 13 1 12 1 9 7 15 13 14 13 11 2
8 3 15 13 1 9 1 9 2
25 9 6 13 1 9 1 9 2 7 3 15 13 0 7 15 15 13 2 3 15 3 1 9 15 2
11 7 15 15 13 0 9 1 10 0 9 2
24 1 9 4 13 9 1 9 7 9 1 9 1 12 9 1 9 1 9 2 0 1 0 9 2
25 9 15 13 2 16 7 4 13 10 0 9 1 9 2 7 14 15 15 4 13 1 9 1 9 2
13 2 12 9 15 13 2 1 1 15 4 13 9 2
26 9 1 9 1 11 13 9 2 15 13 1 9 1 0 9 7 0 9 2 15 13 3 1 0 9 2
7 1 9 13 0 0 9 2
21 2 14 13 9 1 0 9 2 16 15 13 14 13 0 9 2 1 1 13 9 2
16 2 0 9 14 13 9 1 0 9 2 15 13 0 1 9 2
12 0 13 2 16 14 15 13 7 3 0 9 2
13 13 15 9 9 14 13 14 13 3 2 7 6 2
10 9 15 6 13 15 2 7 3 13 2
19 15 3 6 4 13 2 7 9 1 0 0 9 1 0 9 2 15 13 2
15 7 16 15 13 14 13 3 2 15 13 1 0 9 3 2
20 13 15 3 7 9 2 16 1 9 9 13 14 13 9 1 10 9 7 9 2
18 14 16 15 13 9 1 10 0 9 1 9 2 9 1 15 4 13 2
10 2 3 3 3 0 13 9 1 9 2
9 3 15 13 1 9 1 9 3 2
12 15 13 0 9 1 9 1 0 1 9 9 2
6 13 14 4 1 0 2
9 6 15 13 3 2 7 13 9 2
11 10 9 9 2 9 1 9 7 0 9 2
18 9 1 9 13 0 9 1 0 9 7 1 0 9 1 9 1 9 2
7 13 14 9 1 0 9 2
12 9 13 14 3 9 1 0 9 7 0 9 2
9 3 13 1 0 9 1 0 9 2
10 9 9 2 0 9 2 9 2 9 2
12 3 15 13 1 10 9 14 13 1 0 9 2
19 9 1 10 9 1 9 1 9 14 13 9 1 9 1 0 9 1 9 2
19 0 9 3 13 9 1 9 15 1 9 1 0 7 0 9 1 0 9 2
9 16 6 13 9 3 2 9 9 2
2 15 2
4 14 15 13 2
7 14 13 1 9 1 9 2
13 16 13 2 13 15 2 16 13 2 13 15 3 2
6 1 10 9 13 9 2
10 3 1 9 2 3 2 9 6 13 2
21 1 10 9 6 4 13 9 1 9 1 9 1 0 9 2 0 9 2 0 9 2
16 0 9 2 10 13 1 9 7 9 2 1 15 15 13 9 2
17 1 0 15 9 2 1 1 9 2 15 15 13 3 7 1 9 2
17 0 9 1 0 9 1 11 2 11 11 13 3 7 9 0 9 2
12 7 2 0 9 1 9 1 9 13 0 9 2
9 9 1 9 13 9 1 0 9 2
13 9 1 10 9 13 6 4 13 1 0 15 9 2
26 16 13 2 16 9 1 0 9 12 9 3 1 9 4 13 1 9 2 15 13 1 9 1 0 9 2
25 3 13 2 16 1 14 15 13 9 3 2 15 13 3 9 1 9 2 0 1 0 9 1 9 2
12 7 15 13 2 16 0 9 15 13 15 3 2
18 16 1 10 9 15 4 13 1 9 1 10 9 2 15 13 10 9 2
24 16 15 13 1 10 9 2 9 13 6 13 0 15 9 1 10 9 2 3 9 13 0 9 2
9 9 1 0 9 14 13 3 9 2
25 10 9 1 9 1 0 9 1 9 1 0 9 3 13 3 6 15 13 9 7 9 1 0 9 2
26 15 13 0 2 3 9 1 9 1 9 1 0 9 3 15 13 1 9 1 0 9 1 9 1 9 2
42 2 0 13 0 0 0 9 2 9 1 9 1 3 2 9 1 0 0 0 9 2 1 15 3 15 13 9 7 9 7 10 9 2 15 13 9 7 13 1 15 9 2
10 15 15 13 6 13 9 7 0 9 2
14 9 13 2 16 0 9 3 13 6 15 13 1 9 2
14 0 9 1 9 13 9 9 6 4 13 1 0 9 2
13 13 9 9 6 13 9 1 9 7 0 0 9 2
23 0 0 9 2 1 9 1 9 1 9 1 11 2 4 13 3 1 0 9 1 0 9 2
3 0 9 2
3 0 9 2
15 3 9 15 13 1 9 1 0 9 2 0 1 9 9 2
20 1 15 9 13 3 0 2 16 9 14 13 9 1 9 2 16 3 15 13 2
29 2 6 6 4 13 1 14 12 1 9 1 9 2 6 6 13 14 9 2 14 0 9 2 14 6 13 0 9 2
8 1 9 15 13 9 1 9 2
17 9 13 9 1 9 1 9 1 9 15 1 0 9 7 2 9 2
28 9 1 9 1 0 9 1 9 1 0 9 7 9 1 9 7 9 1 0 9 13 0 1 9 1 0 9 2
13 3 9 1 9 14 13 10 0 9 6 15 13 2
18 3 7 3 0 9 13 2 16 9 1 9 13 1 9 1 0 9 2
17 16 10 9 13 9 2 15 13 1 9 1 0 15 9 1 9 2
11 0 13 3 15 6 13 3 0 7 0 2
22 9 1 9 1 0 9 13 1 0 9 1 0 9 2 7 13 13 7 1 0 9 2
9 6 2 6 2 2 13 15 15 2
10 14 7 9 13 9 15 2 3 0 2
26 14 2 13 2 13 15 2 3 16 15 2 9 2 13 1 9 3 1 9 7 1 9 6 15 13 2
21 9 14 4 13 1 0 9 2 1 9 1 9 7 9 1 9 7 9 1 9 2
12 13 13 3 2 3 3 2 15 13 1 9 2
19 1 9 1 9 3 15 13 10 2 15 4 13 6 13 9 1 0 9 2
16 15 13 9 2 13 1 0 9 7 13 12 9 3 1 9 2
6 13 15 7 15 13 2
27 16 6 13 14 3 15 4 13 2 9 3 6 13 0 2 7 14 9 15 1 9 15 13 1 9 15 2
4 15 4 13 2
8 15 13 15 0 1 10 9 2
20 9 1 0 9 1 9 1 9 13 0 9 7 14 4 13 3 1 0 9 2
11 0 9 1 0 9 15 13 1 0 9 2
33 13 15 3 1 0 9 2 16 15 13 1 9 1 0 9 7 0 9 2 7 1 10 9 15 13 9 1 9 1 10 0 9 2
10 15 13 0 9 1 9 1 0 9 2
11 2 13 15 2 3 3 13 7 3 9 2
8 7 15 13 0 2 13 15 2
8 7 15 13 0 2 13 15 2
33 7 1 9 1 9 2 15 13 9 1 15 2 15 3 13 3 15 13 9 1 0 9 7 3 10 9 14 4 13 7 1 11 2
44 1 15 3 1 9 1 9 7 1 9 1 9 2 9 7 9 1 9 1 9 1 0 11 3 3 15 13 9 2 13 15 10 2 15 11 13 14 13 7 14 13 1 9 2
15 9 1 0 9 1 10 9 1 9 1 0 9 1 11 2
9 7 13 14 15 13 14 15 13 2
35 0 0 9 13 11 2 15 9 2 14 13 0 9 1 0 11 2 14 13 9 1 0 11 2 3 16 9 1 0 11 14 13 10 9 2
8 15 2 13 15 2 13 0 2
2 9 2
3 13 3 2
10 13 15 9 2 13 1 9 7 3 2
15 10 0 9 13 0 2 13 15 2 3 1 10 0 9 2
14 16 9 13 0 2 13 9 1 15 3 1 0 9 2
16 9 13 0 9 1 9 15 2 1 1 9 15 15 4 13 2
20 1 0 9 9 13 9 1 9 7 9 2 1 15 9 13 9 7 9 15 2
5 1 9 13 9 2
17 3 2 10 9 15 13 3 7 3 1 15 15 13 14 15 13 2
8 0 1 9 13 9 1 9 2
7 10 9 13 1 10 9 2
12 9 13 2 7 15 15 13 3 1 0 9 2
5 3 13 10 9 2
4 13 0 9 2
6 9 13 1 0 9 2
11 1 9 15 13 9 1 9 7 0 9 2
13 1 10 9 2 0 1 9 2 9 15 13 3 2
7 9 13 10 9 1 9 2
8 9 2 3 9 2 13 9 2
17 9 13 14 13 14 13 1 9 2 1 9 2 1 14 13 9 2
9 9 1 9 15 13 14 15 13 2
19 9 1 9 2 3 1 0 9 2 13 3 0 7 13 3 14 15 13 2
16 1 15 9 15 13 14 13 15 2 7 6 4 13 3 15 2
12 15 13 1 9 1 9 2 1 14 13 9 2
5 9 13 3 0 2
16 10 9 2 15 13 14 13 3 15 2 1 9 6 13 15 2
7 9 13 3 9 1 9 2
6 1 9 3 15 13 2
7 13 7 13 1 0 9 2
11 9 15 13 0 9 2 0 9 15 13 2
7 3 0 13 9 1 9 2
13 3 13 1 15 2 13 2 16 4 13 3 3 2
7 0 1 9 9 13 0 2
10 1 3 9 9 13 9 14 15 13 2
11 0 9 6 13 2 3 0 13 1 15 2
21 9 13 0 9 1 9 7 3 13 3 1 0 9 2 13 0 15 9 7 9 2
13 7 3 13 9 15 1 9 2 15 4 3 0 2
7 9 13 0 9 1 9 2
12 15 13 9 14 13 9 7 9 14 15 13 2
19 1 10 9 2 0 1 9 2 6 13 7 9 2 7 9 2 7 9 2
7 0 6 13 14 13 0 2
19 9 1 10 0 9 2 3 1 10 0 9 2 6 15 13 1 12 9 2
5 9 13 1 0 2
8 3 7 10 0 9 13 0 2
7 9 7 1 9 13 9 2
9 10 9 6 13 0 1 10 9 2
7 0 9 13 7 0 9 2
13 6 2 10 9 13 3 0 2 15 13 3 0 2
10 15 15 13 2 13 2 13 7 13 2
2 9 2
4 13 4 9 2
6 9 13 1 3 9 2
16 9 13 2 13 2 9 2 3 9 3 13 14 13 9 15 2
7 0 9 1 9 13 9 2
5 3 13 1 15 2
12 9 1 10 9 13 1 9 1 9 10 9 2
12 9 15 13 1 9 2 15 15 13 14 13 2
8 1 10 9 13 3 10 9 2
7 9 13 0 1 9 15 2
7 3 7 9 15 15 13 2
9 0 13 0 1 0 9 7 9 2
15 16 0 9 15 13 1 9 2 9 15 15 13 1 9 2
9 3 15 15 13 2 9 4 13 2
12 16 9 13 0 2 13 14 15 13 1 15 2
8 14 9 1 9 1 0 9 2
13 1 9 2 3 15 13 9 2 9 13 3 0 2
6 9 1 9 1 9 2
9 6 4 13 14 13 9 1 9 2
4 13 15 9 2
8 3 13 13 13 7 3 9 2
6 10 0 9 13 0 2
4 9 13 9 2
18 9 2 10 0 9 2 3 9 13 1 9 7 13 14 13 1 9 2
16 3 0 9 13 1 9 2 0 1 9 2 1 15 13 9 2
10 10 9 6 13 3 1 9 1 9 2
18 11 13 1 9 7 13 1 9 2 3 9 15 13 7 13 9 15 2
26 6 15 13 2 13 15 3 1 15 14 1 9 15 7 1 14 13 9 15 2 13 3 2 2 13 2
22 2 6 2 2 13 3 0 9 1 11 2 3 10 9 2 3 3 15 13 14 13 2
61 15 3 6 15 13 2 1 9 15 13 3 0 15 9 2 9 1 0 7 0 15 9 2 0 15 7 0 9 2 9 1 9 15 2 9 15 2 9 15 2 15 3 6 13 2 16 6 15 13 10 3 0 9 2 10 3 0 9 7 9 2
31 15 13 14 9 15 2 9 1 9 15 2 9 1 9 15 2 0 7 0 9 2 9 2 9 2 0 15 9 7 0 2
2 3 2
3 13 15 2
3 1 9 2
5 1 10 7 10 2
4 1 0 9 2
4 1 0 9 2
6 13 14 14 15 13 2
6 11 2 11 7 11 2
4 16 15 13 2
4 9 15 13 2
20 13 9 15 2 13 15 1 9 7 3 13 1 9 2 1 14 15 13 9 2
13 13 2 3 6 13 9 7 15 13 1 9 15 2
9 11 2 0 1 9 2 13 15 2
15 7 6 4 14 15 15 13 2 3 9 13 15 7 9 2
11 15 4 13 15 2 11 4 13 2 9 2
8 6 13 14 15 13 1 15 2
4 13 15 15 2
2 2 3
6 2 6 15 13 9 2
8 2 13 14 15 13 15 2 2
8 3 13 7 15 13 1 15 2
8 2 13 14 15 13 3 9 2
4 13 15 3 2
4 2 15 2 2
8 9 2 9 2 15 14 13 2
15 13 15 15 3 2 1 9 2 3 15 13 1 9 15 2
18 13 15 2 16 13 14 13 0 1 15 7 15 13 3 1 9 15 2
10 6 13 9 2 15 13 1 9 15 2
9 3 1 0 9 13 2 6 13 2
12 13 1 9 2 11 6 15 13 1 9 15 2
3 6 13 2
6 1 9 15 13 9 2
5 0 2 0 9 2
3 0 3 2
2 3 2
24 9 15 13 9 15 2 6 13 14 13 7 9 2 9 15 4 13 2 7 13 9 1 9 2
6 2 9 1 11 13 2
4 2 13 15 2
10 13 9 1 15 7 13 1 0 9 2
20 15 13 1 15 2 13 15 3 2 1 14 13 11 7 15 13 1 15 12 2
4 2 13 15 2
7 15 15 4 13 2 0 2
9 9 15 2 9 2 0 15 9 2
3 13 15 2
9 15 6 13 1 10 4 15 13 2
3 13 15 2
6 2 6 13 1 9 2
14 13 15 11 7 15 13 3 2 15 13 14 15 13 2
9 3 3 13 9 2 14 15 13 2
25 6 15 13 1 9 15 2 13 9 15 1 9 15 2 9 15 13 9 15 2 7 15 15 13 2
6 2 13 15 2 0 2
3 13 15 2
4 7 15 13 2
8 6 15 15 4 13 12 9 2
8 14 3 15 13 14 15 13 2
7 13 7 15 13 1 11 2
5 2 3 14 13 2
12 3 13 14 15 13 2 7 3 15 2 13 2
4 3 14 13 2
6 2 3 6 4 13 3
9 2 13 15 15 2 13 3 9 2
7 9 13 3 1 9 15 2
16 13 15 1 15 2 9 15 15 13 2 13 9 1 15 14 2
6 2 13 14 15 13 2
11 13 1 11 7 11 7 15 3 15 13 2
7 2 15 14 15 13 14 2
3 2 3 2
6 2 13 1 9 11 2
3 2 3 2
9 2 15 12 4 13 14 13 0 9
4 2 1 10 2
5 2 13 15 11 2
13 11 15 13 2 6 15 13 9 15 1 10 9 2
4 3 2 3 2
7 2 13 14 13 0 9 2
5 15 12 7 15 2
9 11 15 13 7 3 13 1 9 2
17 13 2 13 15 14 6 13 1 9 7 9 2 13 14 15 13 2
7 9 15 6 13 1 9 2
7 15 0 9 4 13 9 2
9 7 3 3 15 2 3 13 0 2
4 9 2 7 2
2 6 2
9 13 2 16 13 9 1 15 14 2
14 1 0 0 9 0 1 9 11 15 13 14 15 13 2
7 13 14 15 1 9 15 2
10 3 13 14 13 9 15 7 14 13 2
5 2 6 2 9 2
9 13 4 15 7 3 14 15 13 2
4 14 1 11 2
8 9 1 0 15 13 1 9 2
8 2 7 7 11 2 3 13 2
6 7 1 15 15 13 2
26 9 2 3 0 9 2 9 1 12 7 9 1 0 2 9 1 9 1 9 15 2 3 15 4 13 2
4 9 2 9 2
21 15 13 14 15 13 3 2 7 6 13 14 13 0 2 6 13 14 13 9 15 2
8 7 3 6 13 9 1 9 2
4 6 13 14 2
7 1 0 9 6 4 13 2
6 7 15 13 14 13 2
4 3 2 3 2
3 6 3 2
6 3 13 14 13 15 2
9 1 9 2 1 9 2 1 9 2
16 16 13 1 11 15 13 2 9 13 2 16 13 9 1 9 2
6 3 15 13 7 9 2
11 9 2 0 9 2 9 7 9 2 9 2
2 13 2
7 11 13 7 3 15 13 2
8 13 14 14 15 13 1 9 2
9 2 14 13 2 15 6 15 13 2
11 2 14 13 2 13 15 11 2 2 9 2
6 7 3 6 13 15 2
6 13 14 15 15 9 2
16 11 13 7 0 3 2 13 1 9 1 15 7 3 13 9 2
6 13 9 1 0 9 2
19 11 13 1 9 15 2 13 15 1 15 7 15 13 1 0 15 0 9 2
6 2 9 2 15 13 2
7 2 7 3 6 13 0 2
11 13 2 6 2 16 10 9 4 13 3 2
11 1 14 13 0 2 13 14 13 1 0 2
5 14 13 1 0 2
5 14 13 1 0 2
14 14 13 9 15 3 3 7 14 13 9 15 3 3 2
3 0 9 2
8 0 9 2 1 14 15 13 2
8 3 2 7 13 3 7 3 2
21 9 1 9 1 0 15 15 13 2 3 15 4 13 1 9 7 3 15 4 13 2
6 3 13 3 1 15 2
3 13 15 2
12 13 14 13 9 2 1 14 13 9 7 9 2
18 10 9 4 13 1 3 7 3 9 2 16 15 13 1 3 15 14 2
5 15 3 15 13 2
9 1 12 15 9 15 13 0 9 2
5 2 13 14 15 13
14 0 2 0 9 2 15 16 16 14 13 1 9 15 2
7 3 2 3 2 1 9 2
4 2 1 3 2
18 13 14 15 13 3 2 4 13 1 9 15 7 15 13 9 1 9 2
11 14 15 13 2 16 14 13 0 1 15 2
10 14 15 13 9 2 16 3 15 13 2
10 13 0 9 7 6 15 13 1 15 2
32 7 13 0 2 1 9 1 9 15 2 1 0 9 2 0 7 0 1 0 15 9 2 1 15 4 13 14 13 14 9 15 2
9 3 14 13 9 14 13 3 15 2
6 13 2 3 6 13 2
13 13 1 9 1 11 7 15 13 9 1 1 9 2
7 13 14 13 9 1 9 2
2 11 11
3 9 1 9
9 2 15 6 15 13 1 15 2 2
5 2 15 13 15 2
5 2 13 15 11 2
14 15 13 1 9 2 0 9 1 0 9 1 0 9 2
20 9 15 4 13 1 9 2 3 1 0 9 1 0 9 13 0 9 1 9 2
35 15 15 13 2 13 3 2 13 9 1 0 2 0 9 2 9 1 9 7 0 9 13 9 7 9 13 3 2 3 2 1 0 0 9 2
5 13 7 15 13 2
13 2 15 13 9 1 9 7 10 9 15 13 9 2
13 15 13 0 9 1 0 9 7 0 1 9 9 2
10 2 13 11 7 3 15 13 1 9 2
12 2 6 2 15 14 13 1 10 9 7 9 2
3 13 15 2
4 11 15 13 2
15 2 15 13 9 1 10 3 7 1 9 13 14 15 13 2
7 15 13 0 2 0 9 2
5 11 3 15 13 2
11 2 6 2 6 2 15 6 13 3 3 2
7 13 15 15 3 9 15 2
4 2 9 15 2
2 14 2
6 2 15 3 14 13 2
3 2 13 2
17 9 15 13 2 3 13 12 9 2 7 0 9 1 11 15 13 2
3 2 14 2
6 9 13 7 15 13 2
7 2 7 15 3 15 13 2
5 11 3 15 13 2
2 11 2
6 2 15 3 14 13 2
10 15 14 15 13 0 2 3 0 9 2
10 9 13 3 12 9 7 15 13 3 2
7 2 13 0 15 0 9 2
14 7 15 13 3 0 2 3 13 14 15 13 3 3 2
12 7 1 0 9 15 4 13 1 3 0 9 2
10 1 10 12 9 11 13 10 0 9 2
8 2 0 9 2 12 9 3 2
9 3 3 12 9 7 15 14 13 2
4 9 13 9 2
4 2 9 14 2
2 6 2
5 15 13 3 0 2
7 11 15 13 3 2 3 2
7 2 15 6 13 3 0 2
6 2 3 2 0 2 2
2 7 2
10 0 14 13 2 3 9 7 9 15 2
4 2 14 13 2
3 13 15 2
5 15 13 3 3 2
20 7 3 1 9 15 13 9 2 9 15 13 1 0 9 7 9 15 15 13 2
19 13 2 7 14 9 6 13 1 9 15 2 15 13 0 2 0 2 0 2
5 2 15 13 15 2
12 2 15 13 9 1 9 7 9 15 13 9 2
2 9 0
2 0 9
1 9
19 10 9 13 9 2 0 1 9 2 9 7 9 1 0 9 7 0 9 2
31 9 1 10 9 15 13 7 1 9 1 0 9 7 0 9 1 9 2 15 13 1 0 9 2 1 15 9 13 9 11 2
25 1 0 9 7 0 9 1 0 9 10 9 15 13 1 9 1 9 2 15 15 13 1 0 9 2
13 9 1 9 7 0 9 13 1 9 1 9 15 2
18 9 2 15 4 13 9 7 0 9 2 0 1 9 2 13 10 9 2
20 9 1 9 2 9 2 1 9 1 9 7 0 9 13 1 9 2 9 2 2
26 9 1 9 7 1 0 9 13 9 14 4 13 1 9 2 1 9 7 1 9 1 9 7 0 9 2
1 9
19 9 1 0 9 2 0 1 10 9 2 15 13 1 9 1 0 0 9 2
3 9 1 9
1 9
2 0 9
3 0 0 9
14 9 15 13 1 0 9 2 15 13 0 7 3 0 2
1 9
4 9 7 0 9
17 9 7 0 9 1 0 9 15 13 1 9 1 9 0 7 0 2
2 0 9
24 0 9 1 0 9 15 13 1 9 2 15 13 9 1 9 12 9 2 0 1 9 1 9 2
19 9 1 9 15 13 7 1 0 9 2 3 1 10 9 6 4 13 0 2
2 9 0
2 0 9
7 11 13 9 1 0 9 2
7 0 0 9 13 1 9 2
15 15 15 13 1 15 3 7 1 9 2 0 1 10 11 2
26 10 9 1 9 2 0 9 7 0 9 2 0 9 7 0 9 6 13 14 15 13 9 1 0 9 2
9 9 11 13 0 9 1 0 9 2
7 0 9 1 9 13 0 2
6 9 11 13 0 9 2
10 15 15 13 1 11 7 9 1 9 2
23 9 11 13 9 2 9 7 9 1 9 7 13 9 1 0 9 1 9 7 1 0 9 2
13 11 13 0 9 7 0 9 6 13 14 15 13 2
7 9 1 11 13 0 9 2
14 15 13 9 1 10 9 1 0 9 2 15 15 13 2
6 10 0 9 15 13 2
7 10 9 13 0 1 9 2
40 6 15 13 10 9 1 9 7 9 2 0 1 9 2 9 2 0 9 2 9 2 9 2 9 2 9 2 9 2 0 9 2 0 7 0 9 7 0 9 2
18 9 13 1 9 2 0 1 0 9 7 9 1 10 9 7 0 9 2
16 0 9 13 9 2 9 7 9 1 9 7 13 10 0 9 2
22 9 2 0 7 0 9 15 13 1 9 1 0 2 0 7 0 0 9 1 0 9 2
13 0 9 1 9 11 15 13 1 9 1 0 9 2
16 14 10 0 9 7 9 6 13 14 15 13 7 13 1 0 2
12 9 13 1 9 7 9 1 0 9 1 9 2
4 9 13 0 2
7 0 9 4 13 1 9 2
18 0 9 7 9 2 3 7 0 9 6 13 14 15 13 1 0 9 2
13 9 2 9 7 9 13 1 9 1 9 7 9 2
27 9 11 13 9 7 9 1 0 9 2 9 7 9 1 0 9 7 0 9 1 0 9 7 9 1 9 2
8 9 15 13 7 13 1 9 2
13 9 1 9 7 1 9 15 13 7 13 1 9 2
6 9 13 0 7 0 2
35 0 9 2 0 0 9 2 0 9 2 3 7 9 2 9 7 9 1 0 9 2 0 7 0 9 2 0 1 9 2 13 0 0 9 2
34 9 13 0 9 1 0 9 7 1 0 0 9 1 9 2 9 2 9 2 9 7 9 1 0 2 0 7 0 9 1 10 0 9 2
21 9 13 0 9 1 0 9 7 9 1 0 9 2 0 1 9 11 1 0 9 2
14 0 9 15 13 7 13 1 9 1 9 7 1 9 2
11 9 1 9 11 15 13 1 0 0 9 2
17 9 7 0 9 1 0 7 0 9 7 0 9 15 13 1 9 2
23 9 13 9 1 9 7 0 9 1 9 1 9 7 0 9 1 9 1 0 7 0 9 2
25 9 13 9 1 0 9 1 0 9 1 9 7 13 0 9 7 9 1 0 2 0 7 0 9 2
20 9 7 0 0 9 6 13 14 13 9 1 9 1 9 1 1 9 1 9 2
10 1 10 9 15 13 14 13 9 15 2
25 1 0 1 9 9 9 7 0 0 9 13 14 13 9 1 9 2 9 1 9 7 0 0 9 2
16 9 13 9 1 0 9 1 9 2 9 7 9 7 15 13 2
12 15 15 13 1 9 1 0 0 7 0 9 2
17 0 9 1 9 11 15 13 1 9 1 9 7 9 1 0 9 2
36 0 9 1 0 9 1 9 11 13 0 9 7 9 1 9 2 9 7 0 9 7 9 1 0 9 2 3 7 9 1 9 1 0 0 9 2
2 9 0
11 9 1 0 9 13 0 9 1 0 9 2
13 0 9 1 9 6 13 14 4 13 1 0 9 2
14 0 9 2 0 1 9 2 13 1 9 1 9 11 2
17 9 7 9 1 9 2 9 7 9 1 0 9 15 13 1 9 2
20 9 1 9 11 2 3 7 14 15 13 2 13 10 9 7 9 1 10 11 2
32 9 2 15 13 1 9 11 2 13 10 9 7 9 1 10 11 1 9 1 9 7 9 2 1 15 11 7 9 13 0 9 2
12 9 7 9 1 9 1 9 15 13 1 9 2
6 15 13 9 1 9 2
19 15 6 13 14 4 13 1 0 2 0 7 0 9 1 10 0 0 9 2
9 15 13 9 1 0 9 7 9 2
17 1 9 1 12 9 1 9 9 1 0 9 15 13 1 10 9 2
18 15 13 9 1 0 9 1 9 1 9 15 7 1 9 15 1 9 2
7 9 1 10 9 13 0 2
15 9 15 13 1 0 1 9 1 0 1 0 1 9 9 2
23 1 0 1 9 15 13 9 1 9 1 0 15 9 2 15 6 4 13 1 9 1 9 2
14 9 9 1 9 15 13 3 1 9 2 0 1 9 2
26 15 13 9 1 9 1 0 9 1 0 7 0 15 9 7 1 9 1 10 9 2 9 7 0 9 2
4 9 13 0 2
24 1 9 1 9 15 15 6 13 14 13 7 14 13 1 15 1 1 9 2 3 0 1 9 2
12 9 7 9 1 9 7 1 0 9 13 0 2
25 9 1 10 9 15 13 3 1 9 1 0 9 2 3 15 15 13 1 9 7 9 1 0 9 2
26 10 9 13 14 15 13 3 1 9 2 1 9 1 0 9 2 0 9 7 9 7 9 1 0 9 2
11 10 0 9 13 9 14 15 13 1 9 2
14 9 7 9 1 0 9 13 9 7 9 1 0 9 2
20 9 1 9 2 9 1 9 7 9 1 9 7 1 0 7 0 9 13 0 2
21 9 13 1 9 1 9 7 9 1 0 1 0 9 2 3 7 1 0 7 0 2
15 9 7 0 9 1 0 9 13 0 7 6 13 1 9 2
48 9 7 9 1 0 9 7 1 0 9 1 9 15 13 3 1 9 1 0 9 2 3 15 13 0 9 7 15 13 9 1 0 9 1 3 0 9 2 1 9 1 9 7 1 9 1 9 2
15 16 1 9 1 12 9 6 13 9 2 9 13 9 15 2
11 15 13 9 14 13 2 13 7 13 9 2
14 9 7 9 1 9 1 9 7 9 15 13 1 9 2
15 9 13 9 14 15 13 3 7 1 9 1 9 7 9 2
7 9 13 3 14 15 13 2
62 13 15 9 2 10 9 4 13 1 9 2 0 9 1 9 7 9 1 9 2 1 9 1 0 2 0 2 0 7 0 9 2 1 9 1 9 7 9 1 9 2 3 7 9 2 15 13 0 7 0 9 2 7 15 13 14 13 9 15 1 9 2
21 9 13 9 2 15 13 1 9 2 9 1 10 9 2 3 7 9 15 1 9 2
13 9 13 9 1 9 2 9 7 9 1 0 9 2
9 9 13 0 9 1 9 7 9 2
6 0 13 3 0 9 2
11 9 13 0 9 7 9 1 9 7 9 2
24 9 1 9 2 9 7 9 1 10 9 7 9 2 0 7 0 9 1 9 15 13 1 9 2
19 9 2 0 1 9 1 0 15 2 15 13 1 0 9 1 9 7 9 2
15 9 7 9 1 9 7 9 1 0 9 15 13 1 9 2
6 9 13 9 1 9 2
13 9 15 13 1 9 1 9 1 9 1 10 9 2
17 9 13 9 1 9 1 9 1 9 1 9 1 0 7 0 9 2
11 10 9 3 13 10 9 7 9 1 9 2
11 15 6 13 14 4 13 14 13 0 9 2
2 9 0
9 0 9 15 13 1 12 0 9 2
10 0 9 15 13 1 9 1 12 9 2
17 9 1 0 9 2 15 13 0 9 2 13 9 15 1 9 15 2
7 9 1 0 9 13 3 2
18 0 9 2 0 1 9 2 13 9 15 1 9 2 1 15 13 9 2
12 1 10 9 15 15 13 1 0 1 9 9 2
19 0 9 6 13 0 9 1 0 1 15 9 7 1 9 15 1 0 9 2
13 0 9 13 9 2 10 9 15 13 1 0 9 2
20 16 1 0 9 9 6 13 0 9 2 15 15 13 1 12 0 1 0 9 2
13 0 9 1 0 9 15 13 1 0 0 0 9 2
9 1 0 9 0 9 13 0 9 2
3 13 15 2
12 1 0 9 1 0 9 15 13 9 7 9 2
14 9 1 0 9 13 9 7 13 0 15 1 15 9 2
9 0 9 15 13 1 9 7 9 2
24 0 9 13 9 7 0 9 1 9 3 1 9 1 0 0 9 2 1 3 11 13 0 9 2
13 1 9 0 9 13 14 13 0 9 14 4 13 2
9 1 10 9 15 15 13 1 9 2
11 0 9 13 9 2 9 2 9 7 9 2
17 9 7 9 1 0 9 13 0 1 10 0 9 2 9 7 9 2
12 9 1 0 9 13 10 0 9 7 0 9 2
12 9 1 0 9 15 13 7 13 1 0 9 2
16 9 15 13 7 13 1 12 9 2 15 15 13 1 0 9 2
16 1 9 0 9 13 14 13 12 9 14 15 13 1 12 9 2
17 9 4 13 2 3 1 15 4 13 3 1 9 1 10 0 9 2
18 3 0 9 13 9 1 9 7 1 0 9 2 9 13 9 1 9 2
17 1 9 1 12 0 1 0 9 1 9 13 9 7 15 13 9 2
14 0 9 13 0 9 2 15 13 9 1 9 1 9 2
15 9 2 9 7 9 1 9 1 0 9 15 13 1 9 2
15 0 9 13 3 9 1 9 3 1 9 1 10 0 9 2
17 3 0 1 0 9 9 15 13 1 9 1 0 9 1 9 15 2
14 1 9 1 10 9 9 13 9 2 13 9 7 9 2
16 0 9 13 9 1 9 7 9 1 0 9 1 9 1 9 2
22 16 4 13 2 16 9 7 9 4 13 0 9 7 4 13 11 2 9 15 15 13 2
2 9 0
2 0 9
18 0 9 13 7 13 0 7 0 9 1 9 1 9 1 11 7 9 2
20 0 9 13 0 9 7 0 9 7 13 0 9 1 0 9 7 1 0 9 2
28 0 9 13 9 1 0 9 2 13 9 1 0 9 2 13 2 13 7 13 0 9 1 9 2 0 1 9 2
10 0 9 13 0 7 0 9 1 9 2
11 9 13 0 9 1 16 0 9 13 0 2
7 15 13 9 1 10 9 2
9 0 9 13 9 1 0 0 9 2
17 1 9 1 0 9 0 9 13 9 15 1 9 1 0 0 9 2
22 0 9 13 14 13 0 9 14 15 13 9 1 0 9 2 1 9 7 1 0 9 2
13 9 15 13 1 9 3 1 9 1 0 0 9 2
14 3 0 9 6 13 0 9 2 9 13 9 1 9 2
16 1 9 7 1 9 1 9 0 9 13 9 2 9 7 9 2
11 0 9 13 9 1 9 7 9 1 9 2
2 9 0
6 9 7 9 1 11 2
4 9 1 0 11
20 9 1 9 1 9 7 9 1 11 13 1 12 9 1 0 9 7 1 9 2
21 9 15 13 1 0 9 6 3 1 12 9 7 6 3 1 12 9 1 9 15 2
25 0 9 13 9 1 9 7 9 1 11 1 9 12 9 1 10 0 9 1 12 9 1 0 9 2
29 9 1 9 7 9 1 11 15 13 7 15 13 1 9 1 0 9 1 2 0 9 2 1 0 9 1 9 15 2
16 9 13 9 1 0 0 9 1 0 9 1 9 1 0 9 2
15 1 9 1 9 1 0 0 9 9 1 0 9 15 13 2
23 0 0 9 13 9 1 0 9 1 9 12 0 1 10 0 9 1 12 9 1 0 9 2
15 0 0 9 13 3 10 9 1 11 2 1 15 4 13 2
13 1 0 9 0 0 9 13 9 7 1 0 9 2
13 1 10 9 9 13 9 1 9 2 0 1 9 2
19 9 1 0 0 9 15 13 7 13 1 10 9 1 0 9 1 9 15 2
2 9 0
10 1 0 9 4 13 9 1 9 11 2
19 9 2 1 15 15 13 0 9 7 15 13 0 9 2 15 13 1 9 2
11 9 1 9 11 13 9 2 0 9 2 2
8 9 1 9 11 13 9 11 2
30 3 7 14 13 3 2 12 9 1 9 2 7 3 2 3 12 9 1 9 2 2 10 9 9 14 13 9 1 11 2
4 1 9 6 2
12 3 3 15 13 9 1 11 11 7 11 11 2
23 7 3 12 13 3 3 15 13 2 16 1 12 9 0 9 14 4 13 1 9 1 9 2
11 1 12 9 9 13 9 1 0 0 11 2
6 11 2 9 1 0 9
24 10 9 15 13 3 3 2 3 11 11 7 11 11 13 9 1 9 1 11 7 1 0 9 2
32 3 0 1 10 9 1 9 1 9 7 9 15 0 9 15 13 1 10 9 1 10 9 2 7 14 7 1 9 1 0 11 2
21 10 9 13 1 3 0 9 1 7 1 9 1 0 1 9 9 1 9 1 11 2
19 1 11 1 0 9 15 13 3 3 12 13 14 13 10 9 1 10 9 2
9 1 9 13 3 14 15 13 9 2
28 1 0 11 3 13 9 1 11 2 3 9 1 9 7 9 1 9 13 0 9 1 9 1 9 1 0 9 2
10 3 11 7 11 6 13 14 15 13 2
31 7 1 9 10 0 9 14 15 13 1 9 1 0 2 7 9 3 14 13 6 1 9 7 9 2 7 1 0 7 0 2
3 9 1 9
14 3 1 0 0 9 1 0 9 0 9 14 13 9 2
38 9 1 9 1 9 1 9 1 0 9 13 9 2 3 16 1 3 0 9 4 13 2 7 7 1 9 1 0 9 1 11 14 15 13 3 0 9 2
23 1 0 9 9 1 0 9 14 15 13 1 12 9 7 12 0 9 2 15 3 13 9 2
28 9 1 0 9 7 0 9 2 9 7 0 9 2 9 2 0 7 9 2 9 7 9 13 1 9 1 9 2
15 1 0 9 14 4 13 9 1 9 1 9 7 0 9 2
33 14 9 1 10 9 14 15 13 7 1 9 1 11 2 15 6 13 3 0 1 15 2 1 14 15 13 0 9 14 13 0 9 2
24 0 9 1 9 1 9 1 9 13 9 1 9 1 11 2 0 1 11 2 7 12 0 9 2
14 3 11 2 11 2 11 7 11 14 13 1 12 9 2
11 0 9 9 13 11 7 11 2 1 12 2
14 11 2 11 2 11 2 11 7 11 14 13 1 12 2
16 11 2 11 7 11 14 13 1 1 12 9 1 9 1 9 2
15 11 2 11 2 11 2 11 7 11 14 13 1 12 9 2
39 0 9 13 3 1 10 2 16 1 9 1 9 10 0 9 14 13 1 9 14 13 1 0 9 2 7 14 13 9 1 9 2 14 14 13 0 9 9 2
20 1 0 9 11 2 11 2 11 2 11 7 11 14 13 0 15 9 1 11 2
25 13 15 1 9 14 13 0 9 1 9 1 0 9 1 11 2 15 13 14 13 0 1 10 9 2
22 0 9 3 3 13 9 1 9 1 9 1 9 2 16 15 14 13 9 14 13 9 2
5 12 7 12 7 13
8 9 2 11 11 2 2 11 2
14 1 9 1 15 11 4 13 14 13 1 2 9 2 2
14 3 1 0 9 11 13 1 12 9 9 3 1 11 2
10 15 13 9 15 14 13 0 1 9 2
23 1 0 9 1 12 0 9 15 13 1 10 9 1 9 1 0 9 1 9 1 0 11 2
6 7 15 3 13 9 2
21 1 11 2 11 7 11 1 10 9 2 3 15 14 13 9 2 13 0 11 11 2
14 9 1 11 3 13 0 9 1 9 1 9 7 9 2
29 0 9 15 13 12 9 1 12 9 2 12 2 11 2 2 9 2 9 2 0 9 2 9 2 9 2 9 2 2
17 0 14 13 9 1 11 1 0 9 2 7 1 15 3 13 9 2
26 1 0 9 1 9 1 11 1 0 11 15 13 0 9 10 9 14 13 0 9 1 9 1 0 9 2
13 11 11 4 13 2 16 9 14 13 1 0 9 2
15 7 9 1 11 11 11 14 6 13 0 9 1 0 9 2
14 7 3 10 9 13 0 9 1 9 1 9 1 9 2
40 1 9 1 0 0 9 2 1 9 1 9 1 0 9 7 1 9 1 3 0 15 9 11 3 13 10 9 6 3 1 9 1 0 9 1 9 2 0 9 2
12 7 11 3 13 14 13 9 3 1 9 15 2
28 1 10 9 1 0 1 0 9 0 9 11 13 3 0 9 1 0 9 1 9 14 15 13 3 1 0 9 2
16 11 13 1 0 9 1 0 9 2 7 1 9 1 0 9 2
20 0 0 9 2 0 0 9 1 0 9 1 9 2 4 13 3 1 12 9 2
24 3 11 14 4 13 1 12 9 1 9 1 9 1 11 2 15 3 13 14 4 13 1 9 2
2 0 9
3 11 11 11
17 7 9 2 7 9 2 7 9 1 9 2 7 9 1 0 9 2
6 0 9 7 0 9 2
9 0 9 1 9 2 9 7 9 2
2 9 2
4 9 1 9 2
4 9 1 9 2
13 7 10 9 7 9 1 0 9 7 1 0 9 2
9 13 9 2 15 4 13 14 13 2
9 13 9 2 15 4 13 14 13 2
9 16 13 9 3 2 14 13 15 2
9 16 13 9 3 2 14 13 9 2
31 16 13 1 9 2 14 13 1 9 1 9 1 9 2 1 9 2 1 9 2 14 1 9 1 9 2 15 15 13 9 2
2 3 2
5 10 9 13 9 2
6 6 13 14 15 13 2
5 0 9 13 9 2
8 7 9 6 13 14 13 15 2
8 15 13 3 1 9 7 0 2
11 3 13 1 0 9 7 13 9 1 9 2
13 13 9 7 13 9 2 1 15 14 13 9 15 2
9 10 2 1 10 0 9 1 9 2
9 7 10 9 2 10 9 13 9 2
6 9 6 13 3 0 2
13 0 9 2 7 13 3 14 13 1 9 7 9 2
19 7 1 1 15 13 2 14 15 13 1 3 9 0 2 1 3 9 0 2
5 13 15 0 9 2
12 3 0 2 0 2 0 1 0 9 7 9 2
12 14 13 9 1 9 2 1 14 13 9 15 2
6 3 13 14 13 0 2
14 14 15 13 1 0 9 7 14 15 13 1 0 9 2
5 9 13 14 13 2
5 2 14 13 9 2
4 7 13 9 2
9 14 13 1 9 2 14 13 1 9
22 15 13 1 9 7 15 13 2 16 13 3 0 2 3 15 15 13 14 15 13 0 2
6 3 3 13 3 0 2
9 15 13 14 15 14 15 13 0 2
2 6 2
6 3 15 13 0 9 2
28 1 10 9 14 13 9 3 14 15 13 3 3 1 9 2 14 16 15 13 9 2 0 9 7 9 1 9 2
8 3 4 15 13 1 0 9 2
14 3 3 6 15 4 13 10 15 13 1 9 1 9 2
20 3 4 15 13 1 1 9 1 9 1 9 7 4 4 13 1 0 1 15 2
5 9 6 13 9 2
4 15 13 15 2
13 13 9 1 0 1 11 2 11 2 11 7 11 2
13 13 14 2 16 12 0 1 9 1 9 13 0 2
13 1 3 9 9 13 9 2 9 2 0 1 9 2
5 3 4 13 11 2
14 7 16 13 1 9 2 13 3 14 13 15 13 0 2
22 3 9 15 13 9 2 15 13 9 2 16 9 3 14 15 13 10 9 1 9 15 2
10 12 9 15 13 1 0 9 1 9 2
4 14 13 9 2
2 6 2
13 16 6 13 14 13 1 9 2 13 0 15 9 2
20 3 13 12 9 3 1 10 2 15 15 13 10 9 2 3 9 15 15 13 2
16 1 15 0 9 1 9 1 0 9 13 14 15 13 3 3 2
27 9 15 2 1 7 1 9 2 13 1 15 2 3 14 13 14 13 9 1 14 15 13 15 14 15 13 2
8 0 9 1 9 1 9 1 9
5 7 9 13 9 2
8 3 16 13 14 13 1 9 2
3 7 15 2
29 7 6 13 9 15 2 7 13 14 15 13 2 3 16 2 3 15 13 2 14 13 2 2 1 10 9 13 2 2
9 13 14 15 13 3 1 12 9 2
15 0 9 1 12 13 14 15 13 14 15 13 1 0 9 2
3 13 9 2
11 9 1 9 1 9 15 13 1 0 9 2
8 14 6 13 1 0 0 9 2
3 6 13 2
3 13 15 2
9 13 9 1 9 7 13 0 9 2
17 13 15 14 15 13 1 9 1 0 9 7 15 13 1 0 9 2
40 3 13 1 0 9 1 9 1 9 11 2 13 9 9 14 15 13 1 9 2 9 2 9 2 0 9 2 0 9 2 9 2 9 2 9 2 9 7 9 2
18 13 1 9 0 9 2 1 15 13 9 3 2 1 14 13 1 9 2
9 1 14 13 9 2 13 9 3 2
2 3 2
6 13 3 0 14 13 2
5 13 9 1 9 2
6 3 13 2 3 13 2
12 3 15 13 1 0 2 13 15 7 15 13 2
33 9 13 3 3 2 16 13 9 1 9 7 3 16 14 15 15 13 14 15 13 1 9 7 1 9 15 2 3 13 14 13 3 2
7 13 0 7 0 15 9 2
9 13 0 1 9 2 13 14 3 2
5 6 13 14 13 2
13 13 15 2 16 15 13 9 1 9 1 0 9 2
10 7 15 13 2 16 13 9 1 9 2
10 16 9 15 15 13 2 9 15 13 2
21 6 2 13 14 13 0 2 7 15 13 2 16 6 4 13 9 15 1 0 9 2
6 13 1 9 1 9 2
16 3 15 13 1 10 9 2 3 16 13 14 13 0 0 9 2
4 10 9 13 2
6 3 6 15 13 3 2
7 13 14 13 1 15 14 2
18 3 13 14 15 13 1 9 9 2 16 14 6 13 0 9 1 9 2
16 9 13 2 16 1 9 1 0 0 9 4 13 2 16 13 2
9 13 2 16 9 7 9 13 0 2
22 16 15 13 2 10 9 3 14 15 13 9 2 7 1 10 9 14 15 13 7 13 2
20 4 13 3 1 10 3 0 9 2 13 15 2 16 9 13 9 1 9 15 2
3 13 9 2
8 10 9 13 14 15 13 3 2
23 1 9 3 13 1 9 2 13 1 0 9 7 1 9 2 1 14 13 15 1 0 15 2
8 13 3 15 13 3 14 13 2
8 13 2 3 13 1 0 9 2
14 16 6 13 3 3 1 9 2 13 15 7 13 3 2
15 16 15 13 1 9 9 2 6 13 14 13 15 1 9 2
14 13 15 9 7 13 1 0 9 2 16 15 15 13 2
21 4 13 3 14 13 9 1 0 9 2 1 0 9 7 16 13 1 9 1 9 2
3 6 13 2
17 3 16 13 14 15 13 0 2 3 7 3 13 14 13 1 15 2
4 13 9 15 2
2 13 2
14 9 14 15 13 1 9 1 9 13 14 13 14 13 2
11 3 14 13 1 9 13 3 1 0 9 2
9 3 4 13 9 2 1 14 13 2
20 3 15 13 2 9 15 4 13 7 13 3 14 15 13 3 1 9 1 9 2
12 13 14 9 2 15 14 15 13 0 0 9 2
8 13 14 4 3 0 1 9 2
16 0 9 15 13 14 15 13 3 7 14 13 9 2 3 13 2
19 6 15 13 1 9 1 9 1 9 2 15 13 14 15 13 1 0 9 2
14 15 13 0 9 7 13 2 16 15 13 14 13 9 2
23 1 10 9 14 13 0 9 1 0 9 2 1 15 14 15 13 14 15 13 1 0 9 2
3 13 15 2
13 13 13 4 13 0 9 2 7 3 13 0 9 2
8 2 13 0 9 1 0 9 2
23 7 6 13 9 1 0 9 2 16 9 6 13 0 1 9 2 7 16 9 13 0 9 2
12 1 0 9 2 16 13 9 2 13 3 9 2
18 10 9 4 13 1 11 11 1 2 11 11 11 11 2 1 0 9 2
16 0 7 0 9 1 11 11 3 4 13 2 1 14 4 13 2
6 2 6 2 1 9 2
4 7 1 9 2
10 9 3 13 1 10 9 2 13 11 2
10 16 9 13 3 9 2 13 1 9 2
11 16 9 13 3 9 2 15 13 1 9 2
6 1 12 9 13 9 2
9 6 13 14 15 9 1 10 9 2
15 2 3 2 13 15 15 2 16 0 9 13 9 1 9 2
9 7 15 3 13 7 1 0 9 2
7 15 4 13 1 12 9 2
7 15 4 13 14 15 13 2
14 13 14 9 14 13 10 9 1 0 11 7 1 11 2
2 3 2
9 7 0 2 10 9 9 13 3 2
8 7 15 4 15 13 3 3 2
10 15 4 13 1 10 9 2 3 13 2
13 7 9 13 2 16 0 9 3 15 13 3 3 2
13 15 13 2 3 0 9 3 13 9 1 0 9 2
17 3 11 14 13 10 9 7 0 9 2 15 9 13 14 15 13 2
7 7 9 6 13 1 9 2
5 15 13 1 9 2
24 3 1 9 2 0 15 1 9 1 9 2 9 1 10 9 13 1 9 1 10 9 1 9 2
27 7 10 2 15 13 2 4 13 3 12 0 9 9 2 15 13 2 11 2 1 9 2 3 11 4 13 2
14 3 2 11 2 14 4 13 1 9 1 9 0 9 2
12 1 9 1 10 9 1 9 15 15 13 0 2
7 1 9 1 0 9 14 2
22 7 10 9 6 4 13 3 10 9 2 16 9 1 9 6 4 13 1 9 1 9 2
4 9 13 9 2
9 9 13 9 2 1 14 15 13 2
9 1 14 13 2 9 13 14 13 2
7 2 15 13 12 0 9 2
4 13 0 9 2
12 2 14 9 6 13 0 2 15 13 0 2 2
18 7 9 2 1 15 13 2 13 2 15 7 14 13 2 9 1 9 2
5 11 6 15 13 2
12 15 13 2 16 13 14 15 13 1 10 9 2
15 10 2 15 13 2 15 13 3 3 1 9 1 0 9 2
18 7 13 15 1 9 2 1 1 10 0 9 7 1 9 1 0 9 2
19 7 15 13 3 9 2 16 13 2 16 1 15 13 9 1 9 7 9 2
28 1 9 2 9 1 9 15 13 1 11 2 3 15 13 15 2 1 1 13 2 16 13 14 15 13 3 3 2
16 3 16 0 13 14 13 1 15 14 10 9 1 9 7 9 2
5 10 9 3 13 2
9 15 15 13 9 2 0 7 0 2
20 1 10 0 9 0 0 9 2 10 7 14 13 10 9 2 13 3 1 9 2
17 14 15 13 14 2 1 10 9 3 4 15 13 14 13 10 9 2
14 1 0 9 9 1 10 9 13 9 14 13 1 9 2
24 7 15 6 14 13 10 0 9 1 0 11 2 3 15 13 10 9 1 9 1 3 0 9 2
8 15 13 3 0 2 11 11 2
11 3 3 12 0 9 3 4 13 1 9 2
13 7 15 15 13 14 13 3 0 2 16 13 9 2
15 15 13 2 16 0 9 1 0 9 4 13 1 0 9 2
15 3 7 15 14 15 13 2 10 0 9 13 0 1 15 2
9 7 11 4 13 1 10 0 9 2
18 7 1 9 2 3 0 9 4 13 9 1 0 9 2 15 13 9 2
3 9 13 2
7 3 13 3 9 1 11 2
7 1 11 7 1 10 9 2
27 7 9 13 2 16 13 9 2 15 14 6 15 13 2 1 9 1 11 7 11 2 15 13 9 1 9 2
13 1 10 0 9 15 13 15 13 7 15 15 13 2
10 9 7 9 4 13 14 13 1 9 2
26 3 3 6 13 14 13 0 9 1 2 11 11 2 7 9 1 2 11 11 2 7 2 11 11 2 2
5 7 15 3 13 2
24 7 3 2 3 7 3 2 14 13 3 2 16 9 2 15 13 1 11 2 13 10 0 9 2
10 7 3 6 13 1 9 1 0 9 2
12 15 13 15 2 15 6 13 14 13 1 15 2
8 3 10 0 9 13 9 15 2
6 3 13 14 15 13 2
20 7 3 13 2 0 9 6 15 13 1 9 1 9 2 7 1 9 1 9 2
8 9 1 11 13 0 1 9 2
9 10 9 6 13 0 1 10 9 2
14 15 3 14 13 2 16 13 3 9 1 10 0 9 2
11 3 13 15 3 3 14 13 1 10 9 2
21 9 2 1 15 13 2 15 13 2 7 15 15 13 0 1 0 9 1 10 9 2
1 9
22 9 15 14 15 13 6 4 13 1 9 15 2 15 15 13 7 13 1 0 15 9 2
8 6 13 14 13 0 0 9 2
22 13 15 2 16 10 9 14 15 13 1 9 1 0 9 1 9 1 9 1 10 9 2
16 2 9 1 9 1 9 2 13 3 14 15 13 1 12 9 2
10 13 15 14 13 9 1 9 7 9 2
12 10 1 10 9 13 9 1 0 9 1 9 2
12 0 9 15 13 1 9 2 0 9 7 9 2
22 14 13 3 14 15 13 1 9 1 9 1 9 2 0 1 0 7 0 1 9 9 2
8 1 0 9 13 0 0 9 2
17 1 0 9 13 9 1 10 9 1 9 1 9 1 9 1 9 2
10 13 9 1 0 9 1 9 7 9 2
19 9 13 1 9 1 9 1 9 1 9 1 9 1 10 0 7 0 9 2
15 10 9 13 1 9 1 9 2 9 7 9 1 9 15 2
24 15 13 1 9 1 9 2 2 9 2 7 9 1 9 2 9 2 9 2 9 7 9 15 2
16 15 13 9 1 0 9 1 9 7 1 9 1 9 1 9 2
16 16 13 9 1 9 1 9 15 2 14 13 9 15 1 9 2
17 14 13 1 10 9 1 9 7 1 9 1 9 1 9 1 9 2
7 0 9 13 9 1 9 2
19 3 9 4 13 1 0 9 7 9 2 3 13 14 13 1 9 7 9 2
12 1 10 9 15 13 14 15 13 14 15 13 2
2 0 9
4 15 13 9 2
18 10 0 9 13 2 16 4 13 15 6 3 13 7 3 3 4 13 2
8 3 3 13 10 14 15 13 2
15 3 13 14 13 1 0 9 7 3 14 13 0 7 0 2
25 13 14 13 1 9 14 13 1 9 1 3 9 2 7 14 13 3 14 15 13 1 9 7 9 2
10 7 1 10 9 3 14 15 13 3 2
11 16 9 13 0 2 15 15 13 10 9 2
15 11 13 2 0 2 7 16 13 0 2 14 13 0 9 2
15 11 13 15 3 2 7 13 9 15 2 16 13 0 9 2
2 0 9
7 10 9 15 13 0 9 2
10 1 9 10 1 12 9 13 0 9 2
19 0 9 1 11 15 13 2 16 4 13 1 9 2 15 13 1 10 9 2
15 11 13 2 16 13 0 9 7 15 13 2 0 9 2 2
10 1 10 9 13 14 13 0 0 9 2
7 13 14 13 10 0 9 2
27 14 14 13 1 9 1 9 1 9 7 14 15 13 9 11 7 9 11 2 7 13 13 14 7 9 11 2
17 1 0 9 1 9 0 9 14 15 13 10 9 1 9 1 9 2
3 9 1 9
29 1 1 15 13 1 0 1 10 9 2 14 13 1 9 14 13 0 9 1 9 2 15 13 14 13 1 9 15 2
5 12 0 9 1 9
26 11 7 11 2 11 2 7 11 2 0 2 13 12 0 9 1 9 2 0 1 9 7 0 1 9 2
16 9 1 9 2 0 1 9 2 13 14 4 13 3 7 3 2
19 3 0 9 1 9 13 0 9 2 9 2 9 1 9 7 9 1 9 2
42 3 3 15 13 9 2 0 15 1 10 9 2 13 3 14 13 1 3 0 9 2 11 2 7 11 2 0 2 11 2 11 2 11 2 11 2 7 11 2 0 2 2
17 1 3 9 3 14 13 0 9 1 9 1 10 12 9 1 9 2
31 3 4 13 1 9 2 13 14 15 13 2 16 13 9 2 0 1 9 2 7 13 0 9 1 9 2 0 1 9 2 2
13 9 1 12 9 9 13 0 9 1 9 1 9 2
10 3 14 15 13 1 0 9 1 9 2
5 9 1 9 1 9
11 1 15 13 3 3 4 13 1 0 9 2
42 0 9 1 9 1 10 9 13 1 10 2 14 13 0 9 2 12 2 12 2 12 2 2 0 9 2 12 2 12 2 12 2 7 9 2 12 2 12 2 12 2 2
16 9 1 9 13 2 16 9 13 0 9 7 9 3 1 9 2
12 9 7 9 6 15 13 1 9 1 0 9 2
9 1 15 15 13 7 3 3 0 2
14 2 0 2 13 0 2 0 7 13 1 0 0 9 2
44 1 0 9 1 9 2 1 15 9 15 13 2 1 0 9 15 13 9 1 10 9 1 12 9 1 9 2 9 2 9 2 0 9 7 9 2 11 2 7 11 2 0 2 2
19 15 13 9 1 0 9 1 9 1 9 2 1 15 9 13 1 15 14 2
26 0 9 1 0 9 15 13 1 9 2 15 15 13 0 2 13 15 14 7 15 13 1 9 7 9 2
23 3 0 9 1 9 13 9 2 9 2 9 7 9 9 14 13 7 14 15 13 1 9 2
25 10 2 15 6 4 13 3 9 15 2 13 3 2 3 7 3 7 13 9 2 16 13 9 15 2
14 2 13 9 15 7 15 13 1 10 2 15 13 2 2
9 2 13 15 7 13 15 9 2 2
12 2 13 15 7 13 1 9 1 0 9 2 2
38 1 9 1 9 1 9 1 9 1 9 7 0 1 9 9 9 13 1 0 9 2 0 9 1 9 13 0 9 1 9 2 3 4 13 1 0 9 2
17 0 9 7 9 15 13 3 0 9 2 3 4 13 1 0 9 2
16 0 9 13 0 1 9 9 2 1 15 15 13 12 7 0 2
18 1 14 15 13 3 1 9 1 9 2 13 3 14 13 0 15 9 2
22 13 3 9 1 9 7 14 13 0 0 9 2 1 14 15 13 10 0 9 1 9 2
51 9 1 10 12 0 9 4 13 1 0 3 9 2 11 2 7 11 2 12 2 0 2 11 2 11 2 11 2 11 2 7 11 2 0 2 11 2 0 2 11 2 7 11 2 0 2 11 2 0 2 2
13 9 1 9 1 0 0 9 15 13 1 0 9 2
10 2 3 15 13 7 15 13 0 2 2
8 2 6 13 1 0 9 2 2
13 2 13 15 1 0 2 3 15 6 15 13 2 2
13 2 3 15 15 13 2 15 13 7 15 13 2 2
10 2 13 15 14 4 13 1 9 2 2
11 2 15 13 0 2 0 7 0 9 2 2
7 2 15 13 3 0 2 2
12 2 13 0 9 1 9 15 1 0 9 2 2
12 9 13 0 0 9 2 14 14 6 13 0 2
37 0 9 15 13 1 0 9 1 9 7 9 2 3 7 1 0 9 2 0 0 9 2 0 0 9 2 9 2 9 2 0 9 7 9 1 9 2
25 16 9 13 3 0 7 0 3 2 13 14 13 1 9 2 0 9 2 9 2 9 7 0 9 2
13 9 1 9 1 0 0 9 15 13 1 0 9 2
7 2 15 13 0 9 2 2
9 2 13 15 9 1 0 9 2 2
11 2 13 1 0 9 1 9 1 9 2 2
7 9 13 3 0 0 9 2
11 15 4 13 1 0 9 2 9 7 9 2
17 16 9 13 3 0 7 0 2 13 14 13 1 9 7 0 9 2
13 9 1 9 1 0 0 9 15 13 1 0 9 2
10 2 13 15 14 13 0 1 15 2 2
7 2 13 15 1 0 2 2
11 2 0 15 13 1 0 7 0 9 2 2
24 9 15 13 1 0 0 9 2 9 1 0 2 0 0 9 2 9 2 9 7 9 1 9 2
15 16 10 9 13 0 2 13 14 15 13 1 9 1 9 2
13 9 1 9 1 0 0 9 15 13 1 0 9 2
12 2 13 0 9 1 10 2 15 15 13 2 2
8 2 15 13 3 0 9 2 2
7 2 13 15 0 9 2 2
20 16 9 13 3 0 7 0 2 13 14 13 1 3 0 9 1 9 1 0 2
15 1 0 9 2 13 14 15 13 14 13 9 15 1 0 2
10 13 15 14 13 0 2 0 7 0 2
15 2 3 13 0 2 14 1 10 2 15 13 15 0 2 2
17 2 6 15 13 7 6 15 13 2 3 9 13 0 1 15 2 2
14 2 3 4 13 1 9 2 3 13 0 7 0 2 2
22 9 1 0 9 1 9 4 15 13 14 13 1 9 7 1 15 14 1 3 0 9 2
9 0 9 1 9 13 12 0 9 2
21 13 15 14 1 0 7 0 2 3 13 2 16 0 13 9 1 0 15 1 15 2
17 13 0 7 0 2 3 1 15 15 13 14 15 13 1 15 14 2
9 13 1 0 1 0 7 0 9 2
25 3 2 15 13 9 1 9 15 14 15 13 1 0 9 2 3 4 13 14 13 1 9 1 0 2
20 3 0 4 13 1 0 9 1 0 7 0 9 1 9 2 11 2 0 2 2
13 0 9 1 9 13 3 0 2 11 2 0 2 2
12 3 15 6 13 2 16 6 13 14 15 13 2
27 12 1 0 15 9 13 14 15 13 14 13 0 15 9 2 3 16 3 14 13 7 13 1 0 0 9 2
14 1 9 1 9 9 1 9 13 3 0 9 1 9 2
22 1 14 15 13 1 9 1 9 2 15 13 7 15 13 2 16 15 3 15 14 13 2
10 1 9 3 9 1 9 6 13 3 2
31 1 16 13 14 13 0 9 2 9 3 13 1 0 9 1 0 9 2 3 6 13 3 9 14 15 2 13 1 9 2 2
14 9 13 0 9 1 9 1 9 2 15 13 0 9 2
31 0 9 1 9 1 9 1 9 13 2 16 15 13 1 0 9 1 0 0 9 2 11 2 11 2 7 11 2 0 2 2
11 1 15 0 13 9 7 1 0 0 9 2
23 3 16 4 3 13 1 9 1 0 9 2 15 6 13 14 13 3 9 1 0 13 0 2
8 15 13 9 1 9 7 9 2
10 13 15 14 13 10 14 15 15 13 2
13 10 9 13 2 1 14 13 0 9 1 0 9 2
12 15 13 2 16 9 13 9 2 1 14 13 2
20 9 15 13 1 9 15 14 15 13 1 9 7 9 2 0 1 9 7 9 2
11 10 9 15 13 1 0 9 1 0 9 2
10 15 6 15 13 1 0 1 9 15 2
13 0 13 0 1 9 15 2 3 4 13 1 9 2
12 15 13 14 13 0 7 0 1 9 1 9 2
13 1 14 13 3 9 2 3 13 14 13 0 9 2
18 13 15 0 9 2 3 16 14 13 14 13 9 1 0 9 1 9 2
26 6 13 9 2 15 13 0 15 9 2 7 15 13 9 2 3 15 13 1 15 2 6 2 13 2 2
23 13 15 3 14 2 15 13 9 2 1 9 2 16 13 9 15 7 15 13 1 0 9 2
6 3 9 13 0 15 14
13 9 1 10 0 9 13 14 15 13 14 15 13 2
9 3 0 0 0 9 4 13 3 2
14 9 1 0 9 1 9 6 13 9 1 0 15 9 2
36 15 13 9 1 0 9 2 13 0 9 2 7 3 13 10 2 15 6 13 1 10 9 2 3 9 2 9 2 0 9 7 9 1 9 15 2
19 9 1 0 9 13 9 2 9 1 9 2 9 1 9 2 9 7 9 2
17 9 3 13 2 16 14 13 3 2 3 15 13 1 10 0 9 2
24 9 13 1 0 9 9 2 3 9 13 0 9 7 9 1 0 9 1 9 1 9 7 9 2
45 10 9 1 9 13 9 2 9 2 9 1 0 9 2 9 1 0 9 1 0 9 2 9 1 0 9 2 0 9 2 9 1 9 1 9 7 9 1 9 1 0 9 1 9 2
23 9 3 13 0 9 2 3 6 4 15 13 3 14 15 13 1 9 2 13 0 9 2 2
13 0 9 13 9 1 0 9 7 9 1 0 9 2
10 7 13 9 2 15 6 13 14 13 2
8 0 9 7 0 9 13 9 2
6 13 14 13 0 9 2
18 10 9 4 13 1 9 1 9 2 11 11 2 2 11 2 0 2 2
28 9 1 0 9 14 15 13 13 9 12 2 12 2 12 2 12 7 12 7 6 13 0 1 9 12 7 12 2
21 0 15 13 3 0 2 0 7 0 13 7 13 0 9 1 9 1 9 1 9 2
50 3 13 14 13 0 7 0 9 2 14 13 1 9 7 14 15 13 1 9 1 9 7 0 9 2 11 2 0 2 11 2 7 11 2 0 2 11 2 7 11 2 0 2 0 11 2 0 11 2 2
20 3 16 6 4 13 14 13 9 7 9 1 9 1 0 9 2 3 13 0 2
21 10 9 2 9 2 9 7 9 3 15 13 7 13 14 15 13 1 3 0 9 2
21 16 13 0 15 9 1 9 7 9 2 13 9 14 13 3 7 0 9 1 0 2
7 10 9 1 0 9 1 9
55 3 0 15 4 13 0 12 9 2 11 2 0 2 2 2 0 2 9 2 9 1 9 7 9 1 0 9 2 2 0 2 9 1 9 2 9 1 0 9 1 9 1 9 2 7 2 0 2 9 2 9 1 0 9 2
19 1 16 13 0 9 1 9 1 9 1 9 2 10 15 13 1 0 9 2
20 0 9 0 15 13 1 0 9 1 9 1 9 1 9 1 9 1 9 15 2
15 0 9 6 13 9 1 9 1 12 2 0 1 9 9 2
8 15 13 9 7 9 1 9 2
11 11 11 2 12 9 2 2 9 2 11 2
12 2 13 2 16 1 12 9 4 15 13 3 2
11 11 11 2 12 9 2 2 9 2 11 2
6 2 1 1 12 9 2
11 11 11 2 12 9 2 2 9 2 11 2
8 2 9 15 3 6 15 13 2
8 7 1 12 9 4 13 3 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
15 0 13 15 3 1 12 9 2 1 14 13 0 15 9 2
12 11 11 2 12 9 2 2 0 9 2 11 2
6 2 15 6 13 9 2
11 11 11 2 12 9 2 2 9 2 11 2
11 2 4 13 3 1 1 12 9 1 9 2
11 11 11 2 12 9 2 2 9 2 11 2
12 2 9 6 13 14 15 13 14 15 13 0 2
15 7 13 13 1 0 9 1 12 9 4 15 13 3 3 2
11 11 11 2 12 9 2 2 9 2 11 2
7 12 1 9 2 11 11 2
19 11 11 7 11 11 13 9 1 0 9 1 9 1 11 11 1 0 9 2
9 11 11 2 9 1 2 11 2 2
7 15 13 0 0 9 1 9
21 2 9 11 2 13 14 15 9 1 3 0 0 9 1 9 1 0 9 1 11 2
17 2 15 3 13 0 0 9 2 0 3 1 9 1 2 11 2 2
24 12 9 13 0 15 9 1 0 9 2 12 9 1 15 14 4 13 1 9 1 9 1 9 2
8 1 15 0 15 9 4 13 2
13 2 1 15 13 9 1 9 1 0 9 1 11 2
14 2 1 9 1 9 2 11 2 7 1 2 11 2 2
23 2 13 14 2 16 2 11 2 14 13 14 13 0 15 0 9 1 9 1 9 1 11 2
11 15 13 0 9 1 3 9 1 10 9 2
21 2 10 9 4 13 12 9 1 0 9 1 11 2 11 2 11 2 11 7 11 2
17 1 9 13 7 1 9 2 15 14 13 0 9 1 9 1 11 2
21 1 9 9 14 13 0 2 16 6 4 13 9 1 9 1 9 2 13 3 15 2
17 11 4 13 1 9 2 9 1 9 2 9 1 9 7 0 9 2
9 12 9 1 0 13 2 16 13 9
18 9 13 14 15 13 1 12 9 3 1 0 9 1 0 9 7 9 2
10 12 9 4 13 1 9 1 12 9 2
12 1 0 9 4 13 1 12 9 1 0 9 2
12 1 0 12 9 4 15 13 1 12 9 3 2
21 12 9 1 0 9 1 15 14 13 1 11 2 16 15 13 9 2 13 3 9 2
28 1 11 9 6 13 14 15 13 1 0 9 1 9 2 3 9 15 13 1 0 9 1 3 1 9 1 11 2
11 15 3 13 0 9 1 0 9 1 11 2
12 1 0 13 3 14 13 0 15 9 1 9 2
24 15 14 15 13 1 0 9 1 11 1 0 9 2 3 14 4 13 7 9 1 9 1 9 2
15 0 9 11 14 13 9 1 9 7 14 13 0 15 9 2
10 1 9 10 9 1 11 13 0 9 2
15 1 9 1 11 1 9 0 11 3 6 4 13 9 15 2
24 0 9 1 0 9 1 0 9 13 9 15 14 15 13 1 9 2 13 9 1 11 11 11 2
3 9 13 9
9 9 13 0 9 2 13 14 13 9
21 9 13 0 9 1 12 9 1 9 1 0 9 2 11 11 2 2 13 1 11 2
6 11 11 13 1 9 2
7 9 13 1 9 1 9 2
8 9 13 1 9 1 9 15 2
11 9 15 13 1 12 9 2 13 1 9 2
5 13 1 9 11 2
15 9 1 15 9 13 14 13 9 1 9 7 13 9 15 2
20 2 11 13 0 1 9 9 2 3 9 6 13 3 2 2 13 9 15 11 2
11 15 7 9 15 11 6 13 14 15 13 2
9 9 13 1 0 9 1 0 9 2
5 13 12 0 9 2
16 1 9 9 3 13 9 2 3 16 9 15 13 14 13 9 2
8 1 10 9 13 3 0 9 2
13 3 11 13 9 1 9 2 1 1 9 15 13 2
8 1 12 0 9 13 1 9 2
18 9 2 15 13 0 2 13 1 9 1 9 2 7 9 6 4 13 2
8 11 13 14 13 9 1 9 2
19 1 0 12 9 12 9 4 13 1 9 2 0 1 9 2 0 1 9 2
5 13 7 0 9 2
15 9 1 9 13 0 9 7 15 13 14 13 7 13 9 2
11 15 13 0 9 1 11 11 11 1 11 2
25 1 9 1 9 3 14 15 13 3 0 9 1 9 2 3 13 1 0 9 2 13 3 0 9 2
26 9 2 16 14 13 9 1 11 11 7 11 11 2 15 13 9 1 9 15 1 0 9 2 13 11 2
12 9 1 9 13 9 1 9 7 6 13 0 2
18 1 12 9 9 13 0 12 9 9 2 13 9 15 1 9 9 11 2
28 1 9 15 13 1 12 9 9 1 0 9 7 1 9 12 9 1 9 1 0 9 1 9 2 13 3 11 2
11 3 15 13 9 1 0 9 1 0 9 2
9 0 9 3 13 14 13 1 9 2
10 9 6 4 13 2 13 9 11 11 2
23 12 9 13 1 11 1 12 9 1 9 1 9 2 13 9 1 0 9 1 9 11 11 2
9 1 15 0 15 13 1 12 9 2
2 11 11
5 13 9 1 0 9
23 14 15 13 9 1 9 1 0 0 9 11 11 7 11 11 2 13 1 9 1 0 9 2
15 15 4 13 1 0 9 1 9 1 9 1 9 12 9 2
13 9 15 13 1 9 1 11 1 9 1 12 9 2
10 1 9 1 9 0 9 14 15 13 2
8 9 13 14 13 11 2 13 9
34 7 9 15 13 1 0 9 3 1 9 1 0 9 2 16 0 9 1 9 13 3 9 1 0 9 2 0 15 1 9 2 13 11 2
10 1 9 1 15 4 13 9 1 9 2
13 1 9 13 11 2 11 2 11 2 9 1 11 2
7 0 9 13 1 2 11 2
19 0 9 13 1 2 11 2 1 9 1 0 9 1 11 2 15 13 3 2
2 11 11
5 0 9 13 0 9
25 0 9 11 11 2 15 13 1 0 9 1 0 9 1 0 9 2 13 0 9 1 11 11 11 2
7 0 9 14 13 9 1 11
12 2 11 2 13 9 1 12 0 0 9 1 9
26 0 9 2 11 2 4 13 1 0 9 1 9 2 15 14 13 3 0 9 1 11 2 15 13 3 2
26 9 4 13 1 12 0 0 9 2 0 1 0 9 1 9 1 9 2 0 1 0 9 2 11 2 2
40 1 9 13 0 9 1 9 2 0 9 2 2 1 9 1 0 9 1 11 1 9 1 0 9 2 0 9 1 11 2 3 7 9 1 9 1 9 1 9 2
15 2 11 2 14 13 1 9 1 9 1 9 7 1 11 2
17 13 15 10 9 14 4 13 1 0 9 1 0 9 1 0 9 2
19 2 11 2 13 0 3 1 9 1 9 1 9 2 9 2 7 9 11 2
6 9 1 11 13 1 9
13 9 1 11 1 11 11 13 14 13 3 1 9 2
24 15 13 3 9 1 11 2 11 11 11 1 9 1 0 9 1 0 0 9 1 9 11 11 2
19 0 9 14 13 0 1 0 9 2 3 4 13 9 1 9 1 0 9 2
6 1 0 9 13 1 9
23 1 15 13 3 14 15 13 7 9 1 0 1 10 9 9 2 16 6 13 9 1 9 2
14 1 0 9 2 3 3 13 7 9 1 2 9 2 2
25 9 13 9 1 0 9 1 0 9 2 15 14 13 10 9 2 16 1 10 9 13 9 1 9 2
3 1 10 9
3 1 12 9
13 3 13 0 9 9 11 14 15 13 1 0 9 2
8 9 2 11 2 2 0 9 2
3 1 0 9
9 9 2 0 9 2 2 0 9 2
3 1 12 9
9 9 2 0 9 2 2 0 9 2
24 1 14 4 13 1 9 1 9 1 11 1 0 9 2 9 13 1 9 1 0 9 1 9 2
21 11 13 9 2 7 9 1 0 15 14 4 13 1 0 9 2 1 3 0 9 2
7 0 9 13 9 1 0 9
7 0 9 13 0 9 1 11
23 15 13 3 0 9 2 11 2 7 9 11 2 16 15 13 1 9 1 0 9 1 9 2
28 1 10 9 0 9 1 2 11 11 2 7 0 15 9 9 4 13 1 12 9 1 0 9 3 1 0 9 2
13 1 12 1 9 9 13 3 9 1 9 1 9 2
9 1 0 9 9 3 13 14 4 13
17 0 9 1 9 4 13 1 15 1 9 2 11 2 2 13 11 2
1 11
6 12 9 9 13 0 9
17 10 0 0 9 7 10 0 0 9 1 11 13 1 9 1 9 2
13 10 9 4 13 1 0 9 1 9 2 11 2 2
15 0 9 13 12 9 1 0 9 7 12 9 1 0 9 2
23 1 9 0 9 1 0 9 13 1 12 9 9 3 2 7 12 9 1 0 0 0 9 2
19 0 9 13 9 1 1 12 9 9 2 1 15 3 12 9 13 3 0 2
1 11
1 11
7 11 13 0 0 9 1 11
18 15 13 0 2 1 1 4 13 9 1 9 1 9 2 0 1 11 2
10 9 4 13 1 9 1 9 11 11 2
33 9 1 9 1 0 9 3 6 13 1 0 9 11 11 2 1 0 0 9 1 9 11 11 7 1 9 1 0 0 9 11 11 2
13 9 13 7 1 0 0 9 1 0 9 11 11 2
1 11
19 1 15 13 12 9 1 11 2 11 2 11 2 11 2 11 7 9 12 2
32 9 1 9 13 7 9 1 0 2 11 11 2 2 2 9 1 11 2 2 2 9 1 9 2 7 2 1 9 1 9 2 2
7 3 10 0 9 13 0 2
12 0 9 13 9 11 7 9 1 0 0 9 2
13 9 14 15 13 1 0 9 1 9 9 11 11 2
18 9 1 0 9 2 0 9 2 14 13 9 1 11 11 7 12 9 2
2 11 11
11 11 11 7 11 11 15 13 1 12 9 9
24 11 11 13 9 1 0 9 2 15 15 13 1 10 0 9 1 11 11 2 0 1 0 9 2
14 15 14 13 0 9 14 15 13 1 12 9 0 9 2
15 0 9 4 13 1 11 11 2 7 9 13 1 11 11 2
11 11 11 15 13 14 15 13 1 12 9 2
7 13 9 1 9 1 0 9
23 9 4 13 1 3 2 7 1 9 1 9 1 11 11 11 1 9 15 13 14 15 13 2
18 1 9 1 0 9 1 9 0 9 11 11 14 4 13 9 1 9 2
29 1 9 1 9 13 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 9 11 11 2
10 1 15 14 13 15 0 12 0 9 2
23 16 15 13 1 15 2 15 14 13 11 11 2 1 15 13 0 9 1 0 9 1 11 2
13 1 0 9 14 13 3 14 14 4 13 10 9 2
22 1 0 3 12 1 0 9 1 2 9 2 1 0 9 14 13 1 0 2 11 2 2
1 11
7 2 11 2 13 0 9 2
17 1 9 14 15 13 9 1 2 11 2 7 9 1 2 11 2 2
2 11 11
36 1 9 1 2 11 2 9 1 9 14 15 13 1 0 9 2 1 14 13 1 0 9 11 11 2 11 11 7 11 11 14 15 13 1 9 2
20 1 0 9 9 1 9 1 9 14 13 9 1 9 1 9 1 9 0 9 2
2 0 9
11 0 11 13 1 0 9 1 11 11 11 2
15 15 13 10 11 1 9 1 9 12 9 1 9 1 11 2
13 10 9 15 13 1 0 9 7 13 0 1 15 2
25 13 15 2 16 13 9 1 0 9 11 11 7 4 13 0 9 1 11 2 11 2 11 7 11 2
5 13 9 15 3 2
23 1 9 1 9 6 13 3 14 13 0 9 1 9 1 9 7 9 1 0 1 0 9 2
28 1 9 1 0 0 9 7 1 9 1 9 14 13 0 0 9 1 9 1 1 12 9 1 9 2 11 2 2
26 3 13 14 15 13 7 0 9 1 9 1 9 1 9 2 1 15 4 13 0 9 7 9 1 9 2
17 9 15 13 1 9 1 9 1 12 9 2 13 9 2 11 2 2
13 3 1 10 9 3 11 13 14 15 13 1 9 2
7 1 15 15 13 7 13 2
14 3 1 9 1 0 9 4 13 12 2 0 2 9 2
5 0 9 1 0 9
9 1 9 1 11 14 13 11 11 2
5 0 9 13 1 11
17 0 9 2 15 4 13 0 9 2 13 0 9 9 2 11 2 2
27 15 13 3 0 7 13 14 4 13 7 1 0 9 2 9 7 0 9 1 9 1 9 2 13 0 9 2
30 3 15 13 9 1 9 7 16 15 13 0 2 9 13 14 4 13 1 0 9 1 0 9 2 16 14 13 0 9 2
1 11
3 13 0 9
24 0 9 2 0 1 9 2 15 13 2 16 15 13 10 9 2 7 15 13 2 16 6 13 2
15 1 9 0 9 15 13 14 13 1 0 9 1 0 9 2
1 11
6 9 13 1 9 1 11
1 11
9 11 15 13 1 12 1 0 9 2
16 12 9 14 13 11 1 9 0 9 2 3 9 14 4 13 2
12 15 13 9 1 0 9 2 0 1 9 3 2
15 0 9 14 15 13 7 13 1 0 9 2 0 9 2 2
21 1 9 1 9 7 11 15 13 14 13 1 9 1 9 1 9 1 0 0 9 2
12 1 9 9 1 9 1 2 9 2 13 9 2
17 15 3 13 9 14 13 1 0 15 9 7 1 15 15 13 11 2
17 7 9 2 7 9 14 13 9 1 0 9 13 0 0 9 3 2
14 9 13 11 11 2 11 11 2 11 11 7 11 11 2
12 1 9 6 13 3 1 0 9 1 0 9 2
7 11 15 13 1 9 1 11
19 2 1 9 13 0 9 1 16 15 13 1 10 9 14 13 3 1 12 2
12 13 2 16 15 13 2 16 15 13 1 9 2
13 13 2 16 13 1 9 1 9 1 0 9 7 9
14 11 11 2 15 13 0 15 9 1 11 2 13 0 2
14 0 13 1 9 2 7 6 13 3 2 3 4 13 2
10 1 15 13 9 15 15 13 1 9 2
9 0 13 14 13 2 3 13 9 2
11 3 13 11 2 13 11 2 11 7 0 2
1 11
16 1 15 10 9 9 15 13 3 3 10 9 2 13 3 11 2
8 9 1 9 13 9 12 1 9
27 9 1 9 1 11 13 1 12 9 3 2 16 13 9 1 9 12 1 9 2 12 9 2 2 13 11 2
30 9 1 9 13 0 1 9 1 0 9 1 0 0 9 2 15 13 2 16 9 1 9 1 11 4 13 1 12 9 2
24 1 15 0 9 1 1 9 12 1 9 13 3 0 7 11 4 13 15 14 13 1 12 9 2
2 11 11
23 6 13 0 9 7 6 13 0 9 2 13 9 11 11 1 0 15 9 1 9 1 11 2
18 1 14 13 1 11 2 11 15 13 7 1 11 2 0 9 7 11 2
7 9 3 4 13 1 9 2
17 9 3 13 9 1 9 2 3 13 9 1 9 2 13 3 11 2
5 0 9 14 13 11
9 9 1 9 15 13 2 16 13 9
16 9 2 15 4 13 9 1 0 0 9 2 13 1 9 3 2
17 15 13 9 1 9 1 9 11 11 14 13 9 9 1 0 9 2
17 15 13 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2
27 9 1 11 7 11 1 9 1 11 4 13 1 0 0 9 11 11 1 12 9 1 9 1 9 1 9 2
17 11 11 15 13 1 9 14 13 9 1 11 1 0 9 7 9 2
13 0 2 1 11 2 13 14 15 13 1 0 9 2
10 1 9 1 11 11 13 9 1 9 2
4 11 13 9 2
21 13 15 2 16 12 9 1 11 2 13 2 1 9 2 3 15 13 1 11 11 2
11 3 1 9 1 11 15 6 13 14 13 2
27 1 9 1 9 11 11 15 13 2 16 12 9 1 9 13 0 9 7 13 14 15 13 15 3 4 13 2
4 13 9 1 11
26 9 3 6 13 14 15 13 2 3 9 1 11 13 1 9 2 3 16 15 13 9 1 9 1 9 2
16 0 9 0 9 13 9 15 1 9 2 16 4 13 0 9 2
9 3 3 0 9 13 9 1 9 2
5 11 15 13 1 9
14 1 9 9 2 0 1 0 9 2 15 13 1 9 2
9 9 13 1 9 7 13 1 9 2
12 12 9 7 9 13 1 0 9 7 0 9 2
10 1 9 4 13 0 9 0 1 9 2
8 3 15 13 9 11 11 3 2
16 3 15 13 2 16 3 10 9 6 4 2 13 2 1 9 2
8 10 9 6 13 0 1 11 2
16 3 7 3 2 14 6 15 4 13 1 9 1 9 1 11 2
11 14 9 13 0 9 7 0 9 1 9 2
2 11 11
8 13 15 9 2 13 14 9 2
11 11 11 2 12 9 2 2 9 2 11 2
10 7 3 9 13 2 14 15 13 3 2
8 3 3 13 1 9 1 15 2
11 11 11 2 12 9 2 2 9 2 11 2
10 2 13 15 3 1 9 1 0 9 2
11 11 11 2 12 9 2 2 9 2 11 2
8 7 16 13 9 2 4 13 2
16 13 2 16 10 9 14 15 13 14 15 13 3 14 13 9 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
3 2 6 2
9 7 16 13 10 9 2 4 13 2
14 16 15 13 3 1 0 9 2 4 13 14 13 3 2
11 11 11 2 12 9 2 2 9 2 11 2
14 2 13 15 2 7 1 9 1 12 9 6 13 3 2
11 11 11 2 12 9 2 2 9 2 11 2
5 2 6 2 13 2
4 2 13 15 2
23 0 9 3 4 13 0 15 9 1 9 2 3 3 14 13 1 9 14 13 9 7 6 2
11 11 11 2 12 9 2 2 9 2 11 2
8 2 1 9 6 13 3 9 2
1 11
5 9 1 9 13 11
13 1 0 9 13 9 2 9 7 0 9 1 9 2
19 15 15 13 1 0 9 1 0 9 1 9 1 0 9 2 0 1 11 2
15 0 9 1 10 9 13 3 1 9 2 13 9 1 9 2
1 11
7 11 13 1 12 9 1 11
17 9 11 11 13 1 9 1 9 11 11 1 12 9 1 9 11 2
22 15 13 0 9 11 11 1 9 1 3 0 9 1 0 9 1 9 1 9 0 9 2
17 0 9 1 11 14 13 0 1 9 7 1 9 2 0 1 9 2
1 11
13 0 9 13 0 9 2 0 9 2 1 0 9 2
8 2 6 13 9 15 11 11 2
20 2 0 13 14 6 15 13 9 1 9 2 15 13 1 9 1 2 11 2 2
10 3 3 1 10 9 1 9 13 0 9
2 0 9
8 2 13 14 15 13 0 9 2
26 9 1 11 7 9 1 11 11 11 13 1 9 1 0 9 1 9 1 9 1 11 2 11 11 2 2
9 1 9 15 13 1 9 1 9 2
3 2 3 2
10 2 11 2 13 9 1 2 11 2 2
14 2 9 1 9 15 13 1 0 9 1 9 1 15 2
7 2 15 14 15 13 9 2
15 2 3 15 13 2 16 1 9 14 13 0 9 1 11 2
13 2 13 14 13 9 2 3 3 15 13 1 9 2
12 2 9 1 11 11 11 13 10 9 1 11 2
13 15 13 14 2 16 14 13 7 0 9 1 11 2
8 2 3 14 13 3 10 9 2
1 11
22 12 9 1 0 9 1 11 1 9 14 13 0 15 0 9 1 9 1 9 7 9 2
1 11
2 13 11
3 13 15 9
51 16 15 13 1 0 9 2 14 13 0 9 1 0 1 15 9 2 3 1 0 9 2 2 3 9 14 13 0 9 2 16 15 13 2 14 6 13 15 14 13 9 7 14 15 13 1 10 7 0 9 2
17 3 15 14 13 0 0 9 7 14 15 13 1 9 7 9 15 2
25 1 9 15 13 1 0 2 0 2 0 7 0 2 1 14 15 13 14 13 0 15 9 1 9 2
42 13 9 15 1 15 2 16 15 13 7 1 0 15 9 1 0 7 0 9 1 9 2 7 1 0 15 9 2 1 14 15 13 14 15 13 1 9 7 0 15 9 2
20 16 15 13 0 2 3 14 15 13 1 0 15 9 7 1 3 0 15 9 2
23 1 9 1 9 6 13 3 14 13 0 9 1 9 1 9 7 9 1 0 1 0 9 2
28 1 9 1 0 0 9 7 1 9 1 9 14 13 0 0 9 1 9 1 1 12 9 1 9 2 11 2 2
26 3 13 14 15 13 7 0 9 1 9 1 9 1 9 2 1 15 4 13 0 9 7 9 1 9 2
16 9 13 0 2 16 0 9 1 9 15 13 3 9 12 9 2
33 9 1 0 4 13 1 0 9 1 0 9 2 16 11 11 2 9 1 11 1 0 15 9 11 2 3 13 12 9 9 1 9 2
10 1 11 11 4 13 1 9 1 11 2
18 0 9 11 11 14 15 13 3 9 1 9 1 11 11 11 2 11 2
15 9 14 15 13 1 9 15 1 0 9 2 0 1 9 2
28 9 1 11 11 2 15 13 7 1 9 1 9 2 13 14 13 9 2 11 11 2 2 13 9 2 9 2 2
14 3 12 9 9 15 13 1 9 15 1 9 7 9 2
6 9 13 12 0 0 9
22 0 9 11 11 2 10 0 9 13 1 0 9 2 13 12 0 0 9 2 13 11 2
18 10 1 9 1 11 13 1 0 9 7 4 13 1 0 9 1 11 2
21 1 10 10 9 15 15 13 1 9 7 13 1 0 9 1 0 9 1 0 9 2
31 9 1 9 1 0 9 1 9 1 0 9 13 2 16 1 9 1 9 9 15 13 3 2 3 16 11 13 9 1 9 2
9 9 15 13 1 9 1 9 1 11
11 0 0 9 3 13 9 15 1 0 9 2
21 15 7 0 9 1 0 9 1 11 11 11 15 13 1 9 1 12 9 1 0 2
17 9 7 9 1 9 1 0 9 1 12 9 13 0 9 1 9 2
8 2 9 2 1 9 1 11 13
16 2 9 2 1 9 1 0 9 11 4 13 1 9 1 9 2
21 15 13 9 9 11 11 2 9 1 0 9 1 9 1 0 9 2 11 2 3 2
13 9 13 9 14 4 13 0 9 1 9 9 11 2
14 1 9 0 9 14 13 9 1 3 0 9 1 9 2
13 9 14 15 13 1 9 7 14 15 13 1 9 2
14 3 0 3 12 9 9 1 9 15 13 1 12 9 2
12 1 9 15 13 1 3 9 12 1 9 12 2
5 9 13 9 1 11
7 13 3 9 1 9 1 9
21 9 1 9 14 15 13 1 0 9 2 1 15 14 13 12 9 2 0 1 9 2
6 13 0 9 1 0 9
22 13 0 9 1 9 1 9 1 0 9 1 0 9 2 9 2 2 13 1 9 3 2
16 9 13 2 16 9 1 10 9 1 0 9 13 0 7 0 2
15 13 9 1 9 1 0 9 2 1 9 7 0 0 9 2
9 9 13 9 1 0 9 0 9 2
12 9 13 0 1 0 9 1 9 2 13 9 2
14 9 12 9 13 1 9 7 9 1 2 0 9 2 2
22 3 14 15 13 9 2 15 14 13 12 9 2 7 1 0 9 14 13 3 12 9 2
12 9 1 9 13 0 9 1 11 1 0 9 2
17 13 15 1 0 9 1 9 14 4 13 0 9 1 11 11 11 2
12 11 13 12 9 9 1 9 15 1 0 9 2
12 1 15 13 3 0 1 9 1 9 2 13 9
25 14 7 1 10 0 0 9 3 3 9 14 13 3 0 1 0 9 1 11 2 15 13 1 9 2
31 0 9 2 11 0 9 11 2 2 11 2 7 2 11 2 2 11 2 13 3 9 1 9 1 9 1 0 9 1 15 2
14 9 1 0 9 14 13 1 11 1 11 1 0 9 2
10 9 1 9 1 9 13 12 9 9 2
1 11
21 1 12 9 15 13 12 9 9 9 1 9 2 11 2 1 9 2 15 13 3 2
26 9 4 13 1 0 9 1 9 2 1 9 7 1 0 9 1 0 9 0 9 3 2 9 7 9 2
35 1 0 9 14 15 13 2 16 4 15 13 0 9 9 9 1 11 2 0 9 2 15 13 9 1 9 1 0 9 7 1 9 1 9 2
11 9 13 1 11 3 12 9 2 13 9 2
22 1 9 15 1 9 3 15 13 3 1 12 9 1 9 2 13 9 1 9 11 11 2
6 0 9 1 9 1 11
6 11 13 9 1 0 9
8 9 13 14 13 9 1 9 2
22 3 0 9 13 9 1 9 1 9 2 1 14 13 14 9 14 13 0 7 1 9 2
8 9 13 1 11 7 15 13 2
22 13 15 9 14 13 1 9 2 13 9 11 1 9 15 1 0 9 1 11 7 11 2
19 1 15 15 13 2 16 9 14 13 1 9 1 11 15 13 1 12 9 2
10 15 13 15 14 4 13 1 0 9 2
13 4 13 7 0 9 2 14 4 13 1 0 9 2
30 11 3 13 14 15 13 14 13 9 1 3 0 0 9 1 9 11 2 11 2 0 9 2 0 9 2 9 1 9 2
20 3 9 1 11 11 11 2 15 6 13 1 9 2 15 13 1 9 1 11 2
14 1 15 1 9 13 3 9 2 1 14 13 0 9 2
15 0 13 9 10 9 14 13 1 9 1 9 2 13 15 2
7 11 15 13 1 9 1 11
25 9 11 14 15 13 9 11 11 2 15 13 9 1 9 1 0 9 1 11 2 13 1 0 9 2
13 9 13 1 9 2 7 11 14 15 13 1 9 2
13 0 9 1 10 0 9 13 0 1 9 1 11 2
13 3 1 0 9 3 13 2 16 13 1 0 9 2
8 11 13 0 9 1 9 11 2
14 15 13 0 1 15 1 9 1 9 7 9 1 15 2
6 9 13 1 0 1 9
17 1 9 9 14 13 14 13 1 9 1 9 15 2 13 3 3 2
15 1 14 13 1 0 1 9 2 9 3 14 13 0 9 2
17 1 0 9 14 13 9 2 15 14 13 0 9 2 16 9 13 2
20 3 1 0 0 9 2 0 11 2 15 13 12 1 0 9 1 9 1 9 2
14 11 11 13 1 9 15 11 1 9 1 0 15 9 2
13 12 9 1 0 9 13 2 16 9 13 0 9 2
13 15 13 9 1 0 9 1 9 2 11 11 2 2
7 1 0 0 9 4 0 2
13 1 15 15 13 0 9 2 0 1 9 7 9 2
5 13 9 1 0 9
22 0 13 2 11 11 2 1 9 1 9 1 11 7 9 1 11 11 11 2 13 11 2
22 9 4 13 1 9 1 9 2 11 11 2 1 11 11 1 9 1 12 9 1 9 2
9 0 9 13 0 0 9 1 9 2
4 9 1 9 12
6 0 9 1 9 15 13
6 9 15 13 1 0 9
12 9 3 13 0 9 1 9 1 9 1 11 2
18 13 15 9 1 10 9 2 13 9 1 9 11 11 1 2 11 2 2
12 3 3 4 13 12 9 9 1 12 9 9 2
23 1 9 13 3 9 11 11 2 9 1 11 9 11 11 2 9 1 9 11 11 7 0 2
19 9 15 13 7 1 0 15 9 2 3 16 1 11 11 9 13 3 3 2
15 1 0 9 4 13 7 12 12 0 9 2 0 1 9 2
9 9 1 9 1 2 11 2 13 0
29 1 12 9 9 7 9 1 1 12 9 13 9 1 9 2 11 2 11 11 7 9 1 2 11 2 11 11 11 2
17 1 9 1 9 1 9 12 13 1 9 1 9 1 1 12 9 2
14 9 1 2 11 2 13 1 0 7 0 9 0 9 2
5 9 6 4 13 2
25 15 13 9 2 1 14 6 15 13 15 1 15 7 1 9 15 2 1 16 3 6 13 1 9 2
10 3 2 3 13 14 13 0 15 9 2
14 2 3 13 2 16 13 1 10 9 2 2 13 0 2
15 15 3 13 15 1 9 1 0 9 2 1 15 13 9 2
12 9 3 1 9 15 13 9 1 9 1 9 2
18 0 1 9 1 9 13 2 16 13 1 9 2 7 3 6 13 15 2
12 1 9 0 3 13 0 9 1 9 1 9 2
6 9 13 9 3 1 9
7 3 15 13 1 0 9 2
11 0 9 1 9 1 0 13 1 3 9 2
11 15 15 13 1 15 2 14 7 1 9 2
22 7 16 6 13 14 15 13 2 9 3 14 13 1 9 1 9 1 14 13 1 9 2
21 1 0 9 1 9 0 0 9 4 13 1 9 1 0 9 7 9 1 0 9 2
21 3 13 2 16 1 0 9 9 1 9 1 9 4 13 1 12 9 1 0 9 2
20 3 1 0 9 7 0 9 10 9 13 12 9 2 7 6 15 13 0 9 2
17 3 0 9 15 13 1 9 2 0 1 0 9 1 3 0 9 2
5 7 13 3 9 2
27 9 1 9 1 0 13 3 9 1 9 7 9 1 0 0 9 2 7 0 9 14 4 13 1 0 9 2
27 9 1 9 1 0 13 3 9 1 9 7 9 1 0 0 9 2 7 0 9 14 4 13 1 0 9 2
23 2 7 9 1 9 1 9 1 9 13 0 1 0 11 2 3 16 11 6 15 4 13 2
14 10 9 1 11 13 3 0 9 1 9 1 0 9 2
11 2 3 3 1 9 14 13 0 0 9 2
6 7 13 1 10 9 2
10 2 3 13 1 9 1 0 0 9 2
9 15 13 0 9 7 1 12 9 2
8 3 1 11 0 9 13 0 2
10 7 6 13 15 3 14 13 10 9 2
9 6 13 10 9 14 15 15 13 2
19 7 7 9 7 9 1 9 6 15 13 1 10 14 9 13 0 7 0 2
3 13 9 2
25 16 15 13 2 14 15 13 9 2 16 15 13 2 14 13 9 2 1 14 6 15 13 1 9 2
16 2 9 15 13 3 0 1 9 1 0 9 7 3 0 9 2
16 3 15 13 14 13 14 15 13 7 1 0 9 14 15 13 2
7 0 9 15 13 1 0 9
14 14 13 9 2 16 9 13 0 1 9 1 0 9 2
18 13 15 3 2 16 1 14 15 13 10 0 9 3 13 9 14 13 2
16 3 13 0 9 3 9 13 0 1 14 15 13 9 1 9 2
16 7 16 1 3 9 9 14 13 9 1 9 1 0 15 9 2
8 13 14 9 14 13 1 9 2
12 11 11 2 12 9 2 2 0 9 2 11 2
16 9 13 0 9 7 13 14 13 1 0 9 1 9 1 9 2
8 7 15 13 3 1 0 9 2
11 11 11 2 12 9 2 2 9 2 11 2
8 13 2 16 3 13 3 3 2
11 11 11 2 12 9 2 2 9 2 11 2
16 2 9 3 13 9 14 13 1 9 2 3 15 13 9 9 2
6 9 3 3 13 0 2
12 11 11 2 12 9 2 2 0 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
15 2 4 13 14 13 2 1 14 13 1 10 9 13 9 2
11 11 11 2 12 9 2 2 9 2 11 2
7 2 6 2 15 13 0 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
17 1 10 9 9 14 13 3 13 3 1 9 7 14 13 10 9 2
15 9 4 13 1 0 9 1 9 2 3 13 9 1 9 2
13 13 15 2 16 9 13 9 1 0 0 9 11 2
19 12 9 1 14 4 13 9 1 11 2 1 10 9 1 11 4 13 9 2
12 13 15 2 16 7 10 9 13 9 1 11 2
6 11 13 0 9 1 11
16 9 1 0 9 1 0 9 13 0 9 11 11 2 13 11 2
16 15 13 9 1 11 2 3 15 13 1 0 15 9 11 11 2
37 0 0 9 15 13 1 9 1 9 1 0 11 1 11 2 7 13 2 16 1 15 13 14 4 13 10 0 9 1 0 9 7 9 1 0 9 2
19 15 13 9 2 15 13 14 15 13 2 1 14 4 13 9 2 13 11 2
6 13 15 0 9 11 11
14 9 11 11 13 3 1 12 9 1 0 9 1 9 2
10 7 1 15 2 9 15 2 13 0 2
20 15 13 1 0 9 2 0 1 11 11 2 11 11 2 11 11 7 11 11 2
8 0 9 13 9 1 9 7 9
22 9 13 1 9 2 0 9 1 9 1 0 9 2 7 9 1 0 9 2 13 11 2
20 9 11 11 14 13 0 1 0 1 9 1 9 9 2 11 1 12 9 2 2
13 1 9 9 1 11 11 14 4 13 0 15 9 2
18 9 14 13 1 0 9 1 9 2 9 7 9 2 1 0 11 11 2
4 13 9 1 9
13 11 11 13 9 1 9 1 2 9 9 2 12 2
11 0 9 13 12 0 9 7 12 0 9 2
24 0 9 1 9 15 4 13 1 0 9 2 1 15 15 13 9 1 0 9 7 0 0 9 2
13 9 4 13 1 0 9 1 9 1 9 1 11 2
27 12 9 13 9 2 13 9 7 9 1 0 9 2 1 14 15 13 1 0 9 1 9 1 9 11 11 2
13 1 0 9 11 11 13 1 0 9 2 11 2 2
6 13 11 7 11 1 9
8 9 15 3 13 12 9 0 2
42 9 1 2 0 2 14 4 13 1 0 9 1 9 1 2 11 2 1 9 1 11 3 1 9 2 0 9 2 2 7 14 13 1 9 3 1 3 0 9 1 11 2
15 9 1 9 1 11 1 0 9 4 13 1 9 1 9 2
32 1 0 9 15 13 2 16 0 2 11 2 4 13 0 9 1 9 11 11 2 16 1 0 9 13 14 15 13 7 1 9 2
16 9 1 2 11 2 14 13 9 1 11 3 1 2 9 2 2
26 11 11 13 3 9 1 9 1 9 1 11 2 7 3 3 15 13 1 9 2 11 2 1 0 9 2
18 9 13 1 0 9 7 6 13 9 2 16 9 15 13 1 12 9 2
6 13 15 1 0 9 2
12 9 13 3 1 9 15 1 9 1 11 11 2
22 0 9 13 1 9 1 0 9 1 2 9 2 2 7 13 7 0 9 1 0 9 2
6 13 15 1 0 9 2
15 13 1 0 7 0 9 2 1 9 1 9 7 1 9 2
12 9 1 9 3 13 3 0 7 13 0 9 2
2 0 9
8 0 9 2 0 11 2 9 11
8 0 11 15 13 1 11 11 2
15 15 13 9 7 9 1 0 11 0 7 1 0 11 11 2
5 11 13 9 1 11
23 11 14 15 13 1 11 11 1 9 1 0 9 2 13 9 1 9 1 9 2 11 2 2
21 0 9 13 2 16 3 6 4 13 9 1 9 2 3 16 7 12 13 3 0 2
16 9 13 9 2 16 9 13 14 15 13 1 9 1 0 9 2
10 0 9 14 15 13 14 13 1 11 2
17 9 13 0 9 2 1 1 13 0 1 9 9 1 11 7 11 2
14 11 15 13 9 15 14 13 1 9 1 9 1 11 2
5 9 13 9 1 9
12 0 9 1 0 9 13 9 2 15 13 9 2
10 1 9 0 9 14 13 1 0 11 2
18 9 13 1 12 9 7 12 9 7 14 13 1 12 9 7 12 9 2
19 9 4 13 1 12 9 7 12 9 7 14 13 1 12 9 7 12 9 2
3 9 1 9
4 9 1 9 2
9 2 13 14 15 4 13 0 9 2
4 2 7 0 2
7 9 1 11 13 9 1 9
24 9 1 0 0 9 14 15 13 1 15 1 0 9 2 13 9 1 9 9 11 11 1 11 2
20 15 15 13 2 3 0 9 1 0 9 1 9 15 13 1 9 1 0 11 2
10 9 13 14 15 13 1 9 1 9 2
5 11 13 14 13 9
8 13 15 1 0 9 1 0 9
19 11 13 14 4 13 3 1 0 0 9 2 13 9 1 0 9 1 11 2
21 9 1 11 4 15 13 1 10 9 1 9 15 1 9 9 2 13 9 1 11 2
17 13 15 1 0 9 9 14 13 9 1 9 15 1 0 0 9 2
17 1 9 13 14 13 1 9 2 13 7 9 11 11 1 9 3 2
3 11 15 13
20 0 9 13 2 16 10 9 0 9 15 13 1 9 1 12 9 2 13 11 2
20 16 13 3 9 1 11 2 3 13 14 13 2 16 9 3 14 14 13 3 2
19 1 15 13 3 9 2 15 13 1 0 9 2 15 6 15 13 1 9 2
16 16 3 12 10 9 15 13 3 2 3 13 1 9 1 9 2
5 11 15 13 9 2
19 9 1 0 9 1 9 1 11 7 0 9 13 9 1 11 2 13 11 2
25 9 13 0 9 1 0 9 7 0 9 1 11 14 13 9 15 1 9 14 15 13 0 0 9 2
15 1 0 9 0 9 13 9 1 0 9 7 13 1 9 2
7 9 3 13 9 1 9 2
12 13 4 9 2 15 4 13 0 9 1 9 2
9 11 13 9 1 9 1 2 11 2
26 0 9 4 13 1 9 2 16 9 1 9 1 0 9 13 3 0 2 7 13 9 1 0 0 9 2
13 13 15 11 7 0 9 14 15 13 9 1 9 2
24 1 12 7 12 9 4 13 3 1 9 1 0 9 1 9 1 0 9 1 11 2 13 11 2
19 1 0 1 9 0 9 15 13 2 16 9 4 13 2 1 0 9 2 2
24 0 9 4 13 9 1 9 2 1 9 1 15 4 13 9 1 9 2 11 7 9 1 9 2
6 11 13 0 9 1 11
27 9 1 0 9 1 11 13 14 13 9 1 0 9 1 11 14 4 13 1 9 1 0 9 1 0 9 2
27 9 13 2 16 0 9 3 14 14 13 14 13 0 9 2 16 6 13 0 9 2 16 9 13 7 0 2
13 15 14 13 2 16 9 13 9 1 9 1 11 2
21 3 13 3 2 16 9 1 11 7 9 1 9 11 11 4 13 0 9 1 9 2
14 11 4 4 13 3 3 1 9 15 1 0 9 11 2
13 0 9 13 9 2 9 7 9 1 9 1 11 2
9 11 11 13 9 1 9 2 11 2
17 15 4 13 1 9 1 9 2 11 11 2 6 3 1 11 11 2
24 15 13 9 11 11 1 9 15 1 9 1 9 1 11 7 15 13 1 0 1 9 12 9 2
11 9 13 1 9 2 11 11 2 1 11 2
11 13 15 2 6 15 13 1 9 1 9 2
7 3 6 4 4 13 1 9
9 13 15 9 1 0 9 1 9 15
9 3 14 13 9 1 9 1 9 2
19 1 2 11 2 15 13 1 9 1 9 1 11 11 1 9 1 0 9 2
12 16 9 1 9 13 2 10 14 13 1 11 2
2 11 11
22 9 1 9 1 9 7 9 15 13 1 9 1 9 7 14 4 13 3 1 0 9 2
13 13 15 1 11 14 13 1 12 2 0 2 9 2
2 11 11
2 0 9
7 3 10 9 13 9 15 2
6 15 13 1 12 9 2
5 0 9 2 9 11
1 9
6 3 1 2 0 9 2
14 9 0 1 0 9 1 9 1 0 9 1 0 9 2
18 9 1 0 9 1 0 9 1 9 1 9 11 7 11 2 9 11 2
6 9 13 9 1 9 15
13 9 15 13 1 9 11 2 3 11 13 1 9 2
21 0 15 13 14 13 9 2 7 15 4 13 2 3 16 1 9 15 13 1 9 2
16 9 13 1 9 7 13 14 13 0 2 16 15 13 1 9 2
7 3 3 0 9 15 13 2
2 11 11
8 11 11 13 14 15 13 1 9
22 0 9 1 9 1 11 11 4 13 2 13 15 1 9 1 0 9 2 13 0 9 2
24 1 0 1 9 7 2 0 9 2 9 12 9 1 9 1 11 14 13 3 0 1 12 9 2
8 11 13 14 13 9 1 10 9
13 13 15 9 1 0 9 1 9 1 0 9 7 9
31 3 14 13 9 1 0 9 2 16 6 13 9 1 0 9 2 9 7 9 2 13 3 0 9 1 11 1 15 11 11 2
20 11 15 13 2 3 1 0 9 13 9 1 11 1 3 0 9 2 13 11 2
14 11 11 13 9 2 1 14 13 9 15 14 15 13 2
6 9 14 15 13 1 0
13 9 15 13 1 9 2 16 13 9 15 1 9 2
8 11 14 13 9 1 9 3 9
7 12 9 4 13 1 0 9
15 1 12 9 4 13 9 1 9 1 9 1 0 0 9 2
11 0 9 13 14 13 1 9 1 0 9 2
21 0 0 9 1 9 1 9 14 4 13 1 0 9 1 9 1 3 0 0 9 2
9 9 13 9 1 0 9 1 9 2
6 9 13 12 9 9 2
24 1 15 12 9 9 13 9 1 9 2 12 9 9 13 0 9 7 12 9 9 13 0 9 2
25 3 2 1 12 9 14 4 13 0 0 9 0 9 2 11 2 2 15 14 13 9 1 0 9 2
29 0 9 1 9 13 11 14 13 9 1 9 1 9 1 9 1 12 9 2 3 13 14 15 13 9 1 0 11 2
32 9 13 2 16 11 7 11 13 14 4 13 14 13 2 16 15 15 13 2 16 15 13 14 13 1 9 15 1 9 1 11 2
8 2 11 2 14 13 9 1 11
13 3 12 0 9 13 14 4 13 1 9 1 9 2
14 9 13 9 1 12 9 1 9 7 0 9 1 9 2
8 13 9 12 9 9 1 0 9
5 15 13 9 3 2
2 13 9
19 9 1 0 9 14 4 13 2 1 9 1 0 9 2 15 14 4 13 2
14 15 13 9 1 11 1 9 1 0 9 1 0 9 2
15 9 14 13 1 9 1 9 1 9 7 1 0 0 9 2
14 1 9 9 13 9 1 9 2 0 9 7 0 9 2
4 0 9 13 9
20 1 9 13 0 9 2 7 9 6 13 14 15 13 1 9 2 15 15 13 2
16 1 15 13 3 9 1 9 1 9 1 11 2 9 11 11 2
15 14 13 14 15 13 9 2 13 3 9 1 11 9 11 2
19 13 15 7 9 9 1 9 14 13 3 12 9 3 2 15 13 12 9 2
7 9 13 14 13 1 9 2
18 9 14 13 9 13 9 1 0 7 0 9 2 0 1 9 1 9 2
5 13 9 1 12 9
16 12 9 4 13 1 9 1 0 9 1 9 3 2 13 11 2
15 9 13 1 9 1 9 1 2 11 11 2 1 12 9 2
7 9 13 9 1 12 9 2
3 0 13 2
7 11 2 3 13 15 9 2
22 3 9 1 10 9 13 9 1 0 0 9 1 0 9 2 0 1 0 9 1 9 2
22 0 0 9 14 13 12 9 2 7 1 9 1 0 9 14 13 3 3 1 12 9 2
33 7 10 9 13 0 9 2 3 15 3 2 13 2 9 1 9 1 0 9 1 12 9 7 9 1 0 9 2 12 9 1 9 2
21 1 10 9 13 3 3 3 9 14 13 1 12 9 1 9 1 0 9 12 9 2
23 7 14 7 1 10 15 9 9 14 13 12 9 1 10 0 9 1 9 1 12 9 9 2
6 3 14 13 10 9 2
24 16 0 9 1 0 9 1 12 9 15 13 1 0 9 1 11 2 9 7 1 9 0 9 2
13 3 13 0 9 2 13 14 4 9 1 0 9 2
19 3 6 2 1 1 1 0 9 0 9 14 13 12 9 9 1 15 14 2
33 7 0 13 9 2 16 3 0 9 1 9 1 0 9 13 14 9 9 2 1 15 14 15 13 9 1 3 0 1 0 15 9 2
10 7 16 15 6 13 14 13 10 9 2
13 3 2 6 4 13 9 10 9 13 9 1 11 2
7 7 16 13 1 0 15 2
7 11 2 3 13 15 9 2
27 9 1 9 13 9 1 9 1 3 12 0 9 2 13 9 2 15 13 3 1 9 1 9 1 0 9 2
9 0 9 13 0 9 1 0 9 2
6 11 13 9 1 0 9
12 9 13 0 9 1 11 14 13 9 1 9 2
15 15 13 11 11 1 9 1 0 9 1 0 9 1 11 2
15 1 9 1 0 9 9 1 9 13 0 1 9 1 9 2
15 0 9 13 0 9 1 0 9 1 0 9 2 13 11 2
10 1 9 9 9 15 13 2 13 15 2
8 6 13 9 1 9 1 9 2
9 1 2 9 2 15 13 0 9 2
8 15 13 9 1 9 11 11 2
24 1 9 9 13 2 16 16 15 13 0 9 2 9 13 14 13 9 2 9 7 9 1 11 2
24 9 11 7 0 9 11 11 14 15 13 3 3 2 1 14 13 9 1 9 1 11 1 11 2
3 9 1 9
8 1 9 9 15 13 1 9 2
10 6 13 14 2 16 9 6 15 13 2
4 16 13 14 2
7 13 15 9 1 12 0 9
9 3 15 14 13 2 14 15 6 13
19 2 11 2 14 13 9 1 9 2 15 6 15 13 9 1 12 0 9 2
16 15 13 0 9 1 9 1 9 2 15 14 15 13 1 9 2
28 9 1 9 14 13 1 9 1 0 9 1 9 7 1 9 1 0 9 2 4 13 1 9 1 9 1 9 2
11 9 15 13 1 0 9 1 9 7 9 2
10 9 1 9 13 7 1 9 1 0 9
7 9 4 13 1 0 9 2
28 11 7 11 2 15 13 9 2 11 2 1 0 9 2 15 13 1 12 9 7 3 15 13 1 9 1 9 2
29 2 11 2 13 0 0 9 1 11 2 15 13 9 1 11 1 9 1 9 12 9 1 9 1 9 1 0 9 2
1 11
4 11 14 13 9
29 2 11 2 13 1 9 1 9 7 9 2 15 14 13 1 0 9 1 11 2 13 3 1 0 9 1 9 3 2
19 13 9 7 1 12 0 9 1 9 1 9 2 15 14 15 13 1 11 2
29 1 9 1 12 9 9 1 0 9 14 15 13 10 9 1 0 9 0 2 3 1 0 9 1 9 2 13 9 2
11 9 1 11 13 9 1 0 1 0 9 2
10 11 11 7 9 1 11 2 0 9 2
11 9 1 9 1 11 13 1 9 1 11 2
20 11 6 15 13 1 0 9 2 3 3 14 15 13 3 1 9 2 13 11 2
19 1 9 7 9 15 13 7 0 0 9 2 1 0 9 11 1 11 11 2
6 11 13 9 1 9 2
8 11 13 14 13 9 1 9 2
11 13 15 9 11 14 15 13 1 0 9 2
19 0 9 13 7 13 0 9 1 9 1 11 1 9 7 0 9 1 9 2
21 1 0 9 1 12 9 11 13 9 14 13 1 11 1 0 9 1 9 1 9 2
11 9 1 14 13 9 9 15 13 1 11 2
13 1 9 1 9 2 0 11 11 2 9 13 3 2
9 0 0 9 13 9 1 0 9 2
25 0 9 13 3 3 0 9 1 9 11 11 13 14 15 13 1 9 1 9 2 7 4 13 3 2
6 9 13 14 13 0 9
33 0 0 9 4 13 9 2 1 14 13 0 9 1 11 11 11 7 9 15 2 13 3 3 0 9 2 11 2 2 0 1 11 2
21 1 9 2 0 9 1 9 15 2 0 9 13 2 16 9 1 9 4 13 3 2
13 9 3 15 13 1 9 15 2 3 3 13 9 2
8 9 1 9 4 13 1 9 2
30 9 11 2 0 9 1 11 9 11 11 7 9 1 11 9 11 11 4 15 13 1 9 1 11 1 15 9 11 11 2
10 13 4 15 1 9 1 9 1 9 2
8 9 1 9 13 2 13 9 2
10 13 15 2 16 15 13 9 11 11 2
12 15 13 0 9 11 11 1 11 9 1 9 2
6 9 13 14 13 0 9
33 0 0 9 4 13 9 2 1 14 13 0 9 1 11 11 11 7 9 15 2 13 3 3 0 9 2 11 2 2 0 1 11 2
21 1 9 2 0 9 1 9 15 2 0 9 13 2 16 9 1 9 4 13 3 2
13 9 3 15 13 1 9 15 2 3 3 13 9 2
20 9 2 11 2 4 13 1 0 9 2 9 15 13 1 0 9 2 13 15 2
7 9 13 9 1 9 1 9
23 12 9 4 13 1 9 7 9 0 9 1 11 7 4 13 1 0 9 1 9 1 9 2
13 9 13 1 9 1 0 9 1 11 1 12 9 2
6 13 9 1 11 11 3
17 0 0 9 13 3 14 14 13 9 1 12 9 9 1 11 11 2
11 3 12 9 13 11 11 7 9 11 11 2
7 11 4 13 1 12 9 2
5 9 14 15 13 2
5 3 14 4 13 2
17 3 13 15 4 3 2 7 14 4 15 13 2 3 6 4 13 2
8 7 15 3 15 13 1 9 2
26 7 14 13 1 9 7 9 2 16 6 13 14 13 1 11 11 7 11 11 2 15 13 14 15 13 2
16 9 1 0 9 3 13 1 9 2 3 9 2 3 9 2 2
20 16 1 9 9 15 13 1 9 2 9 15 3 3 14 15 13 7 13 3 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
9 16 15 15 13 2 15 15 13 2
4 6 13 9 2
14 4 13 14 13 0 2 7 15 3 3 6 15 13 2
7 9 3 13 14 15 13 2
11 11 11 2 12 9 2 2 9 2 11 2
12 6 13 2 16 0 7 0 13 0 1 15 2
11 11 11 2 12 9 2 2 9 2 11 2
5 2 3 13 0 2
5 13 3 0 9 2
5 13 3 0 9 2
8 2 3 3 15 13 0 9 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
16 2 0 9 1 15 3 4 13 1 9 7 13 9 1 9 2
7 1 15 15 13 0 9 2
12 11 11 2 12 9 2 2 0 9 2 11 2
10 2 0 13 9 14 13 0 7 0 2
8 14 1 15 13 3 4 13 2
21 0 9 11 11 4 13 1 9 1 0 9 1 11 2 11 2 2 13 0 9 2
23 1 11 2 15 13 0 9 1 0 9 2 13 3 12 9 1 9 1 0 9 1 11 2
19 1 9 1 9 15 13 2 16 13 9 9 14 13 1 0 9 1 11 2
6 9 13 1 0 9 2
6 9 13 1 9 7 9
22 13 15 0 0 9 1 0 9 7 9 15 1 9 11 11 14 13 7 12 0 9 2
16 9 1 11 4 13 1 9 1 0 9 1 0 3 0 9 2
6 9 13 1 9 1 11
18 3 12 9 13 1 9 7 9 2 0 1 0 9 1 0 9 11 2
9 0 9 4 13 7 0 9 11 2
7 9 1 11 13 1 12 9
28 9 1 9 1 11 1 0 9 11 11 13 1 12 9 2 1 1 1 9 11 2 9 11 2 13 0 9 2
18 1 9 2 3 13 9 1 0 9 2 9 11 11 13 3 12 9 2
29 3 9 1 11 4 13 1 12 9 2 7 1 15 15 13 3 1 12 9 1 9 2 0 1 9 2 13 11 2
10 9 7 9 13 9 1 0 9 1 11
15 13 4 12 9 2 13 9 1 0 9 1 11 11 11 2
11 14 15 13 1 10 0 9 2 13 9 2
12 0 9 1 11 3 14 13 0 9 11 11 2
12 3 1 9 14 13 0 9 1 11 11 11 2
13 1 9 1 0 0 9 14 15 13 0 11 11 2
10 11 11 13 1 2 11 2 1 0 9
15 11 11 13 1 0 9 1 9 2 11 2 1 0 9 2
24 9 15 1 0 9 4 13 9 3 2 1 1 0 9 1 2 11 2 13 11 14 13 9 2
7 11 11 13 2 0 11 2
7 13 0 9 1 2 11 2
15 12 1 9 1 9 2 11 2 14 4 13 1 0 9 2
21 9 13 0 0 9 2 15 14 13 0 1 0 9 2 0 9 2 11 7 11 2
14 9 1 9 13 1 0 0 9 1 2 0 9 2 2
7 11 11 13 9 1 0 9
25 1 9 1 9 2 9 1 0 9 2 11 11 7 11 11 3 14 13 9 1 0 9 2 3 2
16 9 13 1 9 1 2 11 2 1 9 2 0 0 9 2 2
9 2 9 11 2 3 14 13 9 2
9 2 14 2 11 2 13 0 9 2
13 2 6 2 13 2 7 14 13 1 9 1 9 2
17 2 1 9 1 11 11 13 0 9 2 15 13 14 13 1 9 2
7 2 13 7 3 15 13 2
5 3 6 4 13 2
12 2 15 13 14 2 16 9 13 1 0 9 2
12 2 6 4 13 2 7 3 13 14 13 9 2
9 2 13 14 15 1 2 11 2 2
7 13 14 9 1 10 9 2
9 2 13 2 7 6 13 14 13 2
15 1 2 11 2 3 6 4 13 0 7 3 9 13 15 2
7 6 13 3 9 1 15 2
5 2 13 3 9 2
9 3 12 9 2 15 13 0 9 2
6 11 13 9 1 9 11
17 15 13 3 14 13 1 2 11 2 7 15 13 12 0 0 9 2
13 3 11 3 13 3 1 9 1 9 1 0 9 2
6 2 11 2 14 13 2
3 1 9 0
11 9 13 1 9 2 7 13 1 0 9 2
11 1 9 14 15 13 1 9 7 1 9 2
11 3 3 13 1 0 9 7 15 13 0 2
3 0 9 13
6 9 15 13 0 9 2
20 11 13 0 9 1 9 15 1 2 9 2 1 9 1 0 1 0 9 9 2
14 3 3 11 13 1 0 9 2 7 11 13 1 0 2
11 11 15 13 7 1 2 11 2 1 9 2
14 11 1 9 7 11 13 0 12 9 1 2 0 2 2
22 1 9 1 9 13 0 9 1 9 7 1 9 1 0 9 1 0 1 9 1 9 2
6 11 11 13 9 1 11
11 9 1 2 9 7 9 2 13 12 0 9
35 9 2 0 1 9 1 9 15 2 11 2 15 13 3 1 12 1 9 15 2 3 13 7 13 1 9 15 1 2 6 2 10 9 2 2
19 3 1 12 9 13 1 11 14 15 13 1 9 1 0 9 1 9 12 2
12 13 15 15 14 13 9 2 14 16 15 13 2
4 11 14 13 9
1 11
22 1 15 13 9 2 9 2 0 9 7 14 9 2 15 13 14 15 13 1 0 9 2
28 0 0 9 1 9 4 13 1 9 1 11 14 13 9 15 1 9 2 13 9 2 11 11 11 11 11 2 2
6 11 11 13 14 13 0
36 1 9 1 9 9 1 0 15 9 2 9 1 3 2 15 13 2 16 3 6 13 0 9 7 4 13 14 13 9 1 11 11 7 11 11 2
20 13 14 13 0 9 1 9 1 11 7 0 9 2 13 0 9 11 11 3 2
19 1 9 1 9 0 9 13 0 2 0 7 0 9 2 3 7 0 9 2
16 3 1 9 3 15 13 3 12 0 9 1 11 7 0 9 2
12 1 15 7 1 0 9 13 3 9 1 9 2
23 9 13 1 9 1 0 9 2 1 0 9 1 3 0 9 2 3 7 1 9 1 11 2
8 9 13 1 0 9 11 11 2
18 14 11 14 13 9 12 12 1 9 1 11 2 14 13 9 1 9 2
19 12 10 0 9 4 13 9 1 9 1 11 1 0 9 2 15 13 3 2
18 15 13 9 1 9 1 9 1 0 9 2 0 9 2 1 0 9 2
16 9 13 1 9 1 0 9 2 16 13 14 13 1 12 9 2
11 9 7 9 15 3 13 14 13 1 11 2
11 11 11 3 13 9 14 4 13 1 10 9
11 1 12 9 15 13 9 1 11 1 9 2
13 1 10 9 9 9 12 3 13 9 14 4 13 2
16 9 1 9 14 13 9 1 12 9 9 1 9 2 13 11 2
27 14 13 9 3 3 2 3 7 3 14 13 9 15 14 15 13 1 9 1 9 1 0 9 2 13 15 2
17 1 0 9 1 9 4 13 12 9 9 1 9 1 9 7 9 2
10 1 12 9 1 10 9 13 1 9 2
15 0 1 12 9 9 13 1 0 9 7 0 9 1 9 2
8 13 9 1 2 9 1 9 2
18 12 0 9 2 0 1 0 9 2 4 13 1 2 9 1 9 2 2
21 9 14 4 13 1 9 1 11 2 11 2 1 0 9 2 13 9 15 11 11 2
31 0 9 14 13 9 2 15 4 13 1 12 9 2 9 2 9 1 3 2 9 7 9 2 9 7 0 9 2 0 9 2
22 1 9 9 4 13 9 1 11 2 0 9 2 2 11 2 2 2 11 2 7 0 2
12 15 13 2 11 11 2 7 2 9 9 2 2
9 2 11 2 14 13 9 7 1 11
25 0 9 2 11 2 13 0 9 1 9 1 9 1 11 1 9 1 9 1 9 2 15 13 3 2
10 9 14 4 13 1 12 9 0 9 2
29 9 1 0 9 14 4 13 1 0 9 1 9 1 9 2 7 9 14 15 13 3 1 0 9 1 0 0 9 2
10 2 11 2 3 13 10 9 1 11 2
12 1 0 9 9 1 11 14 15 13 1 9 2
5 13 10 9 1 11
13 15 13 9 1 0 15 9 1 9 2 13 9 2
15 13 14 4 13 9 3 1 0 7 1 9 1 12 9 2
16 9 1 9 1 0 9 13 3 9 2 9 7 0 0 9 2
13 11 13 9 1 9 1 9 2 9 7 0 9 2
18 0 9 13 9 1 0 9 7 0 0 9 2 13 0 9 11 11 2
2 9 13
12 13 3 9 1 9 1 9 2 15 13 3 2
16 1 12 9 3 9 1 9 11 13 9 1 0 9 1 11 2
6 11 13 0 9 1 9
21 15 13 9 1 11 1 15 11 11 1 9 1 9 1 9 1 9 1 12 9 2
8 11 15 13 1 9 1 11 11
31 1 9 1 9 11 14 13 0 9 1 0 9 2 11 2 2 1 15 13 7 2 11 2 1 9 1 0 9 11 11 2
12 1 9 15 13 3 12 9 7 12 0 9 2
21 2 11 2 14 13 10 9 1 0 9 2 13 9 1 0 9 1 11 11 11 2
5 9 13 0 9 9
7 9 1 0 9 13 1 3
7 15 15 13 1 0 9 2
15 3 1 0 9 15 13 9 1 12 9 2 13 9 11 2
23 12 9 0 9 14 4 13 1 11 2 12 9 1 15 3 13 1 9 2 13 1 9 2
14 9 1 0 9 14 15 13 1 9 1 9 12 9 2
20 1 0 9 13 0 9 1 9 1 9 1 9 1 0 9 2 13 9 11 2
5 11 13 9 1 11
21 12 9 1 11 2 11 7 9 13 3 9 1 9 1 0 9 1 2 9 2 2
4 9 13 1 9
10 9 13 12 12 9 1 9 1 9 15
15 3 9 13 9 1 0 9 1 9 1 9 1 9 9 2
23 11 11 2 12 9 2 4 13 1 0 9 1 9 1 9 7 3 13 1 9 1 11 2
27 9 13 0 9 1 1 12 9 9 1 12 9 9 1 9 12 1 0 9 2 0 9 2 2 13 11 2
20 1 9 1 9 9 15 11 11 2 1 9 11 2 12 9 2 13 14 13 2
9 9 13 9 1 0 9 1 11 2
13 11 15 13 2 7 9 15 4 13 1 12 9 2
7 0 9 13 3 10 9 2
21 16 0 9 13 11 11 2 1 0 9 1 0 9 13 0 9 1 11 11 11 2
4 11 13 0 9
22 0 9 11 2 0 1 0 9 1 11 11 2 13 0 9 1 9 11 2 13 11 2
34 16 15 13 3 3 0 9 2 1 15 13 2 13 9 14 13 2 16 3 3 13 9 7 13 3 3 9 2 13 9 1 0 9 2
32 1 0 12 9 1 9 4 13 12 9 1 11 2 7 9 2 3 1 0 0 9 2 13 14 13 1 0 9 2 13 11 2
3 13 11 11
12 0 9 9 11 11 13 1 11 1 0 9 2
18 11 11 13 1 11 1 0 9 0 9 1 9 1 9 2 11 2 2
1 9
5 11 11 13 0 9
12 2 11 2 13 2 12 0 9 2 1 0 9
24 1 9 1 1 9 9 15 13 1 9 2 7 14 9 13 0 9 2 0 1 0 0 9 2
17 10 2 15 13 2 3 2 1 2 11 2 2 15 13 11 11 2
12 0 13 14 13 10 9 2 3 13 14 13 2
19 15 13 0 0 9 11 2 15 13 9 1 0 9 1 2 0 2 11 2
12 3 14 10 9 1 9 14 13 1 0 9 2
33 11 11 2 3 1 0 9 2 7 9 11 11 13 0 2 16 13 3 12 9 2 1 14 13 9 1 0 9 1 9 1 15 2
9 7 1 12 9 9 13 0 9 2
11 1 0 9 11 7 11 13 1 0 9 2
8 0 9 13 9 7 9 1 9
14 9 1 11 3 13 14 15 13 9 1 0 1 9 2
27 9 13 1 0 9 2 3 16 3 9 3 6 13 1 0 9 2 1 9 2 7 13 0 9 7 9 2
4 13 9 1 11
26 9 13 9 2 11 2 1 0 0 9 11 1 9 15 1 9 2 11 2 13 9 2 11 11 2 2
5 11 11 13 0 9
27 9 1 2 9 11 12 2 13 1 9 2 11 2 2 3 15 13 9 1 0 9 1 9 2 9 2 2
27 9 15 13 2 16 9 1 9 3 13 0 2 1 15 15 6 13 14 13 7 2 9 1 9 12 2 2
18 9 1 3 1 9 13 1 9 2 9 12 2 1 9 2 11 2 2
34 9 1 9 1 0 9 1 12 9 11 11 7 9 11 11 2 2 9 12 2 2 15 13 1 9 1 9 1 11 11 2 11 2 2
6 9 9 1 9 1 9
20 9 0 0 9 4 13 1 9 1 9 1 11 11 11 2 13 1 0 9 2
14 9 4 13 1 9 2 16 13 0 1 9 0 9 2
4 11 13 1 11
20 9 9 9 13 11 11 1 0 9 1 11 11 2 7 15 6 13 9 15 2
11 15 13 0 1 9 2 0 1 11 1 11
9 15 15 13 14 13 1 0 9 2
9 9 1 11 13 0 9 1 9 2
22 15 6 13 0 9 2 3 15 13 1 9 7 13 1 0 9 1 11 2 13 9 2
1 9
9 13 0 9 1 9 1 0 9 2
31 1 0 9 0 9 11 14 13 0 9 1 9 1 11 7 11 2 13 9 1 0 9 1 0 9 2 0 1 0 9 2
21 0 9 13 10 9 1 9 1 10 9 1 0 9 7 9 1 9 1 10 9 2
6 11 13 9 1 11 11
14 9 1 9 13 0 9 1 2 0 0 11 7 11 2
19 11 13 2 16 3 4 13 0 9 1 11 2 7 13 14 13 9 15 2
11 1 0 13 9 1 9 1 9 11 11 2
27 9 1 9 1 11 13 9 1 9 11 11 1 9 1 9 2 11 2 1 2 0 0 11 7 11 2 2
20 1 15 1 9 1 9 1 9 1 0 9 9 4 13 3 0 1 12 9 2
11 9 11 13 3 2 13 1 9 1 9 2
27 9 1 9 13 3 9 2 15 13 0 9 1 9 1 10 9 2 13 1 9 2 0 9 2 1 9 2
20 12 9 1 11 4 13 9 1 9 1 9 1 9 1 9 2 13 11 3 2
13 15 3 13 1 3 0 9 1 9 1 0 9 2
7 10 9 15 13 1 3 2
12 0 9 1 10 9 4 13 3 3 0 9 2
13 1 9 13 2 16 13 14 13 9 1 10 9 2
19 10 9 13 3 1 0 9 7 13 7 1 0 9 2 7 1 0 9 2
7 9 15 13 14 13 0 9
10 11 13 1 9 1 9 1 0 9 2
20 15 13 0 1 9 1 9 11 11 7 9 1 0 15 9 9 9 11 11 2
11 11 13 0 9 1 9 1 9 7 11 2
24 9 1 9 1 9 1 9 1 11 7 11 2 0 9 2 6 4 13 1 15 2 13 11 2
22 3 15 13 9 1 0 9 2 13 14 15 13 9 1 9 1 9 2 13 3 9 2
18 13 9 1 9 1 0 9 7 0 11 2 13 11 7 13 3 9 2
17 3 6 4 13 9 1 9 1 9 1 0 9 2 13 9 11 2
9 3 9 15 13 1 9 12 9 2
12 1 3 9 1 11 3 1 9 13 0 9 2
13 0 9 14 13 1 9 1 0 9 2 13 9 2
10 0 9 13 0 9 7 13 0 9 2
6 13 3 1 0 9 2
6 11 13 9 2 13 9
21 0 9 1 9 1 9 13 9 11 11 2 13 12 9 1 9 1 9 1 11 2
19 1 11 15 13 0 9 11 11 1 12 9 7 9 11 11 1 12 9 2
8 9 15 13 1 9 1 9 15
15 1 9 1 0 9 3 9 13 2 16 6 13 1 9 2
14 1 9 13 9 1 0 9 7 0 9 1 0 9 2
13 9 15 13 3 9 1 0 15 9 2 13 11 2
16 0 9 4 13 7 1 11 11 1 0 15 9 1 0 9 2
19 3 13 0 9 14 15 13 1 9 2 13 15 3 9 1 11 11 11 2
13 15 15 13 1 0 9 1 0 9 2 13 11 2
18 3 11 7 9 11 13 2 16 4 13 2 7 0 9 6 13 15 2
16 0 9 15 13 9 2 1 15 15 13 9 1 9 12 12 2
20 1 0 9 9 3 6 4 13 1 9 2 16 13 1 9 1 9 1 11 2
6 9 11 13 9 1 9
15 1 13 9 4 13 1 9 1 9 1 2 0 9 2 2
15 0 9 9 11 14 15 13 1 9 1 0 9 1 9 2
4 9 13 1 11
24 0 9 4 13 1 9 1 11 1 9 1 0 9 1 9 1 9 1 12 0 9 1 11 2
18 1 0 9 1 0 9 11 13 9 14 13 9 7 1 0 0 9 2
11 9 13 1 9 1 9 2 11 11 2 2
11 1 9 15 13 7 0 3 2 11 2 2
34 9 14 6 15 13 2 13 2 13 2 14 6 13 2 16 6 4 13 3 1 0 9 1 9 1 11 2 3 14 15 13 0 9 2
19 15 13 9 11 11 1 9 2 16 0 15 9 4 13 1 9 1 9 2
7 9 13 14 15 13 9 2
11 15 13 9 1 0 2 0 2 0 9 2
2 13 2
8 1 12 9 9 3 13 9 2
31 13 3 10 0 9 2 3 3 3 15 14 15 13 14 13 9 15 2 1 14 13 1 10 14 13 1 9 1 0 9 2
11 11 11 2 12 9 2 2 9 2 11 2
11 2 13 15 14 15 13 1 9 1 15 2
10 15 13 14 13 10 9 1 10 9 2
11 11 11 2 12 9 2 2 9 2 11 2
10 2 3 4 15 13 2 3 13 2 2
11 11 11 2 12 9 2 2 9 2 11 2
6 6 13 9 14 13 2
10 13 13 15 14 13 1 9 1 9 2
11 11 11 2 12 9 2 2 9 2 11 2
4 2 3 10 2
6 6 15 13 1 9 2
5 13 7 0 9 2
11 11 11 2 12 9 2 2 9 2 11 2
7 2 14 15 13 3 9 2
11 11 11 2 12 9 2 2 9 2 11 2
5 2 6 13 15 2
11 11 11 2 12 9 2 2 9 2 11 2
8 2 13 15 14 15 13 3 2
10 1 9 3 13 14 15 13 1 9 2
11 11 11 2 12 9 2 2 9 2 11 2
2 11 13
7 9 13 1 0 9 1 9
17 14 13 1 9 1 9 1 0 9 2 16 9 13 1 12 9 2
11 3 9 14 13 1 9 1 9 0 9 2
19 11 2 10 0 9 3 4 13 3 2 14 4 13 1 0 9 1 9 2
19 9 1 0 15 9 14 4 13 2 3 9 13 9 2 0 15 1 9 2
20 3 1 15 13 0 9 2 13 9 11 11 2 15 13 1 0 9 3 3 2
17 0 9 13 1 9 7 3 1 0 9 11 11 7 9 11 11 2
16 11 15 13 1 9 2 3 11 11 7 11 11 15 13 9 2
10 11 14 15 13 1 9 1 11 11 2
7 9 13 14 13 9 1 11
12 12 9 1 9 1 0 9 4 15 13 9 2
18 1 9 7 9 0 9 1 11 11 13 3 1 10 1 9 1 11 2
15 9 13 9 1 11 2 13 3 0 9 1 11 11 11 2
17 11 11 15 13 1 9 1 0 1 0 9 2 13 2 11 2 2
15 1 9 11 13 9 1 0 15 9 11 11 7 11 11 2
11 0 9 14 13 1 9 1 9 11 11 2
12 15 13 3 9 1 9 2 3 13 1 11 2
16 0 9 1 0 9 3 6 15 13 7 15 15 13 1 11 2
11 1 10 9 1 10 9 13 14 13 9 2
5 14 0 13 3 2
19 1 9 9 14 13 1 9 1 9 1 9 1 9 1 9 2 11 2 2
12 1 12 9 9 15 13 9 1 0 9 1 9
9 0 3 13 14 13 9 1 9 2
5 14 14 13 0 2
8 11 11 13 9 1 2 11 2
18 0 9 11 11 13 0 9 1 9 1 9 1 9 12 2 11 2 2
4 0 9 9 2
17 11 11 4 13 1 9 2 16 3 15 13 9 1 9 1 11 2
18 1 0 9 9 1 9 13 9 1 9 7 1 1 9 13 3 0 2
7 9 13 11 11 7 11 11
18 9 1 11 11 3 15 13 2 1 16 9 1 9 13 1 12 9 2
31 16 9 15 13 2 1 0 9 14 13 12 9 9 1 9 7 3 12 0 1 9 1 11 2 13 9 2 11 11 2 2
7 9 1 9 15 13 11 11
12 9 1 9 15 13 11 11 1 0 15 9 2
19 1 15 3 9 1 9 15 15 13 3 0 7 15 6 13 14 13 9 2
3 9 1 9
6 9 15 13 1 9 2
13 13 9 2 13 9 2 13 0 9 2 13 9 2
9 2 13 2 16 13 9 14 13 2
6 2 10 9 2 14 2
6 16 13 2 14 13 2
6 6 13 0 9 3 2
10 0 9 13 9 1 9 1 0 9 2
10 1 9 13 0 9 1 10 1 9 2
21 1 9 1 0 9 13 3 3 2 16 3 1 0 9 13 9 7 13 0 9 2
4 1 9 13 9
13 9 15 13 1 9 1 0 9 2 13 1 11 2
5 11 11 13 1 9
20 11 11 4 13 1 9 2 7 11 11 4 13 14 13 3 1 0 0 9 2
9 15 13 7 9 2 15 13 9 2
14 0 9 1 0 9 9 15 13 1 9 2 13 11 2
10 9 15 4 13 1 9 1 0 9 2
9 13 15 2 16 9 13 1 9 2
8 2 3 13 2 13 9 1 11
13 3 1 0 9 9 15 13 9 14 13 0 9 2
19 15 13 1 0 0 9 1 9 11 11 7 9 11 11 2 13 1 0 2
7 9 13 1 9 1 9 2
7 3 9 3 6 13 15 2
6 1 15 13 0 9 2
13 1 9 3 0 13 2 16 4 13 9 1 11 2
13 1 9 9 13 0 2 11 11 4 13 1 9 2
16 1 9 13 3 2 16 0 9 14 13 0 9 1 0 9 2
13 3 9 14 13 0 9 1 0 15 7 1 9 2
3 9 1 9
13 9 13 0 1 9 7 1 9 1 10 9 9 2
3 9 1 9
4 2 7 15 2
4 2 3 15 2
9 15 3 9 13 2 15 9 13 2
5 9 15 13 1 9
21 2 2 9 11 2 15 13 3 1 0 9 1 9 11 2 9 0 9 1 9 2
8 9 13 1 9 2 13 11 2
20 0 11 11 1 9 11 13 9 2 3 13 1 0 1 9 9 2 13 9 2
13 9 15 13 1 9 7 9 15 15 13 1 9 2
8 9 1 11 14 13 9 1 11
11 11 7 11 13 0 9 1 0 1 9 9
17 15 13 3 1 9 2 11 2 2 0 1 9 1 9 1 9 2
9 9 13 1 9 1 9 12 9 2
14 0 0 9 1 9 4 13 1 9 3 1 0 9 2
10 0 9 4 13 3 1 11 1 9 2
16 7 10 9 3 9 4 13 1 0 0 9 1 9 7 9 2
17 1 11 14 1 0 9 13 14 15 13 15 14 13 9 1 9 2
14 9 1 9 15 13 1 9 2 0 1 0 0 9 2
34 1 15 13 3 2 16 12 0 0 9 2 9 7 9 2 13 14 15 13 9 1 9 1 10 9 1 12 9 1 0 1 15 9 2
11 1 9 13 2 16 3 13 9 1 9 2
17 9 4 13 1 11 11 2 9 0 9 1 0 9 1 0 9 2
7 11 13 11 1 0 1 9
7 11 15 13 1 0 9 2
15 3 13 0 9 1 12 2 16 11 14 13 1 0 9 2
13 1 0 10 9 7 9 15 14 15 13 1 9 2
25 0 9 1 9 13 3 0 2 7 7 13 2 16 1 11 13 10 9 2 15 6 15 13 1 15
5 13 9 7 9 2
5 2 0 13 11 2
19 3 9 2 0 2 14 15 13 1 9 2 1 15 13 1 9 1 11 2
5 0 9 13 1 9
29 0 2 0 2 0 7 0 9 1 9 4 13 1 2 0 2 9 1 9 2 1 15 9 13 9 1 0 9 2
10 9 7 9 13 0 9 7 13 9 2
17 1 10 9 9 2 11 2 13 0 15 9 2 0 1 0 9 2
22 9 15 13 1 9 15 2 15 13 1 0 9 1 11 7 14 13 3 1 0 9 2
9 9 13 1 12 9 1 9 3 2
8 9 13 0 9 1 12 9 2
12 12 9 0 9 1 9 13 0 9 1 3 2
14 0 9 14 13 3 1 9 1 9 2 13 3 9 2
4 11 13 1 11
17 15 13 9 1 11 11 11 1 9 9 2 11 2 1 11 11 2
17 3 11 13 9 1 9 7 9 2 0 1 15 2 13 1 11 2
24 3 14 13 3 14 15 13 3 0 9 13 14 13 1 0 9 1 0 9 1 3 10 9 2
11 9 1 10 9 14 13 3 0 1 15 2
7 11 13 9 1 9 1 11
9 11 13 9 1 0 9 1 11 2
20 9 1 11 11 13 1 0 9 0 9 2 7 15 4 13 3 14 15 13 2
11 0 0 9 1 11 11 11 13 1 9 2
12 0 9 1 9 1 9 13 0 9 0 9 2
3 9 1 9
3 2 15 2
23 2 14 3 9 15 15 13 14 13 1 9 2 7 15 15 13 9 2 1 14 13 3 2
7 13 9 1 0 9 1 11
15 9 1 0 9 1 11 14 13 1 9 1 9 1 9 2
15 9 3 3 14 13 2 16 15 13 0 9 1 0 9 2
13 15 13 3 9 1 9 1 9 1 9 11 11 2
11 9 15 3 13 9 1 0 9 1 11 2
15 0 9 1 9 1 15 13 1 12 9 2 13 3 11 2
21 2 11 12 2 13 0 0 9 1 9 2 15 14 4 13 1 9 1 0 9 2
2 11 11
12 9 11 7 9 11 11 13 3 0 1 9 2
20 15 13 9 1 0 9 1 2 11 11 2 2 0 1 9 1 9 1 11 2
12 12 13 0 7 0 9 1 9 1 0 9 2
11 1 15 13 11 11 2 11 7 11 11 2
4 13 9 1 11
6 11 14 13 1 0 9
11 0 9 14 4 13 7 1 11 7 11 2
24 9 1 11 14 15 13 1 9 1 9 1 0 9 9 2 1 14 6 15 13 1 0 9 2
9 9 1 2 0 9 2 13 1 9
12 0 11 11 4 13 1 9 1 0 15 9 2
26 1 9 1 0 4 13 3 12 9 2 9 12 7 9 1 0 9 1 0 9 9 1 0 9 12 2
7 11 11 15 13 1 11 11
17 9 1 11 11 6 13 3 14 13 9 15 7 13 9 1 11 2
28 1 9 1 0 9 11 13 14 15 13 1 9 15 1 9 1 9 1 9 2 13 7 0 2 11 11 2 2
11 9 1 0 9 4 13 1 9 1 9 2
15 3 9 4 13 1 0 9 2 14 4 13 3 12 9 2
3 9 13 11
15 0 9 15 13 1 0 9 1 9 1 11 1 0 9 2
7 9 7 9 13 9 1 11
22 15 14 13 0 9 1 0 9 2 9 1 9 2 9 1 9 2 2 0 1 11 2
25 12 9 4 13 9 1 12 9 9 1 9 1 9 1 9 7 13 14 13 9 1 9 1 9 2
12 1 9 15 15 4 13 7 0 9 11 11 2
6 9 11 11 15 13 2
6 9 3 13 3 9 2
24 11 11 2 11 11 2 11 11 7 11 11 7 11 11 13 9 2 15 9 13 1 0 9 2
12 0 1 15 9 3 14 13 1 9 1 11 2
10 11 13 1 0 1 9 1 9 1 11
40 0 9 1 9 1 11 11 7 11 11 1 0 9 1 0 9 1 9 1 9 7 9 1 11 2 11 2 1 0 9 9 12 9 13 1 9 1 0 9 2
13 11 13 1 0 9 7 13 0 9 1 0 9 2
12 11 14 13 9 12 12 1 0 9 1 9 2
7 13 9 1 2 0 9 2
31 1 9 1 0 9 4 13 9 1 9 1 0 9 2 9 7 0 9 1 11 2 11 2 11 7 11 2 15 13 3 2
14 9 13 1 0 1 11 9 1 9 2 0 9 2 2
15 3 1 15 13 0 9 1 9 1 10 9 2 13 9 2
6 0 9 13 9 1 9
11 14 4 13 7 0 9 1 9 1 9 2
11 0 9 1 9 14 13 9 1 12 9 2
32 16 3 9 13 14 13 9 15 1 0 9 1 0 9 2 9 14 4 13 1 9 2 15 14 13 10 9 2 13 1 9 2
26 9 7 0 9 14 15 13 7 13 1 9 1 9 1 9 2 15 15 13 3 1 9 1 0 9 2
54 9 1 9 7 9 11 11 14 13 9 1 0 0 9 2 1 15 13 9 15 0 9 2 0 11 11 2 2 9 2 11 2 2 2 11 2 2 2 11 2 2 2 11 2 2 2 11 2 2 2 0 9 2 2
15 14 15 13 7 9 1 9 7 9 1 9 1 0 9 2
22 1 9 1 0 9 14 13 9 1 9 9 1 0 0 9 2 9 1 9 11 11 2
4 9 13 1 11
17 3 3 10 13 1 11 7 1 9 13 9 14 15 13 1 9 2
11 11 13 12 3 0 9 1 1 12 9 2
22 13 14 13 1 9 1 9 2 7 3 1 12 9 13 0 15 1 10 9 11 11 2
38 0 9 13 0 9 1 9 1 0 9 2 9 7 0 9 1 0 7 0 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
18 9 15 13 1 0 9 1 9 2 0 9 2 1 10 9 1 11 2
28 3 1 11 13 0 9 1 0 9 1 9 2 15 13 14 15 13 7 1 9 2 16 13 9 1 0 9 2
11 9 13 3 1 12 9 1 3 1 9 2
17 9 13 2 16 2 11 2 13 9 1 9 1 3 1 12 9 2
27 9 1 9 1 9 13 9 1 9 1 0 9 2 3 7 0 9 1 9 1 9 2 13 1 0 9 2
5 13 9 7 1 9
23 1 10 9 9 13 14 15 13 9 7 1 9 2 13 1 2 11 2 2 11 2 3 2
7 9 13 12 9 9 1 9
13 15 13 9 11 1 9 1 0 9 1 11 3 2
13 3 9 1 9 15 1 9 13 1 9 12 9 2
10 1 15 9 13 1 9 1 0 9 2
17 10 0 9 1 9 14 15 13 1 12 9 9 2 13 9 3 2
10 9 13 9 1 9 1 0 0 9 2
38 0 9 13 2 16 9 14 13 9 1 9 2 15 13 1 9 2 9 2 9 7 3 2 13 11 11 2 9 1 9 2 0 9 2 1 0 9 2
22 1 9 1 9 9 1 9 13 2 7 1 0 9 9 6 4 13 2 13 0 9 2
19 11 11 4 13 1 9 1 0 9 2 11 11 2 2 0 3 1 9 2
19 7 9 1 9 1 11 2 11 11 2 15 13 1 10 9 7 15 13 2
10 3 6 13 3 14 9 14 13 0 2
5 9 13 9 1 11
22 9 11 11 7 9 11 11 13 9 1 9 1 0 9 1 9 11 2 13 3 3 2
15 9 13 1 9 1 11 11 7 0 1 0 1 11 9 2
7 9 13 1 9 12 9 2
12 13 15 9 14 13 1 9 7 1 0 9 2
18 1 15 3 9 1 11 13 14 13 0 9 1 0 0 9 1 9 2
15 7 14 3 1 9 9 1 15 3 15 13 1 0 9 2
6 9 1 15 13 3 2
7 1 10 9 2 13 9 2
20 1 0 3 2 0 9 13 7 0 0 9 11 11 2 3 7 0 10 9 2
22 1 9 1 9 15 13 10 0 9 1 9 1 9 2 7 1 9 6 15 13 15 2
8 9 12 9 13 11 1 0 9
31 12 7 12 9 9 13 9 1 11 1 10 9 1 0 9 7 9 1 9 2 13 9 11 2 16 15 13 1 0 9 2
32 0 9 1 9 11 1 0 9 11 11 11 13 9 1 9 1 9 1 9 11 11 1 0 0 9 1 0 9 1 12 9 2
16 1 11 9 1 11 6 4 13 14 13 0 9 2 13 9 2
23 10 9 13 0 9 1 11 2 15 15 13 0 9 14 15 13 14 13 9 15 11 11 2
8 9 13 1 11 1 12 9 2
13 15 13 3 1 10 0 9 1 9 2 11 2 2
5 9 13 1 0 11
21 0 9 4 4 13 3 1 9 1 0 11 2 13 0 9 1 0 9 1 11 2
4 0 9 13 9
8 1 9 13 0 9 11 11 2
21 9 13 7 9 1 9 2 0 9 2 2 15 14 15 13 1 0 9 1 11 2
11 1 9 1 11 11 9 4 13 11 11 2
13 2 11 2 2 11 2 13 9 12 12 1 11 11
25 9 14 13 1 11 1 9 1 9 2 16 1 0 9 14 15 13 1 0 9 1 2 11 2 2
13 9 1 11 1 11 13 1 9 2 13 3 3 2
14 2 9 2 13 0 9 1 9 1 9 1 0 9 2
15 1 9 1 11 15 13 7 14 14 13 1 11 1 9 2
8 13 11 7 11 14 15 13 9
9 9 13 9 1 0 7 9 1 9
26 0 9 11 7 11 2 3 7 0 9 1 0 9 4 13 14 13 9 15 2 13 2 11 11 2 2
13 0 9 1 0 9 1 0 9 13 1 0 9 2
20 0 9 11 11 13 0 9 1 9 1 0 9 2 1 10 9 15 13 9 2
6 13 9 1 9 1 11
24 0 9 1 11 13 3 1 9 1 0 9 1 0 9 7 0 9 1 9 2 13 0 9 2
26 9 4 13 1 9 2 7 1 3 13 1 9 7 9 1 9 2 16 1 15 9 13 0 1 9 2
14 9 13 14 13 9 1 0 1 0 9 7 0 9 2
6 13 9 1 11 1 9
26 9 1 9 1 11 14 4 13 1 1 12 9 2 16 13 3 9 2 13 3 9 11 11 1 11 2
10 15 13 0 9 1 0 9 1 9 2
13 1 0 9 14 13 3 0 9 2 13 9 11 2
24 15 13 9 1 9 2 11 11 2 2 2 11 11 2 2 2 11 11 2 7 2 11 2 2
2 11 11
29 1 9 1 9 1 10 9 1 0 11 7 11 13 9 2 15 13 0 9 2 13 9 1 9 1 11 11 11 2
9 13 9 14 15 13 2 13 11 2
7 11 13 14 13 10 9 2
2 11 11
3 9 1 9
7 0 9 1 0 0 9 2
7 9 11 13 1 0 9 2
5 2 6 2 9 2
6 2 6 2 9 11 2
14 15 13 3 11 11 2 9 1 9 1 9 1 11 2
16 3 9 1 9 13 1 12 9 1 0 15 9 2 13 9 2
13 1 12 9 9 13 9 1 9 1 9 1 9 2
35 11 13 3 1 12 9 9 3 1 9 1 9 7 9 2 3 7 1 9 1 9 1 12 9 1 0 9 1 9 1 12 9 1 9 2
7 1 11 13 12 12 9 2
6 12 9 1 9 1 9
13 3 9 6 15 13 1 9 1 12 9 1 9 2
15 3 3 1 9 1 12 9 14 15 13 12 9 0 9 2
7 13 9 1 9 1 0 9
5 13 0 9 1 9
10 0 9 14 15 13 1 9 1 9 2
16 15 13 1 0 9 1 3 2 15 9 15 13 14 13 3 2
9 3 10 9 15 13 1 12 9 2
25 9 1 9 14 13 9 14 13 9 1 15 2 15 14 13 0 9 2 13 1 9 2 11 2 2
15 9 1 9 1 0 9 13 1 12 9 7 13 12 9 2
12 1 9 14 4 13 7 9 1 9 0 9 2
13 1 10 9 9 15 13 9 15 7 1 0 9 2
16 1 12 9 3 9 14 13 1 9 3 2 13 3 3 3 2
10 1 12 9 9 13 9 1 10 9 2
3 9 13 9
7 9 1 9 13 0 1 9
11 15 13 9 1 11 1 9 1 0 9 2
7 9 14 13 9 2 13 11
10 10 9 14 13 9 15 2 13 9 2
12 15 13 9 1 2 11 2 7 2 11 2 2
8 2 11 2 1 9 1 9 11
6 9 13 9 1 9 15
24 0 9 4 13 1 9 1 9 1 9 1 0 0 9 11 11 2 13 9 1 0 9 3 2
15 15 13 9 1 9 15 2 16 9 15 1 9 13 0 2
18 11 15 13 1 0 9 2 1 14 13 9 15 2 7 3 13 9 2
7 9 13 7 9 11 11 2
16 3 3 6 13 3 10 1 9 4 13 1 0 9 1 11 2
9 3 13 2 16 3 3 13 9 2
7 13 14 3 1 0 9 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
16 2 3 13 1 10 0 9 2 7 3 6 13 14 13 15 2
6 1 9 3 14 13 2
11 11 11 2 12 9 2 2 9 2 11 2
6 1 9 13 12 9 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
10 3 3 6 4 13 14 13 1 9 2
11 11 11 2 12 9 2 2 9 2 11 2
8 1 15 13 3 3 1 15 2
10 13 13 0 9 14 13 14 13 9 2
13 11 11 2 12 9 2 2 9 1 11 2 11 2
3 2 6 2
9 2 6 2 6 4 13 1 9 2
15 3 13 3 1 15 2 7 7 3 6 4 15 13 3 2
12 11 11 2 12 9 2 2 0 9 2 11 2
9 2 6 2 3 3 4 15 13 2
10 3 13 3 14 13 7 14 15 13 2
4 11 13 0 9
20 9 13 2 16 11 13 9 1 0 15 9 1 9 2 15 13 1 0 9 2
14 9 13 3 1 9 1 11 2 11 2 11 7 11 2
6 9 13 14 13 11 11
18 15 3 14 13 2 1 1 9 13 0 9 0 9 7 13 9 15 2
14 15 13 14 13 3 7 0 9 1 0 9 11 11 2
24 11 11 2 9 1 11 2 13 1 10 9 2 16 9 13 14 13 9 15 1 9 1 9 2
21 1 1 9 3 13 9 15 1 11 11 2 9 11 4 13 14 13 1 9 15 2
26 1 9 1 0 9 9 13 9 1 9 15 1 9 2 7 1 0 9 1 11 9 1 11 4 13 2
8 11 11 13 1 0 9 1 11
24 0 15 9 11 11 7 9 11 11 13 3 1 11 2 1 14 13 9 1 0 9 1 9 2
14 1 9 2 9 1 9 2 9 3 13 9 1 9 2
20 0 9 4 13 1 0 0 9 1 9 9 1 0 9 11 2 13 0 9 2
14 11 11 4 13 1 9 2 3 15 13 1 9 15 2
18 15 3 4 13 1 9 7 1 9 9 15 15 13 1 2 0 2 2
14 0 9 0 9 1 0 9 7 9 13 9 1 9 2
22 1 9 2 0 1 11 2 9 13 2 16 10 9 4 13 9 1 2 0 9 2 2
14 15 13 0 9 1 0 9 1 0 9 1 12 9 2
25 3 0 9 2 11 2 13 9 1 0 9 14 13 9 1 9 1 11 7 1 0 9 1 11 2
10 3 3 7 11 13 2 16 13 9 2
11 10 9 13 1 0 9 1 9 1 11 2
15 1 15 13 3 11 2 3 0 2 0 7 3 3 0 2
8 15 13 14 4 13 3 1 9
8 9 3 15 13 1 0 9 2
30 7 16 16 3 6 13 14 13 10 0 9 1 11 7 11 2 3 0 9 1 11 14 13 0 2 13 2 11 2 2
10 9 1 2 11 2 15 13 1 9 11
10 11 11 3 13 1 9 1 9 11 2
19 9 1 0 9 1 9 1 11 14 13 14 15 13 9 1 9 1 9 2
13 9 13 3 0 1 0 9 7 9 1 0 9 2
22 9 2 15 13 14 15 13 9 2 14 15 13 7 9 2 13 9 1 9 11 11 2
11 1 12 9 7 0 9 14 13 1 9 2
7 12 9 14 13 0 9 2
41 1 9 1 9 14 4 13 0 9 1 11 11 2 2 9 2 2 2 11 11 2 2 7 0 9 2 2 7 0 9 1 0 9 1 11 2 0 1 11 11 2
16 0 9 1 9 2 9 7 0 9 14 4 13 1 0 9 2
19 9 14 13 9 1 9 1 9 1 0 9 7 9 1 9 2 11 2 2
13 1 9 14 13 3 12 9 2 13 1 0 9 2
14 9 1 9 1 0 9 15 13 1 0 9 1 9 2
6 13 11 1 9 1 9
18 1 0 0 9 3 14 13 3 9 1 9 0 9 1 0 9 11 2
8 3 14 13 7 9 1 9 2
20 1 9 9 1 0 9 1 2 11 2 13 9 1 9 11 7 11 11 11 2
5 13 15 3 0 2
12 14 13 9 1 9 13 1 14 13 9 1 9
39 0 15 9 11 11 13 1 0 9 11 11 1 0 9 1 0 9 1 12 1 0 9 1 9 1 0 9 9 12 9 2 15 13 1 11 2 11 2 2
13 11 13 1 0 9 2 16 11 3 13 0 9 2
24 3 7 3 13 3 14 13 9 1 9 2 9 7 9 1 0 9 1 3 1 9 1 9 2
4 11 13 1 9
14 11 14 13 1 0 9 3 2 13 1 0 11 3 2
12 9 2 11 2 13 14 4 13 3 1 9 2
20 16 15 13 9 1 0 9 2 0 9 14 13 1 0 0 9 2 13 9 2
7 1 9 9 13 10 9 2
19 9 15 13 1 0 9 1 9 2 13 0 9 1 9 9 9 11 11 2
6 13 0 0 9 3 9
2 11 11
22 9 1 9 1 0 0 9 7 0 9 14 15 13 1 9 1 0 9 2 13 9 2
10 9 1 9 14 15 13 3 12 9 2
15 0 9 1 12 9 14 13 14 13 9 15 2 3 13 2
7 9 13 14 13 12 9 2
6 3 15 13 12 9 2
6 9 4 13 1 11 2
24 1 11 7 9 15 2 11 2 13 7 9 1 11 11 2 11 11 2 15 13 9 1 9 2
9 12 9 9 13 1 11 1 12 9
8 0 9 13 12 9 9 1 9
21 12 9 9 4 13 1 11 3 1 0 12 9 2 13 9 1 9 11 11 3 2
20 1 9 0 9 1 11 13 11 1 9 1 9 1 9 1 0 9 1 9 2
19 9 4 13 1 10 9 7 1 9 13 0 9 2 13 1 0 15 9 2
27 1 1 13 9 1 11 2 11 15 13 7 1 12 9 9 1 10 9 1 15 2 13 3 7 11 11 2
18 9 13 9 1 9 12 9 2 15 4 13 1 0 9 7 0 9 2
12 11 13 2 11 2 1 9 1 2 0 11 2
10 10 9 3 13 12 9 1 0 0 9
17 1 9 1 9 1 9 9 11 13 9 1 2 11 2 1 9 2
22 15 15 13 14 13 1 0 9 1 9 2 15 3 6 15 13 1 9 1 0 9 2
21 3 15 13 1 0 9 1 9 7 9 3 1 3 12 9 1 9 1 0 9 2
8 2 11 2 14 13 9 1 11
10 9 13 1 0 9 2 11 11 2 2
15 3 15 13 9 1 0 9 1 9 1 0 9 1 11 2
11 9 1 10 9 1 9 14 13 12 9 2
21 0 1 9 0 9 1 0 9 14 4 13 1 9 1 0 9 2 15 13 3 2
21 13 9 1 9 1 9 2 16 1 12 9 1 0 9 0 9 3 13 12 9 2
11 12 9 13 0 9 1 0 9 1 11 2
19 9 1 11 13 3 0 2 7 1 11 7 11 9 13 3 1 12 9 2
15 0 9 14 15 13 1 12 9 9 2 1 0 12 9 2
37 9 13 14 13 9 1 9 2 9 2 0 0 9 2 9 1 9 2 9 2 3 0 15 9 4 13 1 0 9 2 13 11 11 1 0 9 2
7 11 13 9 7 13 9 2
12 13 15 3 2 1 14 13 9 1 9 1 9
23 1 10 9 3 9 15 13 9 1 11 2 7 1 0 9 15 13 1 9 7 15 13 2
10 11 11 2 9 1 0 9 1 11 2
8 0 13 14 13 2 16 13 9
1 9
10 11 11 4 13 1 0 9 1 11 2
12 13 7 0 9 1 11 1 9 2 11 2 2
13 2 13 9 14 15 13 2 6 13 1 0 9 2
5 7 6 4 13 2
12 13 1 11 2 1 14 15 13 14 13 3 2
4 3 14 13 2
7 15 13 1 9 1 9 2
9 7 16 13 14 13 2 14 13 2
16 2 13 14 15 15 4 14 13 9 2 1 14 15 13 9 2
3 2 6 2
3 2 6 2
14 3 13 1 9 2 9 13 14 9 13 1 10 9 2
11 16 13 2 3 3 15 15 13 0 9 2
16 2 3 0 9 15 13 2 16 13 3 0 7 3 0 9 2
10 14 0 9 1 9 13 14 13 9 2
6 2 6 2 3 13 2
8 1 9 9 13 9 1 9 2
18 3 3 15 9 13 1 9 2 9 2 9 2 9 2 9 2 9 2
9 2 13 9 2 9 13 14 9 2
10 2 0 13 14 13 2 16 13 9 2
4 2 7 15 2
9 2 7 4 14 13 1 0 9 2
15 3 3 14 13 9 1 12 9 2 9 1 9 2 9 2
12 7 9 13 2 16 9 13 14 6 15 13 2
15 11 13 3 0 9 2 13 9 2 15 13 14 15 13 2
9 2 10 9 13 0 15 0 9 2
13 2 13 14 9 3 9 2 1 14 13 3 9 2
5 7 0 13 9 2
7 2 3 14 13 0 9 2
15 12 12 0 9 13 2 13 7 13 3 3 1 12 9 2
5 13 15 0 9 2
12 3 13 14 15 13 9 1 12 9 1 9 2
12 13 14 13 3 14 15 13 0 9 1 9 2
4 9 1 11 11
4 0 9 13 11
30 9 3 13 14 13 9 2 3 16 13 2 16 9 1 0 9 14 15 13 1 0 9 13 3 0 9 1 10 9 2
14 15 3 6 13 9 2 13 9 2 9 7 9 2 2
16 15 13 14 13 9 1 9 2 16 15 13 3 1 11 11 2
8 0 9 1 11 13 1 0 9
18 3 9 2 0 7 0 15 1 0 9 2 10 13 2 0 9 2 2
25 1 9 3 13 3 2 16 1 10 9 6 13 2 16 6 3 0 9 13 9 2 15 15 13 2
8 0 9 13 2 0 9 2 2
11 11 7 0 9 11 11 3 13 0 9 2
8 9 1 11 13 2 11 12 2
25 9 1 11 11 1 0 2 11 12 2 11 11 13 2 16 14 13 9 1 9 1 9 11 11 2
7 12 13 3 1 0 9 2
3 13 15 9
33 13 14 15 1 0 9 2 14 13 0 9 7 3 1 9 2 3 9 13 1 0 9 7 13 0 9 2 15 14 15 13 9 2
25 16 1 9 15 15 4 13 1 0 15 9 2 15 14 13 9 7 9 15 7 14 13 9 15 2
32 0 2 0 2 0 7 0 2 15 14 15 2 13 2 1 9 1 9 7 9 2 3 9 15 13 7 3 9 15 13 9 2
18 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
2 0 9
21 0 11 15 13 1 9 11 2 11 2 1 9 1 9 2 15 15 13 1 9 2
16 16 13 9 2 13 0 9 2 13 9 7 15 13 1 9 2
8 0 13 1 0 9 1 11 2
7 11 14 13 1 9 1 9
19 1 0 9 3 9 1 11 14 13 9 2 0 1 9 1 9 1 9 2
12 15 13 14 15 13 1 9 1 9 1 9 2
1 9
14 1 9 1 10 0 9 14 13 9 15 1 0 9 2
3 9 1 9
5 2 9 15 13 2
3 2 3 2
5 2 1 12 9 2
8 2 14 2 3 13 1 9 2
9 9 13 1 11 2 11 2 1 9
16 11 13 2 16 14 13 14 15 13 0 15 0 9 1 11 2
16 15 13 7 0 9 2 3 16 3 4 13 3 9 12 9 2
25 1 9 1 12 9 1 11 2 11 2 1 12 9 0 9 1 9 14 4 13 2 13 9 11 2
11 11 11 3 13 14 13 1 0 9 3 2
15 15 13 11 1 9 9 0 0 9 14 13 3 1 11 2
8 6 13 2 16 15 13 0 2
13 1 11 13 9 1 9 11 1 11 2 13 11 2
30 1 15 9 14 13 0 0 9 1 9 1 9 2 15 13 14 13 12 9 2 7 9 1 9 13 14 4 13 3 2
7 9 13 2 16 14 13 2
19 9 1 9 13 9 1 0 9 2 3 1 15 13 9 1 9 1 11 2
14 9 1 11 1 9 1 11 4 13 1 0 9 11 2
15 1 9 1 11 13 2 16 3 14 13 0 9 1 11 2
9 15 14 13 1 11 7 0 9 2
17 1 0 9 14 4 13 0 9 1 9 1 11 1 12 0 9 2
6 14 13 9 1 0 9
29 15 14 13 1 9 1 0 0 9 1 0 0 9 2 9 1 9 2 11 2 1 0 9 2 0 1 0 9 2
17 12 9 1 9 11 4 13 1 9 7 9 1 9 1 0 9 2
15 9 13 2 16 1 11 6 4 13 9 1 0 15 9 2
11 1 10 9 13 7 9 1 11 2 11 2
17 11 7 9 15 11 13 1 2 11 2 1 11 2 7 13 9 2
12 3 15 13 1 9 15 11 7 9 15 11 2
9 1 10 9 13 0 9 1 11 2
14 9 14 15 13 7 13 13 1 9 1 11 7 11 2
24 1 12 4 13 9 1 9 1 0 9 7 9 1 0 0 9 2 15 13 1 12 9 9 2
12 1 0 9 11 13 14 13 3 1 0 9 2
10 11 2 11 2 13 1 11 11 11 11
15 1 0 9 13 0 1 0 9 1 11 1 9 1 9 2
34 1 9 16 15 13 3 3 3 2 1 10 9 1 9 14 15 13 11 2 7 1 15 3 13 14 15 13 9 1 9 1 0 11 2
22 1 0 0 9 1 11 15 13 3 3 12 9 2 16 3 4 13 1 12 9 9 2
5 9 13 0 9 2
9 13 14 9 14 4 13 1 9 2
11 11 11 2 12 9 2 2 9 2 11 2
3 2 6 2
11 11 11 2 12 9 2 2 9 2 11 2
3 2 6 2
13 1 15 9 6 13 14 13 0 1 10 10 9 2
9 0 9 13 14 15 13 1 9 2
11 11 11 2 12 9 2 2 9 2 11 2
3 2 6 2
11 3 13 0 2 7 9 13 0 15 9 2
18 7 3 1 9 2 16 9 13 9 1 9 7 15 13 1 10 9 2
11 11 11 2 12 9 2 2 9 2 11 2
10 2 6 2 13 14 15 13 1 9 2
12 10 9 14 13 0 2 3 9 3 15 13 2
11 11 11 2 12 9 2 2 9 2 11 2
6 2 6 2 6 13 2
11 11 11 2 12 9 2 2 9 2 11 2
10 2 6 2 3 1 9 3 13 0 2
3 2 6 2
13 3 9 13 9 2 15 13 14 15 13 1 9 2
12 9 6 13 9 2 15 13 14 13 10 9 2
11 11 11 2 12 9 2 2 9 2 11 2
3 2 6 2
19 9 13 14 15 13 1 9 2 3 6 4 13 2 16 9 13 9 0 2
11 11 11 2 12 9 2 2 9 2 11 2
3 2 6 2
6 9 1 9 13 0 9
18 3 0 9 11 13 9 1 0 9 1 0 9 2 0 1 0 9 2
30 1 0 9 1 9 2 0 9 2 2 11 11 2 13 2 16 1 12 9 9 1 9 1 9 11 13 0 0 9 2
8 9 13 0 0 9 1 9 2
6 9 1 11 13 0 9
8 9 3 4 13 7 9 4 13
10 15 13 2 16 9 6 13 0 9 2
21 9 13 2 16 1 9 9 1 0 9 11 0 9 13 9 1 0 9 1 11 2
19 1 15 9 13 2 16 13 3 9 1 9 2 3 9 7 12 9 9 2
41 9 1 9 13 11 11 2 15 4 13 9 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2
14 9 15 13 1 0 9 2 0 1 9 9 7 9 2
7 0 9 13 1 11 11 2
15 3 13 14 15 13 3 13 9 7 3 13 9 1 9 2
8 13 15 3 9 7 0 9 2
11 0 15 9 3 14 15 13 1 0 9 2
25 2 11 2 13 9 2 15 0 11 6 4 13 3 1 0 15 9 1 11 1 9 1 0 9 2
24 1 0 9 1 0 9 2 11 2 3 4 13 0 9 1 9 9 11 11 7 9 11 11 2
15 3 1 0 0 9 12 1 0 15 9 13 7 0 9 2
12 1 9 1 9 4 13 0 9 1 11 11 2
13 1 0 9 15 13 9 7 0 15 9 1 9 2
17 1 0 12 9 1 10 0 9 4 13 10 1 0 9 1 9 2
22 3 13 14 15 13 9 1 9 1 11 7 0 0 9 1 9 1 0 9 1 9 2
22 3 1 12 9 10 9 1 11 12 14 15 13 0 9 1 11 2 9 1 9 2 2
14 9 1 9 1 11 11 4 13 1 0 9 1 9 2
13 10 15 4 13 1 10 9 14 13 1 10 9 2
16 11 11 13 0 1 9 1 9 1 0 9 1 9 1 11 2
10 1 9 15 13 12 11 1 0 9 2
8 0 13 11 11 2 11 2 2
14 11 11 15 13 0 1 9 7 0 1 9 1 9 2
7 11 11 13 1 11 1 11
29 1 9 1 9 15 1 11 11 11 14 13 7 1 9 1 2 11 2 11 11 2 9 1 15 13 9 12 12 2
21 16 15 13 1 9 2 11 14 13 0 9 1 0 9 1 9 1 2 11 2 2
9 9 13 1 12 9 1 0 9 2
30 1 9 11 11 1 9 1 11 13 9 1 11 2 11 2 11 2 11 7 11 2 3 13 7 9 1 9 11 11 2
3 13 15 9
32 16 15 13 1 0 9 2 14 13 0 9 2 13 14 9 0 9 2 6 13 14 15 14 13 0 9 7 13 14 15 3 2
18 13 9 7 0 15 9 7 3 15 13 1 10 9 1 0 1 15 2
22 1 9 9 14 13 9 15 3 1 9 2 7 7 14 15 13 9 1 3 0 9 2
26 0 2 0 1 0 9 2 7 1 9 1 9 1 9 2 15 14 15 13 1 15 1 9 7 9 2
24 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
14 15 13 9 11 11 3 1 9 1 0 9 1 9 2
17 10 9 6 13 1 11 7 15 6 4 13 1 15 2 13 11 2
20 10 9 11 14 13 9 1 10 9 1 9 1 9 2 13 0 9 11 11 2
15 15 13 9 1 0 9 7 9 1 9 1 9 7 9 2
14 13 9 1 11 7 11 2 13 9 1 11 11 11 2
4 0 9 13 2
10 13 14 15 13 1 9 2 13 11 2
3 9 13 2
21 3 1 15 13 3 3 2 16 3 9 15 13 1 9 7 13 14 13 1 15 2
6 11 11 13 9 1 9
10 0 9 13 1 0 9 1 9 9 2
13 11 11 15 13 1 9 1 0 9 1 0 9 2
13 1 9 1 0 9 2 0 9 2 13 11 11 2
12 0 9 1 11 1 0 9 13 1 11 11 2
3 9 1 9
6 9 13 9 1 9 2
14 15 13 0 15 9 2 3 4 13 1 9 1 9 2
22 11 13 2 16 1 9 2 1 15 4 13 9 2 15 2 4 13 14 13 9 2 2
5 0 9 13 1 11
5 9 13 1 0 9
10 1 11 13 9 2 15 3 13 9 2
13 15 13 0 9 1 11 7 9 1 11 11 11 2
14 16 15 13 2 15 3 14 13 1 15 2 13 11 2
12 1 15 9 1 9 15 14 13 1 0 9 2
2 11 11
9 9 7 9 13 1 9 2 13 9
17 7 12 9 4 13 9 1 0 9 1 11 2 15 13 9 15 2
20 15 13 7 9 1 0 9 1 9 2 3 7 1 9 1 9 1 0 9 2
19 13 9 7 1 0 0 9 1 9 2 9 7 9 2 0 9 7 0 2
32 9 1 9 2 9 1 9 7 1 0 9 1 9 13 3 12 12 10 9 7 9 1 0 0 9 1 9 2 13 3 3 2
29 9 13 9 1 9 2 16 0 9 13 12 0 9 2 7 1 12 9 2 13 9 1 0 9 1 9 11 11 2
14 9 14 15 13 1 9 1 9 1 0 9 1 9 2
12 0 9 1 15 3 6 4 13 2 13 15 2
7 9 13 1 12 9 1 9
17 0 9 1 9 13 1 9 1 9 3 1 12 9 2 13 9 2
10 9 1 9 0 9 13 1 12 9 2
5 9 1 9 13 9
26 1 12 9 1 0 9 1 9 13 1 3 0 9 2 13 3 9 11 11 1 0 9 2 11 2 2
12 0 13 9 1 0 9 7 1 0 0 11 2
11 1 0 13 10 9 0 9 14 4 13 2
23 15 13 2 16 1 0 9 9 9 14 13 12 9 2 15 13 1 1 12 9 3 3 2
17 13 15 12 12 9 7 0 9 1 3 12 9 9 2 13 9 2
11 9 1 2 0 9 2 13 1 12 9 2
6 13 9 1 9 7 9
17 9 1 3 1 0 9 1 9 4 13 1 12 9 1 0 9 2
5 15 13 11 3 2
12 3 13 9 1 12 9 1 9 1 0 9 2
11 0 9 1 9 4 13 1 12 9 9 2
12 0 9 1 9 13 1 9 7 0 0 9 2
18 1 9 9 1 9 15 4 13 1 12 9 1 0 9 1 0 9 2
11 9 13 7 1 9 1 0 9 7 9 2
6 0 9 14 13 9 15
28 15 13 11 11 2 9 1 9 1 0 11 7 0 11 1 9 2 1 9 15 1 9 11 11 1 11 3 2
13 11 13 9 14 13 1 9 2 9 7 0 9 2
6 13 9 1 9 1 3
2 11 11
35 1 0 9 2 11 2 2 2 11 2 2 11 11 2 11 11 7 2 9 2 14 13 1 3 1 10 2 15 13 14 13 0 9 3 2
10 0 1 9 14 13 11 11 7 11 2
11 9 14 13 9 1 9 3 1 0 9 2
20 14 13 7 0 9 2 1 14 13 14 13 1 9 0 9 2 13 9 11 2
12 3 13 9 1 9 15 2 13 0 9 11 2
20 9 13 1 9 1 11 1 9 1 0 9 1 9 2 11 2 1 12 9 2
13 0 13 1 9 15 2 9 15 7 1 0 9 2
12 1 9 13 9 1 3 2 1 15 0 13 2
7 1 12 9 13 12 9 2
5 15 13 1 9 2
3 11 13 2
9 13 2 13 9 7 15 13 1 9
16 1 9 1 9 15 2 11 13 3 1 0 9 1 0 9 2
4 3 13 9 2
17 9 11 2 12 9 2 15 13 1 9 7 13 9 14 6 13 2
6 3 15 4 4 13 2
11 1 0 11 13 1 9 2 13 1 11 2
10 9 15 13 11 14 6 13 0 9 2
14 1 9 9 1 9 4 13 1 0 9 1 0 9 2
6 9 9 15 13 1 9
10 1 9 9 13 0 15 2 11 2 2
12 13 15 2 16 9 4 15 13 1 0 9 2
13 3 4 13 1 9 1 0 9 7 4 15 13 2
11 1 9 4 13 12 9 7 9 1 9 2
20 9 13 1 9 1 12 9 1 9 1 9 2 11 11 2 7 2 11 2 2
5 11 13 1 9 2
9 11 4 13 1 9 1 0 9 2
15 13 15 2 16 9 4 13 9 1 9 7 15 13 9 2
7 11 11 2 9 1 11 2
10 11 15 13 0 2 7 9 13 15 0
15 1 9 1 9 13 9 2 15 13 14 13 1 0 9 2
12 2 9 11 2 11 13 14 13 9 1 11 2
20 1 0 9 0 9 1 9 1 11 7 11 4 13 9 15 1 0 9 3 2
21 2 16 3 3 15 13 1 9 1 9 1 11 2 13 14 9 14 13 0 9 2
6 2 3 14 13 9 2
11 13 15 3 2 16 13 14 15 13 3 2
9 2 1 0 9 11 4 13 9 2
22 2 1 9 1 9 1 9 9 11 11 15 13 3 14 15 13 0 9 1 0 9 2
2 15 2
8 3 15 13 7 13 0 9 2
14 3 9 6 13 14 13 10 9 2 0 9 1 9 2
16 9 1 9 1 0 9 1 0 9 4 13 9 1 0 9 2
16 1 15 14 15 13 9 1 9 2 15 3 13 1 0 9 2
22 3 0 9 14 13 9 1 0 15 9 2 9 1 9 2 9 2 9 1 0 9 2
11 2 3 13 0 9 1 9 1 0 9 2
9 2 3 13 14 15 13 10 9 2
13 3 0 9 1 15 15 13 1 0 0 0 9 2
16 2 13 14 9 3 0 9 14 2 13 2 9 1 0 9 2
14 2 1 10 9 13 14 3 14 13 9 1 0 9 2
11 2 15 13 9 2 15 13 9 1 11 2
10 6 13 3 14 15 13 7 1 15 2
10 2 1 3 1 9 6 4 13 9 2
28 1 15 13 2 16 13 1 0 9 2 7 3 13 9 2 15 13 14 15 13 1 0 7 0 1 15 9 2
14 3 15 13 12 9 1 0 9 14 15 13 1 9 2
10 10 9 14 13 3 1 9 1 9 2
13 2 10 0 9 3 15 13 7 9 2 7 9 2
10 1 0 9 13 14 13 9 12 9 2
26 16 15 13 9 1 9 14 2 14 15 13 3 0 9 2 15 13 14 13 1 9 1 9 7 9 2
9 2 3 1 15 13 14 13 9 2
11 9 13 0 2 15 13 1 3 0 9 2
18 2 13 15 2 16 1 11 13 14 13 0 9 1 9 1 0 9 2
10 3 14 13 10 9 3 1 10 9 2
9 2 11 6 4 13 1 10 9 2
10 3 3 14 15 13 14 15 13 3 2
12 2 1 9 6 13 9 2 3 3 6 13 2
15 3 16 16 3 13 9 1 0 2 1 9 14 15 13 2
7 11 11 2 9 2 11 2
10 2 9 15 6 15 13 14 13 9 2
10 13 15 9 7 15 15 13 1 9 2
12 11 11 2 2 12 9 2 2 9 2 11 2
5 2 14 13 9 2
12 11 11 2 2 12 9 2 2 9 2 11 2
12 11 11 2 2 12 9 2 2 9 2 11 2
9 2 14 13 1 10 9 1 9 2
12 11 11 2 2 12 9 2 2 9 2 11 2
11 2 6 13 9 7 10 9 13 14 13 2
18 14 7 14 6 13 14 12 9 2 3 13 9 2 1 14 13 9 2
12 11 11 2 2 12 9 2 2 9 2 11 2
14 2 3 4 13 12 9 7 3 1 9 6 4 13 2
12 11 11 2 2 12 9 2 2 9 2 11 2
12 11 11 2 2 12 9 2 2 9 2 11 2
6 2 6 2 13 15 2
9 15 6 15 13 14 15 13 9 2
12 11 11 2 2 12 9 2 2 9 2 11 2
3 2 6 2
6 6 13 9 1 9 2
4 13 3 9 11
16 0 9 11 4 13 3 1 0 1 9 1 9 2 13 11 2
17 0 9 3 13 1 9 1 9 1 11 1 0 9 1 0 11 2
18 0 9 13 2 16 15 13 14 13 1 9 7 1 9 1 0 15 9
16 15 7 14 13 0 9 2 14 15 15 13 0 7 0 1 15
5 11 11 2 9 2
8 6 13 3 14 13 1 0 9
8 3 13 1 2 0 9 2 2
6 13 2 16 13 0 2
10 15 15 13 1 0 9 1 9 3 2
4 2 13 15 2
12 1 11 10 9 13 0 1 0 9 1 9 2
15 7 14 15 13 14 13 3 13 9 2 3 3 3 0 2
10 3 1 10 9 15 13 1 10 9 2
4 3 2 3 2
6 0 13 9 7 9 2
14 10 2 15 14 13 2 6 13 9 1 9 1 11 2
7 2 4 14 13 0 9 2
6 2 6 2 13 15 2
26 16 1 10 9 15 13 15 14 1 9 2 3 15 14 2 13 2 16 14 13 7 9 1 10 9 2
4 15 13 0 2
10 2 13 14 15 4 9 15 1 9 2
13 2 6 2 9 15 1 9 6 4 13 10 9 2
9 13 1 0 9 2 1 0 11 2
14 0 9 2 15 13 3 2 13 0 9 2 0 9 2
12 10 2 15 13 1 9 1 9 2 13 0 2
6 11 11 15 13 1 11
13 15 14 13 1 9 2 11 2 1 9 1 11 2
7 9 1 9 13 11 11 2
17 11 13 3 1 9 1 9 2 15 4 13 1 9 1 0 9 2
8 9 1 11 11 13 9 1 9
27 0 9 1 12 0 9 1 9 2 11 11 2 12 14 15 13 1 9 1 9 7 9 2 0 9 2 2
17 3 9 1 9 13 9 1 0 0 9 7 15 4 13 1 9 2
17 9 1 11 11 11 13 0 9 1 11 9 14 13 1 10 9 2
18 1 15 14 13 0 9 1 11 11 2 13 9 11 11 7 11 11 2
15 1 9 1 9 1 9 14 15 13 0 9 7 0 9 2
15 14 13 9 2 9 2 0 1 0 9 7 0 0 9 2
27 13 4 7 0 9 1 0 9 1 0 9 2 15 13 14 13 12 12 9 2 13 1 9 2 11 2 2
25 11 3 13 9 1 9 1 9 1 9 2 1 15 0 15 9 15 13 1 9 14 13 10 9 2
16 4 15 13 11 14 13 1 15 1 9 2 7 3 15 15 13
13 13 14 13 3 9 1 11 2 11 2 11 2 11
8 6 13 0 9 2 7 15 13
23 0 9 1 2 11 2 11 11 13 9 1 11 1 9 1 9 1 0 9 1 10 9 2
7 1 9 13 12 0 9 2
7 15 13 0 9 1 15 2
14 13 4 2 16 10 9 1 11 7 11 13 1 15 2
10 13 13 9 1 15 13 0 9 1 11
17 9 4 13 1 0 9 1 9 11 11 11 7 0 9 11 11 2
29 1 0 9 1 9 2 11 2 0 9 13 3 9 7 3 13 9 1 12 9 2 15 6 13 1 9 1 9 2
19 0 9 1 9 1 2 0 2 11 11 1 0 12 9 3 13 0 9 2
7 3 13 2 3 13 1 9
7 0 9 15 13 1 9 2
6 3 9 13 9 1 11
10 9 2 11 2 13 1 9 11 11 2
16 15 4 13 1 0 9 2 7 9 15 13 1 10 1 9 2
7 0 9 2 13 2 0 9
27 0 9 2 11 2 13 9 1 9 2 15 3 15 13 0 9 2 9 2 15 13 0 9 2 13 11 2
16 9 1 9 11 11 13 9 1 12 9 9 1 0 15 9 2
13 0 9 1 9 13 1 9 1 9 1 0 9 2
5 9 7 9 13 11
6 9 1 0 9 13 9
23 9 1 9 2 9 9 2 9 1 0 9 7 9 13 11 1 12 9 7 12 9 3 2
18 9 13 1 9 1 9 1 0 9 7 9 1 0 0 9 1 11 2
10 9 13 9 7 15 13 9 1 9 2
8 9 7 1 0 9 13 9 2
10 1 9 1 9 15 13 9 11 11 2
8 3 11 11 15 13 1 0 2
8 0 2 11 15 13 1 9 2
11 9 13 1 9 1 2 0 11 11 2 2
12 1 15 9 11 3 13 1 10 9 1 9 2
13 0 9 15 13 1 0 9 1 9 1 0 9 2
8 15 13 1 9 1 9 11 2
30 1 2 11 2 12 13 11 11 2 11 11 2 9 11 11 2 9 1 11 11 11 2 11 11 2 11 11 7 0 2
8 9 13 1 0 9 1 11 2
6 9 13 1 9 1 9
25 12 9 7 9 2 0 1 9 15 1 11 2 13 1 9 1 0 9 1 11 2 13 11 9 2
11 15 4 13 1 9 1 9 1 0 9 2
12 9 13 9 2 13 9 7 15 13 1 9 2
6 9 1 9 4 13 2
8 3 4 13 12 9 1 11 2
4 9 11 11 2
3 6 13 0
12 15 13 0 9 2 13 0 9 7 13 9 2
6 1 12 9 15 13 2
17 1 12 9 9 3 15 13 7 13 2 16 9 15 13 3 0 2
5 7 12 13 3 2
19 13 15 14 15 13 1 0 9 2 1 14 15 13 1 10 9 1 11 2
9 9 13 1 9 2 13 0 9 2
17 13 9 14 13 2 13 15 1 0 9 7 13 9 1 10 9 2
20 1 11 13 9 1 12 9 2 9 15 13 1 12 9 2 1 14 13 3 2
18 0 14 13 7 1 0 9 2 7 1 9 1 9 2 16 15 13 2
14 16 6 13 14 13 0 0 0 9 2 9 13 9 2
14 14 10 0 15 9 15 13 0 9 7 0 15 9 2
14 9 13 9 1 0 9 9 2 13 1 9 0 9 2
12 9 9 13 1 15 2 13 15 9 11 11 2
10 1 10 9 9 15 13 14 13 9 2
5 13 7 0 9 2
10 1 10 9 15 13 12 9 9 3 2
11 3 13 2 16 0 1 9 13 0 9 2
11 14 13 14 9 9 1 9 2 11 2 2
11 11 11 2 12 9 2 2 9 2 11 2
14 1 9 13 14 13 14 13 2 3 13 3 14 13 2
11 11 11 2 12 9 2 2 9 2 11 2
12 3 1 9 3 4 13 14 13 1 9 15 2
11 11 11 2 12 9 2 2 9 2 11 2
5 2 9 15 13 2
11 11 11 2 12 9 2 2 9 2 11 2
9 2 16 13 0 9 2 4 13 2
4 13 10 9 2
7 9 3 14 13 1 9 2
11 11 11 2 12 9 2 2 9 2 11 2
9 2 6 2 3 14 13 1 9 2
6 9 3 3 15 13 2
12 14 9 2 15 15 13 2 14 15 13 3 2
6 7 15 6 15 13 2
15 13 1 0 9 14 15 15 13 14 13 9 1 9 9 2
11 11 11 2 12 9 2 2 9 2 11 2
8 2 1 11 13 7 14 13 2
17 7 14 7 14 13 3 2 6 4 13 2 3 6 13 10 9 2
12 11 11 2 12 9 2 2 0 9 2 11 2
9 3 13 2 16 13 1 10 9 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
5 2 13 3 9 2
16 7 16 13 14 15 13 2 1 9 4 13 14 13 9 9 2
5 13 9 1 0 9
16 1 9 1 0 9 9 13 2 16 4 13 1 9 1 9 2
11 15 3 13 14 13 3 13 9 1 9 2
34 3 9 2 11 2 13 9 2 16 9 4 13 1 11 2 3 16 11 11 13 9 2 9 2 7 1 9 15 13 9 1 9 11 2
14 12 9 9 13 0 11 2 16 9 15 13 1 0 2
14 6 15 13 10 7 14 13 9 1 9 1 9 15 2
20 9 1 11 1 9 1 9 9 12 1 9 1 0 9 13 11 7 11 11 2
16 11 6 13 7 9 15 1 0 9 3 1 9 2 11 2 2
8 1 9 11 15 6 4 4 13
13 6 4 15 13 1 15 7 6 4 13 1 15 2
4 13 15 3 2
17 7 4 13 3 1 9 2 7 14 15 13 1 15 7 14 13 2
14 11 11 7 11 11 13 2 16 15 13 2 13 11 2
25 9 9 0 7 0 2 15 6 4 13 0 9 1 3 9 2 14 13 9 15 2 13 11 3 2
25 3 6 4 13 0 9 1 1 12 9 7 0 9 1 0 1 9 12 9 2 13 3 1 11 2
21 9 13 2 16 0 9 15 13 1 9 1 0 9 2 15 14 13 9 1 9 2
8 0 9 13 1 12 9 1 9
10 9 13 3 9 1 11 1 0 9 2
30 0 9 2 11 11 2 1 0 11 2 9 1 2 11 2 2 13 9 1 3 2 13 0 9 1 9 11 11 3 2
14 0 9 13 9 1 12 9 0 9 7 3 15 13 2
14 9 1 9 13 1 9 1 9 11 2 1 9 11 2
12 1 9 13 7 0 9 11 2 11 2 11 2
23 1 1 0 9 9 1 9 1 0 9 13 12 9 1 9 1 0 9 2 13 11 11 2
16 0 9 3 13 3 14 15 13 3 9 1 9 1 0 9 2
22 15 14 13 1 9 1 0 9 1 9 15 7 14 13 0 9 1 9 2 13 9 2
31 9 4 13 9 1 2 11 2 1 2 9 2 2 3 1 9 15 6 4 13 0 9 2 0 1 0 9 1 0 9 2
13 0 2 9 2 13 3 9 1 11 2 13 11 2
10 0 9 13 0 9 7 3 13 14 13
18 0 9 13 2 16 1 0 9 1 0 9 9 4 13 3 12 9 2
6 3 3 13 3 1 9
18 12 9 9 1 15 4 13 1 3 0 9 1 9 7 9 1 9 2
1 9
12 1 0 0 9 1 0 9 9 13 1 9 2
13 3 15 13 7 1 9 2 15 4 13 1 9 2
38 7 16 1 9 1 9 12 9 15 13 3 1 12 9 2 1 9 1 0 9 15 3 15 13 1 12 9 2 16 1 9 13 9 7 1 12 9 2
26 3 9 7 9 2 15 13 2 15 13 1 9 2 3 9 1 0 9 15 13 3 1 9 1 9 2
2 0 9
23 7 16 1 9 9 1 0 9 9 13 3 12 9 2 14 1 9 9 15 13 12 9 2
10 9 1 12 9 13 1 1 12 9 2
5 9 2 9 2 9
29 1 0 9 1 9 1 9 1 9 1 9 1 0 0 9 2 0 9 7 0 9 2 1 0 9 6 15 13 2
17 0 9 4 13 2 9 15 13 2 14 7 1 0 9 9 13 2
17 1 9 1 9 13 7 9 1 9 1 9 7 9 1 0 9 2
19 1 12 9 1 9 0 1 9 1 9 1 9 9 3 13 3 12 9 2
9 9 13 9 1 9 1 9 15 2
22 0 9 9 14 6 13 0 13 3 0 9 1 9 2 9 2 9 2 9 7 9 2
28 1 0 15 0 9 9 4 13 14 13 7 9 1 9 2 9 2 9 1 9 2 9 2 0 9 2 9 2
12 0 9 1 15 13 7 15 13 3 0 9 2
15 7 15 13 3 2 1 1 0 9 13 3 1 12 9 2
6 9 15 13 1 0 9
10 9 13 9 15 1 0 9 7 0 11
19 1 0 12 9 9 1 9 1 0 7 0 9 15 4 13 1 0 9 2
15 9 13 0 0 9 2 11 11 2 2 0 1 9 11 2
11 9 13 9 2 1 15 13 3 0 9 2
17 3 12 9 1 0 12 0 9 13 2 16 11 13 9 1 15 2
10 1 12 9 9 13 1 9 1 9 2
15 3 12 9 13 10 2 15 13 2 16 9 13 0 9 2
11 3 12 9 13 2 16 9 13 1 9 2
19 1 9 1 9 12 9 6 4 13 14 9 14 15 13 1 0 15 9 2
21 1 12 9 0 9 2 15 13 14 13 9 2 13 14 6 13 1 0 15 9 2
9 13 9 1 9 1 9 15 1 11
12 15 4 13 1 12 9 1 9 2 11 2 2
5 9 13 1 9 2
9 1 0 9 11 13 3 0 9 2
8 15 13 9 1 0 0 11 2
14 13 15 2 16 13 9 1 0 9 1 11 7 11 2
14 9 2 11 2 13 9 1 0 9 2 11 11 2 2
12 1 11 2 11 11 3 13 0 9 1 9 2
18 9 13 0 9 2 9 1 11 2 7 0 9 2 9 1 11 11 2
13 9 13 0 9 7 9 1 11 3 2 13 11 2
17 9 13 1 9 1 9 12 1 9 2 0 9 2 1 12 9 2
5 0 7 9 13 2
22 9 4 13 1 9 1 0 0 9 1 9 2 11 11 2 7 0 9 2 11 2 2
10 9 1 0 0 9 13 0 11 11 2
4 6 4 13 9
6 13 9 1 9 1 9
24 10 9 1 9 1 9 1 9 14 4 13 1 9 1 0 0 9 2 13 9 15 11 11 2
12 1 0 9 0 15 9 13 1 0 0 9 2
9 14 2 15 13 14 4 15 13 2
21 3 0 9 3 13 7 0 9 1 9 1 9 7 9 1 0 9 1 0 9 2
8 0 3 13 14 13 1 9 2
13 3 1 0 15 9 9 13 3 7 1 0 9 2
20 0 9 1 15 13 2 16 3 12 0 9 1 0 13 9 1 9 1 11 2
23 1 15 3 3 0 9 14 13 0 2 0 7 0 1 9 2 16 13 9 1 0 9 2
30 3 0 1 10 9 13 11 11 2 11 2 2 11 11 2 0 2 2 11 11 2 11 2 2 11 11 2 11 2 2
30 11 3 13 0 9 1 9 9 1 0 9 2 0 1 0 9 2 16 6 15 13 2 13 14 13 2 9 15 2 2
8 1 9 15 13 7 11 11 2
23 9 1 9 2 15 13 9 2 1 9 2 9 2 2 13 3 0 2 7 3 9 13 2
5 13 15 0 9 2
5 13 7 0 9 2
14 15 15 13 2 13 15 1 9 7 13 14 15 13 2
9 16 15 13 9 2 14 15 13 9
22 0 9 3 13 9 1 0 9 1 11 11 11 1 11 2 3 13 14 13 0 9 2
7 3 9 13 12 12 9 2
25 9 7 9 3 14 13 9 1 9 1 0 9 2 3 16 13 9 1 9 1 9 2 13 9 2
12 0 9 0 9 4 13 9 1 12 9 9 2
19 1 12 9 4 13 7 9 1 9 7 9 1 9 2 13 3 1 9 2
26 0 9 13 9 14 13 0 9 2 16 15 14 13 9 1 0 9 2 13 9 1 9 1 0 9 2
9 9 4 13 3 1 9 11 11 2
4 13 9 1 9
20 9 1 9 1 0 9 2 11 2 11 11 4 13 7 13 3 2 13 11 2
18 9 1 12 0 9 1 11 1 0 9 3 14 4 13 1 0 9 2
14 15 13 9 1 0 11 11 2 15 13 1 11 3 2
5 9 1 11 3 0
8 10 9 13 1 9 1 0 9
16 3 0 13 9 1 9 1 11 2 13 1 0 9 1 9 2
29 9 1 0 9 2 0 11 2 4 13 0 9 1 9 1 9 2 1 9 1 0 9 11 2 15 13 3 3 2
5 9 13 1 11 2
17 1 12 9 3 9 1 9 6 4 13 3 0 2 13 0 9 2
14 9 3 13 2 16 9 6 15 13 7 9 14 13 2
14 7 3 0 9 7 9 1 9 13 9 1 0 9 2
14 1 0 0 9 14 15 13 1 3 0 9 1 9 2
19 0 9 13 0 12 9 1 0 9 7 12 9 1 11 1 9 7 9 2
5 13 9 11 2 11
14 0 9 11 2 11 4 13 3 1 9 1 0 9 2
24 9 13 1 0 9 1 0 9 1 9 2 11 11 2 2 11 2 7 2 11 2 2 11 2
13 1 1 9 3 9 13 0 15 9 1 11 9 2
13 9 1 9 7 9 1 9 1 9 13 1 3 2
10 0 9 1 9 1 9 13 0 9 2
14 1 0 9 3 13 9 1 9 1 9 1 0 9 2
22 9 1 10 9 13 0 7 13 14 15 13 1 9 1 0 0 9 1 9 2 9 2
10 9 13 14 15 13 7 1 0 9 2
16 1 12 9 9 15 13 11 2 16 15 13 3 1 0 9 2
15 1 9 9 13 14 15 13 1 12 9 1 9 1 9 2
12 1 12 9 13 9 1 9 1 9 1 9 2
13 1 9 15 13 14 13 0 1 9 1 0 9 2
7 9 1 11 1 0 9 2
8 12 9 1 9 1 12 9 2
11 12 9 7 12 9 1 9 1 12 9 2
11 12 9 7 12 9 1 9 1 12 9 2
5 1 12 12 9 2
12 12 9 7 12 9 1 9 1 12 12 9 2
4 9 3 13 3
13 9 1 0 9 13 1 9 1 12 9 1 9 2
9 13 9 1 9 1 10 9 1 11
32 0 0 9 1 9 1 9 1 15 2 3 7 0 9 1 9 1 11 2 13 1 9 1 0 9 2 13 1 9 1 9 2
11 9 1 11 3 14 13 3 1 0 9 2
18 9 15 1 0 9 1 9 1 11 4 13 1 9 3 1 0 9 2
17 1 9 13 11 2 11 2 11 2 11 2 11 2 11 7 11 2
17 13 15 0 9 1 9 1 0 9 1 0 9 7 9 1 15 2
11 9 4 13 1 0 1 9 9 1 9 2
13 1 9 1 9 14 15 13 0 9 1 0 9 2
15 1 15 14 13 7 9 11 0 2 13 9 1 0 9 2
10 9 13 15 14 13 12 9 1 9 2
8 0 15 9 14 13 11 0 2
14 15 3 13 14 13 11 11 1 9 2 9 11 2 2
15 1 9 1 9 15 13 9 1 11 11 1 9 0 9 2
21 9 11 14 15 13 11 11 2 13 3 0 9 1 11 9 11 11 7 0 9 2
15 9 15 13 1 9 1 9 11 0 1 9 1 0 11 2
17 9 13 9 1 9 7 9 1 9 1 0 9 1 9 1 11 2
18 1 12 12 9 4 13 14 13 0 9 1 3 1 9 2 11 2 2
15 14 15 13 0 9 1 9 2 13 3 3 1 12 9 2
12 9 15 4 13 14 1 9 1 11 1 9 2
17 0 0 9 14 15 4 13 3 2 13 14 13 3 9 7 9 2
12 9 1 1 9 13 11 3 1 14 15 13 2
12 9 13 0 2 3 1 9 13 2 11 2 2
11 9 7 0 9 3 6 13 9 1 9 2
11 3 1 12 9 1 0 9 9 13 11 2
14 0 1 15 3 13 0 9 2 15 15 13 1 9 2
14 1 16 13 0 1 0 9 2 15 6 13 0 9 2
16 6 1 9 1 0 9 2 11 2 3 1 12 9 9 13 2
8 3 1 9 13 2 11 2 2
5 9 13 1 9 2
27 1 0 9 2 15 15 13 2 9 1 9 13 2 7 14 13 9 1 9 1 0 9 15 13 0 9 2
18 1 9 15 15 13 7 9 2 7 9 3 15 13 14 13 1 3 2
13 9 2 9 7 9 13 1 9 1 0 0 9 2
13 11 4 13 1 12 9 1 9 1 9 7 9 2
18 0 11 11 7 0 11 11 13 9 1 9 1 0 15 9 11 11 2
22 1 9 9 13 0 9 2 11 2 1 0 9 2 7 9 1 0 9 15 13 9 2
20 9 1 9 1 2 11 2 11 11 4 13 9 1 1 13 9 1 0 9 2
18 0 9 2 16 9 13 9 15 2 1 15 13 1 0 9 2 13 2
14 11 4 13 1 9 1 9 9 1 1 13 9 15 2
7 9 13 9 1 0 9 2
20 9 1 0 0 9 1 2 11 2 7 9 11 11 3 3 15 13 1 9 2
23 15 4 13 1 0 9 1 9 15 2 7 13 14 13 10 1 9 2 11 11 2 11 2
5 9 1 9 13 11
11 1 12 9 9 13 0 9 1 0 9 2
14 1 12 9 4 13 9 1 9 1 11 9 11 11 2
25 12 0 9 4 13 1 0 9 2 12 9 13 9 7 9 1 12 0 9 1 0 9 11 11 2
11 1 9 4 13 7 9 1 9 11 11 2
33 1 0 9 1 0 9 0 9 4 13 12 9 2 11 11 2 11 2 11 11 2 11 2 11 11 2 11 7 11 11 2 11 2
12 4 13 7 13 0 9 11 11 7 11 11 2
25 15 13 0 9 2 1 1 13 9 1 12 9 2 9 2 0 9 2 9 2 9 7 9 15 2
23 0 0 9 1 9 1 0 9 13 9 1 9 1 11 1 0 9 1 9 1 0 9 2
7 0 11 13 9 1 0 9
11 9 13 1 9 1 0 9 9 11 11 2
7 9 15 13 9 11 11 2
24 11 13 9 15 1 9 0 9 7 1 0 9 1 11 2 7 1 9 3 4 13 1 9 2
5 11 13 0 15 9
19 9 1 9 14 13 1 0 9 7 1 12 0 9 2 1 11 7 11 2
11 11 9 12 15 13 9 9 12 1 11 2
19 9 1 9 13 0 9 14 13 9 1 9 1 9 11 11 1 0 9 2
21 1 16 15 6 13 2 9 13 2 16 0 0 9 14 13 9 1 9 1 9 2
12 1 9 9 13 9 1 11 1 12 9 9 2
10 11 14 15 13 1 2 11 12 2 2
13 1 9 9 1 9 9 15 13 3 9 12 9 2
17 1 1 13 9 1 0 3 15 13 2 16 15 13 12 12 9 2
24 1 11 13 2 0 11 11 2 0 1 15 9 2 9 1 0 9 2 9 7 9 1 9 2
10 9 13 2 16 9 13 0 1 11 2
13 13 15 2 16 3 4 13 9 3 1 12 9 2
17 1 9 0 9 11 13 9 1 9 11 2 15 13 9 1 11 2
4 0 9 13 11
11 9 14 13 0 1 0 9 7 0 9 2
11 9 3 9 13 9 3 1 12 9 9 2
12 1 0 9 1 0 9 13 9 1 9 11 2
12 0 9 11 11 13 2 16 0 9 13 9 2
23 9 9 1 12 9 1 11 13 1 9 2 7 9 15 13 1 9 2 1 14 13 9 2
14 13 15 2 16 0 9 13 9 1 9 1 12 9 2
16 9 3 0 13 9 15 2 7 3 9 4 13 9 1 9 2
5 9 1 9 13 11
18 9 1 9 14 15 13 9 1 9 1 9 7 0 9 13 0 9 2
13 1 0 9 9 13 9 2 9 2 9 2 9 2
4 13 7 0 2
13 7 14 14 15 13 3 9 2 3 13 1 11 2
12 10 9 3 13 12 9 2 0 1 0 9 2
8 14 13 14 14 13 9 15 2
5 9 2 10 0 9
23 0 9 1 0 9 13 10 0 9 2 7 9 7 0 0 9 15 13 1 3 0 9 2
21 9 7 9 13 3 9 2 0 9 1 15 3 3 13 14 4 13 1 0 9 2
7 1 9 3 6 13 9 2
7 1 9 1 15 13 9 2
8 15 15 13 7 1 11 11 2
10 6 13 14 15 13 9 1 0 9 2
12 1 15 3 13 1 9 1 9 1 0 9 2
19 0 15 9 1 9 3 3 14 4 13 14 13 14 0 0 9 1 11 2
21 11 6 13 7 9 1 11 2 1 15 11 11 15 13 9 1 2 9 12 2 2
23 7 2 16 1 9 15 13 3 3 9 1 0 9 2 3 1 3 0 9 15 13 3 2
24 3 0 9 15 13 1 0 9 1 9 1 2 11 2 2 1 15 0 9 3 3 13 9 2
22 9 1 9 7 9 2 11 2 14 6 15 13 2 7 14 9 13 3 3 1 9 2
9 7 2 0 9 15 13 1 9 2
9 7 0 9 7 3 3 0 9 2
8 7 0 12 9 9 0 9 2
7 9 3 13 2 3 13 2
8 15 13 1 9 3 1 9 2
8 7 3 15 13 1 0 9 2
10 1 15 1 9 4 13 3 3 9 2
11 9 2 9 7 9 2 15 13 1 0 9
17 7 16 13 9 1 9 7 9 2 9 13 3 0 7 0 9 2
7 9 1 0 9 3 13 2
18 1 0 9 1 0 9 2 0 9 2 13 9 11 14 15 13 11 2
10 7 15 13 14 13 0 9 1 9 2
13 1 0 15 9 10 9 13 7 9 1 0 9 2
20 3 3 14 13 3 0 9 1 0 9 2 15 4 13 9 15 1 0 9 2
20 3 7 14 13 3 1 9 2 9 1 0 9 3 13 14 13 1 10 9 2
24 13 15 2 13 9 2 16 0 9 13 9 1 9 1 9 15 1 9 1 11 1 0 9 2
9 13 15 14 13 15 14 13 9 2
12 11 11 2 0 9 1 2 11 7 9 2 2
5 9 13 9 1 9
20 2 3 0 2 16 15 13 14 13 1 9 15 1 10 9 2 15 13 9 2
15 3 1 10 9 6 15 13 10 2 15 14 13 10 9 2
10 9 13 3 0 9 2 9 1 9 2
13 0 13 3 9 2 15 6 15 13 2 6 13 2
5 0 9 13 0 2
14 1 0 9 13 3 3 0 9 2 15 3 15 13 2
17 3 3 6 13 14 2 16 3 9 1 15 15 3 3 13 3 2
33 13 15 15 2 16 0 9 1 9 1 9 13 0 1 11 2 3 9 1 0 9 1 9 15 13 2 15 6 13 0 1 15 2
9 3 9 1 9 6 4 13 3 2
20 2 16 13 14 13 0 2 10 15 9 2 13 2 16 15 14 13 3 3 2
37 2 1 16 13 9 1 0 0 9 2 1 9 1 9 0 9 11 11 1 9 1 0 9 13 3 2 16 0 15 9 6 13 1 0 12 9 2
8 7 9 15 6 13 1 9 2
8 3 3 9 6 13 1 9 2
15 1 15 0 9 1 0 9 13 0 2 0 1 0 9 2
16 0 9 13 9 2 3 13 9 1 9 14 13 0 0 9 2
27 3 13 14 15 13 9 10 2 15 13 9 1 9 2 14 13 0 9 1 9 1 0 15 9 1 9 2
10 7 2 13 14 15 13 9 1 9 2
17 15 14 13 9 3 9 1 0 9 14 15 13 1 9 1 9 2
22 1 9 1 12 9 9 7 9 1 12 9 9 1 10 9 15 13 3 1 12 9 2
16 16 10 0 9 13 10 9 2 0 9 3 14 13 1 9 2
19 3 13 14 15 13 12 9 9 1 9 2 1 14 15 13 9 1 11 2
11 11 11 2 12 9 2 2 9 2 11 2
7 2 13 9 14 15 13 2
6 13 3 14 15 13 2
11 11 11 2 12 9 2 2 9 2 11 2
10 2 1 0 9 15 13 1 3 9 2
17 3 2 3 0 2 4 13 9 2 7 9 3 15 13 1 3 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
11 3 14 13 16 13 0 12 9 1 9 2
11 11 11 2 12 9 2 2 0 2 11 2
10 2 14 0 9 14 13 0 7 0 2
17 1 0 9 15 13 14 15 13 9 2 3 3 15 13 3 3 2
12 9 11 2 12 9 2 2 0 9 2 11 2
12 2 13 3 9 2 9 1 11 7 0 9 2
11 13 15 9 15 14 13 3 1 10 9 2
11 11 11 2 12 9 2 2 9 2 11 2
10 2 13 14 13 1 11 1 10 9 2
11 1 15 14 13 14 13 3 0 15 9 2
11 11 11 2 12 9 2 2 9 2 11 2
4 0 9 15 13
20 0 9 11 11 15 13 1 10 9 11 11 2 13 0 9 2 11 2 3 2
20 15 13 1 12 9 0 1 11 2 15 3 4 13 1 11 7 4 13 9 2
6 9 1 9 11 11 11
28 0 9 2 15 4 13 1 9 1 0 9 1 9 2 13 0 9 2 13 9 7 13 9 2 13 11 11 2
4 9 13 0 9
19 1 12 9 4 13 1 0 9 1 0 0 9 11 1 9 2 13 11 2
41 15 15 13 3 0 2 3 0 2 1 0 9 1 9 7 9 2 1 9 7 9 2 1 9 7 9 1 0 9 2 9 2 9 14 15 13 2 13 2 13 2
18 15 15 13 1 0 0 9 2 9 2 9 2 9 2 9 2 9 2
30 15 15 13 1 0 9 7 9 1 0 9 1 0 9 7 0 9 2 1 0 15 0 9 2 1 0 9 1 9 2
15 9 2 3 1 0 9 2 9 2 3 1 9 1 9 2
28 0 9 3 13 2 0 9 7 0 9 1 10 2 0 9 2 7 1 9 10 9 1 9 0 13 3 0 2
23 16 13 9 1 12 9 2 11 13 9 1 9 2 3 1 9 9 1 9 1 0 9 2
16 9 1 9 13 7 0 9 1 0 9 7 0 9 11 11 2
12 9 6 13 9 1 10 9 2 9 13 9 2
4 9 13 0 2
6 13 15 9 1 0 9
22 0 1 12 9 9 1 9 2 11 2 1 11 11 1 0 9 4 13 1 0 9 2
21 15 15 4 13 1 0 9 7 15 4 13 1 0 0 9 1 9 2 14 13 2
23 9 2 15 15 13 1 9 1 2 0 9 2 1 11 2 15 13 1 10 1 0 9 2
34 0 9 13 7 9 1 9 12 2 3 11 11 2 11 11 7 11 11 13 14 13 0 9 1 0 0 9 1 2 9 1 9 2 2
10 0 13 2 16 15 6 13 0 9 2
8 13 15 7 9 1 0 9 2
37 0 9 15 13 3 7 13 2 16 4 13 12 9 2 15 13 1 0 9 7 0 0 9 2 7 0 0 9 2 1 9 2 13 10 0 9 2
18 1 3 0 9 1 15 13 7 0 0 9 1 0 2 11 12 2 2
29 9 13 1 9 1 11 11 0 9 1 0 9 7 9 1 2 11 2 2 0 0 9 1 0 9 1 0 9 2
16 14 9 14 13 15 7 0 15 9 1 10 9 1 0 9 2
7 11 13 9 1 2 11 2
34 1 9 1 9 1 11 1 11 14 9 14 13 7 1 9 1 11 11 2 11 2 2 15 3 14 13 1 9 1 2 11 11 2 2
37 1 0 9 15 13 2 16 1 0 9 1 11 1 9 14 15 13 7 0 9 1 2 11 2 11 11 2 15 4 13 0 9 1 2 0 2 2
14 0 9 1 11 13 3 1 9 1 11 1 12 9 2
15 9 1 2 11 2 13 9 15 1 0 9 1 9 3 2
9 9 15 13 1 0 9 7 13 9
10 1 9 1 9 13 3 3 12 9 2
8 11 13 14 13 1 2 11 2
18 9 1 2 11 2 11 11 13 14 13 1 2 11 2 2 11 2 2
15 10 9 11 4 13 1 11 1 9 7 13 3 12 9 2
12 9 15 1 2 11 2 13 1 9 1 9 2
13 1 0 9 13 7 9 1 2 11 2 11 11 2
20 9 2 15 13 0 15 9 1 9 1 0 9 2 4 13 9 3 12 9 2
14 9 15 13 9 2 7 9 1 11 6 13 3 0 2
6 14 15 13 1 0 9
13 15 13 0 9 1 2 11 2 1 9 1 9 2
10 16 6 13 3 2 6 13 14 13 9
3 13 15 9
31 13 14 15 9 1 0 9 2 14 13 0 7 0 15 1 9 15 9 2 16 9 9 13 0 7 6 13 1 0 9 2
60 0 2 0 2 0 7 3 0 2 9 14 15 13 1 0 15 9 2 1 9 7 9 15 2 15 13 14 13 0 9 2 9 2 9 7 9 2 2 7 14 15 13 1 0 9 1 9 2 1 0 9 7 0 9 7 1 0 15 9 2
16 13 15 1 10 9 7 6 13 9 15 2 16 13 1 15 2
36 1 9 0 9 3 14 13 9 1 9 15 1 0 15 9 2 9 14 13 9 1 9 2 9 7 9 2 7 3 14 15 13 9 1 9 2
23 0 2 0 1 0 9 7 9 1 0 2 0 7 0 2 15 14 13 9 15 1 12 2
14 3 9 15 1 9 7 9 1 10 9 13 3 0 2
18 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
2 0 9
18 9 1 9 11 13 9 1 0 9 7 9 1 0 9 1 10 9 2
7 9 11 11 13 0 0 9
11 11 11 13 9 1 0 9 1 12 9 2
29 1 15 1 9 15 13 11 11 2 12 9 2 2 11 11 2 12 9 2 2 11 11 2 11 11 7 11 11 2
7 9 1 9 13 9 1 11
23 0 0 9 1 11 1 9 1 0 9 13 9 1 0 9 1 9 11 2 13 0 9 2
32 2 9 2 1 9 1 9 11 11 7 9 11 14 13 1 9 1 9 7 9 1 9 2 3 9 7 9 13 14 15 13 2
13 9 13 9 1 12 0 9 7 13 9 12 12 2
8 9 13 14 13 0 9 1 9
17 0 9 13 1 9 11 11 2 15 13 1 12 9 7 12 9 2
15 1 9 15 1 9 11 11 4 13 1 0 9 0 9 2
11 9 1 11 11 15 13 1 9 12 9 2
6 9 13 9 1 0 9
17 11 11 7 11 11 14 15 13 9 1 11 2 11 2 11 2 2
6 9 13 14 15 13 9
14 12 0 9 9 11 11 13 0 0 9 1 9 11 2
29 1 0 9 1 0 9 0 9 15 13 1 2 11 11 2 7 13 1 9 15 2 7 1 9 6 15 13 9 2
17 12 9 3 1 11 12 9 13 1 9 1 9 11 1 0 9 2
14 9 3 9 9 13 1 9 1 9 3 1 10 9 2
31 1 0 9 9 11 11 2 15 13 1 9 2 9 2 2 13 2 16 15 13 1 9 2 1 1 4 13 1 0 9 2
20 9 3 13 3 3 2 12 9 1 9 1 9 11 13 1 0 9 1 9 2
9 1 9 13 9 2 1 0 9 2
18 0 9 13 2 16 9 13 1 9 7 15 13 1 0 9 1 9 2
11 0 0 9 11 2 11 4 13 10 9 2
23 1 16 9 4 13 2 1 9 15 6 15 13 2 3 9 6 13 2 16 9 13 3 2
25 14 13 0 9 1 15 2 13 9 1 11 11 11 1 11 9 1 9 1 9 1 0 0 9 2
14 1 15 13 11 2 11 2 11 7 9 2 11 2 2
20 9 1 0 0 9 2 15 14 13 9 1 9 2 11 2 2 13 0 9 2
22 9 13 0 9 2 0 9 1 0 9 2 7 13 9 2 15 13 14 13 0 9 2
22 13 15 9 2 10 9 3 15 13 1 9 2 14 15 13 1 9 1 9 1 9 2
11 9 1 0 9 13 0 9 1 11 3 2
10 9 13 2 16 9 13 1 9 11 2
11 1 0 9 13 7 9 1 9 1 9 2
6 14 13 9 1 0 9
8 3 9 13 9 1 9 1 9
25 9 2 11 2 13 0 9 1 0 9 7 9 1 9 2 11 2 2 15 13 1 9 0 9 2
31 1 0 9 9 4 13 1 11 2 16 9 1 9 1 9 4 13 1 0 9 1 11 2 11 2 11 2 11 7 11 2
6 0 9 13 0 15 9
17 9 1 9 1 0 9 13 9 7 0 9 2 13 2 11 2 2
18 3 13 3 2 3 0 1 9 1 15 13 1 0 9 2 13 9 2
9 14 13 14 2 9 2 1 0 9
15 2 9 2 6 4 13 1 15 2 3 9 13 3 9 2
21 10 1 0 9 13 0 9 1 11 2 13 9 2 3 0 1 9 1 0 9 2
27 10 12 9 4 13 1 11 7 13 3 3 14 15 13 1 0 2 1 1 13 1 0 9 2 13 9 2
4 15 13 0 2
27 9 2 1 15 15 13 9 1 9 2 15 13 0 9 7 9 3 13 9 7 9 15 2 9 12 2 2
5 9 13 9 1 9
19 7 14 1 0 9 15 13 1 9 14 13 9 7 9 1 0 0 9 2
15 9 13 9 12 7 0 0 9 1 9 1 9 7 9 2
19 10 9 3 14 13 0 9 1 1 14 13 0 9 1 12 3 0 9 2
24 0 1 9 1 9 9 2 9 2 9 2 9 2 9 2 9 7 9 3 15 13 0 9 2
13 7 3 10 9 13 0 15 9 1 9 7 9 2
26 0 9 1 9 1 9 13 2 16 1 12 9 1 9 13 9 2 7 14 2 9 14 13 9 15 2
19 3 13 3 14 15 13 2 16 9 9 14 13 7 13 3 12 9 3 2
22 3 9 7 1 10 9 14 15 13 3 1 9 2 15 7 3 15 13 3 0 9 2
14 13 15 9 1 9 1 0 9 7 0 9 11 11 2
15 1 12 9 15 13 9 15 1 9 1 0 9 1 9 2
3 3 3 2
12 1 10 9 0 9 13 0 9 1 0 9 2
7 2 11 2 14 13 3 9
8 0 9 1 9 14 13 1 9
14 9 1 2 11 2 14 13 1 9 2 13 0 9 2
24 3 15 13 9 1 9 7 3 0 9 2 1 15 15 13 1 9 0 9 2 9 7 9 2
16 0 9 1 0 9 13 9 1 9 1 9 1 9 1 9 2
17 10 9 15 13 7 1 0 9 1 0 9 1 9 1 0 9 2
17 1 9 13 9 7 1 9 2 7 1 0 9 2 7 1 9 2
38 13 14 9 2 16 9 4 13 1 9 1 9 2 3 1 0 9 4 13 2 16 3 9 4 13 0 9 1 0 9 2 9 1 2 11 9 2 2
19 1 15 15 13 7 0 7 0 15 9 1 0 9 7 1 9 1 9 2
40 7 16 6 15 13 9 2 0 2 11 11 11 11 11 2 13 14 13 10 9 2 0 9 7 0 9 1 12 9 9 1 0 1 9 9 1 9 12 9 2
8 7 3 3 9 13 1 3 2
3 13 15 2
13 0 9 1 0 9 4 13 14 13 9 15 11 2
15 15 4 13 1 9 1 0 9 1 11 1 0 9 9 2
15 15 4 13 1 9 1 0 9 1 11 1 0 9 9 2
17 15 13 1 9 2 9 2 9 2 7 13 9 1 9 12 9 2
25 9 13 12 9 1 9 2 9 2 9 7 9 1 9 1 11 7 11 9 2 3 13 10 9 2
4 3 1 9 12
4 9 13 1 9
15 0 11 11 1 9 11 13 1 9 9 1 9 1 11 2
15 1 0 9 11 9 1 9 13 0 9 2 15 13 9 2
5 9 13 0 9 2
10 9 3 13 2 16 4 13 0 9 2
6 13 15 1 9 1 9
10 11 4 13 0 9 1 9 1 9 2
24 15 13 9 1 0 9 2 11 11 2 1 9 1 11 11 2 0 1 9 2 11 11 2 2
8 1 15 4 13 11 7 11 2
27 1 11 15 13 2 16 9 1 0 9 7 9 7 1 11 15 13 1 9 1 9 1 9 7 1 9 2
5 11 13 0 9 2
11 9 1 11 7 11 4 13 1 0 9 2
9 1 9 13 7 0 2 7 9 2
22 9 11 15 13 9 2 15 15 13 1 0 0 9 2 7 13 3 14 15 13 9 2
22 3 3 13 1 0 9 11 11 7 0 9 11 11 2 15 13 9 1 0 0 9 2
8 11 13 9 1 0 0 9 2
8 9 1 9 3 13 1 11 2
16 0 13 9 15 1 9 1 0 9 1 9 1 11 11 11 2
11 3 9 15 13 1 9 1 9 1 11 2
18 0 9 9 9 1 9 11 11 3 13 12 9 1 9 1 0 9 2
6 9 1 11 13 9 2
14 0 9 14 13 14 13 9 1 11 7 0 0 9 2
18 1 11 3 9 1 0 15 9 13 9 1 9 1 9 15 1 11 2
24 0 0 9 13 9 1 0 9 11 11 2 15 13 1 15 1 9 1 9 1 9 1 11 2
10 0 9 1 9 3 3 6 15 13 2
22 13 14 9 0 1 0 9 11 11 2 15 13 0 9 2 11 2 1 9 1 9 2
3 3 3 2
7 9 1 9 14 13 11 2
12 3 7 3 15 13 1 9 3 1 9 15 2
7 9 13 0 2 13 9 2
16 7 3 9 1 9 1 9 7 0 6 13 0 1 0 9 2
15 1 0 9 1 9 9 15 4 13 1 0 0 0 9 2
14 1 0 9 1 12 9 3 15 13 9 1 3 9 2
7 9 1 12 9 13 0 2
13 1 0 9 3 6 13 0 1 0 9 1 9 2
20 1 0 9 3 11 13 2 16 0 9 1 9 14 13 9 1 9 1 9 2
8 3 9 13 9 14 15 13 2
12 0 9 15 14 13 13 11 0 14 13 3 2
12 13 9 14 15 13 9 2 15 6 4 13 2
10 1 0 9 9 13 9 1 0 9 2
16 12 1 9 2 15 14 4 13 2 13 15 14 13 0 9 2
19 9 11 13 2 16 9 13 0 2 1 14 13 2 7 14 13 10 9 2
14 0 9 2 0 9 3 1 9 7 9 1 3 9 2
21 0 9 15 13 7 1 9 3 1 9 9 11 11 11 2 13 9 15 11 11 2
7 9 4 13 1 0 9 2
15 9 13 1 9 1 9 2 1 1 9 11 13 1 9 2
11 13 15 2 16 15 13 0 1 0 9 2
26 11 13 9 1 9 11 1 9 1 9 1 9 2 9 1 9 2 1 9 9 2 7 9 15 13 2
17 7 12 9 13 14 13 14 1 0 9 14 4 13 9 1 9 2
27 0 9 9 1 0 9 4 13 1 9 1 9 2 11 2 1 0 9 11 7 11 11 2 13 3 9 2
19 1 15 9 4 13 1 9 2 15 13 1 9 1 9 7 13 1 9 2
26 1 9 1 9 6 4 13 1 9 1 9 14 4 4 13 9 1 9 9 2 15 4 13 0 9 2
10 15 13 0 9 1 9 2 13 9 2
4 13 9 1 9
22 0 9 13 9 2 11 2 1 9 1 11 1 12 9 1 9 2 13 11 2 11 2
5 13 9 7 0 2
4 9 4 13 2
10 9 13 1 9 2 11 7 11 2 2
22 12 9 13 9 1 9 1 9 1 11 11 1 0 9 1 9 1 9 2 13 11 2
10 3 15 13 0 9 1 9 1 9 2
24 1 9 0 13 2 16 6 13 0 9 2 7 13 9 1 0 0 0 9 2 11 11 2 2
13 15 13 2 16 13 14 13 10 0 9 1 11 2
6 9 4 13 1 11 2
16 0 0 9 13 14 13 0 9 1 9 1 9 1 0 9 2
23 1 12 9 1 9 7 3 9 1 0 11 13 9 11 11 2 1 14 15 13 1 9 2
4 9 13 12 9
9 11 13 1 9 1 9 1 9 2
4 9 4 13 2
24 0 11 11 2 0 1 9 1 0 11 11 1 0 9 2 6 4 13 9 2 13 1 9 2
6 11 13 1 0 9 2
17 3 3 14 4 13 1 9 1 0 9 1 0 9 1 12 9 2
8 11 11 13 9 1 0 9 2
19 15 13 14 13 1 9 15 1 9 2 0 11 2 7 3 6 15 13 2
16 12 9 9 2 9 7 9 13 9 1 0 9 7 0 9 2
12 9 13 9 1 0 9 1 9 7 15 13 2
29 1 0 9 9 13 1 9 1 9 1 9 2 11 2 1 9 11 7 13 1 9 1 0 9 1 0 9 3 2
19 1 0 9 1 9 9 12 1 9 1 9 1 11 13 9 1 0 9 2
15 15 6 13 9 7 3 13 2 6 4 13 14 4 13 2
15 1 15 13 7 9 15 1 9 2 1 15 3 4 13 2
7 9 13 1 0 0 9 2
6 3 4 13 1 9 2
24 1 12 9 1 0 9 4 13 1 9 1 9 2 7 3 16 6 15 13 2 9 15 13 2
10 0 0 9 1 9 13 9 1 11 2
12 1 14 4 13 2 9 4 13 3 7 3 2
14 13 4 2 16 9 4 13 12 9 1 9 1 9 2
9 1 11 0 9 15 13 1 9 2
28 1 12 9 13 9 1 0 15 9 2 7 1 10 9 2 1 15 13 9 2 9 13 14 15 13 0 9 2
4 11 14 15 13
3 9 1 15
8 13 9 2 0 1 0 9 2
28 12 15 13 1 11 2 1 1 4 13 1 9 1 0 0 9 11 11 1 9 1 9 1 9 2 0 9 2
18 9 13 14 13 9 7 9 1 9 2 3 15 13 9 1 9 11 2
5 13 11 1 11 2
9 9 1 9 13 0 9 1 9 2
13 3 9 13 2 16 11 4 13 1 0 0 9 2
14 1 9 15 1 0 9 9 3 4 13 9 1 9 2
16 0 13 7 9 2 16 4 13 9 2 0 1 9 1 9 2
16 11 13 9 3 2 7 9 15 4 13 1 0 9 1 9 2
18 11 13 0 15 9 1 11 2 0 1 9 1 0 15 9 1 9 2
23 1 12 9 11 11 13 7 0 9 2 7 10 9 6 13 0 14 15 13 1 9 15 2
30 3 3 1 9 9 1 11 12 9 4 13 1 9 1 12 9 2 7 6 15 13 9 2 15 14 15 13 1 9 2
22 9 13 1 0 9 2 0 0 9 1 11 11 7 12 9 9 1 9 1 11 11 2
4 9 3 13 2
14 1 12 9 13 1 9 1 9 2 13 11 7 11 2
31 1 1 13 1 0 9 2 0 9 14 13 12 9 2 1 15 14 15 13 3 1 9 2 13 9 1 9 2 11 2 2
12 9 1 2 9 2 9 0 2 13 1 0 9
29 0 0 9 3 15 13 9 3 1 9 1 0 9 1 12 9 2 11 2 11 2 11 7 0 9 2 11 2 2
13 3 2 3 11 13 3 9 7 9 1 0 9 2
23 3 3 3 1 9 1 11 11 6 13 14 15 13 2 16 9 13 12 9 9 0 9 2
24 3 1 15 13 14 13 3 1 9 2 16 13 2 16 15 13 1 0 9 3 1 9 15 2
17 13 15 1 0 9 1 0 9 14 13 9 11 11 7 11 11 2
7 15 14 13 14 13 11 2
15 1 9 1 9 13 7 11 11 2 3 15 1 0 11 2
29 16 13 0 0 9 3 13 3 7 1 0 9 1 11 11 0 9 0 9 14 13 9 1 9 11 0 1 9 2
10 9 2 15 13 14 13 14 4 13 2
4 11 11 2 9
6 11 14 13 9 1 11
17 9 13 9 1 0 9 2 13 15 1 0 0 9 7 0 9 2
9 7 15 13 9 7 9 1 9 2
12 2 0 9 13 2 16 9 1 0 15 13 2
11 15 13 14 13 9 3 1 3 0 9 2
12 9 1 9 1 9 13 9 1 9 1 0 2
15 14 7 1 10 0 9 3 4 13 1 0 1 11 9 2
15 11 6 13 1 9 1 9 2 3 16 13 3 0 9 2
18 9 6 4 13 1 11 7 15 6 13 14 13 10 9 1 9 15 2
17 7 9 11 2 0 1 0 9 2 1 9 6 15 13 1 15 2
5 13 9 1 9 2
20 7 3 13 9 1 9 2 10 9 6 13 14 15 13 14 13 1 10 9 2
18 11 3 13 9 1 0 9 2 13 15 1 0 0 9 7 0 9 2
9 7 15 13 9 7 9 1 9 2
14 3 13 3 2 16 10 9 13 1 0 9 1 11 2
18 7 15 13 2 16 0 9 1 9 1 9 13 9 1 2 11 2 2
6 15 13 0 0 9 2
22 2 9 2 15 9 4 13 1 0 9 2 13 9 1 9 11 2 16 3 13 15 2
6 15 3 6 13 9 2
12 14 15 13 9 2 0 1 11 2 11 11 2
8 0 9 2 1 0 0 9 2
8 2 3 9 1 11 15 13 2
14 3 15 13 2 16 0 9 14 15 13 9 14 2 2
9 14 14 6 13 3 0 0 9 2
15 3 14 13 9 7 1 0 9 14 15 13 9 7 9 2
21 10 2 15 13 14 15 13 1 11 2 13 3 3 7 15 13 1 0 9 9 2
7 15 13 9 1 0 9 2
7 3 7 0 9 3 13 2
11 3 15 3 13 9 1 9 15 1 11 2
17 7 3 1 9 13 0 9 2 1 14 15 13 1 0 15 9 2
14 1 10 9 0 13 9 2 15 13 3 12 9 9 2
21 9 1 15 2 16 10 0 9 13 14 15 13 2 11 14 4 13 1 12 9 2
14 3 15 13 2 16 11 7 11 13 0 15 0 9 2
14 7 16 13 2 1 0 9 14 13 7 1 0 9 2
7 15 13 0 1 15 9 2
12 16 13 2 0 9 15 13 2 13 3 11 2
7 3 13 9 7 13 9 2
5 9 11 15 13 9
18 9 1 9 13 2 16 9 4 13 1 11 2 0 11 2 13 11 2
8 9 6 13 0 2 13 9 2
13 0 9 13 2 16 4 13 0 9 1 0 9 2
10 9 11 15 13 3 7 6 13 9 2
9 3 15 15 13 1 9 15 11 2
15 1 15 15 3 4 13 1 9 1 9 1 9 1 11 2
12 0 9 1 0 9 11 0 3 4 13 9 2
30 1 0 9 1 9 1 9 1 9 15 15 13 0 9 2 7 1 0 9 1 9 1 9 15 13 9 2 13 11 2
19 11 13 9 1 9 0 9 14 13 11 1 0 9 1 9 1 9 11 2
19 0 0 9 1 9 1 0 0 9 1 11 15 13 1 9 2 13 11 2
14 0 4 13 1 9 1 0 9 1 11 1 0 9 2
19 15 13 2 16 1 11 10 9 15 13 12 9 1 9 2 3 1 9 2
6 12 9 1 9 1 9
27 1 9 11 2 15 13 1 9 1 9 1 11 1 0 9 2 13 0 9 1 9 2 11 11 11 2 2
18 3 0 13 9 1 0 1 0 9 2 9 1 11 1 11 11 11 2
14 1 15 13 13 14 13 7 9 1 0 9 1 11 2
37 9 1 9 1 0 2 15 15 13 1 0 15 9 1 9 1 11 11 1 0 9 1 11 2 14 15 13 7 13 1 9 1 0 9 1 9 2
33 6 15 13 14 14 9 11 11 2 0 9 11 11 7 0 9 1 0 0 9 11 11 14 13 1 0 9 2 0 9 1 9 2
20 9 1 0 9 1 11 1 0 9 1 15 14 4 13 1 9 1 0 9 2
37 1 3 10 9 13 9 1 0 1 0 9 7 0 2 13 0 9 1 11 2 0 9 2 11 2 11 2 11 11 7 0 12 0 7 0 9 2
11 15 13 9 1 9 7 9 2 13 11 2
11 0 9 2 15 4 13 9 2 13 11 2
2 1 9
7 11 11 13 11 12 1 9
15 3 15 13 1 9 1 9 1 9 2 9 1 15 2 2
2 11 11
5 11 13 9 1 11
16 14 13 7 0 15 9 1 11 2 13 9 1 11 11 11 2
9 15 13 7 9 1 0 0 9 2
2 11 11
3 9 1 9
26 0 1 0 15 9 2 15 15 13 1 9 2 13 15 1 0 9 11 7 13 14 13 9 7 9 2
9 9 15 13 1 9 1 0 9 2
19 1 9 1 0 9 0 9 1 9 3 13 1 9 1 9 1 9 15 2
10 1 9 9 7 9 13 9 1 0 2
9 9 4 13 1 3 9 1 9 2
31 9 1 11 2 11 2 7 9 1 9 11 11 13 9 15 1 0 9 1 11 1 0 9 1 0 0 9 2 11 2 2
13 9 1 0 9 2 0 1 9 2 13 7 1 0
5 9 15 13 1 9
44 9 11 15 13 1 2 0 0 9 1 0 0 9 2 0 9 1 0 9 9 7 9 2 12 9 2 12 9 2 0 9 2 9 1 0 9 7 3 12 9 1 0 9 2
35 3 16 0 9 13 9 1 9 1 9 2 15 4 13 1 0 1 9 9 1 0 9 7 0 9 2 0 15 9 13 1 9 1 9 2
14 9 15 4 13 1 0 9 2 7 1 9 13 9 2
6 13 4 1 0 9 2
9 3 13 14 15 13 9 1 11 2
22 9 11 15 4 13 1 10 0 9 2 3 13 9 2 13 1 9 7 13 9 9 2
8 0 9 2 0 15 9 11 2
12 11 15 13 1 12 1 0 0 9 1 9 2
8 2 9 13 1 9 1 12 2
7 11 7 11 14 13 3 2
11 11 2 13 15 2 13 14 13 1 9 2
16 2 9 4 13 1 11 2 1 14 13 9 1 9 7 9 2
4 2 3 3 2
10 2 1 15 15 13 14 13 1 9 2
4 2 9 14 2
9 9 13 0 9 1 9 7 9 2
4 3 1 9 2
12 2 9 7 9 6 13 14 15 13 1 9 2
6 13 0 9 1 9 2
7 9 11 13 0 15 9 2
9 10 0 9 13 1 9 1 9 2
13 0 0 9 15 13 2 13 0 15 9 2 13 2
4 11 13 9 2
14 0 9 13 1 0 2 0 9 1 9 7 0 9 2
10 2 13 2 16 9 15 13 1 9 2
20 9 2 11 7 11 15 13 3 1 9 2 0 1 0 9 7 0 1 9 2
7 13 0 9 1 0 9 2
11 11 13 3 0 7 13 0 9 1 9 2
18 9 13 1 9 2 3 3 13 3 3 2 7 15 13 1 0 9 2
25 11 15 13 7 1 0 9 15 13 1 9 15 2 15 3 13 2 13 9 15 7 15 13 3 2
14 9 13 1 9 1 9 7 9 2 9 15 3 13 2
13 2 13 15 2 2 13 7 11 15 13 1 9 2
7 9 11 13 9 1 9 2
15 1 2 6 2 11 2 11 11 13 9 1 0 9 1 9
9 9 13 9 1 0 7 0 9 2
19 1 9 13 0 9 1 0 9 1 0 3 9 2 1 10 9 7 9 2
9 11 11 13 9 1 12 0 9 2
30 0 9 10 9 2 9 1 9 2 4 13 1 0 9 1 12 9 1 9 1 2 11 9 2 7 9 2 9 2 2
5 15 2 10 2 3
5 13 9 1 0 9
17 13 15 1 9 9 1 9 1 9 15 11 7 9 1 10 9 2
12 11 13 9 2 0 7 0 9 1 0 9 2
8 15 13 14 13 1 0 11 2
12 2 9 1 9 2 13 9 1 2 11 2 2
8 9 1 0 13 1 11 11 2
15 9 13 3 9 13 3 14 4 13 1 0 9 1 9 2
19 13 4 10 9 1 9 7 0 15 9 3 1 0 2 3 7 1 13 2
9 11 11 13 9 1 0 9 1 11
19 1 0 15 9 2 1 9 2 11 11 13 9 1 0 9 1 0 9 2
11 2 1 9 2 13 9 1 2 11 2 2
6 9 13 1 11 11 2
6 13 9 14 13 11 2
18 9 1 9 1 0 9 14 13 14 4 13 3 1 9 1 0 9 2
15 1 9 1 0 9 7 1 0 9 15 13 1 12 9 2
19 9 4 13 1 0 11 1 9 0 9 7 4 13 1 0 9 1 9 2
8 11 13 1 2 9 2 1 11
16 9 1 11 11 11 13 1 9 1 2 0 2 1 11 11 2
12 1 9 1 9 11 13 14 13 14 10 9 2
23 3 0 9 1 11 11 11 14 13 9 2 15 14 13 1 9 1 2 11 2 1 9 2
18 9 11 7 3 6 13 1 11 2 1 14 15 13 1 9 1 11 2
21 2 11 2 2 15 6 13 1 0 9 1 0 0 9 1 11 2 13 1 11 2
20 1 16 13 1 3 9 2 2 11 2 13 1 9 11 7 13 3 1 9 2
11 9 11 13 1 0 9 12 9 1 9 2
12 11 13 1 0 9 2 7 1 9 11 13 2
12 9 13 9 15 2 1 16 4 13 9 11 2
27 11 11 7 11 11 13 1 0 9 1 0 9 1 9 1 0 9 1 12 9 1 11 2 11 2 3 2
27 11 11 7 11 11 13 1 0 9 1 0 9 1 9 1 0 9 1 12 9 1 11 2 11 2 3 2
31 1 0 15 9 1 9 7 1 9 11 13 12 9 1 9 7 13 0 1 12 9 1 9 11 2 11 2 1 0 9 2
20 3 3 15 15 13 1 11 2 7 15 13 2 16 6 13 0 2 13 0 9
15 1 9 11 11 14 4 13 1 9 1 11 1 0 9 2
14 0 9 1 10 9 4 13 1 9 1 9 1 9 2
11 1 11 11 15 13 11 11 7 11 11 2
7 15 13 0 9 1 15 2
8 2 15 15 13 1 12 9 2
22 1 9 1 0 9 15 13 3 3 7 1 3 3 13 9 1 0 0 9 1 9 2
5 9 15 13 0 2
12 1 15 15 13 12 3 0 1 10 9 9 2
8 13 14 13 9 1 10 9 2
7 2 3 14 13 3 3 2
12 2 3 4 13 2 16 9 6 13 1 15 2
7 9 13 1 2 11 2 2
12 2 15 15 13 0 9 1 9 1 10 9 2
8 3 15 15 13 1 11 11 2
10 3 13 9 2 3 15 14 6 13 2
15 9 1 11 2 1 11 2 3 1 11 2 3 13 9 2
6 13 3 0 15 9 2
14 3 3 14 13 2 16 1 15 11 11 6 13 0 2
5 13 14 13 9 2
13 13 9 2 13 9 2 13 15 9 14 15 13 2
7 9 13 1 2 11 2 2
17 15 15 4 13 9 2 16 14 13 1 0 9 2 7 15 13 2
11 16 6 13 0 7 0 2 15 6 13 2
15 13 14 13 9 2 7 16 15 13 2 15 13 1 9 2
17 7 15 13 9 12 1 9 1 9 7 13 14 13 10 15 9 2
13 3 12 9 2 1 0 9 11 6 13 0 9 2
16 2 13 14 9 1 11 11 2 16 0 9 13 14 15 13 2
4 2 6 13 2
7 2 14 15 13 3 0 2
8 9 6 4 13 14 13 9 2
18 9 13 14 13 0 2 0 2 0 2 1 15 9 6 13 1 9 2
17 2 0 9 1 9 3 13 1 9 1 11 2 11 7 0 9 2
5 3 15 13 9 2
38 10 2 16 15 13 1 0 9 2 15 13 14 15 13 2 3 10 12 9 15 13 0 0 9 2 15 13 0 9 1 15 14 6 13 9 1 9 2
24 1 9 9 13 1 0 0 9 7 3 9 1 11 15 13 2 1 14 13 14 13 0 9 2
11 1 10 9 3 13 1 9 1 0 9 2
16 14 15 13 0 9 2 15 1 9 1 11 6 13 14 13 2
10 2 3 3 13 9 1 0 0 9 2
17 2 1 10 9 14 13 9 1 0 9 7 3 14 13 0 9 2
9 1 9 1 9 14 13 15 0 2
28 7 12 13 3 0 1 9 1 9 1 11 7 13 2 16 3 9 14 15 13 1 10 9 1 0 15 9 2
20 9 1 11 7 11 1 9 11 12 7 12 13 0 9 1 11 2 13 9 2
28 1 9 1 0 9 3 0 9 13 2 16 1 10 9 13 1 9 1 12 0 9 1 9 11 12 7 12 2
15 13 2 16 15 13 10 0 9 1 11 2 13 0 9 2
17 15 13 2 16 0 9 13 3 0 9 1 10 9 1 10 9 2
20 1 9 1 0 9 1 0 9 1 9 1 9 2 10 9 13 3 0 9 2
26 9 1 9 1 9 1 0 9 13 1 0 9 3 1 10 9 2 3 7 1 10 9 2 13 9 2
17 9 13 2 16 1 11 3 4 13 9 1 0 9 1 10 9 2
18 3 15 4 13 3 10 9 1 0 9 1 0 9 2 13 11 11 2
24 11 13 2 16 13 0 0 9 1 9 15 7 3 13 9 1 11 11 1 0 9 1 11 2
11 9 11 13 0 9 0 1 9 1 9 2
7 9 14 13 1 0 9 2
10 9 11 11 13 9 1 0 0 9 2
38 0 0 9 13 9 15 2 16 0 0 0 9 7 0 0 9 1 10 9 14 13 3 0 9 1 10 0 9 2 3 1 0 9 15 13 0 9 2
30 13 2 3 3 13 1 0 9 1 0 9 2 9 2 15 3 4 15 13 1 9 15 2 15 13 15 2 13 9 2
12 1 9 1 15 15 13 7 1 9 1 9 2
20 10 9 1 2 0 2 9 0 13 12 9 7 12 9 1 9 1 0 9 2
17 9 13 1 9 2 11 2 9 1 9 2 0 1 2 11 2 2
51 10 9 15 13 1 9 2 0 9 1 2 11 2 7 2 0 9 2 2 9 1 2 11 2 2 2 11 9 2 7 2 11 2 2 9 1 2 11 2 7 2 9 11 2 7 9 1 2 11 2 2
7 0 1 9 13 11 11 2
15 9 11 13 3 9 1 0 15 9 1 9 1 0 9 2
17 9 13 9 1 9 7 9 1 2 0 2 3 9 0 9 2 2
20 0 1 0 9 1 9 1 9 13 0 9 1 9 1 9 2 13 11 11 2
10 9 1 9 2 11 11 2 2 0 9
10 9 1 9 1 9 14 4 13 3 2
11 9 13 1 9 1 9 1 0 0 9 2
13 3 1 9 11 4 13 9 1 9 1 0 9 2
22 1 9 1 0 9 1 9 1 0 9 2 0 9 15 13 3 12 9 1 12 9 2
23 9 11 11 13 12 0 9 1 9 1 0 15 9 1 9 1 0 9 1 9 1 9 2
21 15 13 0 15 1 9 1 9 1 0 0 9 1 9 7 9 1 9 1 11 2
38 1 9 2 1 0 9 1 9 2 1 9 3 13 0 9 2 15 13 1 9 2 9 13 2 16 13 15 14 13 3 0 1 10 0 9 1 11 2
10 1 15 9 4 15 13 14 13 9 2
14 7 0 9 3 13 10 7 0 0 9 2 13 9 2
15 3 15 13 0 9 1 9 1 12 9 2 13 11 11 2
38 1 9 0 9 1 0 0 9 1 9 1 9 1 11 1 0 9 11 11 13 2 16 4 15 13 2 16 9 1 11 3 13 14 13 1 10 9 2
21 1 9 1 10 9 13 0 9 14 13 9 1 9 1 10 9 2 13 15 9 2
14 9 7 0 9 13 0 0 9 1 0 0 9 1 11
13 0 9 13 9 1 9 1 9 0 9 1 9 2
19 1 9 1 9 15 1 0 9 9 13 0 0 9 1 9 1 0 9 2
18 1 15 11 11 13 0 9 7 0 9 1 9 7 13 9 1 11 2
26 9 1 9 1 0 9 13 7 9 1 0 9 9 11 11 2 9 1 9 11 11 7 0 0 9 2
15 0 9 2 15 13 1 0 0 9 2 13 10 0 9 2
16 1 0 9 14 13 2 0 9 2 16 6 13 10 9 2 2
28 3 3 15 14 13 9 1 0 9 1 0 9 2 7 1 15 14 13 7 9 1 11 7 14 13 1 9 2
25 1 9 2 0 1 0 9 1 9 2 4 13 9 1 9 9 2 0 1 11 11 7 11 11 2
44 0 9 1 9 1 9 13 1 10 9 14 4 13 10 9 1 9 2 9 2 7 9 1 9 1 15 2 1 14 13 9 3 14 15 13 7 3 14 15 13 9 1 9 2
28 9 1 9 2 11 11 7 11 11 13 9 2 9 2 2 16 13 12 0 9 2 0 1 0 9 1 9 2
58 1 0 9 1 9 4 13 0 9 1 9 7 9 15 1 9 7 9 1 9 2 1 0 9 9 4 13 1 9 1 0 9 2 0 9 13 9 1 9 1 9 1 9 1 9 7 9 2 0 9 13 9 1 9 1 0 9 2
9 2 10 0 9 4 13 1 9 2
16 16 10 9 4 13 1 9 2 15 4 13 9 1 9 2 2
14 0 0 9 13 0 9 2 10 9 4 13 1 9 2
27 3 4 15 13 2 1 14 13 9 1 0 9 1 9 12 9 1 9 1 0 9 11 11 2 13 9 2
23 9 2 15 13 9 1 0 9 1 9 1 0 9 2 13 1 0 9 1 9 11 11 2
14 9 11 11 13 14 13 9 1 9 1 9 1 0 9
15 9 11 11 13 14 13 9 1 9 1 9 1 0 9 2
14 15 13 15 3 1 9 1 9 1 9 15 1 11 2
20 9 13 9 2 16 10 9 1 0 0 9 15 13 1 9 15 14 13 11 2
7 13 4 11 1 12 9 2
22 1 9 14 13 9 1 11 9 13 2 16 0 4 13 14 13 9 1 0 15 9 2
14 1 3 9 13 9 2 9 2 9 2 1 10 9 2
8 3 16 2 14 14 6 13 0
42 1 10 9 0 9 2 1 15 9 9 13 9 1 10 9 2 13 2 16 0 0 9 3 4 13 9 7 1 0 9 2 7 1 0 9 2 13 13 7 1 0 9
11 9 1 11 7 11 13 9 1 9 1 9
22 9 1 9 7 10 9 1 9 13 3 9 1 11 7 1 11 11 11 7 11 11 2
20 0 0 9 13 1 0 9 1 11 7 13 1 9 1 9 1 0 0 9 2
11 15 13 9 11 1 9 1 9 1 9 2
28 1 0 9 9 1 11 1 0 9 4 13 2 16 11 13 0 9 2 15 13 14 15 13 1 9 7 9 2
14 1 9 15 15 13 0 9 1 10 2 15 15 13 2
9 15 13 10 9 1 11 1 9 2
13 11 13 10 0 9 1 0 9 2 13 0 9 2
11 15 13 9 1 9 7 1 9 1 9 11
41 1 9 15 1 9 1 9 1 0 0 9 2 0 1 9 1 11 1 9 1 9 7 9 1 0 0 9 2 9 11 11 13 1 9 1 11 1 9 1 9 2
11 13 4 2 16 9 1 11 6 13 0 2
37 13 9 1 11 7 1 3 12 0 9 2 15 13 0 0 9 2 9 2 0 1 0 9 1 10 9 1 9 1 9 1 0 9 2 13 9 2
26 15 13 0 1 9 1 0 0 9 1 9 1 11 9 2 1 15 11 4 13 2 9 1 9 2 2
12 1 9 11 13 1 10 9 2 13 9 11 2
7 1 11 9 6 13 0 2
9 9 13 0 9 2 0 1 0 9
8 15 13 2 16 13 3 9 2
14 15 13 9 1 0 9 2 1 14 15 13 0 9 2
19 15 13 15 13 9 2 7 15 13 1 9 2 1 14 6 13 1 9 2
12 1 0 9 14 13 2 16 9 13 0 9 2
12 3 9 1 11 13 3 14 15 13 1 9 2
31 3 13 9 1 9 1 0 9 9 1 9 1 9 1 11 15 13 1 0 9 1 9 2 13 0 9 1 11 11 11 2
14 1 11 2 0 11 2 13 10 3 9 14 4 13 2
7 15 15 13 15 6 15 13
4 11 13 9 11
2 11 11
36 11 11 1 0 9 13 2 16 3 4 15 13 2 0 9 1 9 9 1 9 2 7 15 13 1 12 9 2 1 16 11 13 1 12 9 2
13 9 15 13 14 13 7 9 1 9 2 12 9 2
25 9 15 13 1 0 9 1 0 9 2 15 3 6 4 4 13 1 9 1 9 1 9 1 9 2
11 3 13 2 16 15 4 13 1 9 1 11
16 1 0 9 3 9 13 9 2 16 13 14 13 9 1 9 2
8 0 9 4 13 7 0 9 2
25 0 9 1 11 11 11 7 9 1 11 11 11 13 12 9 0 9 7 4 13 1 9 3 9 2
23 11 11 4 13 1 0 9 1 0 0 9 2 1 9 9 15 13 1 1 12 9 9 2
21 9 1 11 11 13 1 3 0 9 1 9 2 0 9 13 1 12 9 1 9 2
4 9 13 1 11
12 13 15 9 2 13 9 7 3 3 15 13 2
8 15 15 13 10 9 1 9 2
11 1 15 1 9 13 14 15 13 0 9 2
4 3 13 9 2
3 3 13 2
16 16 6 15 15 13 15 2 0 15 6 13 7 15 13 1 9
3 9 7 9
3 9 7 9
15 0 9 9 13 1 9 2 0 1 9 2 3 1 9 2
6 15 13 3 1 11 2
8 11 11 3 13 9 1 9 15
13 11 11 13 14 0 15 0 9 1 9 1 9 2
11 9 1 9 13 3 12 0 9 1 9 2
18 9 13 0 15 0 9 1 9 1 9 9 11 1 9 2 11 2 2
10 3 9 15 13 1 0 9 11 11 2
26 1 14 15 13 1 9 15 2 0 11 13 9 1 0 9 2 13 9 7 13 9 2 13 0 9 2
13 0 11 11 15 13 1 11 0 9 1 0 9 2
7 9 7 9 13 12 9 2
13 9 13 2 16 15 14 15 13 0 9 1 9 2
8 13 15 11 11 7 11 11 2
22 11 11 3 13 3 2 7 3 14 10 9 14 15 13 14 13 9 15 2 13 11 2
10 1 9 4 13 12 9 1 0 9 2
29 9 13 2 16 1 0 9 1 11 11 15 13 11 11 2 11 2 11 11 2 11 11 2 11 11 7 11 11 2
15 1 0 12 0 9 13 11 11 1 0 9 7 11 11 2
9 11 13 12 0 9 1 2 11 2
17 15 13 9 1 0 9 1 9 0 9 7 13 2 16 3 13 15
29 0 9 2 15 4 4 13 1 9 1 9 11 7 1 9 1 0 9 2 1 15 13 11 11 2 6 4 13 2
17 1 15 7 9 1 11 7 1 0 9 1 11 6 4 13 9 2
11 6 4 13 0 9 11 14 13 10 9 2
14 13 9 1 10 9 1 10 9 2 14 14 4 13 9
15 9 2 15 13 9 2 13 11 11 2 0 9 1 11 2
4 13 0 9 2
12 13 15 0 9 1 0 9 7 9 1 0 9
40 1 15 3 15 4 2 13 9 1 9 1 10 9 2 7 1 0 9 2 16 4 13 9 1 11 6 4 13 10 9 14 13 9 1 9 1 10 9 2 2
12 3 7 11 6 13 14 13 0 9 1 9 2
14 15 13 1 15 14 13 9 7 13 1 9 1 11 2
14 9 2 15 9 1 11 15 13 13 0 2 13 15 2
5 3 3 15 13 2
39 3 13 15 2 16 10 9 1 11 13 1 0 9 1 0 9 2 15 15 13 1 9 2 16 13 14 15 13 2 1 14 6 15 13 7 14 15 13 9
10 1 15 13 14 13 9 1 10 9 2
7 7 0 9 1 15 13 2
44 13 4 2 9 11 11 2 9 1 0 9 1 0 9 1 11 2 9 11 11 7 9 11 11 2 0 9 1 0 9 2 3 7 9 11 11 2 9 1 9 1 0 9 2
11 1 11 1 9 1 0 9 13 3 3 2
7 15 13 3 0 1 9 2
37 3 13 7 1 10 9 13 0 9 1 11 2 13 0 9 2 15 15 13 0 9 1 0 9 7 6 15 13 3 14 13 14 15 13 1 10 9
14 6 4 13 0 9 1 10 0 9 1 9 1 11 2
4 13 0 9 2
8 13 4 11 2 11 11 2 2
13 1 0 9 13 0 9 1 0 0 9 1 11 2
10 1 9 1 9 4 13 1 0 9 2
11 11 13 9 1 11 2 11 2 11 7 11
13 0 9 14 15 13 3 12 9 1 9 1 9 2
22 1 9 1 9 11 11 9 2 0 1 9 2 13 0 1 10 9 7 13 14 13 2
8 11 3 15 13 3 3 9 2
18 1 9 1 11 9 13 14 13 11 2 11 7 9 1 11 7 0 2
23 3 15 13 2 16 14 15 13 3 9 1 9 2 3 14 15 13 3 10 0 9 1 9
22 1 15 0 9 2 15 15 13 3 13 9 1 0 7 0 9 1 0 9 1 11 2
17 16 4 13 9 1 9 1 11 2 0 15 9 13 14 15 13 9
20 9 1 11 11 11 13 2 16 0 9 1 9 13 9 1 9 9 11 11 2
8 9 1 9 1 9 15 4 13
18 9 1 9 11 7 11 15 13 7 1 9 7 13 14 13 1 15 2
4 9 2 11 11
25 0 9 1 0 9 11 1 9 1 12 9 1 11 7 9 1 0 9 15 13 3 1 9 3 2
28 1 15 1 9 1 1 12 9 15 13 0 0 9 1 9 1 9 2 15 15 13 1 11 2 11 7 11 2
14 1 11 13 0 9 2 0 1 9 1 9 7 9 2
40 1 0 9 9 13 2 16 9 15 13 2 7 13 9 3 2 9 1 0 9 2 9 1 0 9 1 11 7 9 1 9 1 0 9 1 9 1 0 9 2
20 1 11 13 14 13 10 9 1 0 1 9 9 2 3 10 9 6 4 13 2
17 9 15 1 9 2 11 11 2 3 6 13 9 1 9 1 9 2
21 9 1 9 1 11 2 0 1 0 9 1 0 9 2 14 15 13 2 13 11 2
31 3 3 3 6 15 13 14 9 1 11 14 15 13 1 9 1 9 1 0 9 7 14 15 13 1 9 1 9 1 9 2
9 9 3 3 14 13 9 1 0 9
70 1 0 9 4 4 13 12 9 2 9 1 11 1 9 1 11 11 11 2 15 4 13 1 0 15 9 1 11 2 9 1 9 2 0 9 7 9 2 1 11 11 11 2 15 13 1 0 15 9 1 11 2 9 1 9 1 11 11 11 2 15 15 13 1 11 7 0 0 9 2
15 10 9 13 1 9 1 15 1 0 9 1 9 1 9 2
6 9 13 3 1 9 2
26 1 9 15 13 1 9 2 16 7 12 9 13 9 7 3 3 13 2 16 9 13 14 13 1 15 2
9 3 14 15 13 14 13 1 15 2
22 1 15 15 6 13 2 16 3 3 13 9 1 9 1 9 0 9 13 9 1 11 2
6 13 0 9 1 9 2
23 0 9 1 9 2 15 14 15 13 7 13 3 2 15 13 3 1 0 9 1 0 9 2
12 1 9 1 0 0 9 13 9 11 0 9 2
28 1 11 0 0 9 7 10 9 6 13 14 4 13 1 9 1 9 1 9 2 9 2 9 2 9 7 9 2
13 0 9 13 14 13 3 9 1 11 1 10 9 2
10 1 12 9 9 11 11 13 10 9 2
4 9 2 11 11
3 13 9 2
4 14 13 9 15
10 15 4 13 9 1 0 9 0 9 2
11 1 0 9 11 4 13 3 1 10 9 2
27 1 0 9 2 6 13 3 14 15 13 13 9 1 11 1 9 1 9 1 11 1 9 1 11 7 11 2
2 15 2
2 11 2
8 7 1 0 15 15 13 9 2
14 2 13 4 9 1 9 1 9 0 1 9 1 11 2
6 1 10 9 13 9 2
14 2 1 10 9 4 13 9 7 4 13 14 13 9 2
11 2 15 4 13 9 2 13 9 1 15 2
10 2 1 10 9 13 15 14 15 13 2
5 7 15 13 9 2
18 9 1 9 1 11 13 1 9 2 1 14 6 13 0 15 9 9 2
5 3 4 13 9 2
8 2 3 15 15 13 3 13 2
6 15 13 3 1 9 2
10 15 13 9 2 15 15 13 1 9 2
9 10 9 15 4 15 13 10 9 2
11 2 11 11 4 13 1 9 1 0 9 2
8 2 15 6 13 14 13 9 2
16 2 15 13 2 16 4 13 3 0 2 1 14 13 2 2 2
5 3 13 1 11 2
6 13 9 1 9 3 2
19 9 1 12 9 15 15 13 7 13 3 1 12 9 14 13 1 0 9 2
5 15 13 0 9 2
14 1 12 9 15 13 7 1 12 9 15 13 1 9 2
5 13 15 9 9 2
9 3 10 2 13 2 15 15 13 2
7 15 14 13 16 13 0 2
5 7 15 15 13 2
6 9 1 15 13 0 2
5 3 13 1 9 2
10 13 2 16 15 6 13 1 15 14 2
6 13 15 9 1 9 2
4 0 13 3 2
14 3 15 14 15 13 14 13 3 4 13 9 1 11 2
6 2 1 15 4 13 2
4 15 14 13 2
11 3 1 0 9 14 13 12 9 1 11 2
5 15 13 0 9 2
13 13 12 9 2 15 3 13 14 15 13 1 15 2
13 3 13 15 2 13 16 7 3 0 9 13 3 2
14 13 0 9 1 2 10 9 2 2 9 1 9 1 9
3 1 15 13
12 15 13 0 2 3 13 2 3 14 15 13 2
20 2 0 9 1 0 9 2 0 9 1 11 7 0 9 1 9 1 2 11 2
3 7 3 2
4 2 9 1 9
2 2 9
6 2 9 1 9 1 9
5 2 13 1 11 11
6 0 9 13 1 9 2
3 3 3 2
12 14 13 2 3 13 3 2 0 9 1 9 2
17 3 2 14 13 9 1 0 9 2 3 0 9 13 1 0 9 2
10 7 7 1 0 9 3 13 0 9 2
23 7 9 15 13 1 0 9 2 3 0 9 13 0 1 0 9 2 15 15 13 1 9 2
3 7 14 2
6 14 11 13 0 9 2
10 7 0 9 6 4 13 1 9 2 2
11 6 13 1 12 9 2 1 0 9 13 2
7 3 10 13 9 1 9 2
4 1 0 9 2
2 6 2
8 3 0 9 13 9 1 9 2
3 9 1 9
6 6 9 2 7 9 2
26 6 13 3 14 15 13 9 2 9 2 1 9 1 0 9 2 13 3 9 1 0 9 9 11 11 2
6 6 9 2 7 9 2
12 13 9 1 9 2 15 13 9 7 0 9 2
3 11 13 9
18 11 4 13 9 15 1 9 1 0 9 1 9 7 9 1 0 9 2
12 9 13 0 0 9 1 9 2 11 11 2 2
11 1 11 3 15 13 1 0 0 0 9 2
18 1 0 9 1 0 9 15 13 9 1 9 2 9 2 9 7 9 2
12 9 14 4 13 1 0 9 7 1 0 9 2
14 0 9 1 0 9 14 15 13 1 0 9 1 11 2
28 3 9 4 13 1 9 11 0 1 0 9 2 15 13 14 15 13 2 7 13 14 13 9 1 11 1 9 2
29 1 9 1 12 0 9 4 13 1 9 9 2 15 13 1 9 1 9 1 9 1 11 12 1 9 2 11 2 2
7 13 9 14 15 13 3 2
20 13 9 15 1 11 2 7 7 6 13 2 16 9 14 15 13 14 13 1 9
13 0 9 14 15 4 13 1 0 9 2 13 11 2
36 0 9 2 9 1 12 9 2 13 2 16 9 15 4 13 9 1 9 1 2 11 2 2 15 15 13 1 0 0 9 1 9 1 0 9 2
5 0 9 13 1 11
14 0 11 13 0 9 1 9 7 13 1 9 1 9 2
16 9 13 9 1 10 1 9 7 13 1 9 1 3 0 9 2
12 1 9 1 0 9 2 9 1 9 13 3 2
10 9 15 13 1 0 9 11 7 11 2
15 2 11 11 11 11 2 13 1 11 7 14 13 1 11 2
7 2 11 2 13 2 11 2
8 11 13 1 15 1 12 9 2
14 13 14 13 1 0 9 7 3 13 14 15 13 0 9
13 11 11 13 14 13 9 1 11 2 1 14 13 9
21 9 1 11 11 11 13 9 1 0 9 9 1 0 15 9 1 0 9 11 11 2
17 9 1 9 6 13 1 9 15 2 3 3 9 13 9 1 11 2
11 0 15 9 1 11 13 1 0 0 9 2
22 1 0 9 1 9 7 9 1 11 4 13 0 9 2 15 13 1 0 9 1 11 2
6 12 9 13 1 11 2
21 9 14 13 1 12 2 16 9 15 1 9 2 9 11 2 13 1 9 1 9 2
12 13 4 9 1 9 2 1 15 15 13 9 2
9 7 1 0 9 6 4 13 9 2
16 3 1 0 15 13 9 9 12 1 0 9 2 9 11 11 2
16 15 3 13 14 13 1 9 2 3 1 0 9 14 13 9 2
11 11 13 14 13 9 1 9 1 0 9 2
14 11 7 11 13 9 2 3 16 9 6 13 1 9 15
24 1 9 1 11 3 13 9 11 11 7 11 11 2 15 14 13 1 9 1 9 2 11 2 2
7 11 13 0 9 1 11 2
16 12 4 13 1 9 2 11 2 7 1 3 13 9 7 9 2
12 11 15 13 3 7 6 13 14 13 0 9 2
8 9 12 1 9 13 1 0 9
15 15 13 1 0 9 1 9 1 9 2 11 2 1 11 2
10 15 13 3 3 7 6 15 13 10 9
8 0 9 13 9 1 2 11 2
12 9 1 11 13 9 7 15 13 2 13 11 11
18 0 9 11 11 13 0 9 2 15 13 1 9 1 2 11 2 11 2
10 1 9 1 0 9 9 3 13 9 2
14 1 2 11 2 9 15 13 1 0 9 2 15 4 13
12 13 15 3 1 10 0 9 7 9 1 9 2
23 1 10 9 9 1 11 11 2 15 3 13 7 13 0 9 2 4 13 1 3 0 9 2
10 0 9 11 13 0 9 1 11 11 2
14 15 15 13 0 9 7 15 13 1 0 9 11 11 2
20 1 2 11 2 11 13 9 2 16 14 13 0 0 9 1 0 9 1 11 2
5 9 1 9 1 11
27 9 1 2 11 2 11 11 15 13 0 9 1 2 0 2 11 11 14 15 13 1 9 1 2 11 2 2
2 11 11
11 0 9 1 0 9 4 13 1 11 3 2
23 9 1 11 4 13 1 9 1 0 9 11 11 2 16 9 14 13 1 9 1 0 9 2
9 10 9 13 3 9 1 0 9 2
28 1 0 9 13 3 2 16 0 9 1 11 3 13 1 0 9 1 0 9 1 2 11 2 7 2 11 2 2
7 1 15 13 9 1 11 2
25 1 9 1 9 14 13 11 11 2 11 11 2 11 11 7 11 11 2 15 15 13 1 0 9 2
18 3 9 13 7 1 0 0 9 1 10 0 9 1 9 1 0 9 2
13 1 3 3 13 0 9 1 9 2 11 11 2 2
15 0 9 1 9 1 2 11 2 1 2 0 9 2 1 9
2 11 11
11 0 0 9 11 13 9 1 0 15 9 2
22 0 9 1 11 13 14 13 3 0 1 0 9 9 1 9 1 2 11 2 11 11 2
11 3 1 9 11 13 0 12 9 1 9 2
27 3 1 9 2 0 2 13 12 0 9 7 15 13 1 0 9 2 1 15 13 14 13 7 0 15 9 2
30 3 3 1 11 4 13 9 1 9 9 7 9 11 11 14 13 14 13 9 1 9 1 3 0 2 11 2 1 9 2
11 10 1 9 1 11 6 4 13 1 9 2
21 1 0 9 13 3 2 16 9 1 9 1 2 11 2 14 13 1 3 0 9 2
22 13 2 9 2 2 12 9 2 2 9 2 2 12 9 7 2 9 2 2 12 9 2
19 0 14 15 13 9 9 14 13 14 13 15 10 9 1 2 0 9 2 2
18 16 15 13 3 3 0 9 2 13 14 15 13 3 7 1 10 9 2
20 15 15 13 1 9 1 9 1 0 9 7 9 1 9 2 11 2 1 3 2
20 1 9 3 13 0 9 1 9 1 0 0 9 1 11 7 9 1 0 9 2
11 9 14 13 14 13 1 0 2 0 9 2
32 1 11 9 15 13 1 9 2 15 6 13 7 1 9 2 0 1 9 7 9 15 11 11 2 7 1 9 2 0 1 15 2
18 0 9 3 13 1 12 9 9 2 7 3 9 13 1 12 9 9 2
16 1 11 3 13 0 9 14 15 13 0 9 1 9 1 9 2
17 0 9 1 0 9 1 11 11 11 13 9 1 0 9 1 9 2
16 3 9 1 9 7 9 13 0 9 1 9 1 9 1 9 2
15 9 13 9 1 9 2 15 3 4 13 1 9 1 11 2
19 0 9 13 3 9 1 0 9 9 2 1 15 9 13 0 9 7 9 2
5 9 1 9 15 13
1 9
9 9 7 9 14 13 9 1 0 9
13 9 14 13 3 1 11 2 3 3 4 13 9 2
6 9 13 1 9 1 11
23 0 9 2 11 11 11 11 2 4 13 0 9 1 9 14 13 0 9 1 0 0 9 2
17 15 13 14 15 13 1 9 1 9 2 16 13 9 1 9 15 2
19 9 1 0 9 13 12 9 9 2 7 9 1 9 13 1 12 9 9 2
21 16 15 13 9 2 7 14 13 14 13 9 1 11 1 9 1 9 1 12 9 2
1 9
2 11 11
8 0 0 9 13 2 16 13 9
2 11 11
23 15 4 13 1 0 9 7 9 6 4 13 1 14 10 1 9 2 13 9 1 0 9 2
7 9 13 1 12 9 9 2
18 9 15 13 1 9 15 2 7 15 13 9 1 9 1 9 1 11 2
24 13 0 9 2 1 15 3 4 13 2 11 2 2 7 0 9 2 15 15 13 2 13 9 2
1 9
13 16 9 13 9 1 11 2 3 15 3 14 13 2
15 13 2 16 13 14 14 6 13 7 12 9 9 1 11 2
10 6 13 14 13 9 1 9 1 11 2
26 2 11 2 7 11 6 13 14 13 15 1 9 3 12 9 2 1 9 1 2 11 2 2 13 11 2
13 11 1 0 9 15 13 1 9 1 0 0 9 2
7 11 13 9 2 13 11 2
12 1 15 14 13 3 9 1 14 13 0 9 2
10 3 3 12 9 13 14 13 0 9 2
15 2 11 2 13 0 9 7 15 6 13 0 2 13 11 2
1 9
37 6 13 14 13 0 9 1 9 7 9 1 0 9 2 3 16 6 13 9 1 10 9 7 13 9 1 15 2 13 9 1 2 11 2 11 11 2
20 10 9 15 13 9 1 9 2 1 15 15 13 1 12 9 9 2 13 11 2
24 3 1 9 1 0 9 1 9 2 9 14 15 13 7 0 9 2 13 9 1 2 11 2 2
5 11 11 13 1 11
12 9 11 11 13 1 11 2 1 14 13 9 2
16 9 1 2 11 2 11 11 14 13 9 1 9 1 0 9 2
13 1 15 9 3 13 2 3 13 9 1 0 15 9
1 9
9 9 1 0 9 1 0 1 0 9
14 13 9 1 0 9 1 9 1 12 9 1 0 9 2
20 1 9 15 13 1 0 9 1 11 7 13 0 9 1 9 15 1 0 9 2
14 1 9 13 2 16 3 4 15 13 1 15 1 11 2
19 15 14 13 1 9 1 11 2 1 15 9 13 3 2 9 2 3 2 2
16 9 13 12 12 9 2 1 14 15 13 1 9 1 12 9 2
19 2 0 2 7 11 3 13 0 9 1 9 7 3 13 14 13 9 15 2
1 9
28 9 1 11 1 15 11 11 13 3 0 1 9 1 0 9 1 2 11 2 11 11 1 9 1 2 11 2 2
27 3 1 9 15 13 0 9 11 11 1 9 1 11 2 1 14 15 13 1 0 9 1 2 0 2 9 2
26 2 9 11 2 3 14 13 9 1 11 11 1 9 1 9 1 9 9 2 11 2 2 2 11 2 2
26 2 9 11 2 3 14 13 9 1 11 11 1 9 1 9 1 9 9 2 11 2 2 2 11 2 2
18 12 1 12 9 14 4 13 2 7 11 7 11 14 13 14 13 9 2
20 9 11 3 15 13 1 9 2 7 1 9 6 13 14 15 13 1 0 9 2
18 9 1 2 11 2 13 9 7 13 9 15 14 13 9 1 0 9 2
12 13 15 11 7 11 14 6 13 3 0 9 2
11 14 15 13 2 16 3 4 4 13 3 2
9 2 3 14 0 9 13 3 0 2
9 9 3 13 0 9 1 10 9 2
11 14 0 9 14 6 13 0 1 10 9 2
1 9
10 15 13 9 15 1 9 1 9 9 2
14 1 9 1 2 11 2 4 13 14 14 13 0 9 2
18 13 4 14 6 15 13 1 0 9 2 3 3 10 9 14 15 13 3
15 14 13 9 1 9 2 6 13 3 14 15 13 7 1 9
20 9 1 11 11 11 3 15 13 1 9 1 9 2 11 2 2 2 11 2 2
11 15 13 0 1 0 9 1 2 0 2 2
8 13 10 9 14 6 15 13 3
15 11 6 13 14 13 9 1 9 2 3 6 13 1 11 2
13 3 1 0 9 13 9 7 0 9 1 0 0 9
15 11 13 0 9 2 7 1 0 9 2 1 9 13 9 2
21 1 9 1 9 10 9 15 13 12 0 9 2 1 15 13 14 13 15 15 13 2
22 0 9 1 9 4 13 1 9 1 0 9 2 7 1 9 15 13 3 0 7 0 2
12 13 15 3 12 9 1 9 2 11 11 2 2
9 15 6 13 14 13 1 0 9 2
9 15 13 14 13 3 1 0 9 2
11 14 0 9 3 13 1 9 1 9 2 2
6 3 15 4 15 13 2
8 15 6 15 4 13 1 11 2
9 13 9 2 13 9 2 13 9 2
46 3 15 13 10 9 9 14 6 13 14 13 0 9 2 14 13 0 9 2 14 15 13 1 9 2 1 15 13 0 9 2 7 13 9 2 13 9 2 13 9 2 13 9 7 3 2
14 14 3 15 4 4 13 2 1 14 15 13 1 9 2
15 3 15 4 13 1 9 2 3 15 6 13 14 15 13 2
11 6 4 13 1 9 2 15 6 15 13 2
12 9 11 11 13 0 9 1 9 15 11 11 2
13 0 9 4 13 1 9 11 11 2 9 1 9 2
20 9 1 0 9 4 3 13 1 9 2 7 15 15 13 1 0 2 9 2 2
16 13 0 9 1 0 1 9 7 0 9 1 9 13 9 9 2
3 7 14 2
2 13 2
5 1 9 15 13 2
2 13 2
6 10 9 13 10 9 2
14 1 12 9 13 9 1 9 1 9 2 0 9 2 2
4 1 12 4 13
2 11 11
20 3 1 0 9 11 15 13 12 9 2 15 13 9 1 0 9 2 11 2 2
15 1 9 10 9 15 13 1 12 9 2 0 9 7 9 2
30 9 1 9 2 0 9 2 11 11 13 2 16 9 1 0 9 13 0 0 9 1 9 2 7 15 13 9 1 9 2
11 1 0 9 13 9 0 9 1 9 11 2
22 9 13 1 12 9 2 9 2 0 9 7 9 2 9 2 0 0 9 7 0 9 2
1 9
11 15 13 9 2 15 6 13 3 1 11 2
10 0 0 9 1 9 11 11 3 13 2
1 9
6 13 9 1 11 1 9
19 11 13 9 1 9 1 9 9 7 13 2 16 9 13 14 13 9 15 2
6 9 1 9 1 0 9
25 12 9 9 14 13 1 0 9 2 16 0 9 1 9 15 13 2 13 0 9 2 0 1 11 2
19 1 9 3 2 15 13 14 13 9 1 0 9 2 9 13 1 12 9 2
5 9 13 11 1 11
8 0 11 2 0 1 11 11 2
5 13 0 0 9 2
2 11 11
10 9 4 4 13 1 9 12 1 9 2
8 13 4 3 2 7 0 13 2
8 9 4 13 1 0 0 9 2
24 1 0 9 1 9 1 9 15 4 13 0 11 11 2 15 13 1 0 9 1 0 9 12 2
17 11 15 13 1 9 1 0 1 11 9 1 9 9 2 13 9 2
20 15 13 2 16 9 4 13 7 0 15 9 4 4 13 14 15 13 1 9 2
13 1 2 11 2 11 13 2 16 6 4 13 9 2
8 15 13 9 15 1 0 9 2
14 10 9 13 2 16 15 13 0 15 9 1 0 9 2
5 11 13 9 1 9
18 14 15 13 0 9 1 9 7 9 2 13 0 9 1 11 11 11 2
9 0 13 9 7 1 0 1 9 2
10 3 13 14 15 13 0 9 1 9 2
8 15 13 9 1 9 1 9 2
1 9
1 9
4 9 11 13 0
24 1 9 1 9 11 9 1 0 9 2 9 13 12 9 2 2 15 13 3 0 7 0 7 13
12 13 14 13 1 3 2 16 6 15 13 9 2
4 13 0 9 2
18 3 9 11 13 1 0 9 7 13 12 0 9 2 15 15 13 9 2
18 1 1 4 13 1 0 9 2 9 11 15 13 7 13 0 12 9 2
10 3 15 13 3 0 13 1 10 9 2
6 14 15 6 13 9 2
14 13 1 12 9 1 9 2 9 1 9 13 10 9 2
28 13 1 12 9 7 15 13 1 10 15 2 6 4 13 14 12 9 2 3 0 9 2 13 1 9 1 9 2
11 13 4 1 9 7 4 13 1 9 9 2
10 9 2 12 9 11 2 3 15 13 9
36 3 3 13 9 1 0 0 9 14 15 13 9 1 9 1 9 2 11 11 2 2 9 1 9 2 12 9 11 2 2 13 0 9 11 11 2
22 1 12 9 7 9 2 1 9 1 0 0 9 2 9 4 13 2 16 4 13 9 2
17 13 15 2 16 1 9 2 15 3 13 1 0 9 2 13 9 2
21 0 0 9 2 11 2 2 15 3 15 13 1 9 2 15 13 1 9 1 11 2
33 15 4 13 1 11 2 12 9 11 2 2 1 1 13 0 15 9 7 9 3 13 1 9 1 9 7 1 0 9 2 13 11 2
27 1 9 7 9 0 9 13 3 14 13 7 13 9 2 7 1 9 13 2 3 9 15 13 9 1 9 2
5 11 13 3 1 11
5 13 9 1 0 9
8 9 4 13 1 9 1 9 2
14 15 15 13 3 14 13 9 0 9 1 9 7 9 2
12 1 1 12 9 13 12 9 9 1 12 9 2
12 1 15 15 13 0 9 2 15 4 3 13 2
10 1 10 9 9 12 1 9 15 13 2
5 1 0 4 13 2
18 3 15 13 7 0 9 1 0 0 9 2 15 3 13 1 12 9 2
8 0 9 3 13 3 1 9 2
20 13 15 2 16 15 4 13 1 9 2 15 13 9 15 7 13 9 1 9 2
13 12 9 7 0 13 14 15 13 1 12 9 3 2
13 1 9 4 13 12 0 9 2 15 13 12 9 2
14 0 9 2 9 2 13 0 9 1 0 9 1 9 2
15 3 1 9 1 9 13 12 9 1 11 2 11 2 11 2
12 1 12 9 15 4 4 13 2 13 1 11 2
22 0 9 3 4 13 14 13 0 2 0 2 0 7 0 9 2 1 14 13 1 9 2
24 15 13 0 9 1 0 9 1 9 1 9 1 9 1 9 1 9 1 0 9 2 13 9 2
6 0 9 13 12 9 9
8 2 0 9 2 13 9 1 11
17 9 1 2 11 2 11 11 13 9 1 9 1 2 0 9 2 2
4 9 2 11 11
9 0 9 13 0 15 9 1 12 9
5 11 11 2 11 11
18 9 1 2 11 2 3 6 15 13 1 9 1 9 1 9 11 11 2
13 1 2 11 2 13 1 3 12 9 9 1 9 2
11 0 9 3 14 13 9 1 11 7 9 2
19 1 0 9 13 3 0 9 2 13 7 9 1 0 9 1 11 11 11 2
12 1 11 13 12 9 9 1 9 1 0 9 2
20 1 11 2 16 3 15 13 9 3 1 0 9 2 3 14 13 9 1 9 2
24 9 1 9 1 2 0 9 2 6 15 4 13 1 9 1 0 9 2 13 9 9 11 11 2
16 11 15 13 1 0 0 9 1 0 9 2 15 13 10 9 2
22 3 13 14 13 3 0 9 2 7 13 1 9 15 2 3 7 1 9 1 9 1 9
8 13 14 13 3 1 10 9 2
17 15 13 1 9 1 11 1 9 0 9 2 7 1 9 1 9 2
6 3 13 9 1 9 2
14 3 16 13 9 7 6 13 10 4 13 14 15 13 2
14 2 9 1 11 2 0 1 11 13 1 9 2 9 2
28 11 4 13 7 0 9 1 15 11 11 2 13 9 2 11 2 2 16 15 13 1 0 9 1 11 11 11 2
30 1 9 4 13 0 9 1 9 11 7 11 11 2 0 1 0 9 2 11 2 1 0 12 9 1 9 2 13 11 2
12 11 11 6 4 13 1 2 11 2 1 9 2
22 12 2 12 2 12 9 2 9 1 2 11 2 13 1 9 1 9 1 11 1 9 2
8 9 1 9 13 1 12 9 2
16 1 15 12 1 9 14 4 13 2 7 11 7 11 14 13 9
20 9 0 9 1 9 1 11 1 9 15 1 11 11 1 9 0 9 1 11 11
19 11 13 9 1 0 9 2 15 13 3 1 9 1 9 1 2 11 2 2
15 0 9 1 11 14 13 3 15 13 9 1 9 11 11 2
21 9 1 2 11 2 11 11 13 2 16 13 9 1 15 2 7 9 13 1 11 2
6 0 9 13 9 1 11
2 0 9
6 9 7 9 13 1 11
5 11 11 2 11 11
17 1 0 9 1 9 1 9 1 11 1 0 9 13 0 9 1 9
10 15 15 13 1 9 1 0 0 9 2
13 9 15 13 3 1 9 2 0 1 9 1 11 2
11 1 11 9 3 13 14 15 13 1 11 2
11 12 9 1 9 4 13 1 0 9 11 2
19 1 9 1 0 9 1 11 9 11 11 9 6 4 13 1 9 1 11 2
16 9 1 9 1 0 9 1 11 7 0 15 9 6 4 13 2
12 1 11 9 1 9 1 9 6 13 10 9 2
15 9 1 9 1 9 15 13 12 9 3 2 9 7 9 2
17 3 1 0 9 0 9 4 4 13 2 3 9 7 9 4 13 2
11 3 9 14 13 0 9 1 9 1 9 2
7 9 13 0 1 9 9 2
9 9 15 13 3 3 2 13 9 2
8 9 1 0 9 13 1 9 2
8 0 9 13 1 9 7 9 2
17 13 15 9 1 9 2 9 7 9 1 0 9 2 13 1 11 2
10 9 13 0 9 2 0 1 0 9 2
10 0 13 1 12 9 2 13 3 3 2
15 9 3 13 9 1 0 2 9 2 9 2 9 7 9 2
6 9 13 14 15 13 2
17 1 0 11 9 13 1 9 9 9 7 15 13 1 9 7 9 2
25 0 9 11 11 2 9 1 0 0 9 2 13 3 1 9 15 1 11 1 0 12 2 12 9 2
5 13 9 1 9 2
23 9 1 11 13 0 1 0 9 2 1 14 13 2 16 13 14 13 9 7 1 10 9 2
12 1 9 0 0 9 14 13 10 9 1 11 2
34 0 9 13 2 13 15 2 14 13 10 9 1 11 11 2 3 0 9 4 15 13 1 0 9 1 0 10 9 2 0 9 11 11 2
9 15 2 13 15 2 6 13 0 2
7 3 11 13 9 1 11 2
15 11 13 10 0 9 1 9 1 0 9 2 15 9 13 2
28 1 11 11 13 3 3 2 7 3 15 6 15 13 10 9 2 15 6 13 9 2 3 1 14 13 10 9 2
8 1 9 14 13 10 9 3 2
33 1 16 1 3 9 1 11 13 9 2 1 11 11 15 13 9 2 1 14 13 0 9 1 9 1 11 1 9 1 0 15 9 2
24 11 13 0 0 9 2 15 13 14 13 0 1 9 2 7 7 15 3 13 1 10 0 9 2
22 15 3 4 13 9 1 12 9 9 3 7 3 14 6 13 9 1 10 10 0 9 2
16 9 1 9 1 11 7 1 11 4 3 13 7 1 0 9 2
9 15 13 10 11 2 2 4 13 11
25 3 16 2 9 2 1 11 3 13 1 9 1 9 1 11 7 15 3 15 13 1 2 11 2 2
5 14 9 14 13 2
12 7 3 14 9 14 4 13 3 1 0 9 2
21 1 9 0 0 9 1 9 13 1 9 1 10 14 11 14 13 0 9 1 11 2
19 13 15 2 16 15 13 9 2 7 16 11 11 15 13 2 13 12 9 2
15 1 9 1 0 0 9 4 13 0 0 9 1 0 9 2
11 9 1 9 6 13 9 2 16 13 9 2
15 13 3 3 9 1 9 1 10 9 2 3 14 13 3 2
29 3 3 13 2 16 1 9 1 0 9 11 13 10 9 2 7 16 15 13 3 9 1 11 2 15 6 13 0 2
10 0 0 0 9 15 13 14 13 11 2
16 3 14 14 13 9 1 11 2 14 15 13 14 1 0 9 2
9 0 9 1 0 9 13 3 0 2
14 0 13 9 1 11 3 2 3 10 9 13 1 9 2
12 7 3 11 13 1 9 1 0 9 1 9 2
29 3 1 9 2 0 15 1 0 9 2 11 2 2 3 1 9 1 9 2 11 2 2 13 12 9 14 15 13 2
19 0 15 13 0 15 9 1 11 2 9 11 11 2 0 9 1 0 9 2
16 15 13 0 0 9 2 7 1 12 9 3 15 13 12 9 2
16 11 13 2 9 2 2 13 14 15 13 14 13 14 9 15 2
18 0 15 4 13 0 2 7 15 13 1 0 9 1 0 2 13 15 2
31 1 0 9 0 9 13 1 11 1 10 9 2 9 2 10 9 13 1 9 2 11 2 2 0 1 9 1 9 1 11 2
30 6 13 14 13 9 1 9 15 2 3 16 13 9 2 15 14 15 13 1 10 9 7 3 1 0 9 1 0 9 2
16 13 3 7 1 0 0 9 2 1 9 1 9 1 0 9 2
20 13 15 2 3 9 15 13 3 3 1 9 2 13 1 12 9 1 10 9 2
20 0 9 13 1 9 2 10 9 15 13 1 3 9 2 0 9 13 3 0 2
20 0 9 13 1 9 2 10 9 15 13 1 3 9 2 0 9 13 3 0 2
24 1 9 9 1 9 1 9 15 15 13 0 2 1 14 15 13 2 16 13 3 14 13 11 2
11 13 15 14 15 13 1 11 1 0 9 2
20 3 13 1 9 2 9 2 2 9 2 3 0 2 7 15 13 9 1 9 2
35 6 13 1 9 10 9 2 6 15 13 14 13 7 9 1 9 2 7 14 13 1 9 2 3 7 14 13 9 1 3 0 15 9 1 9
37 9 15 13 7 3 9 2 13 15 9 2 13 15 3 7 13 0 9 2 10 15 13 9 2 3 6 13 14 13 3 0 9 2 13 15 15 2
13 1 9 9 1 9 7 9 1 9 9 15 13 2
28 7 9 13 2 1 1 3 13 9 1 9 1 9 2 16 3 13 14 13 1 11 1 9 2 0 1 9 2
7 7 3 15 13 1 11 2
8 3 9 6 13 2 9 13 2
7 15 6 13 15 13 1 9
13 13 3 0 9 1 9 7 9 15 13 1 9 2
14 7 15 4 13 9 2 0 9 1 9 2 1 9 2
20 10 2 16 1 14 15 13 1 0 9 2 15 4 13 14 13 9 11 11 2
6 15 6 15 13 3 9
6 0 9 15 13 3 2
22 16 13 0 9 1 11 9 2 10 9 15 13 1 9 7 9 7 1 9 1 15 2
41 13 15 3 3 1 0 9 2 16 14 13 0 2 13 3 1 9 1 0 9 1 0 9 1 2 0 9 2 1 11 11 2 3 7 1 9 1 9 11 11 2
21 13 3 2 7 1 9 2 7 1 9 1 0 9 7 1 9 15 13 1 0 2
14 9 13 1 9 2 7 1 15 13 7 9 2 2 2
8 9 13 1 9 2 6 15 13
28 1 9 3 13 9 7 1 9 13 0 9 2 9 15 11 11 2 9 1 9 15 2 15 15 13 1 9 2
18 3 13 0 9 2 15 13 1 9 1 11 9 2 13 3 9 15 2
16 3 6 13 14 15 13 9 14 13 1 0 2 7 3 15 13
15 13 3 9 1 9 0 9 7 15 13 1 9 1 9 2
5 3 15 13 1 0
14 14 6 15 13 2 3 1 10 9 1 9 13 9 2
7 7 13 1 9 1 9 2
13 1 0 0 9 13 1 0 9 2 3 1 11 2
13 1 11 6 13 2 7 16 15 13 9 2 13 0
27 2 11 2 8 8 2 2 13 15 9 11 1 0 2 15 13 1 0 2 2 12 9 2 14 15 13 2
10 11 15 13 2 16 0 9 13 11 2
45 1 0 9 9 15 13 14 15 13 9 2 13 12 9 7 15 13 1 9 15 2 9 7 9 1 11 2 0 9 1 9 2 9 7 9 1 11 2 9 1 12 9 1 11 2
8 13 0 9 1 9 1 11 2
38 7 3 16 13 3 14 15 13 1 15 2 11 15 13 1 0 15 9 2 1 0 9 13 10 0 0 9 2 0 1 9 2 9 2 9 7 9 2
8 11 13 0 9 2 6 13 9
12 9 1 11 1 11 13 3 0 1 9 7 9
16 9 1 2 11 11 2 11 13 7 0 0 9 1 3 0 9
14 2 11 11 2 13 0 9 1 0 9 1 0 9 2
20 1 9 9 1 12 0 9 13 3 0 2 7 1 9 15 13 7 0 9 2
12 1 9 1 9 15 13 10 0 9 1 9 2
24 9 1 9 13 1 10 2 16 15 13 9 1 3 0 2 7 0 9 1 9 1 0 9 2
16 7 3 15 13 3 0 9 1 0 15 9 7 0 0 9 2
10 9 1 0 9 1 11 3 13 0 2
10 9 3 14 13 1 9 1 0 9 2
10 0 3 13 9 1 9 1 0 9 2
13 0 9 13 3 0 9 2 7 6 13 0 9 2
22 3 1 15 9 1 9 13 3 0 1 0 9 7 9 1 0 9 4 13 1 12 2
14 15 6 13 0 9 2 7 13 0 1 9 7 9 2
15 1 10 9 15 13 3 0 9 7 9 1 3 9 9 2
7 9 4 13 7 1 9 2
7 1 0 9 3 13 9 2
20 0 1 9 13 0 0 11 0 9 1 1 12 9 1 9 7 9 12 9 2
12 3 0 13 7 0 0 9 1 9 12 9 2
10 1 15 9 12 2 12 13 12 9 2
22 1 15 0 9 15 13 7 1 2 0 2 0 9 1 9 12 9 7 9 12 9 2
19 9 13 14 15 13 3 1 0 9 2 3 7 1 0 9 2 11 2 2
37 1 12 9 1 2 9 2 13 14 15 13 1 9 15 7 15 13 1 9 3 9 2 3 16 11 15 13 1 9 1 0 9 1 11 11 11 2
18 9 13 1 12 9 2 7 1 9 14 15 13 1 9 1 0 9 2
17 11 14 13 0 9 1 2 11 2 1 9 2 15 14 13 3 2
19 9 2 11 2 6 13 1 9 7 3 15 13 15 14 13 14 1 9 2
13 9 7 9 13 2 3 9 2 1 9 2 11 2
16 0 9 13 9 11 1 11 2 9 15 13 1 2 0 9 2
29 9 11 2 9 11 7 9 15 11 2 9 11 11 7 11 11 2 0 9 13 0 1 0 9 7 11 0 9 2
15 12 9 1 9 1 9 14 15 13 0 9 4 13 3 2
12 3 0 9 15 13 1 9 1 9 7 9 2
14 10 0 9 13 9 2 9 2 9 2 9 2 9 2
5 12 13 0 9 2
15 9 1 10 9 13 7 3 13 1 0 9 1 12 9 2
9 3 1 9 3 13 9 1 9 2
7 9 15 13 1 0 9 2
28 1 9 1 9 9 1 9 13 11 11 7 11 2 9 2 11 2 2 0 11 2 11 2 2 11 2 11 2
13 1 9 15 13 7 0 1 9 11 7 11 11 2
8 3 12 9 15 13 3 9 2
12 12 9 1 12 9 15 13 7 9 11 11 2
23 15 4 13 1 9 15 11 2 9 1 9 15 11 11 7 9 15 11 11 7 11 11 2
12 13 12 9 2 15 3 13 1 9 7 9 2
5 14 15 13 1 9
5 3 14 14 13 9
9 12 9 13 2 3 9 2 1 9
17 0 1 9 7 3 0 2 11 7 11 11 3 15 13 1 9 2
12 0 9 13 1 0 9 1 0 9 0 9 2
16 1 9 1 0 9 15 13 3 9 1 9 1 2 11 2 2
30 9 2 9 1 0 9 7 1 0 9 2 9 1 11 4 13 1 0 9 2 9 1 9 2 9 2 9 7 3 2
9 1 9 2 9 13 1 0 9 2
17 3 9 15 13 1 0 2 7 1 3 9 13 2 3 0 2 2
3 0 2 9
7 14 13 1 9 1 11 2
13 7 3 2 7 1 0 9 13 0 9 1 9 2
5 9 13 3 0 2
10 13 15 14 15 13 3 3 7 3 2
7 14 6 13 14 15 13 2
16 0 9 2 0 9 2 0 9 2 10 13 0 9 1 9 2
10 16 15 13 10 9 2 15 13 3 2
6 13 15 3 0 9 2
10 1 0 13 10 9 1 9 1 9 2
11 15 1 10 9 13 0 1 10 0 9 2
9 1 9 6 13 14 13 1 9 2
7 13 14 13 14 15 13 2
7 6 2 15 13 3 0 2
9 3 9 4 13 2 9 13 9 2
10 9 11 7 9 11 15 13 1 9 2
13 9 9 15 13 1 9 2 11 2 14 13 9 2
11 9 13 3 9 2 1 14 13 1 9 2
5 9 15 15 13 2
23 0 9 1 11 1 0 1 9 1 9 9 1 9 1 9 3 6 13 9 1 0 9 2
10 3 13 9 1 0 9 1 0 9 2
16 16 6 13 0 9 2 16 13 10 0 9 1 9 7 9 2
14 3 1 9 0 9 3 6 13 1 9 1 9 15 2
31 9 3 14 15 13 1 9 1 9 2 16 15 15 13 2 16 0 0 9 1 9 14 13 9 1 10 9 2 13 0 2
11 9 1 9 6 15 13 1 9 1 9 2
15 0 9 1 9 1 9 1 9 13 9 1 9 7 9 2
23 16 6 13 14 13 9 15 1 0 9 2 1 1 13 15 14 15 13 7 9 1 15 2
37 7 1 10 0 15 9 7 1 3 0 9 1 0 9 14 15 13 1 9 1 0 9 7 9 3 9 1 9 6 13 1 3 0 9 1 9 2
5 15 14 15 13 2
8 9 2 3 0 1 0 9 2
10 9 13 12 9 9 1 2 0 9 2
9 0 9 13 9 1 9 1 11 11
18 12 9 0 0 9 1 0 9 4 13 1 2 0 9 2 2 11 2
13 11 2 0 9 7 0 9 2 13 9 1 9 2
11 1 9 13 2 16 9 4 13 1 9 2
9 9 4 13 1 0 9 0 9 2
23 1 9 1 2 0 9 2 0 9 13 2 16 1 0 9 0 9 9 4 13 1 9 2
25 0 1 15 9 13 2 16 1 9 2 0 1 2 0 9 2 2 4 15 13 12 9 0 9 2
30 1 0 9 1 9 1 2 11 2 1 11 14 13 12 9 9 2 7 9 1 2 11 2 3 15 13 1 0 9 2
10 0 9 1 9 13 1 12 12 9 2
25 9 1 11 13 14 13 2 0 9 2 1 9 1 9 1 11 11 2 16 3 13 9 1 9 2
15 1 9 1 0 9 0 9 13 9 7 9 3 13 0 2
27 1 9 1 0 9 15 4 3 13 2 16 15 13 2 16 0 9 4 13 1 0 9 7 2 11 2 2
17 9 13 0 9 1 0 0 9 2 7 9 13 0 0 0 9 2
8 7 12 9 13 0 1 9 2
18 9 2 11 2 13 0 9 1 12 9 2 0 0 9 7 0 9 2
18 7 12 9 13 9 1 10 0 9 1 9 2 15 13 3 0 9 2
7 0 9 15 13 1 0 9
10 12 9 9 1 9 2 15 6 13 9
17 1 9 1 12 9 14 4 13 10 2 15 13 9 1 10 9 2
10 15 13 1 0 0 9 2 11 2 2
13 0 9 13 9 2 10 9 13 3 0 1 9 2
15 0 9 13 9 15 1 0 9 14 13 1 12 12 9 2
12 1 9 15 13 3 14 6 4 13 1 11 2
33 9 13 1 9 0 9 2 1 15 15 13 9 2 9 1 9 2 9 1 9 1 9 2 9 7 9 2 3 7 1 0 9 2
22 3 9 13 3 1 9 2 9 15 13 3 1 9 1 9 2 1 15 14 15 13 2
8 9 13 12 9 1 0 9 2
22 9 15 13 3 7 1 0 9 1 0 9 1 9 1 9 7 3 13 9 1 9 2
12 9 13 14 4 13 7 1 9 1 0 9 2
15 14 9 14 4 13 1 9 2 9 15 13 1 0 9 2
12 9 1 10 9 15 13 1 9 1 0 9 2
14 15 14 13 12 9 9 16 1 10 9 13 0 9 2
21 9 15 13 1 0 9 2 1 0 9 7 1 0 9 1 9 1 0 0 9 2
13 9 2 15 14 15 13 1 0 9 1 0 9 2
3 9 1 3
5 9 1 9 1 3
2 0 9
3 9 1 9
5 9 7 9 2 9
3 9 1 9
7 9 2 9 2 9 7 9
12 0 9 2 9 1 0 9 2 0 9 1 9
10 9 1 9 2 0 9 2 9 2 9
7 9 1 9 2 9 2 9
16 9 1 0 9 2 9 2 9 9 2 0 9 2 9 7 9
13 1 0 9 9 15 13 1 12 9 1 0 9 2
23 15 13 9 1 9 1 11 11 2 13 1 0 9 7 15 13 1 9 1 9 11 11 2
25 1 12 0 9 11 13 9 1 0 9 1 0 9 2 7 3 3 2 9 2 13 1 11 11 2
3 0 1 9
3 0 0 9
2 11 11
22 13 9 1 9 1 9 0 9 7 3 13 9 1 0 9 2 9 13 0 1 9 2
9 3 3 0 9 13 9 1 9 2
13 16 13 14 13 9 1 9 7 9 1 10 9 2
17 13 14 15 2 9 1 3 0 9 13 10 9 14 13 7 0 2
16 7 14 13 15 3 2 1 14 15 13 1 9 1 9 15 2
8 3 13 9 2 6 13 3 2
12 9 1 0 9 13 9 1 9 15 1 9 2
8 3 7 15 13 2 16 13 2
10 7 3 1 0 10 9 13 14 13 2
7 13 15 10 0 0 9 2
10 1 15 9 2 1 15 4 13 0 2
14 14 15 13 3 2 14 13 15 14 1 0 0 9 2
7 9 13 0 9 1 0 9
9 9 13 0 0 9 1 0 9 2
31 9 1 11 11 11 7 11 11 13 9 1 0 9 2 11 2 0 9 2 2 0 1 9 2 9 2 11 2 7 11 2
28 1 9 2 1 9 1 2 11 2 11 11 2 13 11 11 2 2 11 2 2 7 11 11 2 11 11 2 2
14 0 0 9 13 1 12 9 2 0 1 1 12 9 2
21 9 4 13 7 1 0 9 1 9 12 2 0 1 9 9 12 1 0 9 11 2
5 0 9 13 1 11
14 1 11 14 13 0 9 11 11 11 7 9 1 9 2
6 2 11 2 13 1 9
7 11 13 9 1 2 11 2
13 1 10 9 9 1 0 9 13 0 9 1 9 2
11 1 12 13 0 9 1 9 1 9 1 11
15 9 13 0 1 9 1 9 0 9 2 1 0 9 2 2
11 0 9 1 0 9 13 9 1 2 11 2
20 1 12 9 0 9 1 11 1 2 11 2 3 4 13 1 0 9 1 11 2
16 9 13 12 9 1 0 9 7 4 13 1 0 2 11 2 2
22 1 1 9 13 1 0 9 1 9 2 9 0 1 10 9 9 1 9 13 1 9 2
10 15 13 0 9 7 15 13 1 9 2
8 1 9 4 13 7 3 9 2
5 1 9 13 9 2
13 9 13 9 3 12 9 1 9 14 13 3 9 2
20 1 10 9 3 9 1 9 11 11 11 11 11 3 15 13 9 14 6 13 2
9 3 9 13 9 1 9 11 11 2
27 1 0 9 1 0 9 4 13 9 1 9 1 9 1 12 9 1 9 2 0 1 0 9 1 10 9 2
7 0 0 9 1 2 11 2
19 1 9 1 0 0 2 11 11 2 13 12 9 9 9 1 0 0 9 2
13 0 9 13 9 1 9 1 0 9 1 0 9 2
19 1 9 1 9 6 4 13 12 9 3 1 0 0 9 7 0 0 9 2
18 3 7 4 3 13 2 1 1 3 9 15 13 1 9 1 12 9 2
22 3 12 9 1 11 2 15 13 14 15 13 3 2 4 13 1 0 9 7 0 9 2
7 11 15 13 1 9 1 11
17 9 15 11 11 15 13 1 0 9 2 3 1 9 13 3 9 2
27 1 1 13 9 1 11 1 9 15 11 2 9 14 13 1 0 2 9 2 1 11 2 9 12 12 2 2
11 3 9 1 0 9 4 13 12 9 3 2
13 1 9 12 9 1 9 15 14 13 9 1 9 2
6 11 13 12 9 11 9
14 0 9 12 1 9 11 11 14 13 9 12 9 11 2
16 9 15 11 13 1 9 1 9 1 9 12 9 7 12 9 2
37 1 0 9 4 13 9 1 11 11 11 1 2 0 9 1 9 1 9 7 9 2 7 15 13 3 9 2 3 13 14 15 13 1 9 1 15 2
7 7 13 7 0 2 2 2
13 0 9 4 13 1 9 1 0 9 1 0 9 2
24 9 15 13 1 9 2 15 13 3 0 9 1 0 2 0 9 2 2 0 1 9 1 9 2
6 13 15 9 1 0 9
25 1 9 1 0 9 1 11 14 11 13 0 9 1 9 1 12 9 1 0 9 3 1 10 9 2
9 9 14 4 13 3 1 9 3 2
19 1 10 9 0 0 9 1 9 13 1 12 9 1 0 9 1 12 9 2
17 9 1 0 9 1 9 4 13 1 9 1 12 9 1 0 9 2
17 9 1 9 1 0 9 0 9 4 13 1 0 9 1 12 9 2
16 0 1 9 9 1 0 9 13 9 1 11 1 0 0 9 2
28 1 0 9 13 7 9 11 0 2 12 9 2 2 11 11 2 12 9 2 2 9 11 0 2 12 9 2 2
42 1 0 12 0 9 13 3 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 2
18 9 1 11 13 2 16 3 1 9 1 9 4 13 9 2 12 9 2
10 1 0 9 1 9 13 9 2 12 2
10 9 3 6 15 13 1 0 15 9 2
10 1 9 3 0 13 11 7 0 9 2
7 1 15 4 13 12 9 2
25 1 9 12 9 15 13 14 14 13 2 12 9 13 0 9 1 11 2 7 12 9 13 0 9 2
19 0 9 13 9 1 12 9 1 0 2 7 1 0 9 15 13 12 9 2
29 1 9 1 9 15 13 12 9 1 0 7 12 9 1 9 2 7 9 13 12 9 1 9 7 12 9 1 9 2
17 1 9 15 13 9 1 9 1 9 1 0 9 1 0 15 9 2
23 9 1 11 9 11 11 13 9 7 13 9 11 11 1 0 15 9 1 9 2 13 11 2
12 11 7 11 13 9 1 0 9 1 0 9 2
11 15 6 4 13 14 3 9 4 13 10 9
12 9 1 9 11 11 1 11 13 1 11 11 2
6 13 15 1 0 9 2
12 13 14 13 3 0 15 9 2 1 14 15 13
23 15 13 9 1 2 0 9 2 2 9 2 0 1 0 9 1 11 2 1 9 1 11 2
14 15 15 15 13 2 15 13 9 14 13 1 11 11 2
6 1 15 9 6 13 2
14 15 15 13 9 11 11 2 2 9 2 1 0 9 2
10 9 11 2 11 13 0 1 9 1 9
8 9 15 13 2 13 2 11 2
11 0 9 3 15 13 2 7 6 15 13 2
20 3 13 9 1 0 9 1 9 7 9 2 15 13 1 9 7 13 3 9 2
10 3 9 15 13 2 15 3 4 13 2
16 1 10 9 9 1 0 9 13 3 0 7 9 13 3 0 2
25 0 0 9 4 3 13 2 16 9 1 9 15 13 14 13 9 1 9 2 13 1 2 11 2 2
10 9 2 11 2 11 2 13 1 0 9
15 1 9 1 12 9 9 14 13 0 9 1 12 12 9 2
8 0 9 1 9 13 12 9 2
33 1 16 9 1 9 13 3 0 2 3 1 9 15 13 9 11 11 2 9 1 0 12 9 2 11 11 2 15 13 1 0 9 2
12 12 3 0 9 1 9 1 9 3 13 3 2
16 15 13 0 9 1 0 9 1 9 11 11 7 9 11 11 2
10 11 11 13 0 9 1 9 1 12 9
10 11 11 13 0 9 1 9 1 12 9
17 3 3 13 10 1 9 11 2 15 13 9 1 9 1 0 9 2
13 15 13 12 9 7 13 0 9 1 0 11 11 2
21 0 0 9 1 9 15 13 1 0 9 3 9 1 12 9 1 2 0 9 2 2
9 15 13 0 9 1 0 11 11 2
12 3 0 13 9 1 0 9 1 9 1 0 2
10 15 13 14 13 3 0 9 1 9 2
22 11 2 15 13 1 12 9 1 0 9 0 9 2 13 9 15 1 0 15 9 9 2
23 1 9 1 3 15 9 2 0 1 0 1 9 9 11 7 11 2 9 14 13 9 11 2
12 9 13 0 9 1 11 3 1 9 1 9 2
7 0 13 3 1 0 9 2
11 3 1 0 9 4 13 7 9 1 0 2
8 0 13 9 1 2 11 2 2
12 15 13 0 9 1 9 1 0 9 1 9 2
17 9 13 9 9 12 1 11 1 0 9 1 9 1 0 9 11 2
21 9 11 11 11 7 11 11 11 11 2 15 13 1 12 0 9 2 13 1 9 2
33 11 13 0 9 1 9 1 9 1 9 7 9 1 11 1 11 1 11 7 11 2 13 0 1 11 0 9 2 11 11 11 2 2
22 1 9 1 0 9 11 13 9 3 7 15 13 14 13 9 1 0 9 1 12 9 2
30 1 0 9 9 11 11 2 0 1 2 12 9 2 2 3 1 9 6 4 13 9 1 2 10 0 9 1 9 2 2
40 1 16 1 0 9 11 7 11 4 13 14 13 0 9 1 11 14 1 0 9 2 1 0 9 1 11 13 9 1 9 1 9 7 9 1 9 1 0 9 2
6 9 7 9 13 0 9
7 0 9 13 1 9 1 9
6 9 13 1 9 7 9
11 1 11 0 9 13 1 9 2 13 11 2
20 3 1 9 9 13 1 0 0 9 11 2 3 1 9 3 9 13 0 9 2
19 1 9 1 9 13 4 12 9 2 1 15 12 9 13 1 9 1 9 2
22 9 1 11 13 2 16 9 13 9 2 16 9 4 4 13 1 0 0 9 1 9 2
23 12 9 13 1 9 1 9 1 0 9 1 0 9 11 1 9 1 0 9 2 13 11 2
23 12 9 13 1 9 1 9 1 0 9 1 0 9 11 1 9 1 0 9 2 13 11 2
9 9 3 15 13 1 9 1 9 2
7 12 9 4 13 1 9 2
18 3 12 9 4 4 13 1 9 1 0 9 1 9 1 0 9 11 2
18 0 9 4 13 7 1 9 11 2 3 9 13 9 1 12 0 9 2
16 1 0 9 1 11 11 1 0 9 15 13 9 1 0 9 2
19 0 9 11 11 13 14 15 13 1 0 2 11 11 2 2 13 0 9 2
22 16 11 13 0 9 2 3 1 0 9 14 13 0 1 9 1 2 11 2 11 11 2
6 7 11 13 9 1 9
9 1 3 11 13 0 9 1 9 2
18 1 9 1 0 0 9 1 9 14 13 14 15 13 9 7 1 9 2
15 1 9 1 9 9 14 4 13 3 1 9 7 1 9 2
16 12 9 1 15 12 9 2 9 7 9 2 14 15 13 3 2
4 3 9 1 9
36 0 9 1 9 4 13 1 9 1 9 1 0 2 3 13 9 2 7 9 1 0 9 3 15 13 1 0 9 1 9 1 0 9 1 9 2
4 2 11 11 2
12 15 3 13 10 3 0 9 1 10 0 9 2
9 7 15 13 0 9 1 9 15 2
10 3 16 9 15 1 10 9 13 0 2
15 0 13 9 2 16 9 15 13 1 0 0 9 1 9 2
7 7 10 9 13 3 0 2
13 3 9 1 9 13 9 7 9 1 0 15 9 2
34 1 3 0 9 1 9 0 9 13 7 9 1 9 2 15 13 9 1 0 9 1 9 1 9 7 13 9 0 0 9 14 13 3 2
22 6 13 14 15 13 1 9 1 0 9 2 15 13 14 15 13 1 9 1 0 9 2
17 3 1 9 7 9 1 9 1 0 9 13 9 1 0 0 9 2
10 2 15 6 13 14 4 13 1 9 2
23 11 7 1 15 13 1 0 9 1 10 0 9 2 3 9 1 9 13 3 0 1 15 2
16 2 13 6 13 2 16 14 13 10 9 3 1 9 1 9 2
5 2 3 6 13 2
23 16 13 9 7 9 1 9 2 14 13 1 9 1 0 9 2 7 15 6 4 13 3 2
20 1 0 9 3 2 15 13 16 10 9 13 0 7 15 15 13 1 10 9 2
15 7 15 13 0 9 1 9 1 0 0 9 1 0 9 2
5 2 15 13 15 2
16 2 11 3 13 1 9 1 0 9 2 7 1 15 13 9 2
11 7 3 9 1 0 9 13 1 0 9 2
22 14 13 2 16 14 13 9 7 0 9 2 13 3 2 7 15 6 13 9 1 9 2
12 0 0 9 13 10 9 1 0 9 14 13 2
21 13 0 9 1 10 9 1 0 9 2 15 13 0 9 2 9 2 9 2 2 2
19 13 14 9 1 9 1 9 1 9 3 14 15 13 1 9 1 10 9 2
11 2 1 9 15 13 3 7 15 13 0 2
28 7 1 1 13 2 16 15 6 13 9 1 0 15 9 2 15 3 15 13 1 15 1 3 0 7 0 9 2
12 2 6 13 9 1 0 9 1 9 1 9 2
43 3 2 15 7 9 15 13 1 0 9 1 0 9 2 3 3 3 15 13 1 9 1 0 9 1 0 9 1 9 7 9 1 0 9 1 9 2 0 1 0 0 9 2
18 7 0 9 1 0 13 0 9 7 9 2 15 13 14 13 0 9 2
16 13 14 9 1 15 14 13 9 1 9 7 1 9 1 11 2
13 0 9 1 0 9 3 13 3 0 9 1 9 2
2 9 2
5 3 13 11 2 9
7 15 3 13 1 9 15 2
7 13 7 14 15 15 13 2
6 13 7 14 13 9 2
13 7 6 13 2 16 10 9 1 9 13 11 11 2
14 15 13 9 1 9 1 9 1 9 2 11 11 2 2
16 3 1 9 3 13 11 11 2 0 1 11 11 7 11 11 2
20 9 13 9 1 9 1 9 2 0 1 0 9 1 11 7 11 1 0 9 2
20 1 9 12 1 11 14 13 9 1 9 1 11 1 2 0 9 2 1 11 2
10 1 9 14 13 7 0 9 11 11 2
26 11 11 2 0 2 0 2 13 9 1 0 0 9 7 9 1 0 9 9 11 11 7 9 11 11 2
8 1 10 9 3 13 9 12 2
15 9 1 2 11 2 13 1 0 9 2 1 15 13 9 2
5 0 2 0 2 0
9 9 13 1 9 2 13 15 1 9
17 11 4 13 3 1 9 2 3 1 0 15 9 6 13 1 9 2
37 9 1 2 11 11 2 11 11 2 1 9 3 2 13 9 12 1 9 1 0 9 1 0 9 2 11 2 2 13 9 1 2 9 2 11 11 2
12 11 13 14 13 12 9 1 0 9 1 9 2
9 0 9 13 3 1 0 0 9 2
15 11 11 7 11 11 14 13 0 9 1 11 1 0 9 2
13 9 15 1 0 9 14 13 1 9 1 12 9 2
18 9 9 12 1 11 13 0 9 1 2 11 2 2 11 2 11 11 2
14 1 9 1 9 2 11 2 13 12 9 7 12 9 2
28 0 9 2 15 13 3 1 9 1 0 9 2 13 1 9 0 9 1 11 11 2 11 2 1 9 1 9 2
15 11 13 1 9 1 0 9 1 9 1 11 2 11 2 2
18 0 9 2 0 15 1 11 2 13 0 9 1 0 9 1 0 9 2
6 9 15 13 1 9 11
23 3 1 10 9 15 13 11 14 13 0 9 7 3 1 9 9 14 13 14 13 9 15 2
26 1 9 4 13 9 7 9 14 13 0 9 2 15 14 13 9 1 10 9 2 7 9 13 1 9 2
10 9 1 11 15 13 3 1 0 9 2
12 0 9 13 0 2 3 3 9 3 13 9 2
14 16 13 9 1 9 2 15 3 6 13 14 15 13 2
20 3 9 7 9 13 14 13 1 9 2 3 15 13 9 7 9 2 13 9 2
3 9 1 9
3 9 1 9
7 3 0 13 0 0 9 2
4 0 0 9 2
5 11 15 13 14 13
21 1 2 9 1 0 9 2 12 2 11 11 13 15 14 2 9 2 11 2 2 2
15 7 1 11 11 4 13 9 1 9 1 11 3 1 9 2
4 0 9 1 9
6 1 11 15 13 7 11
7 1 0 9 3 14 15 13
6 6 2 6 2 3 2
5 15 13 0 9 2
7 13 2 16 13 3 9 2
3 10 9 2
2 13 2
5 3 14 13 0 2
7 14 3 6 13 10 9 2
13 10 2 15 13 3 1 15 2 15 13 10 9 2
9 6 13 14 15 13 1 10 9 2
14 0 9 1 9 7 9 1 9 6 15 13 3 0 2
7 3 13 14 15 13 9 2
2 3 2
10 11 6 13 0 7 9 6 13 0 2
9 9 1 9 7 9 1 10 9 2
2 15 2
10 14 6 13 3 2 15 13 0 9 2
13 13 2 16 6 13 14 15 13 9 1 9 2 2
3 1 9 2
5 1 3 13 9 2
11 9 15 1 9 3 4 13 0 2 2 2
7 2 11 2 13 9 1 9
10 2 11 11 2 13 0 9 1 9 2
14 1 0 9 1 9 13 11 11 2 15 13 12 9 2
15 11 13 7 12 9 1 9 2 7 11 11 13 12 9 2
5 1 9 13 3 2
6 3 9 15 15 13 3
17 9 11 11 6 13 1 9 2 0 15 1 9 1 9 11 11 2
9 0 9 1 9 1 0 9 1 11
14 14 13 7 9 1 0 9 7 0 9 1 0 9 2
29 1 12 0 9 1 0 9 7 9 14 4 13 1 9 1 0 9 1 0 9 1 9 1 9 1 9 1 9 2
14 13 4 7 0 9 1 9 1 12 9 1 12 9 2
15 9 1 0 9 15 13 1 9 2 7 3 1 9 2 2
10 7 0 2 0 9 13 1 0 9 2
13 1 9 9 1 0 11 13 1 0 1 9 15 2
24 2 15 13 7 3 0 9 2 16 3 11 7 11 13 1 0 12 9 1 9 1 9 2 2
13 12 11 4 3 13 1 9 2 9 2 9 2 2
12 0 2 1 0 11 13 3 0 9 1 9 2
12 0 2 1 0 11 13 3 0 9 1 9 2
15 9 3 13 0 11 2 3 3 15 13 9 0 9 3 2
27 1 11 11 14 3 6 4 13 9 1 9 1 9 2 3 13 0 9 1 2 11 11 2 1 0 9 2
10 7 10 9 12 9 1 9 13 9 2
27 1 0 0 9 9 1 9 2 15 13 1 0 9 2 13 3 0 1 9 1 10 2 15 13 0 9 2
9 0 7 3 0 9 3 13 11 2
22 3 7 3 12 9 1 9 7 12 9 1 9 13 1 9 1 0 9 1 0 9 2
10 3 13 2 9 13 0 7 0 9 2
14 12 9 13 2 16 15 14 13 3 0 1 0 9 2
5 12 9 13 9 2
4 0 15 13 2
13 6 13 14 0 15 1 9 1 11 1 10 9 2
11 1 1 11 13 0 9 1 9 1 11 2
19 1 9 0 9 1 0 9 1 2 11 11 2 13 3 9 1 10 9 2
13 1 10 9 9 13 0 9 1 11 1 0 9 2
20 2 9 11 2 10 15 13 1 9 9 1 0 9 2 0 1 2 11 2 2
6 2 15 13 0 9 2
4 9 13 0 2
11 3 16 14 15 13 14 13 3 0 9 2
10 1 9 13 1 9 7 9 1 9 2
5 7 13 1 9 2
12 0 9 3 15 13 14 13 10 9 1 11 2
5 3 14 13 15 2
11 3 13 14 15 13 9 7 1 0 9 2
6 6 13 3 13 9 2
8 1 9 13 0 9 1 11 2
23 13 15 2 13 1 9 2 15 13 10 0 9 7 15 15 13 14 15 13 1 0 9 2
14 2 3 13 9 1 9 1 9 1 0 2 11 2 2
20 2 15 13 9 2 15 13 14 15 13 1 0 9 1 9 2 2 11 2 2
12 13 1 9 11 11 7 1 9 15 11 11 2
7 9 1 2 11 2 13 2
18 13 0 12 9 2 9 12 2 2 1 14 13 14 13 2 11 2 2
6 9 6 13 1 15 2
20 2 1 9 11 4 13 2 16 13 3 14 13 9 1 9 1 2 11 2 2
7 13 14 4 1 10 9 2
7 2 3 3 14 15 13 2
7 13 4 15 9 1 9 2
9 13 3 10 0 9 1 10 9 2
14 3 13 3 2 1 0 9 7 9 1 9 13 3 2
22 3 15 13 9 7 1 11 11 2 7 1 11 11 2 1 11 11 2 1 11 11 2
16 7 1 3 14 10 0 9 6 4 13 1 9 1 11 11 2
29 0 9 6 13 1 9 1 2 9 2 1 9 15 2 1 15 3 13 2 16 6 13 0 1 11 7 9 15 2
16 1 0 9 11 11 4 4 13 2 16 1 9 13 9 15 2
7 3 9 15 13 3 0 2
21 3 13 14 15 13 2 16 9 1 0 9 7 10 9 4 13 1 9 1 9 2
37 3 7 6 15 13 9 1 9 1 3 1 9 7 3 16 9 7 9 6 13 0 9 2 9 4 13 1 0 9 7 3 3 1 9 1 0 2
7 15 13 10 9 7 9 2
6 3 0 9 13 0 2
32 9 1 0 9 13 1 0 9 0 9 1 0 9 1 9 1 11 2 11 11 7 9 15 11 11 2 11 11 7 11 11 2
53 9 13 2 16 2 1 9 15 1 0 9 1 9 1 0 9 1 9 7 9 0 9 12 3 6 4 13 3 9 1 9 2 9 7 9 1 9 7 9 1 0 9 1 0 9 1 9 1 9 0 9 2 2
25 3 12 9 9 1 11 13 9 1 12 12 9 9 2 7 9 2 11 2 15 13 1 12 9 2
15 13 4 3 3 12 9 9 1 9 12 12 12 12 9 2
21 7 9 3 13 15 2 0 9 1 0 2 9 15 1 9 2 0 9 1 9 2
13 9 1 2 11 2 3 4 13 1 12 9 9 2
20 1 9 1 11 2 16 0 9 13 9 1 0 0 9 2 0 6 15 13 2
14 12 9 15 4 13 0 9 1 9 1 11 2 7 13
17 7 14 7 10 1 0 9 1 9 6 13 14 13 15 13 15 2
18 16 2 9 2 13 2 13 14 13 0 9 7 0 0 9 1 0 9
31 1 9 1 0 9 2 9 2 13 9 1 9 2 11 2 1 0 9 1 9 12 9 2 15 13 14 13 1 12 9 2
10 1 10 9 9 13 9 1 9 15 2
8 9 13 0 0 9 11 11 2
18 9 3 6 13 9 15 7 2 9 2 13 1 9 1 9 0 9 2
25 1 9 1 9 0 9 11 13 9 15 11 11 2 16 15 13 1 0 9 1 12 9 9 9 2
5 9 13 0 9 2
8 2 11 2 13 2 11 2 2
11 7 15 6 13 2 16 13 14 4 13 2
7 9 13 11 1 9 1 11
9 3 13 9 1 11 1 9 1 9
21 1 0 9 15 13 9 1 11 1 0 9 7 9 1 9 1 11 1 0 9 2
14 1 9 1 9 4 13 10 9 1 11 2 13 11 2
29 9 1 11 11 15 13 1 9 14 15 13 9 1 0 9 2 3 16 15 4 13 1 9 1 0 9 1 9 2
9 1 15 3 1 9 3 13 9 2
6 13 9 1 9 1 9
16 0 0 9 1 0 9 1 9 1 0 11 13 3 1 11 2
19 15 14 4 13 1 9 1 9 7 9 11 11 7 9 1 9 11 11 2
16 12 9 1 12 9 14 13 0 9 1 9 2 15 13 9 2
21 12 9 0 9 14 4 13 1 0 9 1 0 9 2 15 14 4 13 1 9 2
10 11 13 1 0 9 1 0 9 3 2
25 3 15 14 15 13 1 9 1 9 1 11 11 11 7 9 1 0 15 9 2 11 2 11 11 2
19 11 14 13 3 9 1 9 1 0 9 1 0 9 1 11 1 0 9 2
26 1 9 9 1 9 7 2 11 2 15 13 1 9 1 9 9 15 14 13 12 9 9 0 0 9 2
15 9 1 9 4 13 1 9 7 3 13 1 9 10 9 2
15 0 9 1 11 1 11 1 9 13 12 9 9 0 9 2
15 13 15 1 0 9 14 15 4 13 3 12 9 9 9 2
33 13 9 2 11 9 2 1 0 9 1 10 0 9 1 11 1 0 0 9 1 9 2 9 7 9 1 9 2 13 1 0 9 2
14 0 0 9 4 13 1 9 2 13 1 11 2 11 2
15 13 15 9 1 9 1 9 1 10 9 2 0 1 11 2
15 0 13 9 1 9 2 0 1 11 2 1 12 9 9 2
18 3 1 9 2 15 13 0 9 1 0 9 2 13 0 2 13 11 2
20 15 13 11 7 0 9 1 9 14 13 0 9 2 1 14 15 13 0 9 2
11 9 13 9 1 0 0 9 1 9 1 9
20 9 15 13 3 1 0 3 3 0 9 1 9 1 9 1 0 9 1 15 2
15 9 1 11 4 13 1 9 1 9 1 12 9 1 9 2
18 9 13 9 12 9 1 9 2 7 10 9 13 7 9 1 12 9 2
13 9 1 0 9 15 13 1 9 12 9 1 9 2
13 9 15 13 3 1 14 13 0 2 13 11 11 2
29 1 9 9 1 9 3 6 15 13 1 9 1 9 1 11 2 14 1 0 9 1 9 1 11 1 9 1 11 2
20 13 3 10 9 14 13 0 9 7 11 15 13 2 13 2 11 11 11 2 2
34 3 3 13 9 1 0 9 1 11 1 0 9 2 15 14 13 0 0 9 2 3 3 13 2 16 9 4 13 1 9 2 13 9 2
35 14 15 13 11 1 3 9 13 0 9 2 15 3 13 14 13 9 1 9 2 7 9 13 7 1 10 9 2 13 2 11 11 11 2 2
21 9 1 0 9 1 0 9 2 11 2 14 4 13 1 0 0 9 1 0 9 2
13 15 13 0 9 1 9 2 15 13 1 11 3 2
17 11 13 12 9 1 9 1 2 11 2 2 15 13 1 0 9 2
22 9 1 2 0 0 9 2 11 2 9 13 14 15 13 3 1 3 2 13 1 9 2
20 9 14 15 13 10 9 2 16 3 14 13 9 1 9 1 9 1 12 9 2
49 15 13 2 11 11 2 2 2 11 9 2 2 2 11 9 2 2 2 11 11 2 2 2 11 2 2 2 11 2 11 2 2 2 11 2 2 2 11 2 2 2 0 9 2 7 2 11 2 2
18 0 9 13 12 9 9 7 13 1 0 1 0 9 1 9 1 9 2
15 0 9 13 9 1 9 0 9 7 0 15 9 1 9 2
20 1 3 13 7 0 9 1 9 1 9 2 0 1 11 2 0 0 9 2 2
12 15 13 3 7 13 9 1 9 1 0 9 2
27 12 0 9 1 9 12 9 4 13 1 0 0 9 2 11 2 1 0 12 9 1 9 2 13 3 3 2
11 0 9 1 0 9 14 13 9 1 9 2
22 15 13 3 9 11 11 1 0 9 2 1 15 13 0 15 9 7 9 1 0 9 2
18 1 9 1 9 1 9 14 15 13 3 9 1 9 1 9 1 9 2
15 0 0 9 1 9 3 14 15 13 7 13 3 1 9 2
16 3 9 15 13 1 9 2 12 1 9 7 12 1 0 9 2
12 0 12 0 9 3 14 13 10 9 1 9 2
14 10 9 13 14 13 6 3 1 12 9 2 13 9 2
10 9 13 9 1 9 7 9 1 9 2
20 1 12 0 9 9 1 9 14 15 13 1 0 9 2 0 9 7 12 9 2
10 15 14 15 13 7 13 1 0 9 2
15 11 3 13 14 4 13 0 9 1 9 1 9 1 9 2
18 9 1 0 9 1 11 11 11 6 13 9 1 10 9 2 13 11 2
26 9 14 15 13 1 0 9 2 7 9 14 15 13 1 0 9 7 0 9 2 13 0 9 1 9 2
16 9 14 13 0 9 2 7 14 15 13 1 9 2 13 9 2
18 9 1 11 1 9 11 13 9 1 9 7 15 13 0 2 13 15 2
17 9 13 9 1 0 9 7 9 1 0 9 1 9 2 13 11 2
12 3 14 15 13 7 9 1 9 7 0 9 2
16 11 13 14 15 13 1 9 1 9 7 9 2 13 1 9 2
20 9 14 13 14 13 9 1 9 1 9 7 9 7 9 1 9 1 0 9 2
7 13 9 1 2 0 9 2
9 15 4 13 1 9 1 9 3 2
27 0 9 13 14 13 0 9 1 9 1 9 2 9 11 11 2 3 16 15 14 15 13 2 13 1 11 2
33 13 9 1 0 9 1 0 0 9 7 13 1 9 2 16 9 1 11 11 1 9 1 9 13 0 2 13 9 1 11 11 11 2
24 13 0 9 1 0 9 1 9 2 7 15 4 13 7 15 13 1 9 1 9 2 13 15 2
19 9 1 0 9 15 13 1 0 9 1 9 9 2 3 7 1 0 9 2
28 15 13 9 1 9 1 9 2 9 1 9 7 9 1 9 3 1 9 1 9 2 3 7 1 9 7 9 2
10 3 15 13 1 9 14 13 0 9 2
9 9 13 3 0 9 1 10 9 2
7 9 1 9 13 9 1 11
34 9 6 13 1 9 14 13 7 10 9 11 11 2 13 11 11 2 9 1 0 9 11 11 2 7 11 11 2 9 1 9 11 11 2
21 9 1 0 9 13 14 15 13 1 11 11 2 1 14 15 13 3 13 0 15 2
39 1 1 11 11 7 11 11 13 2 1 0 13 9 7 9 1 9 11 11 2 9 1 11 11 2 9 1 11 11 7 1 11 2 3 7 0 11 11 2
21 12 12 9 4 13 1 0 12 9 1 11 2 13 0 1 11 9 1 0 9 2
9 1 15 9 6 13 3 1 11 2
15 11 13 1 9 9 1 0 9 11 11 1 9 1 11 2
9 11 13 9 1 9 1 11 7 11
23 0 9 14 13 9 2 1 15 9 1 11 7 11 13 0 2 13 0 0 9 11 11 2
6 1 9 15 13 9 2
20 3 0 9 1 0 0 9 15 13 9 1 11 7 9 15 11 11 1 11 2
13 9 1 11 11 3 13 0 9 1 0 15 9 2
15 9 1 9 1 9 14 13 1 9 7 1 0 0 9 2
28 14 15 13 0 9 1 9 1 9 1 0 9 2 7 1 10 9 14 13 0 9 1 9 2 15 13 3 2
11 9 14 13 7 3 3 9 14 13 9 2
5 9 14 13 3 9
13 15 4 13 1 10 9 1 0 9 1 0 9 2
16 1 10 9 9 1 0 0 9 14 15 13 3 1 0 9 2
10 2 11 11 2 13 9 1 9 1 11
30 0 9 1 9 1 9 13 9 1 2 11 11 2 1 9 1 12 9 1 0 9 2 11 9 2 1 9 15 3 2
10 9 15 13 14 13 12 0 0 9 2
9 13 9 1 0 9 1 2 11 2
16 0 9 1 0 0 9 4 13 3 1 9 2 11 2 3 2
13 9 1 9 1 0 0 9 1 9 13 12 9 2
16 1 15 0 11 11 15 13 3 7 1 12 9 14 4 13 2
13 0 9 15 13 3 12 9 3 2 13 9 11 2
15 0 1 9 13 2 16 9 13 7 0 9 1 0 9 2
10 15 13 9 14 15 13 1 12 9 2
5 13 9 1 0 9
21 9 1 9 1 9 13 10 9 1 9 2 1 1 1 9 9 13 1 12 9 2
29 6 4 15 13 1 9 1 0 9 2 14 14 13 1 9 1 9 1 0 9 2 13 3 1 9 1 11 11 2
17 1 9 1 0 9 3 13 14 13 9 1 9 1 11 1 9 2
11 9 1 9 3 4 13 1 9 1 9 2
9 0 9 13 9 14 13 12 9 2
20 16 9 13 9 2 15 14 15 13 1 9 1 0 9 1 0 9 0 9 2
10 9 1 11 13 11 1 9 12 9 2
43 1 9 3 1 9 1 0 9 11 7 0 11 11 4 13 12 0 9 1 11 1 9 1 9 1 9 2 0 0 9 7 0 0 9 7 0 9 1 0 7 0 9 2
6 9 11 11 3 13 2
18 9 13 2 16 9 1 0 9 13 0 1 9 2 10 9 13 9 2
22 9 1 0 9 13 12 9 11 11 2 11 11 7 11 11 2 3 7 9 11 11 2
22 12 13 9 7 9 1 11 1 9 2 11 11 11 2 7 2 11 11 11 11 2 2
16 10 0 9 13 1 9 1 9 12 9 7 12 9 0 9 2
18 1 9 4 13 9 1 9 1 11 1 15 11 11 7 9 11 11 2
16 3 0 9 11 11 3 14 4 13 2 1 14 13 9 15 2
8 0 6 13 2 16 4 13 9
17 6 4 13 9 1 9 1 9 2 3 11 13 9 2 13 9 2
21 10 9 6 4 13 7 1 2 7 1 9 11 2 11 1 9 2 0 9 2 2
25 9 1 12 9 15 13 3 9 1 9 1 9 1 9 2 11 11 2 7 9 2 0 9 2 2
16 1 15 13 9 7 15 13 1 0 9 2 16 9 13 9 2
13 10 1 9 6 13 2 16 13 0 9 1 9 2
13 0 9 15 13 2 16 4 13 1 11 14 13 11
5 3 4 13 3 2
4 13 0 9 2
37 1 0 9 15 13 0 9 7 0 9 1 9 2 11 2 12 1 9 1 9 2 11 11 2 1 9 11 11 2 0 9 1 2 11 2 2 2
22 11 13 2 16 4 13 3 1 11 2 7 6 13 9 1 15 2 7 9 1 9 2
16 3 3 2 3 3 15 13 10 9 1 11 11 7 11 11 2
5 7 15 13 3 0
8 1 15 15 4 13 1 9 2
32 0 9 1 11 13 2 16 9 1 11 6 4 13 3 9 1 0 0 9 7 1 9 1 12 9 4 13 0 9 1 9 2
32 1 15 10 10 9 1 10 9 4 13 2 7 1 9 1 9 7 3 1 0 9 7 1 15 13 3 14 15 13 9 2 2
12 15 13 10 9 1 11 1 9 1 9 9 2
11 3 11 4 13 1 9 1 9 7 9 2
18 1 9 1 2 11 2 9 1 15 13 2 16 11 6 4 13 9 2
18 1 12 0 9 4 4 13 14 13 3 9 2 7 6 15 4 13 2
12 11 13 2 16 13 3 1 0 9 1 11 2
17 3 15 13 1 12 9 7 13 15 2 15 13 1 9 1 0 9
9 9 11 13 9 1 9 1 9 2
6 9 14 15 13 3 2
16 1 0 1 2 11 2 9 1 9 13 2 16 10 9 13 2
5 13 14 15 13 9
13 15 13 10 9 1 12 9 2 11 7 0 9 2
9 3 3 15 13 10 3 0 9 2
3 7 0 2
9 7 10 9 13 14 13 7 0 2
8 9 1 9 13 9 1 9 15
25 0 9 13 2 16 13 0 9 1 9 1 0 9 3 14 4 13 9 1 11 1 9 1 11 2
10 1 10 9 11 13 0 9 1 9 2
13 7 0 9 1 9 13 0 9 1 9 1 11 2
6 3 4 15 13 15 2
6 6 13 7 0 11 2
26 1 15 13 14 15 13 1 12 9 3 2 3 0 9 2 15 15 13 1 9 1 11 13 12 9 2
24 6 15 13 3 15 14 10 2 15 14 13 1 0 9 2 14 13 1 0 9 2 13 11 2
30 3 0 2 16 3 4 13 0 2 0 7 0 9 1 9 1 9 1 9 2 3 15 13 0 0 9 2 13 9 2
23 1 15 0 9 3 13 14 15 13 0 9 1 0 0 9 7 14 15 13 9 1 9 2
19 2 9 11 2 3 14 13 9 1 9 11 11 1 0 0 9 1 11 2
11 2 6 13 14 6 15 13 9 1 9 2
16 0 2 15 13 14 15 13 2 13 14 15 13 0 0 9 2
9 15 13 0 9 1 9 1 9 2
6 9 13 14 15 13 2
8 7 3 14 15 13 0 9 2
12 13 9 1 9 1 0 9 1 10 0 9 2
10 1 10 9 10 0 9 4 13 0 2
6 15 6 13 0 9 2
4 15 13 0 2
19 16 15 15 13 2 16 15 14 13 1 11 1 11 2 15 13 14 13 2
10 15 13 1 0 9 1 10 0 9 2
15 2 14 13 14 9 1 9 1 11 1 9 1 10 9 2
8 2 9 6 13 3 1 9 2
6 9 14 13 3 0 2
18 6 13 3 14 13 2 16 1 12 9 15 14 13 1 9 7 9 2
10 15 15 13 15 14 13 1 0 9 2
21 3 4 15 13 14 13 0 7 0 9 2 13 7 0 0 9 1 11 11 11 2
39 13 2 16 0 9 2 1 15 13 10 0 9 2 13 9 1 0 9 1 9 1 9 2 15 13 0 9 1 9 1 10 9 2 10 0 7 0 9 2
9 15 13 0 9 1 11 11 11 2
9 11 11 15 13 1 2 11 2 12
12 9 13 1 0 9 3 1 9 1 12 9 2
24 0 9 1 2 11 2 12 13 2 16 9 11 4 13 0 9 1 0 9 1 9 11 11 2
18 1 0 9 3 9 13 2 1 14 13 9 1 9 1 9 1 0 2
29 14 13 9 1 10 9 1 9 2 7 15 15 13 1 9 1 0 9 2 0 9 2 13 9 1 9 11 11 2
11 0 9 13 1 9 1 11 7 0 9 2
11 3 15 13 9 1 9 1 9 1 9 2
20 13 2 3 6 13 0 9 1 11 2 9 2 9 7 0 9 2 13 11 2
13 9 11 11 4 13 1 9 1 9 1 11 11 2
15 9 13 1 0 9 0 9 2 16 11 13 9 1 11 2
17 9 13 2 16 11 4 13 1 0 9 2 3 4 13 1 9 2
10 9 13 1 9 1 9 2 11 2 2
10 1 15 4 13 3 12 9 1 9 2
19 13 4 2 16 9 13 12 9 9 9 1 0 7 0 1 9 12 9 2
15 9 15 1 9 4 13 1 0 9 1 11 1 11 3 2
28 11 13 9 14 13 1 2 11 2 7 9 1 12 12 9 14 4 13 1 9 1 9 2 13 9 11 11 2
20 1 10 9 14 4 13 9 1 9 1 9 1 0 9 1 12 9 1 9 2
6 13 3 11 1 0 9
11 12 9 14 13 9 2 13 9 1 0 9
15 0 9 7 0 1 15 9 1 11 14 4 13 3 3 2
15 9 13 14 15 13 1 9 1 0 15 9 2 13 9 2
17 0 9 1 9 14 4 13 1 12 9 11 2 9 2 13 11 2
12 3 0 9 1 9 14 15 13 1 12 9 2
14 3 0 9 1 10 9 13 1 3 0 9 7 9 2
32 11 6 13 3 0 2 16 14 13 12 0 9 2 13 7 9 1 11 11 11 1 9 1 9 1 9 2 11 2 0 9 2
7 11 15 13 1 9 1 11
17 0 9 13 3 1 0 0 9 1 11 2 13 9 1 0 9 2
28 1 9 1 11 4 13 9 1 9 1 9 1 9 2 1 9 2 1 9 2 1 9 7 1 9 1 9 2
12 14 13 0 9 2 16 6 4 13 1 9 2
30 9 1 9 1 11 11 1 0 9 11 11 2 0 9 1 11 11 11 7 11 11 13 2 16 10 9 6 4 13 2
31 9 1 9 1 0 9 1 11 13 0 7 13 14 4 13 2 13 1 9 1 9 2 15 13 1 9 0 9 10 9 2
28 1 9 0 9 11 6 4 13 10 9 1 0 9 7 13 14 6 15 13 1 9 15 2 13 9 11 11 2
7 9 1 11 13 3 0 2
23 10 9 13 14 13 9 15 1 9 1 12 9 2 13 9 1 9 2 11 2 11 11 2
8 3 13 9 3 2 13 9 2
21 1 15 3 1 9 9 1 0 9 7 9 11 11 4 13 9 1 9 1 9 2
21 1 0 9 4 13 9 15 14 13 9 1 9 1 9 1 0 9 1 9 11 2
6 10 9 15 13 3 2
25 1 15 9 1 9 7 9 1 0 9 4 13 1 9 0 9 2 1 14 14 13 9 1 9 2
7 15 4 13 3 1 9 2
16 9 13 7 9 1 0 0 9 2 15 13 0 2 13 15 2
14 3 13 14 12 9 1 9 1 0 9 2 13 15 2
6 9 13 0 9 1 9
16 15 2 9 15 7 9 15 13 0 9 1 9 1 0 11 2
12 16 4 13 2 14 15 15 13 2 13 15 2
12 6 15 4 13 10 9 2 13 1 0 11 2
11 0 9 6 4 13 1 15 2 13 15 2
11 9 13 3 0 9 1 9 1 0 9 2
10 10 9 15 13 1 12 9 1 9 2
21 4 13 3 14 13 10 9 1 0 9 9 2 15 15 13 1 9 2 13 15 2
8 1 0 9 3 15 13 0 2
22 10 0 9 15 13 7 16 4 13 9 2 15 15 13 1 10 9 2 13 9 11 2
19 3 13 9 7 1 9 2 3 9 13 3 9 7 9 7 9 7 9 2
17 3 1 12 9 1 9 3 4 13 0 15 9 2 13 3 15 2
17 9 1 9 1 9 13 1 0 9 1 9 1 0 15 1 12 9
2 11 2
28 12 9 14 2 13 2 12 9 1 12 0 9 2 1 14 13 0 9 1 10 9 7 14 13 1 10 9 2
14 12 1 10 9 4 13 1 9 11 11 1 0 9 2
11 9 13 15 14 13 1 9 1 0 9 2
26 15 14 13 9 15 1 0 9 1 0 9 2 1 0 9 1 10 9 2 16 15 6 4 13 1 9
11 9 13 1 9 1 9 11 1 0 9 2
14 1 15 2 1 9 1 9 2 0 9 13 0 9 2
12 9 13 1 9 1 9 2 0 1 0 9 2
7 9 13 14 13 9 1 11
21 0 9 1 9 11 13 1 10 9 1 12 9 7 13 9 1 9 1 0 11 2
6 15 13 3 0 9 2
35 3 3 2 13 9 1 0 9 1 0 9 2 0 3 9 1 11 13 1 11 11 7 15 13 3 14 13 14 15 13 1 9 1 9 2
8 9 13 1 2 0 9 2 2
9 3 4 13 1 9 1 10 9 2
31 16 15 3 13 14 13 3 3 9 2 1 14 6 13 15 2 15 13 3 0 2 3 14 15 13 1 9 9 1 11 2
15 11 13 9 1 9 1 9 13 0 9 2 9 9 2 2
31 1 9 11 4 13 3 1 2 9 1 9 1 9 7 9 2 0 9 1 11 2 2 1 14 15 13 2 16 13 9 2
11 9 13 9 1 9 1 11 0 1 9 2
17 1 9 1 0 0 9 15 13 2 16 9 1 11 13 12 9 2
10 12 9 13 1 9 1 11 13 11 2
7 9 13 1 11 7 11 2
14 10 1 0 9 1 0 9 11 4 13 1 0 9 2
29 0 9 13 2 16 13 0 1 9 2 0 1 9 1 9 0 9 7 1 9 1 9 1 9 1 9 1 11 2
11 0 0 9 9 1 9 4 13 1 11 2
16 13 4 9 1 0 1 9 0 9 1 0 11 2 13 11 2
10 9 1 15 13 0 9 1 0 9 2
7 0 9 1 9 13 0 2
7 13 9 1 0 2 11 2
12 9 13 0 1 9 1 0 9 1 9 1 9
2 11 2
13 3 13 9 1 9 1 0 9 1 9 1 9 2
15 13 4 0 9 2 0 1 0 2 0 9 1 0 9 2
24 16 15 13 3 2 1 9 7 9 14 13 9 1 0 9 1 0 9 2 13 9 1 9 2
33 9 1 2 11 2 7 10 9 15 13 3 1 0 9 1 9 1 0 9 7 1 0 9 2 13 11 2 3 15 1 0 9 2
19 1 9 1 9 3 1 9 4 13 3 1 9 1 9 1 2 11 2 2
14 15 13 1 9 1 9 12 9 1 0 9 1 15 2
34 0 9 1 0 9 3 13 9 1 0 9 7 9 7 1 9 2 1 9 1 9 2 13 0 9 2 0 1 0 1 0 9 9 2
2 11 2
41 0 9 0 0 9 2 11 2 13 9 1 9 1 9 1 9 1 0 9 2 11 2 7 2 11 2 2 1 0 2 11 11 11 2 7 1 0 2 11 2 2
20 13 15 9 14 13 9 1 0 9 1 12 9 1 11 7 11 1 0 11 2
22 1 9 1 9 11 15 13 1 9 1 11 7 13 2 16 13 14 15 13 1 15 2
20 11 13 7 1 9 1 0 9 1 9 1 10 0 9 2 15 14 13 9 2
18 1 0 9 1 9 1 0 9 14 13 1 12 9 0 9 9 3 2
8 11 13 1 11 1 9 1 11
21 0 0 9 13 1 0 15 9 14 13 9 15 1 11 2 9 1 9 6 13 0
2 11 2
16 13 4 7 9 1 9 1 0 9 2 11 2 2 13 11 2
14 13 14 15 13 0 9 1 9 1 11 2 13 11 2
15 3 1 9 1 0 9 1 11 14 13 7 9 1 11 2
7 11 13 9 1 9 1 11
2 11 2
28 9 13 14 13 1 0 9 1 3 0 9 1 0 9 1 11 2 13 9 1 11 11 11 2 0 1 11 2
9 11 14 4 13 1 9 11 11 2
26 11 13 11 14 15 13 1 0 9 1 0 9 7 13 0 9 1 9 1 0 11 1 10 0 9 2
13 11 14 13 1 11 1 11 10 9 2 13 11 2
34 15 13 10 9 1 9 1 9 1 9 15 3 1 9 11 11 2 15 15 13 1 0 9 2 1 14 13 1 0 0 9 1 11 2
16 1 9 11 9 1 9 1 11 7 11 14 15 13 1 9 2
8 9 3 13 9 1 0 9 2
37 1 11 2 15 13 0 9 1 0 0 9 11 2 15 13 12 9 2 1 14 13 14 13 11 1 9 15 1 11 1 9 1 9 2 13 11 2
5 10 9 13 0 9
2 11 2
17 9 13 0 9 1 0 15 9 1 9 7 9 1 0 0 9 2
5 13 1 9 1 11
19 1 3 3 6 4 13 0 9 1 11 1 9 1 11 7 9 1 9 2
2 11 2
12 1 0 9 9 14 4 13 1 0 0 9 2
20 9 2 0 1 9 2 11 2 2 14 4 13 1 0 9 1 11 11 11 2
14 2 9 13 11 14 13 1 9 1 11 2 9 9 2
8 0 9 13 9 1 9 1 11
42 3 0 9 11 11 13 2 16 11 13 14 13 0 9 1 9 1 0 9 2 16 13 3 9 1 9 1 9 1 9 1 9 1 11 1 9 1 9 2 13 11 2
13 11 15 13 1 9 1 9 15 1 11 1 9 2
32 15 15 13 2 16 14 13 14 13 1 9 1 11 2 7 1 1 0 0 9 13 0 9 7 15 13 1 9 1 0 9 2
6 0 9 1 11 13 9
2 11 2
16 0 9 1 0 0 9 1 11 11 11 13 9 2 13 11 2
36 1 9 9 1 11 1 9 15 13 3 0 2 3 3 16 3 1 12 9 1 9 1 9 0 9 1 9 1 11 15 13 9 1 0 9 2
37 1 11 0 9 1 11 4 3 13 1 9 1 0 15 9 1 9 1 9 1 9 1 9 1 0 9 2 1 15 0 9 13 0 9 11 11 2
7 9 13 7 1 10 9 2
2 11 2
16 13 15 2 16 11 2 11 2 11 7 11 13 3 1 0 9
21 15 4 13 1 9 1 9 1 11 7 3 13 9 1 3 9 2 13 9 11 2
9 1 9 15 11 13 9 1 11 2
13 12 9 13 9 1 0 9 2 13 11 1 11 2
27 0 0 9 11 11 13 2 16 0 0 0 9 4 15 13 14 13 0 9 1 9 1 9 1 0 9 2
30 9 2 15 14 4 13 0 9 2 13 0 0 9 1 0 9 1 9 14 15 13 9 1 0 9 1 0 0 9 2
17 1 0 0 9 14 4 13 7 9 1 0 1 0 9 0 9 2
10 1 9 13 9 1 1 12 9 3 2
28 9 1 9 1 0 9 11 11 13 9 1 9 2 16 1 10 9 15 13 9 1 9 1 9 1 0 9 2
14 11 11 13 12 9 9 2 0 1 9 1 9 1 9
12 3 15 13 0 9 1 0 9 1 0 9 2
13 9 13 1 12 0 9 2 1 10 9 7 11 2
16 7 3 13 0 9 1 10 0 9 2 3 0 13 7 9 2
24 1 9 7 12 9 13 9 1 9 7 9 1 9 2 3 0 0 9 7 3 0 0 9 2
27 1 0 9 0 9 15 4 13 12 9 11 7 13 1 9 15 2 9 1 9 2 1 1 12 9 11 2
16 4 13 2 16 1 11 9 14 4 13 1 9 2 11 2 2
28 1 9 1 9 9 2 11 2 13 14 13 9 1 9 1 9 1 9 1 9 2 0 1 9 1 0 9 2
23 7 1 15 11 11 15 13 1 9 1 0 9 3 1 0 9 1 0 9 1 0 9 2
44 7 1 0 9 2 0 15 1 9 1 9 1 11 2 11 11 13 1 9 1 2 9 1 9 2 9 2 7 3 15 13 7 1 9 0 9 2 1 0 9 2 11 2 2
26 1 10 9 1 9 4 13 9 1 9 1 9 1 12 9 11 2 15 4 4 13 1 9 1 11 2
24 7 3 1 0 15 9 1 3 9 1 0 9 3 6 4 13 2 16 0 11 14 15 13 2
17 1 10 9 0 9 9 2 15 13 11 1 11 2 13 3 9 2
8 1 0 9 15 3 15 13 2
9 1 11 13 2 0 2 9 1 9
13 2 3 3 9 13 10 2 9 2 1 0 9 2
21 3 9 15 13 1 0 9 1 2 0 9 2 2 3 0 1 10 9 1 9 2
24 7 3 13 3 14 15 13 9 1 0 9 9 2 1 1 1 15 15 13 0 9 1 11 2
19 15 14 4 13 1 0 9 1 0 9 2 9 1 0 9 7 0 9 2
29 1 9 1 11 7 9 1 9 1 9 10 9 13 0 9 2 7 3 1 15 3 3 14 14 15 13 1 9 2
15 7 3 1 0 9 9 13 9 1 9 7 9 1 9 2
24 1 1 0 9 1 11 1 10 9 3 9 13 14 15 13 1 0 9 2 7 9 4 13 2
17 1 9 2 9 1 0 9 1 0 11 15 13 14 13 0 9 2
13 1 0 9 0 9 13 3 0 9 1 9 9 2
19 3 14 15 13 1 12 9 1 9 1 0 9 1 9 1 9 1 9 2
6 11 14 13 9 1 11
25 11 11 4 13 0 9 1 0 15 9 14 13 1 9 1 9 2 16 6 15 13 1 0 9 2
10 15 13 11 11 2 1 14 4 13 2
34 1 9 1 0 9 1 11 7 9 1 11 1 0 9 3 11 15 13 7 1 0 9 1 9 7 9 1 0 9 1 9 1 11 2
9 3 9 13 14 15 13 1 9 2
8 11 11 13 1 12 9 1 9
13 1 0 15 0 9 9 13 9 1 0 9 1 11
7 11 11 11 13 3 3 2
13 15 13 11 11 2 9 1 9 2 11 11 2 2
20 1 11 15 13 1 9 7 9 2 9 1 15 4 13 1 9 1 0 9 2
10 9 1 9 13 1 12 9 0 9 2
18 0 9 11 11 11 15 13 1 11 2 1 14 13 9 15 1 9 2
11 13 2 9 1 11 2 3 1 11 11 2
19 15 4 13 1 0 9 2 0 9 2 1 11 7 13 0 9 1 9 2
13 1 9 1 9 9 14 4 13 1 9 1 9 2
7 9 13 9 1 9 1 9
27 1 9 15 13 2 16 3 13 1 9 9 2 10 9 15 13 1 0 2 1 9 7 9 1 0 9 2
16 9 7 9 1 9 2 15 15 13 1 9 2 13 1 1 9
8 2 11 11 2 3 13 1 9
16 9 1 2 11 11 2 3 13 9 12 1 11 2 13 11 2
13 11 4 13 9 1 0 9 1 0 15 9 11 11
15 13 15 3 15 13 1 9 7 15 13 1 10 0 9 2
15 1 12 9 9 1 11 13 9 7 9 1 9 7 9 2
7 0 9 13 1 10 9 2
12 13 15 2 16 3 3 11 11 13 0 9 2
12 9 1 0 9 13 3 9 15 7 15 13 2
7 3 11 3 13 11 9 2
27 3 7 1 0 9 15 13 9 1 9 2 11 11 2 7 9 1 0 0 9 1 9 7 9 1 11 2
20 0 9 1 9 1 9 13 1 0 9 1 9 1 0 9 1 11 11 11 2
13 1 0 9 13 9 15 1 9 7 3 13 9 2
23 1 0 9 3 13 9 1 0 9 1 0 9 2 7 1 0 9 13 1 2 11 2 2
31 13 1 9 1 9 11 11 7 3 13 1 9 1 10 9 3 1 9 1 0 9 1 2 11 2 1 11 1 0 9 2
12 1 9 13 7 1 9 1 2 11 11 2 2
27 3 1 10 0 9 1 0 9 13 1 12 0 9 2 1 9 2 1 9 7 1 9 1 9 1 11 2
33 1 0 9 11 13 9 1 0 9 2 16 9 1 0 9 4 13 1 2 10 9 2 1 11 11 2 7 9 13 1 0 11 2
30 1 0 9 4 13 1 9 1 0 9 1 9 2 11 2 1 11 7 3 9 15 13 1 0 9 1 9 7 9 2
7 15 13 9 1 9 3 2
12 3 3 13 14 13 9 15 1 9 1 9 2
17 15 13 9 1 9 1 0 9 7 0 9 1 0 9 7 9 2
9 9 11 11 13 10 9 1 11 2
12 3 1 9 11 15 13 1 3 1 12 9 2
9 9 13 0 15 9 11 11 11 2
12 9 1 9 11 11 15 13 2 0 9 2 2
17 1 9 9 13 1 11 7 1 11 2 3 0 9 13 0 9 2
21 2 9 1 0 2 14 13 11 1 9 1 0 0 9 1 0 9 2 11 2 2
20 9 1 11 11 13 1 0 9 10 9 7 3 4 13 1 1 12 9 9 2
13 9 3 4 13 1 0 9 1 0 9 1 11 2
9 9 14 15 13 1 9 0 9 2
6 0 9 15 13 1 11
10 1 9 13 12 9 1 10 0 9 2
11 9 1 9 13 1 9 1 11 2 11 2
11 0 13 12 9 2 0 1 9 7 9 2
6 9 13 0 9 7 9
38 10 9 11 11 13 12 0 9 2 15 13 9 1 9 1 9 1 11 1 0 9 1 0 9 1 10 9 2 9 7 9 15 1 9 2 11 2 2
24 0 9 13 10 0 9 1 0 9 2 1 11 14 15 13 1 0 1 15 9 1 0 9 2
13 1 15 4 13 7 0 9 1 9 1 9 15 2
14 1 15 11 13 0 15 9 1 9 1 9 7 9 2
11 15 3 4 13 9 15 7 4 13 9 2
5 10 0 0 11 2
17 14 4 13 14 13 2 16 9 13 3 7 11 13 3 10 9 2
17 10 9 13 0 9 9 1 9 1 11 2 15 13 1 11 11 2
13 0 9 13 7 0 9 7 1 9 1 0 11 2
7 1 9 13 1 0 9 2
4 13 3 3 2
27 1 9 0 9 1 0 9 15 13 11 2 7 11 15 13 1 0 15 9 1 11 11 2 9 1 11 2
4 10 0 9 2
5 9 13 3 0 2
4 6 13 0 2
4 13 9 1 11
23 0 9 13 1 11 1 9 14 15 13 0 9 1 11 1 0 7 0 9 2 13 11 2
10 13 12 9 2 13 4 12 9 9 2
12 0 9 14 13 3 0 1 9 1 0 9 2
16 3 9 4 13 1 12 9 9 2 9 4 13 1 12 9 2
9 0 9 13 3 1 9 7 9 2
16 9 15 13 1 12 12 0 9 2 13 9 1 9 7 9 2
18 0 9 1 9 13 12 0 9 1 9 2 0 9 2 9 1 9 2
30 9 1 9 13 1 9 1 9 1 0 9 2 1 15 13 9 1 11 7 11 3 3 11 15 13 1 9 1 9 2
30 13 4 7 9 1 9 0 9 2 15 13 0 9 2 2 9 2 9 2 2 9 1 0 11 2 0 1 0 9 2
17 0 9 1 9 13 9 1 9 1 11 2 11 2 1 0 9 2
16 6 4 13 7 12 0 0 9 1 0 9 2 0 7 0 2
19 13 4 7 9 1 9 1 9 1 11 11 1 11 11 2 0 1 9 2
9 10 0 9 15 13 1 0 9 2
24 2 0 9 2 1 11 7 2 9 3 2 1 11 11 13 0 9 1 0 9 1 0 9 2
14 9 1 10 9 4 13 1 9 2 15 4 15 13 2
16 1 0 9 0 9 2 11 11 2 3 13 9 15 1 9 2
29 3 0 0 9 14 15 13 1 9 1 0 9 2 1 15 14 13 9 7 9 1 9 15 2 13 11 11 11 2
24 9 1 9 1 9 13 9 1 0 1 0 9 9 1 12 9 2 15 4 13 1 9 9 2
17 3 9 4 13 9 2 15 3 4 13 1 0 9 1 12 9 2
17 13 9 9 1 0 9 2 11 11 2 14 4 13 1 0 9 2
21 11 11 11 4 13 1 0 9 0 9 1 11 2 11 2 7 13 1 0 9 2
39 1 9 15 4 13 0 9 1 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2
14 3 15 13 9 1 11 11 2 3 16 9 13 15 2
16 9 13 3 0 2 1 14 4 13 1 10 9 1 0 9 2
18 1 9 1 0 0 9 9 1 0 0 9 13 1 12 7 12 9 2
32 1 9 9 11 11 13 1 11 3 1 12 9 9 7 9 2 1 15 4 13 2 13 1 9 2 3 15 4 13 0 9 2
5 9 15 13 1 9
29 0 0 9 13 2 16 4 13 9 2 15 15 13 1 9 7 9 15 13 12 9 1 12 9 2 13 11 11 2
19 0 9 1 9 15 13 1 0 9 2 15 15 13 1 0 9 1 9 2
16 9 14 13 14 13 9 1 10 9 1 9 7 14 15 13 2
18 0 9 4 13 1 2 11 11 11 11 2 1 11 2 9 0 11 2
7 0 0 9 13 1 9 2
18 1 9 15 4 13 0 9 2 0 1 0 9 1 11 12 11 11 2
19 9 13 3 0 0 9 1 9 2 0 1 12 9 9 2 13 0 9 2
16 1 11 11 2 9 1 9 2 9 13 1 0 9 11 11 2
11 0 9 4 13 1 12 9 3 1 11 2
6 9 1 0 9 4 13
13 0 9 11 11 13 9 1 0 9 2 13 11 2
34 1 0 9 2 15 15 13 1 11 2 11 11 13 0 9 1 9 2 16 1 9 1 10 9 9 13 14 13 3 3 9 1 9 2
38 16 6 15 13 9 1 9 7 6 13 0 9 1 9 2 14 13 9 1 0 9 2 13 1 9 1 9 0 9 1 9 1 9 1 9 11 11 2
21 1 15 13 14 15 13 9 1 9 1 9 1 9 1 10 9 2 13 1 11 2
9 6 13 1 9 2 1 1 15 13
29 0 0 7 0 9 2 15 3 13 1 15 2 14 13 1 0 9 2 13 9 1 0 9 1 0 9 9 11 11
13 2 13 14 2 9 2 1 0 9 2 9 9 2
3 2 6 2
14 1 9 10 9 0 9 13 9 1 9 1 0 9 2
17 1 0 9 0 9 3 14 13 3 0 7 13 14 13 0 9 2
7 2 13 2 16 13 0 2
9 1 9 2 1 15 6 15 13 2
13 1 15 10 9 13 14 13 1 9 1 0 9 2
10 6 13 1 9 2 1 1 15 13 2
3 2 15 2
22 2 3 0 0 7 0 9 1 9 2 15 6 4 13 0 15 9 2 13 1 15 2
8 3 15 14 13 1 0 9 2
10 14 13 3 9 0 9 2 0 9 2
9 6 13 0 9 1 0 15 9 2
7 12 13 1 9 7 9 2
12 12 13 1 0 9 2 12 13 1 0 9 2
14 12 13 1 9 1 0 9 1 9 2 1 0 9 2
8 1 0 9 6 13 0 9 2
9 2 13 14 3 0 9 1 15 2
9 2 13 14 3 0 9 1 15 2
3 7 9 2
3 2 6 2
17 1 0 1 0 9 15 15 13 14 15 13 1 12 9 1 9 2
18 2 13 2 16 13 9 2 15 14 6 13 14 15 13 1 0 9 2
15 13 9 1 0 9 2 1 14 15 13 1 9 7 9 2
18 1 15 13 9 1 12 9 2 1 15 1 15 13 14 15 13 9 2
6 13 15 9 1 9 2
14 2 15 13 2 13 14 13 1 0 9 1 0 9 2
12 3 12 10 9 7 9 3 13 1 10 9 2
16 2 1 0 0 9 14 13 9 1 9 1 12 12 9 9 2
7 0 9 13 12 9 9 2
30 0 15 9 1 0 9 1 9 13 0 9 1 11 2 9 2 11 2 1 9 1 11 2 9 1 11 2 11 2 2
33 1 9 1 9 15 13 14 13 3 12 12 9 0 9 1 9 11 2 11 2 11 2 11 2 0 11 2 11 7 11 2 11 2
9 9 2 11 2 13 1 9 1 9
16 9 1 0 9 11 11 14 13 9 2 13 0 0 9 11 11
6 3 13 9 1 9 2
15 2 1 9 1 9 9 7 0 9 14 4 13 1 9 2
26 13 2 16 0 15 9 14 4 13 1 9 1 9 1 9 1 9 14 13 0 0 9 1 0 9 2
20 7 13 9 1 0 9 2 15 13 2 16 13 3 6 0 9 2 7 9 2
14 2 16 15 13 9 1 9 2 15 13 14 15 13 2
15 13 4 3 9 1 9 1 9 7 15 3 14 13 9 2
7 2 13 9 2 11 2 2
9 2 1 0 9 15 13 1 15 2
11 13 0 9 1 0 9 1 9 1 9 2
14 1 0 9 13 0 0 0 9 7 15 13 1 9 2
12 11 13 9 2 15 13 0 1 0 0 9 2
21 2 1 9 2 11 2 15 13 2 16 9 1 0 9 4 13 1 9 1 11 2
18 0 9 1 0 9 4 13 1 9 2 9 2 12 9 0 9 2 2
16 2 9 2 0 1 9 2 13 2 16 9 1 9 13 0 2
20 2 16 3 13 10 9 2 15 3 13 1 9 2 15 4 13 3 1 9 2
28 13 2 16 10 9 4 13 1 9 2 16 4 13 3 9 1 9 1 0 9 7 3 14 15 13 7 9 2
17 7 10 9 6 4 13 1 0 9 1 9 7 1 0 0 9 2
12 2 3 0 9 13 14 13 3 1 10 9 2
22 3 3 13 9 1 9 1 12 9 2 1 0 0 9 7 0 9 0 9 7 9 2
19 10 1 9 6 13 14 4 13 2 1 14 15 13 1 15 0 0 9 2
7 2 1 10 14 13 9 2
9 9 13 14 15 13 9 1 9 2
8 11 7 11 13 0 9 1 11
25 6 13 0 9 14 13 1 0 9 1 0 9 2 13 11 11 2 9 1 0 9 1 9 1 11
10 3 7 10 0 0 9 13 0 9 2
14 15 3 13 9 1 11 7 0 0 9 1 0 11 2
25 15 13 0 9 7 3 13 14 13 0 9 1 0 9 1 9 1 9 2 9 1 9 7 3 2
16 2 1 10 0 9 3 13 9 1 0 9 1 9 1 11 2
14 7 0 0 9 13 3 9 9 2 16 6 15 13 2
8 13 1 9 1 9 11 11 2
10 15 15 13 9 1 0 7 0 9 2
15 7 6 13 9 1 9 14 13 1 0 9 1 0 9 2
7 15 13 7 1 0 9 2
12 14 2 13 15 2 0 14 6 13 0 9 2
7 15 13 3 0 1 9 2
8 2 3 15 13 9 1 11 2
19 15 15 13 1 0 9 2 1 9 2 0 9 2 9 2 9 7 3 2
18 7 3 9 13 14 13 0 9 2 15 15 13 1 9 1 0 9 2
29 2 0 2 15 9 13 9 14 13 2 13 14 13 0 9 1 9 2 9 7 9 1 9 1 0 0 0 9 2
12 7 7 10 9 3 13 14 4 13 1 9 2
14 7 1 9 1 0 9 9 13 1 9 1 0 9 2
9 1 16 6 13 9 1 0 9 2
16 7 10 9 13 14 13 9 1 10 9 1 0 9 1 9 2
20 13 15 2 16 1 0 9 13 0 9 2 15 13 1 0 9 1 0 9 2
16 2 15 13 9 1 10 0 9 2 1 15 13 9 7 9 2
20 3 15 13 1 0 9 1 9 11 2 15 13 9 1 9 1 0 0 9 2
11 2 6 2 9 1 9 11 13 3 0 2
12 6 15 13 1 9 1 9 1 9 7 9 2
13 3 10 9 13 3 0 2 3 1 11 7 11 2
11 2 13 14 11 14 4 13 1 0 9 2
8 16 11 13 3 1 15 14 2
8 0 9 13 9 15 2 11 2
12 3 9 15 13 1 9 14 15 13 1 9 2
5 11 15 13 0 9
14 3 13 3 14 15 13 10 9 1 0 9 13 0 2
9 11 11 2 9 1 0 7 0 9
21 0 9 1 0 9 1 0 9 13 3 0 1 10 9 2 0 1 9 1 11 2
24 7 1 10 0 9 15 13 10 0 9 1 9 1 0 1 9 1 11 9 1 9 7 9 2
15 9 1 9 13 1 9 1 0 9 2 0 3 1 11 2
19 3 15 13 0 9 2 15 3 13 9 1 0 9 1 2 0 9 2 2
15 9 2 15 13 1 10 9 14 13 7 13 9 1 9 2
10 15 3 13 0 0 9 1 0 9 2
14 3 3 3 15 13 0 9 2 0 1 0 0 9 2
6 7 15 13 0 9 2
10 1 9 9 1 10 9 13 0 9 2
20 0 9 6 13 14 13 0 9 1 9 1 0 9 1 9 15 1 12 9 2
13 1 10 9 2 13 9 2 15 13 1 0 9 2
19 15 13 9 1 0 9 7 10 2 15 13 3 0 2 7 13 1 11 2
12 1 3 2 11 11 2 2 15 13 0 9 2
8 1 0 9 2 13 0 9 2
5 10 9 13 0 2
11 9 1 10 12 9 13 9 1 0 9 2
18 3 15 13 2 15 15 13 3 0 1 9 1 9 2 9 7 3 2
9 7 9 15 6 13 1 10 9 2
8 3 1 9 9 15 13 3 2
6 14 13 3 0 9 2
10 1 9 15 13 1 12 9 0 9 2
31 0 3 2 1 9 1 12 9 7 9 9 13 9 1 9 7 9 2 9 7 9 1 9 7 9 7 9 1 0 9 2
9 7 15 6 13 0 9 1 9 2
13 1 10 9 9 1 0 9 6 13 14 4 13 2
20 3 16 1 9 9 1 10 9 7 9 6 13 1 0 9 7 9 1 11 2
18 1 9 9 1 0 0 9 1 11 13 1 0 9 1 9 1 9 2
24 10 10 9 2 15 13 1 9 2 4 13 14 13 9 1 9 2 11 2 1 0 0 9 2
22 10 9 3 15 13 1 3 0 9 1 9 2 9 2 0 9 1 0 9 7 3 2
9 14 13 9 1 10 0 0 9 2
16 13 3 12 9 2 15 13 9 1 9 1 9 1 9 15 2
10 9 1 9 15 13 3 3 3 0 2
8 13 9 2 15 14 13 9 2
28 7 0 13 14 15 13 1 9 1 10 10 9 2 15 3 4 13 14 13 1 0 9 1 9 7 0 9 2
7 0 13 9 1 9 1 9
28 10 0 9 13 3 9 1 9 1 9 1 0 9 2 3 7 9 1 0 9 1 9 2 0 1 0 9 2
10 9 1 10 9 13 0 9 1 9 2
17 15 13 7 3 0 9 1 9 1 9 1 9 9 1 0 9 2
19 13 13 9 1 9 13 9 14 4 13 9 1 10 0 7 0 0 9 2
28 15 13 13 14 15 13 1 9 1 9 15 2 7 1 9 14 15 13 1 0 9 1 9 7 0 0 9 2
27 9 1 10 9 1 9 13 9 3 1 0 7 0 9 1 0 9 7 9 15 1 10 0 9 1 9 2
3 11 15 13
12 1 0 9 1 11 4 13 0 0 0 9 2
13 3 15 13 1 9 1 11 1 9 1 11 11 2
20 10 9 13 11 11 2 11 11 7 11 11 2 7 1 9 4 13 11 11 2
6 1 0 9 13 11 2
13 1 9 1 0 9 9 1 0 9 13 3 0 2
12 0 0 9 13 9 0 9 1 9 1 9 2
34 10 0 9 2 11 11 2 3 0 1 9 15 1 11 1 9 1 0 9 7 3 1 9 11 0 2 15 13 3 1 9 1 9 2
18 10 9 13 3 0 9 1 9 2 7 1 15 15 13 9 1 11 2
5 9 13 0 1 9
8 9 1 0 9 6 15 13 2
11 14 15 13 2 16 6 15 13 3 9 2
10 9 13 0 9 14 15 13 0 9 2
13 3 15 13 1 0 9 2 13 14 13 7 9 2
7 9 3 13 1 0 9 2
5 0 9 13 0 2
5 0 13 9 1 9
21 13 15 2 16 9 1 9 2 9 1 0 9 2 14 13 9 1 9 1 9 2
28 9 14 15 13 1 9 1 0 9 7 14 13 10 9 2 7 15 15 13 1 9 1 9 9 14 4 13 2
15 15 3 3 6 4 13 1 9 1 9 2 15 13 0 2
5 9 13 9 1 0
8 0 9 13 9 1 0 9 2
13 9 13 0 7 15 6 13 9 14 13 0 9 2
8 13 10 0 9 1 9 3 2
14 2 13 0 11 11 2 0 9 1 2 11 2 11 2
9 9 3 4 4 13 1 10 9 2
12 1 9 1 0 9 1 0 9 13 0 9 2
15 9 4 15 13 9 1 9 2 7 15 0 13 1 9 2
10 9 14 15 13 9 4 13 7 9 2
10 15 7 14 15 13 2 9 13 0 2
14 10 9 3 12 9 13 1 9 2 13 9 1 9 2
15 15 13 9 1 0 15 9 0 1 0 9 1 9 15 2
8 3 3 13 9 1 0 9 2
18 1 12 9 0 9 9 13 1 12 9 1 0 0 9 1 12 9 2
9 9 13 2 3 15 13 0 9 2
6 0 9 13 0 15 9
16 1 14 13 12 9 2 0 9 3 13 9 1 9 1 9 2
6 3 9 13 9 0 2
18 1 9 1 9 11 11 11 9 1 0 9 1 9 1 9 13 0 2
11 3 12 9 9 13 2 16 0 9 13 2
4 9 13 0 2
10 9 1 9 13 0 7 6 13 15 2
18 1 9 11 13 9 1 0 0 9 2 11 2 1 9 1 0 9 2
13 9 3 3 15 13 1 9 1 9 7 15 13 2
12 3 7 14 15 13 2 15 13 1 0 9 2
11 1 9 2 9 7 9 9 13 1 3 2
16 13 3 0 9 2 7 10 1 9 15 13 7 6 15 13 2
11 6 13 14 13 15 2 13 0 9 1 9
8 15 3 4 13 1 0 9 2
5 0 9 13 9 2
15 0 0 9 1 9 3 13 9 7 15 3 13 1 9 2
9 0 9 4 15 13 1 0 9 2
8 7 9 13 2 7 13 3 2
14 0 13 10 2 15 15 13 2 7 1 9 14 13 2
5 14 13 9 1 9
12 1 12 9 13 1 11 14 15 13 1 9 2
9 7 0 9 1 0 9 15 13 2
18 13 2 16 10 1 0 9 13 1 9 1 9 2 0 9 7 9 2
9 9 1 15 13 0 7 13 1 9
15 0 9 13 0 9 2 15 3 6 13 14 13 9 15 2
21 9 15 4 13 2 7 15 13 1 9 2 3 1 12 9 9 13 14 15 13 2
8 1 10 0 9 9 13 0 2
7 16 13 3 2 14 15 13
11 0 9 13 7 9 1 0 9 11 11 2
15 15 13 1 12 0 9 2 16 3 9 1 15 4 13 2
11 1 9 1 9 9 3 13 9 1 9 2
19 3 1 0 12 9 1 10 9 4 13 12 9 1 0 9 12 12 9 2
12 12 0 9 4 13 1 9 15 1 0 9 2
16 3 13 9 1 0 9 2 3 0 9 13 9 1 0 9 2
12 0 0 9 13 0 9 1 0 9 1 11 2
8 9 13 3 2 7 3 15 13
7 2 13 4 9 1 9 2
7 13 7 9 1 11 1 11
18 9 14 4 13 1 9 1 9 1 11 2 15 15 13 7 1 0 9
15 1 9 15 9 13 9 1 9 7 13 9 1 0 9 2
27 11 13 2 16 14 13 9 15 1 9 1 9 2 3 1 0 9 13 14 13 9 9 0 9 1 11 2
13 9 13 3 7 0 9 1 11 1 11 11 11 2
19 1 11 0 9 1 9 15 14 13 0 9 1 15 13 0 15 0 9 2
13 3 3 6 13 3 15 14 4 13 1 9 9 2
14 1 0 9 1 9 1 11 15 13 12 9 1 11 2
11 13 4 7 9 1 10 1 9 1 9 2
9 11 11 13 14 13 9 1 9 2
9 11 15 13 1 9 1 2 11 2
17 1 11 9 1 9 1 0 9 4 13 1 9 1 11 1 9 2
11 1 10 9 3 4 13 0 9 1 15 2
16 1 9 1 11 9 14 13 9 2 1 14 6 15 13 9 2
9 13 9 1 11 2 13 3 11 2
5 11 13 9 1 11
24 9 1 0 9 3 13 3 14 13 0 9 1 0 1 9 15 9 1 2 11 2 11 11 2
16 9 1 10 9 13 9 15 1 11 11 11 1 9 1 9 2
21 11 13 0 9 2 1 14 13 0 2 7 4 15 13 14 13 9 2 13 11 2
14 15 6 13 14 15 13 2 3 9 15 13 1 9 2
21 11 11 4 13 11 11 14 13 0 9 1 9 1 11 11 2 13 2 11 2 2
10 9 13 3 0 2 13 3 0 9 2
14 3 15 4 13 7 1 11 11 1 9 15 1 9 2
19 9 1 9 1 9 1 11 13 0 15 9 1 0 9 1 11 1 9 2
21 1 9 15 13 9 1 11 1 11 2 9 1 11 7 9 1 11 1 0 9 2
13 0 15 9 1 0 9 14 13 0 0 0 9 2
24 1 9 1 0 0 9 1 9 1 9 4 13 7 9 1 11 11 7 11 11 2 13 0 2
24 11 3 13 2 16 11 13 14 4 13 2 3 16 13 0 1 9 15 1 9 1 0 9 2
7 9 1 11 4 4 13 2
22 9 1 11 13 9 1 11 11 1 0 9 1 9 1 0 9 1 9 1 11 11 2
21 11 11 7 11 11 11 13 9 1 11 1 9 1 0 9 1 9 1 11 11 2
10 0 9 1 11 13 1 12 9 3 2
15 9 1 15 13 7 11 11 2 7 1 12 9 13 9 2
17 1 12 1 2 11 2 12 13 11 11 2 11 11 7 11 11 2
10 11 11 3 6 15 13 3 1 9 2
5 11 11 13 1 11
15 1 9 13 9 1 0 9 2 0 1 9 2 13 15 2
20 0 9 6 15 4 13 3 7 1 0 1 0 9 9 1 0 9 1 11 2
23 9 1 0 9 1 0 9 1 0 9 15 13 1 9 1 0 9 0 9 9 11 11 2
15 3 4 13 1 0 7 9 15 1 9 1 11 1 9 2
25 14 13 9 11 11 3 14 13 0 9 1 0 9 2 13 3 7 9 1 11 1 9 11 11 2
5 0 13 3 0 9
22 1 9 1 11 11 1 0 9 0 9 11 13 14 13 11 3 1 0 9 1 11 2
9 15 13 0 9 2 13 11 11 2
17 9 1 11 13 0 1 11 9 1 12 0 9 2 0 1 9 2
18 1 9 15 13 9 2 16 1 9 13 9 1 0 9 2 11 2 2
14 3 9 1 9 1 11 11 11 13 9 1 0 9 2
16 15 6 13 10 7 14 13 9 1 9 1 11 2 13 15 2
6 11 15 13 1 9 15
29 15 13 2 16 9 1 9 1 11 7 11 13 3 0 2 1 14 15 13 9 1 9 2 3 0 9 13 0 2
34 3 1 15 13 2 16 9 1 0 9 7 9 1 9 1 9 1 11 13 9 2 3 16 13 0 7 0 2 13 1 9 11 11 2
4 9 13 0 9
10 14 13 0 9 1 10 0 0 9 2
20 15 13 9 1 0 9 1 15 1 9 1 9 11 11 3 1 0 0 9 2
25 1 0 9 9 1 11 2 11 2 9 1 9 7 9 1 0 9 1 9 13 0 1 9 15 2
14 3 0 9 13 1 12 9 1 9 15 1 0 9 2
25 9 1 0 9 11 11 13 2 16 9 13 3 14 13 0 9 1 9 1 9 15 1 0 9 2
7 11 13 9 1 11 7 11
12 11 13 0 9 2 13 9 1 11 11 11 2
19 12 4 13 9 1 9 15 1 11 2 13 1 9 1 2 11 2 12 2
9 13 15 1 0 9 1 9 1 9
24 9 13 1 9 1 0 9 2 7 1 9 1 9 2 1 15 15 14 4 13 1 0 9 2
22 1 10 9 14 15 13 1 9 1 0 9 1 0 9 1 9 1 9 1 0 9 2
10 1 9 1 10 9 3 13 0 9 2
13 15 13 14 13 1 0 7 0 9 1 10 9 2
22 3 14 15 13 9 14 13 9 1 0 9 1 11 2 15 14 15 13 1 12 9 2
19 1 11 3 7 3 13 9 1 9 1 9 1 9 15 1 9 1 9 2
6 3 13 14 15 13 9
16 10 9 1 9 13 14 13 0 9 3 1 0 9 1 9 2
9 14 15 13 9 3 13 3 0 2
6 15 13 3 0 9 2
12 4 13 0 2 16 13 1 9 1 11 11 2
3 13 1 11
17 2 9 11 13 2 16 9 1 9 13 1 0 0 9 1 11 2
19 10 9 13 1 9 1 11 7 15 13 7 4 13 2 16 15 14 13 2
19 2 3 14 13 9 1 9 1 0 9 1 11 1 9 1 9 9 11 2
21 2 15 3 13 2 16 6 13 14 13 1 9 11 2 3 13 1 15 3 3 2
14 3 9 1 10 9 13 3 0 9 1 9 1 15 2
16 9 11 3 6 13 2 6 13 14 13 14 13 1 10 9 2
23 1 0 9 4 13 1 10 0 9 1 0 15 3 0 0 9 1 9 1 9 1 9 2
26 9 1 9 11 13 9 1 12 9 1 9 2 1 12 0 9 1 9 2 7 6 13 9 1 9 2
13 0 9 1 9 1 9 13 1 0 9 1 11 2
5 13 9 1 9 2
12 3 1 0 9 3 13 2 16 13 10 9 2
8 15 6 13 0 1 10 9 2
17 9 13 2 16 4 13 3 9 7 1 11 2 7 1 0 9 2
16 11 13 9 1 9 1 9 2 15 13 1 9 1 12 9 2
12 9 1 10 9 3 13 1 9 1 12 9 2
10 1 12 9 15 13 3 9 12 9 2
10 15 2 13 15 2 3 6 13 0 2
8 15 13 9 1 9 1 11 2
12 7 0 9 13 9 2 9 7 9 1 11 2
7 13 9 14 13 0 15 9
7 11 11 2 9 1 0 9
33 9 1 9 1 0 11 13 14 15 13 1 0 9 1 9 1 0 9 1 11 7 1 9 15 1 0 9 1 9 1 0 9 2
16 15 13 0 9 2 15 4 13 14 15 13 1 9 1 9 2
8 3 10 9 4 13 1 9 2
4 11 13 0 9
23 3 13 14 4 13 9 1 11 11 1 9 1 9 1 0 9 2 3 1 9 1 9 2
6 9 1 9 13 0 9
24 2 3 13 9 1 9 1 0 9 1 0 9 11 11 2 13 15 14 13 3 10 0 9 2
15 3 3 15 13 2 16 15 3 3 13 0 9 1 9 2
21 13 0 9 2 1 14 15 13 1 9 2 1 15 6 13 0 2 16 13 9 2
7 2 6 2 13 1 9 2
21 1 9 15 1 15 15 13 2 16 10 9 1 10 9 3 6 13 0 1 11 2
7 2 9 15 13 3 0 2
8 2 6 2 3 13 0 9 2
13 2 14 13 14 11 2 16 13 1 9 1 9 2
13 9 15 1 9 1 9 14 13 0 9 1 11 2
15 3 3 13 7 9 2 7 9 14 13 3 1 10 9 2
7 9 1 9 13 14 15 13
6 11 11 2 9 1 9
6 3 13 9 1 11 0
9 11 11 2 9 1 0 9 7 9
12 15 13 3 9 1 0 9 1 9 11 11 2
15 0 15 9 14 13 3 9 2 16 4 13 1 0 9 2
17 0 9 14 13 1 0 9 7 9 2 0 9 7 9 1 9 2
23 15 4 15 13 3 0 0 9 2 9 1 9 7 0 9 1 9 15 1 0 0 9 2
23 3 13 9 1 1 12 9 2 15 13 2 0 9 2 2 13 9 1 9 9 11 11 2
23 1 14 13 0 9 2 9 13 14 13 3 12 9 2 13 7 9 1 9 9 11 11 2
26 9 2 15 13 1 0 9 7 6 13 14 13 12 9 2 14 13 9 15 7 14 14 13 0 9 2
6 13 9 1 9 1 9
17 1 10 9 4 15 13 0 9 1 9 1 9 2 9 7 0 2
24 9 7 9 1 0 9 14 13 14 15 13 3 1 9 1 9 11 2 1 0 9 1 9 2
7 12 13 1 0 9 1 11
13 9 13 12 9 1 9 2 9 11 13 0 1 11
2 11 2
23 12 9 13 1 0 9 7 0 9 1 11 2 11 2 11 2 11 7 11 2 13 9 2
15 1 0 15 9 13 9 1 9 2 15 15 13 1 9 2
14 3 12 9 13 1 0 9 1 9 1 11 7 11 2
8 1 11 0 9 13 12 9 2
14 1 9 9 1 11 13 12 9 1 9 2 13 11 2
10 1 9 3 4 13 9 1 0 9 2
18 1 0 11 13 0 9 2 3 9 7 0 9 13 9 1 0 9 2
11 1 11 13 9 2 1 9 15 13 9 2
8 9 1 11 7 11 4 13 2
17 12 9 1 9 9 6 13 14 13 1 11 7 13 1 0 9 2
14 1 12 9 1 11 15 13 0 9 1 9 7 9 2
10 9 13 9 1 9 1 11 7 11 2
5 0 9 13 1 9
15 9 14 13 2 0 9 2 1 9 1 0 9 1 11 11
3 11 11 2
31 0 9 13 3 3 14 13 9 1 9 1 9 2 13 9 1 9 1 0 9 1 11 9 11 11 2 0 1 0 9 2
16 9 6 13 3 9 1 0 0 9 1 0 9 2 13 9 2
9 15 13 9 1 9 1 0 9 2
19 15 13 3 0 9 11 11 1 9 1 9 1 9 9 11 2 13 11 2
7 11 13 1 0 9 1 11
2 11 2
13 0 9 11 11 4 13 1 0 9 1 11 3 2
12 9 1 11 15 13 1 0 9 1 0 9 2
10 15 4 13 3 1 0 9 1 9 2
20 9 1 9 11 11 14 13 14 13 9 1 9 1 9 14 13 9 1 9 2
5 3 9 3 13 2
20 11 13 9 1 9 1 9 15 14 15 13 1 9 1 9 1 9 1 9 2
9 9 11 13 2 16 14 13 9 2
7 11 7 11 11 13 11 11
18 9 3 13 0 1 9 1 11 9 2 0 1 11 1 9 1 9 15
16 11 11 11 11 2 2 11 11 11 2 2 3 1 2 11 2
16 1 9 1 2 11 11 11 2 4 13 9 15 2 11 2 2
8 3 9 15 13 2 11 2 2
17 1 9 16 13 2 15 13 0 9 2 7 1 0 9 13 9 2
4 15 6 13 2
23 15 15 13 0 9 14 13 1 9 7 14 15 13 2 16 4 13 14 15 13 0 9 2
20 9 13 9 9 7 13 13 3 6 4 13 9 1 0 9 1 0 15 9 2
7 11 11 13 1 0 9 2
20 7 2 13 15 15 2 9 13 9 14 13 9 1 9 1 10 0 1 15 9
13 11 6 4 13 1 0 15 9 1 3 0 9 2
3 3 14 2
15 15 13 0 9 1 9 9 2 0 1 15 9 1 9 2
16 3 15 13 3 2 11 13 2 16 13 0 9 1 0 9 2
6 9 3 13 1 9 15
5 9 13 1 9 15
15 10 9 15 4 13 12 9 1 3 12 9 1 0 9 2
38 0 9 1 11 3 6 13 0 9 1 9 11 2 7 15 13 1 9 1 0 9 1 0 0 9 7 10 0 9 1 9 1 9 7 9 1 9 2
19 9 1 9 11 1 11 11 3 14 4 13 1 9 3 1 0 15 9 2
21 3 3 7 11 11 6 13 11 14 15 13 1 0 9 7 15 13 3 1 15 2
14 10 9 13 3 1 12 9 1 0 9 9 1 11 2
1 9
11 9 4 13 1 9 2 0 3 1 9 2
20 1 9 4 13 9 1 9 2 7 12 9 4 4 13 1 9 1 0 9 2
8 6 13 3 15 4 13 9 2
15 9 13 0 9 7 13 1 9 12 1 11 2 13 15 9
2 11 2
24 11 6 13 14 13 9 1 0 9 1 11 2 13 9 11 11 1 9 2 0 1 9 11 2
19 11 13 10 0 9 2 13 9 1 0 9 1 9 15 1 0 0 9 2
29 11 6 13 0 9 7 13 9 2 0 1 0 9 2 3 1 0 9 7 9 12 1 9 1 9 1 11 1 11
6 9 1 11 13 1 9
20 0 11 11 13 0 0 9 2 7 1 15 9 15 15 13 2 13 1 9 2
15 6 13 3 3 15 13 3 11 11 7 9 15 11 11 2
5 11 13 9 1 9
24 9 1 9 13 1 0 0 9 9 11 1 9 2 16 15 13 9 1 0 0 9 1 9 2
14 7 12 0 9 1 0 9 13 9 2 0 1 9 2
23 0 9 1 11 2 0 1 0 9 11 11 2 13 3 1 9 1 0 9 1 0 9 2
35 9 12 1 9 1 9 2 0 1 9 9 1 9 1 9 2 13 2 9 1 10 9 9 1 9 9 7 0 9 1 0 9 11 2 2
18 9 1 11 2 15 13 0 0 9 1 11 2 14 13 0 9 9 2
14 15 15 13 2 16 0 9 7 9 14 13 1 9 2
20 9 1 9 13 1 9 1 0 9 2 7 0 9 15 13 1 9 1 9 2
12 1 0 9 11 13 7 0 9 2 11 2 2
10 9 15 13 1 9 1 11 13 11 2
23 9 13 1 9 1 0 1 0 9 9 1 0 9 2 0 9 2 2 13 1 0 9 2
15 12 0 9 2 1 15 12 9 7 12 9 2 13 0 2
12 2 0 9 2 1 11 13 1 12 9 9 2
14 0 9 4 13 1 0 9 1 0 0 9 1 11 2
9 0 12 9 13 9 7 9 15 2
20 9 2 0 1 12 9 0 9 2 13 9 7 13 9 1 0 9 7 9 2
10 3 13 4 9 2 15 15 13 3 2
12 3 13 4 9 15 2 15 4 13 1 9 2
16 13 4 3 1 12 9 2 0 9 1 15 13 9 1 9 2
20 12 13 1 0 9 2 13 1 9 1 0 9 11 11 2 3 4 13 9 2
8 13 1 9 1 0 2 11 2
22 15 13 0 9 1 9 0 9 2 3 11 13 9 1 9 1 0 9 2 13 11 2
2 11 2
25 9 1 0 9 1 11 7 9 1 9 13 0 9 1 9 1 9 1 11 7 0 9 11 11 2
26 9 15 13 1 11 2 1 9 1 11 13 0 9 11 11 2 9 1 9 11 11 7 9 11 11 2
14 11 1 10 9 13 9 14 15 13 9 1 0 9 2
15 11 3 13 11 14 13 11 1 9 1 9 2 13 11 2
8 9 13 9 1 12 9 1 11
23 12 1 9 4 13 14 13 1 0 9 1 0 9 7 13 9 1 9 1 12 0 9 2
13 0 9 1 9 13 0 11 11 2 0 1 9 2
16 9 15 13 2 16 15 13 1 0 2 3 4 13 0 9 2
6 9 13 14 13 9 2
27 11 13 3 2 16 13 9 1 9 1 9 1 0 9 1 11 1 9 1 9 1 0 1 11 1 9 2
6 11 13 0 9 1 9
8 11 11 2 9 2 11 11 2
12 9 1 11 1 0 9 13 0 9 1 9 2
30 14 15 13 9 1 0 9 1 9 9 14 13 10 9 1 0 9 2 0 1 0 9 7 9 1 9 1 0 9 2
19 7 11 2 7 0 9 9 13 1 0 0 9 1 9 2 0 1 9 2
6 0 9 14 13 0 2
20 9 12 2 15 13 9 1 9 1 0 9 2 13 12 9 9 1 0 9 2
12 0 9 13 1 9 1 9 1 9 1 11 2
8 3 3 15 13 2 14 13 2
7 10 1 15 14 13 9 2
13 9 2 13 2 1 12 9 13 9 14 13 0 2
10 15 13 1 9 15 0 9 1 9 2
6 13 1 9 9 9 2
11 3 13 1 9 15 0 9 1 0 9 2
10 9 13 1 9 7 9 15 13 3 2
8 7 0 9 3 7 3 13 2
19 15 3 14 13 7 14 13 9 2 1 7 3 2 1 7 1 0 9 2
5 11 1 9 13 2
7 10 9 1 9 15 13 2
8 9 13 1 9 1 0 9 2
12 11 2 11 7 15 14 13 1 9 1 9 2
8 9 13 9 1 0 15 9 2
6 12 13 2 12 13 2
7 15 15 13 3 1 10 2
15 6 13 14 13 0 1 9 2 15 15 13 1 9 15 2
13 15 13 2 16 15 13 14 13 0 9 1 9 2
14 15 13 14 13 7 14 13 9 1 9 1 10 9 2
11 11 13 14 13 0 9 1 9 1 11 2
12 13 9 14 13 2 16 6 13 9 0 9 2
11 3 1 9 1 0 9 13 14 13 9 2
11 13 4 6 14 13 2 7 14 13 15 2
14 13 4 3 9 2 7 6 13 10 14 13 1 15 2
13 1 14 15 13 2 9 7 9 15 3 3 13 2
12 15 13 3 3 0 2 1 16 4 3 13 2
13 16 13 1 9 1 9 0 9 2 15 13 0 2
11 15 15 13 2 1 14 13 9 1 9 2
8 15 15 13 2 15 14 13 2
15 9 0 9 2 15 13 1 9 2 3 15 13 7 13 2
12 1 9 13 7 9 2 10 1 15 15 13 2
11 6 13 1 9 9 14 6 13 1 15 2
13 3 13 10 14 15 13 1 15 1 9 7 9 2
17 1 15 1 15 7 9 15 13 9 14 14 13 9 3 1 9 2
12 15 3 4 13 0 9 2 14 13 0 9 2
18 15 13 0 9 1 0 9 2 16 14 13 1 15 0 9 1 9 2
10 3 15 13 1 10 9 14 13 9 2
16 9 13 2 15 14 13 9 1 9 1 10 9 7 0 9 2
11 13 3 1 15 2 7 15 1 9 13 2
7 0 9 3 7 3 13 2
16 11 13 1 12 9 14 13 10 0 9 1 0 10 0 9 2
17 13 15 3 1 10 2 16 15 6 13 14 13 1 9 1 15 2
16 15 13 14 13 2 14 13 7 14 13 9 1 0 15 9 2
10 11 13 9 7 13 1 9 1 9 2
13 7 14 13 9 1 15 2 1 9 1 0 9 2
9 7 3 16 13 1 15 10 13 2
10 3 1 0 13 9 1 0 1 9 2
9 14 0 9 1 0 9 15 13 2
9 14 14 13 3 1 9 0 9 2
9 1 0 9 1 11 13 0 9 2
7 9 15 13 1 0 9 2
5 15 6 13 10 2
16 7 10 2 15 13 3 2 3 13 0 15 1 0 9 9 2
13 10 7 14 13 1 11 2 15 13 14 13 3 2
11 13 14 15 13 7 14 15 13 1 9 2
8 3 13 1 9 15 0 9 2
13 10 0 9 3 3 2 3 2 3 7 3 13 2
15 13 15 14 15 13 1 9 7 3 14 15 13 1 0 2
15 7 9 3 3 13 1 0 9 2 1 0 9 2 0 2
7 15 15 13 3 1 10 2
15 1 9 9 11 13 1 9 10 0 9 2 0 1 9 2
19 13 9 1 11 2 13 15 2 13 9 2 13 9 1 9 2 13 9 2
15 0 9 13 2 0 15 9 13 2 7 15 1 9 13 2
16 6 2 9 13 0 2 15 13 15 2 14 3 14 13 3 2
17 1 0 9 13 14 15 13 3 13 7 10 9 2 15 4 13 2
11 13 15 3 2 16 0 9 14 13 0 2
15 15 15 13 1 9 2 15 1 12 9 4 13 1 11 2
10 14 2 14 13 3 10 15 13 9 2
6 2 13 15 15 2 2
6 13 14 9 1 11 2
9 13 15 10 2 15 14 15 13 2
8 13 1 9 2 16 4 13 2
7 15 13 10 2 15 13 2
6 13 9 1 9 15 2
8 13 14 9 1 9 11 3 2
8 13 0 9 1 9 1 9 2
4 15 10 13 2
3 10 13 2
5 13 9 1 9 2
7 9 13 9 1 9 15 2
7 15 15 13 10 1 0 2
7 15 15 13 10 1 0 2
7 15 4 13 2 14 13 2
6 15 13 2 13 10 2
6 13 10 2 15 13 2
9 9 14 15 13 0 3 15 13 2
7 1 9 13 14 13 9 2
8 15 13 10 9 1 10 9 2
15 1 11 7 11 3 14 13 10 7 9 13 9 1 15 2
12 10 13 9 15 1 0 9 1 9 1 11 2
24 1 10 9 15 14 13 0 9 1 9 1 0 9 2 15 3 3 3 13 1 10 0 9 2
12 13 15 9 15 1 9 1 9 7 13 9 2
11 1 9 1 9 13 9 1 9 1 9 2
14 11 13 1 9 2 1 14 15 13 1 9 1 9 2
8 1 9 15 13 9 1 9 2
31 13 0 9 1 0 9 14 15 13 1 11 2 3 16 9 14 13 3 2 16 13 14 13 2 3 13 7 1 12 9 2
17 11 1 10 9 6 4 13 14 13 9 1 9 1 11 7 11 2
17 9 13 2 16 9 2 11 15 13 1 9 1 11 2 13 9 2
28 11 6 13 1 10 9 15 13 10 9 1 10 0 9 2 7 0 15 9 7 0 9 15 15 13 3 0 2
19 11 1 9 13 14 15 13 2 16 9 7 9 6 15 13 7 1 15 2
26 15 15 13 14 15 13 2 14 13 0 9 1 9 15 2 7 15 15 15 13 7 13 14 15 13 2
28 9 15 9 11 2 13 3 1 9 1 11 2 13 15 2 1 0 9 2 1 9 1 9 2 13 7 13 2
18 12 1 3 0 9 13 14 14 13 9 1 9 1 0 9 7 9 2
19 0 0 9 2 15 15 13 1 0 15 9 2 15 13 3 0 1 9 2
13 15 13 1 0 9 0 7 0 1 9 3 9 2
22 2 1 15 13 3 14 13 1 9 2 3 13 3 9 2 1 14 13 14 13 9 2
49 3 2 1 9 1 12 7 0 0 9 2 11 13 9 1 10 0 9 1 10 9 7 3 1 15 13 9 1 0 9 2 15 1 3 9 14 13 9 1 0 0 0 9 1 9 7 0 9 2
14 13 15 3 14 13 9 1 0 0 9 1 0 9 2
16 3 1 10 9 15 13 1 0 15 9 10 12 7 0 9 2
18 9 1 0 9 2 15 3 14 13 0 9 1 11 2 13 3 9 2
13 1 0 9 1 0 9 3 13 0 15 1 9 2
20 7 0 13 9 2 9 14 13 2 16 13 9 14 13 9 1 0 1 9 2
14 0 9 1 11 13 1 9 11 7 15 15 13 3 2
14 4 14 15 13 3 3 1 9 2 0 1 0 9 2
23 1 0 9 3 1 0 9 3 13 3 12 9 2 15 9 3 13 1 9 9 1 9 2
15 0 13 14 13 9 15 2 16 13 10 9 9 1 9 2
35 13 15 2 13 2 9 7 16 13 10 9 15 13 1 9 1 9 1 9 2 9 14 15 13 2 7 10 14 13 2 16 15 13 9 2
11 1 1 9 1 9 13 3 3 1 9 2
14 0 9 1 9 1 12 9 3 13 0 9 1 9 2
37 7 3 1 12 9 1 9 1 15 0 1 9 1 0 9 9 13 1 9 9 1 9 7 3 13 1 9 1 0 9 2 3 1 9 1 9 2
39 0 9 1 9 1 9 14 13 14 4 13 1 9 1 0 9 7 13 3 0 9 1 9 1 9 2 9 1 0 9 2 9 1 0 9 7 0 9 2
21 13 14 14 15 13 2 16 0 9 14 13 9 1 9 7 9 1 9 1 9 2
9 10 1 10 9 14 13 0 9 2
30 7 3 4 13 3 14 15 13 1 10 0 9 2 15 3 13 1 9 1 9 1 9 2 9 1 9 1 0 9 2
10 13 4 3 9 1 10 7 0 9 2
34 10 0 9 13 1 0 9 9 15 2 1 14 13 1 9 1 10 9 2 15 15 13 1 9 15 14 15 13 1 9 1 0 9 2
14 0 2 0 9 1 12 9 15 13 1 9 1 9 2
21 15 3 13 1 15 9 7 15 13 1 0 9 1 9 1 9 9 3 0 9 2
25 9 13 1 15 1 9 2 1 9 2 7 15 1 0 9 13 2 16 3 15 13 14 4 13 2
19 15 13 3 2 16 1 9 9 13 1 9 2 7 7 9 15 13 0 2
32 16 15 13 1 9 1 9 1 0 9 2 13 14 3 14 15 13 1 10 0 9 1 0 9 7 9 1 9 14 13 0 2
34 15 13 2 16 1 10 9 0 9 7 3 10 2 15 13 1 9 1 9 2 13 3 3 1 10 9 2 0 1 9 1 10 9 2
27 0 9 3 13 0 9 2 15 14 13 1 10 9 2 14 13 0 9 2 9 7 3 0 7 0 9 2
18 10 9 1 0 0 9 3 13 9 7 13 1 9 1 9 10 9 2
15 3 13 14 13 0 9 1 15 2 15 3 3 13 3 2
29 2 15 2 13 15 2 14 13 9 1 9 1 0 9 2 1 0 9 7 1 10 9 2 15 13 1 0 9 2
14 9 15 13 3 1 0 15 9 7 13 9 1 9 2
22 1 9 10 0 9 2 9 7 9 13 14 15 13 1 0 9 1 9 1 0 9 2
11 9 1 9 4 13 1 9 1 0 9 2
44 0 1 9 13 2 16 13 3 9 1 10 9 2 1 0 9 2 1 9 1 9 7 0 7 0 9 1 9 1 0 9 1 0 9 7 1 9 1 0 9 1 0 9 2
28 15 13 2 16 11 13 14 15 13 1 9 1 11 2 15 4 13 14 13 0 9 1 9 2 0 1 9 2
34 9 1 0 9 1 0 9 13 2 16 0 9 1 9 13 0 0 9 1 0 9 7 13 1 9 9 2 0 1 0 9 1 9 2
40 1 10 9 9 2 15 3 13 3 1 9 2 13 1 14 10 9 0 1 15 9 2 0 9 1 9 7 3 15 13 14 13 0 9 2 3 15 13 3 2
33 0 9 1 9 13 1 0 0 9 7 1 10 0 1 0 11 9 0 9 13 0 1 9 1 0 1 0 2 15 13 1 9 2
31 13 15 14 13 2 9 9 2 16 15 3 13 10 9 2 3 16 15 13 3 12 9 2 3 12 9 1 0 0 11 2
41 0 3 7 0 3 9 13 14 13 0 9 1 11 1 10 9 1 0 9 1 11 2 15 13 9 11 1 9 1 0 9 1 10 9 7 9 1 0 15 9 2
20 7 13 2 1 15 14 13 14 15 13 2 16 7 1 9 6 15 13 3 2
16 3 4 13 3 0 1 11 7 10 13 9 15 1 0 9 2
9 11 15 13 7 13 9 1 9 2
7 0 9 3 3 15 13 2
10 2 3 9 13 1 10 9 1 11 2
7 2 10 13 9 1 11 2
8 13 9 1 9 9 11 11 2
9 10 9 3 3 13 1 0 9 2
15 3 3 13 9 1 0 0 11 7 6 3 0 0 11 2
16 1 9 1 11 10 14 13 15 2 1 9 2 1 10 9 2
19 14 6 13 2 16 0 14 13 7 1 11 2 1 15 13 0 0 9 2
7 10 13 9 1 10 9 2
17 3 13 14 15 13 9 2 1 14 13 3 2 13 0 9 9 2
17 9 3 4 13 1 9 1 9 2 15 14 13 1 9 1 9 2
25 9 1 10 9 13 3 1 0 9 3 1 9 1 9 1 11 2 3 9 13 1 0 9 0 2
15 9 15 13 9 1 10 9 2 7 9 13 1 10 9 2
30 0 9 1 11 2 15 13 9 1 10 9 13 2 16 15 13 3 1 0 9 1 10 9 14 13 9 1 0 9 2
15 6 13 15 13 2 9 13 15 2 7 13 1 9 9 2
21 3 13 9 1 0 9 2 15 3 14 4 13 1 9 1 9 9 1 0 9 2
20 15 1 9 15 13 3 9 2 15 13 0 15 9 2 16 13 0 0 9 2
45 0 9 13 2 16 1 9 1 0 15 3 1 0 9 9 1 9 1 10 9 3 13 3 2 16 15 6 13 14 13 0 9 2 15 6 13 14 13 0 0 9 2 15 13 2
45 14 15 15 13 2 16 6 13 1 9 14 15 13 1 9 1 10 9 2 3 16 15 14 13 0 9 1 10 9 7 14 13 3 9 1 0 9 1 9 1 9 7 0 9 2
35 9 6 13 0 1 14 12 9 2 7 13 3 3 14 15 13 1 0 1 9 9 2 7 6 14 13 1 9 9 2 15 13 10 9 2
18 14 15 3 13 0 9 1 9 15 1 0 9 2 15 13 11 3 2
7 15 6 13 10 14 13 2
7 10 13 9 1 0 9 2
7 10 13 9 15 1 0 2
8 10 13 9 1 9 1 15 2
8 15 3 3 15 13 1 9 2
8 10 13 0 0 9 1 9 2
6 15 13 9 1 9 2
6 13 9 1 15 15 2
9 2 10 14 13 1 0 0 9 2
9 2 13 14 0 9 1 9 15 2
11 3 2 15 13 1 2 3 13 10 9 2
9 10 13 0 9 1 9 1 9 2
9 10 13 10 9 1 9 1 9 2
10 2 10 13 9 1 9 1 0 9 2
9 10 13 9 1 9 1 0 9 2
9 10 13 9 1 10 9 1 9 2
9 13 3 3 9 1 9 1 9 2
10 10 13 0 9 1 9 1 0 9 2
11 9 15 13 14 6 13 3 3 1 9 2
11 15 13 9 1 15 7 3 13 9 15 2
12 2 10 13 9 1 10 9 1 9 1 9 2
11 10 13 9 1 9 1 0 9 1 9 2
11 14 13 9 1 0 9 1 9 7 9 2
12 2 10 13 9 1 0 9 1 9 1 9 2
11 10 13 10 9 1 0 0 9 1 9 2
13 3 15 13 2 3 13 14 15 13 10 13 9 2
8 13 2 16 13 9 1 9 2
4 2 13 15 2
12 10 13 9 15 1 9 1 0 1 0 9 2
13 3 13 9 2 15 13 14 9 13 9 1 9 2
5 10 13 1 15 2
13 16 15 13 7 13 10 13 9 2 13 15 9 2
13 15 13 2 7 9 15 10 9 15 15 13 0 2
4 3 9 13 2
14 13 14 0 9 3 1 0 9 13 2 16 13 0 2
15 9 1 9 3 13 2 16 13 0 7 14 15 13 0 2
5 10 15 13 9 2
14 15 13 1 0 9 14 15 6 4 13 1 0 9 2
14 13 1 9 1 0 0 9 1 9 1 9 7 9 2
14 1 0 0 9 13 14 15 13 1 9 9 7 9 2
12 0 9 1 9 3 13 2 16 13 0 9 2
15 2 10 14 13 9 1 9 1 9 1 9 1 0 9 2
14 13 10 3 1 9 1 9 7 0 9 1 0 9 2
15 10 13 9 2 3 9 4 13 0 9 1 0 15 9 2
17 2 13 14 0 9 1 0 9 2 10 9 1 9 13 1 9 2
15 15 13 0 0 9 14 1 0 9 2 15 15 15 13 2
8 11 1 9 13 9 1 9 2
16 2 13 14 1 0 0 0 9 0 9 14 15 13 1 9 2
17 2 13 14 0 9 14 13 9 1 10 3 14 15 13 1 9 2
17 7 16 13 1 0 9 0 15 9 2 13 15 1 9 1 9 2
6 10 13 9 1 15 2
16 6 13 3 1 10 9 9 14 13 14 13 9 1 0 9 2
30 11 4 13 1 9 1 0 9 14 15 13 1 9 0 9 2 15 13 0 9 2 7 1 0 9 15 13 1 15 2
40 3 1 12 9 1 0 9 0 15 9 15 13 1 12 9 1 9 7 3 13 9 14 13 9 1 11 7 11 2 15 1 0 9 3 13 1 9 1 9 2
33 0 9 13 0 2 13 4 1 12 1 0 9 1 9 2 15 13 14 13 3 0 2 0 2 14 13 9 2 9 7 0 9 2
19 15 13 0 9 1 10 2 15 3 7 1 9 14 13 9 1 0 9 2
47 9 1 9 1 9 1 9 7 9 1 0 9 14 13 9 1 11 1 10 9 13 3 1 9 9 1 9 7 9 1 9 1 0 9 7 9 1 9 7 9 1 9 1 9 7 9 2
23 3 1 15 0 9 1 0 15 9 13 14 13 9 0 9 2 15 13 1 9 1 11 2
25 15 15 13 9 1 10 9 2 15 2 13 15 2 14 13 10 0 2 0 9 1 9 1 11 2
23 15 4 13 1 9 1 9 3 9 2 7 3 1 0 9 9 15 13 1 9 1 15 2
20 1 0 9 15 13 14 13 3 2 16 9 13 3 3 0 2 0 7 0 2
8 7 15 15 13 10 13 15 2
25 15 13 2 16 13 0 9 7 10 0 9 2 1 15 6 15 13 1 9 1 0 9 1 9 2
13 11 15 13 2 16 4 13 9 1 10 10 9 2
27 3 9 15 13 1 0 15 9 10 0 9 7 13 3 10 9 2 15 1 9 1 9 13 1 9 15 2
16 11 13 3 14 13 1 9 1 0 9 2 16 13 0 9 2
23 13 15 11 9 3 2 13 2 7 13 10 9 2 3 15 13 2 16 9 3 3 13 2
15 13 14 13 2 16 13 3 0 9 1 0 9 1 11 2
27 1 12 9 13 7 4 13 0 9 1 0 9 2 13 4 9 1 15 2 13 0 9 1 9 1 9 2
14 11 15 13 14 13 2 7 15 13 9 1 9 15 2
13 1 10 9 13 0 1 9 9 1 9 1 9 2
22 3 10 9 13 14 13 9 1 9 7 9 1 0 9 2 15 14 15 13 7 13 2
14 3 13 2 13 9 7 13 1 9 1 10 0 9 2
32 2 9 2 16 9 13 1 9 2 3 13 1 9 1 0 9 1 9 2 15 13 14 13 0 9 2 15 14 13 0 9 2
7 10 13 9 15 1 9 2
11 0 9 4 13 11 1 9 1 0 9 2
11 6 13 14 13 2 16 4 13 1 9 2
16 1 11 13 9 1 9 7 3 9 3 13 1 9 1 9 2
9 9 13 10 2 15 13 1 15 2
15 3 13 14 9 1 9 1 0 0 9 7 10 13 15 2
20 7 16 13 9 1 9 2 13 2 13 9 7 9 13 9 15 3 1 9 2
21 7 9 13 7 13 2 13 2 13 7 13 7 13 1 15 0 9 1 0 9 2
21 16 15 13 1 9 1 9 2 15 13 9 15 2 0 0 9 13 9 1 9 2
21 0 0 9 2 1 15 4 13 1 9 0 9 2 15 13 1 9 15 1 9 2
20 10 13 10 9 1 9 1 9 1 0 9 1 10 0 7 3 0 0 9 2
22 13 15 3 3 14 6 13 1 9 1 9 2 15 6 13 14 15 13 10 0 9 2
10 13 10 9 9 1 9 1 0 9 2
4 10 13 15 2
9 3 4 13 3 3 1 3 10 2
7 10 13 9 1 0 9 2
12 13 1 10 0 9 2 16 13 1 0 9 2
15 9 1 0 9 15 13 1 3 0 9 1 9 1 9 2
27 10 13 9 1 9 1 9 2 15 3 13 2 1 9 2 15 13 14 13 7 9 2 15 13 14 13 2
25 0 9 1 0 9 2 15 13 1 9 14 13 9 1 0 9 2 3 13 14 13 7 0 9 2
27 13 15 11 0 9 2 13 15 1 9 15 2 3 13 0 0 9 2 7 13 14 13 7 14 15 13 2
21 13 0 9 2 13 15 2 13 2 13 15 2 13 1 9 9 2 16 15 13 2
25 0 9 1 9 13 9 7 15 14 13 1 9 1 0 9 2 13 1 9 9 1 9 11 11 2
16 13 14 3 14 13 10 14 13 9 1 0 9 1 0 9 2
16 0 9 14 13 1 0 9 9 1 9 1 9 1 0 9 2
16 1 0 9 9 1 0 9 13 1 9 7 9 10 0 9 2
18 2 9 13 9 14 15 13 0 9 1 9 7 9 2 0 1 9 2
18 10 13 9 1 9 1 9 14 6 15 13 9 1 12 9 1 9 2
20 6 13 14 2 16 1 9 1 0 9 13 14 13 10 3 3 0 0 9 2
21 0 9 15 13 2 16 13 14 4 13 0 9 1 9 2 10 9 6 4 13 2
23 14 10 0 9 2 1 15 6 13 9 2 3 15 13 9 1 9 2 0 1 0 9 2
29 14 7 1 9 1 10 0 11 9 1 0 3 13 3 0 7 0 1 9 1 3 0 15 1 0 9 0 9 2
24 1 1 3 4 13 9 1 10 0 9 2 15 13 10 2 16 15 13 9 7 9 1 9 2
20 9 15 3 1 0 9 13 1 9 1 9 7 3 3 13 1 9 1 0 2
11 9 2 2 13 1 9 0 7 0 9 2
11 10 0 9 14 13 14 1 10 1 15 2
14 10 13 9 1 0 9 1 9 7 9 1 0 9 2
25 15 3 4 13 10 9 3 14 13 2 16 15 4 13 10 9 2 3 15 13 9 1 0 9 2
19 10 9 13 0 9 7 15 13 14 13 1 9 1 9 10 0 0 9 2
11 9 4 13 0 15 9 1 0 0 9 2
18 0 9 4 13 3 0 9 7 0 9 1 9 3 4 13 1 9 2
24 0 0 9 3 13 14 13 3 0 15 9 2 1 9 1 15 3 15 13 0 2 0 9 2
24 0 15 13 9 1 0 9 2 10 0 9 7 9 3 7 3 13 14 13 1 0 0 9 2
11 1 10 9 13 14 15 13 0 15 9 2
37 7 13 15 2 7 13 15 2 16 15 13 0 9 2 16 9 9 3 4 13 1 9 1 9 2 3 15 13 9 7 3 15 13 14 13 9 2
27 4 13 14 15 13 3 10 2 15 4 13 1 15 2 14 15 13 0 9 1 9 1 9 1 0 9 2
10 7 15 13 10 13 0 9 1 11 2
28 1 14 13 14 13 0 9 1 15 2 3 3 13 9 14 15 13 3 2 3 3 13 14 13 10 1 15 2
16 4 13 9 1 11 2 7 1 10 9 3 6 13 9 15 2
13 14 10 0 9 15 13 1 10 9 1 0 9 2
36 3 13 9 15 12 7 0 0 9 7 1 15 1 9 1 0 0 9 1 10 9 15 15 13 14 6 13 9 2 3 9 14 15 13 0 2
9 9 3 13 1 3 1 12 9 2
31 13 15 9 14 13 3 7 3 9 1 9 2 9 2 9 2 0 9 2 9 2 9 2 9 7 0 15 0 0 9 2
16 3 13 1 0 9 9 2 13 3 3 14 13 0 0 9 2
26 9 1 0 12 0 9 13 2 16 1 0 9 9 13 3 3 7 3 1 9 1 0 9 7 9 2
8 0 9 13 9 1 0 9 2
18 1 9 16 13 0 2 9 14 13 10 7 9 14 13 1 10 9 2
14 15 1 9 14 15 13 1 0 9 2 15 14 13 2
30 13 0 11 2 3 13 3 14 15 13 3 1 9 2 1 15 9 13 1 0 9 2 3 4 15 13 1 0 9 2
16 13 9 1 0 1 9 9 7 15 13 12 9 1 0 9 2
34 1 9 15 15 13 2 16 0 9 3 15 13 1 9 1 9 2 13 1 10 9 2 13 15 9 7 13 14 13 0 9 1 9 2
32 9 1 0 0 9 7 9 1 0 9 7 9 1 0 9 2 15 13 9 1 9 1 0 7 0 9 2 3 13 0 9 2
15 13 14 15 13 1 9 0 9 14 15 13 1 9 9 2
23 7 0 9 13 3 3 2 16 9 15 13 14 15 13 1 9 7 14 15 13 1 9 2
47 9 13 0 9 1 0 9 2 13 0 0 9 2 13 14 13 0 7 0 9 2 14 13 0 9 1 0 9 1 0 9 2 14 13 9 2 0 7 0 9 2 3 6 13 0 9 2
14 0 9 15 13 3 2 16 9 13 0 9 1 9 2
21 3 14 13 9 2 15 3 3 1 9 15 14 6 4 4 13 14 13 10 9 2
26 1 10 9 10 9 0 9 14 13 9 7 14 13 9 1 9 1 9 1 9 1 9 1 0 9 2
22 13 14 9 2 15 1 9 1 0 9 15 13 1 9 15 14 13 1 9 1 9 2
20 3 16 15 6 13 14 13 9 2 1 15 13 9 1 9 1 10 0 9 2
19 1 14 13 9 13 10 9 7 0 9 1 9 9 1 9 1 0 9 2
21 7 3 10 9 6 13 1 9 15 14 10 9 2 16 15 6 13 9 1 9 2
23 4 13 14 13 10 9 2 7 9 15 13 2 15 3 3 13 10 3 0 9 1 15 2
13 7 3 15 13 14 13 3 7 3 1 0 9 2
16 15 13 3 0 7 13 14 13 3 14 6 13 9 1 15 2
17 9 13 0 9 2 13 3 7 1 14 13 2 13 1 9 9 2
11 3 13 3 3 9 1 9 7 3 13 2
14 13 2 13 2 7 13 1 9 14 13 3 0 9 2
27 15 6 15 4 13 10 14 13 2 3 7 9 6 4 13 14 13 3 0 0 9 2 13 9 1 9 2
12 15 3 1 9 13 14 13 10 0 0 9 2
27 9 1 0 9 2 1 9 1 9 7 1 0 9 1 10 1 12 9 1 9 2 13 3 9 1 9 2
19 13 3 3 1 0 9 7 0 9 1 9 2 15 13 1 9 1 9 2
20 1 9 9 13 9 11 2 7 3 14 13 9 2 7 6 14 13 14 13 2
8 15 13 10 1 9 1 9 2
22 9 9 2 3 3 15 13 1 9 1 9 1 0 9 2 10 13 9 1 10 9 2
23 7 15 2 9 9 2 15 13 2 13 1 9 15 1 0 9 9 1 9 1 10 9 2
31 0 9 2 15 15 13 1 0 9 2 13 6 13 0 9 1 0 9 1 9 2 15 13 9 1 0 9 2 13 9 2
9 15 13 6 13 9 3 6 13 2
28 1 9 7 9 13 6 15 13 9 7 6 15 13 9 2 16 15 13 1 0 0 9 2 3 0 0 9 2
23 9 1 9 1 9 2 9 2 0 9 7 0 0 9 13 9 2 15 1 9 15 13 2
24 15 13 0 9 1 0 9 1 9 1 0 9 7 13 9 2 9 7 9 1 9 1 9 2
26 9 13 7 10 9 2 16 13 14 13 3 3 7 3 3 0 9 2 1 14 13 0 9 1 15 2
22 15 15 13 9 1 15 7 3 3 1 10 9 4 13 7 9 2 15 4 13 3 2
12 7 15 4 13 2 16 1 10 9 13 9 2
19 13 14 13 2 16 1 0 9 0 1 11 1 0 12 9 13 0 9 2
26 13 1 9 14 13 2 16 11 3 13 1 10 12 9 10 0 9 2 15 13 14 13 9 1 9 2
14 15 13 14 13 2 16 15 14 13 10 9 1 11 2
31 15 13 1 9 14 13 3 10 9 3 3 15 13 3 7 13 14 15 15 13 3 2 14 15 13 7 14 15 13 3 2
19 3 11 3 4 13 2 16 16 9 13 1 0 2 9 13 9 1 0 2
13 3 3 13 14 15 13 9 2 16 9 13 9 2
26 15 13 10 9 3 0 9 1 9 15 13 3 3 7 3 2 13 7 15 13 2 3 15 13 9 2
11 1 9 1 9 9 13 0 9 1 9 2
25 1 9 9 1 9 13 0 9 1 9 2 13 0 9 7 9 2 13 0 9 2 13 0 9 2
18 15 13 10 0 2 16 13 2 0 9 1 15 2 15 6 13 9 2
11 9 9 13 1 9 1 0 9 1 9 2
11 6 15 13 14 13 2 13 1 9 9 2
8 0 9 13 3 1 15 9 2
12 7 10 9 13 9 1 10 2 15 15 13 2
20 15 13 14 13 7 3 2 3 3 2 16 14 3 13 1 9 2 3 13 2
12 3 15 13 12 2 15 13 14 13 1 12 2
29 6 13 14 15 15 13 2 10 0 9 4 13 6 3 0 15 9 2 4 15 13 1 3 0 2 0 3 9 2
5 2 13 15 11 2
18 13 1 9 7 13 1 15 0 15 0 9 1 3 3 9 7 9 2
4 2 13 3 2
4 2 13 11 2
11 13 3 3 0 2 13 9 2 3 13 2
6 11 13 9 1 15 2
8 13 1 9 15 9 7 9 2
4 10 13 15 2
7 14 9 15 6 15 13 2
6 2 15 13 1 15 2
30 3 0 6 15 4 13 9 2 4 15 13 1 9 15 2 4 13 14 13 9 1 9 7 1 9 2 7 1 9 2
21 15 13 1 9 2 14 3 2 7 9 15 1 10 14 9 15 13 7 11 13 2
9 10 9 1 9 15 13 1 9 2
33 9 15 6 15 4 13 15 2 7 0 9 1 0 9 2 0 9 2 0 15 0 9 3 15 13 7 15 15 13 3 1 9 2
11 2 1 9 11 14 13 10 2 15 13 2
12 14 12 1 15 6 4 13 1 10 0 9 2
8 7 15 13 14 15 13 9 2
9 6 15 13 3 1 10 1 15 2
22 9 13 2 13 1 9 0 9 2 0 9 3 3 7 3 15 13 1 0 0 9 2
20 1 0 15 9 15 13 0 9 7 13 0 9 1 0 2 0 1 9 9 2
6 2 15 13 10 3 2
15 2 15 13 9 2 15 13 10 2 1 15 14 15 13 2
9 2 13 15 11 7 15 13 9 2
10 13 14 13 3 13 3 3 10 9 2
4 11 15 13 2
24 7 9 13 2 15 13 1 9 15 2 14 14 13 3 7 14 13 1 10 0 9 7 9 2
33 9 2 9 7 10 9 2 15 1 10 9 13 9 14 13 9 1 0 9 2 13 14 13 15 3 7 1 0 9 1 0 9 2
26 9 1 0 9 15 13 1 9 12 1 12 1 0 9 1 9 1 9 2 0 1 9 1 0 9 2
9 0 9 1 9 11 13 0 9 2
37 1 9 13 14 15 13 0 9 1 0 9 2 0 0 7 0 9 2 9 1 0 9 2 9 1 0 9 2 9 2 0 7 3 3 0 9 2
32 0 9 13 10 2 1 15 3 10 9 13 0 9 2 7 15 4 13 1 9 1 9 11 2 16 6 13 0 9 1 9 2
22 9 11 13 9 1 9 2 0 1 10 9 7 9 1 9 1 3 0 9 7 9 2
14 15 13 9 14 15 13 3 1 9 2 15 15 13 2
25 0 9 6 13 14 13 0 0 9 7 14 13 9 2 15 1 9 13 0 1 9 1 0 9 2
18 0 9 13 14 13 7 13 10 9 2 3 13 3 1 9 0 9 2
30 3 0 9 13 9 1 9 1 9 1 0 9 2 0 9 1 9 1 0 9 6 13 14 4 13 1 0 12 9 2
29 1 9 1 9 0 2 9 0 9 13 3 14 13 9 1 0 9 1 0 9 2 15 6 13 14 15 4 13 2
21 9 13 14 13 1 9 9 15 1 9 0 2 9 0 2 0 2 0 7 0 2
16 9 1 0 9 13 1 0 9 9 1 9 0 2 9 0 2
21 9 1 0 9 13 14 13 3 0 9 2 15 13 1 9 1 9 1 0 9 2
23 9 1 0 9 6 13 14 13 9 7 14 13 9 2 15 13 0 1 9 1 0 9 2
23 0 9 13 14 13 7 0 9 7 9 2 15 9 1 0 9 6 13 14 13 7 13 2
16 1 12 9 15 3 1 9 15 1 0 9 13 10 0 9 2
20 1 0 9 1 0 9 11 13 9 1 0 11 3 14 13 9 1 0 9 2
29 0 7 0 9 3 3 15 13 1 9 1 0 9 2 1 14 13 0 0 9 14 13 14 13 1 0 0 9 2
17 15 3 3 1 0 9 14 13 14 13 9 1 9 1 0 9 2
20 3 11 7 0 9 1 0 11 15 13 2 15 13 14 13 9 14 13 9 2
16 11 3 13 1 9 7 9 9 1 9 1 0 7 0 9 2
20 11 2 11 2 11 2 11 7 11 14 13 1 1 12 2 11 14 13 12 2
16 10 1 0 9 14 13 1 12 9 2 16 10 9 13 12 2
21 9 1 0 9 13 14 13 9 1 9 1 0 9 7 14 4 13 1 0 9 2
18 13 7 0 9 2 15 13 14 13 9 1 0 9 7 0 0 9 2
10 9 13 14 13 0 2 14 13 0 2
13 13 14 13 9 9 2 14 13 10 0 0 9 2
11 7 1 9 13 14 13 1 9 15 9 2
16 3 1 15 13 3 4 15 13 1 0 0 9 1 0 9 2
18 3 4 15 13 14 13 10 0 2 0 1 9 3 9 1 9 15 2
36 3 7 3 2 16 13 9 1 9 2 13 9 1 0 9 1 9 2 13 1 9 7 13 9 1 9 2 14 15 13 0 1 9 7 9 2
14 2 13 0 9 1 10 2 16 15 13 9 1 9 2
23 13 15 2 16 13 3 1 9 2 3 15 13 2 16 13 14 13 1 9 2 15 13 2
13 13 15 3 2 13 1 12 7 13 14 13 12 2
12 0 9 13 14 13 9 15 7 14 13 9 2
22 0 9 13 14 13 9 1 9 15 2 14 15 13 2 14 13 9 2 14 13 9 2
19 13 3 2 3 9 13 10 14 13 9 7 3 14 13 3 10 14 13 2
8 13 7 13 10 2 15 13 2
17 6 13 3 0 9 2 15 4 13 12 9 1 14 13 1 9 2
20 13 1 0 9 2 13 15 14 13 2 0 2 7 2 3 2 1 9 2 2
17 9 1 9 13 2 16 15 3 13 15 14 2 13 0 9 2 2
15 14 13 3 0 13 0 2 7 13 7 14 13 3 0 2
33 13 14 15 13 0 2 13 15 1 9 1 9 2 1 15 15 13 12 9 2 7 1 15 3 13 2 16 13 0 9 1 9 2
18 15 13 14 15 13 14 15 13 9 1 9 7 14 15 13 1 15 2
24 3 13 1 9 1 0 12 9 1 9 1 9 2 10 2 15 13 2 13 0 9 1 9 2
11 1 15 13 9 15 1 0 9 7 13 2
22 13 14 13 9 15 1 9 3 7 14 15 13 9 1 9 2 1 14 6 15 13 2
10 15 7 15 3 1 9 14 13 9 2
12 6 15 13 7 1 9 2 16 13 0 9 2
8 3 1 15 15 13 1 9 2
31 3 15 13 3 0 9 7 9 1 10 2 15 6 13 14 15 13 2 13 14 13 3 9 2 0 1 9 9 1 9 2
29 10 0 9 2 3 13 14 4 13 2 13 14 13 2 16 16 9 6 13 0 2 14 15 13 0 3 1 9 2
37 9 2 15 13 0 9 2 14 13 12 0 9 2 6 13 14 13 9 9 14 13 3 9 1 10 2 15 2 1 10 9 2 13 14 13 0 2
14 2 0 9 13 12 9 2 15 13 9 7 0 9 2
20 1 15 15 13 14 13 3 15 13 3 9 1 10 9 2 1 15 13 10 2
25 6 13 14 2 16 15 13 9 1 9 3 3 6 4 13 1 10 15 13 9 1 9 1 9 2
16 7 15 14 13 3 2 14 1 9 2 9 1 0 15 9 2
10 9 13 10 2 15 15 13 1 9 2
27 3 9 15 13 14 13 9 7 14 13 9 2 15 15 13 1 9 14 4 13 7 13 9 1 10 9 2
22 13 14 13 3 0 9 0 9 2 15 4 13 7 15 13 3 7 3 1 0 9 2
42 10 0 9 6 4 15 13 2 16 9 13 9 1 9 2 1 9 1 0 15 9 2 1 0 9 3 1 9 7 9 1 0 9 2 13 15 0 2 0 7 0 2
35 9 15 1 10 9 2 1 0 0 9 2 0 9 2 15 15 13 0 7 0 9 1 9 2 15 13 3 3 1 9 1 10 1 15 2
14 13 14 13 2 16 15 13 11 7 13 0 1 9 2
20 7 15 6 13 14 13 9 7 0 11 13 1 9 15 14 13 1 15 9 2
20 16 13 3 9 2 9 13 14 13 0 2 15 13 10 2 15 13 14 13 2
18 15 13 2 16 0 9 13 0 2 16 1 9 15 6 4 13 10 2
31 7 1 10 9 15 13 14 13 9 1 10 1 10 9 9 2 15 4 13 1 9 1 9 1 10 9 2 15 13 0 2
14 11 6 4 13 10 2 15 15 4 13 1 10 9 2
25 15 13 2 16 0 9 1 10 9 2 2 9 1 11 2 15 4 13 2 2 6 13 10 9 2
23 16 13 3 14 13 2 0 9 2 2 9 3 13 14 15 13 1 11 2 14 10 9 2
14 15 1 10 9 1 9 15 4 13 1 9 7 9 2
19 9 4 13 0 9 1 9 1 10 2 3 9 15 13 1 9 1 9 2
13 15 4 13 9 15 1 9 1 9 1 0 9 2
14 13 14 14 15 13 7 14 15 13 0 9 1 9 2
17 3 13 14 15 13 14 15 13 3 1 9 2 1 15 15 13 2
31 9 15 1 9 1 10 9 13 14 13 1 9 1 10 9 9 2 15 6 4 13 1 0 9 2 0 15 1 0 9 2
10 9 3 13 0 2 7 9 13 9 2
17 13 10 9 1 9 1 9 1 9 7 1 0 15 1 9 9 2
8 14 10 9 1 9 1 9 2
28 9 0 13 0 9 1 10 2 3 14 13 9 1 10 9 1 9 2 7 3 14 13 14 15 13 1 15 2
21 13 14 13 9 2 15 13 9 2 0 15 3 2 1 9 1 0 9 1 9 2
18 0 9 13 14 15 13 14 13 0 15 2 15 4 13 1 0 9 2
14 3 9 13 1 9 7 9 15 1 9 1 10 9 2
6 10 13 14 15 13 2
7 0 2 11 2 15 13 2
23 16 0 15 9 13 2 16 13 9 1 9 2 14 13 14 13 0 9 2 15 13 0 2
32 10 9 13 0 1 9 1 9 2 3 15 13 14 13 0 9 7 9 1 9 7 14 13 10 1 15 13 3 1 0 9 2
28 3 9 15 13 1 0 1 9 9 2 3 13 2 16 13 10 2 15 13 14 13 1 9 7 1 0 9 2
12 2 13 15 15 9 14 13 7 14 13 2 2
22 15 13 14 15 13 1 9 1 9 2 1 15 9 15 13 14 15 13 1 9 15 2
20 2 13 4 2 3 15 13 14 13 0 1 9 2 3 3 6 13 10 2 2
15 3 16 0 13 3 3 1 0 9 2 13 0 9 9 2
23 9 1 9 13 3 14 13 3 13 0 1 9 7 9 1 9 15 2 13 0 9 2 2
9 14 10 9 2 11 2 0 2 2
16 2 13 9 2 1 15 13 14 15 13 14 13 0 9 2 2
14 2 13 14 13 1 9 2 15 13 0 7 0 2 2
16 2 13 9 2 1 15 13 14 15 13 1 9 1 0 2 2
14 2 13 9 2 1 15 9 15 14 15 13 3 2 2
14 2 13 9 2 1 15 13 14 13 1 0 9 2 2
8 2 13 14 15 13 9 2 2
10 2 13 14 15 13 1 0 9 2 2
15 9 13 14 6 13 9 14 15 13 2 3 15 13 0 2
27 3 3 15 13 14 13 0 9 7 14 13 1 0 9 2 9 3 15 13 2 16 6 13 10 0 9 2
21 9 1 9 1 9 7 9 3 15 13 0 7 15 13 1 9 1 2 0 2 2
29 9 2 15 15 13 3 2 13 10 2 2 0 2 1 9 1 9 1 9 7 0 1 9 1 9 15 1 9 2
31 0 0 15 13 0 9 1 9 1 0 9 7 15 13 14 15 13 9 1 9 1 15 1 9 2 9 7 9 1 9 2
29 13 1 9 2 3 9 13 0 9 1 9 15 2 9 2 0 9 7 0 9 2 15 6 13 3 9 7 9 2
11 1 3 3 14 13 14 15 13 0 9 2
16 1 1 12 9 4 13 14 13 3 3 2 1 14 15 13 2
14 6 15 13 1 0 9 12 14 13 9 2 13 9 2
6 13 0 11 1 9 15
18 9 13 1 9 1 9 1 0 9 1 11 2 11 2 1 9 11 2
10 15 13 11 11 1 11 1 11 3 2
18 2 1 9 1 0 9 3 13 9 2 2 13 1 9 15 9 11 11
9 12 9 15 13 1 9 1 9 2
15 13 1 9 12 9 2 13 1 9 1 0 15 7 13 2
27 9 3 13 0 9 2 6 9 7 9 2 7 9 1 9 2 9 14 13 1 9 7 9 1 0 9 2
4 13 9 1 9
6 13 12 9 9 1 9
20 3 15 13 9 1 0 0 9 2 0 9 13 1 9 2 16 9 13 9 2
33 3 0 12 9 0 9 14 13 3 7 1 9 1 0 7 0 9 14 13 9 1 0 9 1 9 2 15 14 15 13 1 11 2
23 1 0 0 0 9 3 13 0 9 7 3 3 13 0 9 1 9 2 13 9 0 2 2
18 3 14 13 2 16 13 1 9 12 9 2 15 13 3 1 12 9 2
6 2 13 2 11 2 2
20 9 1 11 3 4 13 9 1 9 1 11 2 15 3 4 13 1 10 9 2
6 13 11 1 12 1 12
11 9 11 11 13 1 9 10 0 12 9 2
10 2 13 0 3 9 1 0 9 11 2
40 14 13 2 11 2 1 9 1 0 9 2 16 6 4 13 9 7 9 2 0 1 9 1 9 1 2 11 2 2 11 2 2 13 3 9 1 9 11 11 2
25 9 1 9 1 9 4 13 0 9 1 0 9 2 11 2 1 9 9 1 9 1 9 1 11 2
11 2 13 9 1 11 1 9 11 11 2 2
16 9 1 9 1 11 2 11 2 13 0 9 1 0 15 9 2
22 3 9 15 13 1 9 2 1 3 0 9 13 9 1 9 2 3 0 9 13 2 2
24 9 13 1 0 9 14 13 1 0 9 1 11 2 11 2 1 14 6 13 9 1 0 9 2
29 9 13 2 16 12 9 1 0 9 13 9 2 15 3 13 9 2 7 1 0 9 9 1 0 9 13 12 9 2
5 2 13 9 2 2
4 2 13 11 2
17 3 11 15 13 1 12 9 1 0 9 1 11 7 3 13 0 2
18 9 1 10 9 1 0 9 13 14 13 9 1 15 1 0 0 9 2
9 0 9 13 1 9 0 9 3 2
18 16 9 1 0 9 13 0 9 1 0 15 9 2 3 13 0 9 2
20 13 15 1 12 9 14 13 2 1 14 15 13 2 7 1 15 13 0 9 2
14 11 13 2 11 2 2 11 2 1 9 1 2 11 2
27 11 1 2 11 2 13 0 9 1 9 1 9 1 9 1 11 2 11 11 2 2 13 3 1 0 9 2
4 2 13 15 2
10 2 13 4 0 9 1 11 11 11 2
24 1 0 9 13 0 9 1 2 11 2 11 11 2 15 13 1 9 1 9 0 2 11 2 2
26 9 3 14 15 13 2 16 10 0 9 15 13 1 0 0 9 2 1 14 13 0 1 15 0 9 2
6 2 13 9 1 9 2
7 2 13 9 1 0 9 2
27 0 9 2 11 2 3 14 13 6 12 2 7 12 9 1 9 1 9 1 0 9 1 9 1 0 9 2
30 9 1 9 2 11 2 3 14 15 13 1 0 9 2 0 1 9 7 12 9 2 16 7 12 14 15 13 1 9 2
16 0 9 13 9 1 9 1 11 14 13 1 0 9 0 9 2
28 9 14 13 3 9 1 9 1 9 1 9 1 0 9 1 0 9 2 11 2 11 11 1 9 1 9 11 2
24 9 13 0 0 9 1 9 1 12 1 12 1 0 9 1 9 1 9 1 12 9 0 9 2
25 11 2 0 3 9 1 9 1 9 1 11 2 13 0 9 1 9 1 0 9 2 12 1 12 2
26 9 3 13 12 9 9 1 2 11 2 1 9 1 0 9 2 1 14 15 13 9 1 9 0 9 2
21 9 13 1 3 9 14 15 13 7 9 2 15 0 9 13 14 13 1 0 9 2
5 0 13 9 1 9
16 9 13 14 13 9 1 0 2 13 3 9 1 0 1 11 2
20 1 15 14 15 13 3 14 13 1 9 1 9 7 3 14 13 1 0 9 2
19 1 9 1 9 9 13 1 0 9 9 7 0 9 1 9 1 0 9 2
14 1 9 2 3 9 2 13 14 15 13 12 9 9 2
22 11 1 9 13 9 12 1 11 1 9 1 9 2 9 1 0 9 1 9 7 11 2
8 14 12 6 4 13 1 15 2
41 15 3 3 13 9 2 3 1 12 9 2 16 13 0 9 2 0 15 9 13 9 1 9 15 7 15 13 1 0 9 2 1 14 13 2 16 4 13 1 9 2
28 15 13 0 9 2 13 14 13 0 9 2 15 14 13 9 15 2 16 15 13 14 14 15 13 1 10 9 2
28 15 13 0 9 2 13 14 13 0 9 2 15 14 13 9 15 2 16 15 13 14 14 15 13 1 10 9 2
16 0 7 9 3 6 15 13 1 9 3 3 14 15 13 9 2
35 11 11 6 13 14 13 2 16 4 13 3 9 1 9 2 1 14 13 3 9 1 0 9 7 14 14 13 3 1 0 15 9 0 9 2
24 1 9 0 1 9 14 13 12 9 1 11 2 16 1 9 1 0 9 9 13 12 1 12 2
25 9 13 9 14 13 3 3 9 1 9 7 9 2 15 14 15 13 1 9 1 9 7 1 9 2
48 7 1 11 13 2 16 1 0 0 9 9 14 13 1 9 0 9 2 1 12 9 9 2 1 14 13 0 15 9 2 9 7 0 9 1 9 7 9 2 9 7 9 1 9 2 0 9 2
22 16 13 10 9 2 13 14 13 2 16 0 9 14 15 13 3 1 9 1 0 9 2
16 3 9 7 0 9 13 14 13 3 7 14 13 1 0 9 2
21 10 9 13 2 16 13 3 14 15 13 3 0 9 2 15 14 13 1 0 9 2
43 2 0 15 9 13 12 2 6 13 10 9 1 9 2 0 1 9 1 0 9 1 9 1 9 2 14 13 0 7 0 2 3 12 9 1 11 3 15 13 1 0 9 2
21 10 9 13 2 16 13 3 14 15 13 3 0 9 2 15 14 13 1 0 9 2
8 2 10 13 9 1 10 9 2
24 2 6 4 13 3 13 1 0 0 9 2 13 3 2 16 3 0 9 1 0 9 13 0 2
28 16 9 6 13 0 1 0 9 2 14 14 13 9 7 9 14 15 13 9 1 10 9 2 1 15 14 13 2
18 6 13 3 14 15 13 0 9 1 9 2 16 13 9 1 12 9 2
33 1 0 9 13 9 2 15 14 6 13 9 14 15 13 1 0 9 7 14 6 15 13 10 14 13 2 3 9 15 13 1 9 2
18 3 13 14 15 13 14 13 2 16 0 0 9 14 13 3 10 9 2
15 6 13 3 14 13 3 12 2 1 0 9 14 13 11 2
8 3 9 15 3 7 3 13 2
22 0 9 2 0 9 7 0 9 4 13 3 1 9 9 1 2 0 9 2 12 2 2
39 1 0 9 0 0 9 1 11 11 11 13 14 4 4 13 1 9 1 9 1 2 11 2 1 0 9 14 13 1 9 1 0 9 11 1 0 15 9 2
22 0 9 13 0 9 1 0 9 7 9 11 11 6 13 14 13 9 2 0 1 9 2
15 9 13 1 9 1 11 7 13 1 9 11 1 0 9 2
30 9 1 0 9 2 11 2 11 11 13 9 1 0 1 0 2 16 9 15 13 9 7 13 2 14 13 7 9 15 2
7 2 10 1 2 11 2 2
9 2 0 1 11 2 13 3 1 11
12 9 1 9 3 15 13 1 9 1 0 9 2
21 3 3 13 9 7 1 0 9 1 9 2 0 9 2 15 14 13 1 12 9 2
6 11 14 13 9 1 11
33 0 9 1 11 11 11 4 13 0 0 9 11 11 1 9 1 11 14 13 9 2 15 13 9 1 9 1 11 2 13 0 9 2
22 0 9 3 13 1 9 1 11 2 16 9 1 9 14 13 1 0 9 1 0 9 2
10 9 1 11 13 2 16 6 13 0 2
4 2 13 11 2
25 1 0 9 0 0 9 14 13 1 9 1 11 7 11 2 16 0 13 9 9 14 13 15 9 2
15 0 9 14 13 1 11 1 9 1 2 11 2 7 11 2
21 1 10 9 11 13 1 0 9 2 13 1 0 15 9 7 13 1 9 0 9 2
22 9 9 1 0 9 13 0 9 1 11 11 1 11 2 15 4 13 3 1 9 15 2
31 12 9 9 1 9 3 14 15 13 1 9 1 9 1 10 2 15 13 9 1 9 15 2 13 1 2 0 9 2 3 2
22 1 12 9 13 14 13 0 12 9 1 9 2 13 9 1 2 0 9 2 11 11 2
16 15 13 3 1 9 1 9 1 9 9 1 0 9 11 11 2
12 12 13 9 1 0 9 1 9 0 9 3 2
13 12 13 9 1 11 2 13 3 9 1 0 9 2
6 11 13 0 11 1 11
22 9 11 11 13 1 11 9 1 12 9 1 9 1 9 2 13 2 11 11 2 3 2
17 3 1 0 9 13 3 14 15 13 0 9 7 3 14 13 15 2
19 9 15 14 13 9 12 9 9 1 0 9 2 1 15 14 13 0 9 2
8 11 13 1 9 12 9 9 2
23 1 9 9 1 9 1 9 1 9 1 9 11 11 13 1 9 3 0 9 13 10 9 2
33 9 13 2 3 6 13 3 1 9 1 0 9 14 13 3 9 7 0 9 1 9 2 15 3 13 1 11 1 0 15 0 9 2
5 10 13 11 11 2
12 0 9 1 9 1 0 9 13 3 12 9 2
15 1 9 16 9 4 13 9 1 0 9 2 12 1 12 2
34 9 11 11 13 2 16 0 9 3 14 13 1 0 0 9 1 9 1 9 7 9 2 15 13 3 1 12 1 12 1 0 15 9 2
14 2 3 9 14 15 13 14 6 13 0 9 1 9 2
16 2 13 1 2 9 2 0 9 1 2 11 2 11 11 2 2
17 11 11 13 11 1 11 2 16 6 15 13 9 1 2 11 2 12
6 0 13 3 11 11 2
24 15 15 13 2 16 14 13 11 1 11 2 16 0 6 15 13 9 1 9 2 11 2 12 2
21 1 12 9 11 13 9 1 9 2 3 0 9 15 13 1 11 2 13 9 9 2
25 6 13 14 13 0 9 14 15 13 1 9 1 10 9 2 13 1 9 11 2 16 9 13 9 2
10 2 11 15 13 2 15 13 1 9 2
18 11 11 13 10 1 0 1 9 1 0 9 2 11 2 1 0 9 2
18 16 0 9 1 9 1 9 13 2 1 9 13 14 13 14 15 13 2
20 9 7 9 1 0 9 13 1 9 1 9 11 14 13 9 1 0 15 9 2
22 9 1 9 1 1 12 9 13 3 7 9 13 14 13 1 9 3 10 9 7 9 2
13 3 15 3 3 14 15 13 9 1 11 1 11 2
8 9 1 0 9 13 0 9 2
8 13 15 14 13 9 1 9 2
16 2 13 9 7 9 1 2 11 2 1 9 1 9 1 9 2
11 2 10 15 13 9 1 9 1 9 15 2
8 2 13 3 1 9 11 2 2
11 2 13 9 1 2 11 2 11 11 2 2
38 2 0 2 13 1 12 1 12 2 7 13 3 9 1 9 1 9 11 11 2 15 6 13 12 0 1 15 9 1 9 1 0 9 1 11 7 11 2
29 0 9 1 9 12 11 11 13 0 15 9 1 9 7 13 14 13 9 7 9 15 1 0 9 1 12 9 9 2
20 9 1 0 9 11 11 3 13 1 9 2 16 15 15 13 14 13 0 9 2
5 2 13 11 11 2
9 13 1 11 9 1 9 12 12 9
23 11 13 9 1 9 1 0 9 1 11 2 7 13 1 9 9 12 12 2 15 13 3 2
6 13 1 9 11 1 9
14 9 1 13 4 13 1 9 1 0 0 9 11 11 2
23 16 9 13 1 11 2 15 13 14 4 13 1 0 9 7 9 2 7 9 14 13 0 2
20 15 15 13 15 14 13 0 1 0 9 2 1 3 15 4 13 1 0 9 2
14 15 13 0 1 9 1 11 1 11 1 9 1 9 2
16 0 9 15 14 13 1 9 0 9 1 9 15 1 0 9 2
10 1 0 9 13 14 15 13 12 9 2
9 15 13 14 13 0 1 12 9 2
17 9 11 11 14 13 1 9 1 0 9 9 1 0 9 1 9 2
30 10 9 1 0 9 4 13 14 13 0 9 1 9 0 9 0 9 2 3 14 13 1 9 0 0 9 2 13 11 2
25 0 9 13 2 16 13 0 1 9 1 0 9 2 1 14 6 13 3 15 14 13 9 9 12 2
20 13 9 1 9 7 0 9 2 15 13 7 14 15 13 9 7 14 15 13 2
32 0 9 1 11 13 9 15 2 16 13 1 9 15 9 1 9 7 13 9 1 9 1 0 9 2 13 9 2 11 11 2 2
22 11 13 2 16 13 9 2 0 1 9 1 9 2 3 1 9 14 15 13 1 15 2
27 1 10 9 11 3 13 14 15 13 2 16 1 0 9 1 0 9 0 9 14 13 0 9 1 0 9 2
8 0 9 13 9 1 9 1 11
23 9 13 2 16 9 15 1 0 1 0 9 9 13 14 15 13 0 9 7 9 1 9 2
20 1 9 1 9 14 15 13 1 9 9 12 9 2 13 0 9 11 11 3 2
15 9 1 11 13 9 1 12 1 12 1 9 2 13 9 2
27 10 1 9 11 13 1 0 15 9 2 15 13 1 9 15 1 9 1 9 1 0 9 1 11 11 11 2
20 11 13 9 1 11 2 1 14 13 14 9 14 13 0 9 1 0 0 9 2
26 9 1 0 9 9 11 11 4 13 1 9 9 1 9 1 0 9 2 13 9 2 12 9 2 3 2
26 9 1 0 9 1 11 11 11 4 13 0 9 1 9 1 9 11 11 7 11 11 2 13 3 3 2
21 9 1 11 4 13 1 11 11 1 11 2 9 1 11 2 11 2 11 11 2 2
8 10 13 1 0 9 1 9 2
13 15 13 1 9 9 1 0 9 7 9 1 11 2
14 3 13 10 0 9 2 13 3 1 9 9 11 11 2
27 9 6 15 13 2 16 16 0 9 3 13 14 13 1 0 9 1 0 9 2 14 13 3 9 14 13 2
22 1 14 15 13 2 11 14 13 1 9 3 0 3 0 9 1 9 15 2 13 9 2
16 3 9 6 13 14 13 14 1 9 9 1 15 2 13 11 2
5 13 11 11 1 9
16 1 0 9 9 11 11 3 14 15 13 1 0 1 11 12 2
9 2 11 2 13 9 1 9 1 11
11 2 13 9 1 2 11 2 11 11 2 2
30 9 1 10 2 16 11 14 13 3 0 9 1 9 1 9 1 2 11 2 7 11 2 13 1 9 1 2 9 2 2
11 2 13 9 1 2 9 2 11 11 2 2
11 14 13 14 13 0 9 7 14 13 0 9
4 2 13 11 2
4 2 13 9 2
4 9 15 13 2
17 15 13 1 9 2 11 2 1 11 9 1 11 9 11 11 3 2
7 1 9 1 11 11 1 11
25 1 12 9 1 9 1 9 1 12 9 1 11 0 9 9 1 9 13 1 9 2 11 11 2 2
34 11 11 13 1 0 9 11 11 1 0 9 1 0 0 9 1 12 9 1 0 1 11 2 9 2 0 9 1 9 1 9 7 9 2
5 2 13 11 2 2
17 13 1 9 2 7 16 6 13 9 2 6 13 14 13 10 3 2
17 3 3 0 1 9 0 9 13 9 1 9 1 9 1 0 9 2
14 11 7 0 0 9 3 13 14 13 0 9 1 0 2
11 9 13 2 3 1 15 4 13 7 15 2
23 0 9 1 0 2 0 9 2 4 13 2 16 13 1 9 12 9 9 2 13 11 3 2
16 15 13 1 9 1 9 2 9 2 9 1 0 9 11 11 2
24 3 1 9 1 0 9 1 9 13 9 1 11 9 1 11 7 9 1 9 1 10 0 9 2
15 3 15 6 4 13 1 9 0 9 2 13 2 11 2 2
11 11 7 11 3 13 9 14 13 9 3 2
5 2 13 11 11 2
13 1 11 13 14 14 6 13 1 9 1 9 9 2
25 0 0 9 13 1 9 1 11 2 15 13 1 9 14 2 13 2 13 7 13 2 10 0 9 2
11 11 3 13 9 1 9 1 12 1 0 2
12 13 3 1 9 1 9 2 16 13 14 13 3
9 2 13 9 1 9 11 11 2 2
4 2 13 11 2
13 1 9 9 13 14 15 13 3 9 3 13 9 2
21 3 1 12 9 1 10 9 9 15 4 13 1 9 9 12 9 1 9 1 9 2
19 0 2 15 13 3 2 13 2 16 9 13 9 15 1 9 2 13 15 2
7 14 13 1 12 9 0 9
26 0 10 9 0 9 15 13 1 9 1 9 1 9 2 15 13 14 13 9 1 2 11 2 7 9 2
28 1 0 9 0 9 2 0 1 9 1 9 2 13 1 9 9 2 15 6 13 3 3 14 15 13 1 9 2
44 0 0 9 3 15 13 1 9 1 11 2 16 13 9 1 0 9 1 11 1 9 1 9 1 10 9 14 4 13 7 3 0 9 1 0 9 2 0 1 0 9 11 11 2
22 10 0 9 6 13 14 13 9 1 11 1 9 1 9 1 11 7 11 2 13 9 2
33 1 12 9 0 9 11 11 13 1 0 9 9 2 15 13 0 9 1 11 14 13 9 1 0 0 9 2 7 14 13 0 9 2
11 9 1 9 1 0 9 3 3 15 13 2
11 3 9 1 0 9 1 9 13 0 9 2
12 10 9 15 13 3 0 2 13 15 10 1 9
7 1 9 1 11 11 1 11
12 9 1 11 13 14 13 3 9 2 15 13 2
14 9 13 1 12 9 7 0 9 1 9 1 0 9 2
11 9 13 1 12 9 2 16 11 13 3 2
15 1 0 9 0 9 4 13 1 9 7 9 1 0 9 2
18 9 1 0 9 7 3 0 9 13 12 1 3 9 1 9 1 11 2
4 2 13 9 2
23 9 15 13 1 9 2 7 1 2 11 2 13 2 16 14 13 3 0 1 0 0 9 2
13 1 9 9 1 9 1 9 13 9 1 9 11 2
21 3 0 9 4 13 1 9 2 15 6 13 14 14 15 13 9 2 13 3 9 2
22 2 11 2 14 13 1 9 1 9 12 9 9 1 11 2 13 1 0 0 9 3 2
16 1 0 9 3 15 13 14 13 9 1 11 2 9 11 11 2
4 2 13 11 2
4 2 13 11 2
16 15 13 14 13 0 9 7 14 15 13 1 9 9 1 11 2
15 3 13 3 14 13 1 9 2 14 13 7 14 13 9 2
15 13 2 16 1 2 14 15 13 6 13 14 15 13 9 2
14 13 3 14 13 14 15 13 9 7 14 13 1 9 2
11 2 14 15 13 3 14 13 10 13 3 2
8 2 9 6 13 10 1 9 2
11 13 14 13 14 13 15 7 14 15 13 2
22 3 13 14 15 13 7 14 13 1 9 15 2 7 6 14 13 3 14 13 1 15 2
18 2 6 2 1 16 3 13 9 1 0 9 1 9 1 9 7 9 2
37 9 15 13 1 9 1 9 1 0 9 1 1 12 9 1 11 2 15 3 1 12 9 9 13 9 1 9 1 9 1 0 1 9 9 1 9 2
32 0 1 0 9 9 12 1 11 2 11 11 4 13 1 12 9 1 9 1 0 9 2 12 1 0 9 1 0 9 1 11 2
19 6 13 9 1 9 2 0 2 1 9 1 10 9 1 0 9 11 11 2
5 2 13 11 11 2
4 2 13 11 2
29 1 9 1 2 11 2 1 12 1 12 1 9 1 11 11 13 2 16 1 0 0 9 1 9 14 13 9 15 2
14 3 14 15 13 14 13 9 7 14 13 1 0 9 2
31 16 13 3 2 16 15 3 13 14 13 0 2 14 15 13 1 0 9 3 2 3 13 9 7 13 1 9 7 9 15 2
30 11 14 13 1 0 9 9 1 9 1 9 2 15 14 15 13 3 1 9 2 13 3 1 9 1 9 1 9 3 2
8 13 1 12 9 9 1 0 11
6 9 6 13 11 1 9
16 9 6 13 9 11 1 9 2 9 0 2 1 11 3 3 2
18 0 0 9 13 14 13 12 9 1 0 9 1 9 1 3 0 9 2
26 0 9 13 1 9 11 11 2 15 4 13 1 9 1 0 9 11 11 7 9 15 2 13 3 3 2
15 4 14 13 14 13 9 1 9 12 9 7 14 13 3 0
9 0 11 4 13 1 9 1 11 2
19 1 9 13 0 3 9 11 11 2 15 15 13 2 7 12 0 0 9 2
26 1 3 0 9 1 11 9 11 11 13 3 3 14 13 9 1 11 14 15 13 1 11 2 13 9 2
19 9 1 0 9 11 13 1 9 0 15 9 1 0 9 2 13 0 9 2
7 2 13 9 1 0 9 2
39 0 9 3 13 1 0 9 2 7 0 9 1 11 1 0 9 14 13 9 1 9 1 2 11 9 2 3 3 13 9 15 14 13 10 9 1 0 9 2
25 9 2 15 1 9 1 11 13 14 13 7 13 1 11 2 13 0 1 9 15 7 13 12 9 2
17 2 11 2 13 9 1 11 0 9 2 16 13 1 12 1 12 2
30 0 2 0 2 0 2 0 7 3 0 2 9 14 13 9 15 1 9 2 9 2 9 7 14 13 9 1 9 15 2
33 3 15 14 13 2 16 15 13 0 2 13 15 1 9 2 9 7 9 2 1 14 13 9 1 9 15 1 9 2 9 7 9 2
19 11 11 4 13 1 9 1 9 7 13 2 0 9 2 1 9 1 9 2
9 2 13 3 14 13 9 1 9 2
23 0 9 13 1 9 2 16 9 14 13 10 0 9 1 11 1 9 1 0 15 0 9 2
21 1 11 9 14 13 0 9 1 0 9 2 15 6 13 9 1 11 1 0 9 2
12 3 11 1 11 13 1 9 1 9 1 9 2
41 15 4 13 7 1 0 9 11 11 7 11 11 2 16 11 13 9 1 9 1 9 1 0 9 2 1 15 15 13 7 0 9 2 1 15 9 15 13 1 9 2
6 13 1 9 12 12 9
26 9 4 13 1 9 1 12 9 2 7 9 1 9 1 9 3 13 12 1 12 2 13 0 9 3 2
16 0 9 2 11 11 2 13 1 12 1 12 2 1 12 9 2
24 1 12 1 12 2 1 12 9 14 13 9 1 9 1 2 11 2 2 11 2 13 3 9 2
5 2 13 15 11 2
6 15 1 9 13 9 2
9 2 13 0 9 1 2 11 2 2
11 6 13 3 3 10 13 9 1 0 9 2
27 9 1 11 12 9 13 1 9 9 1 12 9 9 1 9 2 11 2 1 9 11 11 2 13 1 9 2
22 0 9 11 11 2 12 9 2 7 11 11 2 12 9 2 1 11 13 14 13 9 2
23 3 9 13 14 13 9 1 11 14 13 10 9 1 9 7 9 15 14 15 13 1 15 2
15 2 9 1 0 9 1 11 1 9 1 9 13 3 0 2
12 9 4 13 1 9 1 3 9 13 14 13 2
12 2 13 14 1 10 9 9 14 13 3 3 2
23 3 9 13 14 13 9 1 11 14 13 10 9 1 9 7 9 15 14 15 13 1 15 2
9 2 10 13 0 9 1 9 3 2
27 14 6 13 2 16 9 13 12 1 3 10 2 1 15 11 3 15 4 13 2 7 3 9 13 3 9 2
14 15 6 15 13 3 14 15 13 2 13 7 14 13 2
7 2 13 2 11 11 2 2
8 2 13 2 11 11 11 2 2
19 2 9 13 1 9 1 9 1 2 11 12 2 11 11 10 14 13 3 2
13 13 2 16 11 13 12 1 0 9 1 10 9 2
11 1 15 1 10 9 13 10 1 10 9 2
5 10 13 9 3 2
13 14 13 2 16 11 1 12 9 4 13 1 15 2
13 13 9 1 9 1 3 0 9 1 10 1 9 2
4 2 13 11 2
12 2 13 11 11 2 1 14 13 9 7 9 2
5 2 13 11 2 2
17 9 1 0 9 13 0 9 1 11 2 15 13 12 9 10 9 2
6 2 13 11 1 9 2
30 1 0 12 3 6 13 9 1 2 11 2 2 12 9 9 1 11 2 7 2 11 2 2 12 9 9 1 11 2 2
18 1 0 0 9 4 13 11 2 15 13 1 12 9 1 9 1 11 2
13 2 13 1 9 9 1 2 11 2 11 11 2 2
7 9 13 0 9 1 0 9
18 1 11 0 9 13 12 9 1 9 1 9 2 1 14 13 0 9 2
20 9 3 1 3 12 9 4 13 1 9 2 3 15 13 3 14 13 1 15 2
21 1 14 6 13 0 15 9 2 15 13 14 13 1 9 15 2 15 15 13 3 2
12 15 13 9 2 15 1 0 9 13 0 9 2
22 1 9 1 9 1 9 3 13 0 2 1 9 1 9 15 13 3 12 9 1 9 2
16 1 14 6 13 9 15 1 9 2 9 3 15 13 1 9 2
9 2 3 13 2 16 13 1 9 2
16 2 13 11 1 9 1 9 15 1 0 15 1 9 9 2 2
5 13 1 9 9 0
24 15 13 3 9 1 2 0 0 9 2 11 11 2 1 10 9 15 13 0 0 9 1 15 2
19 2 11 2 13 1 0 9 0 9 2 1 15 13 2 9 2 1 9 2
20 13 15 7 9 2 7 9 2 7 9 6 13 10 1 0 1 3 0 9 2
8 12 1 15 4 13 1 9 2
8 2 13 11 1 2 11 2 2
16 15 13 1 9 2 16 0 0 9 13 1 9 9 1 11 2
17 1 9 13 3 2 16 0 9 6 13 14 13 9 1 0 9 2
22 1 15 12 1 9 1 0 9 13 2 16 9 6 4 13 9 1 10 1 0 9 2
11 3 1 15 13 14 13 9 1 0 9 2
18 1 11 3 4 13 12 9 2 16 9 1 0 9 13 1 12 11 2
34 1 10 9 9 1 9 7 9 14 15 13 2 1 12 9 2 2 3 1 9 2 1 15 1 9 4 13 9 1 9 1 0 9 2
18 9 4 13 9 1 9 2 13 3 0 9 1 9 2 11 2 3 2
25 9 1 9 13 0 9 1 9 2 3 15 4 13 1 3 0 9 2 13 9 11 1 0 9 2
14 0 3 6 13 1 15 9 1 11 14 15 13 9 2
16 0 15 9 4 13 1 0 9 1 9 1 12 9 1 11 2
21 3 0 9 12 1 15 13 1 0 9 2 7 1 9 1 12 9 9 13 11 2
42 1 0 9 14 15 13 0 9 2 15 13 1 9 2 11 2 2 9 1 11 11 11 7 9 1 9 1 9 1 9 1 0 0 9 7 0 9 1 9 11 11 2
29 1 0 9 2 3 9 3 13 12 9 2 9 1 11 9 12 13 3 12 0 9 2 13 3 9 9 11 11 2
19 0 9 3 15 13 2 16 4 13 1 3 2 3 15 6 15 4 13 2
20 1 15 13 1 9 1 9 9 2 0 1 9 11 11 1 0 9 1 11 2
17 3 9 7 9 15 13 10 9 9 1 0 9 1 9 1 9 2
25 3 0 14 13 9 2 16 3 15 13 1 9 0 9 1 9 2 15 14 13 9 1 0 9 2
15 11 1 0 9 6 13 1 9 0 9 2 9 1 9 2
26 3 1 9 7 9 11 11 13 3 7 1 0 15 9 2 16 6 13 14 15 13 0 9 1 9 2
44 3 9 13 0 9 1 9 2 3 13 1 9 1 11 0 9 2 1 15 3 0 9 2 9 2 13 2 9 15 2 7 9 7 0 9 2 13 2 9 1 0 0 9 2
14 14 2 16 15 13 9 2 13 15 13 14 13 9 2
15 13 15 14 15 13 1 9 2 15 13 9 1 0 9 2
11 7 11 2 7 11 14 13 1 9 0 9
26 3 13 1 0 15 9 2 11 2 2 1 0 9 10 9 11 0 13 9 3 1 14 13 0 9 2
32 11 0 7 1 0 9 13 0 9 2 1 0 9 1 0 9 11 1 0 15 12 9 9 15 13 1 12 9 9 11 11 2
20 2 6 2 3 6 4 13 2 16 15 13 0 9 2 15 13 14 15 13 2
18 1 15 9 1 9 1 9 15 13 12 2 14 13 1 0 15 9 2
8 13 14 13 9 1 0 9 2
17 2 13 2 16 9 1 10 9 1 9 14 13 3 0 1 9 2
6 10 13 1 0 9 2
11 13 7 14 15 13 2 7 14 15 13 2
18 11 13 9 1 0 9 2 9 1 0 9 11 2 0 15 1 11 2
18 9 1 9 4 13 1 9 3 1 9 1 0 9 2 15 13 9 2
37 0 9 1 9 1 9 1 9 2 15 13 3 0 9 1 9 1 10 0 9 7 1 0 0 9 2 6 13 0 9 1 9 1 9 1 9 2
26 3 9 1 2 11 2 11 11 13 0 9 2 13 9 7 13 1 0 9 12 15 0 9 1 9 2
12 2 13 0 9 1 2 0 2 11 11 2 2
7 2 13 9 15 11 11 2
4 2 13 11 2
15 2 13 9 11 7 13 2 16 9 3 13 2 9 2 2
26 9 15 14 13 0 9 2 16 13 9 1 9 15 1 3 0 9 2 1 9 7 0 9 1 9 2
32 9 13 9 15 14 13 1 15 9 1 9 15 2 11 11 11 2 2 15 13 1 0 9 2 13 2 11 11 11 11 2 2
19 1 0 9 0 9 11 11 13 9 3 13 0 9 1 0 9 1 11 2
7 0 9 13 9 1 9 2
28 9 1 0 9 2 9 1 9 2 9 2 0 0 9 1 9 12 9 15 13 3 1 2 11 2 7 11 2
26 1 9 13 7 9 2 15 14 13 1 9 1 0 7 0 9 1 9 2 11 2 2 13 3 11 2
31 0 0 9 2 11 2 13 1 0 15 9 1 9 0 9 1 11 2 1 15 1 12 9 13 9 15 1 10 0 9 2
27 0 9 1 9 2 9 2 9 2 9 7 9 2 13 9 1 0 15 9 2 15 1 9 13 3 0 2
22 0 9 4 13 3 1 11 7 11 2 1 15 15 13 2 16 13 0 9 1 9 2
14 11 1 0 9 15 4 13 3 1 0 9 1 9 2
33 9 13 2 16 13 14 13 0 0 9 1 9 7 13 14 15 13 14 14 6 13 9 1 9 1 9 15 1 9 1 0 9 2
18 10 13 7 2 0 2 9 15 14 13 0 9 2 0 1 0 9 2
17 6 13 14 15 13 2 16 10 2 13 9 1 9 2 13 9 2
17 1 0 9 3 15 13 3 14 13 9 1 2 0 2 0 9 2
22 3 15 13 2 16 1 14 13 2 15 13 14 13 10 9 0 9 1 0 0 9 2
19 14 13 9 1 9 1 9 2 13 0 0 9 2 15 13 9 1 9 2
20 1 0 15 9 11 13 14 13 9 1 9 1 0 9 1 9 11 2 11 2
20 1 9 13 7 0 9 2 15 3 13 14 13 1 9 15 9 1 10 9 2
14 9 15 13 1 9 12 0 9 1 11 1 12 9 2
17 15 13 9 1 0 9 7 9 2 15 1 9 15 13 1 9 2
12 0 9 11 11 13 1 9 0 9 1 9 2
30 11 13 9 1 15 2 16 13 0 9 1 9 1 0 9 7 13 0 9 1 0 9 2 13 1 2 11 2 12 2
10 11 14 1 0 9 13 9 1 11 2
10 1 0 9 9 13 0 9 1 9 2
22 1 9 6 15 13 10 2 15 14 13 9 1 0 9 7 14 13 0 9 1 9 2
16 0 9 1 0 9 14 13 9 11 0 1 15 13 0 9 2
23 9 1 9 7 0 9 13 11 0 1 11 2 15 3 15 13 2 7 15 3 6 13 2
28 11 3 3 4 13 2 16 14 14 13 2 6 13 14 13 9 2 1 1 9 6 15 13 7 13 0 9 2
16 3 13 3 2 16 9 13 12 1 9 1 0 9 1 9 2
28 0 9 1 11 13 1 0 9 9 1 9 2 9 1 12 0 9 2 0 1 9 1 12 0 9 1 11 2
16 9 13 3 1 12 9 2 3 13 13 7 0 2 13 11 2
8 9 4 13 1 9 1 11 2
22 0 11 11 1 11 13 12 9 2 15 15 13 14 15 13 1 0 9 2 13 11 2
11 0 0 9 1 3 3 13 1 0 9 2
17 3 1 2 14 13 9 9 13 11 11 1 0 1 9 1 9 2
9 9 1 9 3 3 6 4 13 2
26 15 13 0 1 0 9 1 9 2 11 2 1 0 9 0 9 2 3 15 13 1 9 1 12 9 2
14 9 1 0 0 9 13 1 0 9 1 9 1 10 2
23 3 1 9 1 9 11 13 1 0 9 1 11 2 3 15 13 9 3 1 12 15 9 2
30 7 3 2 1 1 13 0 9 1 9 15 2 14 13 0 9 1 9 2 11 11 3 13 9 1 0 9 0 9 2
17 3 3 0 9 14 13 14 13 9 2 16 0 9 13 0 9 2
21 1 0 9 14 7 10 2 15 3 13 2 11 2 2 3 13 14 13 12 9 2
20 13 9 1 2 11 2 2 3 0 9 13 14 15 13 9 7 1 0 9 2
11 13 14 10 9 3 1 9 14 15 13 2
25 9 2 16 0 9 1 9 13 9 2 1 1 6 13 11 2 13 10 13 0 9 1 0 9 2
10 1 9 15 3 6 13 14 15 13 2
13 9 2 16 1 15 13 9 1 9 2 6 13 2
11 7 3 11 13 1 10 14 15 13 9 2
24 1 0 9 9 1 9 13 1 9 1 11 2 15 3 13 3 3 7 13 1 9 9 15 2
24 12 13 0 9 1 9 1 0 9 1 11 2 0 9 11 11 7 0 9 1 9 11 11 2
26 11 11 14 13 11 14 13 3 0 9 2 1 15 0 15 14 13 9 2 1 14 15 4 13 9 2
5 13 11 1 0 9
27 1 9 13 14 4 13 9 1 9 2 15 14 15 13 1 0 9 2 0 9 2 1 9 2 11 2 2
26 3 9 1 9 15 15 13 1 0 9 7 13 1 12 9 2 3 1 15 1 9 4 13 1 9 2
5 2 13 0 11 2
23 0 9 11 1 12 9 13 1 0 9 1 9 3 1 9 15 2 15 13 0 1 9 2
11 13 3 2 2 0 9 2 9 11 2 2
14 2 13 9 1 0 9 11 11 1 0 9 1 9 2
23 9 2 11 2 13 1 9 9 2 11 2 1 9 11 11 2 9 1 9 1 0 9 2
20 10 0 9 2 0 15 1 0 9 2 1 3 9 14 4 13 14 13 11 2
23 9 1 9 2 10 9 3 3 6 4 13 2 13 1 9 9 7 9 1 0 0 9 2
5 2 13 11 2 2
34 1 9 1 11 11 1 0 9 2 11 11 2 13 2 11 2 1 12 1 12 1 9 1 9 1 0 9 1 9 1 9 1 11 2
24 9 2 11 2 3 15 13 1 9 2 1 1 13 1 2 11 2 1 12 1 12 1 9 2
5 2 13 15 11 2
14 16 6 4 13 2 11 13 14 13 9 14 13 9 2
19 15 13 9 14 15 13 3 3 7 14 13 0 15 9 1 12 0 9 2
16 3 1 3 13 9 3 2 7 3 15 6 13 2 13 2 2
8 1 15 13 0 9 1 9 2
18 0 9 14 13 9 1 9 7 0 9 2 13 1 9 15 11 11 2
17 11 13 9 1 0 9 1 0 9 7 0 15 9 1 0 9 2
27 9 11 13 9 11 11 1 9 15 1 9 1 9 1 9 1 9 1 0 9 2 3 11 13 0 9 2
4 2 13 9 2
32 1 15 9 13 14 13 3 11 14 15 13 1 0 9 1 0 0 11 2 15 14 13 0 7 0 9 1 9 1 10 9 2
23 9 11 11 7 9 15 11 11 1 0 0 9 13 9 1 0 9 1 9 7 9 1 9
16 3 13 1 9 2 1 10 9 2 13 1 9 15 0 9 2
20 2 13 0 9 1 9 15 1 9 1 9 1 9 1 9 1 9 11 11 2
5 2 13 0 9 2
14 9 1 9 3 2 1 0 0 9 6 13 3 0 2
16 3 15 13 1 9 12 9 2 0 9 7 9 1 9 11 2
27 10 9 13 2 16 0 9 13 14 13 3 2 1 14 13 9 2 15 3 13 2 0 9 7 0 0 9
7 2 13 1 9 11 11 2
26 1 9 1 9 1 0 0 9 9 15 13 2 14 13 9 1 0 9 1 9 2 1 0 15 9 2
24 3 11 13 1 0 9 2 15 13 12 1 0 9 2 15 13 1 9 1 0 2 13 9 2
25 6 13 14 13 10 9 7 14 13 1 9 0 9 1 9 1 3 0 9 2 16 13 0 0 9
4 2 13 15 2
5 2 13 9 11 11
6 2 13 9 11 11 2
5 2 13 11 11 2
5 2 13 0 9 2
12 9 6 13 14 1 10 10 3 13 11 0 2
5 2 13 0 9 2
15 15 3 13 2 16 11 13 1 0 2 15 13 0 9 2
34 15 13 2 16 3 11 13 0 9 14 15 13 1 0 9 1 11 7 4 13 0 9 0 9 7 9 1 10 9 14 13 10 9 2
6 2 13 9 11 11 2
11 3 9 13 14 13 2 16 3 13 3 2
7 11 4 13 9 1 0 9
12 9 13 10 2 3 13 0 9 1 0 9 2
4 2 13 11 2
21 0 9 11 11 13 1 0 9 0 9 2 1 9 2 0 1 2 11 3 2 2
4 2 13 11 2
18 9 15 13 1 9 1 10 9 9 2 15 13 2 16 15 13 9 2
4 2 13 11 2
23 10 13 9 1 3 9 2 0 1 9 1 9 1 0 9 1 9 1 11 2 11 2 2
19 1 7 3 0 1 9 1 9 1 9 2 11 11 6 13 3 1 9 2
18 13 9 2 16 3 9 13 1 9 1 9 9 2 15 13 10 9 2
7 12 1 15 4 3 13 2
12 1 15 9 7 1 12 9 13 7 15 13 2
4 2 13 11 2
4 2 13 9 2
23 1 9 1 9 1 9 11 2 10 9 4 4 13 3 14 13 1 9 1 9 0 9 2
4 2 13 11 2
11 3 15 13 14 13 2 16 4 13 3 2
5 2 13 0 9 2
26 3 7 15 13 9 2 2 15 4 4 13 1 9 1 10 0 9 2 7 6 4 15 13 9 2 2
4 2 13 11 2
4 2 13 15 2
14 15 13 2 16 11 1 9 13 1 9 2 11 2 2
18 9 13 3 0 9 2 7 11 2 7 11 4 13 1 10 9 1 9
4 2 13 11 2
4 2 13 11 2
4 2 13 11 2
9 2 13 9 11 11 3 1 9 2
40 3 3 0 13 2 1 9 1 9 2 14 13 0 0 9 1 9 1 9 2 1 15 14 4 13 0 9 14 15 15 13 2 16 3 13 14 15 13 9 2
10 2 13 9 1 9 1 9 11 11 2
16 2 13 11 1 9 1 9 10 14 13 9 1 0 0 9 2
18 15 13 7 11 3 15 13 2 16 15 6 4 13 2 16 14 13 9
7 2 13 0 1 0 9 2
31 3 11 13 3 12 9 9 7 1 0 9 13 1 9 1 9 7 15 13 2 16 9 3 4 13 9 14 13 0 9 2
32 13 9 9 2 16 9 1 0 9 1 11 4 13 1 9 1 0 9 2 13 3 11 11 2 7 6 13 0 9 1 9 2
4 2 13 11 2
10 2 15 1 9 1 9 6 4 13 2
22 15 13 0 9 7 13 1 0 10 9 2 15 15 13 2 14 13 1 3 0 9 2
8 7 15 13 0 1 9 15 2
5 6 2 15 13 2
19 0 0 9 13 14 13 1 0 9 0 9 1 9 11 11 2 0 11 2
11 2 13 11 11 2 9 1 9 1 11 2
20 0 9 15 13 14 13 9 2 15 15 13 1 12 1 0 9 1 0 9 2
4 2 13 11 2
9 2 13 11 11 1 9 1 9 2
7 11 13 1 9 2 11 2
27 9 1 11 11 11 13 9 1 9 1 2 11 2 1 0 9 1 9 1 9 1 11 1 2 11 2 2
17 13 3 0 9 1 9 11 11 7 13 3 9 1 2 11 2 2
4 2 13 11 2
4 2 13 11 2
9 2 13 11 1 9 2 11 2 2
17 10 9 13 14 13 7 14 13 2 16 9 15 14 15 13 3 2
28 3 9 2 15 15 13 1 0 9 1 2 0 2 2 3 4 13 1 0 9 1 9 1 9 2 9 2 2
30 1 9 1 9 2 11 11 2 13 3 2 16 1 3 3 4 4 13 10 9 1 9 2 9 2 7 2 9 2 2
12 9 14 4 13 3 9 1 0 9 1 9 2
8 11 3 13 0 1 11 1 11
12 0 13 1 2 9 2 9 2 1 12 9 2
9 2 13 0 9 1 2 11 2 2
22 1 12 9 13 3 2 16 12 1 3 0 2 11 11 2 13 9 1 2 11 2 2
15 3 1 9 13 2 16 14 13 1 0 9 9 1 9 2
15 9 7 0 9 14 13 1 0 9 0 9 2 11 2 2
20 1 9 1 10 9 14 15 13 9 12 12 2 0 15 9 13 9 12 9 2
10 0 0 9 13 12 1 0 1 11 2
26 3 13 12 0 9 2 7 0 1 15 4 13 1 9 1 0 9 2 1 14 4 13 2 11 2 2
28 9 1 9 13 9 1 9 14 13 0 7 2 16 13 12 9 9 2 9 14 15 13 1 0 9 1 11 2
31 9 1 0 9 13 9 1 12 9 9 14 13 3 1 12 9 1 9 1 0 9 2 7 9 14 15 13 1 0 11 2
14 13 3 14 13 1 2 11 2 7 14 13 1 9 2
4 2 13 11 2
7 2 13 0 9 11 11 2
21 9 2 11 2 7 11 15 13 14 13 0 9 11 11 2 13 0 1 12 9 2
18 11 13 14 13 1 0 15 9 2 7 13 9 14 13 9 1 15 2
26 3 3 15 6 4 13 3 9 15 1 11 2 15 13 10 9 14 15 13 3 1 11 1 10 9 2
15 2 0 9 13 14 13 1 0 9 7 14 6 15 13 2
4 13 9 1 9
5 2 13 1 9 2
14 15 13 10 9 14 13 9 1 2 11 2 1 9 2
4 2 13 9 2
13 1 15 14 13 9 1 9 1 2 11 2 1 3
4 2 13 15 2
6 2 13 9 1 9 2
12 10 13 9 1 0 0 9 1 9 1 9 2
40 1 9 15 13 2 16 10 9 2 10 9 1 9 1 9 2 0 9 7 9 14 13 0 9 13 3 9 2 15 6 13 0 2 7 4 4 1 9 13 2
5 3 13 14 13 2
33 0 0 9 2 15 6 13 9 15 14 13 7 13 0 1 9 9 2 9 1 9 2 2 14 13 7 1 9 1 11 1 11 2
37 1 9 1 10 9 9 13 9 1 9 1 0 9 1 9 1 9 11 2 7 1 9 14 15 13 1 0 9 1 0 2 0 11 2 1 11 2
37 1 9 1 10 9 9 13 9 1 9 1 0 9 1 9 1 9 11 2 7 1 9 14 15 13 1 0 9 1 0 2 0 11 2 1 11 2
13 1 9 4 13 3 7 0 15 1 9 0 9 2
22 0 9 11 11 13 3 2 16 13 0 9 15 13 1 0 9 2 7 6 15 13 2
20 1 9 0 9 11 11 3 13 2 16 13 0 9 2 15 13 14 15 13 2
20 9 13 2 16 9 1 9 4 13 3 9 1 0 1 9 1 9 1 11 2
18 9 13 2 16 12 9 1 9 14 13 1 9 1 14 13 12 9 2
22 0 9 13 1 9 0 9 11 12 1 0 9 2 11 2 1 12 3 2 13 11 2
9 6 13 14 15 13 10 14 13 2
17 6 4 13 9 7 9 2 7 9 11 3 13 2 13 15 2 2
13 13 14 13 2 16 15 13 0 9 1 0 9 2
17 15 4 13 9 14 15 13 0 9 2 11 2 15 13 1 9 2
20 0 3 1 9 9 1 11 3 15 4 13 2 13 3 1 0 9 1 11 2
26 0 9 2 15 13 7 0 9 2 13 0 9 1 0 0 9 1 9 2 0 9 2 1 9 11 2
37 9 1 11 11 3 3 4 13 1 9 1 2 9 2 1 11 2 1 15 0 9 1 11 13 12 9 9 7 4 13 1 0 9 1 0 9 2
21 15 13 2 16 2 6 13 1 11 2 2 9 1 9 4 13 7 13 0 9 2
13 2 11 2 13 9 2 3 13 9 1 3 0 2
12 16 6 13 1 12 9 9 2 14 13 7 15
4 2 13 11 2
40 10 9 1 0 2 0 9 2 2 15 6 13 1 9 2 1 9 9 1 0 9 1 9 15 13 1 9 15 1 0 9 1 0 1 11 2 11 2 9 2
12 2 13 9 1 0 9 1 0 9 11 11 2
13 15 13 0 0 9 1 10 2 15 13 1 11 2
25 9 13 14 15 13 1 9 2 15 4 13 1 9 0 9 2 1 10 9 2 7 1 0 9 2
19 9 13 0 9 7 0 0 9 14 13 1 0 9 7 10 9 1 9 2
31 0 9 1 2 0 2 11 11 13 1 9 2 16 9 14 13 1 9 1 0 9 7 16 13 2 9 15 14 13 9 2
8 11 13 2 11 2 9 1 9
18 0 2 0 7 0 4 3 13 1 9 1 9 2 15 13 1 11 2
12 1 0 15 9 13 14 13 7 9 1 9 2
5 2 13 0 9 2
25 1 0 9 13 14 6 15 13 9 1 0 9 2 14 6 15 13 9 7 3 14 15 13 9 2
6 0 13 1 12 1 12
23 1 0 9 1 11 15 13 0 0 9 1 9 1 0 9 7 1 9 14 15 13 3 2
13 1 9 1 11 15 13 1 10 11 0 0 9 2
30 1 9 9 1 11 11 11 11 13 1 11 7 3 13 14 13 9 2 16 3 1 11 3 11 14 13 1 0 9 2
16 15 13 3 2 16 11 13 9 2 15 6 13 9 1 9 2
15 13 7 3 3 1 9 1 9 2 3 13 1 0 9 2
18 9 1 0 0 9 1 9 15 13 1 9 2 13 1 0 9 2 2
21 9 1 11 13 1 9 7 1 15 6 15 13 2 9 2 14 15 13 1 11 2
27 14 6 13 2 16 11 3 6 15 4 13 9 1 11 2 7 11 11 1 0 9 13 9 1 3 0 2
46 3 1 9 15 13 2 16 1 0 0 9 1 15 15 13 2 16 1 0 15 9 3 11 7 11 13 14 15 13 10 9 1 9 7 16 11 13 14 15 13 11 1 10 0 11 2
33 1 9 1 11 1 0 9 7 1 9 1 11 7 11 1 9 0 0 9 3 6 15 13 15 13 10 0 9 1 9 1 9 2
22 3 3 9 14 13 9 14 13 10 13 1 15 2 16 15 13 9 14 13 1 9 2
20 0 0 9 6 15 13 3 1 9 1 15 7 1 10 10 13 9 1 11 2
26 3 3 11 13 1 9 7 10 9 13 0 9 1 0 0 9 2 3 1 15 1 9 13 7 9 2
19 2 14 13 15 0 7 0 9 2 2 13 15 2 13 15 14 13 9 2
13 1 9 13 1 9 1 0 0 9 2 11 2 2
23 11 3 13 9 2 15 13 9 1 9 1 9 2 13 15 1 0 9 2 0 1 9 2
15 1 9 1 9 15 13 3 4 13 11 7 3 4 13 2
12 9 13 9 1 0 9 1 9 1 0 9 2
4 2 13 15 2
19 13 15 11 7 15 13 14 15 13 1 11 2 7 1 9 14 6 13 2
12 1 11 0 13 0 2 1 10 9 10 13 2
4 2 13 9 2
15 10 14 13 2 3 1 3 0 13 2 13 4 1 9 3
5 2 13 15 11 2
4 2 13 15 2
8 2 13 1 0 15 9 11 2
4 2 13 15 2
5 2 13 15 11 2
9 2 13 15 7 15 13 1 9 2
4 2 13 11 2
4 2 13 15 2
20 16 13 2 16 15 13 2 1 9 15 13 7 13 0 2 13 1 9 3 2
21 7 13 3 9 15 11 9 15 13 3 9 13 10 11 2 10 15 13 7 13 2
5 2 13 15 11 2
12 1 0 9 1 9 3 13 1 0 9 9 2
8 2 13 15 3 9 7 9 2
18 9 1 10 9 13 10 1 9 1 9 1 2 11 2 1 0 9 2
26 9 3 13 0 9 2 3 4 13 9 9 1 0 9 7 15 13 12 9 3 2 1 9 1 9 2
10 11 11 13 1 9 9 1 2 11 2
34 9 1 2 11 2 2 11 2 11 11 2 15 3 13 9 1 0 2 11 2 2 3 15 13 1 9 1 2 0 2 1 9 9 2
21 13 14 15 13 2 16 9 9 2 9 1 9 13 12 1 12 1 9 1 9 2
32 15 4 13 9 15 3 2 13 14 15 13 1 9 9 9 1 12 9 7 14 13 1 9 1 12 9 7 9 1 12 9 2
16 2 13 15 2 2 3 13 15 7 13 1 9 9 15 9 2
16 11 11 13 9 1 0 15 9 7 2 13 4 11 9 2 2
13 13 14 9 2 1 0 9 13 3 14 13 1 9
29 1 10 9 9 1 11 9 11 7 9 13 0 9 1 9 2 13 15 1 9 2 13 1 15 7 3 13 9 2
21 3 15 13 2 11 13 2 3 13 14 13 9 15 2 13 15 3 1 9 2 2
7 2 13 0 9 11 11 2
6 3 1 0 13 9 2
19 1 9 15 7 9 15 13 10 4 13 2 7 7 1 9 13 10 13 2
35 9 1 0 9 2 11 2 1 9 11 11 13 1 9 2 1 1 0 9 13 1 0 9 1 12 9 1 9 14 15 13 1 9 15 2
23 15 4 13 9 7 15 13 14 13 1 0 9 2 1 14 13 9 14 4 13 1 11 2
50 1 9 1 0 9 1 0 9 1 0 1 9 9 14 15 13 9 1 9 1 9 7 9 13 1 9 2 16 16 6 13 14 13 9 1 9 2 10 2 15 15 13 2 15 13 14 15 13 9 2
18 13 9 9 14 15 13 14 13 0 2 0 7 6 3 0 0 9 2
16 3 1 9 0 9 4 13 14 13 1 0 9 7 0 9 2
21 3 13 0 9 1 0 7 0 0 9 7 9 2 15 3 3 14 13 0 9 2
24 15 13 14 15 13 7 1 9 1 0 0 9 1 9 2 11 2 2 14 15 13 7 13 2
12 1 0 9 9 13 14 13 0 1 0 9 2
9 9 13 9 1 2 11 2 1 11
31 9 11 11 13 12 9 1 9 1 2 11 2 1 2 11 2 1 12 1 12 1 9 1 0 9 1 11 1 0 9 2
31 10 9 13 0 9 2 9 1 9 2 15 13 2 1 9 0 2 2 0 9 7 9 2 16 2 9 6 13 9 2 2
16 13 0 9 1 0 15 9 2 15 14 4 13 1 0 9 2
19 14 0 9 1 0 15 9 14 15 13 3 1 9 14 13 0 0 9 2
28 14 14 13 1 0 9 0 9 2 16 0 15 9 2 15 13 0 9 2 13 10 2 15 13 1 9 15 2
14 1 9 3 1 9 15 13 11 11 1 2 11 2 2
38 2 11 2 2 11 2 2 3 9 13 0 9 11 11 2 13 1 0 9 1 9 1 9 1 11 1 9 1 12 1 12 1 0 0 2 11 2 2
23 0 0 9 11 11 11 4 3 13 1 9 2 0 1 0 11 2 1 0 2 11 2 2
23 0 0 9 11 11 11 4 3 13 1 9 2 0 1 0 11 2 1 0 2 11 2 2
26 1 9 2 11 2 2 15 1 9 1 11 13 9 1 11 2 3 13 1 9 1 9 2 11 2 2
28 1 0 9 14 13 1 11 13 9 11 2 15 13 12 9 1 2 11 2 2 11 2 1 9 1 0 9 2
10 2 13 9 1 2 11 2 11 11 2
25 9 13 3 1 9 1 0 9 1 11 2 9 12 12 2 2 7 3 1 9 15 13 11 11 2
21 3 1 15 1 9 1 11 14 13 9 2 1 16 0 9 6 13 10 1 9 2
24 1 9 1 0 9 14 15 13 3 7 10 9 1 0 9 2 15 15 13 1 9 1 9 2
31 9 1 9 7 9 14 15 13 2 1 10 9 2 2 3 1 9 2 1 15 1 9 4 13 9 1 9 1 0 9 2
27 0 9 11 11 13 1 0 9 9 2 1 15 13 9 7 13 0 0 9 1 0 9 2 13 0 9 2
6 2 4 13 11 11 11
12 15 13 9 1 11 7 4 13 9 1 9 2
8 2 13 1 9 15 0 9 2
4 2 13 11 2
13 10 1 0 9 1 9 13 0 9 1 0 9 2
20 9 15 13 1 9 2 15 13 14 15 13 0 9 2 15 1 9 13 9 2
18 0 0 9 1 11 11 11 13 3 12 9 1 2 11 2 11 2 2
16 1 0 12 9 0 9 11 11 13 9 1 3 1 12 9 2
18 11 11 13 0 9 14 13 0 2 9 3 1 9 15 13 1 9 2
16 2 11 2 13 2 11 2 1 12 1 12 1 9 1 11 2
18 1 9 0 2 1 0 0 9 2 13 9 11 11 1 9 12 9 2
16 3 12 9 2 3 12 9 2 13 3 3 1 9 1 9 2
32 1 9 1 0 0 9 11 11 9 1 9 14 13 9 1 0 9 1 9 7 14 13 1 9 0 9 1 9 1 0 9 2
23 1 9 13 14 13 0 0 9 1 0 9 2 9 2 9 2 0 9 7 9 2 13 9
20 0 9 1 11 1 3 0 9 13 1 0 9 1 10 0 7 0 0 9 2
34 0 9 1 10 9 13 0 7 15 13 2 16 9 13 14 13 7 13 0 9 2 1 14 15 13 9 2 16 15 13 10 4 13 2
24 15 1 0 9 13 9 1 11 7 13 9 1 3 0 9 2 3 1 0 9 1 0 9 2
17 2 10 2 16 15 1 9 13 9 1 9 2 6 13 3 15 2
44 2 13 14 10 9 1 9 1 9 2 1 0 9 7 1 0 9 2 7 1 9 1 9 2 1 9 7 1 9 2 14 13 1 0 1 15 9 0 0 9 1 0 9 2
17 2 6 13 9 2 16 0 9 13 14 13 0 9 1 0 9 2
16 9 1 0 9 3 15 3 13 1 0 15 9 2 1 9 2
15 1 16 9 15 14 13 10 9 4 3 13 1 0 9 2
5 15 13 10 3 2
10 10 1 9 13 2 16 9 13 9 2
20 11 11 13 9 1 2 11 2 2 7 9 13 9 11 11 1 2 11 2 2
9 13 14 13 3 10 1 2 11 2
8 2 13 1 0 9 11 2 2
17 9 13 1 9 9 1 9 1 11 0 9 1 9 1 0 9 2
4 2 13 11 2
40 9 1 0 9 1 0 9 14 13 9 7 1 10 9 2 1 15 14 13 12 0 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 0 11 2
15 12 9 13 0 9 1 0 9 1 0 9 1 0 9 2
26 9 1 0 2 11 2 11 11 4 13 1 0 9 1 0 9 1 10 1 0 9 1 9 1 9 2
19 2 11 2 1 12 9 13 2 12 9 1 9 2 15 15 13 9 2 2
48 9 13 0 9 2 12 12 0 0 9 2 0 0 9 2 9 1 12 9 1 9 2 9 1 0 9 2 9 1 9 1 0 9 1 11 2 9 1 9 1 9 1 11 7 9 1 9 2
10 7 13 14 15 13 10 15 13 3 2
14 15 13 9 7 15 13 9 14 13 2 16 13 9 2
19 14 14 15 13 0 9 2 13 15 14 13 2 16 4 13 9 1 9 2
10 2 13 9 1 2 9 2 11 11 2
5 11 11 13 12 2
16 1 2 11 2 11 11 13 12 9 2 7 11 11 13 12 2
32 0 9 1 0 9 1 0 9 1 0 9 1 11 2 1 0 11 7 0 9 2 14 4 13 1 9 1 9 1 0 9 2
13 9 3 15 13 2 16 1 0 9 14 13 0 2
19 1 9 1 10 9 9 1 9 7 9 13 0 1 9 7 15 13 10 2
17 3 9 1 10 9 6 13 3 0 2 1 14 6 13 10 3 2
18 3 9 7 9 15 13 3 1 15 2 16 14 13 0 1 0 9 2
15 1 10 9 15 13 0 9 1 0 9 1 9 1 15 2
15 15 13 14 13 3 0 0 0 9 10 13 2 11 2 2
11 11 1 9 9 1 11 3 13 0 9 2
16 16 0 9 13 14 13 9 15 2 14 13 9 1 12 9 2
20 3 1 0 9 0 9 1 9 1 2 11 2 13 1 9 11 12 9 1 9
13 2 10 1 10 9 13 14 9 1 2 11 2 2
5 15 13 15 10 2
14 0 9 13 7 1 0 7 0 9 10 0 0 9 2
31 0 9 1 0 9 2 0 9 7 9 1 2 11 2 2 11 13 10 1 0 9 1 9 1 0 9 0 2 0 9 2
17 2 13 1 0 9 0 1 9 1 0 9 9 1 9 11 11 2
16 15 13 9 1 9 2 15 4 15 13 14 13 9 1 9 2
24 12 1 0 9 1 9 2 11 2 13 9 1 2 9 2 2 11 1 9 1 9 1 9 2
26 9 13 1 0 9 0 9 2 3 0 0 9 11 11 3 13 1 0 9 2 16 9 14 4 13 2
4 2 13 9 2
15 15 13 1 2 9 2 3 9 1 9 7 9 11 11 2
19 15 3 13 2 16 11 6 4 13 9 2 1 15 15 13 1 0 9 2
20 1 9 13 3 2 16 9 1 9 1 11 1 0 11 13 1 9 1 11 2
22 3 11 11 13 1 2 9 2 9 2 16 1 9 1 9 4 13 14 15 13 9 2
27 9 1 9 1 9 1 9 3 14 13 7 9 15 1 11 1 9 2 11 2 2 15 13 3 1 11 2
36 0 9 1 9 13 3 3 1 9 1 0 9 1 0 0 9 7 1 10 9 11 11 14 13 9 1 9 2 13 9 2 11 11 11 2 2
27 13 15 7 9 10 0 9 14 13 10 9 1 0 9 1 2 11 2 2 13 0 9 1 11 11 11 2
27 9 1 9 1 9 7 9 15 13 10 9 7 9 3 15 13 1 0 9 2 15 13 1 9 7 9 2
13 1 9 9 13 9 1 9 1 0 9 1 9 2
14 3 12 1 12 1 0 0 9 15 13 1 0 9 2
13 1 9 3 9 13 10 9 1 9 1 0 9 2
12 1 12 9 10 1 15 6 4 13 1 0 2
22 11 13 3 9 1 9 1 10 1 9 1 11 1 9 1 9 2 13 9 1 0 2
18 1 0 12 12 9 13 14 13 14 13 9 15 1 9 2 13 15 2
9 11 1 11 13 0 9 1 11 2
22 0 9 14 4 13 14 15 13 0 9 1 0 9 1 0 9 7 1 0 0 9 2
21 3 11 13 1 9 0 1 9 9 7 13 15 14 4 13 1 0 9 1 15 2
18 9 1 9 2 15 13 1 12 9 1 15 2 15 13 3 0 9 2
4 2 13 11 2
4 2 13 11 2
7 10 9 13 1 9 9 2
4 2 13 11 2
4 2 13 9 2
26 9 13 2 16 1 9 1 9 11 13 9 1 9 1 9 7 15 4 13 14 13 10 1 0 9 2
4 2 13 9 2
34 1 15 13 2 16 10 9 1 11 7 10 9 2 14 13 0 9 1 0 9 1 11 7 0 9 2 15 14 13 10 9 1 9 2
17 13 2 16 11 1 9 15 3 3 13 14 13 9 1 10 9 2
42 11 6 1 9 1 9 2 15 14 13 1 0 0 9 2 7 1 9 1 9 1 11 2 1 9 1 11 2 13 14 13 1 10 0 9 2 1 10 0 0 9 2
21 10 2 16 11 4 13 14 13 0 9 1 9 1 11 13 9 15 1 0 9 2
13 15 13 1 3 0 9 9 1 9 1 0 9 2
27 3 3 7 3 1 9 15 13 1 15 9 14 4 13 3 9 1 9 2 9 1 9 1 9 1 9 2
21 7 1 9 1 10 9 1 9 15 1 9 7 3 13 9 1 9 9 11 11 2
9 15 6 13 1 10 0 9 11 2
16 15 3 4 13 2 16 6 13 14 13 0 9 3 1 11 2
22 13 0 15 0 9 1 0 2 7 0 9 1 9 1 11 13 3 9 2 13 11 2
18 13 9 1 9 1 9 1 15 2 15 13 2 7 9 2 13 9 2
36 16 11 3 15 13 1 9 2 1 15 13 2 15 14 13 1 9 2 1 15 9 2 0 1 9 2 13 1 9 1 0 9 2 13 11 2
11 2 10 13 9 2 15 13 14 13 11 2
5 2 10 13 15 2
41 15 13 2 16 15 4 13 14 13 1 9 7 9 2 16 15 13 3 0 9 1 11 2 16 9 1 9 13 3 14 13 2 7 6 14 13 9 1 0 9 2
13 9 1 9 12 9 13 0 9 0 9 1 11 2
20 0 9 13 14 13 1 0 9 7 14 13 1 9 1 9 1 11 1 9 2
16 9 15 13 14 13 0 9 1 0 9 1 9 2 13 9 2
22 0 9 13 7 1 9 1 11 2 3 15 13 3 7 0 9 2 13 3 9 11 2
24 9 11 2 15 13 0 7 13 14 15 13 1 10 0 10 9 7 14 13 1 9 1 10 9
4 2 13 9 2
14 11 13 14 13 9 1 9 7 9 2 13 3 11 2
8 0 1 9 2 11 11 13 2
14 9 13 1 9 11 2 15 13 0 1 9 1 11 2
11 1 9 1 9 1 9 15 13 7 0 2
14 0 1 0 9 13 12 2 12 1 15 13 0 9 2
32 1 9 11 3 0 1 9 7 0 9 2 0 3 1 9 2 13 1 9 9 1 0 15 9 7 13 1 9 7 0 9 2
36 1 9 1 9 1 9 1 11 4 13 2 16 1 9 1 11 9 6 4 13 10 0 0 9 1 11 2 13 3 0 9 1 11 11 11 2
25 13 14 13 0 9 1 9 2 7 9 1 0 15 9 6 13 14 13 1 9 1 9 15 1 11
4 2 13 15 2
17 1 9 1 9 11 13 14 15 13 2 16 14 13 1 0 9 2
39 0 9 13 14 13 9 1 0 9 2 14 13 9 1 0 9 1 0 1 15 9 7 14 13 1 9 15 1 9 1 9 1 11 2 15 13 1 9 2
31 9 15 13 2 16 0 9 13 14 13 2 16 9 12 1 11 2 1 15 4 13 9 1 11 2 13 9 1 0 9 2
34 1 0 9 2 0 1 0 2 0 0 9 2 2 15 13 2 16 9 1 0 0 9 11 13 9 1 9 14 13 9 1 0 9 2
16 11 13 9 1 10 9 1 3 0 1 0 9 1 9 9 2
29 9 1 9 3 6 15 13 1 9 1 9 1 11 2 14 1 0 9 1 10 9 1 9 1 10 1 0 9 2
69 16 15 6 13 0 9 2 15 14 13 0 0 9 1 0 15 9 13 3 3 1 0 9 2 9 1 9 1 0 0 9 2 10 13 0 15 9 2 15 13 1 10 14 13 9 1 9 10 9 1 11 2 7 15 3 6 13 0 9 1 9 3 14 15 13 9 1 9 2
41 13 15 14 13 11 11 1 9 1 9 1 0 9 11 11 2 15 13 9 2 3 15 1 0 9 2 7 14 13 2 16 9 1 9 14 15 13 1 9 9 2
21 14 15 13 11 1 3 9 13 3 0 9 2 15 3 13 14 13 9 1 11 2
7 11 13 1 9 0 9 2
21 15 13 0 9 2 15 1 9 1 0 0 9 4 4 13 3 14 13 1 11 2
39 3 13 14 13 2 16 1 10 9 11 11 13 0 0 9 1 9 1 10 9 1 9 1 0 0 9 2 0 9 1 9 7 0 9 1 9 1 11 2
21 11 11 15 13 1 9 7 9 1 9 7 15 13 10 1 0 0 9 1 11 2
11 9 2 11 2 3 3 15 13 1 9 2
26 3 11 13 11 11 1 9 1 3 12 9 11 2 15 9 4 13 1 11 1 9 1 9 1 9 2
5 2 13 11 11 2
20 3 13 3 2 10 9 3 3 13 9 1 9 2 15 6 13 9 1 9 2
20 13 14 15 13 2 16 3 0 9 14 13 9 1 9 1 0 9 1 11 2
28 3 6 13 3 14 7 0 15 6 13 0 9 1 9 15 2 16 11 6 4 13 9 15 1 9 7 9 2
13 1 9 0 9 4 13 1 9 1 9 1 9 2
5 2 13 11 11 2
15 12 1 11 7 11 15 13 9 1 9 1 0 7 0 9
11 2 13 9 1 2 6 2 10 11 2 2
13 0 9 3 3 13 0 9 1 11 7 15 13 2
30 10 9 2 3 9 13 0 0 9 1 11 2 15 13 14 13 0 15 9 1 9 1 0 9 1 15 1 0 9 2
15 3 11 11 15 13 2 16 13 10 1 9 1 10 9 2
19 1 11 9 3 13 0 9 2 16 9 1 9 1 11 11 13 3 9 2
33 1 10 9 1 9 15 11 11 2 0 1 9 1 0 15 9 11 1 0 9 2 15 13 9 1 10 9 1 0 7 0 9 2
39 9 2 10 0 9 2 2 4 13 2 16 15 13 1 9 1 9 2 7 3 9 13 9 2 15 3 13 14 13 2 16 1 15 4 13 14 15 13 2
20 10 7 14 13 9 1 11 2 15 3 13 0 0 9 1 11 2 15 13 2
18 1 12 1 9 9 13 2 16 2 13 1 12 1 0 0 9 2 2
15 11 4 13 9 1 10 9 2 10 9 13 14 15 13 2
27 9 4 13 11 11 11 7 13 12 9 1 11 1 12 9 2 16 9 15 13 1 10 1 11 7 11 2
18 13 14 13 0 7 0 9 1 9 1 9 1 9 1 9 1 9 2
8 2 1 15 13 12 0 9 2
15 12 1 12 13 0 2 12 9 13 0 7 0 1 9 2
21 13 14 2 1 9 15 13 7 9 2 15 1 0 9 13 1 0 9 1 9 2
6 2 13 9 1 9 2
20 13 4 9 2 15 13 14 13 1 15 2 1 1 13 2 14 6 4 13 2
9 2 10 14 13 9 1 10 9 2
5 10 13 9 15 2
10 2 6 13 14 13 2 16 13 0 2
33 16 13 0 9 2 13 3 14 13 9 7 1 0 9 2 7 1 9 2 3 6 13 14 15 13 3 1 10 3 14 15 13 2
12 6 13 3 14 13 0 9 1 9 1 9 2
19 3 16 1 9 1 9 2 15 13 1 9 15 12 2 9 2 1 11 2
30 15 15 13 9 2 16 15 13 7 14 13 3 1 10 9 7 13 14 13 1 0 9 2 15 4 15 13 10 9 2
13 7 9 13 9 14 13 9 1 10 7 0 9 2
18 15 15 13 1 0 9 2 15 14 13 9 15 1 10 1 0 9 2
22 7 2 1 14 6 15 13 3 3 1 9 2 13 3 14 13 9 7 9 1 9 2
24 0 13 14 15 13 1 9 1 9 15 2 15 3 4 13 1 0 9 1 0 9 7 0 9
18 1 0 9 9 1 11 4 13 12 1 12 1 9 1 0 0 9 2
23 10 2 16 15 13 6 13 0 15 9 2 9 1 15 3 13 1 11 2 13 0 9 2
16 11 3 3 15 13 1 10 0 9 1 2 9 1 9 2 2
12 10 13 9 7 1 11 2 0 11 7 0 2
24 15 10 9 13 14 15 13 7 14 13 1 9 1 0 9 2 7 13 9 1 9 9 9 2
21 15 15 13 1 9 1 9 1 0 9 2 15 1 9 13 0 9 1 0 9 2
25 0 9 1 9 1 11 1 9 1 9 1 9 13 9 14 13 0 0 9 1 9 1 9 15 2
23 3 0 9 13 9 1 9 2 9 1 9 1 9 2 2 15 1 9 13 1 0 9 2
18 15 3 13 9 1 10 12 9 1 10 9 1 9 1 9 1 11 2
8 1 15 3 12 15 13 0 2
26 9 9 1 0 9 4 13 9 1 9 1 0 9 2 15 3 7 1 0 9 13 1 9 7 13 2
5 2 13 3 11 2
6 2 13 0 11 11 2
21 9 2 15 13 3 1 0 9 2 13 14 15 13 9 2 1 9 14 4 13 2
13 0 9 13 0 2 13 11 7 11 11 1 11 2
5 2 13 11 11 2
5 2 13 15 9 2
18 1 15 1 9 15 13 3 1 9 1 0 9 11 11 1 12 9 2
20 9 1 11 7 2 11 2 13 1 15 9 1 9 1 9 1 9 1 11 2
24 2 11 2 13 9 15 1 9 1 11 14 15 13 9 14 13 9 9 1 1 15 4 13 2
9 2 13 9 1 0 9 11 11 2
22 1 15 15 14 4 13 2 1 14 13 3 9 1 9 14 13 1 0 9 1 9 2
23 15 13 1 0 0 9 1 11 1 11 2 15 13 1 12 9 1 2 11 2 12 3 2
37 9 11 11 7 9 15 11 11 4 13 1 11 1 9 1 9 2 1 15 13 7 0 9 1 0 9 2 13 1 9 9 7 0 9 11 11 2
7 9 1 9 13 9 1 11
31 15 14 13 9 1 9 1 0 9 2 16 15 13 0 0 9 1 9 1 0 9 2 13 15 0 9 1 11 11 11 2
30 11 13 10 9 1 9 9 1 9 1 11 1 9 1 0 9 11 11 11 14 6 13 1 9 9 1 11 7 11 2
41 11 13 3 3 0 15 9 7 9 15 1 9 1 9 1 11 7 6 13 2 16 15 13 1 0 9 1 0 9 2 0 15 3 1 9 1 9 2 13 11 2
24 15 13 1 0 9 9 1 0 9 1 11 1 11 2 11 2 3 7 9 1 9 1 11 2
53 15 13 2 16 1 9 4 13 0 9 1 0 0 9 11 11 2 0 15 1 9 1 9 1 9 1 9 1 9 7 9 1 0 9 2 3 7 16 1 0 9 4 13 1 0 9 1 12 9 9 1 9 2
23 15 13 2 16 1 0 9 0 9 14 13 3 1 10 9 7 3 10 13 10 0 9 2
14 3 13 9 1 0 9 2 13 1 9 9 11 11 2
11 1 2 11 2 12 13 1 9 10 9 2
11 9 13 1 9 7 9 9 1 9 11 2
28 10 9 1 0 4 13 14 13 1 10 0 9 9 7 9 1 9 1 0 0 7 0 9 2 13 1 9 2
21 2 10 13 10 9 1 9 1 9 1 9 1 0 9 1 0 9 9 11 11 2
15 13 2 16 15 3 4 13 2 16 3 15 13 10 9 2
16 15 13 2 16 11 3 13 2 16 13 3 1 3 0 9 2
14 3 13 1 10 9 11 3 14 13 3 3 10 9 2
7 2 1 15 13 9 15 2
18 2 10 13 9 1 9 1 9 1 9 15 1 9 1 9 1 9 2
28 13 3 1 9 15 9 1 9 1 9 2 15 15 15 13 3 2 1 14 13 10 13 9 15 14 15 13 2
25 13 9 1 9 2 11 2 2 15 13 1 0 0 9 2 3 7 1 11 0 1 11 2 11 2
23 1 0 9 1 9 6 4 13 9 1 9 1 9 2 3 16 10 9 3 3 6 13 2
8 12 1 12 1 9 13 1 9
21 13 12 9 1 9 2 15 14 15 13 10 9 1 0 9 2 14 6 13 9 2
21 0 9 11 1 0 9 4 13 1 11 2 1 1 0 9 15 13 1 0 9 2
5 2 13 9 11 2
12 1 0 11 13 1 9 15 1 9 9 11 2
15 15 13 11 11 1 9 1 0 9 7 9 1 0 9 2
11 15 13 9 1 9 1 15 2 13 11 2
19 3 3 15 13 9 14 13 9 1 9 1 9 11 2 15 13 1 9 2
17 3 13 2 16 13 14 13 14 13 9 2 1 14 15 13 9 2
16 10 9 1 0 9 13 14 4 13 0 1 9 1 0 9 2
22 16 9 4 13 1 9 1 9 0 9 2 15 4 13 1 0 9 9 1 9 15 2
21 15 4 13 1 0 9 0 9 2 15 4 13 14 13 1 9 3 12 10 9 2
25 7 15 13 1 10 9 2 1 15 13 9 1 9 15 2 11 2 1 3 0 2 2 11 2 2
7 9 9 3 3 13 11 2
26 9 1 9 1 9 1 9 7 9 4 13 14 1 0 9 2 15 1 10 9 13 9 1 0 9 2
17 3 13 14 13 9 15 1 10 2 3 12 9 13 1 0 15 2
25 2 15 6 13 10 1 9 1 9 2 16 6 13 1 15 1 9 2 2 13 0 9 1 9 2
36 9 2 15 3 3 3 13 9 9 1 10 9 7 14 3 13 2 16 2 13 9 1 9 2 2 6 15 4 13 1 9 1 3 0 9 2
16 9 1 11 3 12 9 13 1 0 9 1 9 12 9 3 2
17 3 12 1 12 1 9 13 0 1 9 2 1 15 15 13 9 2
20 13 9 14 15 13 2 16 1 9 1 2 9 2 1 0 9 9 14 13 2
27 1 15 9 3 12 9 13 9 7 9 1 0 1 9 1 0 9 1 9 9 3 6 13 9 1 9 2
26 10 9 15 13 1 0 9 1 9 1 9 1 11 2 16 0 9 1 11 1 9 13 0 10 9 2
34 1 0 9 1 0 9 1 12 9 1 9 3 13 1 9 1 12 9 1 0 0 9 2 15 1 0 9 14 13 1 15 14 13 2
28 3 12 9 13 1 2 11 2 3 9 2 0 1 9 1 0 9 2 13 3 9 9 1 0 9 1 11 2
23 9 2 3 13 1 9 1 0 9 2 15 13 14 15 13 1 9 1 9 1 11 2 2
4 2 13 11 2
30 9 1 0 0 9 11 11 11 4 13 0 9 1 0 0 9 1 9 2 13 9 2 11 11 2 2 0 1 11 2
52 9 1 9 2 0 1 0 9 10 9 1 0 9 1 11 11 11 7 0 9 1 11 2 3 14 13 11 7 0 9 1 11 7 13 14 13 0 9 1 9 1 11 2 15 13 14 13 0 9 1 11 2
8 0 9 3 3 13 0 9 2
29 11 7 9 1 9 1 11 13 3 1 0 1 9 9 1 11 0 9 2 16 11 13 14 13 0 9 1 11 2
28 7 10 0 0 9 1 11 2 15 13 0 9 1 11 2 1 0 9 13 1 9 0 1 15 9 1 9 2
28 15 13 2 16 9 12 2 3 13 0 9 1 11 2 7 15 6 13 2 16 11 6 13 14 13 0 2 2
22 9 1 9 1 11 13 3 1 0 9 9 7 13 1 9 2 16 15 6 13 9 2
32 11 11 2 9 1 0 9 2 11 2 7 0 9 1 0 0 9 2 13 2 16 4 13 9 1 9 1 0 9 11 11 2
18 11 13 0 1 2 9 2 1 9 1 11 13 3 9 2 11 2 2
9 9 1 10 9 13 9 1 11 2
13 12 1 0 13 9 1 0 9 1 11 11 11 2
16 1 9 1 9 15 13 7 13 1 0 9 1 12 0 9 2
10 2 13 1 9 11 9 1 0 9 2
18 9 13 9 1 0 0 9 11 2 15 1 0 9 13 0 15 9 2
9 2 13 11 11 2 9 1 11 2
4 2 13 15 2
28 9 1 0 9 11 11 13 3 2 16 13 12 9 14 13 0 1 9 1 0 9 1 0 9 2 13 11 2
7 2 13 9 1 0 9 2
11 1 9 9 13 7 13 1 0 9 9 2
28 16 0 9 1 9 1 9 11 11 14 13 1 9 1 9 1 12 9 2 0 9 3 3 15 13 1 9 2
