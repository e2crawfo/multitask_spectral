13000 11
6 11 13 15 0 9 2
13 15 13 1 15 9 4 4 4 2 4 7 9 2
7 15 9 13 15 15 4 2
13 15 13 1 10 0 9 15 15 3 3 13 4 2
12 15 13 3 1 15 1 10 9 4 4 4 2
11 15 13 9 9 4 4 7 13 10 15 2
16 16 15 13 0 1 15 9 3 4 4 1 10 9 1 8 2
27 15 9 1 10 9 13 3 9 9 0 2 15 9 1 10 9 2 13 2 13 7 13 1 10 0 9 2
22 15 4 10 9 4 2 15 7 15 9 13 15 3 7 13 4 7 15 9 1 4 2
12 10 9 16 12 9 0 13 4 4 1 9 2
20 15 9 13 15 9 3 16 15 13 4 2 2 15 13 3 0 2 9 2 2
9 15 9 13 3 1 10 9 3 2
11 15 9 4 4 7 4 1 10 0 9 2
21 11 13 10 9 0 4 16 15 3 15 4 16 10 0 9 1 10 9 7 9 2
23 15 13 10 9 1 15 9 2 13 15 12 9 3 7 13 15 1 10 9 1 10 9 2
18 10 9 4 3 15 16 10 0 9 15 15 13 1 10 0 0 9 2
18 10 9 13 0 1 10 9 7 10 9 1 10 9 13 1 10 9 2
10 15 13 10 0 9 4 4 1 11 2
3 13 15 2
12 7 15 13 0 1 15 12 1 10 12 9 4
4 15 13 3 1
7 3 4 0 4 1 10 9
5 3 13 15 1 4
5 3 13 15 1 4
6 1 10 9 4 0 4
7 0 4 4 3 1 10 9
5 1 4 4 3 15
5 15 4 3 1 4
5 3 4 13 3 15
4 15 13 1 4
8 15 13 3 1 10 12 12 9
5 3 13 15 16 1
5 15 4 15 9 2
6 15 13 15 0 4 2
8 15 4 10 9 1 10 9 2
5 15 9 4 12 9
5 10 9 4 12 9
4 13 1 10 9
4 13 1 10 9
7 12 9 13 4 1 10 9
4 13 1 10 9
9 15 13 0 2 0 1 10 9 3
4 13 1 10 9
12 15 13 3 1 4 1 15 9 1 10 0 9
8 15 13 0 4 4 1 10 9
4 15 13 1 9
7 15 13 15 1 10 0 9
8 15 13 15 1 9 1 10 9
4 15 13 12 9
3 15 4 0
4 15 4 12 9
4 15 4 1 11
9 15 13 13 13 16 15 0 0 0
4 15 4 1 12
4 15 4 1 11
4 15 4 12 9
5 15 13 15 1 11
5 15 13 9 1 11
4 15 13 3 4
3 13 3 4
10 15 13 3 3 3 3 3 3 3 4
6 13 3 3 3 0 4
3 15 13 2
6 15 13 3 0 4 2
4 3 9 15 2
6 15 13 15 3 0 2
6 11 3 4 3 4 2
9 15 13 15 3 10 0 9 4 2
9 1 15 9 13 3 10 0 9 2
5 13 15 15 3 2
3 13 15 2
3 9 0 2
10 13 15 1 9 2 13 15 1 11 2
2 13 15
4 15 13 15 2
5 13 15 3 4 2
10 15 13 15 3 16 15 3 4 4 2
9 15 13 16 15 3 3 4 4 2
10 15 0 1 15 3 4 15 3 13 2
9 3 13 15 15 1 2 4 3 2
10 16 15 15 13 2 13 15 15 4 2
11 16 15 15 13 2 13 15 15 15 4 2
11 13 3 10 9 16 15 16 15 3 13 2
11 15 13 3 1 15 16 15 15 13 4 4
11 13 3 10 9 16 15 8 15 3 13 2
8 15 13 15 16 15 15 13 2
11 15 13 3 1 15 8 15 15 13 4 4
8 15 13 15 16 0 3 1 4
8 10 9 16 10 0 9 1 4
7 8 3 15 4 4 7 9
6 8 15 1 10 9 13
7 15 13 3 4 16 15 4
8 15 13 15 3 4 16 15 4
6 15 13 3 10 9 4
4 15 3 15 9
9 13 9 3 16 15 9 3 3 4
4 3 13 15 2
17 16 15 13 4 7 15 13 1 10 9 2 13 15 3 9 4 2
8 10 9 1 11 15 13 3 4
4 9 4 1 4
6 15 4 0 1 9 2
6 15 4 1 9 13 2
7 15 4 0 16 1 4 2
8 15 4 0 16 15 4 4 2
6 15 4 10 9 0 2
5 15 4 15 13 2
12 15 4 15 13 16 3 1 15 1 4 4 2
4 3 13 15 2
6 15 4 0 16 15 13
5 15 4 0 16 15
7 15 4 9 1 9 16 15
5 15 4 10 0 9
5 15 4 10 0 9
5 15 4 10 0 9
5 8 13 1 15 2
6 8 1 9 1 15 12
4 3 0 16 15
5 3 0 16 10 9
4 15 13 15 2
3 3 0 0
4 9 1 10 9
3 10 9 0
4 0 16 1 13
2 8 13
4 0 1 10 9
2 3 3
3 3 3 3
5 3 13 15 9 1
11 15 9 13 15 16 15 15 9 4 4 2
9 16 15 15 13 16 15 15 4 2
5 15 4 3 3 0
6 15 4 3 12 9 0
4 15 4 3 0
5 15 4 12 9 0
5 1 10 9 3 2
4 1 3 1 2
4 1 3 3 2
7 15 13 3 3 3 4 2
10 13 3 3 16 15 15 3 4 4 2
5 15 13 15 4 2
9 13 3 1 15 3 3 1 4 2
7 15 13 16 15 0 4 2
11 15 9 13 15 16 15 15 9 4 4 2
9 1 11 1 10 9 4 15 13 2
11 1 10 9 1 10 9 0 4 15 13 2
8 1 9 1 9 4 15 13 2
6 10 9 1 10 9 2
5 3 1 10 9 2
4 1 15 3 2
5 12 9 3 12 2
10 15 13 15 3 16 15 3 4 4 2
9 8 15 9 4 15 1 10 9 4
9 8 15 9 13 15 15 3 4 4
9 15 13 3 1 9 1 10 9 11
9 10 9 13 1 10 9 1 15 9
2 3 3
3 3 3 3
4 10 0 9 2
4 15 13 15 2
3 0 9 2
3 15 0 2
3 15 0 2
6 10 9 13 10 0 9
7 10 10 9 13 10 0 9
3 0 12 9
3 0 15 9
3 3 15 9
9 13 15 3 1 15 9 1 15 2
8 15 13 3 1 15 0 9 4
5 15 13 15 0 2
9 15 13 3 1 15 0 9 3 4
7 1 15 8 4 8 8 2
6 8 9 13 15 4 2
5 8 9 13 15 2
7 15 13 15 1 9 4 2
9 15 13 15 16 15 8 9 4 2
2 8 2
2 8 2
10 13 3 11 8 0 9 15 4 13 2
4 15 13 15 2
10 13 3 11 8 0 9 15 4 13 2
3 10 0 9
3 8 0 9
6 8 9 4 15 13 2
7 8 9 13 15 9 4 2
8 15 13 15 9 10 9 4 2
7 9 1 10 0 13 10 9
6 15 13 15 1 15 2
9 15 0 13 1 10 9 1 15 9
7 15 0 9 1 10 9 2
5 9 1 10 9 2
10 15 9 16 10 9 3 1 4 4 2
10 10 9 16 15 3 3 3 4 4 2
10 10 9 7 15 9 1 15 4 4 2
4 10 9 1 9
7 10 9 1 9 1 10 9
4 9 1 0 13
5 10 9 16 1 4
7 15 4 15 0 1 10 9
6 10 9 16 0 1 4
5 10 9 0 9 2
4 0 0 11 2
8 10 15 9 15 15 13 4 2
3 0 15 2
3 15 3 2
3 8 15 2
3 8 15 2
9 3 15 15 13 4 1 15 4 2
11 10 1 10 9 9 13 9 13 10 9 2
5 15 13 15 15 2
51 10 9 13 1 10 9 1 10 0 9 1 10 9 3 10 9 4 4 7 13 1 10 0 0 9 7 2 1 13 9 2 1 10 1 10 1 10 9 13 9 7 9 0 9 3 3 10 0 9 3 2
6 10 0 1 13 9 2
6 10 8 1 13 9 2
5 10 9 15 9 2
5 10 9 10 9 2
3 15 0 2
6 15 9 3 3 3 2
6 9 3 1 10 9 2
5 9 1 10 9 2
4 9 1 9 2
7 15 13 15 1 15 4 2
4 10 9 16 3
9 10 9 1 9 1 11 1 11 2
6 10 9 16 1 13 2
20 15 1 13 13 15 15 3 4 2 7 15 13 9 15 8 1 15 3 13 2
8 10 9 16 15 15 3 0 13
3 11 0 2
3 11 0 2
4 15 3 0 2
3 15 13 2
3 15 9 2
9 15 13 3 0 4 15 3 4 2
7 15 13 15 10 9 3 2
3 15 15 2
7 15 16 9 1 10 11 2
7 11 13 10 9 4 1 9
13 15 13 16 15 10 9 4 16 1 10 9 1 13
6 15 15 13 1 9 3
6 15 13 15 1 9 3
7 16 15 15 1 9 13 9
9 16 15 3 1 9 13 1 15 15
10 16 15 15 16 9 1 10 11 0 13
4 10 9 9 2
11 15 13 15 16 15 3 1 10 9 4 2
14 10 9 2 10 0 9 2 13 15 9 1 10 9 2
15 10 0 9 1 10 9 2 9 13 2 4 3 3 4 2
16 15 9 3 2 8 0 3 1 9 2 4 3 1 9 4 2
11 15 13 11 4 2 10 0 9 1 9 2
2 9 12
2 8 2
4 10 9 11 2
4 10 9 11 2
4 10 9 11 2
3 9 11 2
6 15 13 15 3 15 2
3 10 9 2
6 10 9 1 10 9 2
8 15 0 9 9 13 4 4 2
8 15 13 1 9 1 0 9 2
9 9 13 1 9 11 13 15 9 2
5 10 9 1 11 2
6 15 13 1 10 9 2
10 10 9 1 11 1 10 9 1 8 2
4 9 2 11 2
7 9 2 13 15 10 9 2
4 15 4 0 2
12 15 9 2 11 2 15 13 15 3 3 4 2
3 6 11 2
7 15 4 15 0 2 9 2
6 13 3 3 2 0 2
8 7 9 2 15 13 3 15 2
5 13 3 2 6 2
5 9 2 15 11 2
9 9 15 9 2 13 15 10 9 2
7 13 3 3 2 15 9 2
11 15 13 3 1 15 4 2 15 0 9 2
6 15 13 15 10 9 2
6 15 13 9 1 10 9
5 3 13 15 9 3
3 13 15 15
7 13 15 15 15 15 15 4
9 15 13 15 13 3 15 9 1 9
3 3 10 9
4 15 13 3 15
4 15 13 3 15
7 1 10 12 9 13 9 3
8 15 16 9 9 13 15 9 0
6 15 13 15 3 0 2
1 12
2 12 2
1 8
2 8 2
7 10 9 15 15 13 4 2
7 10 9 15 15 13 4 2
11 10 9 1 15 15 0 13 1 4 4 2
8 10 9 3 15 8 3 13 2
7 15 15 13 13 15 4 2
7 15 15 13 4 15 15 2
6 15 13 10 9 0 2
10 3 15 3 0 4 15 13 15 0 2
10 3 10 9 1 15 15 15 3 13 2
8 13 15 1 15 15 4 13 2
9 15 9 15 3 13 13 15 0 2
7 15 13 3 15 15 4 2
10 15 13 3 3 1 15 15 4 13 2
11 15 13 3 3 1 15 15 15 4 13 2
8 15 13 3 3 1 10 9 2
5 15 13 15 3 2
4 15 4 4 2
5 15 13 15 4 2
7 15 13 15 15 4 4 2
7 15 13 15 15 15 4 2
9 15 0 15 15 4 16 15 4 2
9 13 3 0 3 6 13 2 9 2
8 15 13 15 15 9 4 7 3
11 15 13 3 3 15 9 7 3 8 3 4
7 15 13 15 3 0 7 3
5 15 13 15 4 2
11 15 4 3 4 7 15 13 4 4 7 3
6 7 15 15 4 4 2
14 3 15 4 0 3 0 16 15 3 1 11 4 4 2
9 4 15 3 0 3 10 9 7 2
5 11 13 3 1 9
5 3 13 11 1 9
5 3 11 13 1 9
9 15 13 15 16 15 15 3 13 2
10 15 13 15 2 16 15 15 3 13 2
6 16 15 13 13 15 9
7 15 4 3 0 1 4 2
7 16 15 13 3 13 15 9
10 9 2 15 13 15 3 3 3 0 2
8 15 4 3 3 0 0 2 0
7 15 13 15 3 2 3 2
7 15 13 3 0 2 3 2
7 9 2 15 4 0 3 2
8 9 2 4 15 15 9 4 2
6 11 2 15 4 15 0
9 11 2 13 15 10 9 3 0 2
6 15 4 0 3 2 6
8 15 13 9 4 15 15 0 2
6 15 13 15 8 4 2
12 13 3 2 4 15 3 3 8 15 1 4 2
10 13 2 15 13 3 3 3 3 3 2
8 13 2 3 13 15 15 3 3
13 13 15 4 2 15 4 3 3 1 15 3 4 2
12 3 13 15 15 1 2 4 3 2 13 15 2
11 15 4 3 3 3 0 3 2 13 15 2
12 15 4 3 2 13 15 2 3 3 0 3 2
6 13 15 9 2 15 2
4 9 2 13 2
12 1 10 9 2 11 11 2 8 2 10 11 2
5 15 13 15 4 2
5 0 16 3 9 4
8 15 13 3 0 4 15 3 4
7 15 4 0 4 15 13 11
9 15 13 15 9 4 15 15 9 9
18 1 10 0 9 4 8 15 16 15 13 1 9 4 0 13 9 1 4
28 3 4 3 3 3 4 16 9 7 15 1 10 9 1 13 13 3 13 15 15 3 3 4 6 9 4 1 9
22 15 13 15 3 0 1 15 10 9 9 7 9 16 15 3 3 1 15 9 4 4 2
20 15 13 15 3 0 1 15 10 9 9 7 9 3 3 1 15 9 4 4 2
15 15 13 15 3 0 1 15 15 9 16 15 3 4 4 2
16 15 13 16 16 15 0 4 15 3 10 0 9 1 10 9 13
8 15 13 15 16 0 3 1 4
12 15 13 13 1 10 9 4 15 3 3 3 0
19 13 1 10 9 7 3 3 3 10 9 1 9 15 13 15 3 3 3 0
21 15 13 13 1 10 9 7 3 3 3 10 9 1 9 15 13 15 3 3 3 0
18 1 15 9 15 15 1 15 9 16 15 15 13 4 16 15 15 0 13
18 16 15 13 16 15 16 10 9 9 15 15 4 13 16 15 15 3 13
15 15 13 16 15 15 9 13 4 16 15 4 4 16 15 4
8 15 13 15 16 15 9 1 4
8 15 13 15 16 3 0 1 4
5 15 13 1 15 2
6 15 13 1 10 9 2
5 15 13 12 9 2
5 10 9 13 9 2
4 15 13 9 4
17 1 10 9 4 15 0 0 4 2 1 10 9 9 15 13 9 2
4 15 13 3 2
6 15 13 15 1 9 2
5 15 13 1 9 2
5 15 13 15 3 3
5 16 15 15 3 13
5 15 13 15 3 4
7 15 13 15 3 3 1 4
7 16 15 15 3 3 13 4
7 16 15 15 3 13 4 2
7 16 15 15 9 13 4 2
17 7 15 4 0 15 6 3 10 9 1 9 16 15 13 3 15 2
7 16 15 15 0 13 4 2
8 16 15 3 0 9 13 4 2
5 15 13 15 9 2
5 10 9 13 0 2
6 15 13 15 9 3 2
6 10 9 4 8 4 2
7 3 10 0 9 0 8 13
6 16 0 9 8 1 13
5 15 13 0 3 2
6 15 13 15 3 0 2
11 3 13 15 9 1 9 1 15 0 9 2
4 15 13 0 2
7 10 9 4 4 1 10 9
7 10 9 4 1 10 9 4
7 1 10 9 4 10 9 4
10 10 9 13 1 10 9 10 9 4 2
8 10 9 1 10 9 1 10 9
6 15 1 0 13 1 9
7 10 9 1 11 1 10 9
12 15 13 15 10 9 3 3 3 3 3 4 2
12 15 13 15 3 3 3 3 3 10 9 4 2
11 10 9 3 15 10 9 1 0 9 13 2
11 13 10 9 3 3 3 3 3 3 3 2
6 15 4 3 3 0 2
8 15 13 3 9 10 9 1 15
7 13 15 3 0 16 15 13
7 15 13 15 3 16 15 4
9 15 4 3 1 1 9 12 10 9
7 15 13 3 9 3 4 2
14 15 13 16 15 0 4 16 15 15 9 1 9 8 13
8 10 9 1 9 16 15 8 13
8 10 9 15 10 9 1 3 13
11 15 13 15 13 6 15 13 15 3 4 4
5 15 13 16 15 13
6 3 13 15 1 15 2
5 15 13 15 1 9
6 15 13 0 1 15 9
5 10 9 13 15 0
6 3 13 15 15 3 4
6 15 13 15 1 15 13
7 10 9 13 15 1 15 4
8 3 10 9 15 15 15 3 4
4 3 4 15 3
3 10 9 11
4 9 1 9 8
7 11 2 10 9 2 10 9
8 15 9 2 10 9 13 15 4
4 0 7 0 9
3 0 0 9
3 0 0 9
3 0 1 9
6 15 13 15 1 10 9
6 0 16 10 9 4 4
6 3 13 16 15 15 4
6 15 13 16 15 9 4
5 9 10 9 1 11
6 10 9 15 15 9 4
7 10 9 16 15 10 15 4
10 15 13 1 10 9 16 15 0 4 4
5 15 13 15 0 3
5 15 13 4 7 4
4 13 15 15 2
9 15 13 15 1 4 16 15 3 4
4 15 13 15 3
5 15 13 15 1 4
8 15 13 15 4 16 15 4 4
7 9 9 1 9 11 7 11
6 15 13 15 4 16 9
5 15 13 15 4 4
7 15 13 1 4 1 0 9
9 15 13 15 4 4 16 15 4 4
8 11 4 8 10 9 3 1 4
5 15 13 8 1 4
3 13 3 8
4 15 13 15 8
6 15 15 0 4 13 4
10 15 13 15 3 3 16 15 15 4 4
4 9 11 1 11
3 8 15 9
6 15 4 8 1 15 9
4 4 15 8 2
5 11 4 8 1 15
4 11 4 10 0
5 9 4 3 10 0
3 8 10 9
6 3 16 4 15 10 9
1 12
2 12 12
4 9 1 11 11
1 8
1 8
1 8
4 9 1 10 9
4 9 1 10 9
3 0 10 9
5 15 13 3 15 4
5 15 13 3 15 4
4 15 13 3 15
5 15 4 15 3 0
9 10 9 1 10 9 4 15 0 0
6 15 13 3 15 15 4
9 15 13 3 3 1 15 15 4 13
10 15 13 3 3 1 15 15 15 4 13
7 15 13 3 3 1 10 9
4 15 13 15 3
5 10 9 15 15 13
5 15 4 15 15 4
4 15 13 15 2
5 15 9 13 15 2
6 1 15 9 13 15 2
8 15 4 10 9 1 4 1 11
5 15 13 15 15 4
6 15 13 15 9 15 4
6 10 9 3 9 4 4
6 10 9 15 15 13 4
7 16 13 9 3 0 4 2
6 3 13 15 15 4 2
9 10 9 3 15 3 0 3 4 13
10 3 13 10 9 3 10 9 1 9 13
7 15 4 15 3 15 9 13
8 15 13 0 3 0 16 15 4
5 15 13 1 10 9
3 10 9 15
4 15 13 15 15
9 15 13 10 9 3 16 10 0 9
5 1 12 4 15 0
6 15 9 13 9 16 9
6 15 13 8 0 1 9
9 3 1 15 9 13 15 3 1 11
5 15 13 3 1 11
4 15 13 3 3
9 15 13 3 10 9 1 10 9 4
4 10 9 13 0
8 15 13 1 12 4 15 10 9
2 15 9
11 15 4 10 9 9 16 3 1 11 9 13
7 3 13 9 1 10 0 9
3 10 0 9
2 12 9
3 15 0 9
3 15 0 9
3 10 9 9
3 10 9 9
4 15 4 0 3
3 10 9 9
3 10 9 9
4 10 0 9 9
5 12 0 9 0 9
3 10 9 9
3 10 9 9
3 10 9 9
3 0 12 9
3 0 15 9
3 0 10 9
3 3 1 11
7 15 4 3 16 15 9 13
3 1 15 9
3 8 12 9
3 10 9 0
4 15 9 1 9
3 10 9 9
3 15 9 9
4 10 9 1 9
5 10 9 9 4 0
5 10 9 9 4 12
7 3 4 10 9 1 10 9
4 12 1 12 9
4 12 9 12 9
4 12 7 12 9
5 10 0 0 9 9
5 10 0 0 9 9
4 10 9 1 9
3 9 1 9
3 9 1 9
3 9 1 9
5 10 9 1 10 9
4 15 4 8 4
5 10 9 1 10 9
5 10 9 1 10 9
6 10 9 9 13 9 4
6 10 9 9 13 9 4
5 15 13 3 1 9
5 3 13 15 1 9
8 15 13 16 15 3 1 9 4
6 16 15 1 9 13 2
4 13 1 9 2
6 3 13 15 1 9 2
5 15 13 9 1 9
10 15 9 13 16 8 16 15 10 0 4
15 15 13 16 10 9 15 3 4 4 16 15 3 3 1 13
7 15 9 3 3 15 13 4
10 15 13 15 3 3 15 13 3 1 12
7 15 9 3 3 13 15 4
9 15 13 3 1 15 4 15 3 4
7 15 4 0 1 15 1 13
7 15 13 0 16 10 0 9
10 16 9 13 15 0 4 1 10 0 9
9 15 16 11 13 15 3 4 16 9
5 15 13 3 9 4
9 15 13 15 16 4 15 10 0 9
15 0 9 13 3 3 10 9 4 7 4 1 10 0 9 4
9 10 0 15 0 7 15 0 13 9
4 3 0 16 0
6 15 10 9 16 1 15
8 15 13 16 15 3 0 3 4
11 3 13 10 9 16 15 15 9 1 13 4
8 9 2 15 4 15 15 0 13
6 3 3 2 1 15 9
6 16 15 13 13 15 9
4 15 13 10 9
10 16 15 15 13 2 3 13 15 15 3
11 13 8 10 9 2 3 13 15 8 3 4
15 16 15 0 4 7 15 13 1 9 2 3 13 15 4 6
4 3 10 9 3
3 1 3 1
4 1 10 9 3
3 1 3 3
4 1 10 9 1
6 15 4 10 11 1 8
4 1 11 1 11
4 15 13 15 9
4 1 1 1 3
4 1 9 1 9
4 1 8 1 8
10 7 15 4 3 3 0 2 3 2 11
7 3 0 15 13 2 3 0
5 10 9 2 10 9
10 15 4 3 1 15 7 0 3 1 15
5 13 2 15 4 0
8 1 3 10 9 7 3 10 9
3 8 10 9
6 15 13 15 1 9 11
7 15 13 15 0 16 15 0
4 3 15 13 3
5 7 6 15 13 15
6 15 13 0 10 9 4
5 10 9 13 0 4
7 13 15 3 15 10 9 2
6 15 13 15 10 9 3
7 15 13 15 15 1 10 9
9 15 13 3 15 15 1 10 0 9
6 13 15 15 3 4 2
4 15 13 15 0
4 15 13 10 15
4 15 13 10 9
5 13 0 15 10 9
7 10 9 4 10 15 10 9
5 15 13 0 15 15
7 15 13 3 15 15 1 9
9 10 9 1 13 15 13 3 15 9
8 3 13 15 8 15 3 1 9
5 15 13 9 0 9
3 15 13 9
8 15 13 15 0 16 9 1 13
6 15 4 3 0 3 0
9 10 9 3 15 13 16 15 4 4
8 15 13 3 10 0 9 3 4
5 1 15 13 16 0
8 13 9 4 15 8 1 10 11
7 15 13 15 1 9 1 13
7 3 13 3 15 9 1 9
6 1 9 13 15 3 15
10 15 13 15 3 1 10 9 1 9 2
6 15 13 10 9 1 11
4 10 0 9 11
5 15 13 15 1 13
6 15 13 9 1 15 9
4 3 13 13 15
4 9 13 3 9
5 15 9 13 3 3
7 3 4 4 16 15 0 4
3 3 13 15
7 3 13 3 15 1 10 9
5 3 13 15 1 4
5 3 13 15 4 4
4 15 13 3 12
7 10 0 9 4 8 8 4
5 3 4 3 12 0
10 15 4 3 0 3 4 10 9 1 4
10 15 13 3 3 3 3 16 15 3 4
9 15 13 3 3 16 15 3 3 4
4 15 13 3 4
3 15 9 3
5 1 15 4 15 0
5 9 4 0 1 15
5 0 1 10 9 11
5 15 13 10 9 8
6 15 13 15 1 10 9
7 10 9 4 3 1 10 9
5 15 13 1 10 9
5 15 13 12 9 8
3 1 15 3
5 11 15 9 13 3
7 1 15 12 13 15 1 8
5 1 15 15 12 12
4 15 13 1 9
4 15 4 1 9
5 15 9 16 15 8
4 10 0 0 9
3 9 9 12
4 15 13 0 0
7 3 1 10 9 13 15 9
7 15 4 3 3 0 1 15
9 15 13 15 3 4 5 3 3 2
13 13 15 3 3 3 13 9 2 5 6 2 3 3
8 0 9 4 3 3 3 15 4
3 10 9 8
9 13 15 3 2 5 6 2 3 3
8 15 4 3 3 4 4 0 2
8 3 13 15 3 3 1 9 2
4 3 3 15 13
3 3 1 11
5 3 1 10 0 9
3 10 9 3
3 12 9 3
4 3 1 10 9
4 10 9 3 0
3 10 9 8
8 10 11 4 3 0 16 10 11
7 15 13 3 0 1 10 9
6 15 13 0 1 3 3
4 15 13 0 8
7 15 4 15 8 2 13 15
7 15 4 10 9 3 1 9
6 15 4 3 3 3 3
7 10 9 13 3 3 3 1
8 3 10 9 5 15 13 3 2
10 15 13 3 2 10 11 7 10 11 2
3 10 9 11
9 0 13 3 5 10 9 2 13 15
9 2 3 4 15 3 2 13 10 9
6 13 15 0 11 3 2
7 16 15 3 1 10 9 4
6 11 3 13 1 10 9
5 13 9 16 3 11
9 3 2 15 13 15 7 10 9 13
9 13 3 3 1 10 9 1 9 3
6 15 13 3 3 0 4
10 13 15 3 3 3 15 10 9 4 2
2 9 11
8 15 13 9 1 10 9 8 4
8 15 13 1 10 9 8 1 11
4 15 4 3 0
4 15 13 1 11
7 4 15 3 1 11 4 2
8 15 13 15 3 1 10 9 4
8 13 15 15 3 1 10 9 2
4 15 13 1 9
4 15 13 1 9
4 15 13 9 13
2 9 8
5 15 13 15 9 13
4 15 4 15 13
5 9 4 10 9 13
3 3 3 0
3 15 4 0
6 15 4 3 0 16 15
5 15 4 0 16 15
3 15 4 8
4 15 4 10 0
3 0 16 11
4 8 9 1 9
8 15 9 4 10 9 16 10 0
5 15 13 15 16 15
6 10 0 9 16 10 9
4 15 0 16 15
7 15 13 10 9 9 3 3
2 0 15
2 0 15
4 0 9 7 9
6 15 13 8 4 8 4
7 0 13 9 3 0 3 0
7 3 13 10 0 9 9 2
7 15 9 13 9 1 11 2
9 15 9 4 1 10 9 1 11 2
10 1 15 9 13 10 9 2 11 2 2
14 10 9 4 4 1 10 9 1 10 9 2 11 2 2
8 15 9 13 8 10 9 11 2
5 3 4 8 0 2
11 15 0 9 4 9 1 15 13 1 12 2
5 10 9 13 11 2
9 15 4 10 0 9 1 0 9 2
7 15 4 10 9 1 11 2
7 10 0 9 13 1 11 2
8 15 4 10 9 1 15 8 2
5 15 9 13 8 2
8 3 4 10 0 9 0 4 2
10 1 15 9 13 10 9 1 15 8 2
11 3 0 13 15 1 10 0 9 1 13 2
8 11 9 4 10 2 9 2 2
11 15 4 10 9 1 10 9 1 0 9 2
7 1 15 9 4 11 9 2
7 3 13 10 9 11 3 2
7 15 4 10 9 1 11 2
7 1 15 9 13 15 8 2
7 15 4 10 9 1 11 2
5 3 13 15 8 2
7 15 4 10 9 1 11 2
12 15 4 10 0 9 1 9 2 9 7 9 2
6 15 4 10 0 9 2
6 15 13 10 11 4 2
8 15 4 10 9 1 10 11 2
8 10 9 4 4 1 15 8 2
6 15 9 13 11 8 2
8 1 15 4 10 8 9 4 2
8 10 9 4 3 1 10 9 2
8 3 13 10 0 9 1 11 2
11 15 4 10 9 1 10 9 1 10 9 2
9 3 13 10 0 9 1 10 9 2
6 16 4 15 8 4 2
5 10 9 13 8 2
5 10 9 13 11 2
8 11 4 10 9 1 15 9 2
7 15 9 4 9 1 11 2
9 15 4 10 9 1 10 9 11 2
7 1 15 9 4 15 8 2
6 3 13 10 0 9 2
6 16 4 10 11 4 2
7 1 15 0 9 13 8 2
7 1 15 0 9 13 11 2
7 15 4 10 9 1 8 2
11 1 15 4 8 1 10 0 0 9 4 2
9 1 15 9 4 10 11 8 4 2
6 10 9 9 13 3 2
9 10 9 13 3 1 10 0 9 2
6 3 13 10 0 9 2
18 3 13 15 3 13 9 1 8 15 1 8 2 8 8 8 4 4 2
6 15 13 10 11 4 2
6 3 4 15 8 4 2
7 15 4 10 0 0 9 2
7 1 15 9 4 15 8 2
10 15 0 9 13 9 1 10 9 12 2
6 15 4 10 0 9 2
8 1 15 9 4 15 8 4 2
14 3 0 4 10 9 15 1 10 9 1 11 4 4 2
8 10 9 13 9 1 15 8 2
7 3 13 10 9 11 3 2
11 1 15 9 4 10 9 1 10 9 4 2
6 3 4 10 11 4 2
6 3 4 15 8 4 2
9 1 15 9 13 15 2 8 2 2
8 15 9 13 10 9 1 11 2
9 15 9 1 15 8 13 10 9 2
5 15 13 15 8 2
7 3 13 10 9 1 11 2
11 15 0 9 13 9 1 10 9 1 11 2
4 3 4 11 2
12 1 15 9 13 10 9 1 10 11 9 9 2
12 10 9 13 3 9 10 9 1 10 11 9 2
6 3 13 10 0 9 2
6 11 4 15 8 4 2
10 1 15 9 1 11 4 10 9 4 2
13 15 9 13 10 9 3 10 9 1 11 4 4 2
8 15 0 9 13 1 0 9 2
6 3 13 10 9 9 2
10 1 15 9 4 10 9 1 10 11 2
10 10 0 13 3 1 10 9 1 11 2
4 3 13 11 2
10 1 15 9 4 15 2 8 2 4 2
7 3 13 10 9 11 3 2
6 1 15 9 13 8 2
8 15 0 9 13 10 0 9 2
9 15 9 13 9 1 2 8 2 2
15 1 15 9 4 15 2 8 2 1 9 1 10 9 4 2
10 15 4 10 0 9 1 2 9 2 2
8 1 15 9 13 10 9 11 2
10 15 9 13 10 9 1 11 1 12 2
10 1 15 9 4 10 9 3 3 0 2
5 15 9 13 11 2
7 3 13 10 9 1 8 2
6 15 4 10 0 9 2
8 1 15 9 4 15 8 4 2
5 10 9 13 11 2
5 3 4 8 4 2
7 15 4 10 9 1 11 2
15 15 9 13 10 9 2 8 2 1 9 8 1 15 8 2
9 1 15 9 13 10 0 9 11 2
13 15 9 13 11 16 10 9 13 1 11 1 12 2
17 10 9 13 10 9 16 1 4 1 15 0 8 2 1 10 11 2
9 15 4 10 0 0 9 1 11 2
6 1 15 9 13 8 2
6 15 4 9 1 11 2
5 10 9 13 11 2
14 3 3 4 10 0 9 8 9 9 1 15 8 4 2
9 3 4 10 9 7 9 1 11 2
8 15 4 10 9 1 15 8 2
10 1 15 9 4 10 9 1 15 8 2
10 3 3 4 15 1 11 1 9 4 2
7 1 15 9 4 15 8 2
10 1 15 9 0 11 1 10 9 9 2
9 10 0 9 13 9 1 10 11 2
7 3 13 10 9 11 3 2
7 15 4 10 9 1 11 2
6 15 13 10 11 9 2
13 3 4 10 9 11 1 10 9 16 10 9 4 2
11 1 15 9 1 10 9 4 15 8 4 2
4 15 13 11 2
6 15 9 13 11 8 2
8 1 15 9 9 4 9 4 2
7 15 9 13 10 11 9 2
9 15 9 13 15 9 3 1 11 2
5 15 13 15 8 2
9 15 4 10 0 9 1 10 11 2
6 3 13 10 0 9 2
10 15 0 9 13 10 11 1 11 3 2
14 1 15 9 13 10 0 9 1 9 1 10 11 9 2
9 15 12 0 9 4 8 1 11 2
10 1 15 9 13 10 9 2 8 2 2
12 3 13 10 9 1 10 9 2 8 2 9 2
10 1 15 9 13 10 9 2 8 2 2
14 10 9 4 4 1 10 9 1 10 9 2 8 2 2
14 15 4 10 0 9 1 10 9 1 15 2 8 2 2
14 15 13 10 9 1 10 9 1 10 9 2 8 2 2
18 15 4 10 9 1 9 1 10 9 1 10 9 1 15 2 8 2 2
6 10 0 9 13 11 2
8 15 4 10 9 1 15 8 2
8 10 9 4 9 1 15 8 2
11 1 15 9 4 10 9 1 10 9 4 2
10 3 13 10 0 9 1 15 8 9 2
11 1 15 9 13 10 9 1 10 11 9 2
11 1 15 9 13 10 9 1 15 8 9 2
6 10 9 13 10 11 2
7 15 4 10 9 1 11 2
11 1 15 9 4 10 11 7 10 11 4 2
6 15 4 10 0 9 2
5 10 9 13 11 2
8 15 4 10 9 1 10 11 2
11 15 9 13 11 11 10 0 9 1 9 2
7 15 9 4 1 8 4 2
14 15 0 9 4 4 1 9 1 15 13 1 10 9 2
11 15 0 9 4 1 10 9 4 1 9 2
14 1 15 9 13 8 2 10 0 9 1 9 2 3 2
15 1 15 9 13 10 0 9 10 9 1 9 1 9 3 2
10 1 15 9 4 10 9 1 9 4 2
14 1 15 9 4 1 8 10 9 4 8 9 1 9 2
16 1 15 9 13 10 9 1 11 2 8 2 1 10 0 9 2
6 10 9 13 15 8 2
9 1 15 0 9 13 10 9 9 2
13 10 0 13 8 1 9 1 10 9 2 11 2 2
8 3 13 10 9 1 11 9 2
9 1 10 9 4 10 0 11 4 2
10 10 9 13 4 16 10 9 1 11 2
8 15 9 1 10 9 13 9 2
6 3 0 4 15 8 2
5 3 13 11 3 2
10 10 9 13 10 2 8 2 9 3 2
8 15 4 10 9 1 15 8 2
10 3 13 15 8 10 9 3 1 11 2
6 16 4 10 9 4 2
9 15 0 9 13 9 3 11 11 2
16 10 9 13 16 1 15 13 1 10 11 1 10 9 1 11 2
6 10 9 13 10 9 2
6 16 4 15 8 4 2
7 15 9 4 4 1 8 2
8 3 13 15 8 1 12 9 2
7 1 15 9 4 8 0 2
7 1 15 9 4 15 8 2
16 15 4 4 1 2 8 2 2 10 9 1 10 0 9 8 2
5 10 9 13 11 2
8 1 15 9 4 2 11 2 2
13 15 4 10 0 9 1 10 0 9 2 11 2 2
7 15 4 10 9 1 11 2
5 10 9 13 11 2
7 15 9 13 10 0 9 2
6 1 15 9 13 11 2
9 15 4 10 9 1 2 8 2 2
7 3 4 10 0 9 4 2
10 15 4 9 1 15 8 1 15 8 2
7 3 13 10 0 9 3 2
8 3 0 13 10 9 1 9 2
8 15 9 13 10 9 1 11 2
7 1 15 9 13 10 9 2
10 3 1 11 4 3 10 9 1 9 2
7 1 15 9 4 9 4 2
8 10 9 13 10 9 9 4 2
8 15 4 10 9 1 10 9 2
6 16 4 15 8 4 2
8 15 4 10 9 9 1 9 2
9 3 0 4 10 0 9 1 11 2
7 15 4 10 9 1 11 2
10 15 4 10 9 1 15 2 8 2 2
11 15 0 9 4 3 1 10 0 11 4 2
13 3 13 10 0 9 8 10 9 1 10 0 9 2
14 15 11 9 13 10 9 1 15 9 1 10 0 9 2
10 1 15 9 13 10 9 2 11 2 2
10 10 9 13 15 0 1 9 1 11 2
5 15 4 11 9 2
8 1 15 9 13 8 10 9 2
10 15 13 10 9 1 15 8 0 4 2
7 10 9 4 4 1 9 2
8 15 13 10 9 3 1 11 2
8 15 4 10 9 0 1 9 2
7 3 13 10 9 11 3 2
7 15 4 10 9 1 8 2
5 10 9 13 8 2
6 3 13 10 8 9 2
11 13 10 0 9 15 1 10 9 4 4 2
5 16 4 8 0 2
4 3 13 11 2
7 15 4 15 2 8 2 2
11 10 9 13 16 10 9 11 13 7 13 2
5 3 13 11 3 2
7 10 9 4 3 1 11 2
8 10 9 4 0 4 1 11 2
5 3 0 4 8 2
6 15 4 12 9 0 2
9 15 4 10 9 1 10 11 11 2
7 1 15 9 4 8 9 2
9 13 10 9 3 8 10 9 13 2
8 3 13 10 9 1 10 11 2
5 10 9 13 11 2
8 15 9 4 9 1 15 8 2
8 15 4 10 9 1 10 11 2
8 3 4 10 9 4 1 11 2
6 13 10 9 1 9 2
6 3 13 10 0 11 2
5 3 13 8 8 2
8 15 4 10 0 9 1 11 2
9 15 4 10 0 9 1 10 9 2
7 15 4 10 9 1 8 2
5 13 10 13 9 2
14 3 3 1 15 9 13 10 9 10 9 1 11 4 2
5 3 4 11 4 2
14 10 9 13 10 9 4 16 1 15 8 9 4 4 2
9 3 13 10 9 1 10 9 8 2
8 15 4 10 0 9 1 8 2
7 3 13 11 10 0 9 2
8 15 0 9 13 11 1 12 2
6 13 10 9 1 9 2
8 15 4 10 9 1 15 8 2
7 15 13 10 0 9 8 2
10 15 0 9 13 12 9 4 1 11 2
7 3 13 10 0 0 9 2
8 15 4 10 9 1 15 8 2
6 1 15 9 13 8 2
7 15 4 10 9 1 11 2
10 15 4 3 10 11 1 10 9 4 2
8 15 9 13 1 12 10 9 2
10 3 13 10 9 1 10 9 11 8 2
9 3 0 4 10 9 1 15 8 2
6 3 0 4 15 8 2
7 16 13 10 0 1 11 2
8 3 13 10 9 1 10 11 2
4 3 13 8 2
9 3 13 15 0 8 2 11 2 2
15 15 9 1 10 9 1 9 4 4 1 10 9 1 11 2
11 3 0 4 8 1 10 9 4 1 11 2
6 3 0 4 10 11 2
7 10 9 13 10 9 11 2
14 1 15 9 1 11 13 10 9 1 10 9 0 9 2
9 1 10 0 4 15 8 0 4 2
13 13 10 9 15 1 15 8 2 11 2 4 4 2
8 15 9 13 10 9 11 4 2
11 13 10 9 7 9 3 10 11 4 4 2
13 1 15 9 4 15 13 1 0 7 0 9 4 2
10 15 9 4 3 15 2 8 2 4 2
7 13 10 9 1 15 8 2
7 3 13 10 9 1 8 2
4 3 13 11 2
5 3 13 11 3 2
7 3 13 8 15 0 9 2
11 3 4 13 1 10 9 11 1 9 4 2
5 10 9 13 11 2
9 15 9 13 10 9 2 8 2 2
5 3 13 8 8 2
8 15 4 10 0 9 1 9 2
4 3 13 8 2
5 10 9 13 8 2
7 15 4 10 9 1 11 2
16 15 4 10 9 1 10 9 1 10 9 1 10 0 9 11 2
8 15 4 10 9 1 8 9 2
7 1 15 9 4 13 4 2
5 16 4 11 0 2
11 1 15 8 11 15 11 4 10 9 4 2
7 15 9 13 8 11 11 2
11 15 0 0 0 13 1 10 0 9 11 2
10 15 4 10 0 9 1 10 0 9 2
7 15 4 10 9 1 11 2
10 10 9 13 8 0 9 1 10 9 2
8 10 0 13 4 3 1 11 2
7 15 13 10 2 9 2 2
7 15 13 10 9 1 11 2
7 15 4 10 9 1 11 2
9 15 4 10 9 1 2 8 2 2
10 15 9 4 3 3 2 8 2 4 2
6 3 13 15 10 11 2
12 15 4 10 9 1 10 9 1 10 9 8 2
12 3 0 4 10 9 1 10 9 1 0 9 2
6 13 10 9 1 8 2
12 10 0 9 13 3 1 10 0 9 1 11 2
9 15 4 3 1 10 9 1 11 2
4 15 13 9 2
9 1 15 9 4 10 9 1 11 2
6 15 4 10 0 9 2
7 3 4 10 9 1 11 2
10 15 4 3 10 0 9 1 9 4 2
8 1 15 0 9 13 15 8 2
12 1 15 9 13 10 0 0 9 8 9 0 2
5 15 4 10 9 2
5 16 4 8 0 2
8 15 4 10 0 9 1 8 2
6 1 15 9 13 11 2
5 10 9 13 11 2
10 3 4 10 9 4 1 10 11 8 2
8 15 4 10 0 9 1 11 2
8 16 4 10 0 9 1 11 2
6 1 15 9 13 8 2
6 10 13 9 13 11 2
5 3 4 8 0 2
6 3 13 10 9 11 2
4 3 13 8 2
13 15 9 1 0 9 13 0 1 15 0 0 9 2
5 3 13 8 3 2
8 1 15 9 13 15 8 8 2
10 15 4 10 9 1 10 0 9 11 2
7 15 4 10 9 1 8 2
6 13 10 9 1 11 2
9 15 4 10 9 1 15 0 8 2
6 3 13 11 11 4 2
6 15 13 2 8 2 2
5 3 0 4 8 2
6 3 0 4 15 8 2
11 15 9 13 16 0 9 1 15 8 3 2
11 1 15 9 13 10 0 9 8 9 4 2
17 1 15 9 13 11 1 10 9 16 3 3 1 4 1 15 8 2
6 3 13 8 15 9 2
5 10 9 13 11 2
11 15 4 10 1 12 1 0 9 1 11 2
8 15 4 10 0 9 1 9 2
4 3 13 8 2
8 3 4 10 9 4 1 11 2
7 15 9 13 10 9 8 2
8 15 4 10 0 9 1 8 2
10 15 0 9 13 10 9 1 9 3 2
9 13 10 9 15 1 11 4 4 2
7 15 4 10 9 1 11 2
4 3 13 8 2
7 10 13 1 9 13 11 2
8 3 13 15 8 1 11 9 2
7 15 9 13 15 1 11 2
9 3 3 4 11 9 1 11 4 2
9 15 4 10 0 9 1 9 11 2
8 10 9 13 11 1 12 4 2
4 15 4 9 2
11 3 0 13 15 8 2 10 3 0 9 2
16 1 15 15 9 13 8 1 8 15 8 1 10 9 1 11 2
11 1 15 9 1 11 4 10 0 9 4 2
6 15 9 13 10 11 2
12 3 13 10 9 15 10 9 1 10 9 13 2
10 15 4 8 1 11 1 12 1 12 2
7 15 0 0 13 15 8 2
8 3 13 10 0 0 0 9 2
13 15 9 4 1 12 1 10 9 1 10 9 4 2
14 1 15 9 13 8 2 10 9 0 9 2 9 0 2
10 15 4 10 0 9 1 10 0 9 2
5 10 9 13 11 2
12 3 0 4 8 2 10 0 9 1 10 9 2
12 15 4 10 9 1 10 9 11 1 10 11 2
7 15 4 9 1 10 11 2
7 16 4 10 9 11 4 2
8 15 4 10 9 1 15 8 2
8 3 0 4 8 16 15 13 2
11 15 4 10 9 1 10 9 7 10 9 2
7 15 4 10 9 1 9 2
6 3 0 4 10 9 2
8 10 9 13 9 1 15 8 2
8 1 15 9 4 15 8 4 2
10 1 15 9 13 11 3 1 15 8 2
8 15 4 10 9 1 15 8 2
6 15 4 10 0 9 2
7 15 4 10 9 1 11 2
6 16 4 10 11 4 2
5 3 13 11 3 2
9 15 4 10 0 9 1 0 9 2
6 15 13 10 9 11 2
6 3 0 4 15 8 2
7 3 13 11 1 10 9 2
6 15 4 10 0 9 2
7 15 4 10 9 1 11 2
7 15 9 4 0 9 9 2
13 15 4 10 9 1 10 9 1 10 0 9 9 2
7 15 4 10 9 1 11 2
6 10 9 13 15 8 2
5 10 9 13 11 2
5 10 9 13 11 2
7 3 13 10 9 9 3 2
5 10 9 13 11 2
5 3 4 13 4 2
9 3 13 10 9 1 10 9 9 2
5 3 4 13 4 2
6 10 9 13 10 9 2
7 3 4 10 10 9 4 2
9 15 9 4 10 0 9 1 9 2
10 10 9 4 3 1 9 1 9 4 2
9 15 9 13 10 0 9 1 11 2
6 3 4 15 8 4 2
6 15 13 15 8 4 2
6 3 13 10 0 9 2
7 15 4 10 9 1 11 2
7 1 15 0 9 13 8 2
9 1 15 0 9 13 15 10 9 2
5 10 9 13 8 2
7 15 13 10 9 1 9 2
4 3 13 11 2
7 15 4 10 9 1 11 2
6 3 13 10 0 9 2
4 3 13 11 2
7 15 4 10 9 1 11 2
6 16 13 10 0 9 2
8 15 13 10 9 1 15 8 2
11 3 13 10 11 9 1 10 9 1 12 2
10 15 9 13 11 2 11 7 11 4 2
11 15 9 4 10 0 9 1 9 1 11 2
7 15 13 10 9 9 3 2
10 3 0 4 10 9 1 11 1 9 2
11 1 15 9 13 10 9 1 10 11 9 2
11 10 9 4 3 1 10 9 1 10 11 2
7 1 15 9 13 10 11 2
4 3 13 11 2
7 10 9 13 1 15 8 2
10 15 4 10 9 1 15 8 1 12 2
4 3 13 8 2
7 3 13 2 11 2 3 2
7 15 8 8 9 1 11 2
6 15 9 13 8 4 2
11 15 9 8 1 10 9 1 10 8 11 2
7 10 9 13 10 9 8 2
8 15 13 10 11 1 11 4 2
5 3 4 8 0 2
5 3 4 8 0 2
9 3 13 10 0 0 9 1 11 2
6 15 4 10 0 9 2
8 11 4 10 9 1 15 9 2
9 15 4 10 9 1 11 1 12 2
7 15 4 10 9 1 11 2
5 10 9 13 11 2
10 3 13 10 0 9 1 15 8 9 2
7 1 15 9 4 8 9 2
8 15 9 13 15 12 1 12 2
9 16 4 10 0 9 1 10 11 2
12 15 9 13 1 8 1 10 9 1 10 11 2
4 3 13 11 2
6 3 13 15 8 9 2
6 10 9 13 1 11 2
12 15 4 10 0 9 1 8 2 9 1 11 2
10 10 9 4 3 4 1 10 8 9 2
13 15 9 13 10 0 9 1 15 8 1 15 8 2
9 15 4 10 9 1 2 8 2 2
12 15 13 10 9 1 10 0 9 1 15 8 2
7 3 13 10 9 1 11 2
8 1 15 9 13 10 9 8 2
8 15 4 10 0 9 1 11 2
5 16 4 8 4 2
8 15 0 9 13 8 1 11 2
8 10 9 13 8 4 1 12 2
13 3 13 10 9 1 8 15 0 1 11 4 4 2
8 10 9 13 1 10 11 9 2
6 3 13 8 7 8 2
7 15 4 10 9 1 8 2
11 15 9 1 10 0 9 4 9 12 0 2
8 15 4 10 0 9 1 9 2
7 1 15 9 4 8 9 2
9 3 13 10 0 9 9 1 12 2
8 15 4 10 0 9 1 11 2
6 1 15 9 13 8 2
4 3 13 8 2
4 3 13 11 2
10 1 16 4 3 10 9 1 11 8 2
7 15 4 10 9 1 8 2
5 3 4 15 8 2
4 3 13 11 2
5 3 13 15 8 2
4 3 13 8 2
5 3 4 8 0 2
8 15 4 10 0 9 1 11 2
4 3 13 11 2
8 15 4 10 0 9 1 11 2
6 1 15 9 13 8 2
4 3 13 8 2
6 1 15 9 13 8 2
5 3 4 8 0 2
6 3 13 10 8 9 2
9 15 4 10 0 9 1 15 8 2
4 3 13 11 2
7 15 4 3 0 0 9 2
7 15 4 10 9 1 11 2
7 3 13 10 11 9 3 2
10 1 15 9 13 10 11 1 10 11 2
7 1 15 0 9 13 8 2
4 3 13 11 2
4 3 13 11 2
8 15 4 10 9 1 10 9 2
6 15 13 2 8 2 2
6 15 13 10 9 13 2
7 15 4 15 2 8 2 2
8 15 4 10 9 1 15 8 2
5 11 9 4 8 2
7 15 4 10 9 1 11 2
7 15 4 10 9 1 11 2
8 15 4 10 0 9 1 11 2
6 1 15 4 8 4 2
9 15 4 10 0 9 1 15 8 2
6 15 4 9 1 11 2
8 15 4 10 0 9 1 11 2
7 15 4 10 9 1 8 2
7 15 4 10 9 1 8 2
10 15 4 10 9 1 10 9 1 11 2
8 15 13 10 9 2 8 2 2
9 15 4 10 0 9 1 10 9 2
7 3 13 10 9 1 11 2
7 15 4 10 9 1 11 2
5 15 9 13 8 2
8 1 15 9 4 8 10 9 2
8 15 9 13 15 8 1 9 2
7 1 15 9 4 8 9 2
8 15 9 13 10 9 1 8 2
6 1 15 9 13 8 2
11 15 13 10 11 2 9 1 0 9 2 2
7 10 9 13 10 0 9 2
7 10 9 4 3 1 11 2
5 3 4 15 8 2
5 3 0 4 8 2
8 0 4 15 1 11 1 11 2
6 3 0 4 10 11 2
7 15 13 10 9 1 11 2
7 15 4 10 9 1 11 2
6 10 9 13 15 8 2
9 10 9 13 11 4 1 15 9 2
8 15 4 10 9 1 10 9 2
6 3 4 10 11 4 2
5 16 4 11 0 2
9 3 13 10 9 2 8 2 3 2
5 16 4 8 4 2
4 3 13 8 2
4 3 13 8 2
9 1 15 9 4 11 1 11 4 2
8 3 4 2 8 2 10 9 2
10 1 15 9 13 10 2 0 11 2 2
6 3 4 10 11 4 2
11 15 4 10 9 1 10 9 1 15 8 2
6 15 4 1 12 4 2
5 3 4 8 0 2
6 15 9 4 9 9 2
4 3 13 11 2
10 3 4 11 1 10 0 9 9 9 2
7 15 4 10 0 0 9 2
7 15 13 11 1 10 9 2
8 15 9 4 10 9 1 11 2
6 1 15 9 13 8 2
5 15 9 13 8 2
5 15 9 13 8 2
6 15 4 8 1 8 2
11 1 15 9 4 10 9 1 10 11 4 2
6 15 0 9 13 8 2
5 15 9 13 9 2
6 15 4 10 0 9 2
9 15 4 10 9 1 10 9 9 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
3 15 4 8
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
7 15 4 15 2 8 2 2
5 15 4 10 11 2
5 15 4 10 11 2
4 15 4 11 2
6 3 13 10 9 9 2
10 1 15 9 4 10 9 4 1 8 2
7 15 4 10 9 1 11 2
8 1 15 9 4 10 8 9 2
7 15 4 10 9 1 9 2
8 1 15 13 10 9 15 9 2
8 15 4 10 9 1 9 11 2
12 10 9 4 3 4 1 10 9 1 9 11 2
4 15 4 8 2
5 15 9 13 8 2
9 3 13 8 10 9 1 10 9 2
9 15 4 10 0 9 1 10 9 2
8 10 0 9 4 3 1 11 2
7 1 15 9 13 10 9 2
6 3 4 0 9 4 2
9 15 9 4 10 0 9 1 0 2
8 1 15 9 13 10 9 11 2
6 1 15 9 13 11 2
7 15 9 13 15 1 11 2
10 10 12 9 13 3 16 1 15 8 2
6 3 4 10 9 11 2
12 3 13 10 0 9 1 0 9 1 10 9 2
7 1 15 9 13 15 8 2
5 15 4 11 9 2
6 15 4 10 0 9 2
6 15 13 2 8 2 2
7 15 4 10 9 1 11 2
8 15 9 13 10 2 11 2 2
16 3 13 10 9 1 8 1 1 10 9 8 2 8 7 8 2
9 15 9 13 1 10 9 1 11 2
9 15 4 10 0 9 1 15 8 2
5 15 9 13 8 2
12 15 13 8 1 10 0 9 1 10 12 9 2
14 15 13 8 1 10 0 9 1 10 9 1 15 12 2
6 3 13 10 11 9 2
7 15 13 15 16 10 9 2
13 1 15 9 13 11 2 10 0 9 1 9 11 2
10 1 15 9 13 8 16 15 0 4 2
4 3 13 8 2
7 15 4 10 9 1 8 2
6 1 15 4 8 4 2
13 1 15 9 13 8 1 4 1 15 2 8 2 2
7 1 15 9 13 8 3 2
5 3 13 8 9 2
8 15 4 10 9 1 10 9 2
12 10 9 13 10 11 3 1 9 1 10 9 2
5 15 4 10 9 2
5 15 4 10 11 2
13 15 9 13 8 1 10 9 1 15 2 8 2 2
8 10 9 4 4 1 15 8 2
7 15 4 10 0 0 9 2
9 10 9 13 1 9 1 15 8 2
8 13 10 9 1 10 0 9 2
7 1 15 9 4 11 4 2
6 3 13 10 9 9 2
18 15 9 13 10 12 9 15 10 9 13 1 10 9 1 8 1 12 2
4 3 13 11 2
7 3 4 10 0 9 4 2
7 10 0 4 3 1 11 2
7 3 4 10 9 1 8 2
7 15 4 10 9 1 11 2
6 15 13 9 13 13 2
5 3 4 11 13 2
5 15 13 10 9 2
5 15 13 9 4 2
10 1 15 9 4 10 2 9 2 4 2
6 3 0 4 10 9 2
6 10 0 9 13 3 2
8 10 9 4 3 1 10 9 2
8 10 9 4 3 1 10 9 2
7 1 15 9 4 15 8 2
9 1 10 0 9 4 10 9 4 2
11 10 9 4 3 1 12 1 15 8 4 2
10 1 15 9 4 10 9 4 1 11 2
7 10 9 13 1 10 11 2
9 10 9 13 8 1 10 9 4 2
10 3 4 10 0 9 15 1 9 13 2
9 10 13 13 1 11 1 10 9 2
4 15 4 11 2
9 1 15 9 15 9 0 1 11 2
6 3 4 15 8 4 2
8 13 15 15 1 9 4 4 2
11 1 15 9 4 0 4 1 10 0 9 2
8 10 9 4 3 1 10 9 2
8 15 4 10 0 9 1 11 2
7 3 13 15 1 10 9 2
10 15 9 4 4 1 10 9 1 9 2
11 15 0 9 13 15 3 1 10 0 9 2
4 15 13 9 2
5 3 4 11 4 2
7 10 9 13 11 3 9 2
9 13 4 10 0 9 1 11 4 2
6 10 9 4 3 4 2
8 10 9 4 3 1 10 9 2
7 15 4 10 9 1 8 2
9 15 9 13 10 13 9 1 9 2
10 13 10 9 15 4 4 1 15 8 2
7 3 13 10 9 8 3 2
7 13 10 9 1 10 11 2
5 15 4 15 8 2
6 3 4 15 11 4 2
4 13 10 9 2
8 1 15 9 13 10 0 9 2
4 15 4 8 2
5 3 13 8 3 2
5 3 13 11 3 2
9 1 15 4 10 9 1 11 4 2
4 13 10 0 2
7 1 15 4 10 11 4 2
6 10 0 9 13 3 2
5 15 4 10 11 2
7 15 4 10 9 1 11 2
8 10 9 13 3 11 1 11 2
5 16 4 11 0 2
6 3 4 10 8 9 2
7 13 10 9 16 9 13 2
4 3 13 9 2
6 15 13 2 11 2 2
5 3 4 15 8 2
7 3 4 10 0 0 9 2
7 16 13 9 11 7 11 2
4 3 4 9 2
5 15 13 10 11 2
5 3 4 15 8 2
9 1 15 9 13 10 9 11 3 2
5 15 4 10 11 2
7 15 4 10 9 1 9 2
7 1 15 0 9 13 11 2
10 1 15 9 13 15 8 9 1 11 2
5 3 4 9 4 2
9 15 4 10 9 1 2 11 2 2
4 15 4 8 2
8 3 13 11 15 3 1 11 2
5 13 10 0 9 2
9 3 13 10 9 1 15 8 8 2
5 3 4 8 4 2
4 15 13 9 2
4 3 13 8 2
10 1 15 9 4 10 9 1 11 0 2
7 1 15 9 13 15 8 2
5 3 4 9 4 2
5 3 13 15 8 2
9 3 13 10 9 1 10 11 4 2
4 15 4 8 2
5 15 4 10 9 2
4 3 13 8 2
9 15 13 10 9 1 2 8 2 2
5 15 4 10 9 2
7 3 13 10 9 4 4 2
5 15 9 13 9 2
7 15 4 10 9 1 8 2
5 15 4 10 11 2
8 3 13 9 9 16 1 9 2
5 3 4 15 8 2
11 10 9 13 10 9 1 10 9 1 4 2
7 15 4 10 9 1 11 2
4 3 13 11 2
5 15 9 13 8 2
7 1 15 9 13 10 9 2
8 1 15 9 4 10 11 4 2
6 3 4 0 9 4 2
5 15 13 10 11 2
6 10 9 13 1 11 2
6 8 9 9 13 11 2
5 10 9 13 3 2
7 3 13 10 9 1 8 2
4 13 10 9 2
7 1 15 9 4 15 8 2
9 10 9 4 3 0 1 9 4 2
9 15 4 10 0 0 9 1 11 2
6 15 9 13 1 11 2
7 10 9 1 11 15 9 2
4 15 4 8 2
4 15 4 8 2
6 15 13 2 8 2 2
7 15 13 10 9 11 4 2
5 15 13 10 9 2
8 13 10 9 1 9 1 9 2
9 3 4 11 2 10 9 2 4 2
5 15 4 10 11 2
4 15 4 0 2
5 3 4 8 4 2
5 3 4 15 8 2
14 15 9 13 3 1 10 9 1 10 9 2 8 2 2
9 13 10 0 9 15 8 4 4 2
8 1 15 9 4 9 8 9 2
8 15 13 10 9 11 1 11 2
4 15 4 8 2
5 3 0 4 8 2
4 15 4 11 2
7 1 15 9 13 15 8 2
7 15 4 10 0 0 9 2
7 13 10 9 1 10 9 2
6 3 13 15 9 4 2
4 15 9 13 2
10 10 9 9 3 1 11 1 10 9 2
9 15 13 10 9 1 2 8 2 2
4 3 13 3 2
5 3 4 8 4 2
9 1 15 4 10 9 2 8 2 2
7 1 15 9 13 10 11 2
6 15 9 13 15 8 2
7 15 4 10 9 1 8 2
9 13 10 9 3 10 9 4 4 2
7 13 10 9 15 13 13 2
9 15 9 4 10 0 9 1 9 2
5 15 9 13 8 2
8 3 13 15 2 8 2 9 2
7 15 13 15 2 8 2 2
13 1 15 9 13 11 3 1 10 9 1 12 9 2
9 15 9 13 8 2 8 7 8 2
12 15 9 1 10 9 1 9 4 4 1 11 2
14 10 9 13 3 1 11 7 11 1 10 9 1 12 2
8 10 9 4 13 9 1 11 2
8 15 9 13 10 11 9 3 2
6 3 0 4 10 11 2
15 3 0 13 11 3 1 10 0 9 1 11 3 1 4 2
13 10 9 4 3 4 1 10 9 1 10 9 11 2
11 10 9 4 3 1 9 1 10 0 11 2
12 10 9 13 3 1 9 1 10 9 1 11 2
10 10 9 13 10 9 1 11 7 11 2
8 3 13 10 9 1 10 9 2
11 15 9 13 10 9 1 15 2 8 2 2
7 13 10 0 7 0 9 2
10 15 13 15 4 1 15 2 8 2 2
5 3 4 10 11 2
14 15 9 13 10 16 12 0 7 13 8 1 10 9 2
13 1 15 13 1 15 9 4 10 9 1 8 4 2
5 15 13 8 4 2
10 15 9 4 1 8 1 8 8 4 2
12 15 0 8 13 8 10 0 9 3 1 9 2
6 1 15 9 13 11 2
6 3 4 10 9 4 2
8 3 13 15 8 9 1 12 2
7 1 15 9 4 15 13 2
7 1 15 9 4 10 9 2
5 3 13 9 11 2
4 3 13 8 2
4 3 13 11 2
7 1 15 9 13 10 9 2
8 15 0 9 13 10 11 4 2
7 15 4 9 1 15 8 2
9 15 13 10 0 9 2 8 2 2
11 15 4 10 9 1 10 0 9 1 11 2
6 15 13 2 8 2 2
23 15 13 15 8 11 11 7 0 9 1 15 9 1 10 9 1 10 0 0 9 1 9 2
11 15 13 10 2 8 2 9 8 1 4 2
7 15 13 15 0 8 3 2
10 15 13 10 9 1 15 8 1 11 2
10 15 13 10 0 11 11 2 8 2 2
10 3 13 10 0 0 9 1 10 9 2
10 1 15 9 4 10 0 9 1 11 2
5 16 4 8 4 2
12 1 15 9 4 10 9 1 10 9 1 11 2
6 3 13 10 0 9 2
5 16 4 10 9 2
9 1 15 9 1 8 13 10 9 2
8 16 4 10 0 9 1 11 2
6 3 13 10 11 8 2
6 3 13 8 1 11 2
4 13 10 9 2
4 13 10 9 2
7 1 15 9 4 8 13 2
11 1 15 0 9 13 10 11 0 9 4 2
5 15 9 13 11 2
7 15 9 4 1 8 4 2
10 15 9 13 10 0 0 9 1 11 2
11 15 0 9 13 8 0 9 7 9 4 2
12 15 9 13 0 9 0 1 10 9 1 9 2
19 15 9 4 1 11 2 11 2 11 2 11 2 8 2 11 7 11 4 2
5 15 4 10 11 2
7 15 4 10 2 11 2 2
4 15 4 8 2
4 15 4 8 2
4 15 4 11 2
4 15 4 8 2
4 15 4 8 2
5 15 4 10 11 2
4 15 4 8 2
5 15 4 15 8 2
9 15 4 9 1 15 8 1 12 2
12 1 15 9 4 9 1 15 8 4 1 12 2
8 15 4 9 1 11 1 12 2
8 15 4 9 1 11 1 12 2
7 15 9 13 3 1 12 2
12 1 15 9 2 1 12 2 13 10 9 9 2
9 15 13 10 9 1 11 1 12 2
9 15 9 13 10 0 9 1 12 2
12 15 0 9 13 12 2 8 2 9 1 12 2
18 15 4 10 13 11 9 1 10 9 12 1 15 13 1 10 0 9 2
10 15 4 10 0 9 16 9 1 4 2
10 3 13 10 9 0 1 9 15 4 2
9 3 13 15 8 1 9 4 4 2
10 3 13 15 1 9 4 4 1 11 2
10 3 13 2 1 10 0 9 2 9 2
5 3 4 8 4 2
8 3 13 15 2 8 2 4 2
9 3 13 9 1 10 9 4 4 2
7 3 4 10 0 9 4 2
5 3 9 15 13 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 3 13 11 2
4 15 4 8 2
4 15 4 11 2
4 3 13 11 2
8 15 4 10 9 1 15 8 2
7 15 4 10 9 1 11 2
5 15 4 10 11 2
8 10 0 9 2 15 4 15 2
13 1 15 9 13 10 0 9 15 2 8 2 3 2
6 0 13 1 15 9 2
9 15 4 10 0 9 1 0 9 2
7 1 15 9 4 8 9 2
5 13 10 0 9 2
4 3 13 11 2
6 10 9 13 1 11 2
7 15 4 9 1 10 11 2
5 15 4 10 11 2
6 3 4 10 11 4 2
6 10 9 13 1 11 2
8 1 15 0 9 4 10 11 2
7 15 4 10 9 1 11 2
10 15 4 10 9 1 10 0 9 11 2
7 1 15 9 4 15 8 2
10 3 13 10 9 1 10 0 9 8 2
6 13 10 9 1 11 2
4 15 4 11 2
5 15 4 10 11 2
6 1 15 9 13 11 2
8 1 15 0 9 4 15 8 2
4 15 4 8 2
4 15 4 8 2
7 15 4 9 1 10 9 2
4 15 4 8 2
8 15 4 10 0 9 1 9 2
4 13 10 9 2
7 15 4 9 1 10 11 2
10 15 4 10 0 9 1 10 0 9 2
9 15 4 10 9 1 10 9 11 2
6 1 15 9 13 11 2
4 15 4 11 2
9 3 13 3 10 9 9 1 11 2
5 16 4 8 0 2
8 3 13 10 9 1 10 9 2
11 3 13 10 9 1 10 9 7 9 8 2
7 15 4 10 9 1 11 2
7 15 4 10 9 1 11 2
8 1 15 0 9 4 8 9 2
4 15 4 8 2
5 10 9 13 11 2
4 15 4 11 2
7 15 13 15 8 1 11 2
7 3 13 10 9 1 11 2
10 3 13 10 9 1 10 0 9 8 2
6 1 15 9 13 8 2
7 3 13 10 9 1 11 2
7 15 4 10 9 1 11 2
6 1 15 9 13 8 2
7 15 9 4 9 1 11 2
11 15 4 10 9 1 10 0 9 1 13 2
6 13 10 9 1 11 2
10 1 15 9 4 10 0 9 11 4 2
4 15 4 8 2
7 1 15 9 4 8 0 2
7 3 13 10 9 11 8 2
11 3 13 10 9 1 10 13 0 9 8 2
7 3 4 10 9 8 4 2
4 15 4 8 2
9 3 13 11 1 10 9 1 11 2
6 3 4 10 11 4 2
8 15 4 9 1 10 11 9 2
4 15 4 8 2
8 1 15 9 13 10 9 11 2
8 3 13 10 9 1 15 8 2
8 13 15 1 10 9 1 11 2
8 1 15 9 4 10 11 4 2
5 15 4 8 9 2
4 15 4 8 2
7 15 4 10 0 0 9 2
7 15 4 10 9 1 11 2
7 3 13 10 9 11 3 2
4 3 13 8 2
6 1 15 4 8 4 2
9 15 4 10 9 1 10 9 11 2
8 1 15 0 9 4 8 9 2
8 3 0 4 10 0 9 8 2
7 15 4 9 1 15 8 2
9 3 13 8 15 1 9 1 11 2
4 15 4 8 2
11 3 13 10 9 2 11 2 1 11 3 2
7 1 15 9 13 8 3 2
10 15 13 10 0 9 1 10 0 11 2
9 15 9 9 1 10 9 1 8 2
4 13 10 9 2
6 3 13 10 0 9 2
9 15 4 10 0 9 1 15 9 2
4 15 13 11 2
9 15 9 4 10 0 9 1 8 2
8 15 4 10 0 9 1 9 2
4 15 4 11 2
4 15 4 8 2
4 15 13 11 2
4 15 4 11 2
7 3 13 8 1 10 9 2
7 15 4 10 9 1 8 2
4 16 4 8 0
5 3 4 8 0 2
6 3 13 10 0 9 2
4 15 4 11 2
12 15 4 10 9 1 10 9 1 9 1 11 2
7 10 9 4 3 1 11 2
5 10 9 13 9 2
8 3 13 11 10 9 1 11 2
6 16 4 11 10 9 2
10 15 4 10 9 1 10 9 1 11 2
5 16 13 8 11 2
8 3 4 10 9 1 15 8 2
4 15 4 8 2
4 15 4 11 2
7 15 13 11 11 11 4 2
8 15 9 13 15 9 1 11 2
5 3 4 8 4 2
5 15 13 11 3 2
7 15 4 10 9 1 11 2
4 15 4 11 2
7 15 4 10 9 1 11 2
11 15 4 10 9 1 10 0 9 1 8 2
10 15 13 1 12 4 16 9 1 11 2
5 16 4 8 4 2
5 15 13 8 4 2
7 15 9 13 1 8 4 2
4 15 4 8 2
7 15 13 1 12 10 9 2
3 15 4 8
6 15 4 9 1 11 2
7 15 4 11 0 0 9 2
15 3 0 4 10 9 1 10 0 9 7 9 11 1 12 2
7 3 13 11 10 0 11 2
8 3 4 8 2 11 2 4 2
11 10 9 13 1 11 1 10 9 1 12 2
10 15 9 1 15 9 13 11 1 11 2
4 3 4 8 2
4 15 4 9 2
5 3 4 15 4 2
5 10 9 13 9 2
21 15 13 3 1 12 9 1 4 16 3 1 13 1 10 9 1 0 11 1 8 2
4 15 4 8 2
7 3 4 10 9 1 8 2
5 16 4 15 4 2
7 15 4 10 9 1 11 2
7 10 9 13 3 3 11 2
7 3 4 10 9 1 11 2
5 10 9 13 11 2
4 15 4 8 2
11 16 13 10 9 1 10 0 9 11 3 2
4 15 9 13 8
5 15 9 13 8 2
5 16 4 8 4 2
7 3 4 10 9 1 8 2
7 15 4 10 9 1 11 2
4 15 4 8 2
10 1 15 9 13 11 15 9 1 12 2
4 15 4 8 2
7 15 13 4 4 1 8 2
4 15 4 11 2
9 3 13 11 0 9 1 11 4 2
4 15 4 8 2
9 3 4 15 8 2 11 2 4 2
5 15 4 10 11 2
10 3 13 10 0 9 1 0 0 9 2
4 15 4 11 2
4 15 4 11 2
6 15 13 10 11 9 2
10 3 13 10 0 9 11 1 10 9 2
7 15 9 4 1 8 4 2
7 15 4 8 2 11 2 2
6 15 13 10 9 11 2
4 15 13 11 2
9 3 4 11 1 10 15 9 0 2
8 15 4 10 0 9 1 9 2
8 15 4 10 0 9 1 11 2
7 15 4 10 9 1 11 2
9 3 4 10 11 0 4 1 12 2
10 15 4 3 1 12 4 1 10 11 2
9 15 13 2 8 2 1 11 4 2
7 3 13 12 9 1 11 2
8 15 9 13 15 3 1 11 2
7 3 4 15 11 13 4 2
9 15 4 3 4 1 11 1 11 2
9 15 4 4 1 9 1 15 8 2
6 15 13 10 9 11 2
4 15 13 11 2
9 3 13 12 9 1 15 8 13 2
8 3 4 10 11 1 11 4 2
10 15 4 10 9 1 10 11 1 11 2
6 15 13 8 1 11 2
8 15 9 13 10 9 1 8 2
8 15 4 3 4 1 15 8 2
4 15 4 8 2
4 15 4 11 2
10 3 13 10 9 1 11 9 1 11 2
4 3 4 11 2
8 15 4 10 0 9 1 9 2
11 16 4 10 9 1 10 9 9 1 11 2
4 15 4 8 2
4 3 4 8 2
10 10 9 13 3 8 10 9 1 11 2
5 15 4 15 8 2
4 3 13 11 2
7 16 4 15 8 1 11 2
11 3 13 10 9 15 1 12 1 11 13 2
11 15 13 10 0 9 1 10 9 1 11 2
8 3 13 11 8 9 1 12 2
8 3 4 10 9 1 10 11 2
8 1 3 13 11 3 1 11 2
5 3 13 8 9 2
7 10 9 9 3 1 11 2
4 15 4 8 2
4 15 4 11 2
8 3 13 10 9 1 8 9 2
9 15 4 10 9 1 2 11 2 2
6 3 13 10 0 9 2
4 15 4 8 2
7 15 13 15 8 1 12 2
4 15 4 8 2
6 10 9 13 1 11 2
16 10 9 13 15 1 11 4 1 4 16 10 0 9 1 13 2
4 15 4 8 2
5 15 4 10 11 2
6 3 4 15 8 4 2
4 15 4 11 2
7 3 13 10 9 1 11 2
12 16 1 12 13 10 0 0 9 9 1 11 2
7 15 9 13 8 1 12 2
8 3 4 10 9 1 8 4 2
9 3 13 10 0 9 1 11 9 2
11 15 4 4 1 9 1 15 8 1 11 2
7 1 15 9 4 8 9 2
12 3 13 10 9 1 11 15 1 8 4 4 2
8 1 3 4 9 4 1 11 2
8 15 4 10 0 9 1 8 2
8 15 4 10 0 9 1 11 2
6 3 13 15 8 9 2
6 3 4 15 0 8 2
7 15 4 10 9 1 11 2
8 10 9 13 8 4 1 8 2
8 3 13 10 0 9 1 9 2
4 15 4 11 2
5 15 4 10 11 2
4 15 4 8 2
4 15 4 8 2
9 13 10 9 3 8 3 13 4 2
8 10 9 13 15 1 9 4 2
9 15 9 13 2 8 2 1 12 2
11 15 13 10 9 1 11 16 15 4 4 2
10 15 4 10 9 1 15 8 1 11 2
7 15 13 15 0 8 4 2
11 1 15 9 13 10 0 9 3 1 11 2
5 16 4 8 0 2
8 15 13 10 11 1 11 4 2
5 16 4 8 0 2
14 3 13 11 10 9 1 4 1 10 9 1 10 9 2
8 3 4 10 9 1 10 11 2
7 1 15 0 9 13 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 11 2
5 15 4 10 11 2
10 15 9 13 10 0 9 1 10 11 2
5 16 4 8 0 2
4 15 4 8 2
4 15 4 11 2
8 15 9 13 15 13 1 11 2
5 15 9 13 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
12 1 15 9 13 10 9 11 1 15 0 9 2
12 15 9 4 1 15 0 8 16 0 9 4 2
13 15 9 4 1 12 4 16 9 1 10 0 9 2
4 15 4 8 2
4 15 4 11 2
10 15 9 0 1 9 4 16 0 4 2
9 15 9 13 13 7 9 1 9 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
4 15 4 8 2
7 15 4 10 9 1 11 2
7 15 0 9 13 10 11 2
7 15 4 10 9 1 8 2
11 15 0 9 13 10 9 1 10 11 3 2
6 1 15 4 11 13 2
6 1 15 9 13 11 2
6 15 9 13 1 11 2
8 1 15 9 13 10 9 11 2
4 3 13 11 2
6 1 15 9 13 11 2
6 1 15 9 13 11 2
7 3 13 10 9 11 3 2
6 15 9 13 9 11 2
5 15 13 1 12 2
16 1 15 9 13 10 9 7 11 1 10 9 1 10 9 12 2
4 15 4 8 2
6 1 15 9 13 8 2
5 15 4 10 11 2
7 15 4 10 9 1 8 2
6 15 13 10 9 8 2
5 15 13 9 8 2
11 1 15 9 13 8 12 9 0 1 11 2
7 15 4 10 9 1 11 2
9 1 15 9 4 11 16 9 4 2
8 1 15 9 13 15 0 8 2
4 3 13 8 2
7 3 13 10 9 1 11 2
8 15 4 10 9 1 10 11 2
16 3 4 10 9 15 1 12 4 4 16 10 9 8 1 13 2
8 15 4 4 1 8 1 12 2
11 3 13 10 9 3 15 13 9 4 4 2
5 15 4 10 11 2
8 15 4 0 9 1 10 11 2
4 15 4 11 2
4 3 13 11 2
8 15 9 13 15 8 1 12 2
14 3 13 15 15 9 10 9 1 10 9 1 10 11 2
5 15 4 10 11 2
6 15 13 3 1 12 2
5 15 4 10 11 2
8 15 4 10 0 9 1 9 2
8 15 4 10 9 1 10 11 2
4 15 4 8 2
11 3 0 4 8 16 15 1 9 4 4 2
7 10 9 13 10 9 8 2
4 15 4 11 2
8 15 4 10 0 9 1 9 2
4 15 4 8 2
5 13 10 0 9 2
8 15 4 10 0 9 1 12 2
10 3 4 10 9 1 0 9 11 4 2
5 15 4 15 8 2
5 15 4 15 8 2
5 3 13 15 8 2
7 13 10 0 9 1 9 2
10 15 4 10 0 9 1 10 0 9 2
9 15 4 10 0 9 1 10 11 2
4 15 4 8 2
16 15 4 9 1 10 9 15 10 0 9 2 15 8 2 13 2
8 3 13 10 0 9 1 11 2
7 3 4 11 10 9 3 2
4 15 4 8 2
10 15 9 4 0 1 10 9 1 9 2
11 3 13 10 9 1 11 1 9 1 9 2
5 3 13 10 9 2
10 3 4 10 9 7 9 1 15 8 2
6 15 4 0 1 12 2
5 13 10 0 9 2
4 3 13 8 2
4 3 13 8 2
4 3 13 8 2
5 13 10 0 9 2
4 15 4 8 2
6 3 13 10 0 9 2
6 1 15 9 13 11 2
5 15 4 10 11 2
7 3 13 10 9 1 11 2
4 15 4 11 2
4 15 4 11 2
8 15 4 10 0 9 1 9 2
5 10 9 13 11 2
4 3 13 11 2
7 15 4 10 9 1 11 2
5 3 4 8 0 2
6 15 4 8 0 9 2
7 3 13 10 0 0 9 2
7 15 4 10 9 1 11 2
8 15 9 4 11 0 0 9 2
4 15 4 8 2
10 15 4 10 9 1 15 8 1 12 2
5 13 10 0 9 2
4 15 4 11 2
8 15 4 10 0 9 1 9 2
4 15 4 8 2
8 15 9 4 9 1 15 8 2
4 15 4 8 2
4 15 4 8 2
9 15 4 10 9 1 11 1 12 2
4 15 4 8 2
4 15 4 8 2
9 15 4 10 9 1 11 1 12 2
5 13 10 0 9 2
4 15 4 8 2
11 15 0 9 13 9 1 10 9 1 11 2
9 10 9 13 0 9 1 15 8 2
4 15 4 8 2
7 3 0 4 8 1 12 2
15 10 0 9 1 9 13 3 1 12 7 12 1 10 9 2
7 3 13 15 8 15 9 2
5 15 9 13 8 2
9 15 13 10 9 1 9 1 12 2
4 15 4 8 2
6 3 13 8 0 9 2
5 3 13 8 9 2
9 1 15 9 4 8 9 1 11 2
8 3 13 10 0 9 1 11 2
7 15 4 10 9 1 11 2
4 15 4 8 2
7 15 4 10 9 1 11 2
16 1 15 9 4 11 10 9 16 15 1 12 4 4 1 11 2
10 3 13 10 9 1 10 9 1 11 2
9 1 15 9 4 11 1 11 4 2
5 15 4 10 11 2
5 3 13 9 3 2
9 15 9 4 10 9 1 15 8 2
4 15 4 8 2
4 3 13 11 2
5 15 4 15 8 2
5 15 4 10 11 2
5 13 10 0 9 2
6 15 13 2 8 2 2
6 1 15 9 13 8 2
8 15 4 10 9 1 15 8 2
7 15 4 10 9 1 11 2
7 15 4 10 9 1 11 2
7 15 4 10 9 1 11 2
9 15 9 4 8 0 9 1 9 2
5 15 9 13 8 2
7 15 13 10 9 1 11 2
4 15 4 8 2
4 3 13 8 2
8 3 0 4 8 16 15 13 2
4 3 13 11 2
6 3 0 4 15 8 2
8 15 4 10 0 9 1 11 2
9 10 9 13 1 11 1 10 9 2
7 15 9 13 3 1 8 2
9 15 4 10 9 1 10 9 11 2
8 3 0 13 8 1 10 9 2
5 15 4 10 11 2
9 15 13 15 8 1 12 1 12 2
12 15 4 10 0 9 1 9 1 12 1 12 2
7 1 15 9 13 15 9 2
21 3 13 10 9 9 4 15 4 4 1 10 9 1 10 9 1 10 15 7 9 2
14 3 4 10 0 1 3 0 9 4 15 15 9 13 2
7 15 0 9 13 1 9 2
16 13 10 15 9 1 10 9 15 0 9 13 7 15 9 13 2
8 6 2 15 9 13 3 0 2
8 3 4 10 0 9 1 8 2
9 15 0 9 13 1 11 1 8 2
9 15 9 13 15 1 10 9 13 2
13 1 15 9 13 10 13 9 3 2 2 8 2 2
12 1 10 9 13 15 1 10 9 10 9 4 2
7 1 15 9 4 11 4 2
13 15 0 9 4 10 0 9 1 10 0 0 9 2
11 1 15 9 1 0 9 13 15 8 0 2
9 15 13 9 2 9 7 9 0 2
7 13 10 15 9 1 9 2
9 6 2 15 9 13 1 10 9 2
14 3 4 10 9 7 9 15 13 1 10 9 1 12 2
8 3 4 11 1 10 0 9 2
17 3 13 10 9 4 1 10 9 7 0 9 1 10 9 4 4 2
12 1 15 9 13 10 9 11 1 12 0 3 2
18 1 15 9 1 10 9 1 11 13 10 9 3 0 15 8 4 4 2
9 1 15 9 4 10 11 0 4 2
7 15 0 9 4 8 4 2
13 16 15 13 1 9 2 3 4 15 3 0 3 2
6 3 4 10 9 4 2
9 13 10 0 9 1 2 9 2 2
9 6 2 15 9 9 13 1 11 2
23 3 4 10 9 15 1 10 9 1 12 1 10 11 13 7 15 10 9 16 0 9 13 2
8 1 15 9 13 10 9 11 2
10 15 9 4 3 3 10 0 9 4 2
7 15 9 13 8 1 12 2
13 15 0 9 4 0 1 13 9 2 9 7 9 2
9 3 13 10 9 1 10 0 9 2
14 15 0 9 7 9 4 15 1 10 0 9 1 8 2
8 1 15 13 10 0 9 11 2
9 8 9 4 10 9 11 7 11 2
9 13 10 9 1 10 0 9 9 2
10 6 2 15 9 13 15 1 9 4 2
16 3 13 10 9 15 1 10 0 9 1 10 9 1 8 13 2
9 1 15 0 9 13 10 9 11 2
6 15 4 10 0 9 2
11 3 13 10 3 0 9 1 8 1 12 2
18 10 0 9 8 4 3 1 10 9 1 4 2 15 13 3 10 9 2
10 15 0 9 13 3 4 4 1 9 2
17 15 0 9 13 4 4 16 10 0 9 1 10 0 9 1 11 2
9 1 15 9 13 10 0 9 11 2
18 3 13 15 10 9 15 1 10 9 15 0 2 7 10 0 9 13 2
10 3 13 10 0 9 3 10 9 13 2
9 6 2 15 9 13 1 10 9 2
18 3 4 10 9 3 1 10 0 2 3 13 9 2 9 2 4 4 2
14 15 0 9 4 4 1 10 9 8 2 11 7 11 2
10 15 9 13 1 10 0 9 1 9 2
6 15 9 4 8 4 2
15 15 9 13 10 11 12 2 12 7 12 1 15 9 4 2
13 15 4 10 9 1 10 9 1 11 1 12 9 2
16 15 13 15 1 10 9 7 4 1 12 9 1 11 1 11 2
22 3 13 10 9 7 10 9 1 10 9 7 10 9 4 15 8 1 10 9 4 4 2
11 3 4 9 7 9 4 15 10 9 13 2
14 3 13 10 9 1 10 9 11 7 11 1 15 8 2
7 13 10 0 9 1 9 2
12 3 13 10 0 9 1 10 9 1 10 9 2
9 15 0 9 13 3 8 8 4 2
6 10 9 13 10 9 2
16 15 9 1 8 4 1 12 9 1 11 4 2 13 12 2 2
7 1 15 9 13 10 9 2
9 1 15 9 4 8 10 0 9 2
16 1 15 0 0 1 10 0 9 4 10 9 1 0 9 4 2
13 1 15 9 1 8 1 12 13 8 10 0 9 2
6 8 9 4 10 9 2
14 3 13 10 9 15 13 1 15 13 7 13 1 9 2
7 13 10 0 9 1 9 2
11 3 13 10 9 1 10 0 0 0 9 2
13 15 9 13 1 10 9 1 10 11 7 10 9 2
4 15 4 11 2
8 1 15 9 13 8 4 13 2
8 3 13 10 9 1 10 9 2
7 3 13 11 3 1 12 2
14 15 0 0 1 10 0 9 13 10 9 1 10 11 2
12 3 4 10 0 0 9 2 13 1 0 9 2
8 15 9 13 10 0 9 8 2
10 3 13 10 0 7 0 9 1 11 2
9 13 10 15 9 1 2 13 2 2
15 3 13 10 9 3 10 0 9 8 1 12 15 8 13 2
7 1 15 0 9 13 11 2
8 1 15 9 13 10 9 11 2
11 15 0 9 1 12 4 8 9 16 9 2
12 15 9 13 1 11 12 10 9 1 11 0 2
15 3 4 10 9 15 1 10 9 4 4 1 9 7 9 2
13 15 13 1 12 8 10 0 9 10 9 1 11 2
12 1 15 9 4 1 12 15 8 1 11 4 2
11 15 12 9 13 15 16 10 9 1 13 2
15 3 13 10 0 9 3 10 9 7 15 15 15 9 13 2
10 13 10 15 9 3 13 2 13 9 2
19 3 4 10 9 1 9 8 2 15 10 9 13 1 10 9 2 8 2 2
12 1 15 9 13 10 11 15 1 12 4 4 2
16 15 0 9 13 16 3 15 9 4 16 15 9 0 13 4 2
11 3 4 10 9 3 8 10 0 9 13 2
6 3 4 9 3 4 2
21 3 13 10 9 1 10 9 10 9 1 12 9 3 15 9 2 9 7 9 13 2
6 15 9 13 10 0 2
9 15 0 9 13 10 9 1 11 2
11 15 12 9 13 15 16 10 9 1 13 2
20 3 4 10 9 1 10 9 1 10 0 9 2 13 1 10 9 1 10 9 2
9 13 10 15 9 1 0 7 9 2
7 3 4 10 9 1 8 2
10 1 15 12 9 13 10 9 1 11 2
8 15 9 13 10 0 9 11 2
11 15 9 1 12 13 10 9 1 10 9 2
8 15 0 9 13 15 0 8 2
11 1 15 9 4 1 12 15 0 8 4 2
9 15 4 10 0 9 1 10 11 2
8 1 15 13 10 9 15 9 2
5 3 13 9 9 2
13 3 13 10 9 15 10 10 9 13 1 10 9 2
20 3 4 10 0 2 0 2 13 9 3 1 0 9 3 15 13 15 9 13 2
7 13 10 15 9 1 9 2
18 3 4 10 9 3 10 9 1 10 3 0 9 1 10 9 4 4 2
20 1 10 0 9 4 12 0 9 4 2 8 2 11 2 11 7 2 2 2 2
10 15 13 15 15 0 4 1 10 9 2
10 1 15 9 13 8 1 12 10 11 2
19 15 9 9 2 15 0 1 9 13 2 4 3 15 9 4 2 8 9 2
13 3 13 10 9 4 15 1 12 1 11 9 13 2
11 15 0 9 13 1 12 10 9 1 8 2
19 1 15 9 1 10 11 13 10 9 1 10 0 9 10 9 1 10 9 2
6 3 4 10 0 9 2
12 3 13 10 9 1 0 15 4 4 1 8 2
7 13 10 15 9 1 9 2
21 3 4 10 9 3 9 1 9 4 4 7 10 0 9 1 9 7 9 4 4 2
9 1 15 9 1 11 13 10 9 2
11 1 10 9 13 3 9 1 10 0 9 2
14 1 15 1 15 13 9 13 8 10 9 1 0 9 2
15 15 4 10 9 1 15 8 2 11 2 1 12 1 12 2
20 15 0 9 13 9 16 9 8 1 12 1 0 9 1 11 7 11 0 4 2
12 15 13 1 12 10 0 9 1 9 4 4 2
15 16 15 15 9 13 15 3 1 10 9 15 10 9 9 2
27 3 13 15 10 0 9 1 10 0 9 1 10 9 15 10 0 9 3 13 4 2 7 3 3 1 15 9
9 3 13 10 9 16 11 3 4 2
9 13 10 0 9 1 2 9 2 2
17 3 13 10 9 1 15 9 8 2 15 12 1 15 9 4 13 2
5 15 4 10 9 2
6 10 11 13 15 8 2
11 15 9 1 11 13 8 1 16 9 8 2
7 15 9 4 1 8 4 2
12 15 0 9 13 9 3 1 10 0 0 11 2
16 15 13 1 10 0 9 15 0 9 1 10 9 11 11 2 2
7 1 15 13 8 15 9 2
12 3 13 15 9 15 0 13 8 9 1 9 2
15 3 13 10 9 1 10 9 2 15 4 4 13 1 9 2
16 3 13 10 0 9 15 4 4 1 10 9 1 11 7 11 2
8 3 13 10 9 3 8 13 2
18 3 4 10 0 9 1 10 9 10 9 16 13 15 3 15 4 4 2
7 15 13 10 0 9 3 2
9 15 9 1 11 4 13 1 11 2
12 10 9 1 9 7 13 2 3 4 15 9 2
13 15 9 13 1 12 16 0 9 9 1 10 9 2
12 15 9 4 16 10 9 1 8 10 9 4 2
10 1 15 9 4 0 4 1 10 9 2
11 3 13 10 0 9 1 9 3 3 4 2
16 3 13 10 9 1 10 9 3 10 9 13 0 9 1 4 2
19 3 13 10 1 9 13 9 1 7 1 10 9 3 10 9 13 9 13 2
14 3 4 10 9 3 9 1 10 9 13 1 15 9 2
8 1 15 9 4 11 10 9 2
15 3 4 10 9 4 15 10 0 9 13 1 10 15 9 2
17 1 15 9 1 10 9 1 9 8 2 1 11 4 8 8 0 2
19 1 9 13 15 10 9 4 16 15 13 4 2 1 15 9 13 15 3 2
9 15 4 10 0 9 1 15 8 2
10 15 9 13 1 10 9 1 9 11 2
18 3 4 1 10 9 10 9 1 9 4 15 4 4 1 10 15 9 2
9 3 4 10 13 9 3 3 4 2
8 3 4 10 9 1 10 9 2
10 3 13 10 0 9 1 10 0 9 2
10 3 13 10 9 4 8 1 10 0 2
6 1 15 9 13 11 2
10 3 4 10 9 1 9 7 13 4 2
16 15 4 10 9 1 10 0 9 1 12 9 1 8 1 12 2
13 1 15 9 13 8 10 0 9 0 7 9 4 2
7 15 4 10 0 0 9 2
11 15 0 9 4 4 16 10 9 1 11 2
13 1 15 0 0 9 1 10 9 13 8 7 8 2
14 3 4 1 10 9 1 0 9 10 0 13 9 4 2
16 3 13 10 9 15 10 9 9 8 13 2 16 15 13 4 2
19 3 13 10 0 2 13 9 1 10 9 7 1 10 0 9 1 10 9 2
14 3 13 10 9 1 9 1 12 7 12 3 8 13 2
7 15 4 10 9 1 11 2
17 15 9 13 1 10 9 1 10 0 9 15 1 12 9 8 13 2
11 15 9 1 11 4 4 1 13 0 9 2
10 15 9 13 15 9 1 15 0 8 2
9 1 15 9 13 10 0 0 9 2
14 15 9 4 1 12 10 0 15 15 8 1 9 13 2
20 1 15 9 13 9 8 2 10 0 9 1 11 1 10 11 9 1 12 8 2
12 3 4 9 15 3 1 9 13 3 3 4 2
22 3 4 10 9 1 10 0 9 2 15 10 9 4 1 10 9 11 7 10 9 11 2
12 3 13 10 2 0 2 9 1 10 0 9 2
13 3 13 10 9 3 11 1 10 9 1 8 13 2
7 1 15 9 13 10 11 2
8 15 4 10 9 1 10 9 2
21 8 13 3 1 7 13 10 11 1 10 0 9 1 10 9 1 12 2 15 9 2
14 1 15 9 1 11 4 7 9 1 9 16 13 4 2
17 15 9 13 4 4 16 10 0 9 1 9 2 12 9 1 9 2
13 15 13 9 1 0 9 1 10 9 11 8 2 2
14 15 4 10 9 1 10 0 13 9 15 1 12 13 2
10 1 10 9 13 10 9 1 10 9 2
17 3 13 10 0 0 9 3 0 2 0 9 1 10 9 4 4 2
10 3 13 10 0 9 1 10 0 9 2
10 3 13 10 9 1 8 15 0 13 2
10 3 4 10 9 1 10 9 1 11 2
7 3 13 10 9 11 3 2
9 1 15 9 1 12 13 8 3 2
11 15 0 9 4 0 1 10 0 9 0 2
12 15 0 9 13 10 9 1 10 0 9 11 2
18 15 9 13 9 8 2 2 3 15 13 16 10 9 3 15 9 4 2
16 15 0 9 13 4 1 15 9 1 10 0 9 1 10 9 2
7 3 13 10 9 0 3 2
18 3 13 10 0 9 1 11 2 15 15 3 1 10 9 13 1 12 2
18 3 13 10 9 16 0 2 1 0 9 10 0 9 0 9 1 4 2
23 3 4 10 9 1 9 1 1 10 9 2 10 9 1 10 9 12 1 10 9 7 9 2
12 15 9 1 10 0 11 4 1 10 9 11 2
10 15 9 4 0 10 0 9 1 9 2
25 11 8 2 2 11 8 2 2 11 11 2 7 9 8 2 13 3 10 0 9 2 15 4 10 9
16 3 13 10 9 15 4 4 1 9 15 15 13 4 7 4 2
19 3 13 10 9 9 3 10 0 10 9 15 16 12 9 3 0 0 13 2
20 15 9 13 1 10 9 11 8 2 1 12 7 13 3 8 1 9 8 2 4
11 1 15 9 13 10 9 10 9 11 4 2
11 15 4 8 10 0 9 15 1 9 9 2
7 3 13 10 9 0 3 2
8 3 13 10 9 10 0 9 2
12 3 13 10 1 15 1 0 0 9 1 11 2
19 3 4 15 1 10 0 9 1 11 15 1 4 4 1 10 11 1 11 2
7 15 4 10 9 1 8 2
10 15 9 1 15 9 13 10 9 3 2
13 1 15 9 1 11 13 15 2 8 2 10 9 2
8 3 13 10 0 9 1 8 2
15 1 15 9 4 10 9 16 10 0 9 1 11 13 4 2
14 8 13 1 10 9 1 15 9 4 2 3 4 15 2
8 1 15 9 13 10 9 11 2
6 15 13 10 9 9 2
22 3 13 10 0 9 1 10 11 15 1 11 2 1 9 1 11 2 1 9 4 4 2
19 3 13 10 0 9 3 10 9 1 10 0 9 1 10 9 1 15 13 2
9 3 13 10 9 1 8 1 11 2
9 1 15 9 4 10 0 9 11 2
18 15 0 9 13 3 3 1 9 7 13 10 9 15 2 0 2 13 2
9 15 9 4 4 16 10 0 9 2
21 3 13 10 0 2 0 2 0 0 9 15 3 1 10 9 1 10 9 4 4 2
13 3 4 10 9 1 10 0 9 1 10 0 9 2
13 15 4 2 1 10 0 0 9 10 9 1 11 2
18 16 15 1 11 1 10 2 9 2 13 2 15 13 15 3 3 4 2
9 1 15 0 9 13 10 0 9 2
12 3 13 10 9 1 10 9 1 10 0 9 2
13 3 13 10 0 0 0 9 15 1 10 9 13 2
12 3 13 10 0 9 2 15 4 4 1 8 2
10 1 15 9 4 10 11 10 0 9 2
13 1 15 9 13 10 9 9 1 10 9 1 11 2
18 10 0 9 1 9 4 1 12 4 1 10 9 1 8 2 15 9 2
15 3 13 10 0 9 1 9 2 9 2 9 7 0 9 2
15 1 15 9 4 10 0 9 1 10 11 1 15 8 4 2
10 15 13 8 1 10 9 11 8 2 2
10 1 15 9 13 8 15 1 12 3 2
8 15 13 9 13 3 1 9 2
20 3 4 10 9 2 3 9 7 9 13 13 2 16 15 9 1 11 1 13 2
16 3 4 10 9 3 15 10 9 3 13 7 10 9 13 13 2
18 3 13 10 0 9 1 10 0 9 2 15 3 3 3 1 9 13 2
11 3 13 10 9 1 11 7 10 0 9 2
22 3 4 10 9 1 10 9 3 10 9 3 0 4 15 3 10 9 3 3 13 4 2
17 3 13 10 9 1 8 7 8 1 10 9 1 10 9 1 11 2
7 15 13 15 1 10 9 2
15 3 13 10 9 1 12 4 3 10 9 1 10 9 13 2
12 10 9 1 15 9 4 1 12 4 7 4 2
7 15 4 10 9 1 11 2
11 3 13 10 9 10 9 1 15 9 4 2
11 3 4 10 9 15 10 9 3 13 4 2
11 3 4 10 9 15 3 1 9 4 4 2
13 3 4 15 0 16 4 4 3 7 9 1 8 2
8 3 4 10 9 1 10 11 2
12 15 9 4 10 0 9 1 10 9 1 8 2
10 15 9 1 8 1 12 13 10 9 2
12 1 15 9 13 8 0 9 1 12 1 11 2
14 15 4 10 9 1 10 0 9 15 1 12 4 4 2
16 15 13 10 9 8 8 2 3 1 10 9 1 11 1 12 2
22 3 4 0 9 1 3 10 9 2 15 4 4 1 10 9 1 10 9 7 10 9 2
14 15 9 13 15 9 4 1 15 9 7 10 9 11 2
9 3 13 10 0 9 1 10 9 2
19 3 4 10 0 9 15 15 13 1 9 2 7 15 13 4 1 12 9 2
15 3 13 10 9 3 3 8 15 1 15 9 3 13 4 2
11 15 12 9 4 1 12 9 1 10 11 2
10 15 13 16 0 10 9 1 10 9 2
12 1 15 9 4 1 12 15 8 1 11 4 2
12 1 15 9 13 9 1 11 2 11 7 11 2
8 15 4 10 0 9 1 11 2
6 15 13 10 0 11 2
9 1 15 9 1 11 13 8 9 2
10 3 4 10 9 1 10 9 11 4 2
7 3 4 15 0 9 13 2
15 3 4 10 9 15 4 4 1 9 1 13 9 1 9 2
8 3 13 15 0 9 1 11 2
6 1 15 9 13 11 2
13 3 4 10 0 13 9 15 15 1 10 9 13 2
9 1 15 9 4 10 9 8 8 2
18 15 0 9 13 15 1 15 9 13 2 9 2 9 2 9 7 9 2
14 1 15 0 9 13 10 0 9 11 1 12 9 3 2
15 15 4 1 9 4 3 15 13 1 4 1 10 0 9 2
12 10 9 13 11 1 15 8 1 12 1 11 2
9 1 15 9 13 15 10 9 4 2
16 3 13 10 9 1 11 3 1 10 9 13 7 9 4 4 2
15 3 4 10 0 2 0 9 15 10 15 9 7 9 13 2
15 3 13 10 9 1 8 15 1 12 1 10 9 4 4 2
11 15 12 9 4 1 12 9 1 10 11 2
7 1 15 9 13 10 9 2
16 1 12 13 10 0 9 8 10 9 1 10 11 2 15 9 2
8 1 15 9 13 8 7 8 2
9 3 4 10 9 1 11 1 11 2
11 15 13 8 7 4 10 9 1 15 8 2
11 10 9 13 1 12 9 3 1 10 9 2
20 15 9 13 13 3 16 0 16 15 15 0 7 0 9 0 1 15 9 4 2
17 3 4 15 0 16 9 13 2 13 1 10 9 1 10 9 2 2
8 3 4 10 9 1 10 0 2
10 3 4 10 9 1 11 1 9 8 2
13 15 13 1 12 8 3 16 9 1 10 0 9 2
15 15 9 13 1 15 13 2 10 9 15 9 15 9 13 2
21 10 9 1 8 4 1 12 4 1 8 7 8 1 10 9 2 3 4 15 9 2
12 1 15 9 13 10 9 11 2 11 7 8 2
17 10 9 1 15 9 4 4 7 4 1 10 11 1 12 1 12 2
14 15 0 9 13 1 9 4 7 13 1 12 1 11 2
12 15 0 0 4 1 15 9 1 10 9 4 2
5 15 4 10 9 2
21 3 13 10 9 1 10 9 1 10 9 1 15 8 2 3 3 10 0 9 11 2
12 3 4 10 9 3 15 9 7 9 13 4 2
9 3 4 10 9 1 8 1 11 2
13 13 12 9 15 1 12 3 3 13 1 10 9 2
10 1 15 0 9 4 9 0 15 4 2
11 3 4 10 0 9 15 8 7 8 13 2
7 1 15 9 4 8 0 2
11 15 4 10 9 1 10 13 9 1 11 2
12 15 4 9 1 11 16 11 1 10 9 13 2
7 1 15 9 13 10 11 2
9 3 13 10 9 1 10 0 9 2
8 1 15 9 13 15 10 9 2
23 3 4 15 0 0 9 1 10 0 9 1 10 9 2 15 1 10 0 9 1 11 13 2
15 3 4 10 0 9 13 0 11 2 0 1 10 0 11 2
13 3 4 10 9 15 11 0 1 10 0 9 13 2
7 1 15 9 13 10 9 2
18 1 10 9 1 15 9 13 0 9 10 9 16 1 15 9 1 13 2
14 1 15 9 13 10 9 11 8 2 10 9 1 9 2
20 10 9 1 10 11 9 12 13 15 3 0 1 10 11 4 2 15 4 15 2
7 15 4 15 2 8 2 2
13 15 0 9 13 10 9 1 10 9 1 10 9 2
12 1 15 0 9 13 8 7 10 9 8 3 2
14 15 9 4 10 0 9 1 11 3 10 9 3 13 2
27 3 13 10 9 1 10 0 9 2 15 1 3 10 9 4 2 1 10 9 10 9 7 1 3 10 9 2
16 3 4 10 9 3 10 9 13 4 1 15 1 10 15 9 2
10 3 4 10 9 15 8 1 12 13 2
16 3 4 15 9 1 15 8 2 15 13 1 10 11 7 11 2
14 3 13 15 10 9 3 10 9 3 12 9 0 4 2
16 1 12 13 8 10 11 1 10 0 0 9 2 1 15 9 2
12 1 15 9 13 11 2 11 2 11 7 11 2
14 15 9 1 11 13 15 1 12 3 1 4 1 11 2
10 15 0 9 13 10 9 1 10 9 2
5 15 9 3 13 2
10 1 15 9 13 9 2 9 7 9 2
9 3 13 10 0 9 1 15 8 2
14 3 13 10 9 2 3 15 15 15 4 2 4 4 2
7 3 4 10 9 1 8 2
11 3 4 10 10 9 1 10 0 11 4 2
10 15 9 13 1 9 7 9 1 9 2
17 3 4 10 0 9 1 10 11 15 9 9 12 1 8 4 4 2
9 15 0 9 4 8 4 1 12 2
8 15 4 4 1 10 9 8 2
14 15 0 9 1 10 0 9 13 10 9 1 10 9 2
10 1 15 9 4 10 9 8 3 0 2
12 1 15 9 4 3 12 9 2 9 7 9 2
16 3 4 15 0 9 16 9 2 13 7 9 13 4 7 4 2
15 3 13 10 9 1 10 0 9 15 13 1 0 0 9 2
9 3 4 10 9 1 10 9 8 2
8 1 15 9 13 10 9 11 2
9 15 9 1 10 9 13 10 9 2
9 15 9 13 10 9 11 1 12 2
7 15 9 13 10 0 9 2
12 15 9 4 1 12 4 1 8 7 15 9 2
8 15 0 9 13 1 10 9 2
9 15 4 10 9 1 10 9 11 2
11 15 13 10 9 3 2 3 13 0 4 2
16 3 13 10 9 15 1 10 0 9 7 10 9 10 9 13 2
7 3 4 15 15 9 13 2
13 3 4 10 9 15 10 9 13 1 10 0 9 2
13 3 13 10 9 1 9 3 9 7 9 4 4 2
10 1 15 9 4 10 11 0 10 9 2
7 15 4 15 0 0 8 2
18 15 4 10 9 1 15 9 1 0 9 2 3 9 2 9 7 9 2
15 3 4 10 0 9 7 9 15 4 4 1 10 9 8 2
13 15 9 1 10 0 9 11 4 9 1 15 8 2
8 3 4 10 9 3 3 4 2
10 15 0 9 13 3 16 10 0 9 2
12 3 4 15 13 9 1 10 9 1 10 9 2
11 3 4 1 10 9 10 0 9 7 9 2
11 3 4 10 9 1 10 9 9 1 8 2
18 15 9 13 13 15 3 1 9 1 11 1 1 11 2 11 7 11 2
18 15 9 15 13 13 1 9 7 0 9 1 10 9 4 0 1 9 2
20 3 13 10 9 1 12 3 8 10 0 11 13 16 10 9 0 9 7 9 2
12 15 4 10 0 9 1 10 9 1 10 9 2
13 15 0 9 13 10 0 9 11 1 0 1 8 2
8 15 0 4 1 10 9 4 2
12 15 9 1 8 13 15 9 1 12 1 11 2
9 15 4 10 0 9 1 10 9 2
13 3 4 10 9 1 10 9 11 7 15 9 11 2
22 3 4 10 0 0 9 1 10 9 1 15 9 2 16 1 10 0 9 9 1 13 2
11 3 13 10 9 1 10 13 9 1 8 2
9 15 9 13 1 9 1 15 8 2
9 1 15 9 13 15 13 1 9 2
18 10 9 1 10 9 8 16 9 4 4 1 10 9 1 12 2 15 2
13 3 13 10 9 15 9 4 16 15 12 9 13 2
7 1 15 9 13 8 3 2
12 15 0 9 4 10 0 9 1 10 9 11 2
13 1 10 9 13 10 9 1 13 9 10 9 4 2
6 8 9 4 10 9 2
12 3 4 10 9 1 8 2 15 3 9 4 2
6 3 4 10 0 9 2
21 3 13 15 15 9 2 13 1 10 0 9 2 15 3 4 4 1 10 0 11 2
10 15 4 10 12 9 1 10 0 9 2
10 1 15 0 9 4 10 0 9 0 2
12 1 15 9 13 8 1 12 15 9 16 9 2
14 1 15 0 9 13 9 2 16 7 0 16 9 13 2
23 3 13 15 10 0 9 1 0 9 16 9 13 1 10 9 1 12 1 10 9 1 12 2
10 1 15 13 10 9 8 10 13 9 2
9 1 15 9 13 10 9 15 3 2
10 1 15 9 13 9 1 10 0 9 2
8 3 4 10 0 9 1 11 2
15 3 13 15 10 9 15 3 0 4 1 9 7 0 9 2
14 3 13 15 10 9 1 10 0 9 15 15 9 4 2
15 1 15 9 13 0 10 0 9 1 9 7 0 9 9 2
11 13 10 15 9 1 10 9 1 10 9 2
10 1 15 9 13 10 9 8 1 12 2
8 3 4 15 8 1 12 4 2
6 15 9 1 8 11 2
11 15 0 9 4 0 3 15 2 8 2 2
12 15 0 9 13 1 11 1 15 9 1 11 2
5 15 4 10 9 2
7 3 4 10 9 1 8 2
21 3 13 15 0 10 9 9 3 9 4 4 16 3 1 13 15 10 9 0 4 2
20 3 13 15 10 9 1 10 0 13 9 3 10 9 10 9 1 10 9 13 2
9 1 15 12 9 13 10 9 11 2
8 15 4 10 0 9 1 9 2
18 1 15 9 13 10 11 1 12 7 3 10 9 1 12 10 0 9 2
7 3 4 10 9 1 11 2
12 15 9 4 4 1 10 0 9 11 1 12 2
14 15 1 11 0 0 9 4 10 9 1 10 0 9 2
17 15 0 1 13 9 4 4 1 9 7 9 3 1 13 1 9 2
7 3 4 10 0 9 4 2
16 15 0 9 4 3 1 15 0 9 1 9 1 10 9 4 2
16 3 4 10 0 9 1 10 9 15 1 10 9 10 9 13 2
15 3 13 10 9 10 0 9 1 10 9 13 1 15 9 2
15 3 13 15 10 0 13 9 2 9 7 9 1 0 9 2
13 3 4 10 9 1 0 9 1 11 1 15 8 2
12 3 13 10 0 9 2 16 10 9 0 13 2
13 1 15 9 1 11 13 10 9 3 1 10 9 2
16 15 0 9 4 2 4 2 1 12 1 10 9 8 1 11 2
13 1 15 0 9 13 3 1 10 0 9 1 9 2
10 15 9 4 1 12 1 8 8 4 2
12 1 15 0 9 13 15 10 9 11 8 2 2
12 15 13 10 9 9 2 0 9 7 9 0 2
18 3 4 10 9 15 1 10 9 10 9 13 7 3 9 4 1 4 2
16 3 13 15 9 15 1 15 9 10 9 13 16 15 3 13 2
21 3 13 15 10 0 9 1 9 2 3 9 2 15 4 4 1 0 9 7 9 2
10 3 13 10 0 9 1 10 0 9 2
10 3 13 15 10 9 1 10 9 8 2
7 1 15 9 13 8 3 2
16 3 4 10 9 2 0 9 1 11 15 3 4 4 16 9 2
11 15 0 9 13 1 12 15 9 1 9 2
21 15 9 13 1 10 0 9 1 9 8 3 16 15 9 4 1 15 9 1 11 2
9 15 9 1 10 9 1 10 9 2
4 15 4 13 2
12 3 4 10 9 15 10 0 13 9 9 13 2
13 3 13 15 0 1 0 9 2 8 2 9 2 2
8 3 13 15 10 13 0 9 2
8 15 4 10 0 9 1 11 2
13 15 9 1 10 9 7 10 9 13 9 3 3 2
23 1 12 13 8 10 9 1 10 9 1 10 0 2 0 9 7 9 2 3 13 10 9 2
23 1 15 9 13 15 12 9 1 15 9 4 7 13 10 9 16 12 7 15 9 13 4 2
14 15 0 9 4 0 0 1 10 9 1 10 9 11 2
10 15 13 10 9 1 10 9 1 11 2
15 13 10 15 9 1 2 9 2 2 9 15 16 9 13 2
10 15 4 10 0 9 1 10 0 9 2
11 3 4 10 0 0 9 1 10 9 11 2
17 3 13 15 10 0 9 1 10 9 2 13 16 10 9 1 4 2
12 3 13 15 10 0 7 0 9 1 10 9 2
8 3 13 10 0 9 1 11 2
11 3 13 15 10 0 9 1 10 9 8 2
13 15 9 1 11 13 1 10 9 3 3 0 4 2
13 15 0 9 13 1 9 2 13 1 9 7 9 2
9 15 9 13 9 1 11 1 12 2
9 15 4 10 9 1 10 9 8 2
6 1 15 9 13 11 2
11 8 9 4 9 11 2 10 9 1 8 2
19 3 4 10 9 7 13 1 15 0 8 2 15 3 16 15 10 9 13 2
22 3 13 15 10 0 7 0 9 15 15 13 4 1 15 13 1 10 9 1 10 9 2
13 3 13 15 10 9 1 9 15 1 13 9 13 2
8 1 15 9 13 10 9 11 2
16 15 4 10 0 9 1 15 8 2 10 0 9 1 10 9 2
15 1 15 9 13 10 0 9 7 9 11 1 12 10 11 2
23 15 9 13 10 9 1 10 9 1 13 3 10 9 1 9 13 12 7 15 15 9 4 2
13 15 9 4 11 8 10 9 1 8 1 12 3 2
12 15 9 13 1 12 0 10 9 1 10 9 2
9 3 13 10 9 11 3 1 11 2
11 15 4 10 0 9 15 1 11 4 4 2
7 3 4 10 9 1 8 2
15 3 13 15 10 9 1 9 15 15 13 1 10 0 9 2
15 3 13 15 10 9 16 15 9 13 7 15 3 0 4 2
8 3 4 10 9 11 16 0 2
16 10 9 8 13 9 1 10 9 2 3 4 15 1 10 0 2
11 1 12 13 8 10 9 1 8 2 15 2
11 15 9 4 4 1 10 9 8 1 12 2
10 1 15 0 9 13 10 0 9 8 2
21 15 11 13 1 10 11 10 0 11 7 13 16 11 15 4 4 10 9 1 4 2
12 1 15 9 1 11 13 8 7 8 10 9 2
10 15 4 0 2 9 7 9 1 9 2
9 3 4 10 9 1 11 11 11 2
17 3 13 15 10 9 7 9 1 15 9 1 10 9 9 7 9 2
13 3 13 15 10 9 1 9 7 10 9 1 9 2
8 3 13 10 0 9 1 11 2
16 3 4 15 0 9 1 10 9 1 10 9 3 9 4 4 2
10 1 15 9 9 8 7 8 10 9 2
19 3 13 10 0 9 2 15 13 1 9 7 13 9 13 1 9 7 9 2
10 1 15 9 13 10 9 1 12 8 2
8 15 4 10 9 1 10 9 2
12 10 9 13 15 0 4 1 10 9 1 9 2
8 15 9 4 1 10 9 4 2
11 3 4 10 9 1 11 15 15 9 4 2
17 3 13 15 10 9 1 10 9 7 9 1 10 9 1 10 9 2
15 3 13 15 10 9 1 10 9 2 3 0 9 4 4 2
8 3 4 10 0 9 1 11 2
12 15 0 9 13 10 9 16 10 9 1 13 2
17 1 15 9 13 10 9 11 8 2 1 11 2 11 7 11 3 2
8 15 9 13 15 9 1 8 2
13 15 9 4 1 12 4 1 10 9 2 8 2 2
14 3 4 10 0 9 15 4 13 1 10 11 1 11 2
8 1 15 9 13 10 11 9 2
20 15 0 9 2 3 1 10 0 7 0 9 1 10 9 2 4 3 3 4 2
12 3 4 1 10 0 9 10 9 1 10 9 2
11 3 13 15 10 9 1 15 9 3 13 2
17 3 13 15 10 9 1 0 0 9 2 7 1 9 7 1 9 2
7 15 4 10 9 1 11 2
10 3 13 15 10 9 1 12 0 9 2
15 10 0 9 8 4 3 0 16 10 9 1 12 2 15 2
18 3 13 10 9 3 15 3 0 7 3 0 0 13 4 1 10 9 2
6 15 9 4 0 8 2
9 15 4 10 9 1 15 13 8 2
13 15 4 1 10 9 1 10 9 12 9 1 11 2
11 15 9 13 10 0 9 1 10 9 13 2
6 3 0 13 10 9 2
17 3 13 15 10 9 1 9 7 9 1 9 1 9 2 9 3 2
25 3 13 15 15 13 1 9 2 3 10 9 1 10 9 4 4 1 9 2 3 10 9 4 4 2
8 1 15 9 4 11 10 9 2
11 3 4 10 0 9 1 10 9 1 9 2
15 15 9 1 8 4 4 1 10 9 1 10 0 1 11 2
13 1 15 9 1 13 4 3 15 13 7 9 4 2
16 15 0 9 4 1 12 1 12 10 0 9 1 10 0 9 2
10 15 9 13 15 9 13 1 10 9 2
13 8 4 13 1 10 0 9 2 15 9 13 15 2
7 15 9 13 10 9 0 2
13 15 9 13 8 15 9 15 1 10 9 4 4 2
11 3 13 10 0 9 10 9 1 10 9 2
17 3 13 15 10 9 1 9 15 15 9 13 1 9 7 0 9 2
26 3 13 15 15 15 13 9 1 4 2 7 9 7 13 0 4 2 13 1 10 9 1 10 0 9 2
12 15 9 13 1 10 0 9 1 10 9 11 2
13 15 9 13 10 9 1 10 9 3 1 10 9 2
16 15 9 1 8 1 12 13 10 9 15 13 1 12 0 9 2
12 3 13 15 10 9 15 1 11 0 4 4 2
7 15 0 9 4 0 8 2
11 15 0 9 4 4 1 8 1 10 9 2
22 10 9 1 10 9 7 10 9 4 1 10 9 11 2 15 4 15 9 1 10 9 2
6 15 9 13 10 9 2
23 3 13 10 9 1 10 9 10 9 1 10 9 1 10 9 2 1 10 9 1 10 9 2
12 3 13 15 10 9 16 1 13 9 1 4 2
17 3 13 15 1 10 9 10 13 9 3 10 0 9 10 9 13 2
13 15 9 13 10 0 9 3 2 1 9 1 11 2
12 1 15 9 1 10 9 4 10 13 9 4 2
16 1 15 9 13 9 1 15 9 12 9 1 10 0 9 4 2
10 3 4 10 0 9 1 10 9 11 2
6 3 13 10 9 11 2
14 15 9 13 3 1 8 10 9 1 15 3 0 13 2
16 13 10 13 9 2 2 10 9 13 10 9 1 15 9 2 2
10 15 9 4 10 0 9 1 10 9 2
11 3 13 9 0 10 9 15 0 13 4 2
13 3 13 15 10 9 15 1 13 9 10 9 13 2
11 3 13 15 9 15 0 1 10 9 13 2
8 1 15 9 4 11 10 9 2
8 15 4 10 0 9 1 9 2
15 1 15 9 1 11 13 8 10 9 8 10 9 1 9 2
11 15 9 1 11 13 10 0 9 1 9 2
14 10 9 1 15 0 9 13 0 2 10 0 9 2 2
14 15 4 3 9 10 9 1 10 0 9 11 11 2 2
14 13 10 15 9 1 10 9 2 10 9 1 10 9 2
14 3 13 15 15 4 4 1 10 9 1 9 7 9 2
8 3 13 9 10 9 1 9 2
15 3 13 15 10 13 9 1 10 15 9 2 15 15 13 2
17 3 13 15 9 15 4 4 1 0 9 9 7 0 3 15 9 2
13 15 0 9 13 1 12 1 10 9 1 15 8 2
6 3 0 13 15 13 2
11 3 13 10 0 9 1 10 0 9 11 2
16 15 0 9 13 1 10 9 3 9 10 1 10 0 9 4 2
11 15 9 4 3 4 1 8 2 11 2 2
16 1 15 9 4 8 4 16 15 1 10 9 8 8 4 4 2
9 1 15 9 4 10 9 8 4 2
13 15 9 13 10 9 1 11 7 4 1 12 4 2
8 3 13 9 10 9 1 11 2
23 3 13 15 10 9 15 10 9 1 15 9 13 1 10 0 9 2 3 15 13 9 13 2
20 3 13 10 0 9 4 3 10 9 7 15 12 9 4 4 1 12 0 9 2
7 3 4 10 9 1 11 2
21 15 9 1 9 2 9 7 9 4 4 1 9 7 4 1 10 0 9 8 4 2
5 15 9 13 8 2
16 15 9 4 1 10 0 9 0 1 9 7 3 12 13 9 2
13 15 0 9 4 2 10 0 9 1 11 2 4 2
11 1 15 11 4 10 9 2 2 8 2 2
19 3 4 10 9 3 10 9 7 10 9 1 10 9 1 0 9 4 4 2
7 15 9 13 8 0 4 2
6 3 13 4 9 3 2
13 3 13 15 10 9 15 0 4 1 10 0 9 2
10 3 13 10 9 1 10 9 3 4 2
8 15 12 0 9 13 15 8 2
10 15 13 10 0 9 8 1 12 3 2
8 15 9 4 0 4 1 8 2
18 1 12 4 12 9 4 16 0 9 2 8 2 8 2 8 7 2 2
25 15 9 9 2 15 1 10 9 11 1 10 0 9 13 4 4 2 13 3 3 12 0 1 3 2
14 15 4 10 9 1 10 9 15 9 1 15 8 4 2
9 15 9 13 10 0 9 1 8 2
10 3 13 10 0 8 1 12 10 9 2
8 3 13 10 9 10 0 9 2
15 3 13 15 10 9 1 9 7 9 13 1 10 13 9 2
12 3 13 10 0 9 4 15 10 13 9 13 2
7 1 15 9 13 10 9 2
12 15 0 9 1 10 9 4 0 1 15 9 2
16 15 4 1 12 10 9 13 9 1 15 8 2 11 7 11 2
22 15 9 4 10 0 15 4 4 1 15 1 9 3 1 10 0 13 9 2 15 8 2
12 15 9 13 1 12 15 9 1 10 9 8 2
8 1 15 9 13 8 12 9 2
11 15 4 10 0 9 3 4 4 1 9 2
11 1 15 0 9 4 10 9 11 8 2 2
16 3 13 15 4 10 9 16 10 9 13 15 3 10 9 13 2
11 3 13 15 10 9 16 15 3 1 4 2
21 3 4 10 0 9 4 2 13 1 12 9 9 2 1 10 9 1 10 9 13 2
8 15 4 10 0 9 1 8 2
7 13 10 15 9 1 9 2
24 3 13 10 9 1 12 2 1 10 0 9 8 2 3 9 2 7 3 9 10 0 9 13 2
14 3 13 15 10 0 9 0 2 16 9 13 7 13 2
11 1 15 9 4 10 9 8 1 12 4 2
13 15 4 3 9 1 10 11 7 0 1 15 8 2
9 1 15 9 4 10 0 9 4 2
20 3 13 10 9 1 10 9 7 9 16 10 0 9 7 10 0 0 9 13 2
11 3 13 15 10 0 9 1 8 16 9 2
13 3 13 15 10 9 1 10 1 0 9 13 9 2
24 3 4 10 9 4 2 13 1 10 9 2 3 10 0 9 1 10 9 1 10 9 4 4 2
5 15 13 10 9 2
12 3 13 9 10 0 3 13 9 1 10 9 2
14 3 13 10 9 1 8 1 12 1 10 0 0 9 2
14 15 11 13 2 0 13 2 10 0 9 1 10 9 2
13 15 4 1 12 4 1 9 1 10 9 1 11 2
13 15 4 10 9 1 10 9 1 10 0 9 8 2
14 15 0 9 13 10 9 1 10 0 9 1 15 9 2
8 3 4 10 9 3 3 4 2
22 3 13 15 10 9 13 1 9 7 9 2 3 1 10 9 2 7 9 2 9 13 2
18 3 13 15 10 9 15 13 9 7 13 13 7 4 4 1 0 9 2
21 3 4 10 9 4 1 9 15 9 2 3 1 15 9 1 15 13 1 10 9 2
7 15 9 13 1 15 8 2
17 15 0 9 13 1 12 10 9 7 13 9 7 9 1 0 9 2
9 1 15 9 1 8 13 8 3 2
17 15 0 9 4 4 1 10 9 3 15 1 10 0 9 4 4 2
12 15 0 9 4 0 1 10 9 1 0 9 2
8 1 15 9 13 8 10 9 2
7 15 9 4 4 1 8 2
17 3 4 0 4 15 4 4 8 0 9 15 15 9 13 1 9 2
5 15 13 10 9 2
19 3 13 15 10 9 1 0 9 2 3 1 10 11 0 9 4 1 4 2
12 3 13 15 10 0 9 1 10 0 9 9 2
14 3 4 10 0 0 7 0 9 1 9 3 3 4 2
9 15 9 13 15 1 11 1 11 2
10 15 9 13 15 9 1 15 9 8 2
9 1 15 9 13 8 16 1 12 2
22 15 0 9 4 0 1 13 9 1 10 9 2 15 10 0 0 9 13 2 7 9 2
14 15 0 9 4 4 1 12 1 10 9 1 12 9 2
18 15 9 13 1 10 9 2 2 1 10 9 4 3 3 15 9 2 2
12 1 15 9 4 11 2 10 0 9 2 4 2
4 15 13 8 2
20 3 13 15 10 9 16 15 9 7 9 1 10 9 0 4 4 7 0 4 2
18 3 13 15 10 13 9 1 10 9 2 15 13 1 10 9 7 9 2
16 3 4 10 9 1 13 7 0 9 4 2 13 1 10 9 2
13 3 4 10 0 9 1 10 9 1 10 9 4 2
9 15 4 10 0 9 1 10 9 2
12 1 15 9 13 8 10 11 1 10 0 9 2
11 15 0 9 13 1 11 2 11 7 11 2
15 15 0 9 13 15 9 3 1 13 16 11 4 4 4 2
12 1 15 9 13 10 9 1 10 9 8 4 2
8 3 10 9 2 2 8 2 2
19 3 13 10 0 9 7 9 15 9 1 10 9 11 8 2 1 12 4 2
22 3 13 15 10 9 7 9 15 1 13 9 13 7 10 9 1 9 7 9 13 4 2
9 3 13 15 10 9 15 9 13 2
20 3 4 10 0 9 4 3 15 9 10 0 9 13 3 3 10 9 3 13 2
17 15 4 10 0 9 1 0 9 3 10 9 1 10 0 9 13 2
15 15 13 15 0 1 10 9 7 13 3 9 9 7 9 2
8 3 13 11 2 11 7 11 2
15 15 9 1 9 4 0 1 9 16 8 2 8 7 8 2
13 15 0 11 4 10 9 1 10 0 9 1 11 2
11 1 15 0 9 4 8 3 10 0 9 2
14 3 4 10 9 3 9 4 4 1 10 0 0 9 2
4 15 4 0 2
11 3 13 15 10 9 1 10 8 13 9 2
11 3 13 15 10 0 9 15 15 0 13 2
17 3 4 1 10 0 9 10 0 9 1 10 9 7 10 9 4 2
11 3 13 10 9 1 10 9 7 9 4 2
7 1 15 9 4 9 4 2
13 1 15 9 1 8 13 10 9 11 8 2 3 2
11 1 15 9 13 10 9 1 10 9 9 2
12 15 4 1 12 10 0 9 1 15 0 8 2
11 15 9 13 10 9 1 10 0 9 8 2
8 1 15 9 13 10 9 11 2
6 3 13 10 0 9 2
13 3 13 15 10 9 1 10 9 1 9 7 9 2
20 3 13 15 10 9 1 10 9 15 13 13 7 15 4 4 1 9 7 9 2
12 1 15 0 9 13 8 7 15 9 10 0 2
7 3 13 10 9 11 3 2
8 15 13 1 12 10 9 8 2
13 1 15 9 13 10 13 9 3 2 2 8 2 2
27 3 13 10 9 10 0 2 0 9 1 10 9 1 10 9 2 16 10 9 1 10 9 1 10 9 13 2
13 15 9 1 10 9 4 1 12 4 1 15 8 2
22 15 4 10 0 9 15 9 4 4 1 8 2 15 15 12 4 2 8 2 8 2 8
9 15 9 13 13 1 9 1 9 2
7 8 9 9 4 10 9 2
13 3 13 15 10 1 0 2 0 9 1 10 9 2
8 3 13 15 10 9 1 11 2
11 1 15 9 13 15 4 1 10 9 11 2
8 15 9 13 10 9 1 11 2
13 15 9 13 10 9 16 10 9 1 9 1 13 2
9 15 4 10 0 0 9 1 8 2
11 15 9 8 9 4 4 1 10 9 8 2
11 15 0 0 9 4 1 10 9 11 4 2
17 15 0 9 13 2 10 11 1 4 1 10 0 1 15 9 2 2
12 1 15 9 1 15 9 13 8 15 0 11 2
7 8 9 9 4 10 9 2
15 3 13 15 9 7 9 1 10 0 9 1 10 9 9 2
11 3 13 15 10 9 1 10 0 9 11 2
14 1 15 9 1 8 13 15 1 10 9 1 12 9 2
18 3 13 10 9 4 3 15 9 1 13 9 7 10 0 9 9 13 2
12 15 9 13 1 10 0 9 1 9 1 9 2
13 1 15 9 13 8 7 8 10 9 1 0 9 2
15 3 13 15 15 9 1 15 0 9 1 9 7 15 9 2
15 1 15 9 1 10 9 1 8 4 0 4 1 15 8 2
15 3 13 10 9 1 10 9 10 9 15 9 1 4 13 2
17 15 13 2 0 0 7 1 9 2 0 9 1 10 9 1 12 2
7 1 15 0 9 13 13 2
7 3 13 15 3 10 9 2
11 3 13 15 10 0 9 1 9 7 9 2
9 1 15 9 4 10 9 11 0 2
16 3 4 10 9 16 10 1 10 9 13 9 0 1 4 4 2
9 1 15 9 4 10 9 8 0 2
9 15 4 10 0 9 15 8 13 2
9 15 4 10 0 9 1 10 9 2
16 15 0 9 13 10 0 7 0 1 10 12 9 1 11 4 2
9 3 13 10 9 1 10 9 8 2
11 1 15 9 13 10 9 1 9 1 11 2
15 15 9 2 15 3 13 4 2 4 3 1 11 1 4 2
7 3 13 15 3 0 9 2
11 3 13 15 10 9 13 9 1 10 9 2
11 1 15 9 13 8 15 3 0 9 4 2
10 1 15 9 13 10 9 11 7 9 2
18 3 13 15 10 9 1 10 9 1 10 9 3 10 9 8 4 4 2
10 8 13 3 13 11 2 1 15 9 2
12 1 15 9 4 8 2 8 7 8 0 13 2
19 15 9 4 1 10 9 1 11 4 3 1 12 1 15 9 9 4 4 2
17 1 15 9 4 10 9 4 3 15 9 13 1 15 8 1 11 2
9 15 4 1 10 9 9 1 11 2
6 8 9 4 15 8 2
7 3 13 15 10 13 9 2
14 3 13 15 10 9 1 10 9 1 9 7 9 3 2
14 1 15 9 13 10 9 1 11 3 15 0 9 13 2
6 10 9 13 10 9 2
11 15 9 4 10 9 1 10 9 1 8 2
9 3 13 10 0 9 1 15 8 2
11 1 15 0 9 4 15 8 1 12 4 2
10 1 15 9 13 1 12 10 11 9 2
15 1 15 0 9 13 11 2 8 2 7 11 2 8 2 2
8 15 9 13 10 0 9 8 2
25 15 9 13 1 10 9 10 0 9 3 2 3 10 9 0 1 10 9 13 7 3 1 10 9 1
18 15 4 10 0 9 1 15 8 2 10 0 9 15 3 15 9 13 2
19 3 13 15 10 15 9 1 10 9 7 10 9 1 10 9 1 10 9 2
16 3 13 15 10 15 16 3 0 4 16 15 3 1 4 13 2
9 1 15 9 4 10 9 3 4 2
15 15 9 4 1 12 4 1 8 2 1 0 9 1 9 2
14 15 9 9 1 9 7 9 4 1 10 9 11 4 2
8 1 15 9 13 8 16 9 2
23 15 9 4 4 1 10 9 9 1 7 9 1 15 9 7 1 12 0 7 12 0 9 2
11 15 9 4 1 10 11 11 4 1 9 2
10 15 0 9 13 1 11 1 10 9 2
7 13 10 15 9 1 9 2
15 15 9 13 15 9 10 9 1 10 9 3 16 1 13 2
16 3 13 15 10 1 10 9 13 9 1 10 9 1 10 9 2
13 3 13 15 10 3 13 9 1 0 2 0 9 2
9 1 15 9 4 10 9 8 0 2
19 3 4 10 0 9 15 1 10 0 9 10 0 9 1 9 1 13 4 2
8 15 13 1 12 15 0 8 2
11 1 15 9 1 11 13 10 9 11 3 2
14 1 15 9 4 15 10 9 16 12 9 1 13 4 2
12 15 13 1 10 13 9 13 1 8 7 8 2
11 15 0 9 13 15 9 1 10 9 9 2
9 6 2 13 9 2 12 9 2 2
10 15 9 13 15 9 16 10 13 9 2
16 3 13 15 10 9 13 13 9 2 15 4 4 1 10 9 2
10 3 13 15 10 3 13 9 7 9 2
9 1 15 9 4 8 0 1 12 2
9 1 10 9 13 10 0 0 9 2
17 15 0 9 13 3 1 10 0 9 1 11 16 10 9 3 4 2
23 10 9 8 13 10 9 1 12 1 10 9 11 8 2 2 1 15 9 4 15 9 4 2
18 3 13 10 0 9 1 10 9 1 10 0 11 15 4 4 1 9 2
16 15 0 9 4 3 4 1 8 16 15 1 15 8 4 4 2
20 15 9 4 8 15 9 1 8 2 8 2 4 2 10 9 1 15 0 9 2
8 3 13 10 0 9 1 11 2
18 15 9 4 1 10 9 1 11 4 7 1 10 9 2 8 2 4 2
20 3 13 15 10 9 1 10 0 9 3 10 9 7 10 9 10 15 9 13 2
14 3 13 15 10 9 1 10 0 9 3 10 9 13 2
10 1 15 0 9 13 15 15 11 4 2
12 15 0 9 13 15 9 1 10 3 0 9 2
10 15 9 13 10 9 1 10 0 9 2
11 1 15 0 9 4 10 9 1 9 4 2
8 1 15 9 13 10 9 8 2
19 15 9 9 10 12 9 11 2 11 2 11 2 11 7 11 1 10 11 2
7 15 0 9 4 0 8 2
8 1 15 9 13 10 9 11 2
10 15 0 9 13 15 9 16 10 9 2
12 3 13 15 10 9 15 4 4 1 10 9 2
12 3 13 15 10 9 15 1 10 9 4 4 2
15 1 15 0 9 13 3 1 10 0 9 8 10 9 9 2
12 15 9 13 3 1 10 9 1 10 9 11 2
9 15 9 13 1 12 10 9 3 2
10 15 9 4 1 9 0 4 1 8 2
7 1 15 9 13 15 9 2
15 15 0 9 4 4 1 11 1 10 9 1 8 1 12 2
8 15 13 1 12 10 0 9 2
15 3 13 10 9 4 16 3 1 9 7 13 10 9 13 2
14 11 9 13 15 1 10 9 1 10 9 3 1 9 2
14 3 13 15 10 9 1 10 9 16 9 1 13 13 2
16 3 13 15 10 9 1 10 9 1 9 1 9 1 13 4 2
17 1 15 0 9 13 10 0 9 1 9 8 2 1 8 15 3 2
11 1 15 9 4 10 9 1 10 11 4 2
17 15 0 0 9 13 1 12 1 11 1 10 0 9 1 10 9 2
13 1 15 9 13 10 9 8 9 12 1 15 8 2
16 1 15 9 13 9 15 9 7 9 1 15 13 1 10 9 2
15 15 0 9 13 15 9 1 10 9 1 11 1 12 9 2
21 15 9 1 8 4 16 9 1 15 9 1 10 9 4 1 10 9 1 10 9 12
15 1 15 9 4 13 1 10 9 8 1 10 9 1 8 2
8 1 15 9 13 9 7 9 2
13 3 13 15 10 9 1 10 9 16 15 9 13 2
9 3 13 15 10 0 9 1 9 2
12 1 15 0 9 13 15 15 8 1 11 4 2
16 15 9 13 1 10 9 2 2 3 13 10 9 1 11 2 2
8 15 9 13 3 1 0 9 2
12 1 15 9 4 15 0 8 3 0 1 12 2
19 10 9 7 9 1 10 0 11 4 3 0 2 9 4 3 3 4 16 2
12 15 11 13 0 16 10 0 9 1 10 9 2
13 1 15 9 4 9 8 13 16 15 1 12 13 2
10 15 0 9 4 1 12 1 11 13 2
21 15 9 13 15 3 3 1 9 4 7 13 15 9 1 10 9 15 15 9 13 2
19 3 13 15 15 1 0 9 13 1 2 9 2 15 0 3 4 13 4 2
12 3 13 15 10 9 7 9 1 9 7 9 2
12 1 15 9 13 10 0 9 8 10 0 9 2
20 15 0 9 0 15 0 9 1 10 9 2 2 3 13 15 15 12 3 2 2
9 15 9 1 10 9 13 10 9 2
9 15 9 4 10 0 9 1 8 2
8 1 15 9 13 8 10 9 2
11 15 4 10 9 1 10 0 9 1 11 2
13 1 15 9 13 10 9 11 1 12 10 9 3 2
9 1 15 9 13 10 11 11 3 2
20 1 10 9 1 15 8 13 15 0 9 2 15 4 10 0 9 1 15 9 2
18 3 13 15 15 13 1 9 1 10 15 9 1 10 9 1 10 15 2
11 3 13 15 10 9 15 1 10 9 13 2
9 1 15 9 13 15 15 11 4 2
10 1 15 9 13 15 1 11 4 4 2
11 1 15 9 13 8 10 0 9 1 9 2
22 1 12 13 10 9 8 10 9 1 10 9 1 10 15 9 1 10 9 2 15 9 2
19 15 4 10 9 1 10 0 9 8 15 12 9 10 9 1 15 8 13 2
15 15 4 10 9 1 10 0 9 11 16 9 1 15 8 2
11 15 9 13 1 12 10 0 9 1 8 2
11 1 15 9 4 0 16 15 10 9 13 2
13 15 9 13 1 10 9 1 10 9 7 10 15 2
12 3 13 15 10 9 1 10 9 1 10 9 2
10 3 13 15 10 13 9 1 0 9 2
15 1 15 9 13 10 11 2 15 4 4 1 10 0 9 2
7 15 9 4 1 12 0 2
9 15 9 13 8 1 4 1 9 2
10 1 15 9 13 8 10 9 1 8 2
11 15 9 13 10 10 9 1 10 9 12 2
12 15 9 1 10 11 4 1 12 4 1 11 2
21 1 15 0 9 13 8 1 12 10 0 9 1 10 9 1 10 9 1 10 9 2
9 15 9 13 10 9 11 12 2 2
9 15 9 13 10 9 1 10 9 2
10 15 9 4 10 9 16 15 15 13 2
8 3 13 15 0 9 7 9 2
17 3 13 15 10 9 1 12 9 2 3 10 9 15 10 9 13 2
14 1 15 9 13 10 11 2 10 9 1 10 0 9 2
9 15 9 13 15 1 11 1 9 2
10 1 15 9 4 10 9 1 9 4 2
14 15 0 9 15 1 12 13 4 1 8 7 8 4 2
9 15 4 7 9 13 16 9 12 2
13 15 13 15 9 8 2 1 10 9 1 15 8 2
15 15 0 9 13 1 12 1 15 9 1 15 8 1 11 2
17 13 10 15 9 1 15 9 8 2 2 10 0 9 1 15 8 2
9 3 13 15 15 0 1 10 9 2
18 3 13 15 15 15 8 15 9 0 9 13 4 7 15 9 13 4 2
9 3 13 15 10 9 1 0 9 2
7 1 15 9 13 10 11 2
12 15 13 10 0 9 1 10 0 9 1 12 2
7 15 9 13 0 0 9 2
13 1 10 9 9 8 7 11 1 9 10 9 0 2
6 15 9 13 15 9 2
10 15 13 1 12 10 9 1 10 9 2
6 1 15 9 13 8 2
9 9 2 0 13 2 12 9 2 2
14 3 13 10 0 9 3 11 13 7 15 9 0 13 2
22 3 13 15 1 10 0 9 10 0 9 1 9 15 13 1 15 0 13 1 11 9 2
12 3 13 15 10 9 15 1 13 10 9 13 2
8 1 15 9 13 10 9 8 2
13 15 4 10 9 1 10 9 1 10 0 9 11 2
10 1 15 9 13 15 10 9 1 11 2
13 1 15 9 13 10 9 8 8 1 10 0 9 2
16 8 4 10 0 9 1 0 9 2 3 3 4 15 2 4 2
9 1 15 9 4 8 1 12 4 2
15 3 4 10 0 1 8 1 15 15 3 1 15 9 13 2
19 3 4 10 9 15 15 1 10 9 1 10 0 9 13 1 15 13 8 2
13 1 15 9 1 9 4 10 0 7 0 9 4 2
17 3 13 15 1 10 9 10 0 9 1 15 9 2 9 7 9 2
17 3 13 15 10 0 9 2 15 1 10 0 9 1 10 9 13 2
9 1 15 9 4 10 9 8 0 2
10 15 0 9 4 1 12 4 1 8 2
8 15 9 13 1 12 10 9 2
14 15 4 10 0 9 1 8 2 13 1 9 13 9 2
7 15 9 13 8 1 12 2
11 15 9 4 1 12 4 1 8 7 8 2
14 15 4 1 12 1 10 9 11 10 0 9 1 9 2
10 1 15 9 13 10 11 7 15 8 2
11 15 9 13 10 9 1 10 10 13 9 2
9 3 13 15 1 0 0 10 9 2
20 3 13 15 10 3 13 9 15 4 4 1 10 9 15 10 9 4 1 8 2
10 1 15 9 4 10 9 1 11 4 2
12 1 15 9 13 10 9 1 11 1 12 0 2
11 3 4 10 9 1 10 9 7 10 9 2
10 15 9 1 11 4 4 16 0 9 2
24 3 4 10 0 9 11 4 2 15 8 12 5 1 10 9 1 15 8 13 2 7 3 3 2
15 15 0 9 7 9 13 16 0 1 10 9 1 10 9 2
23 15 0 9 13 3 1 9 1 9 2 2 9 4 3 0 9 16 15 15 9 13 2 2
10 3 4 10 0 0 15 3 9 13 2
19 10 9 1 10 9 9 1 15 8 2 15 4 10 0 9 1 15 9 2
23 3 13 15 1 10 0 10 9 3 1 10 9 13 9 0 4 4 1 9 1 10 9 2
13 3 13 15 10 9 9 1 10 9 1 10 9 2
8 1 15 9 13 15 9 0 2
12 3 4 10 9 1 11 15 1 12 4 4 2
9 15 0 9 13 10 9 1 9 2
14 3 13 10 9 16 1 9 10 15 9 3 1 4 2
27 15 4 10 9 1 10 0 9 1 12 1 10 9 2 8 2 15 1 9 3 1 0 9 0 13 4 2
11 15 4 1 12 10 9 1 10 0 9 2
13 1 15 9 13 15 10 9 1 10 0 9 8 2
15 15 0 9 1 8 13 1 12 10 11 1 0 0 9 2
4 11 2 0 0
15 3 13 15 0 9 2 3 15 13 10 9 1 15 4 2
17 3 13 15 10 0 3 0 9 2 3 10 0 9 3 13 4 2
13 1 15 0 9 13 10 9 1 8 1 10 9 2
10 1 10 9 1 15 9 13 10 11 2
14 13 4 4 16 9 1 9 2 15 4 10 13 9 2
12 1 15 9 4 13 7 9 1 13 9 4 2
21 15 4 10 9 1 10 0 9 8 2 15 12 5 0 7 12 5 9 13 4 2
10 15 4 10 0 9 1 11 1 12 2
11 3 13 10 0 9 1 10 0 9 11 2
9 1 10 9 13 10 9 1 13 2
16 15 9 1 0 9 4 3 1 10 9 0 1 10 0 9 2
18 3 13 15 9 15 13 1 9 1 4 2 1 4 2 7 1 4 2
13 3 13 15 10 9 3 15 13 4 4 7 4 2
7 1 15 9 13 8 3 2
16 15 9 13 10 9 1 10 12 0 9 1 10 0 9 3 2
13 0 13 15 1 10 9 2 1 15 9 13 15 2
21 2 16 15 1 15 13 2 13 15 3 1 15 3 2 4 0 1 10 9 3 2
9 15 4 10 12 9 1 10 9 2
28 15 0 9 13 15 1 9 16 9 11 2 2 11 11 2 2 11 11 2 2 11 11 2 7 9 11 2 2
19 15 0 9 4 4 1 10 9 1 10 9 1 10 9 1 10 9 11 2
8 1 15 9 13 10 0 9 2
10 15 4 10 12 0 9 1 10 9 2
14 3 13 15 9 7 9 1 9 2 3 13 1 9 2
14 3 13 15 10 9 2 13 1 10 13 7 0 9 2
14 1 15 0 9 13 15 10 9 11 11 2 1 8 2
9 1 15 9 4 10 9 11 4 2
9 3 13 15 10 9 1 10 9 2
14 1 15 4 8 10 9 3 1 10 9 11 11 2 2
17 1 15 9 2 15 1 10 9 13 2 13 10 0 9 15 9 2
11 1 15 9 13 10 0 9 8 10 9 2
8 15 4 1 12 9 1 11 2
14 15 0 9 13 1 15 9 1 12 10 0 9 3 2
15 1 15 9 4 3 1 9 10 9 4 1 9 7 9 2
23 3 13 15 13 1 10 9 1 10 9 2 15 15 1 10 9 13 4 1 10 0 9 2
21 3 13 15 10 1 9 2 9 2 9 2 3 2 7 9 2 13 9 7 9 2
13 1 15 0 9 4 10 9 0 7 0 9 4 2
10 3 13 10 0 9 1 10 9 11 2
12 3 4 10 9 3 8 10 9 4 1 4 2
13 3 13 15 10 9 1 8 12 13 1 15 9 2
19 1 15 13 11 9 4 1 15 0 9 1 11 1 10 11 9 1 12 2
10 15 9 4 3 4 16 2 8 2 2
12 15 9 4 3 16 15 9 11 10 13 9 2
3 10 0 9
3 10 0 9
9 3 13 15 1 10 9 3 4 4
7 15 13 15 13 1 10 9
7 1 10 9 3 13 15 3
7 15 13 4 15 15 3 0
7 15 13 4 15 15 3 4
7 10 9 13 11 16 15 0
7 15 13 11 16 10 9 0
10 15 13 11 16 11 4 16 15 4 4
13 11 13 3 4 4 16 11 10 9 3 4 4 4
5 15 13 4 1 4
15 11 13 16 15 3 4 4 1 4 1 10 9 3 1 4
3 10 0 9
16 11 13 16 15 15 3 4 4 1 4 1 10 9 3 1 4
10 15 13 1 4 4 10 9 1 4 4
11 15 13 15 1 4 4 10 9 1 4 4
6 15 13 4 16 1 4
16 11 13 16 15 3 4 4 1 4 16 1 10 9 3 1 4
17 11 13 16 15 15 3 4 4 1 4 16 1 10 9 3 1 4
11 15 13 1 4 4 16 10 9 1 4 4
12 15 13 15 1 4 4 16 10 9 1 4 4
6 15 13 11 4 1 4
6 15 13 11 4 1 4
3 10 0 9
16 11 13 16 15 15 3 4 4 1 4 1 10 9 3 1 4
11 15 13 15 1 4 9 10 9 1 4 4
17 11 13 16 15 15 3 4 4 1 4 16 1 10 9 3 1 4
12 15 13 15 1 4 4 16 10 9 1 4 4
9 15 4 4 16 10 9 3 1 13
10 16 10 9 3 1 13 4 15 0 4
3 15 4 0
4 15 4 10 9
4 0 4 15 3
4 15 13 3 0
3 10 0 9
4 15 13 3 0
4 15 4 15 0
7 10 9 15 15 13 4 13
6 10 9 15 15 9 13
7 10 9 15 15 13 4 13
6 10 9 15 15 13 13
6 9 15 15 13 4 13
5 9 15 15 13 13
7 10 9 16 15 13 4 13
6 10 9 15 15 9 13
3 10 0 9
7 10 9 15 15 13 4 13
6 10 9 15 15 13 13
6 13 15 15 13 4 13
5 13 15 15 13 13
7 10 9 15 15 13 4 13
6 10 9 15 15 9 13
6 9 15 15 13 4 13
5 9 15 15 9 13
7 10 9 16 15 13 4 13
6 10 9 15 15 9 13
3 10 0 9
6 9 15 15 13 4 13
5 9 16 15 9 13
5 10 9 15 9 13
7 10 9 1 15 13 15 13
5 10 9 3 15 13
6 15 13 15 3 13 4
7 15 13 15 15 3 4 4
8 15 13 15 9 15 3 4 4
11 15 0 1 15 9 15 3 4 4 1 11
11 15 0 1 15 13 15 3 4 4 1 11
3 10 0 9
10 15 13 3 10 9 3 4 4 1 11
4 10 9 13 2
9 10 9 2 15 15 13 2 13 2
8 10 9 15 15 13 2 13 2
8 10 9 2 15 15 9 13 2
3 15 13 2
4 15 13 11 4
5 15 13 1 11 4
9 15 13 10 0 11 1 10 9 4
5 15 13 1 9 4
3 10 0 9
5 15 13 15 9 4
6 15 13 15 11 3 4
5 15 13 10 9 4
6 15 13 10 9 4 4
6 15 13 10 9 4 4
7 15 13 10 9 3 4 4
7 15 13 10 9 4 4 4
7 15 13 10 9 4 4 4
9 15 9 13 15 11 4 16 1 4
7 16 15 11 10 9 13 4
3 10 0 9
8 15 11 11 11 10 9 13 4
10 16 11 11 10 9 10 9 13 4 4
13 15 13 16 11 11 11 4 4 16 10 9 4 4
3 3 4 4
6 1 10 9 4 15 4
6 10 9 4 4 1 11
7 3 4 4 10 9 1 4
11 3 4 4 16 3 1 10 9 15 4 4
8 16 8 4 3 1 10 9 4
6 1 10 9 4 1 4
3 10 0 9
4 3 4 1 4
5 10 9 4 1 4
7 10 9 13 1 15 1 4
7 10 9 13 4 3 1 4
8 16 10 9 13 4 3 1 4
8 16 10 9 13 1 15 1 4
8 16 10 9 3 1 4 13 4
7 3 13 10 9 1 10 9
8 3 13 3 10 9 1 10 9
13 3 13 10 0 9 1 10 9 7 10 0 13 3
3 10 0 9
3 10 0 9
4 15 13 15 0
6 15 13 15 1 10 9
5 10 9 13 15 1
6 15 8 13 0 9 4
11 10 11 1 11 13 0 16 10 11 1 12
11 15 13 1 10 9 4 10 9 1 10 9
7 15 13 11 4 1 0 9
7 15 13 15 3 1 10 9
6 10 9 13 1 15 9
5 16 15 1 15 13
3 10 0 9
6 16 15 1 15 3 13
4 15 13 15 0
6 16 15 15 13 1 4
4 15 13 15 0
8 16 15 13 7 15 0 4 4
8 15 13 15 3 3 16 15 4
6 15 13 16 15 0 4
6 15 13 15 16 15 13
10 15 13 15 4 16 11 3 4 1 4
10 10 0 13 10 9 3 2 3 10 9
3 10 0 9
5 15 13 3 1 9
5 7 15 13 11 0
6 10 9 1 15 15 13
7 10 9 1 15 15 13 4
5 10 9 3 15 13
8 15 13 15 3 1 10 9 4
6 15 13 15 15 4 4
6 15 13 3 15 4 4
7 15 13 1 15 15 4 4
6 15 13 3 15 4 4
3 10 0 9
7 15 13 1 15 15 4 4
4 3 13 15 1
6 3 13 15 3 3 4
7 10 9 3 15 3 13 4
5 3 13 15 15 3
4 3 13 15 3
3 3 4 4
4 1 11 4 4
13 15 13 15 15 1 1 9 1 9 1 10 9 11
13 1 9 13 15 10 9 3 1 9 13 15 10 9
3 10 0 9
7 15 13 3 15 3 0 4
10 13 3 3 15 0 16 3 15 0 4
5 8 4 3 8 4
6 15 4 10 9 8 4
8 10 9 4 3 10 9 8 4
6 8 13 8 4 4 4
7 16 8 10 9 8 4 4
6 16 11 8 4 13 4
8 15 13 15 7 0 16 10 9
8 15 13 15 8 13 8 10 9
3 10 0 9
9 15 13 7 1 12 2 7 1 8
10 15 13 2 13 11 2 16 15 3 4
12 15 13 2 3 13 11 2 16 15 3 4 4
9 7 3 13 2 1 15 2 10 9
14 15 13 15 0 2 0 2 0 2 0 2 7 10 9
13 15 13 15 0 2 0 2 0 2 0 7 10 9
13 15 13 15 0 2 0 2 0 2 0 2 10 9
15 15 13 15 7 0 2 0 2 0 2 0 2 16 10 9
14 15 13 15 7 0 2 0 2 0 2 0 16 10 9
13 15 13 10 9 4 15 15 13 7 15 15 3 13
3 10 0 9
7 15 13 1 12 7 16 8
10 15 13 1 15 9 2 7 1 15 9
11 15 13 1 12 7 3 13 15 15 15 13
8 15 13 2 15 13 7 15 13
9 15 4 10 0 2 0 7 0 9
11 15 13 9 2 9 2 9 3 1 15 9
7 15 13 7 11 16 11 4
11 15 13 7 11 2 11 2 11 16 11 4
9 15 13 7 10 9 7 10 9 4
7 15 13 3 3 3 3 4
3 10 0 9
4 15 13 3 4
7 15 13 3 3 3 4 4
9 15 13 3 10 9 3 3 4 4
7 15 13 10 9 3 3 4
5 10 9 4 0 3
5 0 3 4 15 3
8 15 4 10 9 3 15 13 4
6 3 0 13 15 15 9
10 10 9 3 0 15 15 4 4 3 4
6 3 0 13 15 15 9
3 10 0 9
9 15 13 3 0 7 3 0 15 4
7 15 0 1 8 9 15 4
7 15 0 1 8 9 15 4
8 15 13 8 0 9 10 9 4
7 15 13 3 2 13 15 0
10 10 0 0 9 3 10 0 9 4 13
5 15 13 0 0 9
4 15 13 9 4
6 6 2 15 4 10 9
8 9 2 3 13 15 3 3 4
3 10 0 9
8 9 2 13 15 15 9 4 2
6 15 4 15 9 2 6
4 15 13 2 0
4 15 13 2 8
10 13 15 0 4 2 3 13 15 3 4
8 9 2 3 13 15 3 3 3
8 10 1 9 0 9 4 3 0
6 15 9 4 0 1 9
9 10 9 4 0 16 15 1 9 4
5 15 4 0 1 9
3 10 0 9
2 0 9
5 15 4 9 1 9
6 15 4 0 16 1 4
6 15 4 9 16 1 4
6 15 4 0 16 15 13
5 16 15 13 4 0
6 15 4 0 16 1 13
5 16 1 13 4 0
5 3 4 15 0 3
5 15 4 3 0 3
8 9 2 3 4 15 8 0 3
2 0 9
4 10 3 0 9
4 10 15 0 9
3 15 4 8
4 15 4 10 0
4 15 4 8 0
7 15 4 8 0 16 1 4
7 15 4 15 0 16 1 4
4 15 13 8 4
4 15 13 8 4
5 15 4 0 16 15
2 0 9
8 15 4 0 1 11 16 1 11
5 15 4 0 16 0
6 15 13 0 3 3 3
6 15 4 0 16 15 13
9 15 4 0 16 15 13 16 11 4
7 15 4 0 16 16 15 13
10 15 4 0 16 16 15 13 16 11 4
5 15 13 3 16 15
13 15 13 16 15 4 4 7 16 15 15 3 4 4
13 15 13 16 15 15 0 4 7 16 15 15 3 4
2 0 9
12 15 1 9 4 7 15 13 13 3 1 10 9
12 15 13 15 16 15 4 7 16 15 3 4 4
15 15 13 1 9 16 15 3 0 4 7 16 15 3 9 13
5 15 13 3 1 4
8 15 13 3 12 9 1 4 4
8 15 13 3 12 9 4 1 4
7 15 13 12 9 1 4 4
6 15 13 12 9 1 4
7 15 13 12 9 1 4 4
7 15 13 12 9 4 1 4
2 0 9
7 15 13 12 9 1 4 4
7 15 13 15 10 9 1 4
8 15 13 15 10 9 1 4 4
6 1 10 9 4 10 9
8 1 10 9 13 16 11 9 4
9 15 13 1 10 9 16 11 9 4
8 16 11 9 4 13 1 10 9
6 3 13 16 11 9 4
6 15 13 16 11 9 4
7 3 13 3 16 11 9 4
2 0 9
7 10 9 1 11 4 15 0
7 15 4 15 0 16 15 13
6 16 15 13 4 15 0
7 15 4 15 0 16 1 13
6 16 1 13 4 15 0
7 15 13 15 0 16 15 4
6 16 15 4 13 15 0
7 15 13 15 0 16 1 4
6 16 1 4 13 15 0
9 16 15 13 4 13 15 1 10 9
2 0 9
7 16 13 13 15 1 10 9
7 16 15 13 13 15 10 9
9 15 13 10 9 1 1 10 9 4
7 15 4 3 1 1 10 9
7 15 13 3 1 1 10 9
5 15 13 3 1 3
8 15 13 10 9 1 3 1 3
7 15 4 1 3 3 12 9
7 1 9 7 3 4 15 13
8 15 13 1 16 10 9 13 4
2 0 9
7 1 16 0 15 10 9 2
7 15 0 3 3 10 9 4
5 15 13 1 3 3
5 15 13 1 3 3
7 10 9 7 15 4 13 15
8 10 9 15 15 4 4 4 4
9 10 9 13 10 9 15 9 0 4
6 3 13 15 3 1 4
5 3 13 15 1 4
5 10 9 9 12 9
2 0 9
4 10 9 13 9
7 10 9 13 15 10 0 9
8 15 13 1 9 3 4 15 13
13 3 4 10 9 3 3 0 2 10 9 13 15 3
4 15 13 3 9
11 15 13 1 9 16 1 13 7 3 1 13
10 15 13 1 4 7 10 0 9 1 4
8 8 4 4 15 1 15 9 3
6 3 1 4 13 15 15
7 4 13 11 3 1 10 9
2 0 9
6 4 4 10 9 1 4
7 4 4 16 10 9 0 4
4 4 4 3 3
5 1 4 13 3 3
7 3 1 4 13 3 3 15
7 9 4 15 15 1 15 9
5 4 4 16 15 13
7 4 13 11 10 9 10 9
7 4 4 15 16 15 9 4
7 4 13 15 10 9 10 9
3 10 0 9
2 0 9
8 4 4 13 15 10 9 10 9
6 16 15 0 4 16 15
8 16 15 10 0 9 4 16 15
9 16 15 10 0 13 9 13 16 15
9 16 15 10 0 13 9 16 15 13
6 0 16 15 13 15 3
8 10 0 9 16 15 13 3 3
8 15 13 0 7 0 4 16 3
7 15 13 3 0 4 16 3
6 15 4 3 0 16 15
2 0 13
9 16 15 10 15 9 13 4 16 15
7 16 15 15 9 13 16 15
6 15 0 16 15 13 15
7 15 13 15 0 4 16 15
9 15 13 10 9 4 15 15 13 4
13 15 13 10 9 4 15 10 9 13 4 15 3 13
9 15 13 10 9 4 4 15 3 13
9 15 13 9 1 9 4 15 3 13
9 15 13 9 1 9 4 15 3 13
10 15 13 9 1 0 9 4 15 3 13
2 0 9
10 15 13 9 1 0 9 4 15 3 13
10 15 13 10 9 4 16 10 9 15 13
11 15 13 10 9 9 4 15 1 10 9 13
9 15 13 10 9 9 4 15 13 4
11 15 13 15 9 4 16 15 1 10 9 13
13 15 13 10 9 7 10 9 4 15 1 10 9 13
13 10 9 7 10 9 13 15 4 15 1 10 9 13
12 10 0 9 13 15 4 16 15 3 13 1 4
10 12 9 13 15 4 15 1 10 9 13
11 10 9 13 15 4 4 15 1 10 9 13
2 0 9
11 10 9 13 15 4 4 15 1 10 9 13
9 0 9 13 15 4 4 4 16 15
9 0 9 13 15 4 4 4 16 15
8 1 0 9 13 15 4 16 15
11 1 9 13 15 4 4 15 3 1 4 4
7 16 4 4 4 11 9 4
7 16 1 12 13 11 10 11
14 16 11 10 9 13 1 12 2 13 11 10 9 1 12
6 16 13 4 11 9 4
8 15 4 0 4 10 9 1 4
3 10 0 9
6 0 4 15 4 1 4
9 15 4 0 4 16 10 9 4 4
10 0 4 15 3 4 16 10 9 4 4
8 15 13 10 9 4 16 15 4
7 10 9 4 4 16 15 4
8 15 4 10 9 4 15 1 4
7 10 9 4 4 15 1 4
12 15 9 13 3 0 3 3 2 16 15 4 4
10 15 9 13 3 3 2 16 15 4 4
9 15 13 3 3 3 3 16 1 4
3 10 0 9
8 15 13 3 3 3 3 1 4
6 15 13 3 16 1 4
5 15 13 3 1 4
9 15 13 3 3 3 15 15 3 4
8 15 13 3 3 15 15 3 4
8 15 13 3 3 3 16 15 4
7 15 13 3 3 16 15 4
12 15 13 15 3 3 3 4 16 10 9 15 4
11 15 13 15 3 3 4 16 10 9 15 4
7 15 4 10 9 15 15 13
7 11 13 16 11 10 9 4
7 16 15 13 4 3 10 9
8 15 4 15 10 9 16 15 13
8 15 4 15 10 9 16 15 13
7 16 15 13 4 15 10 9
7 16 15 13 4 15 10 9
6 10 9 4 16 15 13
7 10 9 4 15 16 15 13
5 0 4 16 15 13
7 0 4 15 3 16 15 13
9 10 0 9 4 16 3 1 13 4
8 11 13 16 11 10 9 4 4
11 10 0 9 4 15 3 1 3 1 13 4
6 0 4 16 3 1 13
7 0 4 15 16 3 1 13
8 0 13 15 15 3 16 15 4
6 0 13 15 16 15 4
5 0 4 16 1 13
6 0 4 15 16 1 13
8 15 4 3 0 4 16 15 4
8 0 4 15 3 4 16 15 4
7 16 15 4 4 3 0 4
9 11 13 16 11 10 9 4 4 4
7 15 13 16 16 15 15 13
10 15 13 3 9 4 2 1 15 13 9
7 15 4 4 15 15 13 4
8 15 4 4 2 15 15 13 4
12 15 13 1 9 1 15 9 2 7 1 15 9
6 15 15 13 4 15 3
10 15 13 3 4 15 15 0 9 3 13
11 15 13 3 4 2 15 15 0 9 3 13
7 15 15 13 2 4 15 3
8 15 13 2 3 16 15 0 4
10 11 13 16 11 10 9 3 4 1 4
7 15 4 10 9 3 15 13
6 15 13 15 3 15 4
5 15 13 1 3 3
7 10 9 13 2 13 7 13
8 15 13 1 10 9 7 1 9
10 15 13 16 15 4 7 16 15 3 4
13 15 13 1 9 16 15 1 13 2 7 9 1 13
6 16 15 8 13 1 11
6 16 15 1 11 8 4
6 16 15 3 1 8 4
3 10 0 9
11 11 13 16 11 10 9 3 4 1 4 4
5 15 4 3 3 8
8 16 15 8 4 16 11 4 4
10 15 13 1 15 3 16 15 0 4 4
6 15 13 9 1 15 3
6 16 15 10 9 8 13
7 16 15 3 0 8 4 4
9 11 13 8 1 9 2 9 7 9
6 16 15 10 9 3 13
7 16 15 3 10 9 8 13
5 15 13 9 1 9
7 11 13 16 10 9 4 4
5 15 13 3 9 3
4 15 13 3 9
8 15 13 3 9 3 16 15 4
5 16 10 9 8 13
7 16 10 9 3 0 8 13
7 15 9 13 8 1 10 9
6 16 15 12 9 0 13
7 16 15 15 12 9 0 13
5 10 9 4 8 4
8 15 13 15 8 10 9 1 4
7 11 13 16 10 9 4 4
8 10 0 9 13 15 1 15 9
5 10 9 13 3 9
6 10 9 13 9 1 11
5 15 13 3 0 3
7 15 13 3 3 16 10 9
12 15 4 15 3 3 3 0 16 10 9 4 4
12 15 4 15 3 3 3 3 16 0 3 1 4
12 15 4 15 3 0 3 0 16 10 9 4 4
12 15 4 15 3 0 3 3 16 0 3 1 4
6 15 13 15 10 9 8
11 11 13 16 10 9 3 4 1 4 4 4
7 15 13 15 9 1 10 9
5 15 13 15 16 0
6 15 13 3 16 0 3
6 15 13 10 9 16 0
11 15 13 16 1 4 7 16 0 3 1 4
9 15 13 1 4 7 0 3 1 4
9 15 13 16 15 4 3 15 0 4
6 13 15 15 0 4 2
6 15 4 0 15 4 4
6 15 13 12 9 1 4
4 15 0 10 9
4 15 13 15 4
5 15 13 15 4 4
8 15 13 16 15 15 4 4 4
9 15 13 16 15 15 4 4 4 4
5 15 13 15 4 4
6 4 13 15 15 3 4
5 15 13 15 9 4
9 15 15 1 9 13 13 10 0 9
10 15 15 15 3 0 4 9 3 0 1
11 15 13 16 15 15 15 13 1 10 9 4
5 15 13 10 9 4
11 15 13 16 15 1 10 9 4 15 0 4
8 15 15 13 13 16 15 0 4
7 15 13 16 1 15 3 0
6 15 16 9 13 9 0
10 10 9 4 0 1 15 1 10 9 11
4 13 15 4 2
8 15 15 16 8 13 15 4 4
8 15 13 15 15 4 4 16 8
8 15 13 3 15 4 3 1 11
8 3 3 13 15 4 3 1 11
6 15 13 10 9 3 4
8 3 3 13 15 15 9 4 2
10 15 13 3 16 15 0 4 4 1 9
10 15 13 16 15 0 4 1 9 16 15
12 15 13 16 15 0 4 16 15 1 15 0 9
5 15 4 10 9 0
12 15 13 15 3 0 0 4 16 15 3 3 4
12 15 13 15 0 4 16 3 15 9 3 1 4
5 15 13 15 16 3
11 11 13 3 0 4 16 15 1 10 9 13
10 11 13 15 4 16 15 1 10 9 13
7 15 13 10 9 3 4 4
10 10 9 4 15 16 15 1 10 9 13
7 11 13 10 9 4 16 11
7 11 13 15 0 4 16 11
7 3 13 15 3 10 9 1
8 3 4 15 3 9 3 1 4
9 10 9 13 15 3 16 15 0 4
6 15 13 10 9 15 4
7 3 13 3 10 9 3 1
8 3 13 3 10 9 3 1 4
7 15 13 10 9 1 15 4
7 15 13 10 9 3 4 4
7 15 13 15 1 9 1 15
7 10 9 9 13 16 10 9
5 15 13 10 9 4
5 15 4 10 9 0
6 15 4 10 0 9 0
7 0 10 0 9 4 15 0
6 10 9 13 16 3 4
9 10 9 1 15 13 3 10 9 4
4 10 9 13 3
6 15 13 10 9 3 4
4 10 9 13 15
4 15 13 15 3
7 0 13 15 15 9 3 0
6 15 4 10 9 1 4
5 15 13 10 9 3
6 15 13 10 9 3 1
8 11 13 10 9 10 9 3 4
7 3 13 11 15 10 9 3
9 15 13 1 9 3 16 15 0 4
9 15 13 1 9 1 15 3 3 13
6 15 4 3 10 9 8
3 10 0 9
5 10 9 13 15 4
12 15 8 13 12 9 1 3 10 9 1 15 9
6 15 13 15 16 15 4
6 7 15 4 13 15 8
7 15 4 3 4 16 15 4
6 7 15 4 4 3 4
3 15 4 9
5 9 4 15 0 2
11 15 4 1 10 0 9 16 15 9 13 4
7 15 4 1 11 16 15 13
6 15 4 9 15 15 13
6 10 9 13 15 3 4
8 15 4 15 9 15 15 4 13
6 15 4 0 15 15 13
7 15 4 9 15 15 3 13
7 15 13 15 0 16 15 4
6 7 15 4 13 15 0
8 15 4 3 0 3 16 15 4
9 15 4 3 0 1 15 1 4 4
11 15 13 15 3 0 1 10 9 0 1 4
10 15 4 3 1 15 16 10 9 1 13
6 16 15 10 9 4 13
7 10 9 13 15 3 4 4
7 16 15 10 9 3 4 13
8 16 15 10 9 3 3 4 13
4 10 1 13 9
4 10 1 13 9
4 10 1 13 9
10 10 9 15 9 4 4 4 1 10 9
7 15 13 9 13 9 1 11
7 15 13 9 8 10 9 4
11 15 13 3 15 3 4 16 15 3 13 4
5 10 3 1 13 9
7 10 9 13 15 3 4 4
6 16 15 4 13 4 15
5 1 3 4 4 15
4 1 13 4 15
9 16 15 15 9 3 1 10 9 13
8 16 15 1 10 9 15 9 13
7 16 15 15 3 1 9 13
9 16 15 1 9 10 0 9 13 4
7 16 15 1 15 10 9 13
8 16 15 10 9 3 1 15 13
6 16 15 15 10 9 13
5 3 13 15 10 9
7 16 15 10 9 10 9 13
8 3 3 10 9 4 4 15 9
6 3 16 15 0 13 15
11 3 3 3 10 9 15 13 4 4 9 4
7 3 1 11 4 4 1 8
8 15 13 3 4 3 10 9 4
7 15 13 4 3 10 9 4
9 15 4 1 11 4 3 15 3 13
9 15 13 10 0 4 15 10 9 13
6 1 11 0 4 15 0
6 3 13 15 10 9 4
7 1 11 10 9 4 15 0
6 1 0 3 10 0 9
8 15 13 10 9 1 3 10 9
10 1 0 9 1 13 13 15 9 12 9
6 15 13 3 15 15 4
10 15 13 1 3 10 9 15 10 9 4
5 3 4 10 9 2
10 15 13 15 3 3 15 10 9 4 2
8 15 13 15 4 16 15 9 2
7 16 15 9 13 15 4 2
7 3 13 15 10 9 3 4
7 15 13 7 13 10 0 9
7 15 13 7 13 10 9 4
6 15 13 15 4 7 4
6 15 13 15 4 7 4
8 15 13 15 4 4 7 4 4
6 16 15 4 7 4 4
7 16 15 1 4 7 4 4
6 16 15 4 7 4 4
8 15 4 12 9 3 16 15 13
9 16 15 15 9 13 4 12 9 3
8 3 13 15 10 9 3 4 4
6 15 13 10 9 3 15
8 15 13 12 10 9 15 12 15
8 15 13 8 16 10 9 1 13
9 15 13 3 3 8 15 10 9 4
10 15 13 3 3 8 7 10 9 4 4
6 13 15 1 10 9 4
5 13 15 10 9 4
7 15 13 10 3 0 0 9
8 15 13 10 3 0 0 0 9
7 15 13 10 3 0 0 9
8 3 13 15 10 9 3 4 4
5 15 13 3 0 0
6 3 10 0 9 4 4
6 3 10 0 9 4 4
6 3 10 0 9 4 4
5 10 0 9 4 4
6 15 13 3 15 0 4
12 15 13 12 9 2 3 11 2 11 11 11 2
5 15 4 16 15 9
9 15 4 3 2 16 15 10 9 9
9 15 13 10 9 16 10 9 1 13
4 10 9 4 4
10 15 13 15 10 9 16 10 9 1 13
10 15 13 10 9 15 15 9 4 13 4
11 15 13 15 10 9 15 15 9 4 13 4
9 16 15 9 1 13 13 10 0 9
10 16 15 9 1 13 13 15 10 0 9
10 16 15 9 4 13 4 13 10 0 9
11 16 15 9 4 13 4 13 15 10 0 9
8 15 13 15 1 15 16 15 4
8 15 13 15 10 9 3 1 4
5 15 13 8 9 4
3 10 0 9
3 15 4 4
5 15 13 8 9 4
8 15 13 15 1 9 16 15 4
7 16 15 4 13 15 1 9
7 3 4 3 4 16 15 4
8 3 4 3 4 10 9 1 4
7 9 13 13 15 3 1 4
7 10 0 9 2 3 10 9
7 10 9 2 1 15 10 9
4 10 0 9 13
5 10 15 0 9 13
5 3 4 10 9 4
4 15 3 13 13
7 10 0 9 7 3 13 13
8 10 15 0 9 7 3 13 13
7 15 13 15 16 3 1 13
7 16 15 15 13 16 1 13
7 15 4 16 0 2 0 9
7 12 10 9 4 1 15 4
5 15 13 15 9 4
6 15 16 15 13 15 4
6 15 16 15 13 15 4
4 3 4 15 4
7 15 9 16 15 13 15 4
5 3 4 12 9 4
6 3 4 12 9 9 4
5 3 13 12 9 4
6 3 13 12 9 9 4
7 15 4 13 15 16 15 13
9 15 13 15 0 16 3 16 15 4
9 15 13 15 3 0 0 16 1 4
9 10 0 4 16 15 1 15 9 13
6 15 10 0 13 1 3
6 3 13 10 9 4 4
8 8 4 16 15 1 15 9 13
6 8 1 10 9 4 15
6 10 9 15 15 13 4
8 10 9 4 0 15 15 13 4
11 11 2 3 0 16 3 2 13 3 13 9
11 11 2 3 0 16 3 2 13 3 13 9
11 11 5 3 0 16 3 5 13 3 13 9
6 15 13 15 9 0 2
10 15 13 15 9 0 16 9 1 4 2
10 15 4 10 9 0 3 3 0 1 13
5 3 13 15 4 4
11 15 4 10 9 0 16 15 3 1 0 13
5 15 4 10 9 0
9 15 13 15 10 9 0 16 15 4
9 15 13 15 9 16 10 9 1 13
9 15 4 15 9 16 10 9 1 13
9 15 4 0 15 16 10 9 1 13
6 10 9 16 15 15 13
5 13 9 11 13 15
6 15 13 1 13 9 11
4 15 13 0 11
4 15 13 11 3
5 15 13 1 0 11
10 15 13 1 16 9 16 10 9 3 4
6 3 13 13 15 1 11
3 15 9 3
6 15 4 0 1 15 9
10 15 4 3 0 1 1 15 1 4 4
9 15 4 3 0 3 16 15 3 4
5 15 13 15 16 0
8 15 13 15 16 0 16 1 4
8 15 13 15 16 0 16 15 4
4 15 13 11 4
11 15 16 10 9 1 10 9 13 1 10 9
11 15 16 10 9 1 10 9 13 1 10 9
7 10 10 16 12 9 13 15
11 15 13 10 9 2 3 10 9 2 11 2
13 1 10 12 9 1 0 9 13 11 3 2 12 2
7 15 16 3 13 15 10 9
6 15 13 10 9 16 3
7 15 13 12 9 15 16 3
6 15 13 3 0 16 11
6 15 13 3 12 9 3
5 15 13 11 3 4
5 15 13 15 1 9
5 15 13 8 1 9
11 15 13 15 1 15 9 9 1 9 1 4
10 15 13 15 3 3 3 16 9 0 4
8 15 13 15 9 15 13 13 4
9 15 13 1 10 9 16 9 4 4
7 15 13 8 16 9 0 4
5 7 9 13 15 8
8 15 13 10 9 4 13 1 13
6 9 13 3 10 9 0
6 15 13 11 3 4 4
4 15 13 13 3
5 10 9 13 0 3
6 10 9 13 15 0 3
7 15 13 0 3 16 15 13
8 15 13 15 0 3 16 15 13
8 15 13 15 9 16 15 4 4
7 15 9 9 16 15 4 4
5 15 13 9 1 11
9 12 9 10 9 13 15 10 9 3
11 13 9 16 9 1 13 13 15 15 9 3
7 15 13 11 3 3 4 4
9 15 13 8 16 15 0 9 1 13
3 15 13 8
9 15 4 3 0 1 10 9 1 4
2 3 13
8 16 15 15 9 13 4 1 11
10 16 15 10 9 1 15 9 13 1 11
8 16 15 10 9 4 1 15 9
10 16 15 10 9 1 15 9 4 1 11
10 15 13 2 13 15 2 10 9 4 2
11 15 13 2 3 13 15 2 10 9 4 2
3 10 0 9
6 15 13 11 3 4 4
10 15 13 2 3 13 15 2 15 3 4
10 15 13 15 2 3 13 15 2 3 4
10 15 13 15 3 2 3 13 15 2 4
9 15 13 2 13 15 2 15 3 4
9 15 13 15 2 13 15 2 3 4
9 15 13 15 3 2 13 15 2 4
6 15 13 2 15 0 2
8 15 13 2 15 13 15 4 2
6 15 13 2 1 3 2
8 15 13 1 15 2 13 15 2
7 15 13 11 3 3 4 4
9 15 13 1 15 2 3 13 15 2
13 15 13 1 15 2 3 13 2 13 15 2 10 9
10 15 13 3 2 13 15 2 3 4 2
8 16 15 2 13 15 2 13 2
12 4 15 0 2 3 13 15 2 16 15 13 2
11 4 15 0 2 13 15 2 16 15 13 2
10 13 15 2 13 15 2 10 9 3 2
12 15 13 2 3 13 15 2 13 15 2 4 2
8 15 13 2 15 13 15 3 2
9 15 13 15 2 15 13 15 4 2
4 13 13 15 3
11 15 13 15 3 3 15 13 4 2 9 2
11 16 15 15 3 13 2 15 13 15 4 2
12 15 9 2 13 10 9 3 2 13 12 9 2
13 15 9 2 3 13 10 9 3 2 13 12 9 2
15 16 15 15 9 13 4 1 10 9 7 10 9 15 13 4
9 15 13 2 3 11 2 0 4 2
4 10 3 13 9
4 10 3 13 9
4 15 0 9 13
5 10 9 7 9 8
4 11 13 15 4
10 15 4 8 2 10 0 9 7 9 2
14 10 9 7 10 9 2 9 1 11 2 13 1 3 2
11 9 2 11 2 11 2 11 2 11 2 11
11 9 2 11 2 11 2 11 2 11 7 11
12 9 2 11 2 11 2 11 2 11 2 7 11
12 7 11 2 11 2 11 2 11 2 11 16 11
13 7 11 2 11 2 11 2 11 2 11 2 16 11
6 0 2 16 15 3 13
5 0 16 15 3 13
5 3 16 15 13 2
5 3 13 15 3 4
5 15 13 15 3 2
7 15 13 15 3 8 9 2
7 15 13 15 3 1 15 2
5 10 9 4 3 2
7 11 1 15 9 8 4 13
8 15 13 10 9 7 15 9 8
11 15 13 15 9 1 0 9 2 3 0 8
10 15 4 1 10 0 9 2 16 15 13
10 15 4 1 0 9 2 8 3 1 13
7 10 0 4 1 10 0 9
6 11 13 15 3 4 4
10 15 13 15 10 9 0 16 15 3 4
9 16 15 3 4 13 15 10 9 0
14 15 13 15 1 10 0 9 16 9 7 9 3 1 4
12 9 7 9 3 1 4 13 15 1 10 0 9
8 15 4 10 9 1 3 15 13
6 8 2 3 13 15 9
4 8 10 9 2
6 0 16 15 3 13 2
4 15 4 9 2
8 0 9 4 15 3 10 9 2
6 3 13 15 3 4 4
8 3 4 0 16 15 9 13 2
13 16 3 0 3 3 1 13 2 7 15 13 3 2
3 15 9 2
6 15 16 15 1 13 2
6 15 12 1 10 0 2
5 12 1 15 9 2
6 15 13 3 16 15 12
5 6 2 10 0 9
7 3 2 1 11 13 15 3
7 3 1 11 13 15 4 2
5 3 13 15 11 3
9 3 16 15 15 9 13 15 3 3
8 3 16 15 3 13 4 15 4
4 3 3 15 9
5 3 13 9 1 9
7 3 13 9 3 16 8 4
6 15 4 15 3 1 4
7 15 4 15 16 15 13 4
8 15 13 1 4 16 15 4 4
8 15 4 3 1 4 16 15 4
8 15 4 3 1 4 16 15 4
5 3 13 15 11 4
6 16 15 4 13 1 4
7 7 15 4 13 3 1 4
7 16 15 4 13 3 1 4
9 15 13 3 1 4 4 16 15 4
10 15 13 15 3 0 1 4 16 15 4
4 15 8 4 0
9 3 1 11 11 11 13 15 10 0
14 10 9 7 9 1 0 7 0 9 13 15 9 7 9
7 3 7 11 13 10 9 4
11 9 2 2 15 13 3 10 9 0 4 2
6 3 13 15 11 3 4
5 15 13 3 4 4
5 15 13 3 4 4
6 15 13 3 4 1 4
4 15 13 4 3
6 15 13 4 9 15 9
4 15 13 4 3
3 3 15 2
4 3 1 11 2
3 3 0 2
3 3 3 2
3 10 0 9
7 3 13 15 11 3 4 4
5 3 15 0 13 2
5 3 15 9 13 2
6 3 10 9 1 13 2
7 15 1 13 1 15 9 2
6 11 13 1 15 12 2
5 15 13 3 16 2
9 15 13 16 15 15 3 0 4 2
6 15 13 16 15 13 2
11 15 9 13 16 3 10 9 1 15 9 9
7 15 13 3 16 15 9 4
7 3 13 15 11 3 4 4
8 15 4 10 9 2 9 7 9
5 15 4 15 0 3
9 15 13 15 13 3 16 3 1 13
8 15 13 15 0 3 16 15 13
11 15 13 16 3 1 13 7 3 16 1 13
10 15 13 12 7 16 0 1 4 12 9
6 15 13 3 7 0 3
8 15 9 4 0 7 0 10 9
10 15 13 1 10 9 7 0 1 10 9
12 15 13 16 15 4 7 0 16 15 3 4 4
3 11 4 4
5 15 13 15 12 9
7 10 9 4 15 12 9 4
6 10 9 4 12 9 4
8 1 10 9 9 13 15 9 4
11 1 12 9 13 13 15 1 10 9 12 4
8 15 13 1 15 4 16 1 4
8 15 13 1 15 1 16 1 4
10 10 0 2 2 2 9 13 11 1 12
9 15 4 10 9 15 15 13 7 13
10 13 2 2 15 4 15 0 9 2 2
3 15 4 4
7 15 4 3 0 16 1 13
10 15 4 15 3 0 9 16 3 1 13
11 15 13 3 0 4 16 10 9 1 13 4
4 15 13 1 3
5 15 4 0 1 3
7 15 13 3 8 15 13 4
7 15 4 3 0 3 1 13
6 13 3 3 16 15 13
7 0 13 3 3 16 15 13
6 0 13 4 16 15 13
4 3 4 11 4
7 15 13 15 0 16 15 13
6 16 15 13 13 15 0
6 13 13 15 16 15 13
7 3 13 15 15 16 15 13
9 15 13 15 0 16 3 4 1 4
8 15 13 15 0 3 4 1 4
8 16 3 4 1 4 13 15 0
7 3 4 1 4 13 15 0
9 0 13 15 15 1 3 4 1 4
8 0 13 15 15 3 4 1 4
4 3 4 15 4
8 0 13 15 1 3 4 1 4
7 0 13 15 3 4 1 4
11 15 4 15 10 9 0 16 10 9 1 13
11 15 4 15 10 9 0 16 10 9 4 4
8 15 12 10 9 13 15 9 1
8 0 9 4 16 10 9 0 4
7 1 15 9 2 15 13 3
11 15 4 10 9 3 11 13 16 15 4 4
12 15 13 3 0 11 4 16 10 9 4 4 4
5 15 13 8 15 4
5 3 13 11 4 4
7 15 13 15 16 3 4 4
7 15 13 15 16 3 4 4
7 15 13 15 8 3 4 4
7 3 13 15 10 9 0 3
7 3 13 1 11 10 13 9
6 13 15 2 15 13 3
6 6 2 3 13 10 9
9 15 13 15 16 1 15 9 0 9
6 10 9 13 12 9 1
5 10 9 13 12 9
5 3 13 15 4 4
11 15 13 3 10 9 16 10 9 3 10 9
5 11 13 12 9 9
8 15 13 10 9 1 8 1 9
5 10 9 4 1 9
7 10 9 13 15 8 10 9
4 15 13 15 8
9 1 10 9 1 9 13 15 3 4
5 15 13 1 10 9
6 9 10 9 13 10 9
6 15 13 1 15 4 3
6 15 13 1 10 9 3
4 15 13 1 3
8 15 13 3 15 1 15 4 3
5 15 4 10 9 4
6 15 13 15 10 9 4
6 15 13 15 10 9 4
7 10 9 4 12 9 3 4
5 10 11 13 9 1
5 10 11 13 9 1
6 3 0 16 15 3 13
4 11 2 0 9
8 3 13 15 1 10 9 3 4
8 10 9 13 10 9 1 12 9
6 1 12 8 13 10 9
8 0 3 1 3 7 3 10 9
9 1 15 9 3 13 15 10 0 9
4 15 0 7 0
7 15 12 4 4 16 12 8
8 1 15 12 9 13 15 12 9
7 15 4 1 4 4 1 11
8 15 13 1 4 4 4 1 11
8 10 9 13 15 0 1 10 9
3 10 9 8
3 15 8 2
4 10 15 13 9
8 10 9 10 9 13 13 10 9
11 10 15 8 13 9 13 10 15 8 13 9
4 10 15 13 9
11 10 9 1 11 7 10 9 13 1 10 9
6 1 11 7 3 13 11
6 3 7 15 4 3 0
7 0 0 7 15 4 3 0
5 15 2 16 15 13
4 15 16 15 13
5 1 12 9 1 11
5 15 16 3 1 13
6 15 2 16 3 1 13
5 15 1 15 0 9
6 15 2 1 15 0 9
9 15 9 2 0 7 0 13 4 2
7 3 0 3 15 4 15 0
7 3 0 15 4 2 3 0
9 3 0 15 4 2 8 0 15 4
9 8 0 15 9 2 8 0 15 4
7 8 13 10 9 1 15 8
4 0 9 1 11
12 10 9 1 11 2 7 10 9 13 1 10 9
7 1 11 2 7 3 13 11
7 3 2 7 15 4 3 0
8 0 0 2 7 15 4 3 0
8 0 3 3 1 13 13 15 0
6 15 4 10 9 11 0
6 15 13 16 1 4 2
4 9 11 13 4
4 13 15 13 4
4 16 15 9 4
7 16 6 2 15 13 3 2
3 15 4 4
4 15 4 3 4
3 15 4 4
3 15 4 9
4 15 4 4 4
6 15 13 15 3 4 3
5 15 13 15 4 8
3 15 13 3
8 15 13 3 16 15 0 1 13
5 1 3 4 15 0
6 15 2 8 2 13 9
5 3 0 13 15 2
10 3 0 13 15 16 15 0 1 13 2
7 15 13 3 13 16 15 13
8 15 13 3 0 13 16 15 13
4 15 13 15 8
8 15 4 15 9 3 3 4 4
9 3 0 10 9 2 3 0 15 9
7 3 0 10 9 2 3 0
9 3 0 10 9 2 3 0 15 4
8 3 0 10 9 4 2 8 0
13 15 5 3 0 16 10 9 5 13 15 9 3 4
9 15 13 10 9 3 2 4 2 4
8 15 13 3 3 16 15 3 4
7 15 13 3 3 0 1 4
5 15 13 3 9 3
6 3 4 10 9 3 1
3 15 13 3
4 15 13 3 3
5 3 3 13 15 3
4 0 13 15 3
4 15 13 1 3
9 15 13 10 9 15 0 0 1 4
5 15 13 1 3 3
5 15 13 3 4 4
4 15 13 4 4
4 15 13 4 4
6 10 1 13 0 9 13
6 10 9 13 13 9 13
5 10 1 13 12 9
5 10 16 13 12 9
8 3 13 3 1 4 16 15 4
8 3 13 3 1 4 16 15 4
10 10 9 4 0 2 15 13 3 1 11
7 15 15 13 4 16 15 13
8 15 15 15 0 4 16 15 13
7 15 13 15 1 10 9 4
8 15 13 15 3 4 1 15 9
10 16 15 15 9 13 4 2 4 15 0
4 1 3 3 0
5 11 2 3 13 15
6 10 9 2 3 4 15
7 15 13 2 2 3 13 15
12 3 13 15 15 1 15 9 16 15 1 4 2
7 6 2 11 13 3 3 2
9 15 13 15 12 9 8 16 1 4
4 15 4 11 0
4 3 13 13 15
5 15 4 3 13 2
8 15 4 2 3 2 2 3 0
8 15 4 2 3 2 2 3 0
8 15 4 2 3 2 2 3 0
8 10 9 4 3 3 0 3 2
9 15 13 10 9 3 3 0 3 2
5 15 13 11 16 8
5 15 13 9 13 2
5 15 13 11 16 8
7 3 1 2 3 7 3 2
12 15 13 1 9 2 13 11 2 7 15 4 0
16 2 15 13 1 9 2 2 13 11 2 2 7 15 4 0 2
9 15 3 16 11 13 15 4 4 2
7 15 3 13 15 4 4 2
7 10 9 3 2 7 15 13
9 15 9 13 15 1 13 1 10 9
8 15 9 4 16 0 3 1 4
9 15 9 13 15 3 16 3 1 13
9 1 11 7 3 3 4 15 10 0
6 15 8 13 3 3 2
6 15 16 15 13 10 9
6 3 13 15 9 9 11
10 8 2 9 10 11 2 13 1 10 9
6 15 4 3 0 3 0
6 15 13 3 0 3 0
9 15 13 3 2 15 13 16 15 4
8 15 4 0 7 1 0 7 9
8 15 4 0 7 1 9 16 9
7 15 4 15 0 16 15 13
9 15 4 15 0 16 1 11 1 13
7 11 15 9 15 9 13 2
6 10 9 13 15 3 3
6 15 13 10 9 3 1
6 1 0 3 1 4 2
4 10 8 9 2
5 15 4 10 9 4
7 3 13 0 0 7 9 13
4 3 4 1 3
5 3 13 15 1 3
5 15 13 3 1 0
4 15 13 1 3
5 15 15 9 13 2
7 15 13 4 1 3 15 13
7 15 13 3 16 15 4 4
5 15 9 4 15 9
7 10 0 3 1 13 9 2
8 15 9 13 3 1 4 4 2
10 15 13 10 0 9 16 0 0 4 2
6 15 13 3 1 0 13
7 10 0 9 13 9 9 1
10 16 15 15 10 9 1 10 9 13 2
9 16 15 15 15 1 10 9 13 2
7 3 13 1 15 9 0 9
8 3 15 3 13 4 16 15 4
8 3 15 3 13 4 16 1 4
7 3 15 3 13 4 1 4
10 3 15 15 3 13 4 4 16 15 4
10 3 15 3 0 1 4 4 16 15 4
9 3 15 15 1 9 4 16 15 4
13 3 15 15 3 13 4 4 4 4 4 16 15 4
8 15 13 0 7 16 15 4 4
8 15 13 16 7 3 15 4 4
10 15 13 3 7 3 15 15 0 4 4
6 1 15 9 13 0 9
10 15 13 0 7 3 15 15 0 4 4
8 15 13 16 7 3 15 4 4
8 15 13 3 7 16 15 4 4
10 15 13 16 15 0 4 4 16 15 13
7 15 13 8 10 9 1 9
5 15 4 10 0 9
6 15 13 1 3 12 9
13 15 13 1 3 0 1 13 9 1 10 1 13 9
9 15 13 1 10 3 0 1 13 9
9 10 9 15 15 3 3 3 13 4
5 3 13 0 9 1
10 15 13 15 10 9 3 4 16 15 4
11 15 13 15 1 10 9 3 4 16 15 4
7 15 13 2 15 13 3 2
8 15 13 11 1 11 7 3 15
9 16 15 3 13 16 13 15 10 9
6 8 16 13 15 10 9
6 15 13 4 15 15 13
6 15 13 13 15 1 9
7 10 9 13 0 4 16 4
8 16 15 15 13 2 13 3 3
6 0 13 3 0 9 1
8 3 4 15 1 4 16 15 4
4 15 3 9 2
8 16 15 13 2 13 1 15 2
9 16 15 4 4 1 15 1 4 2
9 3 16 1 13 7 16 3 1 13
10 11 2 1 9 10 9 2 13 12 9
6 0 9 13 3 0 1
3 8 12 9
4 8 12 12 0
9 15 13 7 7 8 16 15 4 4
10 15 13 7 7 8 1 15 15 4 4
8 15 13 7 7 8 15 15 4
8 15 13 10 9 3 8 15 9
3 15 13 9
6 8 0 13 15 4 2
7 13 4 9 7 0 4 0
7 15 13 1 15 9 10 9
3 15 13 8
4 15 13 3 4
6 16 15 3 3 13 4
6 15 4 15 15 9 0
7 15 4 15 15 10 9 0
7 15 4 15 0 1 10 9
9 15 4 15 3 0 1 16 15 4
8 15 4 15 3 16 15 4 4
10 15 4 15 3 3 3 0 16 15 4
10 15 4 15 3 3 3 3 16 1 4
7 1 15 9 13 15 10 9
7 15 4 15 0 1 15 13
8 15 4 15 3 1 9 1 4
10 4 15 15 3 7 0 1 10 9 2
11 4 15 15 3 7 0 16 10 9 4 2
4 9 9 12 2
6 15 13 15 8 4 2
8 15 13 10 9 1 10 9 4
8 15 13 2 0 7 0 9 2
8 10 13 9 4 1 12 4 2
8 10 9 4 15 1 12 4 2
6 15 13 0 13 1 3
6 15 13 3 10 9 1
8 10 9 9 13 1 12 4 2
10 10 9 9 13 15 9 1 12 4 2
4 15 0 13 2
7 15 13 15 9 1 15 9
8 15 13 15 10 9 1 15 9
6 15 4 4 1 15 9
6 15 13 4 1 15 9
8 15 13 10 9 4 1 15 9
8 15 4 10 9 4 1 15 9
12 1 10 9 2 15 13 3 3 10 9 4 2
10 10 9 16 15 3 0 3 13 4 0
13 1 10 9 2 2 15 13 3 3 10 9 4 2
8 15 12 13 15 12 1 15 12
6 15 13 12 13 15 3
9 1 8 3 15 12 10 9 3 13
12 15 13 10 9 1 9 16 2 15 4 0 2
14 15 13 1 9 16 2 2 15 4 0 2 2 10 9
13 1 10 9 2 15 13 3 3 10 9 4 2 2
11 1 10 9 2 15 13 3 3 10 9 4
5 15 13 3 0 8
5 3 4 0 8 9
9 10 9 15 3 0 3 13 4 0
7 15 13 15 10 0 9 4
7 15 13 15 10 0 9 3
8 3 13 15 16 15 15 9 13
13 10 9 15 15 10 0 9 13 4 13 15 9 3
8 15 13 15 1 0 16 15 4
8 15 13 15 1 0 3 1 4
5 15 13 15 1 0
9 15 13 15 1 10 9 15 15 4
9 15 13 15 1 10 9 3 1 4
6 15 13 15 1 10 9
4 15 8 13 13
8 15 13 15 1 10 9 7 0
6 9 11 9 4 3 4
6 9 11 9 4 3 4
8 3 13 3 3 15 0 3 13
9 3 4 3 3 1 4 15 15 13
7 15 13 3 15 15 3 13
9 15 13 0 4 13 15 1 9 4
11 15 13 0 4 2 13 15 3 1 9 4
7 15 13 3 13 15 0 4
10 10 9 2 13 15 0 4 2 13 3
8 10 9 13 2 15 2 1 11
5 15 13 10 12 9
8 15 13 10 9 7 1 10 9
7 16 15 1 15 3 9 13
7 15 13 16 16 15 1 13
9 15 9 2 13 9 2 4 15 0
6 15 13 10 0 3 0
14 1 10 9 1 16 11 3 11 2 11 2 11 7 11
6 10 9 13 15 3 2
6 15 9 13 15 3 2
8 3 0 13 15 3 3 0 2
10 10 9 13 2 3 0 2 1 10 9
7 3 3 13 15 1 0 2
7 15 13 10 9 16 15 4
11 15 13 10 9 15 9 15 15 1 11 4
10 15 4 3 10 9 1 10 9 1 13
7 15 1 13 13 15 3 4
9 13 15 15 1 13 7 1 13 2
1 2
4 15 0 13 2
3 15 13 0
9 16 15 15 3 1 10 9 0 4
7 15 13 10 9 16 1 13
8 16 15 15 3 16 1 0 4
11 16 15 15 3 3 1 0 4 16 15 4
10 16 15 15 3 3 1 0 4 1 4
10 16 15 15 3 3 0 4 16 15 4
9 16 15 15 3 3 0 4 1 4
7 10 9 0 13 15 3 3
8 16 15 15 16 10 9 0 4
9 15 10 9 0 13 15 1 10 9
9 10 15 10 9 0 9 13 3 3
4 10 3 0 9
13 15 13 15 3 10 9 1 3 15 10 9 4 4
10 10 15 3 3 1 0 9 13 10 9
8 15 13 12 0 7 10 0 9
7 15 13 10 9 3 7 3
7 10 15 16 15 13 3 4
8 15 13 0 10 15 3 15 2
8 15 4 0 16 7 8 15 13
10 15 13 10 9 15 9 12 9 4 2
5 13 4 13 9 13
6 15 13 1 11 13 2
6 10 12 1 0 9 13
8 15 13 15 9 3 1 15 9
8 10 15 1 0 9 13 10 9
5 10 12 1 0 9
7 10 15 1 0 13 10 9
5 4 10 0 0 9
8 1 15 7 15 4 15 9 2
10 15 13 1 15 7 15 15 0 4 4
9 15 13 3 13 16 15 3 4 4
11 16 15 3 3 13 13 16 15 3 4 4
10 15 13 15 3 3 3 13 16 15 4
10 15 13 15 3 13 16 1 15 1 4
8 15 4 16 10 9 15 15 13
8 15 13 15 3 13 16 15 4
10 15 9 4 0 16 1 10 9 1 4
8 15 9 4 0 16 3 1 4
9 15 9 4 3 0 16 3 1 13
9 15 9 4 0 15 16 3 1 13
11 15 9 4 0 15 1 4 16 3 1 13
7 16 15 9 13 15 3 3
9 1 15 9 4 8 3 3 1 2
13 0 13 0 16 10 9 3 4 3 15 13 9 2
6 10 9 3 3 15 13
9 15 13 2 0 16 3 0 1 4
7 15 4 1 9 16 15 13
12 16 3 15 3 13 2 13 10 9 3 0 0
6 15 13 3 10 9 3
7 3 3 4 0 15 3 13
9 3 3 4 15 8 1 3 4 2
11 3 13 4 16 10 9 1 10 9 13 2
15 3 13 15 15 9 3 2 13 10 9 0 2 7 13 2
7 10 9 13 9 3 3 12
6 15 9 13 3 3 3
8 15 13 1 15 9 3 4 2
5 15 2 0 2 13
5 15 4 15 15 13
5 10 2 0 2 9
6 15 4 2 0 2 13
6 2 7 15 3 2 2
6 2 7 15 3 2 2
5 2 7 15 3 2
3 2 2 2
6 15 13 2 12 2 9
9 15 13 10 9 2 7 15 9 2
10 15 13 10 9 2 7 3 15 9 2
13 15 13 10 9 2 7 2 16 13 2 15 9 2
7 4 15 16 15 3 13 2
12 15 13 10 9 4 2 15 15 3 0 13 2
7 10 1 11 9 7 13 9
8 15 4 10 0 9 1 10 9
16 15 8 13 10 0 9 3 2 15 3 4 4 1 13 9 2
12 10 9 11 4 10 9 2 9 4 15 3 4
8 10 2 1 15 3 0 2 9
6 15 4 2 3 2 0
6 15 13 4 2 4 15
6 15 13 4 2 4 15
7 15 13 4 2 13 15 1
7 4 15 16 15 3 13 2
8 10 12 9 13 3 1 10 9
4 15 4 9 9
6 15 4 8 9 1 9
5 8 13 10 9 4
9 3 3 1 15 9 4 15 3 0
8 3 1 15 9 4 15 3 0
6 15 15 4 16 15 13
10 7 15 4 15 15 16 0 3 1 13
7 13 1 10 0 13 15 4
7 12 1 10 0 13 15 4
7 15 4 15 15 3 13 2
7 13 1 10 0 13 15 4
7 12 1 10 0 13 15 4
4 11 15 3 2
7 10 9 3 2 3 2 11
7 10 9 3 2 3 2 11
7 10 9 3 2 6 2 11
10 15 0 8 2 7 2 10 0 9 2
8 10 9 1 3 2 0 9 2
7 15 4 15 15 3 13 2
8 15 4 15 4 15 15 13 2
9 15 4 15 1 4 15 15 13 2
8 15 4 10 9 1 3 4 2
7 10 15 13 1 10 9 2
8 15 4 10 0 9 1 11 2
9 15 9 3 1 10 9 13 8 4
9 10 9 1 12 9 3 13 15 0
7 1 15 3 4 1 8 4
8 10 0 9 3 13 10 9 4
11 15 13 16 16 10 9 13 2 10 9 4
5 10 8 12 0 2
4 15 12 0 2
4 15 12 0 2
4 15 0 12 0
10 10 9 13 12 2 12 2 12 9 2
10 15 13 1 9 2 15 13 3 4 2
11 10 9 13 12 2 3 12 2 12 9 2
8 10 0 9 1 10 9 4 8
6 15 0 13 13 16 9
12 10 9 13 1 15 12 7 15 12 12 9 2
10 10 9 13 1 12 7 12 12 9 2
11 10 9 13 1 15 12 7 12 12 9 2
2 6 2
10 2 13 15 3 2 2 2 13 15 2
8 15 13 3 2 2 13 15 2
9 15 13 10 9 7 9 16 0 4
11 15 4 1 11 2 12 9 2 15 9 2
6 15 13 0 9 12 9
6 15 4 15 9 0 2
11 15 4 15 15 0 16 15 16 1 13 2
11 15 4 15 15 0 16 15 3 3 13 2
7 15 13 3 2 13 15 2
7 15 13 3 3 1 4 2
7 15 13 1 9 4 10 9
6 15 9 13 4 10 9
6 15 1 11 13 13 15
7 15 13 1 11 4 10 9
6 9 5 9 1 10 9
8 15 13 16 10 9 4 4 9
7 15 13 3 1 4 13 3
6 15 0 4 4 15 0
9 15 15 1 11 9 9 4 10 9
7 15 9 13 4 4 3 9
9 15 10 0 9 13 4 13 15 9
10 15 10 0 9 1 13 4 13 15 9
7 10 3 0 9 4 8 9
11 10 8 0 9 4 3 0 16 0 1 4
9 15 9 13 7 13 13 15 0 15
5 11 3 1 15 8
8 15 0 13 1 10 9 13 9
14 15 3 3 13 13 7 3 15 9 13 13 13 4 2
6 15 13 1 15 7 3
5 15 13 12 1 11
5 15 10 9 13 9
4 10 15 13 9
5 10 9 8 13 9
4 10 0 13 9
4 10 0 13 9
5 10 15 9 13 9
10 15 8 10 0 0 9 1 10 9 2
22 10 9 13 3 16 3 10 9 1 12 9 3 10 0 9 4 8 10 3 13 9 2
22 15 13 3 9 4 4 3 13 13 15 15 13 2 3 15 15 13 2 15 3 13 2
13 10 9 13 1 10 9 1 15 13 1 15 8 2
18 10 9 11 2 9 1 10 0 9 2 4 12 9 3 9 1 11 2
18 10 9 1 10 9 8 2 8 2 7 8 2 0 2 4 8 4 2
11 15 4 10 9 1 0 9 8 7 8 2
18 10 9 11 13 16 9 1 11 7 10 9 11 4 13 1 10 9 2
21 1 15 9 13 15 4 16 3 9 4 1 10 9 7 10 9 3 0 4 4 2
25 10 9 1 10 9 1 10 9 13 9 1 15 9 4 2 15 1 10 9 1 10 9 13 4 2
8 15 9 4 3 0 1 4 2
12 0 4 15 3 1 10 9 1 15 8 13 2
22 10 9 13 3 3 15 9 10 9 1 13 2 16 3 10 9 9 1 9 13 4 2
16 8 13 15 13 9 3 1 10 0 9 1 10 9 4 4 2
12 10 9 12 3 10 9 1 15 9 3 0 2
6 10 9 13 0 3 2
7 10 8 9 13 12 9 2
21 1 10 9 4 10 9 1 10 0 9 1 10 9 7 13 10 9 12 9 3 2
15 16 10 9 3 3 3 3 0 4 2 4 10 9 0 2
9 12 9 13 9 1 12 10 9 2
12 9 4 10 0 13 7 3 0 13 9 9 2
10 15 4 10 9 15 3 15 9 13 2
48 8 2 10 0 2 7 0 9 1 10 0 0 9 2 13 1 12 3 4 2 16 11 10 9 4 16 2 0 9 1 0 9 2 1 4 7 3 2 10 9 1 15 15 9 2 1 4 2
18 1 8 2 10 9 1 10 0 0 9 2 4 15 9 3 0 4 2
10 11 13 10 1 15 13 9 0 0 2
45 10 13 9 7 9 1 10 9 2 15 13 13 1 0 9 13 1 10 15 9 3 1 10 9 1 10 9 4 2 16 15 1 10 13 9 9 1 10 9 3 15 13 13 4 2
22 15 4 15 9 15 13 9 1 9 1 10 2 0 2 2 15 13 9 4 13 4 2
9 3 4 11 9 1 15 9 0 2
35 15 9 13 10 9 10 9 16 10 9 10 9 1 15 13 2 15 1 3 0 9 4 16 15 0 4 2 1 10 0 9 3 1 13 2
8 3 13 15 3 1 10 9 2
49 11 4 3 10 9 1 4 10 9 3 15 1 10 9 1 13 7 3 10 9 1 13 1 10 9 1 10 9 16 8 0 13 9 1 9 0 3 3 0 13 9 1 9 1 13 7 1 13 2
5 0 13 15 3 2
20 10 9 8 15 1 11 2 10 0 9 2 4 2 13 3 10 0 9 3 2
24 10 0 0 9 4 3 15 0 2 3 3 10 9 1 15 13 1 10 0 9 1 10 9 2
9 2 1 11 13 10 9 3 3 2
24 11 4 15 0 0 1 10 0 9 5 16 15 1 11 13 2 15 13 3 1 10 0 0 2
10 15 13 10 9 3 7 13 15 9 2
19 3 13 3 10 0 4 4 4 16 10 0 9 15 15 1 10 9 13 2
13 15 4 13 2 0 2 13 3 15 1 15 9 2
22 1 10 9 9 7 9 4 10 0 9 1 4 1 8 7 10 9 1 10 0 9 2
35 10 9 4 16 1 11 10 0 0 9 3 10 9 4 4 2 8 15 15 13 4 1 4 1 10 0 9 15 1 15 15 9 4 4 2
29 1 10 9 1 10 9 4 15 1 4 16 0 10 0 9 2 10 0 9 1 10 0 9 2 8 7 8 4 2
30 15 0 0 9 13 1 10 9 1 15 15 1 10 9 7 10 1 15 9 3 0 9 2 9 7 9 3 1 4 2
37 15 13 15 3 3 2 7 3 13 15 11 0 9 1 9 1 10 0 9 2 7 3 1 10 0 2 0 0 0 2 15 1 11 3 13 4 2
23 1 11 2 15 15 1 10 0 9 13 4 1 10 0 9 2 4 15 15 3 1 4 2
24 3 3 1 11 13 1 10 0 9 8 2 0 1 15 8 2 10 9 8 2 9 8 2 2
17 15 11 13 11 1 15 9 3 9 7 9 1 9 7 9 4 2
19 1 10 9 13 10 0 9 5 3 3 1 10 9 5 1 10 13 9 2
13 15 0 13 9 13 10 9 1 15 9 1 13 2
25 3 13 3 3 10 0 9 1 10 0 9 1 8 2 8 2 8 2 11 2 9 8 2 4 2
14 1 15 13 1 9 4 3 3 1 10 0 9 4 2
15 10 9 0 9 4 2 9 4 7 10 0 0 9 4 2
27 1 10 9 3 3 4 3 10 9 1 10 9 4 3 10 9 0 13 4 4 1 15 9 1 10 9 2
11 9 2 9 2 9 2 0 9 7 9 2
23 3 1 10 9 2 3 2 3 2 2 7 0 1 0 9 1 10 9 1 10 15 9 2
21 15 13 15 3 3 3 1 10 9 1 10 0 2 15 0 9 7 9 15 13 2
23 10 9 1 15 8 2 8 2 9 1 11 2 13 11 1 9 11 9 7 10 9 4 2
22 10 0 9 2 8 2 13 9 2 3 1 10 0 9 2 10 9 4 1 9 11 2
7 3 4 12 0 9 4 2
16 15 13 3 15 0 9 3 1 10 9 1 10 0 0 9 2
13 10 13 0 13 3 0 9 2 3 10 9 8 2
27 10 9 13 3 10 9 1 12 12 9 2 3 0 12 1 12 12 4 4 1 10 9 7 10 0 9 2
24 15 13 3 1 0 9 1 15 9 16 10 13 0 2 15 15 9 3 3 1 9 13 4 2
12 10 13 0 13 8 15 1 15 9 7 9 2
35 16 1 10 0 3 13 9 4 10 0 9 2 15 1 11 0 9 4 2 1 10 11 13 9 0 1 10 0 9 0 1 10 13 9 2
16 1 10 9 11 13 10 9 1 12 1 12 1 10 12 9 2
14 9 4 16 1 10 9 3 10 9 7 3 10 9 2
13 10 9 13 1 10 9 3 1 12 1 12 9 2
19 7 1 10 0 13 10 9 3 3 0 4 3 3 15 7 3 15 4 2
13 15 13 15 1 9 7 9 1 10 9 11 3 2
20 15 2 16 10 9 1 10 9 3 0 4 7 15 7 15 10 0 9 13 2
20 1 0 9 13 10 9 10 9 16 15 1 10 9 1 15 9 0 13 4 2
22 10 9 1 15 9 4 1 15 9 3 1 8 12 1 12 4 1 8 12 1 12 2
4 3 15 9 2
31 10 13 9 13 2 8 10 1 15 0 9 2 11 10 9 1 9 1 9 7 9 2 3 10 9 0 3 4 2 4 2
25 1 10 13 11 13 11 3 10 9 4 16 2 1 10 9 1 15 9 2 10 13 9 1 4 2
7 7 3 13 10 9 3 2
41 3 4 9 8 9 10 2 13 2 9 4 2 13 3 1 10 9 0 9 2 9 2 9 2 9 2 9 7 9 2 15 0 0 4 16 15 0 9 1 4 2
27 16 15 9 1 10 0 9 2 15 15 3 10 0 9 4 2 1 10 9 4 4 2 4 3 0 3 2
3 3 8 2
15 2 10 0 9 7 3 10 9 1 8 13 15 1 15 2
14 15 1 10 0 9 1 15 9 2 4 10 0 9 2
22 8 15 15 9 1 0 9 3 3 0 13 13 1 15 11 11 0 9 1 15 9 2
26 1 8 13 15 3 5 7 15 1 3 13 9 5 10 9 3 16 15 1 10 0 9 0 1 4 2
23 1 15 0 9 13 3 10 9 4 3 15 0 9 2 9 12 2 15 15 9 4 4 2
13 15 13 9 4 0 1 10 13 9 1 10 9 2
15 3 13 10 9 1 11 2 15 11 3 3 13 4 4 2
5 8 13 11 8 2
7 15 13 10 9 3 3 2
17 15 13 15 3 0 4 2 7 10 0 9 4 0 4 1 8 2
16 11 2 15 16 9 3 15 9 4 2 13 3 15 3 0 2
11 7 1 11 15 4 10 0 9 3 0 2
15 15 13 10 9 1 8 1 7 13 10 0 9 1 11 2
18 11 13 1 10 0 9 1 11 0 3 7 13 10 0 9 1 12 2
17 11 13 0 3 1 10 9 1 12 1 10 9 1 10 9 11 2
22 8 10 0 9 13 8 2 15 0 13 2 12 2 1 11 2 11 1 10 0 9 2
12 11 13 3 12 9 1 11 7 11 15 12 2
18 10 0 9 8 13 10 0 9 1 10 0 9 2 12 2 1 8 2
16 10 9 13 3 1 0 1 11 2 15 10 0 9 8 13 2
33 11 13 12 9 1 9 10 9 15 0 1 10 9 2 12 2 7 11 13 1 10 0 9 1 10 0 9 3 0 2 12 2 2
22 1 10 0 9 4 12 2 2 2 9 3 15 1 11 16 8 10 15 9 1 4 2
14 11 4 15 9 1 10 0 9 4 1 3 13 13 2
23 3 0 10 9 3 13 4 2 16 15 4 4 4 1 10 0 9 1 0 9 0 0 2
32 16 10 15 9 15 13 2 13 7 13 2 16 1 10 9 8 1 11 2 13 15 0 0 9 3 1 3 10 9 9 4 2
27 15 4 16 10 0 9 1 10 9 1 10 0 9 1 10 1 8 13 9 2 1 12 0 1 15 8 2
30 15 13 3 3 3 4 16 10 9 15 9 8 15 3 4 4 2 3 13 10 9 10 0 9 15 0 1 10 9 2
18 1 10 9 2 3 13 10 0 9 8 4 10 11 1 12 9 13 2
12 11 2 11 7 16 0 9 11 7 10 9 2
15 0 0 13 15 4 1 10 9 1 9 1 11 7 11 2
29 1 10 9 4 3 3 1 9 1 0 9 1 10 9 10 9 3 4 16 10 3 0 9 1 0 9 1 13 2
21 1 0 9 1 11 4 1 10 13 9 3 12 9 7 10 0 9 9 13 4 2
17 12 9 1 10 0 9 13 1 10 0 9 1 10 9 4 4 2
7 3 4 3 12 9 4 2
9 15 4 3 8 1 15 0 8 2
33 10 0 9 4 10 0 9 2 15 11 13 13 4 2 7 3 4 3 3 10 9 1 9 15 1 10 9 10 0 9 13 4 2
22 10 9 4 8 4 7 10 9 0 4 2 7 1 10 9 1 9 7 9 0 4 2
11 9 1 10 9 7 10 9 4 0 4 2
24 12 9 2 15 15 1 9 9 2 13 9 1 11 7 11 1 10 9 1 3 12 9 4 2
35 10 9 1 11 13 11 3 2 16 9 1 11 7 1 11 10 9 2 15 1 11 10 9 13 2 9 4 4 2 15 15 1 9 13 2
12 10 9 1 10 9 4 3 1 0 9 4 2
12 16 10 9 10 9 13 4 10 9 3 4 2
13 15 13 16 10 9 4 4 16 3 15 9 4 2
12 10 9 13 3 0 4 2 7 10 9 13 2
8 2 10 9 13 1 4 2 2
16 10 9 8 13 15 3 16 15 3 3 3 0 4 1 11 2
18 12 0 9 13 1 10 9 1 10 0 9 10 9 1 15 9 4 2
16 3 13 3 3 15 9 7 10 9 4 3 3 2 13 15 2
13 1 10 9 1 11 13 15 3 15 0 9 3 2
15 10 15 0 9 4 15 0 13 1 0 9 1 10 9 2
31 1 10 0 9 2 1 9 7 9 2 13 3 3 3 3 0 9 2 15 16 10 9 0 8 9 2 10 0 9 4 2
16 15 4 1 9 15 3 3 15 0 15 1 10 9 4 4 2
9 0 13 3 1 15 9 0 9 2
11 10 9 4 4 1 10 0 7 0 9 2
26 1 15 12 7 12 12 9 13 8 7 8 4 1 10 0 9 1 9 1 10 9 1 10 0 9 2
9 3 13 15 1 15 9 3 9 2
17 10 9 13 1 10 12 9 0 9 1 11 7 8 1 10 11 2
34 9 13 10 0 9 1 10 2 9 9 2 2 16 15 0 0 4 2 16 9 8 7 10 9 11 15 3 3 3 1 15 13 4 2
12 1 10 16 12 9 9 13 10 9 4 4 2
8 10 9 13 9 12 4 4 2
6 3 10 9 4 4 2
17 12 9 1 12 9 4 1 15 0 2 3 12 9 13 9 0 2
34 10 9 8 1 11 13 3 0 8 2 13 1 15 13 1 10 9 1 10 0 0 9 7 13 10 9 1 10 9 0 4 1 4 2
8 2 10 9 4 8 9 2 2
21 1 15 13 1 10 9 1 12 1 12 13 15 16 10 9 10 9 0 0 4 2
10 11 13 15 3 16 15 1 9 4 2
17 12 9 0 13 15 15 15 4 7 12 9 4 15 9 3 4 2
7 15 9 4 15 0 3 2
23 15 9 3 2 7 12 9 13 0 15 9 1 10 9 2 3 10 0 9 8 13 4 2
3 3 8 2
14 12 9 1 15 9 1 11 13 10 9 3 0 0 2
16 15 13 7 13 15 3 7 13 1 15 9 1 9 4 4 2
19 2 15 13 3 16 10 9 2 0 3 3 11 2 0 2 2 13 15 2
11 11 13 1 10 9 1 10 0 0 9 2
43 1 15 9 2 3 15 10 9 13 1 10 9 1 10 11 1 10 0 11 2 13 11 1 10 9 3 10 15 9 1 10 0 9 4 16 1 12 8 1 10 9 13 2
27 11 2 15 1 9 10 0 4 2 13 0 3 1 10 0 0 9 11 2 15 15 3 3 0 3 13 2
21 10 0 9 1 15 4 16 10 9 1 10 15 9 1 10 11 13 3 1 4 2
18 3 3 13 10 0 9 9 1 10 0 9 1 15 8 1 11 4 2
34 10 9 1 15 9 4 16 11 3 1 4 10 0 9 1 4 7 10 1 11 13 9 1 10 0 0 9 1 15 9 0 1 4 2
34 10 9 4 10 9 1 10 0 9 3 3 4 2 16 8 1 10 9 1 10 9 11 10 9 13 15 0 13 2 13 16 10 9 2
7 1 3 15 9 1 8 2
24 1 12 9 13 10 0 11 3 0 8 2 7 3 2 16 1 11 13 2 1 10 0 9 2
14 10 0 9 16 10 0 9 15 1 15 9 4 4 2
13 16 3 15 9 13 13 10 11 3 3 4 4 2
11 8 2 10 3 13 9 2 13 1 3 2
22 3 3 1 10 11 13 15 16 3 3 1 13 1 10 9 1 13 9 1 10 9 2
24 16 11 4 11 4 1 10 9 11 2 3 15 3 1 11 0 9 1 9 2 8 4 4 2
4 3 10 9 2
46 10 9 13 10 0 9 1 15 13 1 15 1 9 13 9 2 3 10 9 2 7 8 10 0 9 8 13 2 2 7 10 0 0 9 8 13 15 9 1 10 9 7 10 0 9 2
22 1 15 10 9 0 13 4 15 0 0 2 15 13 3 0 15 1 10 9 4 4 2
18 15 13 0 3 2 7 15 13 3 3 10 9 15 1 4 4 2 2
11 3 13 11 3 3 1 9 4 1 4 2
19 15 13 3 1 10 9 2 15 15 3 0 13 2 4 1 11 7 11 2
25 10 9 13 15 1 10 9 8 4 1 10 9 2 16 10 9 1 11 10 0 0 9 4 4 2
15 1 10 9 13 10 9 0 9 4 1 10 9 10 9 2
14 3 13 10 0 9 1 11 15 16 3 3 1 13 2
18 10 0 9 4 12 9 2 10 9 4 1 10 9 8 0 12 9 2
42 1 10 0 9 4 4 12 9 9 2 10 9 7 9 1 10 0 9 7 1 0 9 2 10 9 2 10 9 0 9 2 10 9 8 2 10 9 7 10 0 9 2
9 1 9 13 10 9 1 12 9 2
19 15 8 2 12 9 2 13 16 0 9 13 4 1 10 9 1 15 9 2
17 1 15 9 13 10 9 2 10 9 2 3 0 9 2 3 8 2
16 8 4 3 0 3 4 2 16 9 7 9 0 1 15 4 2
20 2 3 3 4 15 3 3 0 1 9 7 0 9 10 13 0 9 1 13 2
13 3 3 13 15 10 0 9 1 9 7 9 2 2
25 8 13 3 2 16 10 9 1 0 13 0 3 0 4 4 16 15 9 13 1 15 9 1 9 2
25 3 13 3 10 9 16 10 9 10 9 4 2 3 15 10 9 3 1 13 16 15 3 1 13 2
13 15 13 0 9 4 2 15 9 2 9 7 9 2
20 10 0 9 4 15 3 15 15 13 1 10 9 1 15 15 8 13 4 2 2
8 15 0 9 4 3 0 13 2
22 10 0 0 9 1 10 9 4 1 3 0 9 4 1 10 0 9 2 13 8 3 2
29 10 0 9 13 3 10 9 4 2 7 15 13 10 9 3 3 1 15 0 16 15 15 1 9 1 10 9 13 2
8 15 13 3 3 10 0 9 2
19 2 3 4 3 10 9 3 2 16 10 0 9 7 11 15 3 8 4 2
37 7 16 10 9 1 11 2 1 10 9 1 12 9 1 8 2 9 1 15 9 2 2 1 10 9 1 9 9 13 4 3 4 15 10 9 3 2
31 10 9 15 16 9 1 9 13 2 4 8 8 8 3 1 4 1 10 9 16 16 15 3 3 10 0 9 1 15 13 2
35 9 7 9 13 10 9 4 2 16 1 10 9 11 8 9 4 1 10 9 7 9 1 10 0 9 7 1 10 9 1 10 11 1 11 2
15 3 13 10 9 10 9 16 10 9 1 8 0 1 4 2
26 1 10 9 1 15 9 13 3 10 9 1 8 2 11 2 8 2 11 2 11 7 8 4 4 4 2
37 1 10 9 8 2 15 8 10 0 9 10 9 13 4 1 10 9 1 10 9 1 10 0 9 2 4 10 0 9 8 1 15 9 0 8 4 2
19 15 4 4 1 9 7 13 15 15 1 10 9 4 7 15 9 15 13 2
19 10 9 13 10 9 2 10 9 11 2 1 15 8 3 1 10 9 4 2
59 16 0 9 4 4 8 2 7 8 15 9 2 3 10 9 16 10 9 10 0 9 4 4 7 16 15 0 4 16 10 9 1 10 9 13 7 16 10 0 0 9 10 0 9 4 1 9 2 2 3 4 15 9 3 15 9 1 4 2
21 10 9 4 3 16 10 9 1 15 2 0 0 2 13 3 1 0 9 0 4 2
23 15 4 15 4 1 10 9 1 11 2 7 15 13 15 0 4 16 10 9 1 10 9 2
12 1 10 9 1 11 4 10 15 9 1 4 2
59 8 13 0 9 3 4 2 16 1 8 10 9 1 15 4 4 2 7 1 10 9 1 10 0 9 1 10 9 1 10 9 2 3 8 3 3 9 13 2 13 15 10 0 9 10 4 16 15 1 10 9 1 10 9 1 10 11 13 2
42 3 3 2 8 2 10 9 1 15 8 7 0 0 3 15 0 9 2 13 10 9 1 10 9 1 10 9 3 0 9 4 2 16 15 10 9 1 9 1 13 4 2
27 7 10 9 1 8 2 3 3 3 0 1 11 9 2 13 1 10 0 9 4 4 4 16 11 3 13 2
17 10 9 5 3 15 1 10 0 9 5 4 3 3 3 0 4 2
22 1 12 9 1 10 9 11 4 3 1 8 10 9 1 10 9 11 2 11 2 4 2
21 10 9 13 0 1 10 9 2 3 10 0 9 13 2 7 13 3 1 15 9 2
26 10 9 2 10 0 9 8 2 2 12 0 7 13 2 1 11 2 13 15 8 15 9 1 9 4 2
25 10 9 13 3 16 10 9 15 1 12 1 11 4 4 7 15 1 12 1 11 13 4 2 13 2
11 15 4 3 1 15 12 0 10 9 4 2
24 10 9 1 11 2 15 15 10 13 9 16 2 9 2 13 4 2 13 15 3 0 8 4 2
13 10 9 13 3 10 9 2 10 9 1 12 9 2
36 16 10 9 15 9 1 1 10 9 13 4 16 3 0 1 10 0 9 1 13 2 13 15 10 9 3 1 10 9 2 15 1 10 9 13 2
28 10 9 13 3 9 1 10 12 9 2 15 15 1 9 1 10 9 13 4 7 1 9 1 15 9 13 4 2
24 15 13 1 9 1 9 4 15 9 7 15 13 3 4 16 15 3 0 0 1 10 9 13 2
51 15 13 3 10 9 7 10 9 7 15 9 8 2 7 15 13 1 11 7 11 7 15 13 10 9 9 1 15 1 10 9 7 3 13 15 3 3 13 2 16 3 1 15 0 9 10 9 4 4 2 2
14 3 2 3 1 10 9 2 13 15 12 9 1 11 2
14 7 3 13 3 10 9 10 0 9 4 1 10 11 2
8 0 9 8 10 9 12 9 2
8 0 2 10 9 13 9 4 2
19 15 13 3 3 1 10 9 1 9 10 0 9 2 7 10 9 13 3 2
21 10 9 15 15 3 10 9 13 4 1 9 7 15 3 15 15 15 13 2 13 2
10 15 13 9 2 9 2 9 2 9 2
27 10 9 13 10 9 3 16 3 3 3 12 9 9 1 4 4 2 7 15 13 10 9 3 1 15 8 2
20 1 9 8 1 10 11 1 11 4 3 1 12 10 0 9 1 10 9 4 2
10 8 3 13 4 4 4 3 15 4 2
30 1 10 1 9 13 9 13 15 12 9 9 2 15 1 10 9 1 10 9 1 15 9 2 1 0 9 2 4 4 2
9 10 9 4 1 15 9 3 4 2
13 0 2 15 4 4 1 10 9 2 13 10 9 2
22 1 11 4 10 9 4 2 15 15 8 13 9 3 1 4 16 10 9 1 10 9 2
22 10 9 4 4 1 10 0 9 7 9 2 8 2 15 1 12 1 11 13 7 13 2
45 9 4 10 9 1 15 9 2 15 2 0 2 13 1 10 9 1 12 9 2 7 10 15 0 4 1 2 10 0 7 13 9 2 1 9 2 15 1 11 9 13 4 1 9 2
63 15 13 3 8 4 1 10 9 1 10 0 9 2 1 10 9 1 9 7 15 9 2 15 15 1 3 0 9 13 2 1 10 9 1 9 2 1 10 9 1 9 2 7 3 1 10 9 1 9 2 1 10 0 9 2 3 15 9 7 9 3 13 2
12 7 15 13 3 1 10 0 9 9 16 4 2
14 1 10 9 1 9 2 9 7 9 13 15 4 4 2
10 15 4 13 1 10 9 1 10 9 2
24 10 9 1 15 1 15 8 13 9 1 0 7 9 4 10 0 9 16 16 9 1 4 4 2
15 1 15 9 13 15 8 11 2 11 2 11 7 11 13 2
11 2 1 11 13 15 3 8 12 12 4 2
13 3 13 15 3 3 9 16 1 10 9 1 4 2
13 15 4 3 10 9 13 7 15 4 9 0 8 2
25 15 9 13 8 10 9 1 11 7 11 1 11 0 3 1 10 9 1 11 16 1 15 1 11 2
13 8 13 1 9 12 9 3 7 11 4 8 0 2
15 11 13 12 9 7 0 4 3 0 8 2 11 7 11 2
11 6 2 15 13 15 9 2 9 7 9 2
8 3 13 8 12 9 1 3 2
13 10 0 9 4 1 10 9 15 0 16 1 9 2
48 10 9 1 15 9 16 11 10 9 1 10 9 1 9 4 2 13 1 10 13 9 15 13 9 2 16 4 15 9 4 1 15 1 10 9 13 1 11 2 15 10 9 1 10 9 11 13 2
30 1 12 9 4 10 9 1 11 0 1 4 2 7 10 9 1 11 13 12 9 0 10 9 16 10 9 1 10 9 2
15 10 0 9 1 11 4 1 15 3 3 0 8 3 15 2
4 2 12 2 2
17 8 13 3 1 15 15 9 11 10 9 4 1 10 0 13 9 2
20 11 13 9 3 1 10 9 1 12 9 15 3 10 0 9 13 1 10 9 2
20 10 9 13 1 10 9 3 1 10 9 1 8 2 15 10 9 3 3 13 2
10 1 10 9 4 15 3 0 1 8 2
4 1 9 3 2
14 0 0 1 15 9 4 8 2 15 10 0 9 13 2
21 3 8 13 1 10 9 8 15 9 3 3 2 16 13 15 9 10 9 0 8 2
10 10 9 13 1 3 0 9 1 11 2
26 8 13 15 9 16 9 2 16 3 1 10 9 2 11 1 10 0 9 13 7 10 0 0 9 13 2
46 10 13 9 13 3 15 2 9 2 1 10 9 2 15 10 9 8 1 10 0 9 13 7 10 9 1 9 1 10 0 9 11 2 15 1 10 9 1 12 9 3 0 0 4 4 2
8 10 9 13 15 3 3 0 2
32 8 1 10 2 0 2 9 2 8 1 10 0 9 1 10 9 1 10 9 1 10 9 2 15 1 10 0 9 13 4 4 2
35 1 9 1 9 10 13 9 13 10 9 1 11 15 1 15 9 1 10 11 12 0 9 2 12 8 2 10 9 7 10 0 9 4 4 2
25 10 3 13 9 13 0 16 10 9 7 10 9 1 10 0 9 10 9 7 10 9 4 4 4 2
23 10 9 13 1 10 9 1 15 9 3 7 15 4 1 10 9 1 10 9 1 10 9 2
18 3 13 15 3 3 1 10 9 1 4 2 1 13 2 3 1 13 2
20 8 2 9 1 10 9 1 15 8 2 13 0 16 9 3 1 4 1 8 2
15 15 9 4 4 1 10 9 1 10 9 1 10 9 8 2
30 8 13 3 16 10 0 0 9 1 10 12 9 1 15 9 15 15 9 1 9 4 4 1 15 0 13 1 15 9 2
26 10 9 13 16 0 7 13 0 9 1 0 9 4 4 1 10 0 9 7 15 13 1 10 0 9 2
7 1 12 9 4 15 13 2
8 15 13 10 9 3 3 4 2
9 10 9 13 1 13 9 1 3 2
13 10 9 1 10 9 4 3 4 2 13 9 11 2
23 10 9 13 3 1 10 9 1 11 1 10 9 11 3 2 3 15 1 13 9 4 4 2
15 13 1 9 2 7 15 4 1 10 9 1 10 9 4 2
10 15 13 15 15 9 3 3 3 2 2
18 1 9 11 2 2 15 4 15 9 0 2 2 4 15 10 0 9 2
15 8 1 11 13 11 1 9 1 8 7 1 9 1 8 2
10 8 13 1 11 10 9 1 9 8 2
29 10 9 1 10 9 1 10 9 4 3 0 2 16 3 3 0 9 1 15 8 1 11 13 16 10 9 8 13 2
15 3 1 10 0 9 1 15 8 4 3 10 9 3 13 2
8 11 13 3 3 10 0 9 2
11 9 4 3 0 0 1 10 9 7 9 2
15 15 4 9 2 15 1 15 13 9 4 4 1 15 9 2
12 15 13 16 9 1 9 7 3 9 1 9 2
10 1 10 9 13 15 9 0 16 9 2
20 9 8 2 15 15 1 8 3 0 1 11 13 0 2 13 3 1 10 9 2
15 15 4 15 3 1 10 0 9 4 2 7 13 15 9 2
15 3 13 3 9 13 1 10 9 1 10 9 15 15 13 2
9 15 13 9 2 9 2 3 4 2
35 10 9 1 15 9 13 3 15 3 16 3 15 15 3 1 15 9 1 15 9 4 4 2 16 15 5 1 15 9 13 5 1 3 13 2
5 15 13 0 4 2
25 4 15 0 2 3 13 15 2 16 10 9 11 1 15 9 10 3 0 9 13 4 1 15 9 2
4 9 11 13 2
21 15 13 8 1 15 9 13 15 2 15 13 3 10 0 9 1 10 0 9 9 2
11 12 0 9 13 15 9 1 9 1 11 2
14 15 13 10 9 4 15 3 1 10 9 11 4 4 2
21 2 15 4 9 15 3 4 4 2 2 13 15 2 2 15 4 3 0 1 11 2
10 9 7 9 4 1 0 12 9 4 2
16 15 1 10 9 13 3 9 1 15 13 7 13 1 15 9 2
22 15 4 8 2 15 0 9 8 13 2 16 15 3 1 8 1 10 9 1 11 13 2
13 10 0 9 8 1 11 4 3 1 9 8 4 2
21 10 9 13 1 4 1 10 9 1 10 9 8 2 15 1 10 11 1 11 13 2
16 10 9 1 10 9 4 13 4 2 3 10 9 13 1 4 2
21 16 9 8 3 16 15 13 15 9 13 2 13 15 15 9 1 10 9 0 9 2
5 10 9 4 4 2
21 9 8 2 15 9 1 2 8 2 1 11 2 13 3 15 0 9 1 15 4 2
19 15 13 15 0 9 1 11 16 2 3 13 15 3 2 15 9 1 13 2
10 0 13 3 3 3 9 1 10 9 2
11 1 12 13 10 9 1 9 1 15 8 2
13 3 13 10 11 1 10 9 10 0 9 1 4 2
17 3 13 10 9 2 15 3 1 10 9 4 4 2 10 0 9 2
24 12 9 4 4 1 9 1 10 0 9 1 10 13 9 2 3 9 1 0 9 1 9 13 2
4 15 12 4 2
20 11 2 11 2 11 2 8 2 9 2 8 2 11 2 11 2 11 7 11 2
15 8 12 13 15 0 9 4 2 3 15 12 9 13 4 2
10 3 13 4 4 16 10 9 0 4 2
20 10 9 13 4 4 1 10 9 2 15 1 10 0 12 9 1 10 9 13 2
9 3 13 10 0 9 1 9 11 2
17 15 4 3 0 1 15 0 9 2 7 9 4 3 0 3 4 2
16 15 13 8 11 1 4 1 10 9 1 10 11 1 10 11 2
10 15 13 10 9 4 1 0 0 9 2
39 15 15 15 13 4 1 10 9 13 1 9 9 4 2 7 10 9 4 3 4 1 10 9 2 3 15 13 10 2 0 9 2 1 10 9 13 4 4 2
11 11 13 3 0 9 4 1 10 9 2 2
27 3 13 3 10 0 9 9 2 3 3 3 3 3 15 13 7 5 16 15 0 3 3 13 5 15 13 2
23 15 13 3 3 15 4 4 2 16 13 15 4 2 16 10 0 13 9 3 13 4 4 2
6 3 15 0 2 6 2
43 16 15 3 3 10 0 9 4 2 13 15 13 1 15 9 15 3 4 4 2 7 0 1 10 9 13 10 9 3 10 0 2 16 3 1 13 2 0 9 1 15 9 2
24 10 0 9 8 13 10 9 1 0 9 4 10 9 3 1 4 1 9 8 1 10 0 9 2
26 10 9 11 13 10 9 3 2 15 0 8 1 11 1 9 1 15 9 1 10 0 9 1 4 4 2
35 10 0 9 15 10 9 13 4 16 15 9 1 4 1 10 9 1 10 9 1 10 9 4 10 0 9 1 10 9 1 0 9 7 9 2
18 3 4 15 3 3 13 2 16 10 9 1 11 15 3 9 13 4 2
21 8 4 1 10 9 8 4 2 16 15 3 0 9 13 2 16 15 10 9 4 2
7 15 13 10 9 15 4 2
13 0 1 0 9 2 0 1 0 9 2 3 0 2
24 3 0 10 9 1 15 0 9 13 4 4 2 13 15 0 13 9 9 3 9 0 9 13 2
25 15 13 3 5 16 0 5 3 7 13 3 3 0 2 16 0 2 7 3 0 2 1 10 9 2
32 15 13 1 15 0 9 9 2 7 15 13 15 4 2 15 13 3 10 15 16 10 9 2 7 9 2 3 15 8 9 13 2
16 7 15 9 5 15 13 3 12 5 13 3 1 10 9 4 2
7 15 4 8 1 15 9 2
9 0 11 13 10 0 9 15 4 2
3 9 11 2
14 1 10 9 15 4 10 0 9 3 8 2 1 4 2
8 15 13 3 3 15 12 3 2
6 7 15 4 3 0 2
18 8 13 15 15 0 1 10 9 3 2 3 0 15 15 9 3 7 2
15 3 4 9 4 2 0 9 2 9 2 9 7 0 9 2
11 3 4 4 0 9 7 9 1 4 4 2
15 10 9 13 0 3 1 4 1 9 1 10 9 1 9 2
15 1 10 9 13 10 0 9 9 7 9 0 1 4 4 2
20 10 9 13 3 2 16 10 9 10 9 1 10 9 1 10 9 1 13 4 2
10 4 4 10 9 9 3 1 4 1 2
9 9 2 9 2 9 2 9 9 2
28 10 0 9 1 11 13 15 2 16 15 8 1 10 0 9 1 9 8 13 4 2 3 0 4 1 10 9 2
13 1 8 13 10 0 9 8 1 10 9 10 9 2
4 10 9 13 2
13 10 9 13 10 9 4 2 3 10 9 13 4 2
23 10 9 13 10 9 1 12 9 7 13 9 1 10 9 1 10 9 7 10 9 1 4 2
21 9 8 1 15 8 13 3 9 4 10 9 1 10 9 1 10 9 11 1 4 2
6 15 13 10 9 3 2
13 1 11 13 15 9 4 1 9 16 9 1 9 2
25 12 0 9 13 3 4 4 7 1 10 9 1 10 9 13 15 12 9 4 1 15 13 1 9 2
15 3 2 3 13 8 2 4 4 1 10 9 1 10 9 2
22 9 13 15 0 9 16 9 7 9 7 15 8 13 1 10 9 3 13 1 10 9 2
7 10 9 13 15 3 0 2
32 15 13 9 1 10 9 1 10 9 2 15 4 4 1 10 9 16 3 10 9 1 13 2 3 15 13 15 9 1 4 4 2
7 15 9 4 1 9 4 2
20 1 10 9 1 10 9 4 15 2 16 15 9 4 4 1 9 7 9 3 2
14 3 4 10 9 1 15 9 1 10 9 1 4 4 2
23 10 12 9 0 2 1 9 7 9 13 9 1 10 0 9 8 4 3 0 4 1 11 2
28 10 9 4 8 7 4 10 9 1 10 9 11 1 15 9 2 13 8 10 9 1 10 0 9 1 15 8 2
25 8 2 15 1 10 9 1 10 9 9 13 2 13 1 11 1 15 9 2 15 0 1 3 1 2
6 15 13 15 1 8 2
41 10 9 8 13 10 0 9 1 10 10 0 12 9 13 13 9 0 1 9 7 13 3 10 9 3 16 10 9 1 11 3 3 3 0 0 1 10 9 4 4 2
13 10 9 0 13 0 1 10 12 9 1 10 9 2
16 1 10 9 1 10 9 4 3 10 12 0 12 9 0 4 2
10 15 13 1 15 9 1 10 9 9 2
6 8 13 10 9 15 2
7 2 9 4 3 3 9 2
7 10 0 13 3 9 2 2
16 3 0 7 0 4 3 10 0 9 16 9 3 15 3 13 2
10 10 0 9 16 15 0 9 1 4 2
13 1 8 4 3 9 1 4 1 8 1 10 11 2
20 15 4 3 0 7 0 4 7 3 13 9 2 9 7 0 9 3 8 4 2
16 15 13 1 9 1 0 9 7 3 13 3 10 0 9 3 2
28 2 15 13 16 3 1 10 0 9 10 9 1 9 4 2 7 3 13 15 15 9 1 10 0 9 8 2 2
13 10 0 9 13 3 1 12 1 0 9 11 12 2
24 10 0 9 8 1 11 13 3 1 15 9 1 10 9 1 10 0 9 2 8 2 15 9 2
20 15 13 3 16 15 1 12 0 9 0 15 9 1 10 11 1 11 8 13 2
10 8 13 10 9 1 11 1 12 4 2
12 15 4 10 0 9 1 12 9 1 10 11 2
23 10 9 1 10 0 9 1 9 2 8 4 3 3 1 10 9 4 1 10 9 1 11 2
19 15 4 10 12 9 2 15 15 4 1 11 16 15 1 4 1 10 9 2
11 10 0 9 1 12 9 4 1 12 4 2
10 15 13 15 3 3 1 8 3 4 2
4 9 15 9 2
6 2 6 2 13 11 2
8 1 10 0 9 4 12 4 2
5 2 15 13 0 2
27 2 15 4 9 1 10 9 7 15 9 4 3 3 3 0 1 13 2 16 15 15 9 13 16 1 4 2
18 15 13 8 1 10 9 0 3 12 9 4 7 3 4 15 3 4 2
15 3 13 15 0 4 7 8 3 3 10 0 9 4 4 2
25 1 12 13 15 10 9 3 2 3 10 0 9 7 9 1 10 9 16 9 1 10 9 4 4 2
27 1 10 9 4 3 1 10 9 1 11 4 2 7 1 10 0 9 13 10 9 1 12 10 9 3 4 2
15 1 9 1 10 9 13 10 9 1 10 9 15 9 4 2
16 1 10 9 3 4 15 1 11 4 2 3 16 15 1 13 2
37 10 9 15 1 10 9 3 9 7 3 9 1 9 3 13 4 13 1 10 9 16 10 9 3 9 4 4 4 1 15 0 2 0 7 0 9 2
6 9 3 4 3 15 2
5 10 9 4 0 2
36 8 2 9 1 10 9 1 11 7 11 13 16 1 9 7 9 10 0 9 0 4 4 4 2 3 16 10 0 9 1 9 7 9 8 13 2
10 10 9 8 13 16 9 1 15 9 2
19 15 13 15 9 10 13 9 1 3 12 9 4 7 3 10 9 3 13 2
32 10 9 13 3 10 9 4 1 0 1 13 16 0 9 1 10 9 2 1 10 9 15 13 2 3 1 10 9 4 4 4 2
8 8 13 10 9 1 9 4 2
9 3 4 1 15 9 0 9 8 2
14 15 13 3 15 12 9 2 12 9 2 0 1 9 2
29 15 13 0 3 4 4 16 15 12 9 3 13 16 1 3 1 13 7 16 15 3 3 3 15 9 3 13 2 2
5 10 9 4 0 2
22 9 13 15 3 3 2 10 9 13 3 15 2 7 10 9 4 3 0 1 15 9 2
15 0 13 10 9 3 8 9 15 3 1 0 12 7 12 2
7 12 9 7 15 9 3 2
21 2 15 13 2 13 15 3 2 2 10 0 9 4 1 10 9 7 9 1 11 2
33 9 1 12 13 8 1 15 9 2 13 1 10 9 0 9 2 1 10 9 1 10 9 2 8 2 2 9 1 15 3 13 9 2
3 15 13 2
12 2 1 15 13 15 15 9 1 12 4 2 2
8 8 4 0 1 10 0 9 2
27 2 15 4 0 2 13 15 0 3 4 4 2 7 13 15 4 16 15 9 0 3 15 0 9 4 2 2
33 10 9 13 3 2 16 3 1 9 12 0 9 1 10 2 13 9 2 4 4 4 2 16 15 12 0 12 9 1 3 1 9 2
14 10 9 2 8 2 2 15 3 9 13 4 2 13 2
26 1 10 0 9 13 8 1 10 2 1 15 9 1 11 2 9 1 10 9 1 9 1 12 7 12 2
8 3 10 0 9 4 0 13 2
27 1 10 0 9 2 7 3 0 13 2 13 10 9 1 12 4 2 10 9 2 13 9 2 3 1 4 2
15 10 0 9 8 13 9 1 15 9 1 10 9 1 11 2
19 15 0 9 13 0 0 10 9 1 15 12 9 2 12 12 9 2 4 2
31 1 10 9 11 13 10 9 3 10 9 4 1 10 9 1 9 11 2 3 15 15 9 13 16 2 0 15 1 4 2 2
12 15 13 16 15 13 4 7 15 0 0 4 2
16 10 9 13 3 1 12 3 0 9 4 1 10 0 0 9 2
23 10 9 2 15 10 11 1 13 9 13 2 13 12 9 2 7 10 9 4 3 10 9 2
18 15 13 16 10 9 15 9 2 1 9 3 2 2 1 12 9 4 2
16 10 0 9 1 10 9 13 1 12 12 3 1 12 12 9 2
20 3 13 10 9 2 8 2 3 1 15 9 1 10 9 12 15 0 9 4 2
30 15 13 3 2 16 2 16 3 10 9 15 8 13 2 3 15 0 13 4 2 1 15 15 9 10 9 0 0 4 2
15 10 9 1 9 4 4 1 10 0 9 8 2 12 2 2
14 10 9 1 10 9 4 10 9 15 0 9 1 13 2
48 10 9 13 4 16 15 4 2 3 13 10 3 0 9 3 2 1 10 9 4 10 3 13 9 4 2 15 8 13 2 16 15 10 9 2 15 3 0 13 4 2 1 10 9 4 4 4 2
11 7 15 13 10 9 1 9 1 12 9 2
38 15 13 3 2 16 10 0 9 2 10 16 12 9 2 4 1 10 2 0 9 2 2 15 1 15 0 9 15 9 10 9 13 4 1 10 15 9 2
24 2 7 15 2 2 3 11 2 2 13 15 15 9 2 7 9 7 15 4 15 3 3 2 2
23 15 13 16 10 9 1 10 0 9 0 10 9 10 9 4 16 15 9 0 3 1 4 2
14 8 1 11 4 3 1 11 13 9 1 11 9 4 2
34 10 9 3 4 2 16 8 1 11 2 15 15 9 0 0 8 13 2 16 15 0 3 1 13 4 10 0 9 3 1 9 4 4 2
21 1 11 2 3 3 10 2 13 9 2 13 2 13 15 9 1 10 0 9 3 2
15 15 13 3 0 16 10 0 9 1 8 7 8 1 11 2
16 15 13 10 9 2 8 2 1 15 0 9 8 2 12 2 2
13 13 10 13 9 1 10 0 9 1 11 15 9 2
16 16 6 2 4 10 9 1 10 0 13 9 1 11 0 13 2
13 9 2 15 1 10 9 3 3 0 1 4 4 2
30 3 3 2 16 10 9 1 11 13 16 10 9 3 1 4 1 10 9 2 15 15 9 8 10 9 0 13 2 8 2
18 10 9 1 11 4 3 0 1 10 1 10 9 13 9 1 15 9 2
18 3 13 3 16 10 9 3 0 4 10 9 1 8 1 9 1 4 2
14 3 13 10 9 9 1 10 11 1 15 1 13 13 2
4 10 9 13 2
23 15 10 9 8 1 10 0 9 13 2 4 16 15 3 1 15 9 10 13 9 13 4 2
26 9 13 3 3 3 1 10 9 1 10 0 0 9 8 2 15 9 1 10 9 1 15 9 4 4 2
18 15 0 9 1 9 13 1 12 1 9 8 1 11 1 11 4 4 2
37 10 0 9 8 15 1 10 9 1 10 9 1 10 9 1 15 8 10 9 8 13 7 13 2 4 9 1 12 8 1 10 9 1 15 9 4 2
9 10 9 4 1 10 9 8 4 2
20 8 13 1 15 8 4 5 8 8 10 0 9 5 10 9 1 11 1 4 2
33 10 9 1 15 8 13 15 10 9 4 1 10 9 1 10 9 2 3 15 10 9 13 9 3 13 4 7 15 15 15 9 13 2
28 15 13 1 15 9 3 1 10 9 2 15 11 1 11 1 10 9 1 10 11 4 4 1 9 1 10 9 2
36 10 9 1 15 8 7 15 12 9 8 7 8 1 10 0 11 13 1 10 9 15 0 9 4 2 3 13 10 9 1 9 1 11 4 4 2
17 1 10 9 13 10 12 9 4 4 1 10 9 1 10 0 9 2
14 10 9 1 9 13 1 10 9 10 9 1 10 9 2
10 1 11 7 10 9 13 3 12 9 2
10 15 13 3 9 1 10 9 1 9 2
30 10 12 9 4 4 1 10 9 1 12 9 1 15 0 9 8 9 2 9 1 0 9 1 10 9 1 0 9 2 2
30 11 8 1 10 9 1 10 11 13 12 9 4 15 13 1 9 2 3 9 7 15 9 13 2 8 10 9 1 4 2
7 10 2 9 2 4 4 2
17 15 13 3 1 9 1 10 0 0 9 1 12 1 3 12 9 2
20 10 13 9 13 1 15 9 3 1 10 9 3 7 4 0 1 10 9 4 2
19 10 15 12 9 0 9 8 1 11 4 1 10 9 1 11 1 11 4 2
9 1 10 9 4 10 0 9 13 2
16 1 10 9 1 10 9 4 10 9 7 9 4 1 15 8 2
11 1 10 9 13 10 0 9 8 0 9 2
7 1 15 15 4 15 3 2
10 10 9 8 13 1 15 13 15 4 2
35 15 13 3 2 16 10 9 1 15 9 10 9 13 4 2 3 13 15 0 9 15 3 10 9 9 3 4 2 3 3 8 3 4 2 2
18 1 10 11 1 11 4 1 10 9 1 11 1 11 4 10 9 8 2
27 15 4 0 1 9 16 9 1 11 7 1 10 9 16 9 1 10 9 11 7 16 0 9 1 15 8 2
6 8 4 12 9 4 2
32 15 9 13 3 0 9 15 8 3 2 16 15 15 3 13 4 7 15 0 9 3 9 13 4 1 10 9 1 10 9 11 2
31 1 10 9 15 1 10 9 1 11 13 13 1 15 9 10 9 1 10 9 16 15 9 7 9 1 10 9 3 1 13 2
10 15 16 15 13 1 10 9 1 13 2
8 8 4 15 10 0 9 4 2
14 11 13 1 10 12 13 9 3 10 0 0 9 3 2
10 10 0 9 13 10 13 9 1 4 2
9 1 10 0 9 4 11 0 8 2
14 10 0 13 1 3 10 9 1 10 9 1 10 9 2
15 10 9 13 10 9 15 9 1 10 0 9 1 4 4 2
13 3 1 9 4 15 3 12 2 3 8 9 11 2
9 1 10 0 9 4 11 0 0 2
13 10 9 4 15 8 2 3 16 0 3 1 13 2
16 0 13 8 1 9 15 0 9 7 4 11 13 16 9 4 2
28 1 10 9 4 9 11 0 2 7 10 9 1 10 9 13 3 3 15 9 3 4 2 16 10 9 0 4 2
25 11 13 11 1 0 9 2 12 2 7 11 13 1 15 9 3 3 3 9 1 11 2 12 2 2
7 8 13 1 12 0 3 2
12 8 13 4 1 10 9 1 10 9 1 9 2
33 8 2 1 0 9 1 12 8 12 11 2 13 4 4 1 9 1 12 9 2 16 13 9 3 2 3 4 11 1 10 9 4 2
9 9 13 15 0 9 1 15 9 2
10 12 9 13 3 10 9 1 15 4 2
29 10 9 1 10 11 13 15 11 3 4 1 10 9 9 2 16 10 9 3 4 4 1 9 7 9 1 10 9 2
22 2 15 13 3 3 0 9 1 10 9 1 10 9 2 2 13 10 9 1 10 9 2
19 2 8 13 15 3 4 7 3 13 15 15 1 10 9 1 9 8 4 2
16 15 13 1 9 13 15 0 3 4 16 15 13 1 9 2 2
22 12 1 10 9 13 10 13 9 3 1 10 9 16 15 3 3 3 1 10 9 4 2
13 3 8 2 15 8 13 1 10 9 1 12 3 2
25 16 12 2 0 9 2 13 8 2 8 2 8 2 8 2 8 2 8 7 8 1 10 9 4 2
29 15 13 9 4 8 9 2 9 7 9 2 15 9 8 10 9 2 9 2 9 7 9 1 10 13 9 13 4 2
13 15 8 4 1 10 9 2 11 2 1 11 4 2
9 1 9 1 9 13 15 1 4 2
8 12 9 13 2 3 2 4 2
6 8 2 8 7 8 2
18 3 4 8 2 12 2 10 13 9 1 10 9 1 15 8 1 11 2
11 15 4 10 0 9 1 10 0 9 12 2
29 7 3 13 15 16 0 0 9 12 9 1 11 2 3 12 9 1 15 9 1 10 9 4 4 1 9 7 9 2
5 3 13 11 9 2
16 2 15 13 15 9 4 16 15 9 10 0 9 4 4 2 2
12 11 13 1 15 9 10 9 2 1 9 2 2
32 10 0 9 1 15 8 13 15 9 2 9 7 10 9 10 9 16 15 15 9 3 13 9 4 4 1 10 9 1 10 9 2
8 2 16 15 0 9 4 4 2
20 15 13 10 9 15 15 0 13 2 3 3 13 15 10 9 4 2 1 4 2
32 3 10 9 15 0 1 10 9 7 10 0 12 9 4 4 8 1 10 0 15 9 2 13 15 15 3 2 2 3 10 9 2
15 10 0 9 1 10 9 13 1 15 9 4 1 0 9 2
25 10 11 4 1 10 9 1 15 9 3 3 0 4 2 16 10 0 9 15 1 10 9 13 4 2
20 7 8 9 13 10 9 8 2 15 1 10 9 1 11 1 15 9 4 4 2
13 15 13 15 9 10 0 9 10 9 3 1 13 2
4 15 13 3 2
4 0 7 3 2
13 15 13 1 15 9 12 3 3 3 3 3 3 2
6 15 13 11 1 11 2
22 1 10 9 7 13 3 1 10 9 2 13 13 15 0 0 4 4 2 0 15 9 2
13 6 2 15 4 10 9 1 15 9 10 9 0 2
18 1 11 13 15 0 2 16 11 0 4 10 11 1 4 1 11 2 2
24 9 8 4 3 15 3 0 2 16 10 0 12 0 15 3 1 11 13 2 15 8 4 4 2
26 15 13 15 1 15 0 9 9 4 2 10 0 9 3 1 4 7 3 9 3 1 4 1 15 9 2
4 3 10 9 2
8 7 15 13 1 10 9 2 2
7 15 4 10 9 2 6 2
2 8 2
21 2 16 15 1 9 1 10 13 9 13 2 13 15 9 2 15 13 15 3 3 2
17 7 15 13 3 16 9 3 4 2 16 10 9 1 15 9 4 2
21 15 4 0 1 10 9 7 10 9 2 15 13 4 2 16 3 3 4 4 2 2
22 9 7 9 4 3 10 0 9 3 1 10 9 10 0 9 13 2 13 1 0 9 2
39 10 9 4 16 15 9 0 1 13 16 15 3 0 4 4 16 1 10 11 1 13 4 16 16 3 3 4 1 4 15 9 1 2 8 2 1 4 4 2
4 10 0 9 2
18 15 1 10 9 4 15 0 13 2 16 11 3 13 1 10 9 11 2
7 7 10 9 4 3 0 2
12 15 8 1 11 13 1 12 9 15 0 13 2
7 15 9 4 0 7 13 2
10 15 1 15 9 13 15 15 0 9 2
7 3 3 4 10 9 0 2
24 8 3 13 10 9 7 10 9 2 13 1 8 7 8 2 7 1 2 11 2 3 10 9 2
22 3 4 10 11 3 0 8 1 10 9 1 10 9 1 9 2 11 7 15 0 9 2
21 11 13 0 10 9 2 15 11 5 0 0 16 9 1 4 5 1 10 9 13 2
18 6 2 15 13 16 15 0 12 9 11 4 16 12 9 11 1 11 2
29 10 12 9 0 13 9 13 15 3 7 10 13 9 13 10 9 8 4 15 3 1 11 7 10 9 4 4 2 2
13 3 4 10 9 0 15 16 3 1 9 1 13 2
19 12 0 9 13 15 1 15 9 1 0 3 1 11 3 10 9 4 4 2
17 2 11 2 13 15 1 12 0 9 2 10 9 1 10 12 9 2
29 1 10 0 13 12 9 10 9 3 8 16 15 12 4 2 0 9 2 12 9 2 13 15 3 1 9 1 12 2
10 15 0 9 4 0 1 9 11 4 2
23 9 8 2 15 12 9 3 1 10 9 1 15 0 7 0 9 1 11 13 4 2 13 2
7 2 11 13 9 1 4 2
19 1 15 9 1 10 9 13 15 0 8 10 9 8 11 3 1 4 2 2
14 1 11 13 9 1 11 4 16 11 9 4 1 11 2
21 15 0 8 2 1 12 12 7 12 11 1 10 11 2 13 3 15 9 1 4 2
26 10 9 3 9 8 13 1 10 9 1 15 9 8 2 13 1 12 0 2 13 9 8 10 0 9 2
27 1 10 0 9 1 10 9 11 2 1 12 0 2 13 15 9 8 15 9 1 11 1 15 1 10 9 2
37 15 13 15 1 15 0 9 1 11 0 3 4 1 4 1 0 9 2 16 15 0 9 1 10 9 0 4 1 9 7 16 10 9 10 9 4 2
23 0 4 16 10 9 11 3 10 9 8 13 15 10 9 1 12 9 1 10 11 13 4 2
18 1 15 9 13 15 16 12 0 9 8 15 9 3 10 0 9 2 2
17 1 10 9 1 11 13 15 1 10 9 1 10 11 1 12 9 2
15 15 13 1 12 9 1 10 11 2 3 0 1 12 9 2
12 11 4 4 16 9 1 0 7 3 0 9 2
9 7 3 13 11 2 11 7 8 2
22 15 13 10 9 4 15 1 10 9 1 10 11 13 7 10 9 13 9 7 9 4 2
18 3 0 4 10 9 3 4 10 15 0 9 1 15 1 4 15 9 2
13 3 13 1 11 7 11 1 12 9 1 15 9 2
6 15 13 3 3 15 2
16 15 4 3 0 2 16 0 9 3 3 9 13 4 16 9 2
16 15 13 3 3 1 15 9 1 10 13 7 13 9 9 4 2
35 2 10 9 15 8 13 4 2 2 3 13 8 1 15 1 10 0 9 2 8 2 2 2 10 0 9 1 9 2 0 1 0 9 2 2
22 10 0 11 4 4 1 10 0 9 8 2 12 2 15 1 0 3 2 8 2 13 2
6 2 3 15 9 2 2
40 11 4 1 9 3 0 7 0 2 7 8 15 9 13 15 3 15 10 9 4 1 10 0 0 9 2 3 2 8 2 1 10 0 9 2 1 15 9 13 2
22 8 2 12 2 10 0 9 2 13 1 10 3 1 10 9 11 13 9 15 9 4 2
32 15 0 16 10 13 9 1 8 2 15 15 1 10 0 9 13 2 13 3 10 9 3 2 15 10 9 1 0 9 13 4 2
31 10 0 1 10 9 2 15 1 15 15 8 1 10 15 13 2 13 1 10 11 10 0 9 4 1 10 9 1 0 9 2
17 15 13 15 3 16 15 15 1 0 13 1 10 9 4 4 4 2
16 1 10 0 9 15 1 10 9 4 4 2 4 11 10 9 2
9 15 4 10 9 9 1 13 9 2
24 16 15 1 10 11 2 3 11 2 4 4 2 13 15 12 9 2 15 1 10 9 4 4 2
10 8 13 15 9 4 16 15 9 4 2
15 1 10 9 12 9 1 10 11 4 10 9 4 7 4 2
7 1 10 9 13 10 11 2
14 2 15 4 3 8 1 11 7 10 9 1 0 9 2
11 1 15 8 13 15 3 15 9 4 2 2
21 3 10 9 1 10 9 1 11 2 8 1 10 9 2 16 15 3 1 11 13 2
15 16 10 0 9 15 9 4 4 2 13 1 10 0 9 2
22 15 13 10 15 9 1 10 15 7 13 3 10 9 1 8 2 10 9 1 10 11 2
22 10 9 1 15 9 2 15 13 4 1 10 9 7 9 1 10 9 9 13 3 0 2
15 11 7 11 13 4 2 8 1 10 9 1 10 12 9 2
22 15 13 1 11 10 9 4 1 10 9 1 9 2 10 9 1 7 0 7 0 9 2
25 9 4 4 1 9 1 10 9 7 10 9 1 10 9 2 1 9 2 1 9 7 1 10 9 2
19 15 4 2 3 3 10 9 1 11 1 11 2 15 1 10 0 13 9 2
22 2 15 13 15 1 10 9 11 8 4 2 13 10 9 1 10 9 11 1 15 9 2
35 10 9 1 9 4 1 8 1 10 9 4 2 16 10 9 2 10 11 7 10 11 2 3 10 11 9 13 2 15 9 2 3 2 4 2
17 10 9 13 10 11 15 9 7 10 9 3 1 4 1 10 9 2
31 15 9 13 1 15 9 12 9 3 15 12 9 4 2 15 13 1 12 9 1 10 9 2 7 15 13 15 9 1 9 2
22 1 10 0 0 7 0 9 1 10 9 7 10 9 13 3 10 13 9 1 10 9 2
17 11 7 3 3 10 15 9 2 8 2 13 9 1 0 9 3 2
28 15 13 3 1 9 1 9 2 16 10 0 9 1 10 9 10 9 1 10 11 2 3 3 9 13 4 2 2
12 15 9 3 2 13 15 12 9 4 1 9 2
29 9 8 2 3 2 2 15 1 9 15 9 1 10 0 9 8 13 4 2 4 4 1 10 1 15 8 0 9 2
12 15 9 8 2 3 2 2 13 15 1 4 2
12 3 13 13 10 0 9 8 1 10 0 9 2
8 1 10 0 9 13 15 0 2
13 2 3 4 4 1 9 7 9 1 0 9 2 2
24 3 13 15 3 4 2 16 15 10 0 9 4 2 10 9 9 15 3 1 3 1 9 0 2
9 15 13 15 3 2 4 10 9 2
19 15 8 13 0 1 10 9 1 10 9 1 12 1 12 1 10 13 9 2
56 10 0 9 2 15 15 1 15 13 2 4 10 9 2 3 10 13 2 9 2 9 2 9 2 15 3 0 3 3 3 7 3 0 1 0 9 0 4 2 16 10 9 7 10 9 15 3 2 8 13 2 1 10 0 9 2
21 11 2 15 9 13 2 13 3 2 16 15 9 2 10 9 10 9 2 4 4 2
5 11 4 15 9 2
15 10 11 13 15 10 9 1 10 9 1 10 0 9 8 2
25 8 13 10 0 9 4 1 2 11 13 1 11 2 10 0 9 8 15 12 9 0 9 13 4 2
27 11 13 2 16 15 0 4 4 1 9 7 16 15 9 4 4 2 3 15 15 4 13 1 10 0 9 2
26 1 12 9 0 1 10 9 1 13 4 4 10 0 9 8 3 1 10 9 1 10 0 9 11 4 2
17 1 10 9 1 11 13 15 10 0 9 15 11 1 9 13 4 2
23 8 4 1 12 1 11 1 10 0 9 4 1 9 2 16 15 8 13 4 0 1 4 2
18 15 2 9 2 4 15 0 8 15 15 16 9 1 15 9 13 4 2
32 9 8 2 9 2 4 7 1 10 11 7 1 10 11 1 9 4 10 9 9 1 9 1 12 1 15 9 1 4 1 12 2
26 10 9 11 2 9 1 15 8 1 11 2 13 15 12 9 2 16 1 9 1 13 2 15 0 4 2
10 9 13 1 15 9 0 1 9 4 2
16 1 15 8 13 15 2 15 1 10 9 0 9 4 4 4 2
37 1 10 9 11 13 15 8 2 16 10 11 2 3 11 4 4 2 15 9 13 16 15 1 10 9 1 10 9 7 9 2 1 9 2 1 13 2
34 10 0 9 13 4 2 16 1 10 9 1 9 8 2 3 0 9 10 0 9 8 13 4 4 2 3 10 9 7 10 9 4 4 2
9 15 13 1 10 9 1 10 9 2
20 3 0 4 1 10 9 1 9 11 10 9 2 10 9 7 10 0 9 4 2
15 10 9 13 3 3 8 1 10 9 1 10 9 13 9 2
16 10 9 1 10 9 16 10 9 1 11 13 15 15 9 3 2
5 11 13 0 8 2
18 15 9 5 8 10 11 5 13 15 0 9 1 10 9 1 10 9 2
19 11 13 3 0 7 3 3 0 4 2 3 16 1 0 0 9 1 13 2
21 10 9 4 15 0 4 16 1 13 16 11 4 2 16 16 1 13 16 11 4 2
20 10 0 0 9 2 13 10 9 1 12 2 4 3 3 10 9 1 10 9 2
26 3 10 9 1 15 8 13 3 1 0 9 4 9 1 4 16 3 1 13 1 10 9 1 9 11 2
16 1 10 9 1 10 9 13 10 2 9 2 10 3 13 9 2
28 3 4 15 1 10 9 16 10 10 9 2 10 9 0 2 13 4 2 8 1 4 4 2 15 10 9 4 2
25 10 9 10 9 13 3 3 10 9 1 9 2 2 1 10 9 2 4 7 4 3 10 9 9 2
23 10 9 2 15 0 2 4 1 15 9 3 3 4 16 10 9 1 10 9 4 1 13 2
19 3 4 10 9 1 10 9 1 10 13 9 1 15 9 3 0 0 4 2
22 15 13 5 8 5 16 10 9 1 9 1 9 7 1 10 15 9 0 1 10 9 2
4 3 13 15 2
24 3 13 1 15 8 10 9 1 11 4 4 16 1 13 1 9 2 9 7 9 1 10 9 2
24 3 13 10 0 9 1 11 2 3 15 0 8 0 9 4 2 7 1 11 1 11 9 4 2
11 13 15 15 9 3 3 1 15 9 4 2
15 10 0 9 13 3 1 10 9 3 10 0 2 0 9 2
17 1 10 9 1 9 4 3 7 1 10 9 7 1 10 9 4 2
15 15 10 0 9 1 10 8 2 11 2 11 4 8 4 2
23 1 12 2 16 10 9 11 1 15 8 4 4 2 13 10 11 10 9 4 1 15 8 2
24 10 13 9 13 3 10 9 4 1 10 9 1 9 11 16 10 0 9 1 11 0 1 4 2
13 15 9 4 4 1 15 1 11 13 2 12 2 2
9 15 8 1 11 13 10 11 4 2
10 1 11 7 11 4 3 3 3 4 2
10 8 1 10 9 1 10 9 13 15 2
15 7 1 10 0 9 1 3 8 13 15 3 1 9 2 2
13 10 9 11 13 10 9 1 10 9 1 9 4 2
22 2 10 10 9 13 2 3 13 15 3 4 4 2 7 15 4 13 1 10 9 2 2
7 10 9 11 13 15 3 2
11 2 10 0 1 10 12 9 9 13 3 2
17 1 10 12 9 13 3 3 12 1 10 9 2 2 3 13 15 2
28 10 9 15 15 1 8 13 2 4 13 2 7 4 3 4 1 10 9 1 0 7 0 9 1 0 0 9 2
23 15 0 13 9 4 10 9 2 15 1 13 9 10 9 1 15 0 2 7 0 9 13 2
38 0 4 3 10 9 1 8 7 8 7 10 10 9 7 9 15 1 8 9 8 13 1 10 0 9 3 11 13 2 10 9 15 0 7 0 9 4 2
18 1 9 4 10 9 8 10 9 1 10 9 15 11 1 11 4 4 2
38 2 1 11 0 4 10 9 1 15 9 7 15 1 11 4 7 3 4 3 1 15 9 1 11 0 4 1 0 9 2 15 9 0 13 1 15 9 2
18 10 2 0 9 2 13 1 11 4 4 2 3 0 15 9 13 4 2
22 10 1 2 9 2 0 0 4 11 13 2 1 10 0 9 1 10 9 2 1 8 2
17 3 1 10 9 13 4 4 4 16 10 9 1 10 9 0 4 2
9 1 9 4 11 1 10 9 4 2
45 1 10 9 1 10 9 1 11 13 11 1 9 12 1 10 9 1 10 9 9 9 16 0 1 4 1 11 15 1 12 9 4 4 7 3 3 3 12 9 9 13 1 10 9 2
18 11 13 1 11 1 9 12 1 12 1 11 16 15 13 8 13 13 2
15 1 15 9 13 11 3 1 12 9 1 12 9 10 9 2
18 10 9 11 1 11 13 1 8 10 9 1 15 8 8 10 0 9 2
11 15 9 13 1 10 11 1 11 4 4 2
23 10 9 13 15 9 4 1 10 3 0 0 9 2 16 3 15 0 0 15 9 13 4 2
17 9 1 11 13 3 12 1 12 9 2 15 0 16 8 1 11 2
8 10 9 1 10 9 1 9 2
17 8 2 8 2 8 2 8 2 9 11 2 9 10 2 11 2 2
17 3 13 3 2 0 2 9 2 15 1 15 0 9 0 9 13 2
19 15 13 3 3 8 3 2 1 10 13 9 2 16 15 9 8 0 4 2
20 15 4 10 3 13 9 2 15 15 1 10 9 2 0 13 2 9 0 13 2
26 10 9 13 1 15 8 1 15 9 2 7 15 13 3 3 3 2 16 10 7 15 9 0 0 4 2
7 7 11 4 3 3 11 2
12 15 13 3 12 2 3 3 12 9 1 9 2
30 10 0 9 1 8 1 10 9 2 15 3 3 11 1 11 4 2 10 9 1 9 2 15 1 10 0 2 0 9 2
6 15 9 13 15 3 2
14 10 0 9 1 9 2 8 2 13 15 3 3 4 2
7 2 13 15 15 3 2 2
5 9 1 13 0 2
10 2 0 9 2 15 4 15 3 2 2
19 15 9 13 15 9 3 1 15 7 15 9 1 10 9 1 10 0 9 2
34 3 4 10 0 9 1 11 2 7 11 5 3 1 9 11 0 13 5 13 10 13 9 11 7 13 1 10 0 9 3 8 15 9 2
20 2 15 13 3 12 9 0 4 2 7 3 12 9 13 2 2 13 9 11 2
13 2 0 9 13 11 3 0 7 13 3 3 3 2
7 15 13 15 3 4 2 2
6 15 4 0 13 0 2
24 1 10 0 9 1 10 9 1 10 0 9 13 10 9 1 3 10 9 9 12 0 9 4 2
32 2 15 13 15 3 3 2 2 13 15 2 2 16 3 3 15 9 4 4 1 10 9 7 10 9 1 9 1 11 7 11 2
26 10 9 3 13 10 0 9 1 11 10 0 9 7 13 11 7 11 4 10 9 1 11 0 10 0 2
40 16 1 10 9 13 10 9 15 2 8 2 3 1 10 9 2 15 1 10 1 12 13 0 9 1 10 0 9 2 1 10 2 0 2 9 1 10 9 13 2
8 10 0 0 1 11 4 8 2
28 10 9 4 3 4 1 10 0 9 3 10 9 3 3 1 15 0 4 2 11 13 1 10 0 9 3 3 2
22 15 13 3 0 1 10 12 9 1 12 9 7 3 13 10 9 7 9 13 9 3 2
14 3 10 9 1 10 0 9 4 0 1 10 0 9 2
11 11 13 0 7 13 12 9 1 12 9 2
13 1 10 9 11 4 11 10 9 11 1 11 4 2
51 10 9 13 15 1 10 9 3 2 13 0 13 9 3 1 12 2 3 10 9 1 8 2 12 7 8 2 12 4 4 7 13 3 1 11 2 12 2 11 2 12 7 8 12 8 2 0 12 1 12 2
18 1 11 13 11 12 1 12 2 8 2 2 8 2 13 12 1 12 2
12 10 9 13 1 10 9 3 10 9 9 4 2
31 10 0 9 13 9 0 4 1 0 9 2 3 10 0 9 4 4 1 0 9 1 10 9 9 7 9 7 13 0 9 2
27 8 10 9 1 9 13 10 9 1 9 16 0 9 4 4 4 7 3 8 9 1 10 0 9 7 9 2
20 1 10 9 1 10 11 13 0 9 0 1 4 1 0 2 0 7 15 9 2
11 3 1 11 4 1 10 9 10 9 4 2
11 15 9 13 1 8 2 10 9 1 8 2
17 3 11 4 1 15 9 8 1 10 9 1 11 1 8 1 8 2
11 10 9 1 10 9 4 0 1 15 0 2
28 4 4 16 3 3 9 4 1 10 0 0 9 2 15 3 4 4 1 10 0 9 1 10 0 12 11 9 2
4 15 13 9 2
4 9 7 9 2
31 10 12 9 1 11 7 11 13 0 9 4 4 1 10 9 11 7 11 16 9 1 9 10 9 1 13 4 16 0 4 2
26 15 9 3 13 4 2 13 0 4 1 15 13 1 9 15 3 16 1 9 1 10 9 4 13 4 2
14 15 1 9 13 2 13 10 9 4 15 10 9 13 2
12 15 4 10 0 9 2 3 15 0 9 13 2
23 15 4 10 9 15 10 9 16 10 11 13 4 1 3 10 0 9 2 15 15 9 13 2
17 3 10 2 9 2 2 15 9 10 0 9 13 1 9 1 9 2
28 3 0 4 3 15 0 1 8 13 8 1 11 2 16 4 15 3 3 1 10 0 7 1 15 0 9 4 2
23 10 9 4 4 1 9 1 15 0 8 2 0 0 2 0 13 7 0 2 7 0 13 2
25 15 13 15 1 11 8 1 8 7 0 12 0 9 1 8 2 3 3 10 9 3 1 9 11 2
34 10 0 9 1 8 13 9 4 4 1 12 9 1 10 9 2 15 8 13 4 1 10 9 1 10 0 9 1 10 0 9 1 11 2
23 10 9 1 10 9 1 8 13 16 15 9 4 4 16 11 3 10 9 13 1 12 9 2
32 10 0 9 8 13 10 9 1 8 3 4 16 15 3 8 4 2 16 3 3 13 4 4 1 10 9 1 10 9 1 11 2
28 15 9 4 4 16 11 10 9 1 10 9 1 8 2 12 2 7 8 2 12 2 16 10 9 3 13 4 2
18 3 13 3 3 10 9 1 10 0 9 7 3 13 9 11 3 4 2
20 1 9 13 10 15 11 1 10 9 2 3 0 2 7 11 4 4 1 11 2
38 15 9 13 0 3 16 10 9 1 10 9 15 10 9 3 1 4 2 7 10 9 13 1 15 3 0 9 15 11 9 13 1 10 0 9 1 4 2
38 10 9 8 2 9 2 13 9 11 1 9 0 4 16 15 9 4 4 1 10 9 16 10 0 9 1 9 0 1 9 1 9 15 9 4 4 4 2
29 4 4 16 10 9 10 9 4 16 15 9 3 0 9 4 16 2 3 3 1 9 2 10 9 1 9 1 13 2
28 10 9 13 4 16 10 9 0 4 1 4 16 10 0 9 10 9 4 1 10 9 1 10 9 1 10 9 2
21 0 10 9 3 13 1 10 9 1 10 9 12 9 1 3 2 3 1 10 9 2
38 10 8 10 9 1 11 13 9 13 3 2 16 15 3 13 4 16 16 10 9 1 10 9 7 1 10 15 9 1 10 9 1 10 0 9 1 13 2
23 1 10 9 4 15 3 4 2 0 9 1 15 12 9 2 2 7 1 10 15 9 3 2
16 1 15 8 4 4 2 16 10 9 11 15 9 0 4 4 2
40 10 9 13 3 10 9 16 15 9 15 0 0 7 0 9 1 11 4 4 2 15 0 7 0 9 1 15 9 4 4 2 7 15 9 7 9 3 4 4 2
24 10 9 16 11 7 11 15 1 9 4 13 1 15 3 4 16 10 9 10 0 9 4 4 2
6 10 0 9 4 0 2
16 1 10 1 9 8 0 13 9 4 11 3 9 1 10 9 2
43 1 10 0 9 4 8 3 10 0 2 7 3 10 9 1 11 4 4 1 10 15 15 13 13 9 7 3 3 4 4 1 9 2 13 8 10 0 9 15 9 1 4 2
22 1 9 1 9 13 11 10 9 4 16 1 4 7 15 4 0 1 9 16 0 9 2
19 3 3 4 3 1 10 13 9 10 0 9 1 4 1 15 13 1 9 2
29 10 9 2 15 10 9 1 15 8 2 13 1 10 9 1 10 9 2 1 10 15 9 13 2 13 10 9 8 2
7 2 15 4 10 0 9 2
5 0 9 13 15 2
14 10 9 4 3 3 10 0 9 1 15 9 1 4 2
9 3 0 13 10 9 0 9 4 2
22 10 9 1 10 0 9 1 10 9 2 10 9 0 9 1 3 12 9 9 2 13 2
17 1 12 8 12 4 1 15 8 1 11 10 9 4 1 10 9 2
3 11 11 2
12 15 9 13 12 9 1 8 1 15 15 9 2
23 15 4 10 9 15 8 10 9 4 4 7 15 10 9 13 1 10 9 1 11 0 9 2
8 10 9 4 8 3 3 4 2
7 1 10 9 1 10 9 2
10 2 1 11 4 10 9 3 3 0 2
9 3 0 15 4 2 3 15 13 2
9 15 9 13 3 0 1 10 9 2
31 3 13 10 9 11 10 9 10 9 4 1 10 2 9 1 9 8 16 15 1 10 9 1 15 13 1 9 1 13 2 2
29 7 16 15 13 4 10 0 9 3 1 4 1 15 15 9 2 3 13 15 15 9 2 1 9 2 3 4 2 2
3 1 9 2
18 2 3 4 2 7 13 2 1 10 0 9 8 10 9 10 9 1 2
8 15 13 15 9 0 3 9 2
7 3 4 15 15 3 0 2
27 10 9 3 10 0 9 1 15 9 15 9 3 1 10 0 9 8 4 4 2 13 3 10 3 13 9 2
14 15 4 10 9 1 9 8 2 9 1 10 0 9 2
12 1 15 13 10 9 15 3 1 10 9 13 2
22 2 1 9 1 9 2 2 13 15 15 3 2 2 13 15 10 9 1 12 9 0 2
10 8 13 1 15 9 3 12 9 2 2
30 8 2 12 2 2 15 9 11 7 15 9 11 1 12 9 4 1 10 9 1 10 0 9 11 1 10 0 11 4 2
20 3 10 9 1 10 0 9 16 9 1 10 0 9 1 10 9 2 13 9 2
20 10 9 13 3 16 9 4 4 5 9 7 9 4 1 0 9 3 0 9 2
24 1 10 0 9 4 10 9 3 13 1 10 15 9 1 9 2 3 13 12 1 12 0 9 2
10 15 9 13 3 1 15 0 9 4 2
21 2 15 4 15 10 9 1 10 11 7 10 0 9 1 10 9 8 10 0 9 2
19 1 11 13 15 10 9 1 10 9 0 1 10 9 1 10 0 0 9 2
14 15 13 15 3 3 0 1 10 9 3 15 15 13 2
11 10 9 15 0 4 13 9 3 1 4 2
20 8 13 11 1 10 0 9 1 15 9 10 0 9 1 11 1 15 9 4 2
21 1 10 9 1 15 8 13 15 1 12 2 12 2 12 2 12 1 10 9 11 2
15 15 13 15 13 1 10 13 9 1 9 7 9 1 11 2
14 10 9 1 10 0 9 4 4 1 10 9 1 11 2
14 10 9 13 3 1 10 9 1 10 0 9 15 9 2
12 3 13 15 11 12 9 0 0 0 9 4 2
38 1 10 9 8 2 15 3 10 0 9 8 13 4 4 2 13 3 15 9 8 1 11 10 0 9 2 2 12 9 2 10 9 4 4 1 10 9 2
2 11 2
33 11 13 3 10 0 9 1 12 9 1 15 9 4 2 3 15 4 13 9 2 9 2 9 7 9 1 10 0 9 3 1 4 2
18 10 10 9 4 9 2 9 5 10 9 3 0 5 13 3 3 15 2
56 1 15 9 13 15 9 2 8 10 9 1 10 9 1 10 9 1 11 2 12 2 2 2 3 3 1 8 2 10 0 9 1 12 2 8 2 12 2 2 9 1 15 9 2 0 7 0 9 1 8 2 8 2 8 2 3
11 1 12 13 8 10 0 9 1 11 4 2
10 15 4 0 9 1 10 9 1 11 2
13 2 15 13 3 4 16 15 15 9 8 13 4 2
32 8 1 11 7 11 1 11 4 10 9 4 16 10 9 8 10 9 1 9 2 9 7 9 1 10 0 7 0 9 1 13 2
16 1 10 9 1 12 9 13 10 9 15 9 2 3 10 9 2
41 10 9 8 4 10 12 9 0 9 7 4 13 1 10 9 1 9 7 9 3 1 9 1 11 7 11 4 10 0 9 1 11 2 10 0 9 1 9 1 9 2
46 16 10 9 11 3 3 3 4 4 13 1 15 9 3 10 1 12 1 8 13 9 2 15 3 3 1 15 9 4 4 2 3 13 3 12 9 3 2 7 15 1 12 9 4 4 2
29 3 1 11 7 11 4 15 9 1 10 0 9 5 10 1 10 15 15 3 1 10 9 1 15 9 13 5 4 2
14 15 1 10 0 9 3 10 9 4 4 4 10 11 2
18 10 0 9 13 3 9 16 10 9 8 1 10 0 9 4 4 4 2
39 11 13 10 9 3 4 16 15 1 10 0 9 10 9 13 4 16 10 1 15 3 0 8 1 8 1 11 1 10 9 1 9 13 9 3 4 4 4 2
9 10 9 4 3 4 1 0 9 2
23 3 4 15 0 9 4 7 15 13 3 10 0 9 16 11 10 9 1 12 1 15 13 2
7 3 13 11 15 9 3 2
15 2 1 15 9 4 15 3 0 1 15 2 2 3 11 2
7 11 13 15 9 9 3 2
13 2 1 15 9 13 11 15 15 3 0 4 2 2
17 1 10 9 4 10 0 9 2 12 9 2 10 9 1 10 9 2
5 11 13 12 9 2
26 10 0 11 13 7 1 0 7 1 15 9 3 0 2 7 10 12 13 9 13 15 12 0 9 4 2
14 2 10 9 13 1 15 9 1 3 12 9 9 2 2
5 9 1 15 13 2
12 9 2 9 2 9 2 4 0 4 16 13 2
25 10 9 2 2 9 2 13 15 10 9 5 3 1 13 1 9 5 2 13 16 10 9 1 11 2
9 15 13 16 15 9 1 9 4 2
32 10 9 13 15 1 9 8 2 15 10 0 9 2 15 1 12 1 10 9 1 11 4 4 2 1 12 3 1 9 0 13 2
47 16 15 15 1 9 13 7 3 0 0 4 2 1 15 9 1 9 4 4 2 4 1 0 3 8 1 10 0 9 0 4 2 7 15 4 3 0 0 1 15 13 1 9 1 0 9 2
12 1 10 0 9 13 11 10 0 9 1 4 2
11 10 0 9 1 8 13 10 9 1 8 2
23 1 9 4 1 10 9 4 1 10 9 1 10 0 9 2 15 1 10 9 4 0 4 2
18 8 10 9 1 15 9 1 8 13 10 9 1 8 8 3 1 8 2
19 11 13 15 0 9 1 10 9 1 15 9 0 13 8 2 3 4 4 2
37 10 9 1 11 13 15 1 10 0 9 1 15 1 4 2 7 10 9 2 3 13 2 4 3 15 15 16 0 2 3 10 0 9 0 8 13 2
30 10 0 9 2 15 1 12 9 10 9 3 12 9 13 2 13 3 1 13 9 4 4 7 0 3 13 10 9 3 2
32 10 9 1 9 1 0 13 9 5 3 8 1 9 5 1 0 9 1 4 4 4 1 11 2 10 9 7 11 4 0 4 2
16 3 4 15 1 11 4 2 3 15 9 13 2 2 13 11 2
27 16 15 9 1 13 4 13 0 0 9 1 4 4 2 15 3 3 10 9 1 10 9 1 10 9 13 2
22 9 7 9 13 11 3 1 9 2 16 3 16 15 13 4 1 10 9 1 15 9 2
46 10 9 13 16 15 0 2 8 2 2 10 9 15 10 9 1 15 0 7 0 9 1 9 13 2 3 4 1 10 0 1 15 9 2 1 10 9 2 7 3 12 9 4 4 4 2
43 10 9 1 10 9 1 0 9 15 1 10 9 13 1 12 1 12 9 2 1 10 9 2 13 1 12 9 2 1 10 9 2 2 3 1 10 9 10 9 1 12 9 2
33 7 3 13 10 3 13 9 15 0 3 2 1 10 9 0 9 3 10 9 1 10 0 3 3 1 10 9 1 10 9 8 13 2
11 10 0 9 11 4 1 3 3 1 9 2
35 10 9 1 10 9 7 9 13 3 7 15 1 10 9 3 15 9 0 4 2 16 15 1 10 11 10 9 13 4 1 10 9 1 12 2
44 3 15 9 13 10 0 7 0 0 3 1 10 9 1 10 9 15 0 12 1 10 11 2 16 15 13 16 7 10 13 9 1 11 16 10 0 9 10 9 3 0 4 4 2
23 7 10 9 13 3 4 1 3 3 9 4 1 15 9 1 10 11 7 15 1 10 9 2
25 11 7 11 3 13 10 0 9 7 11 7 11 13 1 10 9 15 0 9 3 1 10 9 4 2
4 7 15 9 2
9 13 15 15 9 7 15 15 9 2
11 13 3 10 0 9 16 1 9 1 4 2
16 3 13 3 10 9 1 11 2 15 8 1 9 1 9 13 2
23 15 13 15 13 10 9 0 0 9 2 16 15 13 15 1 15 9 1 10 9 1 4 2
16 15 4 10 3 13 9 2 7 15 13 15 7 15 13 15 2
4 16 15 13 2
12 6 2 7 3 13 15 15 3 4 7 4 2
31 2 13 15 3 4 2 9 2 16 15 1 10 15 9 0 4 4 2 13 15 15 3 13 4 3 9 3 1 4 2 2
4 2 10 9 2
5 13 15 9 4 2
29 15 13 15 3 3 1 10 0 9 1 10 0 2 0 0 7 0 0 9 1 15 9 2 2 13 10 0 9 2
8 3 1 11 2 15 9 2 2
8 3 3 6 2 1 15 9 2
10 3 13 15 4 3 15 3 1 4 2
9 16 15 3 15 3 13 4 2 2
22 7 13 15 3 3 3 15 1 9 9 4 4 2 7 3 13 15 3 1 10 9 2
17 16 9 3 1 15 1 9 13 2 3 13 15 3 3 1 9 2
29 15 9 13 3 1 10 9 1 10 9 2 16 15 15 9 13 2 10 9 1 10 9 13 2 15 13 3 0 2
7 2 6 2 13 2 9 2
9 15 13 0 9 7 15 13 2 2
5 15 4 10 9 2
13 7 3 13 15 3 8 3 3 10 0 9 3 2
5 10 9 8 13 2
16 10 12 9 3 16 0 0 9 13 11 13 3 3 15 9 2
26 12 9 3 13 15 9 3 4 2 15 1 10 12 9 8 10 9 1 10 9 2 8 2 4 4 2
11 1 10 0 9 13 15 1 10 9 9 2
13 7 3 13 15 3 4 2 16 11 3 4 4 2
9 7 3 15 9 13 15 10 0 2
5 3 13 15 9 2
6 15 13 15 9 4 2
3 6 3 2
20 10 9 7 9 13 3 3 2 13 7 13 8 3 1 10 0 9 1 9 2
23 11 0 9 1 10 3 9 13 9 15 15 3 1 15 3 0 9 13 4 4 13 3 2
19 2 1 15 0 9 13 15 0 4 2 16 15 9 1 10 9 4 4 2
2 11 2
22 2 3 4 15 0 3 0 2 16 15 16 0 1 10 12 9 1 10 9 4 4 2
9 10 9 13 15 1 15 9 4 2
39 7 3 16 10 9 12 9 3 13 15 1 10 0 12 9 15 13 9 1 10 9 1 10 9 5 10 9 13 8 3 12 9 2 5 3 3 3 4 2
10 2 15 4 0 15 3 4 4 2 2
50 15 4 10 0 9 1 10 13 9 2 16 15 15 1 15 15 15 0 13 5 7 15 4 3 15 1 15 0 9 1 10 0 0 9 5 1 13 9 13 9 1 10 12 9 1 13 9 13 4 2
5 10 9 13 4 2
32 8 2 10 9 1 11 2 13 10 9 1 15 0 9 3 1 12 9 1 10 9 3 3 0 10 9 1 9 11 1 13 2
15 9 11 13 10 9 0 7 13 10 9 1 10 12 9 2
9 2 3 2 11 2 9 7 3 2
32 16 10 9 15 9 4 4 13 15 3 4 16 10 9 2 16 15 15 1 10 9 4 4 7 4 4 1 10 0 9 2 2
9 3 13 15 2 16 15 3 13 2
10 2 13 9 8 1 9 1 0 9 2
38 10 9 1 12 9 1 15 8 7 15 2 8 2 2 4 9 1 10 13 9 8 1 13 4 5 1 10 9 1 10 9 1 15 8 1 11 4 2
35 1 10 9 4 9 4 2 3 10 9 2 15 11 8 4 4 2 4 4 1 10 9 1 9 1 10 9 2 9 7 9 1 10 9 2
20 1 3 12 9 4 10 0 9 1 15 8 4 7 4 1 10 9 1 11 2
16 3 13 11 1 15 9 2 15 15 15 1 10 9 13 4 2
19 15 4 0 16 10 9 15 9 13 4 7 15 13 10 9 10 9 2 2
19 1 10 9 7 1 10 9 1 10 9 4 10 0 9 10 9 1 9 2
18 3 4 10 9 1 10 9 12 9 2 16 10 13 9 12 9 4 2
19 0 13 3 12 9 1 9 7 1 10 9 1 0 9 4 3 9 4 2
16 15 8 13 15 1 12 13 9 12 4 1 10 9 1 8 2
12 1 10 13 9 4 3 10 9 1 8 4 2
14 16 0 4 4 10 9 2 3 12 9 2 1 4 2
23 10 9 13 3 10 0 0 9 3 1 8 2 16 1 9 3 8 2 3 12 2 13 2
29 1 9 1 8 2 12 2 1 9 7 10 0 9 1 9 1 8 2 12 2 13 3 10 9 1 0 12 9 2
29 3 13 3 10 0 9 4 4 1 9 1 10 9 2 16 0 1 10 0 9 8 4 4 4 0 9 1 4 2
7 2 3 13 10 9 8 2
36 10 9 13 3 1 10 9 1 10 0 9 10 9 1 10 0 9 4 2 8 10 0 9 16 15 3 3 1 10 9 1 12 4 4 4 2
28 10 9 13 3 3 3 2 16 15 1 10 9 12 9 0 10 9 4 4 16 1 10 9 12 9 7 0 2
9 8 13 16 0 10 9 7 13 2
11 2 4 15 9 3 4 1 10 9 2 2
8 15 13 16 9 10 0 9 2
5 10 9 4 0 2
6 3 13 15 3 3 2
17 1 10 12 9 0 9 1 11 4 15 0 16 3 15 8 13 2
17 4 4 1 10 11 13 15 4 16 3 3 13 1 10 0 9 2
32 1 15 13 15 3 7 15 13 1 0 16 0 7 1 11 1 10 9 2 7 1 10 9 15 9 0 7 0 1 4 4 2
19 0 3 13 15 0 1 15 4 2 7 15 13 3 2 16 15 4 4 2
11 15 13 15 7 15 4 15 1 11 13 2
32 7 3 4 3 3 10 9 9 7 9 5 10 10 3 0 16 10 15 5 0 2 0 2 4 15 3 3 13 0 3 3 2
10 0 0 2 7 3 0 0 1 9 2
19 1 11 13 15 3 3 1 10 9 1 4 2 16 15 0 4 1 4 2
8 15 13 3 15 15 9 4 2
8 15 13 15 9 15 9 3 2
9 15 13 3 10 0 9 3 4 2
7 15 13 15 3 0 4 2
16 10 9 1 8 13 8 2 7 15 13 3 8 15 9 0 2
9 10 9 13 15 1 12 9 3 2
28 15 13 10 9 2 15 3 0 12 9 4 2 7 15 13 15 3 3 0 4 16 15 3 12 4 4 2 2
27 10 9 1 10 0 9 2 8 2 2 13 3 9 4 1 10 9 1 10 9 1 15 8 1 10 9 2
27 3 15 9 13 3 0 9 1 10 9 2 3 15 8 2 15 8 7 10 9 2 7 15 8 4 4 2
21 8 2 9 1 3 15 8 2 13 11 0 10 9 1 9 7 10 9 1 11 2
9 9 11 4 8 11 3 1 4 2
18 1 15 9 13 15 3 10 9 1 11 4 3 9 11 15 13 4 2
15 10 9 13 15 16 15 3 9 13 4 1 15 9 8 2
8 1 15 9 1 11 13 15 2
23 2 15 4 15 3 1 15 9 0 4 7 10 9 1 15 4 0 16 1 10 9 2 2
15 3 11 13 15 0 1 10 9 1 10 9 1 12 9 2
36 1 10 1 10 11 13 9 1 0 12 9 2 3 13 7 13 1 10 9 7 1 15 9 13 2 4 10 11 16 10 3 0 9 8 4 2
15 16 15 9 3 4 4 13 11 3 3 2 7 13 15 2
21 12 9 1 15 13 13 10 11 10 3 0 9 2 12 9 13 0 1 10 11 2
32 10 11 13 1 12 9 1 10 0 9 2 10 11 1 12 9 1 10 0 7 10 11 5 1 12 9 5 1 10 0 9 2
34 11 13 10 9 4 1 15 9 2 15 15 1 11 1 0 9 1 11 2 11 7 8 13 1 10 9 2 15 8 11 3 4 13 2
31 15 3 13 15 0 13 3 1 10 0 9 1 15 0 0 9 2 15 1 10 9 12 8 10 0 9 11 1 11 13 2
18 15 4 10 1 0 9 13 9 1 11 8 2 3 11 9 4 4 2
13 6 2 10 9 4 3 0 2 3 1 0 9 2
52 3 13 9 7 9 2 3 13 10 9 1 0 9 7 9 1 9 7 9 2 3 13 0 9 16 0 1 9 2 3 13 10 0 7 0 2 3 13 0 9 1 9 7 3 13 10 9 1 9 7 9 2
17 3 13 10 0 9 2 10 0 9 2 10 0 9 1 9 12 2
39 2 15 4 10 0 9 2 15 3 3 3 13 16 15 1 15 9 15 3 1 15 0 4 2 7 3 10 9 1 9 13 15 0 9 1 15 13 4 2
16 3 16 15 15 3 8 1 15 0 4 1 15 15 9 2 2
8 2 9 13 15 0 10 9 2
30 11 4 3 8 10 9 1 11 1 10 0 11 2 10 9 15 3 1 12 13 7 3 15 9 1 9 1 4 4 2
10 10 9 13 1 15 3 0 11 9 2
9 2 6 2 11 4 10 0 9 2
13 0 4 15 3 16 15 3 13 3 15 1 4 2
17 10 9 1 3 11 7 8 4 0 7 13 10 9 1 10 9 2
15 16 11 3 1 0 13 9 13 4 4 3 9 4 2 2
14 8 2 12 2 2 9 1 15 8 1 11 2 13 2
3 15 13 2
8 2 3 15 13 15 3 4 2
9 8 13 15 9 3 3 4 4 2
15 10 9 1 11 13 9 1 2 9 2 1 10 9 4 2
24 15 13 10 9 1 10 0 12 9 9 15 3 0 2 3 15 3 3 10 0 9 13 4 2
16 2 7 3 13 15 1 12 9 3 3 1 2 2 13 8 2
17 2 13 3 16 11 8 10 9 4 4 7 3 1 9 4 4 2
10 15 13 13 15 3 0 4 4 2 2
31 10 9 1 8 13 3 0 9 4 2 1 10 9 2 16 10 9 1 15 8 1 15 0 8 3 1 10 0 4 4 2
31 10 9 1 10 8 0 4 1 9 1 10 16 12 9 13 2 16 1 10 0 9 1 11 3 3 15 9 7 12 13 2
32 10 9 4 3 15 0 16 10 0 9 2 15 13 1 10 9 1 1 12 12 9 2 7 3 12 12 15 16 10 0 9 2
32 1 10 0 9 1 9 7 9 13 3 15 0 8 1 11 2 11 2 15 3 12 9 0 9 11 1 10 9 1 11 4 2
28 1 10 0 9 1 15 15 9 13 15 3 1 10 0 9 15 9 4 4 2 16 15 15 7 10 9 13 2
21 0 1 10 9 13 10 9 2 15 3 1 9 3 1 10 9 3 4 2 3 2
15 10 9 2 0 2 4 1 15 15 9 3 3 0 0 2
13 10 10 9 1 3 1 4 9 1 9 7 9 2
24 0 9 2 15 3 1 0 9 3 13 2 13 15 0 4 1 10 0 13 1 15 9 2 2
15 3 0 4 10 9 1 10 9 15 9 1 10 9 13 2
9 2 12 1 12 9 1 10 9 2
5 15 13 3 3 2
14 1 10 9 4 10 0 9 1 12 9 1 9 0 2
16 10 9 1 10 9 15 0 4 13 1 10 12 7 12 9 2
20 10 9 1 10 9 8 16 15 13 1 4 2 13 10 9 11 2 0 2 2
17 10 9 13 3 3 10 0 9 4 4 7 3 13 10 9 3 2
24 15 13 1 10 0 9 10 0 9 1 10 9 15 8 10 9 1 10 9 10 9 4 4 2
35 15 13 3 4 10 9 1 9 16 11 2 11 2 2 8 2 11 2 7 11 2 11 2 5 15 2 3 16 11 2 9 1 10 9 2
12 1 10 0 9 13 1 10 9 3 9 9 2
26 9 8 1 10 9 1 10 9 11 1 15 8 1 11 13 3 1 8 0 1 10 9 1 10 9 2
21 10 9 2 8 12 9 2 13 0 3 8 1 10 9 7 13 13 1 10 9 2
20 10 9 11 13 0 3 15 9 2 15 1 10 9 1 10 9 10 9 13 2
20 15 8 4 10 0 9 1 11 7 1 10 9 1 10 9 13 3 10 9 2
11 3 10 0 9 13 7 13 15 3 4 2
18 15 13 1 10 9 0 10 9 1 10 9 1 10 11 7 0 9 2
13 3 4 10 9 1 10 0 9 1 10 11 4 2
25 3 13 9 1 10 9 1 10 11 1 10 9 2 10 0 9 4 3 0 1 10 0 9 2 2
6 3 13 15 3 0 2
6 15 13 10 15 9 2
22 9 2 9 7 9 13 15 9 4 4 2 15 10 9 1 10 9 7 10 9 13 2
5 11 4 3 4 2
26 15 0 8 2 8 2 15 3 15 9 1 0 9 13 2 13 15 16 10 0 9 4 4 16 9 2
13 16 15 3 15 9 1 10 9 13 16 10 0 2
31 2 15 13 3 10 9 1 10 9 2 2 13 10 0 9 1 10 0 2 16 15 11 2 1 10 9 9 2 4 4 2
8 13 7 13 13 15 10 9 2
31 13 10 9 1 11 10 9 4 7 3 4 10 0 9 2 0 7 9 2 1 11 0 9 7 9 8 7 11 9 8 2
19 1 15 9 13 3 10 0 9 4 4 2 16 10 9 1 11 4 4 2
27 10 0 9 3 13 3 10 11 4 2 15 1 15 3 13 8 15 9 3 1 10 9 1 11 13 4 2
9 10 9 13 3 3 16 0 9 2
12 15 4 3 3 9 7 8 9 1 0 9 2
20 1 15 9 13 15 10 9 4 4 2 16 8 3 1 15 9 9 13 4 2
21 10 0 9 4 9 2 7 13 15 0 4 4 2 16 15 3 1 9 4 4 2
14 3 0 13 1 11 10 9 2 3 10 9 15 4 2
6 3 0 4 10 9 2
13 10 11 13 3 1 10 0 9 2 15 8 13 2
23 10 9 1 9 4 0 16 11 1 4 2 16 15 9 1 10 9 1 13 7 1 13 2
23 15 13 15 1 15 9 4 7 1 10 0 15 15 3 3 13 2 13 15 15 0 9 2
15 15 13 15 16 10 0 0 9 1 10 9 0 1 13 2
24 7 16 15 3 13 16 10 9 3 0 3 4 1 10 9 1 4 2 4 15 0 1 15 2
12 15 4 0 0 16 15 15 9 4 4 2 2
7 3 13 15 15 13 8 2
46 1 10 9 13 3 12 9 3 2 10 9 11 2 10 0 9 2 13 1 10 0 0 9 2 15 1 15 15 9 0 9 13 1 10 2 9 2 2 3 9 1 15 9 4 4 2
11 2 8 2 2 8 1 10 9 1 8 2
10 1 3 8 2 8 2 8 7 8 2
2 0 2
7 1 11 2 8 7 11 2
20 8 4 0 7 15 9 13 3 1 10 9 16 10 9 1 0 2 0 9 2
20 15 13 3 10 0 9 1 10 0 9 1 11 11 2 15 3 0 4 4 2
19 2 10 0 9 1 10 0 9 3 15 15 0 9 3 0 4 4 2 2
48 3 4 1 15 9 15 9 1 9 1 4 1 10 9 2 15 3 1 0 9 13 4 16 3 9 4 4 1 9 2 3 15 8 7 10 9 2 10 9 15 1 10 0 9 3 0 4 2
23 0 4 15 9 3 3 10 9 1 0 9 2 3 10 9 1 9 1 15 9 4 4 2
11 3 4 3 1 15 9 15 9 1 9 2
30 1 10 9 2 0 16 15 1 15 9 13 4 2 13 10 0 0 9 2 11 2 3 2 15 1 10 15 11 13 2
32 8 13 3 1 10 0 9 1 10 9 3 0 4 1 10 9 1 10 9 2 10 9 15 15 15 9 13 4 3 1 4 2
16 3 13 9 8 10 9 7 9 7 8 10 9 8 4 4 2
30 15 9 4 15 3 3 0 2 16 9 1 15 15 13 4 16 15 0 9 1 10 9 1 0 13 9 3 1 4 2
5 11 13 10 9 2
20 10 9 13 16 16 10 9 9 1 10 9 13 2 15 10 0 9 4 4 2
25 15 4 4 1 10 9 1 10 9 1 9 2 7 10 9 4 13 1 10 15 9 9 1 4 2
29 15 13 0 15 15 9 1 10 9 2 7 15 4 3 1 10 9 10 9 10 9 0 1 13 2 3 10 9 2
31 1 10 9 15 3 10 9 1 9 4 13 1 10 15 9 1 10 9 7 10 9 1 10 9 2 4 15 10 9 4 2
15 3 13 15 1 10 15 9 1 10 0 9 1 10 9 2
29 16 15 3 4 13 7 16 3 10 9 13 4 4 4 0 13 2 16 13 15 10 0 3 0 15 3 1 13 2
21 11 13 15 11 3 1 4 2 7 10 9 4 3 3 1 15 9 3 1 4 2
23 1 10 0 9 4 10 9 1 12 9 3 0 1 4 2 16 3 15 0 9 4 4 2
12 10 0 9 1 11 13 3 3 10 13 9 2
43 3 10 9 1 15 8 4 1 15 3 3 0 0 2 16 4 10 15 0 15 3 3 3 0 16 15 11 4 10 11 1 9 1 4 5 3 0 10 0 9 8 4 2
12 8 1 10 0 9 11 2 3 11 4 0 2
25 3 13 3 12 9 10 9 7 13 1 10 9 1 10 9 9 3 16 1 9 7 9 1 13 2
14 15 0 12 9 13 3 8 4 16 10 9 1 13 2
10 12 9 4 4 7 10 9 4 4 2
10 12 15 9 13 3 12 9 9 3 2
15 1 8 1 11 4 3 12 9 1 10 0 9 8 4 2
34 16 9 4 4 10 9 1 10 9 2 16 3 10 9 3 9 11 10 9 1 10 9 1 9 13 4 4 2 9 1 9 13 4 2
22 1 10 11 13 9 8 2 15 2 1 15 9 1 9 1 10 9 2 10 9 13 2
26 10 9 13 8 10 9 0 4 4 2 7 10 9 13 3 8 3 8 10 9 0 1 9 1 4 2
24 10 0 9 13 3 1 10 13 9 15 9 1 10 1 9 8 13 0 9 1 0 9 4 2
23 12 9 13 3 7 12 3 2 1 15 10 9 1 10 0 9 7 1 10 0 0 9 2
23 10 9 1 10 0 9 8 2 11 7 11 13 15 9 3 1 11 9 1 10 13 9 2
12 15 4 3 10 9 7 10 9 0 13 4 2
31 1 8 2 9 1 11 15 16 9 10 9 13 2 13 10 9 1 10 0 9 3 1 12 9 1 10 9 1 10 9 2
32 2 16 15 2 10 9 11 2 10 0 9 1 11 2 9 13 4 4 16 15 0 9 1 13 4 2 13 15 15 3 4 2
10 15 4 0 16 15 9 15 12 13 2
18 7 15 4 3 3 0 0 16 10 9 7 15 8 2 2 13 15 2
25 3 13 10 9 1 11 7 11 5 3 0 7 3 0 16 0 1 4 5 1 10 9 1 11 2
32 1 15 9 13 15 10 9 3 15 15 16 9 15 13 4 16 16 9 7 15 13 4 16 11 1 15 9 10 0 9 13 2
16 10 9 7 0 9 4 1 10 9 10 0 9 1 10 9 2
34 1 15 9 1 10 9 1 9 13 15 8 10 0 9 2 15 8 4 16 1 15 9 7 8 10 0 2 9 2 13 9 1 4 2
30 1 10 9 1 10 9 13 10 9 1 10 0 3 0 4 4 16 15 1 10 9 1 10 9 1 9 10 9 4 2
19 3 1 10 0 9 1 10 9 13 15 9 1 10 9 1 9 4 4 2
29 1 10 9 1 10 9 13 10 9 3 1 10 9 1 0 9 1 10 9 4 2 16 9 4 4 1 10 9 2
10 15 13 16 15 9 3 0 0 13 2
37 0 4 1 15 9 10 3 1 11 13 9 1 10 0 0 9 8 3 13 16 3 15 15 9 4 4 2 15 4 4 1 10 0 9 1 11 2
17 10 9 13 0 4 4 1 10 0 9 1 10 9 1 10 9 2
33 10 9 13 1 15 10 9 1 10 0 9 1 10 9 7 10 9 1 15 8 4 2 16 10 9 0 15 13 0 9 13 4 2
28 7 3 4 15 0 15 9 2 15 1 10 9 8 2 1 12 7 12 9 1 15 9 7 15 9 4 4 2
21 15 9 13 3 3 0 1 10 9 2 8 2 1 11 1 9 2 9 7 9 2
34 15 13 3 15 9 3 7 15 4 2 0 3 2 15 13 3 3 15 0 4 4 2 10 0 2 0 10 0 3 15 9 3 13 2
7 3 4 0 15 4 3 2
5 8 13 0 9 2
22 8 7 8 13 3 1 8 2 3 3 10 9 2 10 3 13 9 15 15 9 13 2
13 10 11 13 1 10 0 9 15 15 9 9 4 2
30 1 3 1 4 1 10 9 11 2 15 1 0 9 1 10 11 7 11 4 4 2 3 4 1 8 2 9 2 9 2
18 9 1 10 11 7 11 13 3 4 16 1 13 4 1 10 0 9 2
34 10 0 9 7 0 3 10 13 13 9 1 11 7 11 13 13 9 3 1 10 9 4 1 4 16 1 12 1 11 10 9 4 4 2
38 9 11 13 15 9 1 10 9 1 10 0 9 11 4 2 16 15 7 9 11 1 11 4 4 16 3 10 9 1 10 0 7 10 0 9 1 4 2
16 3 4 3 4 1 10 9 1 15 9 2 7 1 0 9 2
24 1 10 0 9 1 10 9 4 15 0 2 3 16 10 9 1 15 9 10 0 9 3 13 2
33 3 4 11 0 2 11 2 1 12 3 15 0 2 10 0 9 1 10 9 7 10 9 1 10 13 9 7 10 13 9 16 9 2
4 12 0 9 2
22 1 9 11 13 9 1 9 1 9 15 15 9 13 2 1 4 4 1 10 0 9 2
35 10 9 1 9 1 10 0 9 2 7 1 9 7 1 0 9 2 13 10 0 9 2 3 13 8 1 10 9 1 10 3 13 9 8 2
27 10 9 15 1 15 8 1 15 13 9 16 11 7 11 3 9 4 2 7 1 11 3 10 9 4 4 2
24 10 0 9 2 7 3 10 9 1 15 9 7 1 10 0 9 13 10 9 1 0 9 8 2
17 1 10 0 9 8 4 10 13 11 0 10 0 7 15 0 9 2
20 15 13 15 9 2 9 7 9 4 4 2 15 0 9 13 0 7 0 9 2
46 15 13 10 9 8 5 10 0 9 1 12 0 13 9 5 7 3 10 9 1 10 3 13 9 1 15 9 1 12 2 8 2 10 9 4 15 9 2 7 13 3 15 0 1 4 2
28 15 13 10 0 9 4 16 8 15 0 9 1 10 9 12 2 15 15 0 9 1 11 13 2 3 13 4 2
47 0 16 11 2 11 2 8 7 11 13 3 3 1 10 9 3 1 4 2 4 10 9 1 11 2 15 15 10 0 9 1 15 0 1 15 9 3 3 1 10 9 13 4 2 3 0 2
20 1 10 9 1 10 0 11 4 1 15 13 1 10 2 9 2 10 9 4 2
3 12 9 2
28 15 13 2 16 3 0 0 1 10 9 1 10 9 4 4 4 16 1 10 0 9 7 10 0 9 1 13 2
42 10 9 11 2 15 13 1 10 0 9 1 10 9 7 10 9 1 10 9 1 10 0 9 2 13 1 2 8 3 0 9 2 15 4 13 4 1 10 9 7 9 2
21 10 9 1 10 0 9 4 1 10 9 11 8 4 1 15 13 1 10 0 9 2
12 3 1 9 7 3 1 15 9 1 12 4 2
4 5 15 8 2
14 5 15 8 2 10 0 9 15 0 16 3 0 13 2
9 5 10 11 2 10 0 0 9 2
10 5 10 0 9 2 1 15 10 9 2
39 13 1 10 9 1 10 9 4 15 10 0 9 3 4 2 3 13 1 4 4 16 9 1 10 9 3 1 9 4 1 4 4 2 7 1 2 9 2 2
3 0 9 2
64 10 9 1 8 1 11 13 15 15 2 13 2 4 4 2 7 1 0 12 9 9 13 10 9 13 10 9 1 9 11 4 16 11 5 15 9 13 5 3 3 8 4 13 7 3 10 9 4 4 16 16 2 0 2 1 9 3 1 10 9 1 13 4 2
2 9 2
5 10 9 4 13 2
21 10 9 11 13 15 3 13 9 1 10 9 1 10 11 4 1 10 9 1 11 2
17 15 13 3 8 10 9 11 10 9 1 10 0 9 1 10 11 2
11 1 10 9 13 3 10 9 1 10 9 2
20 11 13 9 1 10 9 15 13 4 1 9 1 10 9 1 10 13 0 9 2
7 4 4 1 9 7 9 2
16 2 9 2 2 5 1 15 0 0 2 5 2 6 9 2 2
23 15 4 3 0 0 2 7 3 15 1 11 13 15 10 9 4 2 8 3 15 3 4 2
17 1 0 9 4 10 9 0 4 16 15 1 8 1 9 13 4 2
30 10 0 9 1 15 9 13 1 10 9 1 8 1 11 2 7 10 9 1 10 0 11 4 3 0 16 11 15 9 2
10 15 9 13 3 1 10 9 12 9 2
26 15 13 15 4 16 16 15 10 9 13 2 7 10 9 3 15 13 13 3 4 16 16 15 0 4 2
26 15 8 13 10 1 12 13 12 9 13 9 8 1 9 4 1 10 9 1 10 9 11 2 11 2 2
21 10 9 2 1 9 1 12 9 2 4 1 12 1 10 0 9 4 1 10 11 2
28 10 9 1 10 11 2 15 10 9 1 10 9 11 1 10 9 13 2 13 16 15 8 0 0 1 4 4 2
14 1 10 9 1 15 9 13 10 9 15 9 1 4 2
6 10 9 4 9 13 2
12 3 4 10 0 12 0 9 8 4 1 12 2
9 16 15 13 4 10 9 12 9 2
10 3 4 15 8 8 1 15 9 4 2
20 9 8 13 3 0 3 2 7 3 0 13 13 3 10 9 1 3 0 9 2
8 10 9 4 4 1 12 9 2
9 3 4 9 1 15 9 1 4 2
10 1 10 0 9 4 11 12 9 0 2
7 3 11 13 15 9 4 2
20 3 13 3 3 15 9 16 15 15 9 1 9 7 9 1 11 0 4 4 2
14 13 1 15 9 1 4 13 10 9 2 10 9 13 2
15 2 15 13 4 16 15 16 15 13 10 0 9 4 2 2
17 1 15 9 13 10 0 9 10 9 4 1 10 0 9 8 11 2
10 3 4 15 3 1 10 0 9 4 2
20 9 8 1 10 0 11 13 15 3 1 10 0 9 3 4 4 1 15 9 2
16 1 10 9 13 5 7 15 4 15 13 5 10 9 0 8 2
34 3 13 15 3 4 1 15 9 1 0 9 2 15 3 10 9 13 4 16 9 1 13 1 10 9 15 15 1 10 9 13 4 4 2
27 10 9 1 9 1 8 8 13 10 0 9 3 2 3 10 9 3 0 13 1 10 9 8 13 4 4 2
22 10 11 13 0 4 9 0 1 4 1 10 0 9 1 10 11 7 1 15 0 9 2
23 15 9 13 10 9 1 15 9 4 4 2 3 10 0 9 1 0 7 11 13 4 4 2
19 15 9 13 3 10 0 9 1 0 9 2 11 2 1 10 9 1 11 2
12 1 11 13 11 3 3 4 4 16 10 9 2
15 11 13 3 3 16 1 10 0 9 10 0 9 1 4 2
25 3 16 1 13 16 15 1 10 13 9 1 10 9 4 1 4 13 10 0 9 10 9 11 4 2
20 3 4 15 3 1 10 9 4 16 10 9 1 11 13 3 3 10 9 3 2
17 15 13 16 10 0 9 16 9 1 10 0 9 0 9 4 4 2
25 10 9 1 8 2 12 2 4 8 3 0 16 10 0 9 1 11 2 0 7 11 3 1 13 2
27 1 15 9 1 15 9 15 11 4 13 4 3 3 4 2 16 1 10 9 1 10 9 15 3 8 13 2
22 15 3 3 13 1 4 2 16 10 9 1 10 9 3 3 3 3 10 9 4 4 2
16 3 13 3 15 10 0 7 0 9 1 11 13 3 15 8 2
24 10 9 8 2 0 16 9 7 16 9 1 10 9 1 10 9 1 8 2 4 1 8 4 2
5 15 4 12 9 2
12 8 2 0 11 2 4 0 1 11 1 11 2
45 15 13 2 1 0 9 1 13 4 1 10 0 9 8 2 1 12 1 11 9 2 3 15 2 1 10 9 1 3 12 9 1 2 15 13 3 10 15 9 2 2 3 4 4 2
29 1 10 0 0 9 1 10 11 5 10 9 4 12 1 12 5 13 11 10 9 1 0 9 4 4 1 10 9 2
24 3 15 4 10 9 1 15 3 3 1 3 4 4 1 10 9 10 9 15 3 13 4 4 2
17 3 13 15 9 10 9 10 9 4 4 2 3 10 9 1 4 2
15 7 15 12 13 9 7 9 15 9 8 15 9 0 4 2
21 10 9 1 15 9 13 3 10 9 3 4 16 3 15 13 1 10 9 3 13 2
30 12 9 1 10 0 9 10 0 9 2 13 2 1 11 2 8 7 8 2 4 13 2 3 13 10 9 1 11 4 2
22 10 9 4 1 10 0 9 8 4 1 15 9 2 16 1 10 11 1 3 4 4 2
12 15 9 13 9 1 9 3 10 9 4 4 2
35 1 10 9 1 10 9 13 16 10 9 3 9 13 1 10 9 1 10 9 2 7 15 13 10 15 9 4 4 2 15 15 1 10 9 2
17 10 0 9 13 3 4 16 9 7 9 12 9 1 15 9 4 2
20 16 3 1 10 9 9 0 4 2 13 15 3 3 10 9 1 9 4 4 2
26 15 9 4 8 10 9 1 12 0 3 2 4 2 1 16 0 9 2 16 3 3 15 4 1 4 2
7 1 12 13 15 3 3 2
21 3 13 8 12 9 2 15 15 3 13 4 4 2 16 4 15 0 9 3 0 2
36 1 10 9 1 11 13 15 8 8 2 8 2 10 9 4 1 10 9 8 2 15 15 3 13 15 1 10 11 0 1 10 9 1 4 4 2
32 16 15 5 1 12 5 1 0 9 1 10 11 13 4 11 3 1 15 8 7 1 15 8 2 9 1 15 8 2 13 4 2
16 1 15 9 13 15 15 1 10 9 1 10 9 13 4 4 2
36 0 13 15 15 2 16 15 3 10 9 13 2 1 10 9 1 10 9 2 7 15 13 3 3 9 2 9 7 9 2 9 7 2 9 2 2
17 15 13 3 2 3 2 10 9 4 7 3 0 10 9 3 4 2
52 10 0 9 2 15 3 4 4 1 10 9 3 3 10 0 7 3 1 10 9 1 10 9 3 15 0 0 9 1 4 1 10 9 1 15 9 2 13 8 1 10 0 9 4 1 10 9 1 12 0 9 2
8 11 1 8 7 8 1 11 2
23 16 9 1 15 9 13 4 10 9 8 2 10 9 8 2 10 9 8 7 10 9 8 2
40 10 9 4 15 1 10 9 3 3 2 16 10 0 9 10 0 9 4 1 10 0 9 7 9 2 16 1 15 15 9 1 10 9 13 2 15 3 4 4 2
13 1 10 0 13 9 4 3 3 10 9 8 4 2
25 10 9 13 3 3 13 3 16 15 9 0 1 4 1 10 9 7 3 1 4 1 10 0 9 2
10 10 9 13 10 9 1 0 9 3 2
18 15 13 1 10 9 11 15 1 8 1 12 9 0 1 10 9 13 2
25 1 15 13 10 9 11 1 8 3 0 1 10 9 7 10 9 1 10 9 13 15 3 3 4 2
13 15 12 13 15 3 1 10 0 1 10 0 9 2
47 11 7 11 2 10 15 0 9 1 10 9 2 13 11 3 3 1 10 0 9 1 4 7 1 12 13 10 9 3 10 0 9 2 7 10 0 9 13 3 10 9 7 13 12 9 3 2
15 10 0 9 4 3 3 0 4 1 10 9 1 15 8 2
36 10 9 0 0 8 8 13 1 15 9 1 9 1 0 9 10 9 4 3 15 9 1 10 0 9 3 12 9 0 8 4 2 10 0 9 2
26 1 10 0 13 9 1 10 0 13 3 12 13 9 4 2 15 10 0 0 9 1 15 9 13 4 2
17 10 9 1 10 9 2 9 7 9 2 13 4 4 1 12 9 2
14 10 9 1 8 2 11 7 11 13 10 9 3 8 2
40 1 10 13 9 4 15 0 10 9 8 10 9 1 13 2 16 1 15 9 10 9 0 4 2 10 0 9 4 4 7 9 4 4 1 15 3 1 9 13 2
28 7 3 13 2 1 10 9 8 2 3 9 2 9 7 15 9 2 15 15 15 9 1 2 8 2 13 4 2
14 3 13 11 1 10 9 1 10 9 1 10 0 9 2
8 1 15 12 9 13 4 4 2
31 3 13 10 9 1 10 9 11 15 9 4 2 16 1 13 2 16 10 9 3 12 9 1 10 9 1 10 9 4 4 2
42 10 9 4 15 0 2 7 0 3 0 2 0 1 10 9 1 15 9 2 15 0 16 10 9 1 10 9 7 10 9 2 12 9 3 0 2 16 15 1 10 9 2
17 3 13 3 12 9 0 4 16 15 1 15 12 9 3 1 4 2
23 15 13 4 4 16 3 1 13 2 16 10 9 10 0 9 4 16 15 3 10 9 13 2
45 1 10 9 1 10 11 1 10 9 1 7 10 9 1 10 0 9 1 10 9 2 10 9 7 1 10 3 13 9 13 9 7 9 10 3 0 9 2 0 12 7 12 9 2 2
20 12 9 13 10 9 8 0 2 12 9 10 13 9 7 12 9 13 15 9 2
17 3 10 9 15 3 1 10 9 11 1 10 11 1 11 4 4 2
28 2 15 13 3 3 4 2 15 3 2 2 13 8 1 10 9 7 11 1 15 1 10 9 9 4 4 4 2
3 2 8 2
32 15 13 10 9 3 1 8 2 9 1 15 8 2 2 15 15 1 15 9 3 13 8 1 4 4 15 1 10 9 1 4 2
32 15 4 3 0 3 4 1 4 2 2 13 11 2 16 10 9 15 13 4 1 10 9 1 4 2 3 10 9 1 9 13 2
15 7 11 13 13 3 2 16 10 9 15 1 15 9 13 2
9 3 4 10 9 3 1 10 11 2
32 10 9 15 8 13 1 12 1 10 13 9 10 9 4 1 12 9 2 1 12 9 1 10 13 9 2 3 13 1 10 9 2
11 8 4 10 9 1 9 2 8 1 9 2
17 10 9 1 10 9 4 1 10 9 4 1 8 12 1 8 12 2
21 10 10 9 4 4 1 9 1 9 2 16 10 0 9 1 15 9 15 4 4 2
6 1 12 1 12 9 2
6 10 9 13 1 3 2
11 1 11 13 9 0 10 9 8 0 3 2
22 2 1 13 1 11 1 10 0 1 11 2 2 13 10 9 1 15 9 1 10 11 2
27 10 9 2 15 3 0 4 4 2 13 1 10 9 15 4 7 13 1 4 16 12 13 9 1 9 4 2
9 10 9 4 4 1 8 10 9 2
12 11 13 10 9 1 10 11 1 11 0 3 2
7 10 9 4 1 8 4 2
5 10 9 4 0 2
37 7 3 13 15 1 10 15 0 13 9 1 11 2 15 1 10 0 7 3 3 0 9 1 11 2 7 8 10 9 1 10 0 9 10 12 9 2
18 10 9 13 1 9 11 15 3 1 10 9 13 16 11 3 13 4 2
15 10 9 1 0 1 10 13 9 11 7 10 9 4 4 2
10 10 0 9 13 0 10 0 13 11 2
17 1 10 9 1 4 8 15 15 16 10 9 3 15 9 9 13 2
17 7 0 13 13 15 15 10 9 2 16 15 3 3 4 4 2 2
22 15 4 10 1 10 0 9 15 0 9 2 3 9 1 12 7 12 9 8 13 4 2
31 13 2 9 2 13 2 13 2 9 13 2 13 2 9 2 9 2 15 0 9 4 3 0 2 7 9 11 13 16 9 2
6 15 13 16 15 13 2
19 3 0 3 4 15 4 1 10 9 8 2 3 9 1 10 9 7 9 2
12 1 15 0 9 13 15 3 3 3 1 4 2
31 11 2 15 16 10 0 9 9 4 4 2 13 3 0 10 9 1 10 0 9 2 3 10 0 9 3 10 0 9 4 2
11 10 9 1 10 9 13 15 2 8 2 2
34 10 0 9 1 10 13 9 1 0 9 7 9 13 10 0 0 2 0 9 4 2 13 1 0 2 0 2 0 2 0 7 0 9 2
19 0 9 4 3 8 7 0 9 1 4 1 10 0 9 1 10 12 9 2
15 10 0 9 13 15 3 1 0 9 10 0 9 1 4 2
24 8 2 10 0 9 13 15 9 3 1 11 2 3 3 0 16 15 15 7 10 9 13 4 2
16 10 9 4 3 3 3 4 16 10 9 9 1 11 4 4 2
26 16 10 9 3 10 0 9 13 4 4 13 10 0 9 3 1 15 9 16 10 0 0 9 1 13 2
9 15 9 13 15 15 16 15 9 2
16 1 8 13 15 2 1 10 0 9 1 9 2 2 8 2 2
6 15 13 10 13 9 2
17 11 13 1 11 7 13 10 9 1 4 16 15 10 0 11 4 2
14 15 13 3 3 13 2 0 7 0 2 7 0 9 2
13 15 13 15 3 16 15 15 3 3 0 4 4 2
14 1 10 0 0 9 15 15 13 13 15 9 7 9 2
17 1 10 0 9 8 2 12 2 4 8 12 9 1 10 0 4 2
35 2 15 13 15 4 2 0 0 1 9 1 4 1 10 0 9 7 9 11 2 15 15 8 13 7 15 0 13 15 15 3 7 3 13 2
20 10 0 3 4 10 1 12 13 9 8 2 8 2 11 12 2 9 8 2 2
27 11 4 0 1 15 0 3 1 10 0 13 9 7 15 9 4 1 9 1 15 0 9 0 13 1 4 2
27 10 9 13 10 9 1 8 2 10 3 13 9 2 15 1 10 0 9 0 1 10 15 13 9 4 13 2
16 10 0 0 9 13 8 0 4 10 9 3 1 15 1 4 2
9 1 10 9 13 11 0 4 4 2
7 3 4 4 1 12 9 2
19 10 9 1 9 1 10 9 1 9 7 9 2 10 9 1 10 0 9 2
18 10 9 1 9 7 10 9 1 10 9 1 10 9 1 9 7 9 2
18 12 0 9 13 10 9 4 2 10 9 8 2 8 2 8 7 8 2
26 10 0 0 9 1 10 0 9 4 1 12 10 0 9 2 15 1 12 1 12 11 1 11 4 4 2
14 8 2 9 1 15 8 2 13 1 15 9 15 9 2
45 15 0 9 5 2 0 2 16 3 10 9 1 10 0 9 4 4 5 13 4 4 16 10 9 1 9 1 10 9 1 10 0 9 2 3 1 15 0 8 3 1 9 4 4 2
20 10 0 9 1 11 7 10 9 4 4 1 10 12 9 1 10 2 9 2 2
20 10 9 1 10 9 15 3 1 10 9 1 11 1 11 4 4 2 4 12 2
6 3 13 3 12 9 2
19 10 9 13 2 1 10 9 1 11 2 3 12 9 1 10 9 8 4 2
13 8 2 10 0 9 1 10 9 2 13 0 3 2
15 10 9 13 1 9 11 3 2 3 8 0 0 13 4 2
24 10 9 9 1 11 13 1 10 9 9 4 16 15 1 10 9 1 10 9 10 9 4 4 2
12 1 10 0 9 4 10 9 3 1 0 9 2
29 10 9 1 3 12 0 13 1 8 1 10 9 10 9 9 1 12 9 2 15 4 4 16 15 9 13 4 4 2
25 2 13 10 13 7 0 9 1 10 9 4 4 1 9 2 16 9 2 9 3 3 3 13 4 2
15 10 9 13 3 1 9 3 7 13 10 9 10 9 3 2
43 0 13 10 0 9 1 8 2 8 2 10 0 9 1 11 4 10 9 9 11 2 15 0 4 13 16 15 9 0 1 10 9 9 4 4 2 1 15 9 3 1 4 2
16 9 1 11 13 10 9 15 10 0 9 9 4 13 0 4 2
27 4 4 16 3 0 10 2 0 7 0 2 9 4 15 11 1 10 9 1 10 9 1 10 11 13 4 2
33 10 0 9 13 12 9 3 5 0 9 12 9 5 2 7 13 16 10 2 0 9 2 1 11 2 3 2 9 1 10 9 4 2
14 10 0 9 4 1 11 4 2 16 15 1 9 13 2
13 10 9 4 3 10 9 9 9 1 15 1 4 2
19 1 10 1 10 9 3 3 0 9 11 1 11 4 15 3 15 9 0 2
16 15 0 9 13 3 10 0 9 2 15 15 0 13 16 3 2
15 10 9 8 2 9 1 10 0 9 13 10 0 9 3 2
12 10 0 2 9 2 15 3 7 3 3 13 2
18 15 4 0 16 10 9 3 3 3 4 7 16 3 0 10 9 4 2
9 15 13 3 3 3 3 3 4 2
12 10 9 8 13 3 0 3 4 1 10 9 2
8 3 4 3 10 9 3 4 2
11 15 4 3 16 15 8 10 0 9 4 2
12 15 4 15 0 2 3 13 15 8 9 3 2
11 15 0 4 13 10 9 1 15 15 13 2
9 15 13 13 15 15 1 9 13 2
8 15 13 3 1 9 3 4 2
11 13 9 2 7 3 13 15 9 1 9 2
28 3 13 10 9 1 10 9 2 15 3 10 0 9 1 9 2 2 2 4 4 1 10 9 4 4 7 4 2
11 15 13 7 0 9 7 13 7 3 13 2
22 10 0 9 13 10 9 2 3 10 1 10 0 13 9 2 15 13 1 10 9 8 2
11 13 2 13 2 13 1 10 0 9 8 2
2 9 2
10 10 9 13 1 10 9 1 10 11 2
23 15 4 3 3 4 1 10 9 11 2 15 13 16 15 9 1 10 9 7 10 9 4 2
19 10 9 1 15 9 13 1 13 1 10 9 16 15 1 15 9 4 4 2
30 15 12 1 10 9 11 2 3 10 9 3 1 12 1 12 9 4 4 2 7 12 1 10 1 12 9 13 9 9 2
25 10 0 9 1 11 13 3 3 3 1 9 9 2 7 15 13 3 15 9 1 10 8 0 9 2
27 15 13 3 3 3 3 2 3 3 16 3 3 15 9 1 10 9 13 2 16 2 8 2 10 13 9 2
8 16 15 0 9 3 1 13 2
17 7 13 3 10 9 9 7 9 16 3 1 2 4 2 13 4 2
17 1 10 0 9 13 15 3 0 16 10 9 1 10 9 1 13 2
9 7 10 9 4 3 1 12 0 2
15 10 0 9 8 13 10 9 4 1 15 9 1 0 9 2
14 15 1 12 13 2 8 2 4 3 3 9 4 4 2
34 3 13 10 0 9 1 10 0 0 9 1 11 10 9 2 3 10 9 4 4 3 0 0 1 10 2 9 1 10 9 2 1 4 2
15 1 10 9 4 1 11 12 0 4 1 2 0 9 2 2
26 10 13 9 1 9 13 9 4 1 10 9 1 8 1 15 9 1 10 9 1 9 1 10 0 9 2
15 1 10 9 4 10 9 4 1 10 1 10 9 13 9 2
19 3 8 13 10 13 9 1 4 4 16 0 10 13 9 8 4 4 4 2
2 12 2
11 1 12 1 10 9 4 11 10 0 9 2
15 10 9 1 10 9 1 9 8 10 0 9 1 15 9 2
18 2 15 13 15 3 10 9 9 1 4 2 2 13 15 1 10 9 2
22 2 16 10 9 1 15 9 0 4 13 2 13 15 15 3 10 9 1 9 1 4 2
23 15 13 15 3 3 0 16 3 10 0 0 9 4 4 15 0 3 1 9 13 4 2 2
16 3 10 9 3 8 1 10 9 13 15 9 1 10 9 13 2
11 0 9 13 3 0 1 10 9 10 9 2
31 15 13 3 16 15 3 3 10 9 4 1 10 9 16 15 9 9 3 1 13 2 16 15 1 13 13 1 10 0 9 2
27 2 15 13 16 10 0 9 1 10 0 9 15 9 9 4 2 3 13 1 9 8 9 2 9 7 9 2
36 16 15 3 13 16 4 15 0 9 3 3 0 2 2 3 8 2 15 13 15 0 1 4 4 1 10 9 1 1 10 0 15 1 4 4 2
34 10 9 1 10 9 12 7 12 13 1 15 10 0 9 1 10 0 9 2 10 13 9 16 2 9 2 1 10 3 0 7 13 9 2
21 7 1 10 9 2 1 10 9 2 4 15 12 9 3 16 1 13 1 9 8 2
10 7 1 15 13 15 3 0 16 15 2
23 16 10 2 9 2 1 9 2 9 7 9 0 4 13 15 3 1 10 9 1 10 9 2
9 0 13 15 9 1 10 0 9 2
21 3 2 1 10 9 1 10 1 15 8 13 0 9 2 13 10 9 3 3 8 2
22 12 0 0 0 9 1 10 9 11 13 8 15 8 11 3 3 1 9 1 4 4 2
26 1 9 1 10 9 1 12 1 12 13 1 9 1 10 0 9 4 4 16 10 9 1 15 12 13 2
22 15 0 9 13 0 3 12 9 8 4 4 16 10 9 8 4 16 15 3 4 4 2
11 12 9 4 3 1 8 1 10 9 4 2
23 15 10 9 2 3 1 0 0 9 2 1 8 13 2 13 1 15 9 10 0 9 4 2
20 3 4 15 2 8 2 2 10 0 9 1 9 7 9 2 16 10 9 13 2
40 10 9 13 1 10 9 1 0 2 0 7 0 2 15 3 15 9 13 4 1 10 0 9 2 7 15 3 10 9 2 3 10 9 1 10 9 2 13 4 2
28 0 9 1 11 9 4 3 10 9 2 1 15 9 8 2 2 10 2 9 2 2 3 15 13 15 13 4 2
8 11 7 11 1 2 8 2 2
16 3 10 2 9 2 2 3 11 10 9 13 4 3 0 4 2
7 3 13 0 3 12 9 2
50 7 10 0 9 4 1 15 15 9 4 2 16 15 13 2 16 3 11 15 1 11 3 4 2 3 3 1 10 0 0 9 4 4 2 7 15 4 3 0 2 16 11 15 3 3 3 1 9 13 2
20 1 15 1 10 0 0 9 1 15 8 2 13 11 10 9 16 10 0 9 2
19 1 10 0 9 13 10 9 1 0 9 1 4 2 15 12 9 0 4 2
26 3 4 9 0 2 2 10 0 9 1 15 9 13 3 1 12 9 2 7 12 9 4 10 0 9 2
10 10 9 13 3 3 3 8 3 4 2
27 15 4 1 15 10 0 9 9 1 10 9 2 3 16 15 13 8 0 9 15 9 1 8 15 4 4 2
18 15 9 13 0 12 9 4 1 0 9 2 15 8 13 4 16 9 2
18 10 0 9 1 11 2 8 2 4 8 12 4 1 0 9 1 11 2
29 8 2 10 0 7 0 9 15 1 11 7 11 10 9 13 2 13 3 8 3 2 15 1 11 9 1 11 4 2
11 10 9 1 9 1 11 4 3 0 4 2
13 0 9 11 13 8 10 9 1 9 11 1 8 2
19 2 15 1 10 9 1 10 9 1 15 9 2 4 0 1 10 0 9 2
25 10 9 2 16 3 3 13 13 15 9 1 4 2 3 10 9 3 1 10 15 0 4 13 4 2
25 15 13 3 3 3 7 15 4 3 0 2 16 15 10 9 4 16 1 15 9 9 1 4 2 2
28 3 9 8 2 1 10 9 15 10 9 2 11 2 3 1 10 9 1 10 11 1 11 13 8 15 0 9 2
16 15 4 13 1 10 9 15 9 1 10 13 9 4 13 4 2
28 10 9 13 15 3 3 3 4 2 3 16 10 9 10 0 9 13 7 3 3 3 1 10 9 13 4 4 2
36 10 9 13 1 15 1 5 3 1 9 3 1 13 5 9 2 13 9 2 9 2 9 7 10 9 15 9 2 10 0 9 1 10 0 9 2
20 15 4 3 0 16 10 13 9 3 0 13 7 3 13 4 16 2 8 2 2
26 3 13 9 15 15 13 4 2 3 10 9 1 10 9 1 16 9 10 9 2 10 9 7 10 9 2
22 1 10 3 0 9 4 3 10 0 0 9 1 10 9 1 15 8 1 11 8 4 2
29 1 10 9 1 9 13 8 2 9 1 15 1 12 13 8 2 15 3 10 9 3 13 9 2 10 9 1 8 2
9 10 11 4 4 1 10 9 8 2
30 15 4 10 0 2 0 9 4 2 3 16 10 0 9 2 15 1 9 4 13 4 9 2 9 7 10 9 4 4 2
22 15 4 1 8 0 3 15 0 9 2 16 15 15 3 0 13 9 0 13 1 4 2
30 2 13 9 13 1 9 1 9 4 4 7 1 10 9 1 12 13 10 9 1 10 11 3 1 10 1 9 13 9 2
18 15 13 15 3 3 3 2 7 1 12 9 13 15 3 4 3 2 2
29 2 15 4 3 0 0 16 10 9 1 10 9 3 0 13 4 2 16 15 3 1 13 13 4 1 10 9 2 2
22 13 10 9 1 15 9 1 9 1 0 9 8 3 0 9 2 3 13 10 9 4 2
25 8 10 9 1 10 9 1 15 8 2 13 8 12 3 10 9 7 10 9 1 10 9 4 4 2
22 3 4 10 9 1 4 1 10 0 9 3 10 9 8 12 4 4 1 8 1 8 2
13 10 9 1 8 7 8 4 4 1 8 3 8 2
35 12 0 9 2 9 1 10 11 1 9 1 9 7 9 2 4 3 1 8 1 10 9 1 11 4 2 16 15 1 12 3 13 4 4 2
28 12 9 0 13 10 9 2 10 9 9 7 10 0 9 9 10 9 4 1 10 9 7 9 1 10 0 11 2
23 1 12 9 13 15 9 15 8 10 9 4 1 10 9 1 12 9 2 15 1 9 4 2
26 10 9 8 1 11 2 0 1 15 8 1 11 2 4 1 8 4 1 10 0 9 13 1 15 8 2
15 10 9 4 15 4 1 9 11 1 10 9 1 10 9 2
18 10 9 8 2 13 8 13 1 12 16 0 9 1 10 9 1 9 2
15 15 13 3 1 13 9 7 13 1 12 16 9 1 11 2
12 1 10 0 9 2 13 15 10 0 9 4 2
12 11 13 15 1 11 7 1 11 15 9 4 2
7 7 15 4 10 9 3 2
7 15 13 3 10 9 2 2
20 3 2 13 15 1 15 0 9 2 13 15 9 9 1 4 1 10 0 9 2
10 15 13 2 16 15 9 3 0 4 2
23 11 2 3 3 15 1 12 15 9 1 11 13 4 2 13 15 10 9 8 3 0 0 2
18 10 9 1 11 13 15 3 1 0 9 4 1 10 1 11 13 9 2
32 10 9 1 10 9 13 3 10 9 2 16 10 2 0 4 2 9 3 10 16 12 9 0 4 4 16 1 10 9 1 4 2
7 10 9 11 2 11 2 2
15 2 15 4 15 9 2 15 10 12 9 16 0 13 4 2
17 1 10 0 9 4 15 10 0 13 11 15 10 9 1 11 13 2
22 10 9 13 1 10 0 9 15 12 9 4 7 3 13 15 10 9 3 0 3 4 2
16 8 13 1 15 9 1 10 9 1 15 8 7 8 15 9 2
15 15 13 15 9 1 15 2 3 4 12 9 1 15 4 2
19 1 15 9 13 15 15 15 9 2 15 0 8 2 15 13 9 1 4 2
17 0 1 10 9 4 10 15 9 1 11 2 10 0 9 8 4 2
11 11 4 8 10 9 11 3 3 0 4 2
14 15 13 16 9 7 9 1 10 9 10 9 4 4 2
25 0 9 4 1 10 9 3 0 1 10 0 9 2 3 10 9 2 7 15 13 1 10 9 3 2
23 15 9 7 9 13 10 0 9 9 3 7 13 9 1 10 9 1 10 9 2 13 15 2
28 10 9 13 10 13 0 1 12 9 8 10 0 9 10 9 4 1 9 1 9 7 9 1 12 9 1 9 2
39 0 0 13 11 15 9 2 16 0 11 0 13 4 16 11 15 0 1 8 13 7 16 11 0 3 13 4 16 11 15 1 10 9 0 1 10 9 13 2
28 1 11 11 2 1 10 11 1 10 11 4 3 10 9 4 2 3 12 9 2 15 10 9 13 2 13 4 2
9 10 9 1 10 1 15 4 0 2
9 15 4 4 1 15 8 1 11 2
33 1 9 12 2 15 4 4 2 13 10 9 1 11 2 8 2 15 9 11 3 1 10 9 1 10 11 1 11 15 9 13 4 2
9 10 9 13 1 10 9 1 8 2
26 10 9 1 11 2 13 1 12 9 2 4 3 1 11 1 8 1 10 9 1 10 9 4 7 4 2
11 15 16 10 9 1 10 9 4 3 4 2
16 10 9 2 15 3 4 1 10 9 2 13 3 10 0 9 2
18 10 9 2 3 10 9 0 4 2 13 10 0 9 3 1 10 9 2
38 1 10 0 9 13 9 8 4 1 10 9 1 9 11 1 10 1 10 9 0 9 1 10 0 9 1 10 9 2 15 9 8 1 12 1 15 13 2
14 2 0 2 7 2 0 2 15 0 9 1 15 9 2
30 12 0 9 3 1 11 1 10 0 9 2 3 8 15 4 13 4 1 10 9 1 10 9 2 15 3 10 9 13 2
18 10 9 11 13 16 10 9 0 4 4 7 16 15 15 4 4 4 2
20 10 9 1 10 9 4 0 0 2 7 0 13 3 0 2 3 10 9 11 2
21 10 9 13 3 0 7 1 11 13 15 10 11 9 4 16 3 15 3 1 4 2
11 1 3 15 9 13 15 15 9 4 2 2
16 1 8 13 15 9 10 11 4 10 9 1 12 3 1 4 2
7 3 4 3 15 9 4 2
36 1 15 9 4 10 9 1 10 11 4 16 15 9 2 3 15 1 10 9 2 10 9 8 1 11 2 3 1 4 1 10 9 1 10 9 2
24 3 13 10 0 9 1 10 9 10 0 11 2 10 0 11 2 10 0 11 7 10 0 11 2
24 10 0 9 0 9 1 11 2 11 2 11 2 11 2 13 3 10 9 1 10 0 9 11 2
45 1 10 9 13 15 16 10 9 1 11 1 8 2 11 2 11 2 11 7 11 1 4 4 16 1 15 9 11 10 9 4 4 2 16 3 10 1 11 13 9 16 9 1 13 2
15 10 0 9 2 15 10 9 13 2 13 3 10 0 9 2
7 15 4 15 9 1 9 2
11 10 0 9 2 15 15 13 4 10 0 2
7 15 4 0 0 1 9 2
15 15 13 0 16 15 10 9 13 9 1 10 9 3 3 2
10 3 13 10 9 3 3 1 15 9 2
12 15 13 10 9 1 9 7 3 10 0 9 2
22 15 13 3 1 10 9 4 4 16 15 15 9 3 1 13 3 10 9 0 4 2 2
15 10 0 9 1 15 9 4 0 4 1 0 2 9 2 2
16 10 9 13 5 1 0 9 13 5 10 9 1 10 9 9 2
9 10 0 9 4 1 15 9 4 2
20 8 1 10 9 4 15 10 9 4 9 1 10 0 9 1 10 9 1 4 2
21 13 15 1 15 15 15 12 9 0 2 3 13 15 10 9 3 9 10 9 13 2
16 16 10 9 3 1 9 13 13 15 9 12 9 1 15 9 2
14 15 4 10 9 1 10 9 1 11 2 11 7 11 2
6 11 13 3 11 4 2
9 10 12 9 13 3 3 0 3 2
21 0 11 13 3 1 0 9 7 13 10 9 1 15 9 2 15 9 15 0 13 2
11 2 15 13 0 0 2 2 13 8 0 2
8 3 13 11 11 1 11 4 2
17 11 2 15 3 13 16 15 13 9 0 3 1 10 9 4 4 2
27 10 9 4 3 4 1 10 9 1 3 10 9 7 1 10 0 9 0 9 2 0 9 1 3 10 9 2
12 8 13 13 10 1 0 9 13 9 4 4 2
31 11 13 12 9 3 1 10 2 9 2 1 10 9 2 13 1 10 0 9 8 11 2 3 2 10 0 9 0 4 4 2
16 10 9 13 4 4 1 10 3 3 0 9 13 9 7 9 2
3 11 13 2
9 9 1 0 9 2 8 1 9 2
3 0 9 2
4 2 9 2 2
3 10 9 2
2 9 2
19 10 9 1 10 11 4 1 10 0 9 1 9 2 3 10 9 3 13 2
17 3 13 3 10 0 9 1 13 9 2 3 3 0 9 13 4 2
26 2 16 10 9 0 4 2 13 15 1 10 9 3 1 0 9 10 9 0 9 4 2 2 3 8 2
10 9 1 10 11 4 3 3 0 4 2
12 1 10 9 1 11 13 3 3 3 9 3 2
26 1 11 7 11 4 1 10 9 10 9 1 10 9 4 2 3 1 10 9 7 1 10 9 1 11 2
38 11 13 15 9 0 4 2 2 9 13 10 9 1 2 2 16 15 0 13 4 16 10 9 3 1 10 9 4 4 7 3 1 10 9 13 4 2 2
12 16 15 1 13 4 13 11 1 10 0 9 2
8 10 2 9 2 4 10 9 2
16 11 13 4 2 3 13 15 9 4 16 15 15 1 9 13 2
5 7 3 1 11 2
23 2 1 11 13 10 9 9 4 2 7 1 11 13 15 15 1 9 4 2 11 2 2 2
8 3 4 10 9 9 0 0 2
9 10 9 4 1 10 13 9 4 2
40 1 12 9 1 10 0 9 13 11 10 9 1 11 8 1 10 9 7 4 10 9 1 0 13 1 8 2 15 10 0 13 9 13 2 1 10 12 9 4 2
24 16 10 11 0 1 9 8 9 2 13 3 1 10 9 0 9 2 15 1 10 9 4 4 2
18 1 12 9 4 11 0 10 0 9 1 9 1 10 9 1 10 9 2
9 11 13 1 10 0 9 1 11 2
16 10 9 1 11 7 11 4 1 10 0 0 9 1 11 4 2
15 11 13 0 9 16 1 10 0 9 1 9 8 1 13 2
12 11 13 0 1 10 9 1 10 9 1 8 2
16 1 10 9 1 11 13 10 9 11 0 0 16 2 8 2 2
25 1 15 9 7 1 15 1 2 10 0 2 5 16 15 15 3 1 10 9 13 5 13 15 15 2
25 2 8 2 13 15 10 9 11 3 16 15 1 15 9 16 9 1 10 11 0 9 7 9 13 2
20 10 9 1 10 9 1 0 9 13 1 9 1 10 9 1 10 9 1 9 2
20 15 13 10 0 9 4 2 3 16 4 9 8 10 0 9 1 15 9 4 2
21 15 13 3 13 9 1 9 1 10 12 9 1 11 7 11 7 1 11 7 11 2
36 12 9 13 0 0 7 4 3 8 1 10 9 16 15 12 1 15 13 1 10 0 9 1 0 15 9 3 13 7 15 9 3 3 13 4 2
17 2 13 15 15 4 2 13 3 3 12 1 11 1 0 9 2 2
8 1 15 9 4 10 9 4 2
21 8 13 10 9 1 11 4 7 15 13 3 15 9 4 3 10 0 3 1 4 2
26 3 13 15 10 9 7 9 0 4 1 15 9 2 3 1 15 10 15 11 0 1 15 9 13 4 2
21 15 13 15 3 0 8 0 1 4 4 7 16 9 1 10 15 13 9 1 4 2
10 10 9 11 1 11 13 10 15 9 2
6 10 9 1 15 8 2
14 10 9 1 10 9 13 1 10 0 9 4 1 4 2
22 3 13 10 9 1 10 0 9 2 3 10 11 0 13 4 1 15 9 1 15 8 2
19 10 9 11 13 5 16 15 3 13 5 1 8 7 4 1 12 9 13 2
18 15 8 15 9 9 7 13 1 10 9 4 1 15 10 0 13 9 2
9 13 9 11 13 10 9 11 4 2
16 15 13 1 9 1 10 0 9 13 1 11 10 9 1 4 2
30 15 9 13 3 9 1 0 9 2 16 10 9 16 9 9 4 7 3 16 15 1 10 9 13 2 10 9 1 13 2
15 10 0 9 13 3 10 9 1 9 4 2 8 10 9 2
10 0 12 9 7 9 13 3 3 4 2
10 10 9 4 4 1 10 9 1 11 2
20 2 10 0 2 0 10 9 0 2 9 2 1 15 3 9 1 9 13 2 2
24 10 9 1 10 11 1 10 1 11 13 9 7 10 9 2 3 15 9 4 4 2 4 0 2
22 3 13 10 9 8 1 12 0 1 10 0 9 15 8 2 16 15 9 12 9 4 2
14 3 4 0 4 2 16 15 15 16 10 0 9 4 2
32 10 9 11 13 15 9 16 9 1 10 9 7 15 4 3 3 1 3 15 0 2 16 15 3 4 13 15 9 3 1 4 2
14 1 8 13 15 10 9 1 11 7 11 4 7 4 2
5 3 8 7 11 2
22 3 13 15 4 1 10 1 10 0 9 13 13 9 8 2 16 10 9 1 9 13 2
14 10 0 9 2 15 0 10 9 1 15 13 0 4 2
11 10 11 4 10 9 3 15 15 13 4 2
19 1 10 9 0 1 10 9 13 7 10 0 9 13 15 10 0 9 4 2
46 10 9 1 10 9 11 13 2 13 1 15 3 0 9 1 4 2 16 10 9 3 0 4 4 1 16 9 16 15 1 10 0 9 3 4 4 4 7 3 10 0 0 9 4 4 2
27 15 4 1 15 9 1 16 10 9 11 1 11 13 1 10 9 1 13 1 15 9 1 9 1 15 9 2
9 7 15 13 3 1 10 0 11 2
25 16 15 1 10 9 4 4 4 3 15 0 9 0 4 7 3 4 15 9 1 15 9 4 13 2
17 1 10 13 12 9 13 3 0 3 12 1 12 9 0 9 4 2
27 10 1 10 9 0 9 1 0 9 1 10 0 9 2 3 1 10 9 10 9 13 2 13 1 10 9 2
12 1 10 0 9 13 1 10 9 3 0 9 2
40 9 13 11 1 8 9 11 16 9 8 2 3 1 9 13 3 1 12 7 12 9 10 0 9 1 10 9 11 1 8 1 8 9 11 2 11 8 9 11 2
15 11 13 3 10 9 9 3 1 10 0 9 1 12 9 2
27 10 0 9 9 1 10 9 2 10 9 1 12 9 2 3 10 0 11 15 3 13 4 1 15 0 8 2
16 15 4 1 10 0 9 3 0 7 13 3 1 11 0 9 2
13 8 13 3 1 15 9 9 3 3 1 10 9 2
14 8 8 9 7 9 2 8 1 15 1 9 7 9 2
24 15 4 1 15 9 2 16 10 9 11 13 1 10 0 9 3 11 7 11 1 9 4 4 2
13 15 13 4 2 7 9 8 13 15 9 0 8 2
38 9 11 1 11 7 10 0 9 11 13 15 13 9 11 2 12 2 1 11 2 10 12 9 13 9 1 10 11 2 15 0 3 1 11 7 11 13 2
36 10 9 3 4 3 1 10 0 9 1 10 13 9 1 11 4 1 10 0 9 2 16 9 11 15 11 0 13 4 9 11 1 11 1 4 2
53 9 11 2 8 2 13 13 9 10 9 1 15 8 4 1 10 9 1 10 11 2 3 3 4 4 10 13 9 3 1 4 2 9 7 0 9 3 1 4 1 15 8 7 10 9 1 10 0 9 3 1 4 2
24 2 15 4 0 16 1 10 0 9 1 10 9 15 9 1 9 4 4 2 2 3 9 11 2
14 2 15 13 16 10 11 1 10 0 9 4 4 2 2
16 3 13 15 3 3 3 16 10 11 1 10 13 9 13 4 2
2 8 2
20 15 13 15 3 2 7 16 15 3 4 2 3 4 10 9 3 3 0 3 2
25 1 10 0 9 13 15 1 9 7 3 13 15 13 15 3 15 15 1 0 13 9 1 10 9 2
26 16 15 9 15 1 11 0 7 8 1 15 8 13 4 1 10 9 1 11 1 10 9 1 10 11 2
13 15 13 3 3 16 10 9 0 1 15 13 4 2
8 13 3 3 15 3 3 3 2
30 10 9 13 7 13 3 3 1 11 1 10 9 7 15 4 3 10 0 9 1 15 15 1 11 3 3 0 1 13 2
11 3 13 3 15 2 16 15 3 3 13 2
21 15 4 10 9 2 15 10 9 9 8 13 4 16 11 3 3 1 11 1 13 2
20 3 13 3 0 15 0 9 4 2 7 1 11 13 15 0 3 4 4 4 2
35 10 0 13 9 1 0 12 9 0 2 15 1 10 11 1 10 11 1 9 15 9 13 4 2 13 3 9 4 1 12 12 9 0 9 2
18 15 9 13 1 10 11 2 7 13 8 4 1 10 9 1 10 11 2
19 15 13 10 12 9 3 3 1 4 2 7 15 1 10 11 3 1 4 2
27 10 9 13 3 4 16 1 15 13 1 10 0 9 8 10 9 15 9 4 4 4 16 1 10 0 9 2
48 16 8 15 9 3 0 4 4 2 7 8 15 9 10 9 13 4 2 13 15 15 9 4 4 4 1 15 15 2 10 9 1 10 9 2 7 2 11 11 9 1 11 2 13 4 4 4 2
26 13 10 9 3 4 10 9 1 9 8 10 0 9 3 4 4 2 2 13 10 0 9 1 10 9 2
27 16 13 2 13 1 9 1 9 10 0 1 10 9 12 2 15 1 12 3 3 4 4 1 15 0 9 2
8 7 15 4 1 15 15 4 2
27 10 9 4 2 16 10 9 1 10 9 1 10 11 3 3 13 4 16 10 9 1 15 9 3 1 13 2
16 10 9 13 3 10 0 9 4 15 4 4 1 10 0 9 2
29 15 13 3 1 10 9 1 10 9 4 7 15 13 3 2 16 15 9 3 1 15 9 13 4 2 15 9 3 2
6 3 4 15 3 4 2
13 16 1 11 0 9 10 9 13 1 11 11 11 2
15 10 9 13 1 10 9 1 11 11 11 3 3 15 3 2
13 7 12 9 0 13 10 9 1 11 1 15 9 2
27 1 10 9 1 9 11 13 10 9 10 9 1 10 0 9 1 2 8 2 3 1 10 0 7 0 9 2
22 1 10 9 12 9 2 13 2 16 15 4 13 10 9 1 10 0 9 3 1 4 2
4 10 0 9 2
25 10 0 9 1 10 2 9 2 1 10 9 1 11 7 11 2 3 10 9 15 3 1 13 13 2
23 1 10 9 1 10 9 1 9 1 15 9 13 9 7 9 4 4 4 7 9 4 4 2
37 16 1 8 0 1 12 15 9 1 10 9 4 4 2 13 10 9 0 3 2 16 10 9 0 4 2 3 15 15 13 4 1 0 1 13 13 2
17 1 3 4 10 9 4 1 10 9 3 1 15 13 1 10 9 2
28 10 0 9 13 3 10 9 1 10 9 15 1 10 9 1 11 1 11 1 11 13 8 9 1 9 2 4 2
11 15 4 10 0 9 8 1 10 0 9 2
21 1 10 9 1 10 11 13 15 10 0 9 8 1 11 1 10 9 1 10 9 2
14 8 4 0 13 1 10 11 4 2 3 0 4 4 2
36 3 0 7 0 16 10 9 2 16 15 0 10 0 9 4 2 3 1 15 2 16 15 3 3 13 4 7 0 15 9 1 4 13 4 4 2
9 10 9 13 3 3 3 1 9 2
12 2 15 12 2 12 9 4 15 3 3 0 2
14 3 13 1 9 4 4 2 1 9 2 9 2 9 3
16 7 15 13 15 3 3 10 15 9 16 3 15 0 13 2 2
19 16 9 7 3 10 9 0 4 13 4 2 13 10 9 3 3 0 8 2
15 10 9 8 2 12 2 2 9 1 15 0 8 2 13 2
29 2 15 1 15 13 15 1 10 0 12 9 2 3 15 8 12 9 1 15 9 13 4 7 10 11 12 9 2 2
32 16 10 9 1 11 7 11 1 10 9 1 10 9 1 10 9 3 3 0 4 4 2 13 3 0 16 3 10 9 4 4 2
20 16 10 9 8 13 2 13 11 10 9 11 4 1 11 1 10 9 1 9 2
30 10 9 13 3 1 12 9 1 15 13 1 10 9 4 4 2 15 10 0 9 1 10 9 1 10 9 3 13 4 2
12 1 10 11 1 8 13 10 9 1 8 8 2
40 12 13 9 1 9 1 15 8 2 9 2 1 0 9 1 11 13 1 10 13 9 1 10 0 9 9 4 1 10 9 1 15 15 7 15 9 1 10 9 2
32 1 10 9 4 4 1 10 13 7 9 1 10 9 2 15 13 1 9 16 13 9 3 1 1 4 7 15 0 13 1 9 2
12 8 10 9 4 10 9 4 2 15 3 13 2
14 10 9 1 15 0 8 1 11 2 11 2 4 4 2
30 15 0 8 1 11 13 3 1 10 9 1 11 4 1 10 9 1 8 10 9 1 10 0 9 1 4 4 7 4 2
11 11 4 3 4 1 10 0 9 1 9 2
9 15 4 4 1 15 8 1 11 2
17 11 4 0 9 11 4 2 13 1 9 1 10 0 9 1 11 2
35 10 9 1 3 12 0 9 7 9 2 15 1 10 13 9 9 1 9 1 8 2 11 2 13 2 13 0 16 10 13 9 1 4 4 2
5 16 0 1 4 2
20 2 8 2 2 13 1 10 9 1 8 7 12 9 3 13 8 10 0 9 2
26 15 4 3 12 15 9 13 4 2 15 12 15 4 3 1 12 2 16 1 10 12 9 3 12 13 2
21 10 0 9 13 1 10 0 9 1 10 12 9 2 15 4 4 1 10 0 9 2
20 10 13 11 1 10 0 9 2 15 15 9 3 0 16 0 13 2 4 8 2
12 1 12 9 4 15 9 1 10 0 9 11 2
24 15 4 3 12 9 0 2 9 1 10 9 1 10 9 1 11 7 9 1 15 8 1 11 2
17 1 12 13 15 10 0 9 1 10 0 0 11 2 1 16 9 2
29 2 10 0 9 1 10 9 2 2 15 15 10 9 1 11 7 10 0 9 1 10 0 9 1 10 15 9 13 2
24 10 9 11 1 10 11 2 9 9 1 15 0 2 13 10 0 9 1 10 9 8 13 4 2
15 1 9 13 3 3 15 4 4 2 16 10 0 9 13 2
19 10 9 1 10 9 2 13 1 10 9 11 1 11 2 4 4 1 8 2
25 16 15 1 10 11 11 1 13 9 3 3 13 1 9 2 3 13 15 1 15 9 4 1 9 2
21 10 9 13 0 3 3 15 16 8 4 2 16 10 9 1 0 9 13 4 4 2
29 1 10 11 13 8 3 15 0 9 1 11 2 3 4 1 11 10 0 11 4 2 1 12 9 13 9 8 4 2
25 10 9 1 10 9 2 3 3 8 9 8 13 2 4 4 1 10 9 8 1 11 7 9 8 2
15 8 13 3 10 9 9 2 15 4 4 1 0 0 9 2
21 1 10 1 12 9 13 9 4 12 2 9 2 4 2 13 1 15 9 7 9 2
6 1 3 10 9 11 2
26 3 10 9 1 15 0 9 1 11 2 10 3 0 0 9 2 15 3 4 4 1 9 3 2 8 2
31 15 13 16 10 0 9 1 9 3 4 1 9 2 7 15 13 3 0 3 16 10 9 2 1 15 2 0 7 0 4 2
11 2 7 3 0 7 0 2 2 13 15 2
12 15 13 1 0 9 4 1 15 1 10 9 2
36 10 9 13 12 9 2 8 10 9 1 0 9 7 9 7 3 10 9 1 10 9 1 10 12 9 2 15 3 15 4 4 1 10 0 9 2
8 2 3 4 15 4 7 4 2
34 1 10 11 1 11 13 3 1 8 9 11 15 0 9 7 15 0 9 2 10 9 1 10 9 8 2 0 1 10 9 1 10 9 2
9 10 9 4 8 1 10 9 4 2
13 1 10 9 13 10 9 3 15 0 9 1 3 2
15 15 13 16 15 9 1 9 4 4 7 3 0 4 4 2
26 15 9 13 3 4 0 9 11 12 0 9 1 0 9 1 10 9 1 4 4 7 3 1 4 4 2
16 10 0 9 13 15 3 3 4 16 3 1 10 9 1 4 2
17 15 1 10 12 2 13 2 9 13 9 4 1 11 3 1 4 2
29 15 13 10 9 8 4 16 10 0 9 1 13 16 15 1 11 1 12 0 9 8 4 4 7 1 9 4 4 2
13 10 0 9 4 13 1 10 3 0 9 1 9 2
49 9 8 15 1 15 9 1 11 3 13 4 1 12 8 1 11 7 1 10 9 10 9 1 10 10 9 1 8 4 2 13 15 13 1 15 11 16 10 0 9 1 10 1 10 13 9 13 9 2
9 1 13 9 13 3 9 13 4 2
16 10 9 1 10 9 9 1 10 9 4 3 1 4 1 9 2
32 10 0 9 13 3 3 0 1 15 9 4 16 1 10 15 9 0 4 15 9 1 15 13 1 15 9 4 7 10 9 4 2
21 10 0 9 13 1 10 0 9 2 8 2 3 3 10 9 1 10 9 4 4 2
36 10 9 1 10 9 13 3 3 15 10 9 1 10 0 9 1 10 11 15 2 3 13 15 2 1 12 2 0 2 10 9 1 10 11 13 2
41 15 13 3 3 0 3 2 7 3 13 1 15 9 2 3 1 15 13 1 10 9 2 1 9 11 9 3 15 9 1 10 11 2 7 8 10 9 1 10 11 2
33 7 9 11 2 16 15 10 9 13 1 11 1 4 2 13 1 10 9 15 0 15 15 10 11 3 7 15 8 3 1 9 13 2
36 11 4 0 2 15 4 0 2 15 13 10 0 9 1 10 0 9 2 7 15 13 11 9 7 11 9 2 7 15 13 10 3 0 9 3 2
19 15 0 9 4 1 10 0 9 3 3 0 16 10 0 1 15 13 9 2
22 7 15 13 15 3 2 7 3 8 13 4 4 3 3 3 0 7 13 3 3 9 2
10 15 2 0 9 2 13 15 9 4 2
30 2 0 4 3 10 0 9 1 15 8 1 9 7 10 9 1 9 2 7 10 9 4 3 3 3 3 3 0 3 2
19 1 10 13 9 7 9 13 15 10 9 7 0 9 16 13 9 1 13 2
5 10 9 4 4 2
27 15 13 3 3 1 10 9 7 9 10 9 4 16 3 3 1 13 4 7 15 1 9 7 9 1 13 2
27 10 9 7 10 9 2 3 1 15 13 0 1 13 9 7 15 0 13 9 2 13 1 10 9 4 4 2
10 1 15 9 13 12 9 7 12 9 2
28 10 9 13 3 1 10 0 9 4 4 7 3 4 3 7 1 10 9 7 1 10 9 10 9 7 9 4 2
16 10 9 1 15 1 10 9 0 9 13 3 1 10 13 9 2
20 1 9 8 1 15 8 1 11 13 12 10 9 4 4 1 15 3 13 8 2
13 10 9 13 1 15 9 15 9 7 15 9 4 2
31 0 4 1 10 9 1 10 9 2 10 0 9 2 10 9 7 9 2 10 9 7 9 2 7 10 9 1 10 9 4 2
8 15 0 9 4 0 0 4 2
14 10 9 13 3 3 9 4 1 11 2 11 7 11 2
31 15 8 4 1 10 0 9 1 15 9 4 1 8 2 9 1 15 8 1 9 7 9 2 1 15 0 9 1 10 9 2
16 10 9 13 3 1 10 9 1 11 2 3 13 10 11 3 2
20 10 9 4 10 9 1 10 9 7 10 0 11 9 2 7 4 0 9 4 2
50 10 9 8 2 12 2 1 11 2 9 1 0 9 1 15 8 2 9 7 9 1 11 7 9 1 10 0 9 2 4 1 10 9 4 16 9 1 10 0 9 2 1 9 8 2 1 10 9 8 2
18 10 11 13 0 3 10 0 9 2 8 10 9 1 10 9 1 11 2
29 1 15 9 2 15 0 4 4 1 8 2 11 2 4 10 9 8 2 9 1 15 8 1 11 2 1 3 4 2
30 16 10 9 1 10 9 11 1 10 11 10 13 9 0 1 4 13 1 10 0 9 2 13 3 3 0 9 1 4 2
16 0 3 1 10 9 13 8 1 10 0 9 12 1 10 9 2
9 10 9 13 3 3 12 9 0 2
13 15 8 13 10 9 1 12 0 4 1 12 9 2
21 1 10 9 13 11 1 12 15 9 1 10 9 1 8 7 10 13 9 1 11 2
12 10 9 1 15 9 13 3 3 15 9 3 2
19 4 4 16 15 9 9 13 1 10 9 16 15 0 1 9 7 9 4 2
12 3 10 9 1 13 9 4 15 8 1 4 2
11 15 4 3 10 9 16 10 9 4 4 2
33 9 15 10 9 13 16 1 10 13 9 1 9 1 4 7 10 13 9 3 1 9 1 4 13 3 1 15 9 3 4 1 4 2
33 15 8 13 1 10 0 9 8 1 11 2 11 2 4 1 10 0 9 2 8 2 15 4 4 1 11 2 3 13 1 15 8 2
19 10 9 1 10 9 4 10 9 1 7 10 9 1 9 1 10 0 9 2
14 10 9 13 4 4 1 10 9 11 7 8 1 11 2
7 8 13 4 1 10 9 2
13 1 12 4 12 9 4 7 1 12 3 12 9 2
7 10 9 13 4 1 8 2
25 10 0 9 7 15 9 4 0 8 11 1 10 9 11 8 1 10 9 1 10 9 1 10 11 2
19 10 13 9 2 15 1 9 1 15 8 4 4 2 13 1 12 4 4 2
29 16 15 13 1 10 9 7 15 13 1 9 1 10 9 13 3 15 13 1 12 9 9 1 10 9 1 10 9 2
17 1 15 9 13 10 9 3 3 10 9 9 8 15 12 9 4 2
17 1 11 1 10 0 9 3 4 8 1 10 0 9 13 8 4 2
23 7 1 9 1 0 9 15 10 9 1 15 9 0 9 13 4 2 4 15 3 8 4 2
28 10 0 9 4 3 0 3 16 10 9 1 10 0 9 1 15 9 13 9 1 11 1 11 1 11 4 4 2
49 8 2 12 2 13 1 15 10 9 10 0 9 13 2 10 9 4 10 9 0 7 10 9 4 3 0 2 16 3 15 7 3 0 13 1 10 9 1 8 2 1 10 9 1 10 9 1 11 2
26 7 3 1 9 2 12 9 2 4 15 10 0 9 1 4 2 10 3 0 9 1 10 11 1 3 2
24 10 9 13 1 10 13 9 1 8 12 3 3 15 0 3 16 15 8 12 1 10 13 9 2
22 3 13 15 3 2 13 8 10 9 11 3 10 9 1 10 9 7 10 0 0 9 2
11 1 10 10 15 9 4 3 15 9 3 2
6 3 4 13 8 0 2
4 10 9 13 2
22 2 15 13 16 3 15 9 3 13 1 10 9 7 3 13 10 9 1 9 7 9 2
10 15 13 1 12 9 1 10 9 2 2
6 10 0 9 4 0 2
19 13 10 9 1 10 9 2 7 15 13 3 3 1 15 12 1 10 9 2
17 10 0 9 4 3 3 1 0 9 7 15 9 4 9 1 11 2
17 3 15 3 16 0 9 1 10 11 1 10 9 1 9 4 4 2
31 16 1 10 9 11 10 9 1 9 0 4 2 13 3 10 0 0 9 1 10 9 4 4 1 8 2 3 12 2 12 2
2 11 2
27 2 15 4 10 9 15 15 3 0 4 4 7 15 13 0 16 15 10 11 0 3 3 10 0 9 13 2
14 15 4 0 15 9 3 1 3 9 1 9 7 9 2
12 1 10 9 1 10 9 10 9 10 9 13 2
16 9 2 9 7 9 13 7 10 0 12 9 1 10 9 13 2
6 10 9 0 0 13 2
19 10 13 9 1 12 9 9 7 12 9 13 9 13 7 3 9 3 13 2
2 9 2
22 13 0 9 1 10 9 1 9 2 9 2 3 10 13 9 2 9 2 9 7 9 2
2 9 2
42 2 16 15 3 15 9 13 2 4 15 15 0 2 16 3 9 4 1 9 2 2 13 3 10 9 1 10 9 2 15 3 12 9 1 15 0 8 13 1 10 9 2
15 9 9 2 1 10 9 1 9 2 9 2 9 7 9 2
22 1 11 13 10 0 9 8 15 3 0 0 2 11 7 15 9 9 13 3 10 9 2
27 15 4 8 4 16 15 9 15 9 1 10 9 7 15 9 13 2 7 15 13 10 9 7 3 10 9 2
28 10 9 4 2 1 11 2 3 15 0 4 16 15 10 9 9 4 4 4 2 7 16 9 13 15 15 3 2
15 3 13 1 8 1 10 9 1 12 1 11 10 13 9 2
6 10 0 9 4 8 2
4 10 0 9 2
17 1 15 9 9 13 10 9 1 9 1 9 2 1 9 1 9 2
12 0 4 3 4 3 0 15 13 4 1 11 2
17 1 10 9 1 12 1 12 9 1 9 13 15 1 12 3 4 2
23 1 10 9 2 3 1 10 9 1 15 8 2 4 12 9 4 2 15 15 0 4 4 2
10 10 9 13 3 2 16 15 9 13 2
15 15 9 2 1 11 9 2 4 10 9 1 15 15 13 2
19 1 10 9 1 10 9 13 3 0 10 9 1 10 9 16 9 1 9 2
32 16 15 1 10 0 9 9 13 4 13 10 9 2 10 0 9 2 3 3 3 0 1 4 7 13 15 1 10 9 4 4 2
12 3 13 3 1 15 9 1 0 9 9 4 2
14 10 9 1 10 9 9 4 10 0 9 8 0 4 2
34 1 8 3 4 15 1 10 9 1 10 11 1 11 4 1 15 0 8 1 11 2 15 15 8 10 9 1 15 9 13 1 10 9 2
19 11 11 13 3 1 10 9 10 9 1 10 9 0 4 15 13 1 4 2
8 10 9 13 10 9 1 4 2
11 15 13 9 3 1 4 2 7 13 3 2
36 0 4 2 16 16 10 9 3 13 2 7 1 10 9 2 7 1 10 9 9 13 2 16 1 10 9 1 10 9 15 1 9 4 1 4 2
6 8 4 10 13 9 2
45 1 10 9 1 8 2 3 15 13 1 15 9 1 11 2 1 15 15 12 9 13 2 13 11 10 13 9 10 13 9 2 3 15 15 9 1 10 9 1 10 9 10 9 13 2
12 3 13 8 10 9 1 10 9 1 10 9 2
5 2 0 9 2 2
20 11 13 1 15 9 15 9 1 10 13 9 2 3 15 3 3 0 13 4 2
8 3 13 10 9 3 10 9 2
29 7 3 4 15 3 0 16 10 9 16 10 9 1 15 1 4 2 3 1 10 9 2 1 3 1 10 9 4 2
24 11 4 3 1 10 9 1 10 11 4 7 15 13 16 15 8 15 3 3 0 0 4 4 2
15 16 11 13 4 1 10 0 9 3 13 15 3 0 4 2
27 8 12 9 1 13 9 4 3 1 10 11 4 4 1 10 9 7 15 13 13 1 10 9 8 1 11 2
44 10 0 9 4 16 10 0 9 2 15 1 8 4 4 2 10 0 9 1 12 0 9 1 9 4 13 16 9 7 9 3 1 13 7 1 10 9 15 0 9 3 1 13 2
7 10 0 9 1 12 9 2
17 1 10 15 9 15 9 2 1 10 15 13 10 9 1 9 0 2
13 8 2 9 1 10 11 2 9 7 9 1 9 2
8 2 15 13 10 9 0 3 2
7 7 15 13 3 3 3 2
40 16 10 9 1 15 13 9 3 0 13 4 2 15 4 0 4 2 4 15 9 3 1 4 1 10 9 1 10 0 2 10 9 13 2 9 16 0 3 13 2
17 3 13 15 1 4 1 10 0 13 2 9 2 1 10 0 9 2
23 13 1 15 0 9 16 8 7 8 4 10 0 9 1 10 9 0 7 4 15 3 4 2
18 15 0 13 8 13 3 4 4 16 0 16 1 4 1 9 7 9 2
12 0 9 13 3 3 0 1 10 9 4 4 2
11 15 13 1 0 2 0 2 0 7 0 2
21 15 13 16 1 10 9 1 3 10 9 9 2 3 15 1 10 0 9 3 13 2
13 10 9 13 4 1 10 9 1 10 0 13 9 2
40 15 9 13 4 3 1 4 1 10 9 15 1 10 13 9 4 4 2 16 15 13 1 15 9 2 16 15 8 10 9 2 10 9 7 10 9 1 10 9 2
29 15 9 4 4 1 10 9 1 10 9 1 9 2 8 2 1 10 9 1 10 9 1 15 8 2 15 8 2 2
22 1 10 9 13 11 15 15 3 15 1 10 9 4 4 2 16 15 15 3 0 13 2
21 1 10 0 9 13 15 3 3 3 7 1 10 9 13 15 15 9 1 4 4 2
18 15 13 3 0 11 4 2 15 0 0 4 7 3 0 9 13 2 2
17 2 1 10 9 13 15 15 9 0 4 1 10 9 1 10 11 2
9 15 13 15 4 16 15 1 13 2
36 16 10 0 9 2 8 2 3 3 1 15 9 8 7 8 0 4 16 10 13 9 8 1 13 1 9 13 3 10 9 8 2 8 2 8 2
20 9 2 16 8 3 1 10 0 9 1 10 9 1 11 1 10 9 4 4 2
5 3 3 10 9 2
34 7 1 10 0 9 1 10 0 9 13 3 10 0 0 9 15 9 2 7 10 0 9 13 15 0 9 2 8 2 3 1 15 9 2
32 8 2 0 9 9 1 11 2 13 3 1 10 9 1 11 3 15 8 1 10 0 9 1 11 4 2 13 1 10 9 9 2
24 10 9 1 8 13 1 15 9 11 0 9 4 1 10 9 8 2 9 1 10 9 1 11 2
4 8 4 0 2
17 10 0 9 13 10 9 1 10 9 3 1 12 9 9 1 11 2
11 8 13 1 15 9 0 3 10 9 4 2
14 10 9 4 3 3 15 16 10 9 7 13 10 9 2
10 12 9 1 10 9 13 11 10 9 2
15 1 10 9 1 10 9 13 10 9 1 10 9 1 11 2
3 9 12 2
18 15 13 1 10 0 9 3 10 9 1 15 12 1 12 9 1 9 2
19 1 10 9 13 11 10 9 9 2 7 9 11 1 8 13 10 0 9 2
26 10 9 1 15 9 4 15 1 10 0 9 15 1 10 9 1 10 11 11 13 1 10 13 0 9 2
18 10 9 13 3 2 16 15 15 9 9 4 2 15 8 3 4 4 2
54 15 13 3 9 4 1 10 9 2 13 1 10 9 11 2 11 2 2 11 2 11 2 7 11 2 11 2 1 10 9 2 3 4 4 16 2 10 9 10 0 9 4 4 1 9 1 10 1 13 9 13 9 2 2
33 15 4 15 1 10 0 9 1 10 9 1 10 9 3 9 3 1 13 2 15 4 15 1 10 9 1 10 9 1 15 9 0 2
16 7 3 4 15 0 1 15 9 9 15 0 1 10 9 4 2
23 10 15 9 2 15 1 15 16 0 4 4 2 4 10 0 9 1 9 1 8 7 15 2
10 10 1 15 9 13 9 13 15 3 2
3 15 4 2
20 8 2 12 2 2 8 2 12 2 2 8 2 8 7 8 2 15 12 2 2
25 16 10 9 1 8 2 8 2 3 0 13 2 13 10 0 9 1 9 7 9 1 12 4 4 2
34 10 9 2 16 10 0 9 7 10 0 9 15 3 10 9 1 10 9 1 15 9 4 4 2 13 15 0 10 9 1 12 1 4 2
13 3 13 7 13 10 9 3 10 9 1 10 11 2
33 16 9 1 10 9 1 15 9 13 15 8 10 3 13 9 8 4 2 3 10 9 13 1 10 9 1 12 1 10 12 13 9 2
21 15 0 9 13 1 2 6 2 1 10 9 2 7 10 9 13 15 3 3 13 2
17 9 11 13 15 3 1 8 1 10 9 10 0 9 1 10 9 2
7 10 9 4 3 1 4 2
38 10 13 9 13 10 9 8 16 15 3 3 10 9 4 7 15 9 7 9 1 11 3 3 13 4 2 3 16 13 2 15 9 2 15 3 3 0 2
22 15 13 2 15 9 16 12 4 15 4 1 15 9 16 3 10 0 9 1 12 4 2
14 1 9 15 15 3 13 13 15 15 15 3 3 4 2
9 3 16 9 3 8 1 4 13 2
23 15 13 3 1 9 2 15 1 10 9 5 0 5 4 4 2 16 3 3 15 3 4 2
19 15 9 13 3 3 1 10 9 7 1 9 1 9 1 0 9 4 4 2
7 1 10 9 13 9 12 2
5 11 13 15 3 2
9 2 0 13 2 6 2 9 2 2
13 6 2 13 10 2 11 2 2 15 4 0 13 2
8 11 13 3 3 3 1 4 2
18 15 9 13 1 15 0 9 7 15 13 1 15 13 1 15 0 9 2
15 2 6 2 15 13 15 4 2 7 15 13 3 4 4 2
11 10 9 13 15 3 3 3 0 16 0 2
13 7 15 13 3 3 10 0 9 4 1 10 9 2
14 10 0 9 1 10 13 9 13 10 11 3 4 4 2
16 2 3 13 15 3 3 3 9 3 2 15 9 12 9 13 2
7 7 15 13 8 6 2 2
27 0 4 10 9 1 8 2 13 1 10 9 2 15 1 10 13 9 3 3 3 15 9 13 1 15 13 2
7 2 15 13 3 1 15 2
7 3 13 15 15 0 3 2
6 13 3 3 15 3 2
19 0 8 13 15 0 9 7 3 2 7 3 4 10 9 3 3 3 3 2
20 1 15 0 9 13 15 3 1 10 9 4 16 1 10 9 1 11 1 4 2
10 3 13 3 1 11 3 10 9 3 2
14 1 11 4 15 0 10 0 7 3 0 9 1 13 2
12 15 13 13 3 15 9 1 10 9 4 4 2
16 1 10 9 16 3 3 15 15 9 4 2 13 15 7 13 2
12 2 15 13 10 9 1 15 9 10 9 4 2
6 3 4 15 0 0 2
11 3 3 13 0 8 10 0 9 9 3 2
23 15 4 10 1 11 3 0 9 2 3 1 10 9 11 10 9 0 3 1 10 9 13 2
28 10 3 0 9 8 15 1 8 7 12 13 4 16 3 0 1 10 9 10 0 9 1 0 9 13 1 13 2
34 1 11 1 11 7 1 11 1 11 4 10 9 3 15 9 0 4 16 10 9 13 4 1 10 9 15 8 10 9 7 9 4 4 2
20 3 13 10 11 10 9 3 1 10 11 10 0 4 15 3 1 10 9 13 2
17 1 11 13 3 1 10 9 3 15 9 1 10 9 4 4 4 2
10 7 16 9 13 15 3 3 3 3 2
30 10 0 11 13 13 9 2 1 15 16 10 13 9 1 10 9 10 9 13 2 16 10 1 11 12 13 9 4 4 2
12 2 10 9 1 10 13 9 4 3 15 0 2
29 15 8 13 10 9 2 3 1 10 9 2 16 10 0 9 3 15 15 13 1 10 9 4 7 3 3 15 13 2
27 11 8 2 15 1 10 12 15 0 9 1 9 2 13 3 3 7 0 3 0 4 10 9 1 15 8 2
23 10 9 1 10 9 1 11 2 8 2 13 10 9 2 15 15 3 1 15 13 15 4 2
10 2 6 2 15 13 3 3 3 4 2
19 0 13 15 3 9 16 15 0 4 2 7 15 13 3 15 15 9 3 2
24 10 9 1 10 9 4 0 3 0 2 16 15 3 16 0 9 15 3 3 3 13 4 2 2
25 9 8 2 12 2 7 9 8 2 12 2 1 11 13 4 3 0 10 9 1 10 9 3 4 2
15 10 15 9 4 16 10 9 15 3 3 0 3 13 4 2
42 13 4 2 16 10 11 10 9 13 16 10 11 2 3 3 2 16 10 11 3 3 3 0 4 1 4 2 16 10 11 3 10 9 1 8 3 3 16 10 9 13 2
36 10 9 1 15 0 0 8 1 11 13 3 3 15 9 0 4 4 2 16 9 8 1 10 0 9 15 0 9 1 15 15 0 9 13 4 2
6 15 13 3 3 3 2
3 15 13 2
29 9 2 3 10 9 1 15 9 13 3 3 0 3 4 7 13 16 10 11 4 16 15 2 3 16 15 2 4 2
30 10 13 9 13 0 10 0 9 2 7 15 1 10 9 4 3 3 3 13 2 16 10 9 2 8 12 0 2 13 2
10 10 12 15 9 4 1 10 9 4 2
11 10 9 13 3 16 10 9 3 1 13 2
13 10 9 4 3 0 9 8 4 15 9 1 4 2
9 1 8 13 9 4 4 1 9 2
13 15 8 13 10 0 9 4 1 10 9 0 9 2
29 1 10 9 13 1 10 13 9 15 13 3 1 9 1 0 9 7 9 4 4 10 9 1 10 9 3 1 4 2
32 3 13 10 9 11 0 9 7 10 9 15 9 3 4 4 1 10 0 9 2 1 10 9 13 2 16 11 9 8 3 13 2
25 0 13 10 9 1 15 9 1 9 1 12 7 12 4 4 2 1 9 1 10 9 1 10 9 2
25 1 10 9 13 3 9 1 4 4 1 9 2 9 2 9 7 9 2 1 10 9 2 11 2 2
33 10 0 13 0 9 8 1 11 4 3 1 15 2 8 2 2 10 0 9 1 11 2 1 10 9 4 1 15 13 1 10 9 2
22 16 3 0 10 9 4 4 7 4 13 11 1 10 9 1 10 9 11 1 11 4 2
11 10 9 13 15 3 0 0 1 8 8 2
17 10 9 11 13 1 9 1 10 9 0 9 1 10 0 9 4 2
10 15 13 15 1 15 9 15 13 9 2
20 0 4 15 3 3 4 2 15 15 9 4 2 16 13 10 9 15 3 4 2
24 16 15 15 9 3 3 4 13 4 15 1 9 7 9 1 15 2 15 13 4 1 15 9 2
14 4 15 3 3 2 1 0 9 2 2 16 15 13 2
18 1 10 15 9 4 3 1 10 0 9 10 0 13 9 7 9 0 2
40 10 9 1 8 2 8 2 13 0 9 1 10 9 7 9 1 9 4 16 0 3 1 13 2 16 10 9 15 3 1 15 9 13 4 1 9 3 1 4 2
3 3 3 2
20 10 9 15 15 9 1 10 9 13 2 15 13 16 9 7 16 9 15 9 2
33 3 13 10 0 9 11 1 10 9 1 10 9 15 9 3 4 4 1 11 2 16 10 0 9 3 1 15 3 13 9 13 4 2
38 8 2 9 1 15 8 2 13 3 1 10 9 1 10 9 1 11 15 9 4 1 15 3 4 4 16 10 9 1 10 9 13 1 10 9 1 8 2
45 9 8 2 8 2 13 1 10 9 1 15 8 4 16 15 4 16 10 9 1 10 9 1 0 9 1 12 3 3 4 4 16 3 15 9 4 4 1 10 0 9 1 10 9 2
21 10 9 13 1 15 9 0 4 1 10 9 1 10 9 16 16 3 9 4 4 2
24 10 13 9 13 3 1 3 8 10 9 4 1 10 9 1 10 9 1 15 8 1 15 8 2
28 15 4 0 4 1 10 9 1 3 12 9 16 10 9 2 10 9 8 2 12 2 2 4 4 15 1 4 2
21 15 4 10 0 9 1 0 9 16 10 13 9 1 10 9 1 15 8 4 4 2
24 7 3 3 13 10 9 0 4 4 7 10 0 9 1 0 9 4 4 1 10 0 0 9 2
36 15 13 13 3 1 15 13 1 9 1 10 1 9 13 1 10 9 1 10 9 2 16 10 9 1 10 9 2 10 11 9 1 10 9 13 2
40 10 0 9 9 13 3 3 0 9 3 3 16 10 9 1 10 0 9 1 10 9 3 1 4 7 0 1 4 16 10 0 0 9 1 11 0 9 4 3 2
26 9 11 13 15 9 3 3 1 15 15 9 1 9 4 2 16 15 3 8 4 1 4 1 10 9 2
27 8 2 8 7 8 13 5 1 15 9 5 16 0 1 10 9 1 10 11 1 11 1 10 9 1 12 2
9 15 13 10 9 1 15 12 9 2
13 10 9 13 0 4 4 1 10 0 9 1 11 2
10 10 9 13 1 9 12 9 9 4 2
15 12 1 15 13 10 9 1 10 9 4 1 4 3 3 2
27 9 7 9 13 15 9 1 9 7 9 2 13 10 9 1 4 2 16 15 1 15 9 1 13 9 9 2
16 9 8 1 11 13 3 1 9 2 16 15 3 0 0 4 2
30 15 9 4 3 3 13 2 15 1 10 9 10 0 9 9 7 9 1 15 13 2 16 15 9 1 10 9 13 4 2
17 4 15 3 15 3 4 1 10 0 7 0 0 9 10 9 4 2
54 8 15 1 13 1 0 9 7 9 2 15 15 10 9 13 1 15 9 7 15 9 2 13 10 9 15 1 0 9 16 10 0 0 9 2 9 7 9 2 15 8 9 7 9 8 13 4 4 7 8 4 13 4 2
17 3 1 10 1 10 9 13 9 13 15 10 3 0 7 0 9 2
17 10 0 11 13 10 9 1 10 9 1 15 8 3 3 3 4 2
30 8 10 12 9 1 9 11 7 10 9 1 9 8 1 11 13 10 9 2 1 3 12 9 1 13 2 3 12 9 2
10 16 11 1 0 9 4 2 13 8 2
12 1 10 12 9 4 10 9 1 0 9 4 2
14 11 13 15 3 1 9 8 10 0 11 2 12 2 2
28 12 9 1 15 8 2 11 2 13 15 0 12 9 4 1 10 9 1 10 9 11 1 11 1 10 13 9 2
22 10 9 11 13 11 0 3 4 4 2 7 13 10 9 15 10 11 3 13 3 0 2
29 10 11 4 3 3 1 0 1 9 4 1 10 9 10 9 1 9 3 1 4 16 3 10 9 3 8 1 13 2
26 10 0 9 4 0 3 3 16 10 9 1 15 9 15 4 1 10 0 9 3 15 3 10 9 13 2
40 10 9 1 9 1 11 2 11 7 11 4 0 1 10 9 13 2 3 8 15 13 16 10 11 9 15 9 15 9 15 1 10 9 3 4 4 0 4 4 2
17 2 10 9 13 1 15 0 9 9 4 4 2 2 3 13 8 2
23 10 0 9 1 11 2 10 0 9 1 15 9 2 4 0 0 1 10 9 1 15 8 2
23 8 2 9 1 10 9 11 2 13 1 8 9 4 1 10 0 9 1 10 9 1 11 2
26 15 13 4 16 10 9 11 16 9 4 4 1 10 0 9 7 15 10 9 4 16 11 3 13 4 2
21 10 9 11 4 3 3 3 13 1 4 16 11 15 1 10 13 9 4 4 4 2
25 16 15 13 13 9 11 13 2 13 1 10 0 9 1 10 9 10 9 2 1 9 2 4 4 2
18 1 9 13 10 9 16 12 9 4 7 0 12 9 1 10 9 4 2
16 1 10 9 13 10 11 12 9 4 16 1 15 4 1 4 2
18 9 15 3 4 4 2 13 0 1 10 9 1 10 0 9 4 4 2
25 7 3 13 15 3 2 15 0 13 0 9 13 1 0 0 9 2 15 10 9 3 3 3 13 2
9 10 9 1 15 9 13 1 12 2
27 15 0 8 2 15 8 1 11 2 11 7 11 13 15 10 9 1 8 15 0 8 8 7 15 8 8 2
15 10 9 1 8 13 15 1 10 9 2 8 2 1 11 2
11 1 15 9 16 15 15 4 4 13 4 2
14 10 0 9 1 10 9 13 10 9 4 1 15 9 2
17 10 9 2 3 12 9 13 2 3 12 1 11 2 13 1 12 2
15 2 3 1 10 9 4 3 3 10 0 9 2 15 13 2
7 2 3 4 10 9 8 2
3 8 2 2
15 10 9 4 1 15 15 0 2 3 3 3 13 4 4 2
43 15 13 0 10 9 1 10 0 9 16 10 9 16 15 8 13 16 15 0 9 13 10 9 1 11 8 3 1 13 2 16 15 13 1 10 9 1 10 15 9 1 11 2
28 15 13 10 0 9 3 2 2 13 15 2 2 16 15 10 9 1 0 1 10 9 1 10 9 4 4 2 2
20 1 15 13 10 9 2 15 0 13 3 15 12 2 16 10 0 9 0 4 2
28 8 4 10 9 1 15 8 15 10 11 9 1 10 11 13 1 10 9 15 3 1 10 9 4 13 4 4 2
16 3 10 0 9 13 10 9 1 10 0 9 1 10 0 9 2
26 10 0 9 4 2 16 11 3 3 3 11 7 11 13 2 7 15 3 1 10 9 0 9 1 8 2
16 10 9 8 1 11 13 3 4 1 10 9 9 1 4 4 2
12 15 13 4 16 10 9 13 9 15 9 13 2
24 1 10 0 9 1 10 0 9 2 0 1 12 2 13 10 9 11 3 3 4 7 4 4 2
8 15 13 0 3 3 9 4 2
13 10 0 9 4 4 1 15 13 1 10 0 9 2
20 3 13 15 3 8 15 3 2 7 1 10 9 1 10 9 7 1 10 9 2
5 12 0 9 13 2
21 15 4 0 2 16 10 11 10 13 9 10 9 2 8 2 1 10 9 13 4 2
11 10 9 4 3 16 10 11 4 1 8 2
15 3 15 9 1 10 11 13 3 1 15 2 8 2 4 2
15 10 0 9 13 1 10 9 1 8 2 9 1 10 11 2
10 11 13 3 3 15 10 9 8 4 2
4 15 13 8 2
22 12 9 3 13 10 0 0 9 3 1 0 9 1 11 16 10 9 9 3 1 13 2
14 15 9 13 9 11 7 9 11 15 0 1 10 11 2
18 1 10 13 9 13 15 3 1 10 9 7 9 3 10 9 4 4 2
41 16 15 12 9 4 2 13 15 3 1 15 9 1 10 9 1 15 9 2 7 15 13 10 9 5 1 15 15 3 3 10 9 13 5 16 15 15 15 13 4 2
22 10 9 15 1 15 9 1 10 9 13 1 4 2 13 15 0 1 15 9 4 4 2
5 8 13 15 3 2
3 15 13 2
28 2 10 9 4 10 9 1 10 9 2 16 10 2 0 9 2 10 9 4 1 9 7 0 9 1 10 9 2
22 15 4 1 10 9 0 2 0 2 1 4 1 10 11 16 15 0 9 1 13 4 2
16 10 9 2 10 11 2 10 9 1 11 2 1 11 7 11 2
11 8 13 3 1 11 1 10 9 1 8 2
13 10 9 9 1 10 0 9 10 9 1 12 9 2
35 8 13 3 3 16 8 4 2 16 10 9 10 9 1 11 1 11 2 3 15 4 4 16 15 9 3 4 4 2 16 10 0 9 13 2
12 8 13 10 9 1 10 9 1 10 11 4 2
14 15 4 10 3 0 7 0 9 15 15 3 4 13 2
24 8 7 8 1 11 13 9 4 1 10 9 1 9 1 11 1 10 0 9 1 11 1 11 2
7 10 9 13 0 12 4 2
10 1 9 13 12 12 9 9 4 4 2
9 10 9 13 10 9 1 12 9 2
13 10 9 13 1 10 11 4 4 1 9 1 11 2
11 1 10 9 1 15 9 13 11 12 9 2
16 1 0 9 13 9 1 10 11 15 4 1 9 1 10 9 2
26 10 9 4 4 1 15 9 7 13 4 4 2 13 12 9 1 10 12 9 15 1 15 9 13 4 2
8 1 15 12 9 4 12 9 2
16 1 10 9 1 9 13 3 9 1 10 9 3 9 4 4 2
31 15 13 1 10 9 8 4 2 16 11 7 11 10 13 9 9 4 4 2 3 15 1 10 0 9 13 4 1 15 9 2
22 0 12 9 13 16 10 0 9 0 4 7 0 12 9 12 3 0 9 1 15 9 2
19 3 10 11 2 11 7 10 0 9 8 13 1 9 1 10 9 1 11 2
27 12 1 12 4 3 10 9 2 7 0 1 10 0 4 3 13 10 0 1 10 9 3 1 10 0 9 2
11 10 9 13 3 0 10 9 3 1 4 2
17 12 0 13 15 1 10 9 2 13 10 9 7 13 1 10 9 2
16 10 9 13 10 9 0 2 16 3 9 1 10 9 4 4 2
10 10 0 9 13 3 1 11 9 3 2
17 1 10 0 9 2 16 3 3 10 9 1 10 9 13 4 4 2
19 3 10 9 2 15 0 1 10 0 9 1 10 9 13 2 13 15 9 2
7 3 13 10 9 9 8 2
32 9 8 2 8 2 13 1 10 9 1 15 0 9 5 15 12 0 13 5 1 10 9 9 4 1 10 0 9 1 10 9 2
25 2 16 3 10 9 13 2 13 15 10 0 9 4 1 0 0 2 15 1 10 9 1 11 13 2
42 1 10 0 9 1 10 12 9 15 3 3 10 2 8 2 13 16 10 9 1 10 9 2 3 12 9 9 1 9 2 13 10 9 3 1 15 9 1 10 9 4 2
29 15 0 9 4 2 16 10 9 1 10 9 1 10 0 13 9 3 10 0 9 13 4 1 10 9 9 1 4 2
12 10 15 9 4 3 3 1 10 9 1 4 2
47 16 9 11 3 15 9 2 3 12 9 2 1 0 9 1 0 9 4 13 4 2 13 3 15 9 1 15 9 2 9 7 12 9 2 1 10 0 9 1 10 9 1 10 9 4 4 2
17 10 13 9 1 10 0 9 13 0 9 10 9 8 3 0 4 2
14 10 9 1 10 9 1 11 13 8 1 15 1 12 2
19 1 10 0 12 9 1 15 9 4 10 9 1 10 0 9 13 1 4 2
29 10 9 7 9 1 12 4 1 9 1 8 4 1 10 0 9 1 8 2 15 12 9 15 4 16 10 13 9 2
26 10 9 1 10 11 1 9 7 9 7 0 9 2 11 1 11 2 4 4 16 16 3 9 4 4 2
9 10 9 13 3 15 9 8 4 2
32 10 9 2 15 13 1 10 2 0 2 9 2 13 3 8 9 7 9 13 4 4 2 2 3 15 1 10 9 1 10 9 2
21 15 1 15 10 9 13 4 13 1 12 9 4 1 9 15 10 9 13 4 4 2
21 3 13 1 10 9 1 9 7 9 10 9 1 11 7 11 3 1 10 9 4 2
14 2 3 13 10 9 8 10 9 1 9 1 11 4 2
7 1 15 9 4 3 4 2
23 3 13 10 9 9 2 15 1 10 9 1 10 0 9 3 3 9 1 15 9 13 4 2
13 7 10 9 13 15 1 10 9 8 8 4 4 2
19 15 9 13 10 9 1 10 9 1 15 9 7 3 12 9 10 0 9 2
14 1 15 9 4 3 1 10 0 9 3 3 15 4 2
18 0 1 10 9 1 11 13 10 0 9 8 10 0 9 1 15 9 2
14 15 1 10 9 2 9 7 10 0 9 1 15 9 2
46 16 10 9 1 15 0 13 1 11 5 0 8 5 1 11 7 10 9 1 10 0 9 3 13 2 13 10 12 9 0 9 3 3 10 0 9 4 2 16 10 0 3 3 11 13 2
10 10 9 13 3 10 0 9 1 9 2
15 15 13 1 10 0 9 15 1 11 3 0 2 13 9 2
18 11 13 15 9 15 0 1 10 9 2 3 15 15 3 3 13 13 2
32 8 15 0 9 1 4 4 2 13 15 10 9 1 10 9 7 13 11 3 10 9 1 0 9 3 3 1 0 9 1 4 2
20 0 9 1 10 0 0 9 4 11 2 15 0 3 10 9 1 11 9 13 2
21 10 9 1 10 9 2 15 0 9 3 4 4 2 13 11 0 9 0 4 4 2
18 1 10 9 1 10 9 9 4 3 3 1 10 9 10 0 9 4 2
9 1 10 0 11 13 10 0 11 2
12 10 9 13 15 9 1 11 1 12 1 13 2
11 10 9 4 12 2 12 2 12 7 12 2
11 15 0 9 13 3 3 1 10 9 4 2
15 11 13 1 10 9 10 0 11 1 12 9 2 12 2 2
20 10 0 9 13 15 3 4 1 10 9 1 8 7 8 2 15 13 1 11 2
35 1 10 8 12 9 13 9 13 12 9 1 10 9 1 11 1 11 9 4 1 8 12 9 1 9 7 9 1 4 1 10 9 1 11 2
16 15 13 12 9 1 10 9 7 13 1 10 0 9 1 3 2
22 10 9 13 1 12 9 7 1 10 9 1 10 1 3 0 13 1 10 9 13 9 2
45 1 15 9 13 9 8 3 16 15 0 9 1 10 9 2 9 7 15 0 1 10 9 4 4 16 10 13 0 3 1 9 12 7 15 9 1 9 1 9 7 9 4 4 4 2
25 2 15 13 15 15 9 1 4 2 16 3 1 13 1 10 9 1 10 13 0 2 2 3 11 2
22 16 9 13 15 10 9 1 10 1 10 9 9 13 9 16 1 10 15 9 1 4 2
16 10 9 4 3 2 8 1 2 1 10 9 1 10 9 4 2
21 16 15 0 13 4 10 9 1 10 9 1 10 9 1 4 13 15 10 11 3 2
12 10 9 1 11 4 3 0 2 3 13 4 2
11 10 3 13 9 13 15 8 1 10 9 2
20 10 9 13 3 1 10 9 2 16 10 9 1 10 3 13 9 3 1 13 2
15 10 9 1 10 11 13 15 3 7 13 1 10 9 8 2
20 11 13 10 12 9 4 1 10 0 9 1 11 15 15 1 11 13 0 4 2
20 3 10 15 9 4 3 1 9 2 13 1 9 8 2 1 10 9 8 4 2
34 8 10 0 9 2 15 13 1 15 9 1 11 2 13 0 10 0 9 9 7 9 10 9 7 9 3 16 3 10 9 3 1 13 2
11 3 4 1 10 9 15 13 9 1 9 2
9 15 13 15 10 9 8 1 8 2
31 1 10 0 9 1 10 9 13 10 0 9 16 15 9 8 1 15 0 9 1 10 0 9 4 16 3 10 9 1 13 2
17 0 4 15 3 0 2 7 10 9 1 12 4 3 3 0 15 2
27 10 9 13 15 3 3 15 15 1 0 9 4 2 16 15 3 3 0 0 9 3 1 0 9 0 4 2
24 15 13 2 16 15 15 3 3 13 2 16 15 1 10 9 4 4 16 15 10 9 13 4 2
6 0 13 15 1 11 2
9 11 13 1 10 9 8 3 0 2
11 3 13 11 15 3 3 1 15 9 3 2
12 15 13 3 1 15 9 10 3 0 9 4 2
7 15 4 3 10 3 0 2
6 11 13 3 15 3 2
25 2 12 9 3 10 9 1 10 9 1 10 0 1 11 2 13 10 0 9 10 9 1 10 9 2
25 1 10 9 7 10 0 9 1 8 4 10 9 4 1 10 0 9 1 11 2 10 0 1 8 2
13 15 4 4 1 10 9 2 9 2 11 2 2 2
19 1 15 0 9 8 13 1 10 0 3 13 9 12 9 1 10 9 4 2
16 10 9 13 4 4 16 10 9 2 15 4 3 3 10 9 2
10 10 9 4 12 9 13 1 10 11 2
15 10 9 4 16 9 1 10 9 4 2 3 16 2 8 2
12 11 13 15 9 10 9 1 12 9 1 4 2
7 15 4 4 1 10 9 2
16 10 9 13 3 0 2 7 13 2 16 4 4 2 0 4 2
14 1 12 13 11 12 9 1 10 0 9 1 9 9 2
23 10 9 1 10 9 4 3 1 12 9 1 9 4 7 10 9 1 15 9 4 3 4 2
38 15 9 2 1 10 9 3 10 9 1 15 9 13 4 2 13 3 3 2 16 10 13 9 1 9 4 4 7 16 10 9 0 1 12 9 4 4 2
13 15 0 9 13 1 9 8 7 13 3 4 4 2
24 15 13 3 1 15 13 13 2 15 4 4 1 10 0 9 2 8 2 2 10 0 9 9 2
21 1 15 0 9 2 7 1 10 13 9 2 13 10 0 11 11 15 3 0 4 2
29 10 0 9 1 10 9 1 11 7 11 2 8 2 13 10 9 3 1 10 9 1 10 9 1 10 0 9 11 2
37 1 10 9 1 10 0 9 2 15 9 3 2 4 15 3 3 4 2 16 10 9 1 10 0 7 0 9 1 10 0 9 1 10 9 4 4 2
12 15 1 15 4 0 13 10 15 4 8 4 2
7 15 9 4 12 9 0 2
10 15 4 9 7 3 2 15 4 9 2
23 9 4 8 15 1 9 1 10 9 13 1 12 9 1 12 9 1 10 9 3 1 11 2
27 16 10 9 13 2 16 10 0 9 3 9 3 4 2 3 13 15 4 2 16 15 0 0 9 0 4 2
3 2 2 2
30 10 9 1 9 1 10 9 13 3 1 10 0 9 2 15 1 10 11 2 15 15 13 4 4 16 13 0 9 2 2
9 1 9 13 15 3 3 0 9 2
11 10 9 13 15 3 0 1 10 9 4 2
22 10 0 9 3 2 13 3 1 13 9 7 3 1 9 15 15 0 7 3 13 13 2
22 10 9 1 10 0 9 4 8 2 16 15 0 4 13 4 1 10 9 1 10 9 2
11 15 13 10 0 9 8 2 3 10 9 2
25 10 11 13 3 16 15 9 4 4 4 1 10 9 1 10 9 1 9 7 9 1 10 0 9 2
6 3 13 15 3 4 2
24 10 9 1 10 13 9 13 15 8 1 15 8 4 4 2 16 3 10 9 1 8 4 4 2
16 10 0 0 9 1 15 9 13 10 9 1 11 0 4 4 2
12 10 9 2 8 10 0 11 2 4 3 4 2
9 7 3 15 13 1 11 4 4 2
13 8 13 11 3 15 9 3 1 4 7 15 9 2
20 10 9 2 16 10 9 1 10 9 1 10 11 15 15 9 4 4 3 0 2
23 1 15 15 3 13 4 2 13 10 9 7 9 0 4 2 16 10 9 3 0 13 4 2
17 10 9 13 10 0 9 1 10 0 0 9 0 9 1 4 4 2
12 10 9 1 9 13 15 9 3 3 0 4 2
16 11 2 11 2 11 7 11 13 10 15 0 9 16 0 9 2
13 3 13 15 10 9 1 9 3 3 3 0 4 2
16 10 9 13 10 9 1 9 4 2 15 1 10 9 9 13 2
26 0 13 15 0 4 2 1 10 9 1 10 9 15 1 1 10 9 3 1 13 2 15 16 9 13 2
10 15 9 13 10 9 1 10 9 4 2
14 10 9 4 3 10 0 9 7 13 1 10 9 9 2
33 15 13 15 0 8 10 0 9 15 10 9 8 2 15 15 0 13 1 10 9 1 9 1 10 9 7 10 9 2 8 13 4 2
31 2 3 13 9 2 2 3 13 15 2 2 3 0 16 10 9 15 3 4 4 2 13 15 3 9 4 8 1 4 2 2
23 10 9 13 15 3 2 13 3 1 10 9 7 13 15 16 3 15 3 15 1 13 4 2
7 7 15 4 10 9 8 2
6 15 13 10 9 3 2
29 15 13 1 15 9 3 15 9 16 10 9 15 9 1 15 0 9 13 1 10 9 1 9 7 9 1 10 9 2
22 2 15 13 15 3 2 2 13 15 10 13 9 1 10 9 1 10 9 1 10 9 2
16 7 15 16 15 15 9 13 3 13 3 1 4 1 11 2 2
19 10 9 16 10 9 15 3 1 9 4 4 2 13 11 0 1 10 9 2
22 2 16 15 10 9 13 4 3 1 9 1 15 9 1 4 2 13 15 15 0 4 2
28 15 4 15 9 12 9 1 10 11 4 2 15 4 1 9 0 1 10 9 1 10 9 1 10 9 1 9 2
11 1 0 9 4 8 8 10 0 9 4 2
21 15 8 13 1 10 13 9 10 0 9 1 9 1 10 0 0 9 7 10 9 2
35 3 13 15 8 10 9 9 1 10 9 0 3 1 13 1 15 13 1 13 9 7 15 13 1 9 7 9 1 9 1 10 0 0 9 2
27 16 15 9 1 0 9 10 0 13 9 13 4 2 4 10 9 1 10 9 1 10 0 9 10 13 9 2
24 1 10 9 8 4 10 11 10 9 1 10 9 1 10 0 7 0 9 1 10 9 8 4 2
6 3 3 3 1 11 2
34 2 10 9 1 15 9 15 10 0 9 13 7 15 9 13 16 1 13 16 10 11 3 0 7 0 4 7 11 3 0 7 0 2 2
32 3 13 10 9 8 3 10 9 1 11 7 11 16 15 10 9 13 4 4 1 2 10 0 0 9 3 10 9 9 13 2 2
19 1 11 13 10 9 15 1 12 1 10 9 4 4 2 3 3 4 4 2
34 16 10 9 1 0 9 10 9 1 10 0 9 1 15 8 13 4 2 13 10 9 1 10 0 9 11 16 3 1 9 4 4 4 2
16 10 15 9 1 10 11 4 1 12 9 1 7 12 3 4 2
24 9 3 13 10 9 1 10 9 7 9 1 10 9 9 4 1 10 9 2 3 15 9 13 2
24 10 9 13 3 0 1 10 9 4 4 2 16 3 3 10 9 1 15 0 9 13 4 4 2
22 3 4 15 9 3 11 16 9 4 2 3 10 9 15 3 1 15 9 13 4 4 2
28 1 10 9 2 8 10 9 13 15 10 0 9 2 1 10 9 7 9 1 10 9 13 10 9 15 0 4 2
13 13 9 13 3 3 1 9 1 10 9 1 4 2
29 10 3 13 11 15 15 1 10 9 1 10 9 1 10 9 1 9 13 1 4 2 13 1 9 1 15 9 9 2
39 1 10 9 13 15 1 10 9 7 10 9 10 9 3 0 8 1 13 2 16 10 9 2 15 15 3 3 0 13 13 4 2 1 10 9 13 4 4 2
18 9 4 15 0 8 1 11 1 10 9 1 10 11 1 11 8 4 2
21 10 9 2 3 10 9 13 2 4 1 10 15 9 2 15 15 9 13 2 4 2
16 8 4 1 10 9 4 2 16 10 9 1 10 9 4 4 2
5 15 4 8 0 2
23 15 9 7 9 13 0 13 1 10 9 1 11 4 4 2 16 12 0 1 10 15 9 2
30 10 11 13 0 4 3 1 0 10 9 1 9 4 4 4 7 3 10 9 1 10 9 1 9 7 0 4 4 4 2
19 15 13 15 3 16 15 3 12 4 4 4 2 16 15 9 4 4 2 2
10 9 8 13 3 3 3 1 10 9 2
27 1 0 9 1 15 13 8 4 2 16 11 7 3 11 2 15 1 12 7 12 13 2 3 10 9 4 2
9 15 13 3 15 9 15 9 4 2
9 15 2 16 10 9 3 3 13 2
10 3 0 13 12 3 3 1 10 9 2
12 1 10 0 9 13 3 0 9 1 9 8 2
14 10 9 4 8 4 1 9 1 8 2 4 12 2 2
28 10 9 13 1 10 0 8 2 12 9 2 0 9 3 1 15 4 4 2 16 4 4 1 10 9 1 8 2
15 0 13 10 0 9 1 8 2 3 12 9 15 4 4 2
15 16 11 0 1 10 9 13 2 13 15 9 1 12 9 2
14 10 9 13 3 3 4 2 13 15 7 13 3 3 2
36 3 1 10 9 13 15 2 7 1 10 9 3 2 15 10 0 9 1 10 9 4 13 2 13 15 3 15 15 9 4 1 10 15 0 9 2
8 10 9 13 15 3 0 4 2
11 11 13 8 9 15 1 10 9 13 4 2
8 15 4 3 13 1 10 9 2
21 15 4 10 9 8 7 10 9 4 3 3 4 1 3 10 9 1 10 9 3 2
30 9 11 13 3 4 2 16 15 12 9 15 8 8 13 2 3 15 3 4 2 16 15 1 11 3 1 10 9 4 2
27 15 13 3 15 3 2 7 15 4 15 1 15 9 9 4 4 2 15 1 10 9 0 3 13 4 4 2
18 3 1 15 9 1 10 0 9 2 8 2 3 0 2 13 15 9 2
16 13 15 9 2 16 15 3 13 8 2 16 15 9 3 13 2
6 3 4 15 9 4 2
9 15 13 15 4 2 16 15 0 2
6 15 4 13 1 4 2
20 15 13 15 9 1 11 3 3 4 4 2 7 15 9 4 3 13 7 13 2
14 7 3 3 13 15 1 10 0 2 15 10 0 13 2
9 7 15 1 15 13 15 9 4 2
8 15 1 10 9 13 15 9 2
32 16 11 10 9 4 2 13 15 15 0 9 2 15 11 13 1 0 9 2 9 7 9 2 16 10 9 15 13 4 1 11 2
39 10 1 11 13 9 4 3 3 3 0 2 7 15 1 10 0 9 1 11 4 10 0 9 1 9 1 9 7 9 7 9 2 3 9 7 9 1 9 2
15 3 13 10 9 10 9 4 16 10 0 9 1 10 9 2
32 15 13 3 0 9 4 2 15 0 4 4 1 10 9 2 10 0 9 15 9 2 9 2 9 7 15 9 13 1 15 9 2
17 1 12 0 13 11 15 9 1 10 9 1 9 1 10 0 9 2
22 3 13 3 10 15 9 9 13 1 0 7 0 9 2 15 0 0 13 1 10 9 2
29 15 13 15 1 10 9 5 10 9 5 15 1 10 9 1 15 8 13 2 7 3 3 4 4 1 10 0 9 2
16 10 0 9 11 1 8 13 15 16 9 7 15 9 1 13 2
26 8 12 13 10 0 9 2 8 2 9 2 15 0 9 2 7 10 9 9 15 15 8 1 4 13 2
44 1 12 9 13 3 15 9 7 9 10 2 0 9 1 10 9 2 10 15 0 9 1 10 0 15 9 2 15 12 9 13 4 8 10 9 1 10 3 13 9 2 8 2 2
14 8 13 15 4 16 3 1 10 9 0 9 4 4 2
9 2 15 13 1 10 9 0 4 2
12 7 1 0 9 2 13 15 3 3 3 4 2
13 10 9 13 3 10 0 9 4 1 10 0 9 2
5 15 13 3 9 2
21 3 13 15 16 10 0 9 2 15 1 10 9 1 10 9 13 2 3 1 13 2
16 3 13 15 3 16 3 1 15 9 10 9 1 4 4 2 2
30 15 9 1 10 9 8 2 2 10 9 1 9 1 8 8 10 9 1 10 0 9 1 10 0 9 2 13 16 9 2
9 0 8 11 8 1 8 7 8 2
29 1 10 0 9 1 8 2 3 10 9 7 15 8 1 15 1 15 9 9 13 1 3 11 2 11 0 11 2 2
10 11 2 11 2 11 2 11 2 11 2
17 10 9 1 9 1 9 1 10 0 7 1 10 0 9 15 9 2
8 8 9 13 10 9 3 4 2
6 11 13 15 15 0 2
44 3 16 3 0 8 2 12 9 3 2 2 10 0 11 2 15 1 10 0 9 1 10 9 7 15 2 8 2 13 4 2 0 8 10 9 2 15 3 10 0 9 3 13 2
11 10 9 1 15 8 13 10 9 3 4 2
31 11 13 16 15 9 3 9 4 7 3 15 9 13 15 15 13 8 0 3 16 10 0 9 10 9 1 10 9 1 13 2
17 3 0 13 11 3 1 11 1 8 3 15 9 1 11 7 11 2
8 15 13 9 13 3 15 4 2
19 15 4 3 0 1 10 9 1 13 16 10 0 9 3 1 11 4 4 2
11 10 9 1 10 0 9 13 3 15 9 2
19 1 10 9 1 8 13 10 0 9 8 3 1 10 9 7 15 9 4 2
8 3 13 15 1 10 0 9 2
16 15 4 10 9 1 11 1 15 9 3 10 9 3 1 13 2
10 2 8 2 4 10 0 0 9 4 2
11 16 15 1 10 9 1 9 8 1 13 2
16 2 10 9 1 15 9 7 3 13 15 0 9 3 3 2 2
26 3 4 3 3 15 15 3 3 1 9 13 2 15 13 10 0 9 4 15 10 9 3 15 13 13 2
26 3 1 10 0 9 1 10 0 9 13 12 9 7 9 3 1 15 9 7 9 7 9 3 3 4 2
25 15 4 10 9 1 9 8 7 9 8 10 9 1 10 0 11 1 15 0 2 0 9 1 13 2
38 8 2 0 0 0 9 1 1 10 9 13 1 9 8 1 10 0 9 3 1 10 9 5 10 9 1 0 9 5 15 1 15 0 9 9 13 4 2
8 10 9 1 15 4 0 8 2
30 1 10 9 13 8 9 1 15 8 1 10 9 1 10 1 10 9 15 9 1 11 13 4 2 11 1 10 15 9 2
26 1 10 13 9 2 10 0 1 10 11 1 15 9 2 13 15 10 9 4 1 10 9 1 9 11 2
11 1 10 9 4 3 3 12 0 9 4 2
29 1 10 11 8 2 10 9 1 10 0 9 2 0 16 15 0 8 4 2 7 1 10 11 10 9 8 1 11 2
21 13 4 3 3 3 2 16 2 1 10 9 3 2 1 15 9 0 10 9 4 2
47 3 13 15 12 9 1 10 11 7 15 13 10 9 1 15 15 9 7 10 0 9 1 15 9 2 15 3 1 13 9 1 10 9 4 4 7 3 13 15 15 3 4 15 15 4 4 2
18 10 9 13 2 16 3 3 4 4 2 1 0 9 2 13 1 12 0
9 11 13 1 12 10 0 9 3 2
32 1 10 0 9 13 15 9 16 15 10 9 1 10 0 9 13 4 2 10 0 9 3 15 3 3 3 1 10 9 13 4 2
18 15 16 1 10 9 3 2 3 9 13 10 9 1 15 1 1 4 2
13 3 13 1 15 9 3 15 3 15 8 4 4 2
30 10 9 4 1 10 0 9 4 5 9 2 0 9 7 0 9 1 10 9 5 15 15 3 13 7 3 0 9 13 2
22 10 9 4 3 13 2 16 10 9 1 10 9 1 10 9 15 3 0 7 0 4 2
12 15 13 1 10 13 9 7 13 10 9 3 2
32 1 11 2 3 1 10 9 1 11 9 10 9 4 4 2 13 16 10 0 0 9 3 3 10 0 9 15 9 1 10 9 2
35 15 3 0 8 15 10 0 9 1 15 9 1 15 9 13 2 13 15 3 1 10 9 1 15 9 1 10 1 3 1 13 9 1 8 2
23 9 3 8 2 9 8 2 9 8 2 8 7 0 9 1 11 8 1 10 0 9 13 2
14 15 12 0 15 11 1 3 13 4 4 0 8 4 2
11 1 10 9 2 10 9 1 9 7 8 2
28 3 10 9 1 10 9 15 10 9 8 13 16 1 11 2 1 11 11 7 11 1 10 11 1 8 1 4 2
23 9 2 15 15 8 13 7 13 2 10 9 1 10 0 9 1 9 2 13 0 4 4 2
11 15 13 3 0 4 0 10 9 1 13 2
13 1 10 0 9 13 10 12 9 0 9 1 9 2
15 11 13 3 3 15 1 9 2 15 4 3 10 0 9 2
31 1 15 8 1 12 1 11 13 15 12 0 9 7 1 15 8 1 12 1 11 13 15 3 1 9 11 3 3 12 3 2
24 1 10 9 4 11 9 1 10 9 1 4 1 10 9 11 7 8 1 10 9 2 8 2 2
14 10 13 9 4 3 1 10 0 9 15 9 9 4 2
20 12 9 2 15 9 1 10 9 11 8 13 15 8 3 4 1 10 0 9 2
9 1 15 4 3 12 9 0 13 2
21 15 15 16 10 9 1 10 9 15 9 1 10 9 13 4 3 15 9 13 4 2
16 16 15 3 13 16 15 3 4 2 13 15 15 1 15 13 2
17 10 9 1 15 12 13 2 15 1 10 9 4 4 4 3 0 2
9 3 13 9 7 9 7 15 9 2
5 16 9 1 13 2
16 15 13 3 2 16 10 0 9 1 10 9 1 10 9 4 2
40 10 0 9 3 2 7 10 0 9 1 10 9 2 3 9 10 0 9 1 15 9 13 7 10 13 9 13 2 13 3 1 10 9 7 1 10 9 15 2 2
22 1 15 13 9 2 12 9 5 9 12 1 8 2 13 8 10 9 1 13 13 9 2
15 8 16 0 1 13 2 16 10 0 15 9 1 9 13 2
27 1 10 9 1 10 0 0 9 13 10 0 9 9 16 15 8 2 8 2 8 2 8 2 8 7 8 2
25 8 8 2 13 2 3 12 0 9 11 3 16 10 11 3 2 16 15 10 9 1 15 8 13 2
29 10 9 1 10 0 0 9 2 1 10 0 2 9 7 9 4 3 4 2 16 3 1 0 9 3 13 9 13 2
31 15 13 3 1 15 9 11 3 2 7 15 13 3 16 15 1 10 0 9 1 11 1 10 9 1 15 0 13 4 2 2
32 1 15 0 9 16 9 1 10 11 2 10 9 1 10 0 7 0 9 1 15 0 8 13 11 10 9 1 10 0 9 4 2
29 3 13 15 3 2 16 10 0 0 9 1 10 0 9 15 4 1 10 0 0 9 1 10 9 1 10 0 9 2
28 0 4 15 4 2 0 2 15 4 0 2 7 15 9 4 9 2 3 15 1 10 9 10 0 9 13 2 2
11 1 9 13 3 1 10 9 12 9 4 2
13 1 15 8 4 15 1 10 0 9 4 7 4 2
12 1 10 9 13 15 16 9 1 10 0 9 2
12 1 10 9 13 3 3 3 15 16 15 9 2
8 2 15 13 3 3 4 2 2
27 8 13 15 15 9 2 16 15 15 13 7 13 1 10 9 1 11 1 10 9 1 10 0 9 9 13 2
17 10 9 4 1 10 9 1 10 0 9 9 1 10 9 8 4 2
7 2 15 4 0 3 0 2
4 11 4 13 2
8 2 15 4 3 15 9 2 2
6 15 13 12 9 3 2
9 2 15 4 0 0 1 15 9 2
10 15 13 1 3 1 3 1 10 9 2
24 3 0 13 10 9 1 10 0 9 2 15 3 10 9 13 4 1 10 9 1 10 0 9 2
25 10 9 1 10 11 4 1 10 9 1 9 1 12 4 7 10 9 4 0 2 0 7 0 9 2
23 10 9 5 10 0 9 1 10 9 5 13 11 1 12 2 7 15 12 9 9 13 15 2
22 10 9 13 3 12 9 10 9 7 4 1 10 9 8 3 3 0 1 10 13 9 2
9 3 4 10 9 0 1 9 4 2
12 15 13 15 3 9 2 2 4 15 0 9 2
7 10 9 4 3 1 11 2
14 15 4 3 3 0 15 3 3 1 10 11 13 4 2
9 16 3 13 13 4 15 0 4 2
12 7 15 4 3 0 16 10 11 1 11 13 2
16 1 15 9 13 9 1 10 9 1 15 12 7 12 9 4 2
12 9 11 1 11 13 10 0 9 4 1 12 2
8 10 9 9 10 9 1 8 2
7 3 12 13 3 0 4 2
18 15 13 1 10 9 15 0 4 16 10 9 1 10 9 3 1 4 2
9 10 9 4 1 10 9 3 0 2
34 7 10 0 9 1 11 13 15 3 4 16 15 15 8 4 4 2 16 15 0 9 3 1 13 7 10 15 9 1 15 1 13 2 2
14 10 9 4 1 9 12 1 15 9 0 1 9 4 2
8 4 4 10 9 3 1 4 2
20 10 11 13 1 10 13 9 10 9 1 10 9 1 10 9 1 10 0 9 2
38 1 10 9 15 10 9 13 7 1 10 9 1 0 9 13 10 9 3 2 16 10 11 13 1 12 1 12 9 2 7 1 12 1 12 9 15 4 2
32 10 9 13 15 2 0 9 2 1 10 9 1 10 9 1 10 9 2 15 0 4 10 0 9 1 10 9 12 3 1 4 2
40 1 10 0 9 1 15 8 1 11 2 15 1 10 9 1 9 1 11 1 15 1 10 0 12 9 4 4 2 13 15 1 9 1 9 1 9 7 9 3 2
9 10 9 1 10 0 9 11 13 2
27 2 10 9 13 1 3 0 9 10 15 9 1 11 4 16 15 15 3 0 16 9 1 15 9 13 2 2
21 9 7 9 13 10 0 9 1 10 12 1 12 9 15 10 9 0 1 4 13 2
36 1 10 0 9 1 10 9 1 11 7 11 2 13 1 10 0 9 2 15 9 10 0 9 8 1 11 7 10 0 9 8 1 8 8 4 2
17 1 15 0 15 2 0 2 9 13 13 9 11 3 1 11 3 2
20 10 9 1 9 11 7 15 0 9 11 4 0 13 1 10 9 1 11 4 2
7 15 9 4 3 3 0 2
15 10 15 13 15 9 2 3 1 11 4 1 10 0 9 2
14 11 13 3 2 15 3 10 0 2 0 9 8 4 2
37 15 0 9 13 10 9 1 11 4 4 2 15 1 10 9 13 16 10 0 9 2 15 10 0 9 1 10 9 13 1 10 0 9 1 10 9 2
18 2 15 4 15 0 16 9 2 2 13 11 16 15 15 13 9 13 2
21 10 9 13 15 1 15 9 3 1 10 9 3 1 10 0 9 0 9 4 4 2
13 3 10 9 1 10 9 1 0 9 4 0 4 2
8 0 13 15 9 1 15 9 2
31 1 10 9 1 10 9 1 10 0 9 13 15 12 0 9 8 4 2 15 1 15 9 0 12 7 12 9 0 13 4 2
16 3 13 15 7 15 9 12 9 9 4 2 15 9 12 9 2
20 3 4 15 10 9 1 15 8 7 15 8 2 1 15 9 15 15 9 13 2
16 0 4 11 9 1 15 8 7 9 1 15 9 1 15 9 2
19 10 10 9 13 8 3 16 9 1 15 9 1 15 8 2 10 0 11 2
19 15 4 9 1 10 0 9 9 2 1 10 9 11 7 9 1 10 9 2
8 7 15 13 15 3 3 4 2
16 15 13 15 3 4 16 15 9 4 7 15 3 0 9 4 2
24 3 1 9 13 15 0 9 3 2 7 0 13 15 13 15 3 3 0 4 16 3 1 11 2
11 0 2 15 13 3 3 3 1 15 9 2
10 7 15 13 15 3 3 3 15 4 2
11 3 13 15 15 9 7 15 13 0 4 2
43 3 4 10 9 2 15 13 1 10 15 9 15 1 11 4 4 1 10 11 1 11 4 2 7 9 11 2 1 10 9 1 9 2 13 1 10 9 7 13 15 0 9 2
25 10 9 1 10 0 9 1 12 9 13 3 15 9 1 0 9 16 11 2 11 2 11 7 11 2
20 10 0 9 13 11 2 10 0 9 1 10 9 1 8 2 0 1 15 9 2
32 11 2 10 9 1 10 13 9 1 10 0 9 2 13 1 9 4 2 1 0 9 13 15 1 10 13 9 1 11 3 3 2
19 1 10 9 1 3 12 9 13 11 1 12 9 1 13 4 1 10 9 2
20 15 4 8 1 12 2 16 15 0 8 3 1 10 11 1 10 11 4 4 2
16 3 13 15 1 10 1 10 9 13 9 1 11 15 9 3 2
12 3 12 1 10 12 13 9 9 10 9 3 2
21 1 10 9 1 10 11 1 11 13 3 10 11 1 10 9 1 11 15 9 4 2
5 15 13 1 11 2
10 11 13 8 1 8 1 10 0 9 2
14 10 2 8 2 11 2 15 10 0 9 1 11 13 2
33 10 9 1 11 7 10 0 9 1 10 9 1 10 9 2 8 8 2 13 3 10 9 2 15 10 9 13 1 15 15 0 9 2
20 8 4 11 1 10 9 1 15 3 10 9 0 7 3 13 9 8 16 0 2
24 1 10 0 9 13 8 3 10 9 1 12 9 2 13 1 8 1 12 7 8 1 12 9 2
41 10 9 13 3 1 10 9 4 16 10 9 1 8 2 9 1 10 9 11 1 10 9 3 4 1 0 9 2 3 1 0 9 7 3 1 10 0 9 1 9 2
15 8 13 16 15 8 4 16 10 9 4 4 1 10 9 2
35 1 9 1 10 9 9 1 9 13 15 12 9 3 13 9 1 3 4 7 15 4 8 9 1 9 7 9 3 3 0 2 3 13 8 2
22 15 0 8 2 10 0 0 9 2 15 0 10 13 9 13 2 4 11 0 0 4 2
44 10 9 4 10 0 9 1 10 9 4 1 9 1 9 1 10 11 2 8 2 1 10 0 7 0 9 1 10 9 10 11 2 15 15 9 13 1 0 9 1 9 7 9 2
26 16 1 10 9 1 10 9 3 1 13 13 10 9 9 8 4 2 3 4 13 4 1 9 7 9 2
20 3 13 3 10 9 0 2 15 3 4 13 7 1 10 9 1 10 11 13 2
15 7 3 13 3 3 15 15 10 9 1 10 11 13 2 2
10 3 4 3 10 9 1 12 9 8 2
20 2 6 2 1 10 9 2 10 9 2 13 3 0 15 9 1 10 11 13 2
18 1 15 13 1 10 9 1 10 0 9 13 15 10 9 1 9 2 2
43 1 10 0 9 3 1 10 9 8 2 9 1 15 8 2 13 15 4 2 16 11 4 4 10 0 9 1 4 4 1 15 13 2 9 2 9 2 9 2 9 7 9 2
31 1 10 9 1 10 9 7 10 9 1 8 2 4 5 8 1 10 9 5 15 0 2 8 3 13 9 2 8 2 4 2
24 10 13 9 2 8 2 2 13 1 12 9 2 4 3 0 16 1 10 0 11 1 4 4 2
14 15 13 15 15 13 2 4 1 10 9 1 13 9 2
12 7 2 9 1 10 9 2 15 13 3 15 2
14 10 9 13 2 15 13 1 3 2 16 3 1 3 2
23 15 13 15 9 2 13 15 3 2 13 1 10 9 1 15 12 9 7 13 10 0 9 2
23 1 15 9 13 16 10 9 9 2 15 16 12 9 2 16 15 1 13 2 4 15 4 2
6 15 13 10 0 9 2
24 1 0 9 1 10 9 4 10 9 1 11 9 1 0 9 0 4 1 10 9 1 15 8 2
13 3 13 15 8 1 10 9 11 3 10 9 3 2
14 10 0 9 13 15 4 1 9 15 9 13 1 9 2
10 15 13 15 8 10 9 8 10 9 2
23 15 13 3 3 1 15 0 9 1 4 2 7 3 0 9 13 0 9 7 9 0 4 2
28 1 10 0 9 8 1 8 13 15 15 9 3 3 4 7 15 13 3 3 3 4 1 10 9 1 10 9 2
22 10 9 3 4 3 16 10 9 2 3 11 10 9 9 13 4 2 0 7 0 4 2
17 15 13 1 10 9 2 15 1 11 10 9 13 2 2 8 2 2
26 15 13 3 10 3 1 10 0 9 13 0 9 11 2 8 2 2 15 15 1 10 9 13 13 4 2
52 10 9 13 1 15 9 3 9 1 4 1 10 9 2 16 15 13 10 15 13 9 16 10 0 9 4 4 2 16 15 15 3 0 0 1 15 13 12 2 7 13 16 15 10 9 4 2 15 15 3 13 2
10 2 15 4 15 0 9 7 10 9 2
16 10 9 13 10 9 1 10 9 1 10 9 1 13 1 9 2
20 15 0 8 13 5 15 13 1 0 0 9 5 13 1 15 9 0 1 9 2
7 10 9 13 10 9 8 2
20 2 15 13 15 4 16 15 3 3 3 0 4 1 15 9 1 9 7 9 2
22 16 1 15 9 10 9 13 4 2 4 10 9 16 15 3 3 1 4 3 0 0 2
19 7 15 9 1 8 4 3 9 3 4 7 13 3 0 0 0 8 2 2
6 15 4 3 10 9 2
26 11 9 8 2 0 7 16 15 0 9 13 1 10 0 0 9 2 13 1 10 9 1 11 15 9 2
26 0 13 15 0 4 16 3 15 1 10 12 9 2 15 1 10 0 9 1 8 4 4 2 4 4 2
12 10 9 8 13 3 4 16 9 1 4 4 2
32 15 4 10 0 0 7 0 9 1 15 13 9 1 10 9 7 10 9 2 15 3 1 11 13 4 2 2 3 10 0 9 2
18 2 4 15 15 15 2 3 13 15 15 10 9 1 10 9 11 4 2
16 7 3 13 15 3 10 9 4 2 7 15 13 10 9 2 2
37 1 10 9 1 10 0 9 4 1 0 9 10 9 1 9 4 2 15 4 4 1 10 9 1 10 11 7 1 10 13 12 9 2 15 0 9 2
31 10 9 13 15 0 16 15 1 10 9 4 4 7 3 2 10 0 9 2 4 4 1 10 9 1 10 9 7 10 9 2
26 2 15 4 1 15 0 2 2 3 10 9 2 2 16 0 9 1 15 8 3 16 9 4 4 2 2
24 9 2 15 11 1 10 9 1 9 9 13 1 10 9 1 15 13 2 13 15 9 3 4 2
17 15 13 3 15 0 13 8 10 9 1 10 9 16 10 9 4 2
13 10 9 4 10 9 0 1 9 1 12 9 4 2
39 10 9 13 10 9 0 1 10 9 1 10 9 4 2 13 3 3 2 13 3 3 1 2 13 15 1 10 9 1 10 9 3 7 13 3 1 10 9 2
34 9 1 10 0 9 11 2 15 1 12 8 12 11 1 11 4 4 2 13 15 4 3 0 10 9 1 10 9 1 10 9 4 4 2
17 9 11 13 10 9 1 3 1 10 9 7 13 1 10 9 0 2
27 10 9 11 4 1 10 11 3 0 1 10 0 9 2 15 10 9 9 1 10 9 1 10 11 13 4 2
21 3 1 15 9 13 10 9 11 10 9 1 10 11 4 1 9 2 3 1 9 2
13 15 4 10 9 7 10 9 9 1 10 9 11 2
18 10 12 0 9 13 15 9 15 9 1 10 9 1 12 9 1 15 2
57 1 8 1 4 3 3 3 9 4 1 10 9 1 11 2 10 9 15 1 12 0 4 4 2 12 9 13 7 5 0 10 9 1 10 9 16 15 15 9 4 4 5 10 0 9 1 9 3 0 0 4 2 9 8 12 2 2
15 8 13 3 10 0 9 1 15 9 1 10 9 1 4 2
9 11 13 8 1 0 9 8 4 2
17 10 1 11 3 0 13 9 4 3 1 10 0 0 9 8 4 2
9 10 0 9 13 3 10 0 9 2
8 11 4 3 10 9 0 3 2
2 12 2
2 8 2
8 2 15 13 3 15 1 9 2
16 15 13 3 10 9 2 10 9 2 15 1 10 9 13 4 2
2 8 2
24 9 1 11 3 1 8 2 10 0 1 8 13 9 2 15 3 10 9 13 1 15 0 9 2
17 8 4 1 11 4 16 1 10 3 0 9 1 10 9 1 13 2
7 11 13 0 1 15 9 2
11 0 13 13 15 10 3 0 9 8 3 2
20 11 13 3 2 3 2 12 9 2 12 1 7 12 1 10 9 2 3 0 2
13 15 13 3 3 12 3 0 9 3 1 9 8 2
17 8 13 15 1 15 9 2 15 3 12 9 1 10 9 3 13 2
26 11 2 15 9 1 11 15 13 1 10 9 11 2 13 8 15 9 16 0 9 8 2 11 7 11 2
52 2 10 9 16 11 15 8 4 4 7 0 9 16 8 7 11 4 4 2 4 1 15 10 0 9 16 10 0 9 3 0 4 2 2 3 11 2 15 3 13 4 16 15 11 10 0 7 0 9 4 4 2
18 1 10 9 1 10 0 9 1 10 9 1 11 13 15 0 3 4 2
28 10 0 0 9 8 2 13 15 12 9 3 2 12 9 3 13 1 10 11 1 12 9 9 0 3 0 4 2
19 10 1 9 1 15 8 13 11 13 1 8 2 1 10 0 9 9 4 2
6 11 12 2 8 12 2
19 8 4 3 9 1 10 13 9 1 10 1 9 13 11 3 1 9 4 2
23 10 9 2 15 11 7 11 3 1 10 9 13 2 13 8 8 1 12 9 1 12 9 2
19 9 4 11 1 12 2 11 1 12 2 8 1 12 7 8 1 12 9 2
11 8 13 3 3 3 1 10 9 1 4 2
22 9 11 13 10 9 0 1 11 15 9 1 8 3 1 10 13 9 1 11 4 4 2
14 0 13 13 3 10 9 1 10 9 1 10 0 9 2
39 12 1 10 12 9 13 1 11 13 3 1 10 9 4 2 1 10 0 9 10 0 13 3 10 0 9 9 1 10 15 9 16 10 9 8 9 4 4 2
27 1 8 7 8 13 11 3 3 4 2 16 10 0 9 2 10 15 9 1 9 2 3 0 13 1 4 2
15 12 9 2 15 10 0 9 13 2 13 15 9 0 3 2
13 10 9 8 13 3 3 15 9 1 9 7 9 2
15 10 9 4 4 16 15 9 11 11 11 1 11 4 4 2
29 16 15 4 4 1 9 1 9 8 1 9 11 4 9 4 1 9 15 13 10 0 9 1 10 9 11 1 4 2
66 10 9 8 7 8 13 9 11 2 11 11 7 9 2 7 9 8 2 11 11 2 4 1 10 9 1 10 9 1 10 9 8 11 2 3 10 9 13 16 10 9 1 10 9 9 2 3 0 4 4 4 1 0 9 7 1 9 2 3 9 1 9 4 4 2 2
29 10 12 9 13 1 0 9 3 10 9 4 2 16 10 9 1 15 9 3 3 0 4 4 1 10 9 1 9 2
17 7 16 15 9 0 0 4 7 1 8 9 13 4 2 13 8 2
40 15 4 3 3 10 3 0 9 1 11 2 7 16 15 10 9 0 10 9 13 4 16 11 11 3 13 4 2 13 11 10 9 1 10 0 9 1 10 9 2
9 1 15 9 13 0 9 8 4 2
14 15 4 10 9 2 8 10 13 9 1 10 0 4 2
22 7 15 4 15 0 2 16 15 1 15 9 10 9 2 9 2 10 15 13 9 13 2
22 7 15 13 10 9 2 7 0 9 1 10 3 15 0 2 0 9 4 4 16 0 2
6 8 13 1 10 9 2
27 15 13 0 16 15 0 1 11 3 2 7 3 3 2 15 9 4 1 10 9 7 1 15 10 9 13 2
9 1 15 13 10 9 1 10 9 2
8 1 15 1 9 1 10 9 2
19 15 13 2 3 13 8 2 16 2 9 2 10 9 4 1 2 9 2 2
15 1 10 0 4 10 9 10 9 1 10 9 1 10 9 2
22 13 1 10 9 1 12 9 4 10 9 12 9 0 16 15 8 7 3 12 9 0 2
22 16 10 15 9 1 10 0 11 1 11 10 15 9 4 13 4 2 13 0 3 8 2
40 15 4 10 9 2 15 10 11 2 10 9 1 10 13 9 2 13 7 13 13 2 16 10 0 9 8 10 9 1 10 15 9 10 0 9 1 10 9 13 2
16 10 9 4 3 0 3 0 13 1 10 9 1 10 0 9 2
17 3 1 10 9 1 11 4 11 4 1 10 0 9 1 0 9 2
18 1 15 9 4 10 9 9 0 4 15 10 11 13 4 4 1 9 2
6 15 3 4 10 9 2
9 10 0 9 4 4 1 12 9 2
13 10 11 13 0 9 1 11 15 9 1 15 9 2
23 10 9 1 0 9 7 10 9 15 9 1 11 0 1 4 2 16 10 9 3 4 4 2
12 15 9 13 3 1 4 4 2 16 11 13 2
28 10 0 9 1 15 8 1 10 9 1 15 12 9 1 15 0 8 13 10 9 1 9 15 1 15 9 4 2
36 3 13 8 10 1 10 9 1 8 13 12 9 3 1 4 2 7 1 9 1 8 2 8 7 3 11 4 10 0 9 3 3 0 2 12 2
27 15 13 3 15 9 1 15 3 7 8 13 1 10 0 9 8 7 15 4 3 0 1 10 9 1 3 2
7 0 13 8 1 10 9 2
12 8 13 3 1 11 10 9 4 1 9 8 2
28 10 9 13 10 1 12 9 1 3 12 9 1 8 2 1 11 2 11 7 10 9 1 15 8 1 9 8 2
10 1 15 9 13 10 11 7 10 11 2
40 10 9 13 1 1 15 0 0 9 15 9 1 4 1 0 2 9 7 9 2 15 15 0 3 15 0 1 15 9 13 13 4 4 1 10 9 1 0 9 2
39 16 10 9 1 10 9 8 4 13 10 9 9 1 10 9 10 9 1 10 9 2 15 10 9 13 4 2 1 9 4 7 1 15 9 0 1 8 4 2
29 9 2 13 1 9 1 8 2 13 3 0 4 4 2 16 9 1 10 9 1 10 9 16 15 0 1 13 4 2
21 10 9 1 10 9 1 15 8 2 15 3 15 9 13 2 13 3 0 1 4 2
47 1 9 1 10 9 8 2 11 2 5 0 9 1 10 11 5 13 15 9 8 10 0 9 4 16 3 13 1 10 9 15 10 12 0 9 2 10 11 7 10 11 2 1 10 9 13 2
19 3 13 8 0 10 9 2 7 3 13 8 0 10 9 0 2 12 2 2
8 1 9 11 4 15 9 0 2
15 10 9 1 0 9 13 15 9 1 15 9 3 8 4 2
26 1 10 9 1 9 7 9 1 8 1 10 11 1 11 4 10 9 1 10 11 4 10 9 1 4 2
16 8 7 9 8 13 1 10 0 9 1 15 13 3 1 4 2
19 15 9 13 0 1 15 13 1 9 16 15 9 3 1 9 13 4 4 2
36 2 15 9 13 3 3 15 9 15 4 2 7 16 15 15 9 1 10 9 13 2 13 15 3 13 3 3 2 2 13 15 1 10 9 0 2
14 11 2 9 1 11 7 10 0 9 2 13 12 9 2
35 3 4 3 12 9 1 9 1 10 9 4 2 15 16 3 15 9 1 10 9 1 10 9 5 15 3 4 4 1 10 9 5 1 4 2
9 10 9 4 4 1 10 9 8 2
19 1 10 9 4 10 9 4 1 0 9 2 3 7 3 13 13 1 9 2
10 3 13 3 15 9 3 1 15 8 2
21 3 13 12 9 3 1 10 9 1 10 9 4 4 2 16 11 1 8 4 4 2
4 11 13 3 2
20 3 13 3 3 10 9 4 4 16 15 0 13 4 8 11 10 9 13 4 2
24 7 1 15 9 13 8 15 15 9 4 1 10 9 1 15 9 16 15 10 9 1 11 13 2
10 13 4 2 16 11 15 15 9 13 2
33 7 7 11 12 16 11 12 4 10 9 1 10 9 15 1 10 9 12 3 3 10 0 0 9 1 10 9 1 11 13 4 4 2
34 15 4 0 16 10 0 9 10 0 9 8 10 0 9 1 9 1 11 7 11 10 0 9 13 4 1 10 9 10 9 1 15 8 2
18 1 9 1 10 0 9 1 12 4 10 9 1 11 1 10 9 0 2
16 10 9 11 13 3 3 16 10 9 15 15 3 3 0 4 2
20 0 13 3 3 15 1 10 9 2 10 13 9 13 15 1 15 9 15 0 2
45 2 15 13 15 11 3 0 4 2 2 13 9 8 2 0 9 1 11 2 7 1 10 13 9 11 9 1 10 0 9 2 8 10 1 15 9 1 12 13 9 1 10 9 9 2
17 10 9 11 13 2 16 10 11 1 15 9 1 10 0 9 4 2
16 1 10 9 13 10 9 8 8 16 10 9 3 3 8 4 2
32 8 10 9 1 9 7 10 9 1 10 9 13 15 0 9 1 11 2 16 1 10 9 1 10 9 0 9 4 4 4 4 2
17 3 13 10 1 1 10 9 13 9 16 9 3 9 1 10 9 2
11 15 13 16 10 9 1 9 4 4 4 2
9 15 9 4 3 0 1 10 9 2
47 10 9 1 11 13 16 12 9 2 15 13 1 10 9 2 8 4 1 15 0 9 7 0 1 10 9 9 4 4 1 10 0 9 1 10 9 7 10 11 2 15 1 0 9 4 4 2
27 3 13 10 0 9 2 15 0 3 0 9 9 7 9 1 15 13 2 13 1 9 7 1 9 13 9 2
14 3 13 10 9 13 2 3 15 15 3 0 9 13 2
30 10 0 9 13 15 0 8 2 10 9 13 9 2 3 15 9 1 15 8 4 4 2 0 1 9 15 3 13 4 2
22 2 1 0 9 7 0 9 13 15 10 9 1 10 9 1 10 12 0 9 0 3 2
21 1 11 1 11 2 3 15 9 15 9 13 2 13 11 3 15 1 15 9 4 2
33 3 13 15 8 15 12 9 15 0 1 11 7 9 4 4 1 15 0 9 2 15 10 9 1 0 9 1 15 15 9 13 4 2
17 10 0 9 1 9 4 1 9 4 1 9 1 12 9 1 8 2
26 12 9 13 8 1 10 9 1 11 2 15 15 3 3 3 1 10 9 1 3 12 9 13 0 4 2
19 1 9 13 15 1 10 9 2 1 10 9 7 1 15 0 7 0 9 2
26 10 9 2 15 3 1 10 9 1 9 1 11 4 4 2 13 1 11 1 15 9 11 16 9 4 2
13 8 15 9 13 10 9 1 8 15 15 9 4 2
30 15 4 1 10 9 3 3 15 16 10 9 2 16 10 11 15 9 1 15 9 0 13 4 4 1 9 1 0 9 2
18 2 16 15 15 1 10 9 3 0 4 2 13 15 15 3 0 4 2
6 0 2 16 15 13 2
8 7 2 3 13 10 9 4 2
20 3 12 12 9 4 4 1 0 7 0 9 1 0 9 2 7 1 0 9 2
19 1 11 2 11 7 11 13 15 1 0 9 7 1 9 1 10 0 9 2
32 10 9 1 10 0 9 2 2 11 2 2 13 9 1 10 9 4 16 1 13 2 16 3 2 3 10 0 0 0 9 4 2
23 1 10 9 4 3 0 4 16 10 9 0 1 13 7 10 0 9 1 11 1 13 2 2
23 3 4 1 10 9 9 7 9 10 9 4 1 10 9 1 10 9 1 9 1 10 9 2
28 10 0 9 9 4 8 16 10 9 3 10 9 4 4 2 7 3 15 9 9 13 15 9 3 3 3 4 2
15 3 4 10 9 1 9 10 9 1 4 16 15 1 9 2
23 0 0 9 7 10 13 9 1 10 9 13 15 8 0 10 3 13 7 0 9 1 4 2
17 1 10 9 13 15 10 0 9 8 10 0 0 9 7 0 9 2
22 10 9 8 2 10 9 1 0 9 2 13 3 15 9 16 10 0 9 0 1 13 2
16 16 15 3 3 1 9 13 2 13 15 3 3 15 3 4 2
7 11 13 15 9 16 3 2
13 13 4 10 0 9 3 8 15 2 8 2 13 2
9 8 13 15 9 13 1 4 4 2
17 15 13 1 10 9 1 11 13 10 9 10 0 9 10 0 9 2
19 2 13 15 9 4 2 3 13 10 9 1 11 9 15 0 4 4 2 2
43 15 13 3 3 3 16 10 9 1 10 3 1 11 13 9 2 1 9 1 10 9 3 10 9 2 3 9 7 0 3 3 12 9 13 2 0 2 0 2 4 4 4 2
25 1 0 9 1 10 9 1 10 9 2 15 8 7 10 9 4 9 15 8 2 11 2 8 4 2
40 1 10 0 11 1 10 11 2 1 10 9 3 0 10 9 1 8 13 2 4 1 10 13 7 13 10 0 2 0 9 4 15 15 13 4 16 10 9 3 2
24 11 4 3 10 0 13 9 1 15 15 1 10 9 4 4 2 3 8 1 10 0 4 4 2
20 11 13 3 10 9 1 12 9 4 2 16 11 10 9 1 12 9 13 4 2
4 10 12 9 2
44 11 4 3 0 10 0 9 10 9 3 1 4 7 15 13 3 8 10 9 1 12 9 7 1 15 9 8 3 1 13 2 7 10 9 1 13 1 9 1 9 7 0 9 2
8 3 13 9 2 10 9 8 2
20 10 9 2 11 2 4 0 1 0 9 1 15 9 2 10 11 7 10 11 2
34 10 9 13 11 2 15 9 1 10 11 16 13 1 4 2 2 16 10 9 1 10 12 9 13 1 2 13 1 10 0 0 9 2 2
10 10 9 1 10 11 13 3 10 11 2
30 10 9 1 10 11 13 15 1 15 1 10 12 9 2 15 0 9 11 10 0 9 13 1 15 8 2 15 11 13 2
9 8 3 4 9 2 1 15 3 2
15 15 13 10 9 1 10 11 8 4 2 7 9 11 2 2
10 2 3 13 15 15 9 11 8 4 2
18 15 13 16 0 9 10 0 9 1 15 15 1 10 0 9 4 4 2
13 11 2 11 2 8 7 8 15 0 9 1 11 2
14 15 13 8 1 15 3 15 15 9 3 13 4 4 2
19 3 13 8 11 10 9 2 3 15 1 11 1 8 7 11 1 11 13 2
27 10 9 13 2 15 3 1 15 9 13 1 10 0 9 2 4 1 10 9 15 15 13 4 10 13 9 2
22 15 13 16 9 4 1 11 7 4 13 1 10 9 2 3 3 15 0 9 4 4 2
9 0 4 15 3 1 15 9 4 2
21 10 9 7 9 1 10 9 13 3 1 0 9 0 9 4 1 10 0 0 9 2
26 1 10 0 9 2 3 9 7 9 15 3 0 4 2 4 3 3 1 10 9 15 9 10 9 4 2
19 3 13 3 10 0 9 1 9 2 9 7 9 1 9 2 9 7 9 2
8 10 9 1 10 9 13 0 2
14 10 9 4 15 16 3 1 10 9 1 10 9 4 2
19 15 13 10 0 9 1 10 0 9 9 7 4 1 10 0 9 9 4 2
15 11 13 8 11 0 12 1 10 9 7 9 1 15 8 2
46 10 0 12 9 1 10 9 2 11 2 13 10 0 9 1 12 9 2 15 13 2 16 3 0 12 12 9 1 12 9 7 0 2 1 15 9 4 10 9 4 2 1 15 9 4 2
13 15 9 4 13 1 15 9 1 15 9 0 0 2
9 10 9 4 3 0 2 3 12 2
8 15 13 1 9 1 15 8 2
14 10 9 1 2 11 2 4 1 10 0 9 0 4 2
34 1 15 9 13 11 10 9 2 3 15 4 1 10 9 15 15 8 1 15 13 16 1 4 10 9 1 10 9 7 10 11 1 4 2
24 15 9 4 4 2 16 11 7 11 1 10 12 9 13 1 10 9 1 10 9 1 15 8 2
26 11 7 11 13 15 9 3 1 10 9 2 15 15 3 13 1 10 9 1 10 0 9 1 10 9 2
6 3 13 15 3 15 2
7 10 9 0 9 13 2 2
15 8 4 3 4 1 10 9 1 10 8 9 11 1 11 2
51 11 2 0 2 0 2 13 2 9 1 8 2 0 1 0 9 5 15 13 10 16 12 9 3 5 2 0 9 2 4 0 0 1 10 9 1 9 11 2 15 15 1 10 9 1 11 1 10 9 13 2
14 2 15 13 2 16 15 3 1 9 3 4 4 2 2
4 15 0 13 2
4 8 3 13 2
6 2 10 9 4 0 2
10 8 4 10 3 0 9 1 10 9 2
6 10 9 4 15 13 2
11 12 10 9 7 9 15 9 1 10 9 2
31 12 8 13 1 0 13 1 10 9 10 9 3 1 10 9 2 7 4 1 10 9 1 10 9 8 10 9 1 10 9 2
26 12 16 10 9 10 9 13 13 15 2 0 1 10 9 2 1 15 9 1 15 15 9 4 4 4 2
20 10 0 11 4 0 9 1 11 4 2 3 13 16 10 0 9 1 11 13 2
53 9 7 9 1 10 0 9 13 3 1 10 9 1 10 0 9 3 3 2 16 3 10 9 4 4 2 3 10 12 9 1 9 7 9 2 0 9 2 0 7 0 9 7 10 9 0 7 1 0 9 4 4 2
13 1 15 9 13 3 9 1 10 9 9 4 4 2
13 10 9 13 15 9 4 1 10 9 1 10 9 2
48 10 0 9 1 10 9 2 8 1 10 0 9 2 8 7 8 1 10 0 9 2 2 13 15 3 3 4 2 16 9 1 10 9 1 9 13 2 16 15 8 15 1 7 1 11 4 4 2
10 2 15 13 10 0 9 1 15 9 2
15 7 16 15 3 1 11 13 4 2 13 15 15 8 4 2
12 15 13 3 1 11 0 4 2 2 13 8 2
15 12 13 1 10 9 1 10 0 0 9 16 0 9 4 2
14 3 13 10 0 9 1 11 3 10 9 1 10 9 2
12 15 9 13 16 9 10 9 1 10 11 3 2
33 1 10 0 9 11 4 10 9 2 10 9 11 2 12 2 2 15 9 2 12 2 7 10 9 11 2 12 2 1 0 9 4 2
53 1 10 3 3 13 9 13 10 9 1 10 12 13 9 10 9 3 2 16 15 1 10 9 15 9 9 16 3 2 12 2 4 4 2 3 3 15 2 16 10 0 1 9 13 12 9 3 4 4 1 10 11 2
18 2 15 13 16 15 10 9 4 4 2 15 15 13 7 13 4 2 2
33 2 3 4 15 2 3 3 2 7 3 3 3 2 16 15 10 9 13 16 10 0 9 1 9 10 0 9 1 10 0 9 4 2
24 3 10 9 15 3 13 4 10 0 7 0 9 0 7 1 3 3 0 0 9 8 1 4 2
27 13 15 0 3 4 16 3 1 11 12 9 4 2 16 15 3 15 13 7 13 1 9 1 10 9 2 2
19 11 7 1 10 9 3 11 13 3 0 4 4 1 10 9 1 15 9 2
20 1 9 15 3 0 1 15 1 12 9 4 4 13 3 10 0 9 4 4 2
22 15 13 9 11 2 9 7 9 2 3 1 4 1 10 0 9 1 15 8 1 11 2
22 2 1 10 9 13 15 10 0 9 16 10 15 9 3 1 4 1 10 0 0 9 2
15 13 8 2 10 0 9 1 10 0 9 11 3 1 11 2
25 10 9 15 9 10 9 13 4 13 10 12 9 1 13 9 1 10 9 7 10 9 1 10 9 2
4 11 13 3 2
28 10 9 13 10 9 16 9 1 15 8 1 11 4 2 7 15 13 3 3 4 4 1 15 0 9 1 11 2
32 8 2 15 1 12 9 1 11 4 1 10 9 7 13 1 15 8 1 11 13 1 12 10 0 9 4 1 15 9 1 11 2
6 15 4 10 0 9 2
6 9 4 0 3 0 2
6 15 13 0 10 9 2
15 15 9 13 10 9 1 12 9 1 9 1 15 9 4 2
6 3 13 15 3 4 2
8 1 15 13 15 0 4 2 2
17 8 2 12 9 2 3 12 1 11 7 12 1 10 0 9 3 2
11 3 13 15 3 15 15 9 1 10 9 2
8 0 9 1 11 1 10 9 2
2 11 2
19 2 16 15 15 3 13 3 13 15 0 0 4 4 16 9 1 9 2 2
35 16 15 1 10 9 1 11 3 15 4 1 0 9 2 10 9 3 2 13 16 2 15 3 1 15 10 0 9 4 4 2 2 13 11 2
9 2 15 4 3 10 9 0 3 2
18 15 4 3 3 16 10 11 8 1 15 9 10 3 15 9 13 2 2
2 11 2
8 2 15 13 3 3 0 3 2
8 0 9 1 15 9 13 15 2
6 2 15 4 3 13 2
13 15 9 3 13 10 9 11 10 9 4 3 13 2
8 15 13 10 0 9 0 4 2
23 15 9 4 15 9 3 7 16 15 3 3 15 0 9 13 4 2 13 15 3 4 2 2
32 8 2 12 2 13 1 15 9 10 9 0 1 15 0 9 2 15 3 0 10 9 13 1 10 0 13 9 1 10 0 9 2
22 10 0 0 9 1 8 4 16 15 10 9 9 2 16 15 9 13 4 2 0 13 2
13 1 3 1 13 1 9 15 9 10 15 9 4 2
28 3 4 10 9 4 2 16 15 13 1 9 3 0 9 1 15 13 2 9 15 3 1 15 9 13 4 4 2
20 8 13 15 0 9 8 4 16 15 10 1 9 11 13 9 3 3 13 4 2
27 10 0 9 13 15 4 16 10 9 9 2 0 9 2 15 15 1 9 13 7 15 3 1 10 9 13 2
18 15 13 10 9 1 9 2 3 3 12 1 10 9 1 10 9 13 2
25 15 13 15 1 15 13 1 10 9 1 15 9 2 15 3 13 4 1 0 9 2 10 9 4 2
12 2 16 15 15 9 13 2 13 15 15 2 2
7 10 9 4 0 9 4 2
18 15 13 2 3 2 3 3 15 4 1 4 2 7 11 9 13 3 2
3 1 11 2
17 15 9 13 15 1 10 9 9 4 1 10 9 1 9 1 11 2
24 0 13 10 9 1 10 9 3 15 8 4 7 15 13 9 7 9 15 4 1 10 13 9 2
6 13 4 16 15 3 2
17 3 4 15 0 1 13 16 12 1 10 12 13 9 0 9 4 2
23 10 12 13 9 5 15 1 10 9 8 10 9 1 11 13 4 5 13 15 9 3 4 2
15 8 13 9 7 9 1 15 9 4 1 10 0 9 8 2
23 15 9 4 1 4 4 1 10 0 9 8 5 3 1 11 1 9 5 15 10 9 13 2
21 10 1 11 12 1 8 13 0 9 8 13 3 12 9 1 10 9 1 8 4 2
11 9 8 1 8 13 3 9 1 9 4 2
18 3 15 4 9 4 1 10 9 2 3 8 10 9 1 8 4 0 2
13 7 15 13 15 3 4 3 10 9 1 15 13 2
21 13 1 10 9 13 10 9 1 15 2 10 9 1 10 13 7 10 0 13 9 2
10 0 1 10 9 13 13 2 8 2 2
17 15 13 3 16 15 0 9 3 1 4 4 1 9 1 15 9 2
17 2 15 3 3 2 2 13 8 2 2 11 4 10 0 9 2 2
9 0 9 0 13 15 15 1 11 2
25 15 9 11 13 15 3 0 10 9 3 2 15 1 10 0 9 10 0 9 13 1 15 0 9 2
30 7 3 3 13 3 15 9 6 3 1 4 7 3 13 15 9 1 10 9 2 10 0 9 1 0 9 2 15 3 2
7 10 9 4 1 9 4 2
11 2 9 15 13 3 12 9 0 1 2 2
9 15 15 9 3 3 10 9 13 2
10 3 13 15 3 3 15 3 3 4 2
7 3 4 15 10 9 0 2
8 3 13 15 10 9 0 4 2
19 15 4 12 9 1 10 9 0 7 12 7 12 9 0 2 3 4 15 2
12 15 4 15 0 9 16 15 13 1 15 9 2
16 15 4 0 16 15 3 3 4 2 7 15 9 4 3 0 2
49 10 9 1 0 9 1 10 0 9 1 15 8 1 11 2 1 10 9 2 8 2 2 13 10 0 9 2 8 10 9 0 9 1 10 9 1 10 9 2 0 7 0 9 2 15 10 9 13 2
26 15 4 10 9 1 0 9 1 10 9 1 15 8 1 11 2 10 9 1 11 7 15 8 1 11 2
6 10 9 13 9 3 2
18 1 15 9 13 15 8 3 10 9 1 10 0 9 1 9 7 9 2
21 10 3 0 9 2 15 10 0 9 13 1 10 2 9 1 15 13 2 1 11 2
16 15 13 3 0 9 1 4 2 7 3 4 15 9 3 2 2
5 9 2 9 8 2
9 2 15 15 13 4 10 9 9 2
15 15 13 9 1 9 4 4 7 15 3 1 15 4 4 2
22 7 15 4 3 3 9 1 0 9 2 1 15 15 9 2 3 2 1 15 0 9 2
5 15 4 0 2 2
3 9 8 2
17 2 0 13 0 15 3 0 2 7 15 4 3 10 13 0 9 2
6 1 4 13 3 15 2
10 10 0 9 1 11 13 3 8 12 2
21 10 9 13 1 10 15 8 2 15 13 3 1 9 2 3 13 3 15 1 4 2
22 3 13 15 0 9 1 9 2 15 9 2 3 4 15 9 2 15 9 1 10 0 2
15 10 9 9 15 2 1 15 9 2 0 0 1 10 9 2
7 15 13 3 15 1 9 2
14 15 13 15 4 1 10 9 2 10 9 1 10 9 2
14 2 8 2 13 15 9 3 0 9 4 1 15 9 2
15 3 1 10 9 4 1 15 9 10 9 7 9 0 4 2
7 15 13 0 1 9 4 2
9 15 13 10 9 0 10 13 9 2
28 3 13 1 4 16 15 2 3 1 15 9 4 4 1 15 9 1 9 2 7 1 15 0 9 8 9 4 2
15 11 13 15 9 1 8 1 11 2 7 10 9 1 11 2
22 10 13 9 13 9 1 10 9 2 13 1 10 9 1 9 2 9 13 15 0 3 2
11 10 9 1 9 13 7 13 1 10 9 2
15 13 3 10 9 1 10 9 7 13 3 10 9 9 3 2
15 13 1 10 9 10 9 9 7 13 3 12 9 9 3 2
7 13 10 9 1 13 9 2
25 10 9 9 13 1 10 0 9 1 10 9 4 4 7 3 1 10 9 4 2 16 15 15 13 2
14 10 9 7 10 9 1 11 13 10 9 1 8 4 2
18 15 13 0 1 10 9 1 10 9 1 10 0 13 9 1 10 9 2
18 10 9 1 10 13 9 2 10 9 2 10 9 7 3 15 0 9 2
9 16 10 0 9 1 10 9 13 2
6 10 9 13 12 9 2
25 2 13 15 9 3 2 3 13 3 9 2 2 13 10 9 16 15 15 1 10 9 1 13 4 2
47 10 0 9 4 10 2 9 2 2 3 10 9 10 9 1 10 9 13 2 10 0 9 13 7 1 10 0 9 10 13 9 13 2 3 2 3 15 15 13 3 15 15 3 13 7 13 2
12 3 13 15 9 10 13 9 7 4 15 0 2
4 7 3 3 2
35 8 13 10 9 1 10 9 1 0 9 2 15 13 16 15 3 3 4 16 10 9 15 13 4 16 15 10 0 9 1 10 9 4 4 2
21 15 13 3 0 9 0 4 7 0 0 9 13 4 1 0 9 1 3 0 9 2
19 10 9 1 9 2 9 7 10 0 9 13 4 1 11 2 11 7 11 2
23 10 9 13 3 1 11 4 2 7 3 5 13 10 9 0 5 13 11 3 0 3 4 2
22 8 3 13 9 13 11 15 15 0 4 1 4 1 9 2 9 7 3 3 3 9 2
10 1 12 13 11 1 12 12 9 4 2
19 15 4 3 3 4 7 3 4 11 2 3 13 15 3 2 8 13 4 2
19 13 15 10 9 1 9 4 16 15 2 16 11 2 0 1 0 9 13 2
3 0 3 2
23 13 15 9 4 1 10 9 16 12 13 2 3 7 8 13 1 9 2 1 9 13 13 2
15 9 11 13 15 8 16 9 10 0 9 4 1 0 4 2
10 2 15 4 3 3 0 1 10 9 2
8 15 4 3 3 0 3 4 2
21 3 13 3 15 13 9 2 3 3 0 9 4 13 4 16 10 13 9 1 13 2
7 15 9 4 4 1 11 2
16 15 13 10 0 9 4 2 16 0 9 1 10 9 4 4 2
11 16 10 12 13 9 4 3 3 15 4 2
20 2 1 15 9 4 15 3 3 3 4 7 3 13 15 15 3 0 3 4 2
16 15 13 15 3 3 0 15 4 4 16 10 9 1 13 4 2
8 0 13 10 9 8 15 0 2
17 1 11 13 15 3 15 4 2 16 15 3 3 1 9 4 4 2
6 9 1 10 9 9 2
22 10 9 15 15 1 10 11 13 1 2 8 2 2 10 0 9 2 13 15 0 3 2
11 0 13 2 3 10 9 4 3 0 13 2
12 3 13 15 1 15 9 3 1 10 0 9 2
20 11 4 4 1 13 1 8 8 1 10 9 2 15 4 3 10 9 8 11 2
18 8 2 3 13 15 15 3 1 9 4 16 15 0 4 0 1 13 2
24 11 13 3 8 4 2 15 13 10 10 9 1 10 0 9 1 10 3 3 13 9 1 8 2
6 15 10 0 9 13 2
14 15 4 3 0 2 16 12 9 0 4 1 15 9 2
6 3 13 9 4 2 2
24 3 3 13 10 0 9 15 9 1 9 2 16 8 15 11 10 9 1 9 1 10 9 13 2
11 2 15 13 3 3 3 2 16 15 13 2
7 3 13 15 3 4 4 2
16 15 13 3 1 15 16 15 3 3 1 15 9 3 4 4 2
8 15 13 4 15 15 13 2 2
7 11 9 4 0 1 9 2
25 16 10 9 1 9 15 0 4 16 1 11 2 7 9 13 4 2 13 10 9 15 9 15 9 2
4 13 4 13 2
9 15 4 3 3 0 1 15 9 2
12 10 9 4 1 10 9 7 1 10 9 4 2
12 9 2 1 9 3 2 4 1 11 3 4 2
17 3 0 15 0 0 11 3 13 4 2 1 13 9 4 3 4 2
18 1 15 8 4 3 10 0 9 8 1 10 11 1 10 13 9 4 2
28 10 9 4 0 10 9 1 9 3 1 4 1 15 1 9 4 8 2 16 10 9 2 13 1 9 3 13 2
15 10 9 13 1 9 1 10 9 1 10 9 3 4 4 2
11 1 9 1 10 11 4 15 1 4 4 2
28 15 4 12 7 12 9 3 16 12 9 1 10 9 2 3 9 1 3 0 9 2 9 13 4 1 10 9 2
19 16 9 13 15 10 9 1 15 9 1 10 0 4 7 15 15 9 4 2
20 15 13 15 3 2 7 11 13 10 9 4 7 4 3 4 16 9 1 13 2
13 15 13 16 15 3 13 1 11 12 9 8 4 2
12 8 16 10 9 15 1 15 13 9 4 4 2
19 10 9 11 13 10 3 0 9 3 2 8 1 2 9 2 3 9 4 2
6 10 9 13 3 4 2
23 16 10 0 9 1 10 9 3 3 4 4 2 3 13 10 9 3 4 1 10 15 9 2
18 13 15 9 7 13 15 15 3 4 13 2 7 1 15 13 2 4 2
6 10 0 1 15 9 2
13 11 9 13 1 15 9 1 15 9 15 0 9 2
57 15 13 3 1 10 3 3 0 11 3 1 9 7 3 13 0 9 15 2 1 10 9 2 15 3 9 4 2 16 1 11 2 2 3 12 9 13 4 4 16 15 15 3 3 3 13 1 10 9 1 12 9 1 9 1 4 2
28 11 13 13 1 10 1 15 8 13 9 1 10 0 9 2 10 0 11 2 7 1 15 9 13 15 15 4 2
19 15 13 15 8 4 1 15 0 8 7 13 1 10 15 9 15 9 3 2
29 15 13 16 15 15 9 15 3 4 4 2 3 13 15 0 13 1 11 7 13 15 3 3 3 3 3 10 9 2
34 10 9 4 11 1 9 4 1 10 9 1 10 9 8 2 10 3 13 9 13 3 4 4 16 15 4 4 1 15 1 11 0 9 2
45 1 13 9 13 15 1 15 9 5 8 2 8 2 2 8 2 11 2 2 8 2 8 2 2 8 2 8 2 7 10 9 1 10 0 13 9 13 5 1 9 5 3 0 0 2
31 10 9 7 15 0 8 1 11 2 15 10 9 9 1 10 9 13 2 4 0 4 1 15 9 1 10 3 0 0 9 2
47 16 10 9 9 1 10 11 2 13 1 10 9 1 0 9 1 10 9 3 13 1 15 13 1 15 0 9 2 13 10 0 9 1 10 9 9 1 10 9 1 10 9 9 1 4 16 2
7 2 15 13 11 11 11 2
7 15 2 15 2 15 2 2
17 15 9 2 2 13 8 2 15 1 10 9 16 9 7 9 13 2
7 2 10 9 4 9 4 2
9 10 9 13 3 15 3 0 3 2
16 13 15 10 0 9 1 10 9 4 4 7 0 10 9 4 2
12 3 13 1 12 9 9 7 12 9 4 4 2
24 0 9 13 2 13 10 9 3 1 8 1 12 10 9 1 10 9 1 10 9 1 15 8 2
12 10 0 9 1 10 9 13 1 12 1 9 2
16 2 10 9 2 15 10 9 13 13 1 10 9 3 7 13 2
21 1 10 9 1 11 1 11 4 1 10 9 1 10 9 8 1 11 12 9 4 2
6 10 0 9 4 0 2
18 10 0 9 8 13 15 9 1 10 0 9 8 2 3 10 9 13 2
10 12 13 1 9 1 10 9 1 9 2
14 10 9 1 11 4 0 4 2 15 1 8 0 4 2
14 1 15 8 13 9 10 9 1 10 9 1 10 9 2
33 1 7 1 15 1 1 10 9 3 15 15 13 2 13 10 9 9 7 9 15 15 1 15 10 9 13 1 10 9 15 11 4 2
10 15 4 9 2 9 2 9 2 9 2
11 15 13 1 9 1 12 1 10 0 9 2
12 15 4 15 15 0 10 9 1 10 9 13 2
37 1 15 9 13 8 4 1 10 0 2 0 2 3 0 9 2 3 15 1 15 9 13 16 3 10 15 9 9 2 15 1 10 9 2 8 4 2
21 10 9 13 10 9 10 9 1 9 7 9 4 3 10 9 3 0 3 13 4 2
36 10 0 9 2 15 8 10 9 13 2 15 1 15 13 13 4 2 13 15 4 7 8 4 1 10 11 2 15 0 4 1 13 7 0 13 2
12 3 1 10 9 9 4 10 0 1 9 4 2
12 15 4 3 1 10 9 13 1 10 0 9 2
16 8 11 13 9 1 10 0 9 1 11 10 9 1 10 9 2
9 10 9 13 15 9 13 1 12 2
13 8 13 0 15 0 2 7 10 9 4 3 8 2
24 11 13 3 10 0 9 1 10 13 9 7 10 0 9 2 3 8 15 9 1 0 9 13 2
27 9 4 1 8 1 12 1 12 10 0 9 1 4 1 10 9 1 15 8 1 10 9 11 1 15 8 2
21 1 10 0 9 13 8 1 10 9 1 8 10 9 0 1 10 9 2 12 2 2
9 10 9 13 15 0 0 3 4 2
21 10 9 1 10 9 2 3 15 13 15 15 3 4 2 13 15 3 16 15 13 2
10 10 9 0 4 10 9 4 1 9 2
20 10 9 4 15 9 1 9 4 7 13 1 10 0 9 1 10 9 1 4 2
9 15 1 10 0 9 13 15 4 2
22 15 4 3 1 15 0 9 5 10 9 4 3 4 1 1 12 5 16 9 4 4 2
17 1 10 0 9 13 10 0 3 15 4 16 15 9 1 13 4 2
18 15 13 3 3 2 7 1 10 3 0 9 13 10 0 9 1 12 2
19 11 13 1 10 0 12 9 0 10 9 2 7 15 4 3 0 0 12 2
20 1 8 4 15 9 1 12 1 12 1 8 7 8 10 9 1 15 9 4 2
14 8 13 3 10 9 3 1 4 2 3 1 0 9 2
20 15 4 12 1 10 9 2 7 1 10 9 13 11 3 10 9 1 10 9 2
9 0 9 1 10 9 13 8 3 2
15 3 0 1 9 2 0 13 2 13 15 3 1 10 9 2
12 1 15 1 13 0 9 2 15 1 8 13 2
6 2 11 2 11 2 2
8 2 3 2 11 2 11 2 2
14 10 0 2 0 9 1 11 2 13 3 1 10 9 2
9 15 4 3 0 1 15 0 9 2
5 15 13 15 3 2
21 3 4 15 15 1 15 0 2 16 15 0 1 15 9 4 2 15 9 1 13 2
14 2 2 13 15 1 9 2 2 7 3 13 10 9 2
19 10 9 16 9 1 10 9 7 15 4 1 4 2 7 15 13 0 4 2
15 15 13 1 10 15 3 2 15 13 15 2 9 2 4 2
10 9 4 2 3 2 1 9 7 13 2
7 9 4 15 4 16 0 2
12 10 0 9 4 3 1 3 0 7 0 9 2
15 10 0 9 1 0 7 0 2 0 7 0 13 0 9 2
16 10 9 13 10 9 1 10 9 4 1 10 0 9 1 8 2
14 10 9 1 10 0 9 13 9 11 1 10 9 4 2
18 1 15 9 13 11 1 11 16 1 15 8 3 1 13 1 0 9 2
10 7 15 4 9 2 7 15 4 4 2
9 15 13 13 4 4 1 10 9 2
11 3 4 3 3 10 9 4 1 10 9 2
6 9 1 9 7 9 2
7 2 11 11 11 11 2 2
13 12 9 0 3 13 8 2 10 9 2 15 9 2
8 2 3 4 15 15 13 3 2
16 15 13 3 0 4 7 3 13 10 9 0 3 1 10 9 2
9 2 10 9 13 3 3 3 2 2
7 2 15 4 3 10 0 2
19 15 13 3 3 3 1 11 4 16 3 1 13 2 7 15 13 3 3 2
7 3 13 15 3 9 3 2
15 7 15 13 3 1 10 9 1 11 4 2 8 10 9 2
8 15 13 3 1 10 0 9 2
17 2 11 4 10 0 9 2 15 1 10 0 3 15 3 13 4 2
11 3 11 2 15 4 10 9 1 10 9 2
16 15 13 15 3 4 4 2 8 2 15 13 0 10 0 9 2
3 10 9 2
12 7 15 13 10 9 2 15 10 0 9 13 2
13 13 11 3 3 3 4 1 10 0 9 1 4 2
20 15 8 13 8 15 8 4 1 10 1 15 13 0 9 10 0 9 2 8 2
32 10 9 11 4 3 1 10 9 10 9 2 8 4 15 8 1 10 11 1 4 2 0 16 15 1 15 9 1 9 13 4 2
11 15 13 1 3 10 9 9 1 15 9 2
36 15 9 3 13 10 9 10 9 2 10 9 8 2 8 10 9 1 8 15 1 13 4 2 16 15 8 4 4 16 15 3 15 9 13 4 2
34 1 9 13 9 7 9 10 0 9 3 4 16 10 9 0 3 13 1 9 1 10 0 2 3 3 0 9 13 1 10 9 1 9 2
31 10 9 13 3 1 10 9 1 10 9 2 0 13 16 10 9 1 10 0 9 11 1 13 2 10 9 1 10 9 3 2
16 3 1 10 9 13 10 9 3 3 2 7 1 10 9 0 2
16 11 7 11 13 9 11 10 9 4 1 10 0 9 1 9 2
24 3 4 2 13 1 12 9 2 15 0 8 4 2 15 15 3 3 13 4 1 10 0 9 2
27 10 9 2 15 0 12 1 9 2 13 1 10 9 10 15 9 4 4 2 3 15 3 0 0 13 4 2
8 10 0 9 13 15 9 4 2
11 3 13 8 2 12 2 15 9 0 13 2
6 15 13 4 2 6 2
8 9 15 15 3 13 4 4 2
15 1 10 11 4 10 9 1 8 12 9 4 1 10 9 2
13 11 2 11 2 7 10 0 9 7 3 12 9 2
28 8 2 12 2 7 8 2 12 2 4 10 9 2 7 15 13 15 9 7 1 15 9 4 15 2 0 2 2
7 16 15 15 13 4 4 2
9 15 4 3 0 16 15 1 13 2
14 10 9 1 10 9 4 15 3 1 15 4 1 4 2
13 10 9 13 15 9 1 3 7 13 1 10 9 2
13 7 3 13 15 3 8 1 10 9 1 9 8 2
18 15 13 10 9 1 15 13 7 15 13 16 15 3 13 4 1 4 2
13 3 15 9 13 3 1 10 9 9 8 10 9 2
11 3 13 15 16 15 15 0 4 7 0 2
31 2 15 9 4 3 12 3 3 15 0 0 4 4 1 10 0 2 0 2 0 9 1 0 9 2 2 3 13 10 11 2
16 1 0 9 13 3 2 1 10 11 15 0 9 4 4 4 2
14 3 13 3 10 9 4 3 9 9 7 9 13 4 2
18 3 13 3 10 9 4 4 16 13 9 10 0 9 1 4 1 9 2
36 15 13 15 0 9 2 7 10 9 1 11 0 9 1 10 0 9 2 2 15 1 10 9 1 10 9 7 10 9 1 12 9 4 4 2 2
39 3 1 10 0 9 2 15 0 1 10 0 9 1 10 9 13 2 13 10 9 1 10 9 10 9 1 10 0 9 1 10 0 9 2 13 9 1 11 2
12 1 11 13 15 0 4 1 10 9 1 11 2
5 15 13 15 3 2
35 10 9 1 11 4 3 15 1 10 12 13 0 2 8 2 12 2 2 8 2 8 2 12 2 2 8 2 12 2 7 8 2 12 2 2
34 10 13 9 2 15 1 8 2 7 3 1 10 9 1 3 2 9 2 1 8 0 9 8 2 4 4 2 4 3 15 1 15 9 2
36 1 10 9 1 11 1 10 11 1 8 4 1 11 10 9 4 2 7 1 9 0 3 13 10 9 15 3 1 10 0 0 7 0 0 9 2
22 15 13 0 1 9 2 6 2 7 15 13 3 16 10 9 4 2 16 15 0 4 2
16 15 13 3 9 4 1 15 15 2 1 15 3 0 0 9 2
16 10 11 13 15 9 3 1 10 9 0 4 1 9 1 11 2
19 8 8 7 8 13 10 0 9 1 10 2 9 1 10 0 9 2 4 2
32 1 9 15 3 3 8 4 1 15 9 9 13 10 9 10 9 2 7 16 15 3 13 1 4 4 4 2 13 15 1 4 2
8 15 13 15 0 10 9 0 2
18 12 13 9 2 12 0 13 1 10 9 1 11 2 13 10 9 0 2
30 3 13 9 11 1 11 3 10 9 2 1 9 2 3 2 7 15 13 5 13 8 5 15 15 9 1 10 9 4 2
9 8 13 10 2 15 2 9 3 2
32 16 10 9 8 3 0 13 2 4 10 9 1 0 11 15 15 9 1 10 0 9 1 10 0 9 3 3 3 2 13 2 2
18 1 10 9 1 10 9 12 13 15 3 10 9 1 11 1 10 9 2
11 10 9 8 2 12 2 1 11 13 15 2
9 15 9 4 1 9 3 3 0 2
41 8 2 10 9 2 7 1 0 9 3 3 10 0 9 2 9 7 1 15 9 3 3 13 1 10 9 1 10 9 2 7 1 10 9 1 10 9 1 10 9 2
14 10 3 0 0 11 13 15 1 7 1 10 9 3 2
13 3 13 10 9 1 15 8 1 11 15 9 4 2
17 15 4 10 9 8 1 8 2 15 9 13 1 10 9 1 11 2
6 0 9 13 9 8 2
22 10 13 9 13 3 8 10 9 1 10 0 9 3 10 9 1 0 9 8 4 4 2
17 10 9 13 0 2 16 10 9 3 1 13 2 10 9 4 4 2
9 10 0 9 13 12 12 9 4 2
11 15 13 12 9 9 1 9 1 12 9 2
15 3 11 4 4 2 11 7 11 0 13 13 9 9 4 2
18 1 10 9 1 0 12 9 4 9 1 10 9 1 12 9 1 9 2
21 3 13 12 0 9 2 10 0 9 1 15 13 7 13 1 9 7 3 10 9 2
20 10 0 9 4 1 10 0 13 9 8 4 1 11 1 15 9 8 0 9 2
20 10 9 12 0 7 0 7 13 2 13 15 9 1 10 9 2 0 7 13 2
28 15 4 10 9 16 15 7 15 2 1 9 9 7 9 2 15 13 1 0 9 2 4 15 0 3 4 2 2
11 8 2 15 13 3 4 3 15 15 4 2
9 1 15 9 13 15 1 0 9 2
9 1 8 1 11 4 15 3 4 2
12 15 13 3 0 1 10 9 4 1 15 9 2
38 3 16 10 9 15 7 15 13 9 3 3 3 13 3 4 4 1 10 9 1 10 9 2 13 10 9 1 10 9 7 15 1 10 9 3 4 4 2
3 15 13 2
30 15 2 1 10 9 1 15 0 9 15 0 9 13 10 9 1 15 8 8 1 10 9 1 10 9 1 10 9 12 2
18 10 9 13 4 16 15 1 12 3 12 9 1 10 0 9 4 4 2
14 11 13 1 10 9 1 10 9 10 9 1 11 4 2
20 10 0 9 13 1 10 9 1 9 10 9 1 10 0 9 11 1 15 3 2
22 10 9 1 11 13 1 10 0 9 9 2 16 15 1 1 9 0 9 10 9 13 2
9 8 4 1 12 9 10 0 9 2
8 8 13 1 10 12 15 9 2
25 1 10 0 9 13 8 3 10 0 9 1 10 9 16 1 10 9 1 8 3 1 13 2 12 2
17 10 9 13 0 16 8 7 8 1 0 13 1 9 8 13 4 2
24 10 9 4 16 8 2 10 9 1 11 2 13 16 15 0 8 1 4 1 10 0 9 8 2
16 2 13 15 3 9 4 1 10 0 9 1 10 9 1 11 2
15 1 10 0 9 13 8 9 10 9 1 12 3 1 4 2
13 1 11 13 15 1 0 13 10 9 0 1 4 2
20 1 11 13 10 0 9 3 16 10 12 9 7 10 9 10 9 8 13 4 2
22 1 11 13 10 9 2 16 15 3 1 10 15 9 1 10 9 1 10 9 4 4 2
24 10 0 9 13 1 10 0 9 15 1 10 0 9 4 4 3 1 10 9 3 10 9 13 2
49 7 10 15 13 1 15 9 2 10 15 13 0 3 1 15 9 1 9 2 10 0 13 15 9 3 1 4 1 15 15 9 11 12 9 1 10 0 9 1 10 9 10 15 2 0 9 13 4 2
16 0 16 15 1 10 0 9 1 9 3 15 9 13 4 4 2
12 13 15 4 1 10 9 1 10 9 1 8 2
19 2 15 13 16 11 0 1 15 4 4 16 15 1 9 11 4 4 2 2
25 11 13 15 1 0 9 4 4 2 7 1 15 9 1 13 7 16 15 1 13 9 3 1 13 2
18 2 6 2 11 13 3 9 16 3 5 1 15 5 10 10 9 13 2
22 15 4 10 9 1 10 0 9 1 10 2 9 2 1 11 15 11 1 11 4 4 2
32 11 13 15 0 4 2 13 15 1 10 9 4 4 2 9 1 10 9 4 0 16 9 1 10 9 2 2 4 15 13 9 2
28 1 15 9 13 9 11 0 3 1 10 9 1 9 11 2 3 5 8 10 9 5 10 11 0 9 4 4 2
27 2 15 13 10 9 2 2 3 10 9 11 2 2 16 10 9 15 4 4 16 10 9 9 1 10 9 2
32 2 16 10 9 13 16 9 1 10 11 3 8 13 9 4 2 3 13 15 10 9 1 10 9 2 15 1 15 9 8 4 2
19 8 13 3 3 0 1 9 2 15 15 0 3 13 7 3 13 4 3 2
10 3 13 15 15 16 15 2 8 2 2
30 15 13 10 0 9 9 2 3 10 9 9 0 13 1 4 16 15 0 9 2 3 15 0 13 10 0 9 1 4 2
15 0 4 15 3 3 3 1 15 0 0 9 1 15 9 2
8 15 4 9 3 2 13 15 2
23 1 12 9 13 9 8 2 8 2 8 2 11 2 10 9 1 15 1 12 13 0 9 2
20 15 4 3 3 0 2 7 15 15 2 9 2 3 13 4 15 13 10 9 2
7 15 13 15 3 12 3 2
19 10 0 9 7 10 0 13 9 2 15 10 9 1 10 0 9 13 4 2
25 10 9 15 10 9 1 10 9 10 0 9 1 9 13 4 13 1 10 9 15 0 0 9 4 2
23 7 10 9 13 3 10 0 9 16 15 9 4 1 10 13 9 1 9 2 9 2 9 2
9 0 4 3 10 0 9 8 4 2
9 15 9 13 15 3 15 9 4 2
31 15 8 1 11 2 10 9 1 10 9 2 9 10 9 11 2 16 15 15 9 4 4 16 15 1 9 3 8 1 13 2
29 1 10 13 9 13 10 9 11 2 15 9 1 10 9 2 1 10 9 1 10 11 3 3 10 9 1 10 9 2
15 10 0 9 1 10 9 13 1 8 15 13 1 10 9 2
38 2 15 13 1 15 9 0 1 2 2 13 3 10 0 0 9 8 1 11 2 15 15 9 16 0 10 12 9 1 10 9 1 10 9 0 13 4 2
44 16 9 8 1 11 13 2 3 0 1 4 16 10 9 4 4 2 2 7 15 1 15 9 4 4 16 10 9 1 10 9 1 4 2 13 11 16 11 3 10 0 9 4 2
22 3 13 15 8 3 10 9 1 10 9 2 15 3 3 1 9 1 10 9 4 4 2
19 10 9 1 11 13 1 8 10 9 1 10 9 1 10 9 1 10 9 2
14 10 9 13 8 1 12 9 1 10 9 1 10 11 2
26 10 9 8 1 10 9 13 3 10 0 9 1 10 9 1 9 7 9 2 3 10 9 9 13 4 2
8 10 9 1 10 9 4 4 2
17 8 1 11 2 9 2 13 10 9 3 1 4 1 10 0 9 2
19 0 9 5 3 13 15 5 13 3 13 1 0 9 7 13 10 9 3 2
25 15 9 13 3 1 10 9 2 16 9 10 9 4 2 15 0 4 1 10 9 1 10 9 2 2
20 7 16 3 3 3 4 13 4 2 3 0 1 9 16 1 9 2 13 8 2
18 9 1 12 13 15 3 1 10 9 16 15 10 12 9 0 4 4 2
17 1 10 9 1 10 9 15 15 9 13 2 13 10 9 3 3 2
14 10 0 9 3 2 16 10 0 9 10 0 9 4 2
16 10 0 9 2 3 15 10 0 9 4 1 10 9 2 13 2
5 9 1 10 9 2
18 15 4 16 9 0 7 13 3 10 9 16 15 9 9 4 4 4 2
14 7 2 9 2 1 10 9 7 2 9 2 1 0 2
6 15 4 8 9 4 2
14 0 1 15 4 1 15 9 10 13 7 0 9 4 2
9 15 13 1 10 9 16 15 13 2
26 16 9 11 13 15 9 1 9 1 4 4 2 13 15 15 9 1 0 15 9 12 9 3 0 3 2
12 15 13 1 9 3 16 3 0 9 13 2 2
14 1 0 9 7 13 9 4 10 9 13 3 1 4 2
28 1 15 10 9 3 3 13 9 1 2 9 2 9 2 9 7 9 2 13 3 10 0 9 2 0 7 0 2
19 15 4 3 15 0 0 9 2 0 3 16 15 15 13 1 10 0 9 2
24 10 9 2 10 0 9 2 10 15 0 9 7 3 10 9 13 10 11 10 0 0 9 4 2
52 7 3 13 12 9 1 11 2 10 9 7 10 9 13 0 4 16 15 12 9 1 9 13 2 10 9 1 12 9 1 9 4 10 9 1 15 9 5 7 15 16 10 9 3 0 4 2 3 1 0 9 2
17 10 9 2 15 0 4 16 0 1 4 4 15 15 8 13 2 2
33 10 9 9 2 15 9 2 2 15 13 15 9 16 1 15 13 9 3 3 10 9 3 1 4 2 2 13 11 3 1 15 9 2
23 1 10 9 9 4 15 0 10 9 3 1 4 1 9 2 15 8 10 9 13 4 4 2
45 16 15 15 9 4 1 10 9 2 13 15 3 2 7 1 15 9 13 15 8 1 10 0 9 1 10 9 2 1 0 3 16 9 3 10 0 2 0 9 2 3 11 4 4 2
24 16 15 15 12 4 4 7 15 15 8 13 4 2 4 0 9 10 0 9 1 9 7 9 2
16 2 15 4 3 3 4 2 16 15 12 9 1 10 9 4 2
13 1 15 0 9 13 15 3 3 9 7 9 3 2
23 10 9 8 2 0 9 1 10 0 9 1 11 2 4 3 0 13 1 15 9 1 9 2
22 0 13 15 1 15 9 4 7 3 3 13 15 1 4 2 16 3 15 3 3 4 2
19 15 13 15 3 4 15 9 1 4 2 7 15 13 15 1 15 4 2 2
21 8 13 1 10 13 9 1 10 9 11 15 1 15 8 13 8 1 15 9 4 2
11 11 13 1 9 12 12 9 1 12 9 2
7 11 4 0 1 12 9 2
20 11 13 5 1 10 13 9 1 8 2 11 2 5 1 12 9 10 12 9 2
20 8 13 15 3 1 15 15 0 9 2 16 15 1 10 0 9 9 13 4 2
12 15 4 3 15 15 0 2 10 9 4 0 2
44 10 0 9 1 10 9 1 15 8 2 13 1 8 13 8 15 9 1 10 0 9 2 11 2 2 0 10 9 2 7 3 10 16 3 10 9 16 2 8 2 4 4 4 2
31 15 13 2 16 10 0 9 1 10 11 0 12 9 4 4 13 3 3 1 4 16 1 13 15 15 1 10 0 9 4 2
20 1 11 2 10 9 1 10 0 9 1 10 0 9 2 13 15 3 3 0 2
21 7 7 8 2 7 10 11 13 0 10 0 1 11 2 3 13 11 3 3 4 2
10 9 3 3 16 15 11 15 9 13 2
12 15 13 8 12 9 16 15 9 0 1 13 2
22 8 2 15 13 15 3 4 1 11 2 16 15 3 3 3 1 11 4 16 15 13 2
15 11 13 3 12 12 1 15 2 15 4 12 9 1 9 2
14 7 3 13 15 3 9 4 1 10 0 9 7 9 2
11 13 3 3 1 10 0 9 0 9 3 2
8 10 9 13 10 9 1 9 2
17 10 9 4 3 2 16 15 3 3 0 4 2 16 10 9 13 2
8 13 4 3 13 1 0 9 2
9 7 2 15 13 1 0 9 4 2
15 3 4 1 11 7 11 12 9 2 15 15 1 13 13 2
18 10 9 1 9 1 11 13 0 3 7 3 10 9 4 1 10 9 2
14 15 9 1 9 8 13 3 10 9 1 10 0 9 2
37 1 10 9 1 10 9 2 15 1 0 3 13 2 4 10 9 13 1 10 9 4 16 1 10 0 9 1 13 1 15 0 1 10 9 13 9 2
2 7 2
43 2 16 15 9 4 1 10 0 0 11 2 7 1 10 9 1 13 1 10 9 2 4 15 3 15 9 16 10 13 9 1 10 0 9 2 15 1 15 0 9 13 2 2
2 7 2
20 10 9 13 0 4 4 2 7 16 15 15 9 4 4 2 13 10 9 3 2
27 2 16 2 9 10 9 2 3 8 2 4 4 2 13 3 1 15 9 4 2 7 3 1 15 3 2 2
15 3 4 10 9 13 2 3 9 9 13 2 3 3 4 2
25 15 9 13 3 1 10 9 1 10 0 2 0 2 9 1 11 2 8 2 1 10 9 1 11 2
26 1 10 0 9 13 10 0 9 2 15 15 9 7 3 3 10 9 15 13 16 15 9 3 1 13 2
22 10 0 2 0 9 2 15 13 1 10 9 13 2 7 3 13 1 10 9 1 9 2
20 2 15 4 0 1 10 9 5 15 13 3 9 2 6 9 5 1 10 0 2
13 10 9 13 0 4 2 7 0 4 15 0 2 2
17 10 0 9 4 3 0 3 1 4 1 10 9 1 11 1 12 2
23 7 10 9 2 1 15 9 13 2 13 15 3 4 1 10 9 3 1 13 1 10 9 2
8 10 9 13 10 11 3 4 2
8 15 13 9 1 15 3 16 2
11 10 0 9 13 1 10 9 1 10 9 2
10 11 13 10 0 9 1 10 9 0 2
32 15 4 3 10 9 2 15 13 3 15 12 9 3 2 7 15 13 3 13 3 16 15 15 9 0 3 1 10 9 13 4 2
16 15 13 0 3 4 16 15 3 13 0 10 0 9 1 4 2
27 3 13 15 9 1 15 8 2 10 0 9 15 15 9 4 2 7 3 3 8 2 10 15 16 15 8 2
29 3 4 0 9 11 1 10 9 1 10 9 15 4 2 3 15 13 4 16 3 2 3 0 2 13 15 9 4 2
7 10 11 4 10 0 9 2
6 10 9 1 0 9 2
20 10 0 9 3 2 7 3 15 15 9 13 2 3 10 15 3 3 1 13 2
30 3 4 15 3 3 16 15 15 0 16 15 0 4 2 7 15 1 4 13 2 13 4 16 0 9 1 9 1 4 2
15 0 13 7 13 2 10 9 13 0 4 2 15 4 0 2
33 11 4 0 10 9 2 10 9 4 10 9 2 2 7 15 4 3 1 10 0 11 4 2 16 15 3 13 3 15 3 4 4 2
20 10 9 9 4 1 10 0 9 10 9 1 10 3 0 9 11 2 12 2 2
12 11 4 1 3 0 9 3 9 1 8 4 2
15 15 4 0 2 16 10 9 1 15 9 10 0 9 13 2
26 3 16 15 15 13 1 10 0 9 2 3 13 15 11 10 10 9 4 2 1 10 0 9 1 11 2
30 11 13 10 0 2 0 1 10 9 4 1 10 13 7 0 9 2 7 15 13 1 11 0 9 8 3 3 4 4 2
8 10 9 4 15 9 1 15 2
9 10 0 9 13 11 1 10 9 2
17 11 13 7 3 4 2 11 2 11 7 11 2 7 15 4 9 2
19 16 3 15 13 9 4 2 13 15 10 9 3 12 12 9 1 9 4 2
10 3 15 0 13 1 11 0 9 4 2
27 15 4 15 3 3 0 2 16 10 9 10 9 1 15 9 13 1 9 8 15 9 2 2 3 10 9 2
21 8 2 11 7 15 8 13 15 9 3 4 1 10 0 9 1 0 9 7 9 2
22 10 0 9 8 2 3 11 2 13 15 3 3 13 9 4 1 12 9 8 1 13 2
21 15 1 8 2 9 1 9 7 9 2 7 15 8 2 9 3 13 1 9 2 2
17 8 4 10 3 0 9 2 15 15 8 4 13 10 9 1 4 2
38 15 13 15 4 16 1 15 9 1 10 9 2 1 10 0 9 1 10 9 2 0 9 1 13 2 15 10 9 1 10 9 1 10 9 3 13 4 2
24 0 1 12 1 12 9 13 1 10 0 9 7 15 13 3 1 10 0 9 3 3 1 13 2
28 15 4 3 1 4 16 10 9 1 10 9 2 15 3 0 0 4 1 10 9 2 1 10 9 3 4 4 2
21 10 0 9 1 9 13 15 13 1 10 11 1 0 9 1 10 13 9 1 9 2
16 3 4 3 4 1 10 13 9 2 15 10 13 0 9 13 2
25 10 0 9 13 1 9 10 15 9 1 10 15 1 10 11 7 13 15 9 3 0 0 4 4 2
16 15 13 4 3 10 9 1 8 4 2 2 3 10 9 8 2
12 1 10 9 4 10 9 1 9 4 2 8 2
30 2 10 0 9 7 9 2 0 0 9 1 15 0 9 2 9 1 10 9 7 9 1 10 9 1 10 0 9 2 2
32 10 9 13 16 10 9 10 9 1 10 11 4 4 2 2 16 3 1 15 8 10 9 16 0 9 1 15 9 13 4 2 2
46 3 13 15 2 13 1 10 13 9 1 10 0 9 2 3 15 9 3 3 2 16 15 9 15 4 4 4 1 0 9 1 10 13 9 7 16 16 15 9 9 1 0 9 13 4 2
24 15 13 1 10 0 9 15 1 10 9 4 4 7 1 10 13 9 1 10 9 1 10 9 2
19 0 4 1 10 9 4 1 10 9 1 10 0 9 1 10 13 0 9 2
29 0 7 0 13 15 9 4 4 1 0 9 1 10 9 1 11 13 0 9 7 1 10 9 1 10 11 1 11 2
10 16 15 9 4 4 13 10 9 4 2
10 1 3 13 10 0 0 9 0 2 2
19 15 13 16 16 10 0 9 3 1 11 4 4 2 10 15 3 4 4 2
15 10 9 1 15 8 13 1 15 8 10 13 9 1 11 2
19 15 13 3 3 0 4 16 11 15 0 13 1 11 7 15 15 0 9 2
32 10 10 16 12 9 15 8 1 15 12 9 13 7 15 1 12 1 4 4 1 10 11 1 11 2 4 3 4 1 10 9 2
24 15 2 15 15 0 9 1 10 9 4 13 2 13 3 5 1 12 5 3 1 8 1 11 2
33 10 0 0 9 1 8 2 3 15 9 13 1 10 9 1 15 8 1 11 2 4 3 2 1 12 2 1 15 8 1 11 4 2
25 10 1 10 9 0 9 0 9 4 1 9 1 9 1 10 15 9 4 7 1 10 13 9 4 2
12 15 3 3 0 9 2 9 3 4 3 4 2
12 1 10 9 1 10 13 0 9 15 9 13 2
12 10 9 7 9 1 10 9 0 9 4 13 2
22 1 9 1 15 9 5 1 9 1 10 9 13 15 0 4 2 1 15 9 13 4 2
27 3 13 10 9 1 10 0 9 1 11 10 0 9 1 15 9 2 15 3 1 10 9 9 3 3 13 2
38 15 4 3 0 2 16 15 8 1 0 9 0 13 4 1 10 9 3 9 11 13 4 2 9 3 1 4 1 0 9 15 4 4 1 10 0 9 2
11 3 13 1 15 9 12 0 9 4 4 2
35 3 13 10 9 1 15 0 9 5 15 0 4 16 2 1 9 2 10 0 9 10 9 1 9 3 13 4 4 5 1 12 9 4 4 2
33 3 13 10 9 3 2 3 13 16 15 2 16 10 9 1 15 1 13 2 2 10 9 13 2 11 2 8 2 1 10 9 2 2
10 9 13 15 3 10 9 9 3 4 2
27 10 9 1 8 13 10 9 2 10 9 13 1 10 9 7 3 13 3 10 9 1 2 10 0 9 2 2
11 1 10 9 1 10 9 4 10 11 4 2
26 1 12 8 13 10 9 10 9 1 10 9 1 10 11 1 15 8 1 10 9 1 9 1 10 9 2
5 12 9 4 4 2
12 3 4 10 0 9 9 1 9 7 9 4 2
18 15 13 15 3 2 9 1 10 11 7 0 7 0 9 15 15 4 2
8 2 6 2 3 13 10 0 2
12 1 15 9 4 10 9 1 10 13 9 4 2
17 10 9 13 3 10 9 4 3 9 4 4 1 15 13 1 9 2
28 10 9 1 11 2 3 15 3 9 13 1 12 9 1 9 2 4 0 1 10 1 3 0 9 13 0 9 2
28 10 11 13 3 10 9 4 1 15 9 1 9 1 10 9 10 9 1 11 1 4 2 7 3 0 1 4 2
20 1 9 3 1 10 13 9 2 1 10 9 0 13 2 13 15 13 4 4 2
12 11 13 10 0 9 1 10 9 1 12 9 2
17 10 9 13 15 3 0 2 8 2 15 2 8 2 1 4 4 2
7 3 4 3 15 0 9 2
2 8 2
7 10 0 9 1 10 9 2
22 16 15 0 10 9 13 4 1 15 9 2 4 15 15 3 10 0 9 1 15 0 2
43 6 2 10 9 1 2 15 4 12 1 11 2 7 3 2 1 9 1 11 2 11 7 11 2 1 9 0 10 9 7 10 9 3 2 1 10 9 1 2 0 2 9 2
13 10 2 0 2 9 1 11 4 3 3 0 0 2
25 1 10 9 4 1 9 12 9 11 4 1 10 1 10 9 2 11 2 1 11 13 9 1 11 2
21 15 13 4 16 1 10 12 0 9 2 15 0 12 3 15 2 0 9 2 13 2
53 1 10 9 1 8 5 15 2 11 2 13 8 10 9 1 0 9 8 5 13 15 16 15 9 3 3 1 10 9 4 4 4 7 3 13 3 3 15 13 16 0 15 9 15 9 1 10 0 9 13 1 11 2
12 9 13 15 12 9 1 10 11 10 0 4 2
8 1 12 9 13 10 0 9 2
7 8 13 1 15 9 8 2
18 2 15 4 1 10 9 4 2 7 3 1 10 9 1 10 13 9 2
24 15 13 1 10 0 9 2 15 3 0 13 13 4 7 3 13 13 4 1 0 13 7 13 2
22 15 13 0 10 0 9 4 1 10 0 9 7 15 0 4 1 15 9 1 10 9 2
12 1 15 9 13 15 15 15 15 9 13 2 2
22 3 8 2 15 5 16 15 13 5 15 1 10 9 1 10 9 10 0 13 2 13 2
24 2 15 13 16 16 15 3 1 11 0 13 4 2 15 10 13 9 3 1 15 8 4 4 2
5 15 9 13 11 2
22 7 16 15 13 1 10 9 2 15 15 10 0 9 3 1 11 13 2 3 13 15 2
6 3 4 15 4 2 2
11 2 11 13 3 1 10 9 4 4 4 2
14 15 13 3 10 9 3 4 4 7 9 1 15 4 2
28 7 15 13 15 0 1 10 9 2 7 15 9 7 9 13 0 1 15 9 7 3 13 15 15 0 15 4 2
7 15 4 4 1 10 9 2
28 7 10 9 4 3 13 4 1 15 0 9 2 15 0 1 3 4 13 4 4 5 10 9 4 0 7 0 2
7 15 13 0 4 4 2 2
34 8 7 8 2 10 9 9 2 15 3 3 1 10 9 13 2 1 8 7 1 11 2 13 3 1 11 15 9 1 10 0 0 9 2
36 10 9 1 15 8 2 15 10 9 1 10 9 13 2 4 1 15 0 8 1 0 9 4 1 10 9 1 10 13 9 2 15 1 12 13 2
14 3 4 10 9 15 0 7 0 4 7 10 9 0 2
23 10 0 9 13 1 10 9 1 12 9 2 3 1 12 9 2 1 12 9 7 3 0 2
19 10 15 9 1 10 12 9 9 2 3 9 4 4 2 13 15 0 9 2
8 11 4 3 9 1 11 4 2
22 1 10 0 9 1 10 9 1 10 9 13 10 9 1 15 9 10 3 13 11 12 2
5 10 9 4 12 2
9 8 11 9 1 11 15 0 9 2
43 4 4 10 9 1 10 9 12 3 1 4 16 15 3 1 10 0 9 15 1 11 13 9 1 11 4 4 2 1 13 7 10 9 1 10 9 1 10 9 4 4 4 2
7 11 13 10 9 1 12 2
16 9 8 13 3 0 16 0 15 9 11 1 10 0 9 4 2
10 9 11 13 0 1 11 1 11 4 2
11 15 16 1 13 16 3 3 0 9 13 2
24 1 0 9 13 15 12 9 1 10 0 9 4 7 15 13 3 12 12 9 1 9 4 4 2
14 10 9 13 10 9 1 10 0 9 0 16 10 9 2
20 15 1 10 9 4 10 9 1 11 11 2 15 3 0 4 1 10 0 11 2
48 10 9 8 2 10 9 1 10 9 15 3 3 12 9 1 10 9 13 1 10 9 1 10 0 9 11 2 13 1 10 9 1 11 10 9 4 1 10 0 11 2 9 1 15 2 8 2 2
27 10 9 13 10 9 3 0 2 16 15 8 13 4 4 10 9 1 3 8 1 10 9 11 3 1 4 2
20 16 1 10 9 15 9 4 4 2 13 11 15 11 1 10 9 1 11 4 2
23 16 10 9 10 3 0 9 1 9 1 3 15 9 13 2 13 1 15 9 10 0 9 2
17 7 15 10 0 9 13 2 10 9 1 10 9 13 15 3 4 2
26 2 15 4 3 2 16 10 9 13 2 7 15 10 9 13 2 15 13 16 10 9 3 9 3 4 2
35 10 9 2 16 3 1 10 9 3 10 9 4 1 10 0 0 9 2 13 9 8 1 15 3 4 2 7 15 13 8 3 3 0 4 2
23 15 9 4 2 4 15 2 3 0 1 4 1 15 9 9 8 1 11 13 1 10 9 2
23 2 10 9 4 15 10 9 3 0 13 2 15 11 4 2 15 15 3 13 7 13 4 2
13 15 9 1 12 13 15 7 15 13 15 3 2 2
36 1 10 9 1 10 11 13 15 9 0 7 1 11 4 2 3 13 15 2 11 7 3 4 1 9 2 15 0 3 1 9 11 13 4 4 2
13 10 9 13 15 1 15 9 3 10 15 1 11 2
16 3 8 9 8 2 15 1 10 0 9 10 9 9 0 9 2
19 11 13 15 9 16 15 1 10 9 1 10 0 9 1 10 9 1 4 2
19 3 10 9 13 1 0 9 9 1 10 9 15 9 2 8 1 11 3 2
24 13 13 3 3 3 15 1 11 2 7 1 0 13 4 1 10 0 9 10 9 1 12 13 2
11 3 8 13 1 12 9 1 10 0 9 2
10 15 13 11 9 1 11 1 9 4 2
17 15 13 2 16 15 9 0 10 9 1 10 2 0 2 9 4 2
16 15 13 15 10 9 4 7 3 13 10 9 0 9 3 4 2
11 11 13 15 1 10 0 9 4 4 2 2
5 11 13 11 4 2
3 0 3 2
14 7 10 0 1 10 9 13 3 15 0 1 10 9 2
39 1 3 0 9 13 3 1 10 0 9 1 10 9 1 10 9 1 11 2 11 2 10 9 4 1 15 12 0 0 9 2 15 3 1 12 10 9 13 2
53 1 15 9 1 15 0 7 0 9 1 10 9 1 15 9 2 1 15 15 3 1 11 10 13 9 13 2 4 10 0 0 7 3 0 11 0 1 10 9 4 16 10 0 9 7 10 15 2 0 9 1 13 2
35 15 13 10 9 3 1 10 9 1 15 9 15 8 2 3 10 9 1 10 1 15 0 9 4 4 2 4 4 1 10 0 9 7 13 2
16 9 13 15 13 1 10 9 1 15 8 3 15 8 4 4 2
24 12 0 13 0 9 2 15 1 10 9 1 10 9 1 9 13 2 13 10 9 1 11 9 2
31 15 13 12 9 1 9 2 8 7 8 2 7 4 1 15 9 4 1 7 10 9 2 7 12 2 12 7 12 9 9 2
12 3 0 10 9 4 15 4 4 2 4 9 2
5 10 9 4 13 2
9 3 13 15 9 1 9 7 9 2
2 8 2
10 2 10 9 13 15 9 1 10 9 2
23 10 0 9 2 15 13 1 10 9 9 13 11 1 11 10 0 9 1 11 1 12 4 2
7 15 13 3 1 15 9 2
11 1 10 9 13 10 9 10 9 1 12 2
24 10 9 1 11 4 4 1 11 2 0 7 0 9 2 7 1 11 1 11 2 0 9 2 2
5 3 4 12 9 2
16 1 11 13 10 9 1 11 7 11 1 15 0 2 12 2 2
9 15 9 4 3 1 10 9 4 2
28 1 10 0 9 1 11 13 15 4 16 9 15 1 10 13 9 9 13 2 3 0 10 9 1 15 9 4 2
16 15 13 0 10 9 1 9 7 10 3 13 9 1 10 9 2
38 10 0 9 16 9 3 9 4 16 9 2 13 1 15 9 4 4 1 15 3 15 13 1 9 7 9 2 3 13 9 11 3 1 10 0 9 11 2
12 11 13 15 9 12 9 16 9 1 15 9 2
21 15 13 10 9 1 10 9 1 2 10 9 1 9 1 10 0 2 7 15 15 2
7 2 15 13 15 0 0 2
24 15 13 15 1 15 9 0 1 10 2 0 9 2 15 4 4 1 10 9 1 10 9 3 2
14 1 15 9 13 15 10 9 1 10 9 0 9 4 2
23 10 9 4 3 0 7 10 9 4 3 1 4 2 7 10 9 13 16 15 15 0 4 2
22 8 2 15 15 0 9 13 16 10 0 9 2 4 3 3 15 15 9 1 9 4 2
12 13 15 0 15 0 8 3 1 10 0 9 2
2 11 2
3 2 8 2
11 8 13 3 1 9 7 13 15 0 4 2
9 15 13 15 3 0 3 0 4 2
11 15 0 13 15 9 3 3 0 4 2 2
32 15 13 3 3 0 8 1 11 15 3 10 9 13 4 16 9 1 4 4 1 10 9 15 1 11 0 1 11 13 4 4 2
31 1 10 9 13 10 9 1 11 2 10 9 1 11 7 10 9 1 11 1 11 16 1 13 15 15 3 4 4 4 2 2
5 8 1 15 9 2
15 2 15 13 10 9 16 15 4 4 1 10 9 1 8 2
24 1 10 1 9 13 9 4 3 15 9 1 3 4 7 15 13 3 8 10 12 0 3 3 2
15 15 0 4 8 1 10 9 1 11 7 8 1 15 8 2
24 15 15 15 13 4 13 4 4 1 15 9 15 8 15 13 1 10 9 1 10 9 1 11 2
27 2 15 13 15 3 15 3 4 1 10 9 2 3 15 15 8 13 16 15 15 3 1 15 9 3 4 2
27 1 10 9 13 15 9 1 15 9 7 13 15 16 15 0 4 4 4 3 3 10 9 1 15 1 13 2
27 1 10 9 3 2 7 1 10 9 1 10 9 13 15 4 16 9 7 15 9 15 3 4 4 4 2 2
10 15 13 3 10 10 9 1 4 4 2
12 10 9 13 0 7 15 13 3 0 9 2 2
13 11 13 15 9 10 0 9 1 10 9 1 8 2
10 9 11 1 11 13 1 10 9 3 2
5 2 15 3 0 2
5 15 4 0 2 2
22 10 9 13 3 1 10 9 15 15 3 0 0 1 10 9 1 10 9 8 13 4 2
39 10 13 0 9 1 10 9 1 10 0 9 13 15 9 1 9 2 7 3 3 1 9 4 2 7 1 15 9 1 13 13 3 8 0 9 10 9 4 2
41 10 9 1 10 12 9 13 9 11 2 15 0 8 1 11 7 10 0 9 8 4 1 12 1 8 4 2 13 1 10 9 12 9 0 9 10 9 3 1 4 2
27 15 4 12 4 7 10 9 2 12 9 7 10 9 2 15 1 15 3 12 9 0 4 2 4 8 4 2
21 10 9 1 10 9 2 9 8 13 9 11 0 9 0 1 9 1 15 9 4 2
7 15 4 10 9 3 2 2
8 3 13 3 15 9 1 11 2
8 15 13 1 15 9 7 9 2
7 3 13 3 15 16 8 2
3 8 13 2
11 2 15 13 3 3 4 10 9 1 4 2
24 15 13 3 3 10 0 9 4 1 1 15 0 0 7 0 9 15 15 3 0 3 13 4 2
32 7 15 13 3 4 10 9 3 16 15 10 9 4 2 3 13 15 1 15 9 10 0 9 1 10 9 16 15 0 13 4 2
18 3 13 1 10 9 2 3 3 15 12 9 4 4 2 8 1 4 2
14 2 15 13 1 4 16 10 11 15 3 15 4 4 2
9 1 15 9 13 3 15 1 3 2
16 10 0 15 15 13 4 4 15 13 7 9 13 1 15 9 2
12 13 9 3 15 13 2 13 10 9 2 13 2
41 15 0 7 0 13 1 8 1 15 8 1 12 2 3 15 16 2 9 1 10 9 2 1 2 11 11 2 9 13 2 13 3 3 16 15 1 11 15 4 4 2
20 16 1 11 1 4 2 3 15 9 1 0 9 2 9 2 9 2 9 2 2
34 15 15 3 1 3 1 1 8 4 4 2 4 8 3 3 10 0 9 1 10 9 15 3 13 4 1 10 9 15 11 15 4 13 2
2 11 2
15 2 15 13 0 12 9 8 2 7 3 0 13 15 9 2
29 0 2 16 15 15 9 3 10 9 13 16 3 1 4 16 10 9 2 13 15 15 0 9 4 16 15 1 13 2
15 8 4 15 12 9 3 16 8 9 1 9 1 11 13 2
26 10 9 13 1 10 9 2 11 2 1 10 3 1 9 13 11 7 13 1 10 11 1 11 1 11 2
22 1 15 9 4 11 10 9 2 3 15 15 1 9 7 9 1 13 13 10 9 13 2
17 3 13 9 9 7 9 2 3 4 9 4 7 3 13 10 9 2
16 15 13 8 9 7 4 13 1 15 10 0 9 1 10 11 2
30 2 15 13 3 0 4 16 1 11 9 1 13 2 15 4 3 3 0 1 10 9 1 9 1 11 7 11 2 2 2
24 15 4 10 9 8 1 11 2 8 7 8 1 11 2 8 1 11 2 8 7 8 1 11 2
41 10 13 9 13 15 3 1 10 9 3 10 9 8 5 1 10 0 9 1 10 13 9 13 16 9 1 10 0 9 10 9 1 10 9 8 7 11 8 13 4 2
29 10 9 1 10 9 1 11 2 3 9 2 13 1 10 9 1 10 9 8 1 10 9 9 1 4 9 1 4 2
17 10 9 13 4 10 9 1 10 9 1 4 16 10 9 4 4 2
19 10 9 1 10 9 4 15 3 3 3 0 7 13 10 9 0 1 4 2
22 10 9 13 1 15 9 10 9 1 0 9 1 4 2 10 9 16 10 9 15 13 2
36 10 9 1 15 9 1 3 1 10 9 1 10 9 9 1 10 11 2 10 0 9 1 10 11 2 13 2 8 10 9 10 0 9 4 4 2
25 10 9 13 15 3 0 2 16 1 10 9 1 10 0 9 3 3 10 9 1 10 9 4 4 2
15 15 0 4 10 9 1 10 9 1 9 2 3 10 9 2
22 15 9 3 13 15 1 11 10 9 1 12 9 5 0 9 2 10 9 8 7 8 2
20 2 15 9 13 15 0 16 15 10 9 9 1 10 13 9 1 10 9 4 2
26 10 9 1 9 13 0 7 0 3 1 10 9 1 10 9 2 7 15 13 3 3 3 3 4 4 2
44 16 15 15 0 9 7 9 13 15 15 4 7 4 2 16 15 10 0 9 13 1 10 9 1 8 2 13 15 1 0 9 2 16 15 9 1 15 3 3 0 1 15 4 2
13 3 1 0 9 13 10 9 7 10 9 15 0 2
18 3 13 8 15 9 0 2 7 10 9 9 0 2 10 9 1 0 2
15 15 0 13 10 9 1 15 9 3 7 9 4 0 4 2
31 1 15 9 13 10 9 7 9 0 9 1 9 2 3 10 9 1 0 7 0 9 2 8 0 9 2 10 0 9 4 2
8 3 13 10 9 1 15 12 2
14 15 13 1 10 9 1 9 7 9 2 9 7 9 2
9 1 10 9 9 13 15 9 4 2
8 15 13 3 2 15 9 4 2
8 7 15 0 3 3 0 3 2
46 1 9 13 3 4 4 2 16 10 9 3 15 0 4 13 2 16 3 15 9 2 3 10 9 3 2 10 9 13 4 2 16 10 9 3 0 4 2 16 15 3 3 4 13 4 2
23 0 4 2 16 10 9 1 0 9 1 10 9 10 9 3 13 4 10 9 3 1 4 2
37 1 10 0 9 13 12 0 9 1 10 9 9 3 2 3 0 4 4 16 1 10 9 1 9 1 10 9 10 9 1 10 9 4 4 1 4 2
11 3 4 9 7 9 1 10 13 9 4 2
8 3 13 10 9 10 9 4 2
39 8 4 3 3 1 10 0 9 1 11 3 10 9 1 15 1 12 4 2 1 11 2 11 7 11 2 4 15 3 3 12 2 1 11 5 12 9 11 2
28 15 4 0 9 4 2 15 15 9 13 7 10 9 1 12 9 1 11 7 11 13 1 10 9 3 1 4 2
9 7 15 4 1 10 0 9 4 2
23 8 4 10 9 2 13 1 10 9 15 1 10 0 9 1 0 9 1 10 9 4 4 2
12 1 10 0 9 2 7 3 1 15 0 9 2
19 15 4 3 3 15 0 7 15 9 4 3 0 2 16 15 13 4 2 2
25 11 9 13 10 9 5 7 3 1 10 9 1 13 1 0 0 9 2 10 2 0 2 9 2 2
17 15 9 13 3 8 2 15 13 2 10 9 1 10 2 9 2 2
11 15 13 10 0 2 13 7 3 0 9 2
17 10 9 1 10 0 9 1 8 13 12 9 1 9 10 0 9 2
13 15 13 1 9 15 10 0 9 9 8 13 4 2
16 10 9 4 3 13 2 16 1 8 15 0 9 1 9 13 2
12 10 0 9 1 10 9 4 9 2 9 2 2
35 15 13 1 15 9 1 10 0 9 13 1 10 0 9 4 4 1 10 9 1 10 11 2 15 9 16 9 1 10 9 1 15 9 13 2
39 9 2 7 0 15 15 1 10 9 4 4 2 4 16 1 10 13 9 3 12 7 12 9 1 9 4 4 2 15 1 9 3 3 3 10 9 0 13 2
13 10 0 9 1 10 9 9 13 3 0 4 4 2
15 15 4 3 3 10 0 9 15 15 10 10 9 13 4 2
10 1 15 9 13 10 9 3 15 9 2
2 8 2
18 2 0 13 10 9 9 1 10 9 7 10 9 3 15 9 4 4 2
19 16 9 3 3 10 15 9 13 4 2 13 1 10 9 1 10 15 0 2
39 3 4 10 9 1 10 9 1 9 1 9 3 0 0 16 1 9 1 9 2 7 4 10 0 0 3 1 0 9 1 10 9 1 10 1 1 13 9 2
9 15 13 8 2 9 9 1 8 2
14 10 0 9 1 10 9 1 10 9 4 3 3 0 2
12 15 13 15 8 10 13 9 1 10 9 9 2
5 10 9 13 13 2
9 15 13 16 15 9 15 3 4 2
20 2 15 4 1 15 0 9 3 15 13 4 3 15 3 0 1 15 9 4 2
2 9 2
13 10 9 13 15 9 10 0 15 0 1 10 9 2
10 10 9 13 13 9 3 1 10 9 2
31 1 15 13 1 10 0 9 7 9 1 10 9 1 8 2 13 10 11 15 9 1 10 0 9 1 10 9 1 10 9 2
33 1 10 15 13 9 1 12 2 9 2 12 9 1 12 9 2 13 10 9 1 10 9 1 10 9 1 12 10 0 9 1 4 2
22 1 11 1 15 9 4 3 12 9 4 7 3 10 9 0 4 10 9 1 12 4 2
17 11 1 11 9 13 9 8 10 0 9 1 11 10 9 1 9 2
14 15 4 10 0 9 1 11 3 10 0 9 4 4 2
6 1 11 4 10 9 2
26 15 13 1 10 0 9 1 10 0 9 13 4 1 10 0 9 1 15 8 7 10 9 1 10 9 2
11 10 0 9 11 4 4 1 15 9 11 2
41 16 15 9 1 12 13 4 4 2 4 3 1 4 1 10 0 7 0 9 1 10 9 2 15 15 13 1 10 0 13 9 15 10 0 9 13 1 4 1 8 2
15 3 13 11 3 10 0 9 8 2 8 10 11 1 11 2
10 1 9 4 0 3 9 4 1 11 2
7 11 7 11 2 11 2 2
11 11 13 1 9 3 1 3 12 9 4 2
43 11 4 3 0 3 2 16 15 1 10 0 9 5 16 15 9 3 13 16 3 15 3 0 4 5 10 0 9 13 2 8 2 15 3 1 10 9 15 9 1 15 13 2
6 15 13 15 3 4 2
5 7 15 13 15 2
20 11 13 15 3 1 10 0 9 2 7 3 13 9 8 15 3 3 4 4 2
26 15 13 15 3 0 0 2 0 16 3 10 9 9 13 9 1 13 2 7 0 0 4 15 3 3 2
20 7 16 11 7 11 8 1 10 9 13 4 4 3 0 1 15 0 0 9 2
27 15 9 1 11 13 12 9 3 1 15 0 9 10 9 3 2 15 15 3 1 0 9 0 13 4 4 2
33 3 13 3 0 0 10 9 10 0 9 4 7 3 10 9 1 11 2 16 15 1 10 9 1 12 1 10 0 9 15 12 0 2
23 3 13 11 10 9 4 1 9 0 3 1 4 7 10 9 13 1 12 7 13 3 0 2
9 15 13 3 3 3 15 4 2 2
11 1 10 0 9 13 15 15 13 9 3 2
9 3 3 13 10 9 10 0 9 2
9 8 13 1 10 9 10 9 8 2
9 10 0 9 13 12 10 0 12 2
21 10 11 2 15 15 9 0 0 3 4 4 2 13 11 10 9 1 8 1 12 2
16 3 4 3 3 15 15 9 2 16 1 11 2 16 8 2 2
13 10 9 1 8 13 1 12 8 15 8 12 4 2
16 1 15 9 4 10 9 1 8 12 9 1 10 9 4 4 2
9 10 9 13 3 3 1 8 12 2
8 1 12 4 1 8 9 4 2
18 4 4 16 10 9 15 1 12 8 12 13 2 3 8 12 4 4 2
14 10 9 4 1 10 13 9 4 1 12 1 12 9 2
7 10 9 13 0 8 12 2
10 10 9 8 2 11 2 13 10 9 2
13 2 15 2 8 2 4 3 16 15 8 1 13 2
8 15 13 15 16 9 0 2 2
30 15 9 13 2 16 8 0 4 4 2 16 3 3 7 0 13 10 9 1 10 9 2 9 12 9 2 3 1 13 2
9 1 15 15 13 8 10 9 4 2
26 9 8 2 12 2 7 9 8 2 12 2 13 3 16 15 1 10 9 4 4 4 1 10 0 9 2
10 2 15 13 0 4 1 9 13 2 2
11 10 12 9 0 9 4 3 15 9 4 2
13 15 9 13 9 16 15 0 1 10 9 4 4 2
15 1 11 4 1 10 9 3 12 9 4 2 1 11 12 2
8 15 13 1 9 7 0 9 2
26 10 0 9 1 10 0 9 2 11 12 1 12 9 5 2 13 15 3 1 8 1 11 1 11 3 2
13 15 8 2 9 2 13 10 9 1 9 11 4 2
21 3 4 4 2 16 10 11 3 1 10 9 1 10 9 11 15 9 0 4 4 2
4 10 9 13 2
10 2 10 9 13 10 9 1 15 9 2
19 8 4 8 4 1 10 3 0 9 2 16 15 13 4 4 1 15 8 2
18 10 9 7 9 1 10 9 11 13 9 3 1 15 9 1 10 9 2
21 15 4 0 10 9 0 1 13 1 10 9 2 15 9 13 13 1 10 9 2 2
34 9 2 0 1 9 13 3 1 10 9 1 9 1 10 0 9 2 16 10 9 1 9 11 3 1 9 1 10 9 1 9 13 4 2
42 2 10 0 9 2 3 1 0 9 10 9 15 13 4 2 13 15 10 9 11 1 15 8 11 1 10 9 2 8 10 0 9 1 10 9 1 10 9 13 4 4 2
20 10 9 1 15 9 2 3 1 11 1 11 7 1 8 2 4 3 3 4 2
15 3 13 15 10 9 1 10 0 9 0 1 10 9 4 2
17 3 10 0 9 13 0 4 1 15 13 1 10 0 9 1 11 2
12 1 8 7 8 13 10 9 3 0 9 3 2
32 9 7 9 4 1 11 3 3 0 4 16 10 9 2 16 12 1 15 12 9 15 9 13 16 1 9 1 13 1 10 9 2
18 7 15 13 3 15 1 10 9 2 15 10 9 1 10 0 9 13 2
17 3 15 9 8 2 13 1 0 0 1 9 2 4 10 9 4 2
10 1 15 9 13 3 1 10 9 9 2
11 15 16 9 13 1 15 9 3 4 4 2
21 15 13 3 15 8 10 0 9 4 16 16 9 1 10 9 1 10 9 1 13 2
23 15 4 15 15 15 0 9 4 4 2 15 0 9 13 7 15 13 15 3 8 4 2 2
25 10 15 9 4 10 0 9 15 1 0 9 10 0 9 13 2 10 9 1 9 2 10 0 9 2
8 1 10 0 9 4 9 4 2
9 15 13 1 10 9 15 0 2 2
10 15 13 9 1 9 15 13 9 13 2
4 10 9 11 2
6 2 3 13 0 9 2
23 15 0 13 13 3 3 3 10 9 4 1 9 8 2 15 10 0 9 1 10 9 13 2
18 10 9 4 0 4 1 0 9 1 8 11 2 8 2 11 7 11 2
14 10 9 1 10 9 1 15 8 4 3 3 0 2 2
19 10 9 8 13 3 2 16 10 0 9 0 4 1 9 1 10 0 9 2
15 10 9 4 2 3 4 1 9 9 0 2 3 12 9 2
11 15 4 1 9 1 10 0 9 10 0 2
2 8 2
9 2 10 9 13 3 15 9 4 2
10 1 15 9 4 10 9 10 9 2 2
26 3 13 3 3 16 10 9 2 15 3 15 4 4 1 0 0 9 2 1 9 2 3 0 9 13 2
20 1 10 0 9 4 15 0 2 0 9 1 10 9 1 13 1 10 0 9 2
13 0 13 2 8 2 3 10 9 1 15 8 3 2
22 1 11 2 15 12 9 0 8 13 2 13 0 2 0 7 0 9 16 10 13 9 2
12 1 15 9 13 11 8 3 12 9 8 4 2
20 2 15 13 0 3 1 10 9 15 15 13 2 2 3 10 9 11 1 11 2
13 11 13 3 10 9 15 10 9 0 9 13 4 2
29 10 9 1 8 9 2 10 9 8 2 12 2 1 15 15 1 15 0 9 10 9 13 2 13 1 10 0 9 2
7 15 4 3 0 10 9 2
4 10 9 11 2
10 2 15 4 3 0 7 3 15 0 2
8 10 9 13 3 3 9 3 2
18 1 10 9 4 15 4 1 12 9 9 1 9 7 9 1 10 9 2
45 15 13 3 3 3 16 15 1 15 2 0 0 9 2 3 12 9 4 2 7 12 2 15 5 1 15 9 8 5 15 1 9 13 10 0 9 1 0 9 1 12 1 4 2 2
21 10 9 1 10 9 13 2 7 1 12 13 15 0 2 16 3 15 9 3 4 2
13 0 8 4 10 9 4 7 1 8 4 15 4 2
9 1 10 9 15 4 3 15 4 2
16 1 12 7 12 4 3 13 1 15 8 4 1 9 7 11 2
10 10 9 13 15 9 1 10 9 8 2
16 10 9 13 1 10 9 1 13 1 10 13 1 9 13 9 2
9 10 3 0 4 9 13 10 9 2
10 1 15 15 15 15 1 9 13 4 2
22 3 13 3 1 10 9 8 11 2 10 9 2 8 2 1 8 7 8 2 8 2 2
29 15 4 12 9 15 16 10 9 2 15 10 0 9 15 1 0 9 13 4 2 3 1 10 9 1 12 9 9 2
8 1 8 7 8 2 8 2 2
23 15 4 10 9 1 10 9 2 11 1 10 9 2 8 2 1 8 2 15 1 12 13 2
2 8 2
31 9 5 10 9 13 8 1 11 4 10 9 9 1 9 1 4 7 1 0 9 1 4 1 10 9 1 9 1 15 9 2
25 10 9 13 12 9 7 9 4 1 4 7 3 2 1 10 9 9 3 2 0 9 1 4 4 2
10 10 1 9 13 9 4 15 3 0 2
12 10 9 4 2 10 9 1 15 9 2 4 2
15 1 10 9 4 10 2 0 9 2 1 10 13 9 4 2
20 16 15 11 3 13 4 13 15 3 3 3 15 3 4 16 15 3 13 4 2
13 1 15 13 1 10 9 13 15 3 10 9 2 2
19 3 15 4 10 9 15 0 1 10 9 1 10 2 9 2 3 13 4 2
25 10 0 9 13 13 2 16 2 8 2 10 9 1 10 0 9 8 7 9 8 1 11 4 4 2
42 8 1 11 13 1 15 3 13 1 10 9 1 10 9 11 7 10 9 1 11 2 16 15 1 10 2 9 10 9 2 13 4 4 2 3 1 13 0 9 4 4 2
3 3 13 2
40 10 9 2 8 3 13 2 13 15 1 10 0 9 2 3 1 10 9 1 15 0 9 2 7 10 9 1 11 13 15 3 4 16 10 2 9 2 1 13 2
35 8 10 0 4 1 10 0 9 4 16 15 1 10 0 2 0 7 0 4 4 1 10 0 9 8 4 2 7 15 15 1 15 9 4 2
14 3 4 12 9 1 10 0 9 7 12 0 9 4 2
27 15 13 2 13 1 10 0 9 2 3 15 12 9 4 7 10 9 4 1 0 9 2 1 9 7 9 2
31 16 10 9 3 3 3 0 1 13 13 10 11 15 5 0 5 9 3 4 1 10 0 9 7 1 10 0 13 0 9 2
17 10 9 13 1 15 9 15 15 8 3 15 9 3 1 9 13 2
13 10 0 0 9 2 8 2 13 10 0 9 4 2
12 3 13 10 9 1 10 15 9 3 3 3 2
45 15 13 16 15 2 16 10 0 9 2 0 0 4 2 16 15 0 4 1 15 15 0 13 9 1 4 16 15 1 11 0 8 3 3 0 15 13 3 1 10 0 3 1 4 2
17 8 2 10 0 9 9 1 11 13 3 0 9 1 10 0 9 2
25 11 4 10 9 2 15 16 0 1 15 9 0 9 13 4 1 10 9 1 15 0 8 1 11 2
31 8 15 9 2 15 10 9 1 10 9 2 7 3 3 3 2 0 1 9 13 2 13 15 15 9 0 9 4 16 9 2
35 10 9 10 9 8 2 1 12 9 13 1 10 0 9 1 10 0 9 1 11 2 4 1 9 1 10 9 1 10 11 1 15 9 4 2
28 9 8 2 3 9 1 10 9 1 11 7 9 1 10 0 9 1 15 9 2 13 9 8 4 1 10 9 2
23 3 10 9 10 9 8 2 13 1 10 0 9 2 4 4 1 10 9 10 9 1 11 2
26 9 13 10 9 1 9 15 0 2 7 13 3 7 8 10 9 7 8 10 9 10 9 15 9 4 2
22 1 10 9 2 15 3 1 10 0 9 13 4 4 2 4 0 9 1 11 3 13 2
9 15 9 13 10 13 9 1 9 2
13 10 9 1 10 11 1 11 4 1 8 8 4 2
24 11 13 3 3 0 3 1 15 2 7 15 4 0 13 1 10 9 7 10 9 1 15 9 2
15 10 0 9 4 1 11 0 7 13 15 9 1 15 9 2
11 1 10 9 1 10 9 13 11 15 4 2
13 10 9 4 3 16 10 9 15 1 11 13 4 2
3 7 13 2
13 15 4 3 0 2 16 15 11 8 13 4 4 2
16 7 15 13 10 9 10 9 4 10 9 1 11 3 1 4 2
7 7 15 13 15 15 4 2
6 3 4 15 3 9 2
17 10 9 13 1 10 10 9 1 15 9 1 9 10 9 8 4 2
14 3 13 9 3 2 15 1 15 16 10 9 13 4 2
16 1 12 9 9 13 11 2 1 12 9 2 12 9 1 11 2
20 10 9 1 11 1 11 2 15 3 8 12 9 13 2 13 3 0 12 9 2
24 1 10 0 9 1 10 9 4 10 9 1 9 15 0 16 0 2 15 3 10 0 9 13 2
15 0 12 9 1 10 9 13 10 9 1 10 16 12 9 2
15 3 12 9 1 10 9 13 10 9 1 10 16 12 9 2
10 15 12 9 13 10 9 1 12 9 2
11 11 3 13 1 12 9 3 9 4 4 2
37 16 10 0 9 1 10 9 4 4 1 15 9 13 1 10 9 13 2 10 0 9 2 7 0 1 10 9 2 7 1 10 9 2 3 4 4 2
4 10 9 13 2
27 2 10 13 9 13 3 16 15 3 3 4 3 15 3 1 4 13 15 9 15 1 15 9 8 4 4 2
28 9 2 15 0 16 0 4 4 2 8 1 10 9 2 4 3 1 10 0 9 1 10 9 1 4 4 9 2
10 8 2 11 2 8 2 8 7 11 2
24 9 1 10 9 2 3 1 10 0 0 9 4 1 15 9 4 16 0 7 0 1 15 9 2
24 1 10 1 9 13 2 0 0 7 8 0 9 1 11 8 13 8 4 0 9 3 3 4 2
36 15 1 10 9 1 10 9 13 9 7 10 1 1 15 9 13 9 13 1 8 7 10 9 10 9 16 3 15 13 1 0 9 3 8 13 2
14 10 9 1 10 9 1 9 2 9 7 9 4 0 2
25 16 3 12 9 8 4 4 15 1 9 13 2 4 7 1 10 9 7 1 10 9 15 9 4 2
26 10 9 4 16 3 15 1 9 11 10 0 9 13 2 3 3 10 9 1 10 9 9 1 4 4 2
6 11 9 8 1 9 2
10 2 1 9 13 15 15 15 1 13 2
12 1 15 9 13 15 15 13 0 4 2 13 2
7 15 4 0 1 10 9 2
41 15 13 4 1 15 1 11 13 9 4 3 10 9 1 4 1 10 0 9 11 1 10 9 2 15 0 4 16 10 12 9 15 2 11 2 1 10 0 9 13 2
2 8 2
9 2 15 4 0 16 15 3 13 2
10 1 10 12 9 13 15 15 9 4 2
5 15 13 11 4 2
5 15 4 0 2 2
27 15 0 4 4 10 9 1 8 16 11 1 10 0 9 0 1 4 2 16 3 15 9 1 10 9 4 2
12 10 9 13 1 15 0 9 10 0 9 3 2
2 11 2
14 2 15 13 3 1 10 9 16 15 15 0 13 2 2
43 8 2 15 1 10 0 9 1 10 9 1 11 7 11 2 1 12 1 11 2 12 2 2 1 9 11 1 10 9 4 4 1 9 2 4 1 10 11 1 12 9 4 2
10 11 13 15 9 3 1 11 4 4 2
15 10 9 1 11 13 11 1 11 1 10 9 3 3 4 2
19 15 9 4 0 4 1 8 2 15 11 3 1 10 9 1 10 9 13 2
21 10 9 8 2 9 1 10 9 2 13 10 0 9 4 1 10 9 1 15 8 2
19 1 15 4 10 9 1 15 1 15 9 1 11 3 13 1 10 11 4 2
10 15 13 3 3 15 9 1 0 9 2
28 10 9 11 13 16 15 4 4 4 10 0 9 1 1 10 9 15 13 1 4 16 13 1 9 1 13 4 2
17 2 0 13 1 10 9 1 11 13 15 15 10 0 9 1 4 2
25 1 15 15 0 9 7 9 13 15 10 1 15 0 13 9 3 16 0 9 1 15 9 1 4 2
6 7 10 9 4 4 2
7 15 13 11 4 4 2 2
28 8 2 15 9 13 10 9 1 15 9 1 11 0 3 1 4 2 13 10 1 11 13 9 1 10 13 9 2
39 10 15 0 9 1 10 0 13 9 1 15 0 9 13 1 10 9 0 1 3 2 3 10 12 9 1 10 0 9 2 8 2 8 7 8 15 13 13 2
21 10 9 8 13 10 9 16 10 0 9 4 4 4 1 11 7 11 3 3 8 2
26 10 9 13 10 9 15 4 16 12 9 13 13 4 1 12 9 1 10 9 16 10 9 1 13 4 2
12 10 9 13 4 16 12 1 10 9 13 4 2
11 0 9 13 3 0 15 4 2 13 8 2
17 15 15 3 1 15 9 3 13 4 10 0 9 7 10 0 9 2
31 10 9 7 9 2 15 15 3 3 13 2 4 1 0 9 7 0 9 2 16 0 9 2 9 2 9 2 9 7 9 2
8 1 15 9 4 13 9 4 2
15 16 1 11 4 15 9 3 4 1 10 9 8 7 11 2
10 1 10 9 11 13 3 10 15 9 2
6 10 9 4 3 3 2
18 10 10 9 1 9 4 1 4 1 15 13 1 15 9 1 10 9 2
17 3 4 3 10 9 4 15 15 1 15 9 1 10 9 13 4 2
36 15 9 2 3 10 13 9 15 3 3 13 13 2 13 15 9 4 1 10 9 2 10 9 2 10 9 7 10 9 16 9 2 9 7 9 2
11 1 10 0 9 1 10 11 13 11 0 2
17 2 16 15 1 11 13 4 7 4 2 3 13 15 15 9 0 2
9 13 15 3 3 3 3 4 2 2
7 6 2 3 13 15 2 2
25 10 9 2 3 1 10 11 1 10 10 9 1 10 0 9 4 4 2 4 15 15 9 3 4 2
14 10 9 13 10 9 1 11 1 10 9 1 0 9 2
7 3 13 15 10 0 9 2
12 11 13 3 1 12 9 1 4 1 10 11 2
55 10 3 0 9 2 10 0 9 15 3 3 0 0 4 4 7 3 9 2 9 7 9 16 9 13 2 13 8 1 10 0 9 2 15 3 10 0 13 7 13 2 7 3 3 0 9 7 0 9 1 10 9 3 13 2
15 1 15 9 13 15 10 9 1 8 4 7 3 15 9 2
10 15 4 3 9 1 10 0 9 4 2
4 1 15 9 2
40 10 9 1 15 15 0 8 2 0 2 11 2 2 10 0 2 9 9 2 16 5 1 15 15 13 5 1 10 0 9 0 1 15 9 13 16 1 15 9 2
37 1 2 8 2 1 11 13 10 9 1 10 9 1 10 9 2 8 2 2 8 4 0 1 15 0 13 9 1 10 9 1 10 9 1 10 9 2
9 9 13 3 3 3 2 13 15 2
41 8 10 0 9 1 10 9 1 11 13 9 11 10 0 9 1 2 8 2 2 10 13 9 1 11 1 9 2 13 1 10 9 7 9 8 7 13 8 15 8 2
8 15 0 9 13 3 12 9 2
25 15 13 10 9 1 10 0 9 1 8 8 10 0 9 1 8 2 15 1 11 15 9 13 4 2
5 10 0 9 3 2
11 15 13 9 8 3 0 1 10 0 11 2
16 10 9 13 10 9 3 3 4 1 4 1 9 4 1 4 2
11 15 13 3 10 9 4 16 10 9 15 2
10 3 10 9 15 9 3 3 1 4 2
16 10 9 15 1 0 9 4 4 13 12 9 1 10 9 9 2
6 0 15 1 10 9 2
12 10 9 13 10 9 2 10 9 13 0 9 2
3 1 0 2
14 10 9 13 10 0 9 7 10 9 13 10 9 3 2
45 2 1 10 9 1 10 13 9 3 1 12 7 12 9 4 15 13 2 1 15 9 11 2 9 11 2 9 11 7 9 11 1 15 9 4 7 4 15 10 9 1 10 9 4 2
31 1 10 0 13 9 1 10 9 1 10 9 13 15 2 16 15 15 9 13 2 9 11 2 13 1 0 9 1 15 11 2
40 11 13 2 16 15 15 3 0 4 1 10 9 10 9 2 8 2 15 1 10 9 1 10 9 13 4 16 11 3 1 12 7 12 1 10 11 4 4 4 2
19 10 9 3 15 0 0 9 0 9 7 0 1 9 13 13 15 8 4 2
50 2 9 4 3 3 0 16 9 2 2 13 8 2 12 2 2 15 1 10 12 5 15 9 11 2 9 1 0 9 2 9 7 9 2 4 10 15 5 9 1 10 0 9 2 8 2 2 11 2 2
12 10 9 2 15 15 2 3 15 9 13 4 2
2 3 2
15 3 3 3 16 15 2 8 2 10 0 13 9 1 13 2
28 16 11 0 1 0 9 13 2 2 15 13 3 4 2 15 4 15 0 2 2 4 15 0 9 1 0 9 2
11 15 13 1 10 9 2 1 15 9 8 2
20 15 13 4 16 1 10 0 9 3 3 15 9 13 15 10 9 1 9 13 2
14 3 13 15 4 16 0 9 4 4 7 0 0 9 2
10 3 0 15 4 13 15 4 1 11 2
33 1 10 9 1 10 10 9 16 15 10 9 4 4 2 16 13 4 16 10 9 1 10 9 3 0 4 2 13 10 0 9 13 2
15 15 13 0 9 0 7 13 0 1 9 1 9 4 4 2
22 3 13 15 0 7 15 13 16 3 15 9 4 3 13 9 1 11 3 13 4 2 2
17 1 10 9 1 8 2 16 15 13 9 3 3 4 1 10 9 2
12 2 15 4 0 1 13 16 15 3 3 4 2
22 3 13 15 1 11 2 15 10 9 13 1 10 9 16 11 2 7 15 4 3 15 2
23 10 2 9 2 4 12 9 7 16 15 15 1 10 0 9 3 13 4 4 2 13 4 2
21 10 0 12 9 1 15 9 13 8 15 9 1 12 10 9 1 12 9 1 4 2
12 0 0 1 10 9 4 10 0 2 9 2 2
26 10 0 9 13 15 0 9 1 10 9 2 9 7 9 2 16 10 9 0 9 7 3 13 9 13 2
8 10 9 13 15 3 1 11 2
16 15 9 11 2 15 15 0 9 3 13 4 4 2 13 3 2
15 1 12 9 4 0 9 4 16 15 15 15 9 13 4 2
11 1 12 1 15 4 15 9 0 3 4 2
9 1 12 9 4 10 0 9 4 2
20 10 9 13 2 16 15 13 1 9 1 9 3 1 9 4 1 10 0 9 2
20 1 15 9 13 2 16 9 12 9 10 9 13 4 16 10 9 3 1 13 2
19 0 16 0 10 0 13 9 1 10 9 1 13 4 2 13 10 0 9 2
28 15 13 15 3 1 10 9 4 16 10 11 3 15 9 4 4 16 1 9 1 10 9 1 9 8 1 13 2
17 7 3 4 1 10 9 4 16 10 15 13 9 0 8 4 4 2
7 9 7 9 13 10 9 2
10 1 3 13 1 15 9 1 9 9 2
20 10 0 0 7 0 9 2 0 9 1 8 2 13 0 13 3 1 15 9 2
34 16 10 9 1 10 0 9 9 13 2 15 1 10 9 1 15 9 13 7 15 10 9 13 16 9 1 4 2 13 10 9 0 0 2
20 2 10 9 4 3 3 13 16 10 9 4 1 10 9 2 2 13 8 3 2
7 2 10 9 4 3 3 2
19 1 12 13 10 9 3 1 10 9 1 9 10 9 3 15 10 9 13 2
24 1 10 12 9 13 12 3 13 2 15 3 3 0 1 10 9 8 4 0 4 7 12 3 2
14 3 10 0 9 1 10 9 4 1 15 10 0 9 2
19 2 15 2 2 13 10 9 11 2 2 13 0 3 3 1 10 0 9 2
6 15 4 3 3 0 2
27 15 0 4 8 10 9 1 10 9 2 16 10 0 9 4 4 7 16 15 1 15 9 3 0 4 2 2
18 15 13 3 1 10 9 3 10 9 1 10 15 9 7 9 4 4 2
12 10 9 13 1 11 16 3 10 9 1 13 2
33 10 3 1 10 9 3 0 9 2 8 2 13 10 9 1 10 9 1 10 9 1 0 13 16 15 8 13 4 10 9 1 4 2
17 1 10 9 13 10 9 11 1 10 9 1 10 9 1 10 9 2
13 8 2 10 9 1 15 8 1 11 2 13 3 2
31 2 10 9 1 10 0 9 7 10 9 1 15 8 13 16 1 10 9 1 10 9 3 3 3 1 3 1 15 4 4 2
27 15 13 16 16 10 9 10 9 13 4 2 15 1 9 1 15 8 4 4 2 15 9 0 4 4 4 2
20 15 13 16 10 9 2 3 0 4 4 2 3 1 10 9 4 4 4 2 2
17 15 13 2 16 10 9 1 10 9 10 0 9 1 10 9 4 2
18 15 13 3 3 3 2 16 10 10 0 9 15 15 16 15 9 4 2
18 10 0 9 1 0 9 4 15 3 1 0 9 10 9 1 10 9 2
21 3 4 10 9 2 10 13 9 7 2 16 15 4 13 2 3 3 10 9 3 2
22 0 13 15 3 3 8 3 16 0 4 1 13 16 10 9 1 9 10 0 9 4 2
12 15 8 13 3 3 1 10 13 11 4 4 2
11 1 10 9 13 10 9 1 11 4 4 2
19 1 10 9 4 10 9 10 0 0 11 15 1 10 0 9 13 4 4 2
25 1 10 9 1 9 2 9 2 1 10 11 13 10 0 9 15 1 9 1 15 9 3 3 0 2
12 0 9 4 0 12 9 4 1 12 1 12 2
27 8 13 15 2 1 10 9 2 3 3 9 3 3 3 13 5 9 13 4 2 1 10 0 9 4 2 2
20 10 9 1 10 9 4 15 9 3 3 3 0 2 7 3 0 4 15 3 2
10 3 13 15 15 9 1 15 9 4 2
11 3 13 10 9 10 9 12 9 0 4 2
8 15 0 2 13 15 3 3 2
15 2 10 9 13 15 9 2 3 13 15 15 0 1 15 2
17 8 2 15 15 1 11 4 13 2 13 15 0 1 10 9 4 2
25 1 10 0 9 13 10 9 15 9 1 9 7 9 2 16 9 16 9 7 9 1 10 9 13 2
16 1 10 0 9 1 10 0 9 4 10 0 9 1 9 4 2
42 1 10 13 9 16 1 10 9 1 15 8 10 9 3 1 4 2 13 10 9 1 9 8 9 4 1 15 9 16 1 10 9 15 9 1 4 2 15 3 3 13 2
24 4 15 2 3 10 9 1 10 9 15 0 9 13 4 2 3 0 16 3 3 3 1 13 2
17 2 6 2 2 13 10 9 11 2 2 15 4 15 15 3 3 2
10 10 9 1 15 9 4 3 3 13 2
8 3 4 15 3 3 15 0 2
15 3 1 10 9 1 10 0 9 4 3 10 9 1 11 2
11 15 9 4 3 3 2 8 9 2 4 2
13 3 1 10 9 1 11 13 15 10 0 9 4 2
13 8 2 0 1 10 9 2 4 3 0 3 0 2
21 2 15 4 11 1 10 9 10 9 4 7 15 13 3 3 3 0 3 4 2 2
2 11 2
16 2 11 13 3 10 0 0 7 0 9 1 10 9 4 2 2
4 7 15 3 2
6 11 7 11 4 9 2
7 4 10 9 3 0 0 2
49 0 2 8 4 1 15 9 3 1 10 9 4 4 2 15 13 15 15 15 0 1 2 8 2 8 2 7 1 15 13 15 9 2 10 9 7 10 9 1 10 9 2 3 0 16 0 1 3 2
28 11 7 11 13 3 3 0 3 7 16 15 13 16 15 1 10 9 3 1 13 9 4 2 13 16 15 9 2
6 15 13 15 3 4 2
5 3 2 0 9 2
16 15 10 9 2 8 2 13 2 15 13 10 0 9 13 4 2
21 15 9 13 3 1 15 1 10 0 9 1 10 0 9 1 9 1 9 4 4 2
21 11 13 3 1 10 0 9 1 10 0 9 2 3 13 9 11 3 1 8 4 2
51 2 3 13 15 10 0 9 1 10 9 3 3 3 4 2 2 13 10 9 2 2 15 4 3 15 16 12 1 12 9 1 10 0 9 15 0 13 4 2 7 15 13 3 10 15 9 4 1 15 9 2
35 15 0 9 1 9 7 9 1 9 1 10 9 7 15 9 3 2 4 15 0 8 1 15 8 2 3 9 1 12 9 7 9 8 13 2
9 10 9 4 3 15 9 8 4 2
23 15 8 13 9 1 9 10 13 9 16 15 5 16 0 5 1 13 1 9 1 10 9 2
18 15 13 3 10 9 1 9 2 15 1 15 0 9 0 13 4 4 2
27 1 10 11 4 3 10 9 4 2 16 1 10 0 9 9 1 9 7 9 9 4 4 1 10 0 9 2
11 8 9 12 1 11 13 4 10 0 0 2
23 15 4 10 9 2 15 4 4 16 15 15 9 3 3 15 9 7 10 0 9 13 2 2
32 2 10 9 1 15 9 4 3 0 0 2 7 1 3 1 4 10 9 1 10 9 1 15 9 7 9 1 10 9 4 2 2
20 10 11 13 10 9 3 1 10 0 0 9 10 9 9 1 4 1 10 9 2
34 1 12 13 15 15 1 10 0 9 10 0 9 4 1 9 1 15 3 10 15 15 9 1 15 9 1 10 9 1 10 9 13 4 2
19 1 9 1 10 1 15 8 3 1 13 9 2 13 9 11 10 9 4 2
19 1 15 9 4 10 9 4 1 10 11 2 8 1 11 2 1 9 12 2
13 9 4 3 1 0 3 4 1 9 2 8 2 2
20 2 3 13 3 16 0 9 4 4 2 16 10 0 9 16 10 0 4 4 2
22 15 13 1 15 9 16 15 1 15 4 4 2 16 10 9 1 0 9 1 13 2 2
33 3 10 9 1 15 8 2 8 2 15 15 1 10 9 1 15 8 3 13 2 16 10 0 9 16 9 8 16 9 4 4 4 2
22 3 8 2 0 9 1 10 9 1 8 7 1 10 9 9 1 10 9 1 15 8 2
28 2 1 15 9 2 3 0 3 8 2 12 2 7 8 2 12 2 1 10 0 13 2 13 10 9 13 4 2
49 1 10 9 11 2 15 3 9 13 1 10 9 1 10 1 10 0 9 1 11 2 15 8 1 11 2 13 15 10 9 1 10 9 1 10 9 1 10 9 1 9 2 16 15 0 8 4 4 2
7 8 1 10 9 1 11 2
13 2 0 9 13 15 3 3 3 4 9 1 4 2
9 8 7 15 13 15 15 3 4 2
12 7 15 13 16 11 3 3 0 0 3 4 2
8 15 13 10 0 0 9 4 2
14 15 9 13 11 3 15 3 4 16 15 9 1 13 2
10 15 13 13 4 1 10 9 0 9 2
11 3 13 11 10 0 11 15 0 9 4 2
24 1 13 0 9 4 10 0 9 10 9 1 10 0 9 15 1 9 11 10 0 0 9 13 2
12 16 0 9 13 15 15 2 16 3 1 13 2
8 3 1 15 13 11 1 12 2
24 1 10 9 13 11 11 1 10 9 4 9 2 7 15 13 3 0 1 10 13 9 1 11 2
14 15 11 13 3 0 10 0 9 13 4 1 9 11 2
32 0 9 3 1 11 2 3 10 9 1 9 8 2 1 9 8 2 10 9 1 9 0 3 13 1 10 0 9 2 12 2 2
22 1 10 0 9 7 10 0 9 13 10 9 15 7 13 1 12 7 12 10 12 9 2
25 10 9 4 3 3 0 3 7 1 8 16 0 9 7 8 7 8 16 13 9 13 15 8 4 2
25 1 10 9 13 3 1 15 9 3 10 9 2 7 4 10 9 1 15 9 3 3 15 3 0 2
15 10 9 11 13 11 8 10 0 9 8 10 13 9 4 2
8 1 10 9 13 9 4 4 2
31 15 13 1 0 9 1 10 9 2 15 3 13 4 1 15 13 1 10 9 1 10 9 2 13 3 3 3 0 0 4 2
18 3 13 15 9 2 3 15 3 1 10 9 13 4 2 10 0 9 2
16 8 10 9 11 1 12 1 10 0 11 4 12 9 0 13 2
10 10 0 9 13 1 10 9 4 4 2
7 12 9 13 0 1 15 2
12 10 9 1 10 12 9 4 0 15 0 4 2
13 10 9 13 1 10 9 1 10 11 7 15 8 2
26 12 9 1 9 12 2 15 13 1 10 9 7 10 15 1 11 2 13 15 1 10 9 0 4 4 2
27 15 8 1 10 9 13 10 9 4 4 1 10 0 9 2 7 15 4 1 13 9 1 10 9 3 4 2
6 10 9 1 8 13 2
21 12 9 0 2 0 9 2 0 9 2 0 9 2 9 13 2 3 0 9 2 2
11 15 4 1 15 9 13 1 10 0 9 2
11 15 13 15 3 10 0 7 0 9 4 2
23 15 15 9 13 4 1 10 9 1 8 4 4 15 8 1 4 1 10 0 9 1 9 2
27 10 9 13 10 0 9 2 13 1 9 2 10 0 9 13 15 2 8 1 9 2 3 1 9 7 0 2
15 2 16 9 3 4 0 15 2 3 1 9 2 0 2 2
29 7 15 2 3 10 9 8 2 16 10 0 9 1 0 9 1 10 9 15 16 15 4 16 1 15 9 1 4 2
22 7 10 0 9 4 3 8 10 9 2 1 10 13 9 1 10 0 9 4 1 9 2
18 10 0 9 1 10 9 1 10 13 11 2 3 8 13 10 0 9 2
12 2 15 0 3 2 15 13 11 4 4 2 2
4 0 13 3 2
11 2 15 3 3 3 13 4 10 11 2 2
9 10 9 4 3 15 3 3 1 2
15 3 13 15 0 4 16 15 1 10 0 9 1 13 4 2
10 2 7 15 13 11 3 3 4 2 2
22 11 2 10 0 9 1 15 8 2 1 12 2 2 13 3 1 10 0 9 1 8 2
54 1 10 11 13 0 9 1 10 11 13 10 9 8 2 9 1 15 8 7 0 9 1 15 8 2 4 1 10 9 1 10 9 1 13 0 9 2 3 10 9 10 9 13 1 4 1 15 1 13 13 1 10 9 2
30 10 9 8 13 2 16 10 0 9 1 9 8 4 1 10 0 9 1 10 0 9 7 15 13 15 0 1 10 9 2
17 2 11 13 3 0 4 4 4 2 7 0 0 4 15 15 3 2
10 15 13 15 4 16 10 9 8 4 2
23 3 2 16 15 10 9 1 15 0 12 9 0 13 4 4 2 3 13 15 15 3 4 2
11 7 15 0 12 9 13 15 3 3 15 2
20 16 11 3 3 0 13 13 15 0 3 16 3 3 15 3 1 4 4 2 2
19 0 13 4 1 15 2 8 2 1 8 7 3 1 15 12 9 9 4 2
5 15 13 15 4 2
15 15 4 10 9 3 4 1 10 9 1 10 9 1 13 2
20 1 10 13 9 13 15 10 9 0 2 3 9 7 15 9 0 13 1 4 2
20 1 10 0 9 4 10 0 9 4 1 10 9 1 10 9 2 10 9 8 2
11 10 9 2 10 9 7 10 9 4 4 2
32 7 15 4 0 16 10 9 1 15 9 0 4 4 2 3 16 15 10 9 13 4 1 15 1 3 10 13 7 10 0 9 2
23 8 10 9 1 15 0 9 0 7 15 0 13 1 10 9 1 10 12 9 9 10 9 2
25 1 10 9 13 15 10 2 13 2 9 3 16 10 9 8 10 9 1 15 0 0 9 0 4 2
21 0 13 15 3 9 1 10 0 9 7 9 2 15 15 9 1 10 0 9 13 2
23 15 9 9 13 15 1 10 9 2 16 15 10 0 9 1 10 9 1 2 8 2 13 2
40 10 0 0 9 2 15 1 12 1 10 9 1 8 15 9 13 2 4 15 3 1 10 0 9 1 4 4 2 16 15 0 1 15 9 10 9 13 4 4 2
17 7 0 3 13 15 0 9 13 9 3 3 1 0 9 4 4 2
19 10 8 4 9 1 10 9 1 11 7 11 13 0 9 1 0 9 3 2
25 10 3 0 9 4 10 12 9 1 11 7 11 1 12 7 10 12 9 1 11 7 11 1 12 2
21 10 0 9 13 11 1 12 7 10 0 9 11 13 1 12 1 11 15 15 4 2
15 10 0 9 1 10 9 4 1 12 1 11 7 8 4 2
18 10 9 11 13 16 10 9 1 10 9 1 0 9 10 0 9 4 2
14 3 8 0 9 15 3 1 15 0 9 0 0 13 2
30 10 9 1 10 9 16 9 4 3 4 1 10 0 9 8 9 2 15 10 9 1 10 9 4 2 3 10 9 11 2
14 2 10 9 4 1 15 9 3 7 3 15 0 2 2
8 8 13 8 1 10 0 9 2
16 11 7 11 13 15 8 2 11 8 2 8 8 7 11 3 2
24 15 0 3 12 9 0 8 2 13 3 15 0 9 4 2 1 1 15 10 0 0 9 11 2
9 1 8 4 3 12 9 0 4 2
11 8 13 8 2 8 12 7 11 12 9 2
9 8 7 11 13 15 12 9 9 2
8 8 13 12 7 8 12 9 2
26 2 3 13 15 10 9 1 10 9 15 4 4 2 7 4 4 7 10 9 3 1 10 9 4 4 2
10 15 13 1 10 9 4 1 0 9 2
13 15 13 3 3 10 9 4 3 10 9 1 4 2
26 6 2 3 13 10 9 11 2 2 15 1 11 13 15 10 9 1 10 9 13 2 3 3 15 4 2
24 9 11 13 3 1 10 9 1 15 9 10 9 2 10 0 0 9 2 3 16 10 9 8 2
17 2 10 9 2 15 4 10 9 1 10 9 2 2 13 9 11 2
4 15 0 9 2
13 0 13 15 16 11 10 9 1 15 8 4 4 2
24 2 15 13 15 3 8 10 9 1 9 1 15 9 4 2 2 13 10 0 9 15 9 3 2
33 10 9 13 15 9 3 3 7 16 1 10 13 9 3 3 15 7 15 13 13 2 13 3 1 0 9 1 15 3 9 4 4 2
21 15 13 3 3 4 7 3 9 4 1 10 0 0 9 2 15 13 15 15 4 2
30 3 13 3 3 16 11 3 10 9 13 1 10 9 15 15 9 1 10 9 15 4 16 10 9 1 10 9 1 4 2
41 1 10 0 9 13 10 0 9 8 7 8 15 3 1 10 9 9 1 9 11 1 10 13 9 1 10 13 9 3 1 4 16 1 10 9 1 8 9 4 4 2
26 0 9 1 10 9 4 3 1 12 13 1 10 0 9 2 3 13 15 0 9 15 1 4 4 4 2
12 7 10 13 9 13 15 9 1 10 0 9 2
32 1 10 9 1 10 0 9 4 15 0 3 0 16 10 9 1 10 0 9 11 7 10 9 1 11 1 10 0 9 1 11 2
50 10 9 3 11 3 13 4 3 10 9 1 10 9 1 12 9 16 15 0 9 3 1 4 1 10 9 1 10 9 2 3 10 9 3 13 2 7 3 16 3 9 1 13 1 10 9 1 10 9 2
12 10 0 9 13 11 2 8 2 3 9 4 2
14 10 0 2 0 9 2 1 15 10 9 10 0 4 2
12 7 3 10 9 15 1 10 0 13 9 13 2
15 10 0 0 9 13 0 10 9 1 9 8 2 4 2 2
13 10 9 13 8 8 1 10 9 1 9 0 4 2
17 10 9 13 15 9 4 16 10 9 1 2 0 9 2 13 4 2
26 3 13 2 13 15 2 3 9 4 7 3 13 15 1 4 16 10 9 1 10 9 0 3 0 4 2
10 10 9 1 10 9 4 15 9 3 2
36 15 13 15 4 1 9 1 10 9 0 13 9 2 3 13 8 1 15 9 1 10 3 13 0 9 12 1 10 0 9 1 9 1 0 9 2
20 8 13 15 3 3 10 9 15 1 10 1 15 13 9 4 4 1 10 9 2
14 10 0 9 7 3 10 9 13 15 3 3 4 4 2
40 9 8 2 11 11 2 13 3 1 10 9 1 10 11 15 3 3 0 1 4 16 15 3 3 0 1 4 1 10 9 3 10 0 9 1 10 9 4 4 2
22 8 13 15 10 0 9 1 10 0 9 4 2 16 15 0 9 1 11 13 4 4 2
18 15 13 3 3 3 3 1 10 0 13 9 16 3 1 9 4 4 2
27 3 16 10 9 1 15 13 1 10 9 4 13 4 2 13 15 9 4 1 10 9 2 3 13 9 8 2
26 10 11 13 2 16 15 10 0 9 1 11 7 11 4 4 2 3 10 9 2 8 2 1 8 4 2
18 11 13 1 9 1 10 9 1 11 15 3 8 1 15 8 4 4 2
17 3 4 15 10 9 1 11 16 15 9 1 10 0 9 1 13 2
26 10 9 15 3 9 13 1 15 9 2 8 2 2 3 1 10 11 13 2 13 10 0 15 9 4 2
22 8 13 1 15 9 1 10 9 16 10 9 1 15 9 0 1 4 1 10 0 9 2
41 0 4 3 3 4 2 16 15 9 3 8 4 4 4 1 9 1 9 2 9 7 0 9 2 16 3 3 15 9 1 9 4 13 4 1 15 13 1 15 9 2
8 10 9 4 3 3 2 8 2
10 15 13 16 15 9 0 7 0 4 2
7 15 15 1 15 9 13 2
5 15 13 15 9 2
7 15 9 13 1 10 9 2
10 15 13 1 10 0 7 1 10 9 2
16 15 13 3 15 0 9 7 10 9 4 7 13 15 3 4 2
18 15 13 10 9 1 10 9 1 4 7 3 4 15 1 10 9 4 2
9 15 4 15 10 0 9 4 2 2
22 10 9 1 10 0 9 13 10 9 0 4 4 7 15 13 3 10 9 4 4 2 2
24 1 15 1 15 9 13 9 13 10 11 3 1 0 9 15 9 4 1 10 9 1 15 8 2
11 3 13 9 8 10 9 1 15 9 4 2
27 2 9 13 9 4 2 2 3 10 9 2 7 16 11 11 13 2 13 15 15 16 15 9 1 13 2 2
10 15 13 15 1 15 12 9 7 9 2
23 0 2 3 10 9 15 15 1 10 0 9 1 11 4 4 2 13 15 3 3 15 2 2
51 7 3 11 13 15 16 10 9 1 10 9 1 11 13 4 2 10 9 0 1 4 4 2 10 9 1 10 0 9 3 1 4 4 7 10 0 9 1 10 0 9 13 4 1 15 8 7 10 0 9 2
18 3 13 10 0 9 3 3 15 9 3 4 11 10 9 3 1 4 2
42 10 0 9 13 10 0 9 8 4 1 12 9 9 1 9 1 10 9 1 9 1 10 9 1 10 11 2 16 15 1 12 10 0 8 15 9 1 10 9 13 4 2
14 10 9 4 1 10 9 9 1 9 7 0 9 4 2
10 3 13 12 9 1 9 1 11 4 2
14 8 10 3 0 9 1 10 9 4 10 0 9 0 2
12 8 13 3 10 9 3 4 12 2 12 2 2
23 10 0 9 1 11 2 13 1 10 9 2 13 0 3 9 4 1 10 0 9 1 8 2
14 4 13 4 16 15 9 1 10 3 0 9 3 4 2
14 15 9 4 3 0 7 13 3 1 15 10 9 4 2
19 11 13 0 1 12 7 0 3 13 10 0 9 3 1 12 2 12 2 2
28 3 3 13 15 3 1 11 1 0 9 8 1 10 0 9 1 9 1 12 9 1 11 7 12 9 1 11 2
16 10 9 3 4 10 9 1 10 11 1 10 9 1 12 9 2
25 15 4 1 10 0 9 15 13 15 9 4 1 9 1 10 9 1 10 9 7 15 4 13 0 2
8 15 13 8 3 1 10 9 2
11 15 13 16 1 10 9 10 9 4 4 2
30 10 9 1 10 13 0 13 3 3 3 3 16 15 15 9 4 2 7 3 1 10 9 16 15 3 3 13 0 4 2
15 10 9 1 9 13 10 9 1 10 9 1 10 9 3 2
9 1 12 13 10 9 1 10 9 2
17 10 9 13 3 4 1 10 0 0 9 7 3 10 9 1 9 2
15 15 4 1 12 9 1 9 4 7 4 3 1 10 9 2
39 10 9 1 9 1 10 9 1 11 2 8 2 13 1 10 0 9 8 1 11 12 9 12 9 9 1 9 4 1 12 9 1 12 9 1 11 7 9 2
24 10 9 0 1 11 0 12 9 1 9 1 11 2 11 7 11 3 15 3 8 13 4 4 2
16 1 9 3 3 1 10 9 1 4 4 15 1 11 8 4 2
16 1 9 1 15 8 4 10 9 11 4 1 10 9 1 9 2
35 10 11 13 15 8 4 7 9 1 15 7 15 9 4 3 3 4 11 13 3 1 10 0 9 3 3 1 11 4 16 1 13 1 11 2
22 16 10 9 10 0 9 1 15 13 4 13 15 1 10 9 3 16 0 9 4 4 2
14 7 15 4 3 3 15 2 3 15 15 9 4 4 2
35 15 9 4 15 2 3 3 3 0 13 1 10 9 2 3 10 9 16 15 0 0 2 7 3 15 0 2 8 0 3 3 3 0 13 2
15 15 9 13 3 4 4 1 9 1 10 9 0 9 11 2
11 0 8 10 0 9 13 11 15 1 4 2
14 10 9 15 4 4 1 0 0 9 2 15 0 13 2
26 1 10 0 9 2 13 1 9 16 10 0 9 1 9 13 2 4 4 10 9 1 15 9 1 4 2
4 9 11 3 2
8 2 15 0 9 13 15 0 2
6 15 13 15 0 13 2
13 0 0 2 7 1 15 9 13 15 0 0 2 2
3 7 8 2
17 2 1 15 9 13 15 10 9 2 16 8 4 3 1 4 4 2
29 3 10 9 3 4 4 13 8 16 15 10 9 4 16 10 0 9 10 9 7 0 8 3 1 10 9 4 4 2
29 10 9 4 4 1 10 9 2 15 10 9 0 3 13 4 2 7 15 4 1 10 9 3 16 10 0 9 4 2
30 16 15 12 9 3 1 0 9 1 13 13 15 1 10 9 8 4 4 7 8 13 15 3 15 10 0 9 1 4 2
10 15 13 15 10 9 1 9 4 4 2
5 15 13 11 3 2
15 10 0 11 13 10 9 1 10 9 3 3 2 4 15 2
21 1 10 0 9 1 10 0 9 2 11 2 8 7 8 13 3 3 0 9 2 2
22 3 3 13 11 1 15 1 15 13 9 2 7 8 2 10 0 0 11 2 13 0 2
9 11 13 3 0 1 10 0 9 2
11 7 3 13 11 15 0 9 1 10 9 2
18 9 1 9 13 10 7 0 9 16 9 15 15 9 1 10 9 4 2
33 1 15 9 4 10 9 9 7 9 1 10 0 9 4 2 1 10 9 2 15 1 10 9 12 4 4 1 10 0 9 1 9 2
27 10 9 4 4 1 10 9 1 12 0 9 1 10 9 2 10 9 15 1 10 9 0 0 4 13 4 2
28 10 9 13 3 0 10 9 0 3 4 4 7 15 3 0 13 1 15 9 1 15 13 4 3 15 13 4 2
10 7 9 16 0 4 10 9 0 11 2
29 15 10 0 13 2 13 10 9 4 4 1 8 2 15 10 0 9 1 10 9 7 10 9 8 3 4 1 4 2
10 1 15 0 9 4 10 9 10 0 2
12 11 13 8 12 1 15 9 1 15 8 4 2
22 15 13 9 1 10 9 1 3 8 12 2 15 1 10 9 1 10 0 9 13 4 2
23 10 9 13 3 1 15 15 11 1 10 9 1 10 11 0 13 4 1 9 1 15 9 2
23 1 15 13 1 10 9 4 1 10 9 15 0 9 0 7 10 9 13 3 1 4 4 2
19 10 9 1 15 0 7 0 9 13 15 1 12 1 10 13 9 0 4 2
23 10 0 9 2 15 1 15 9 13 2 7 3 3 1 10 9 1 10 9 13 2 4 2
16 15 13 15 0 9 1 12 9 7 15 9 9 13 9 4 2
32 9 13 4 2 15 8 10 9 2 15 1 10 0 9 3 13 4 4 2 1 12 1 12 9 2 12 1 9 2 3 4 2
13 10 9 0 2 0 2 0 7 0 4 0 4 2
36 11 9 1 8 2 10 9 11 2 4 1 9 0 9 9 1 10 9 2 15 13 3 10 9 2 10 9 2 3 15 0 3 12 9 13 2
19 15 9 2 15 15 9 13 7 10 9 12 13 2 13 15 3 16 9 2
11 3 15 13 3 3 3 15 1 9 3 2
28 15 9 1 10 11 13 15 8 13 9 1 10 9 1 15 8 2 10 0 9 2 10 9 1 9 7 9 2
11 1 10 9 1 10 11 13 3 3 9 2
18 0 13 12 9 1 15 4 2 16 16 10 15 10 15 15 13 4 2
9 0 9 7 9 13 0 10 9 2
48 3 1 10 9 4 0 3 4 1 0 9 16 9 16 1 10 9 1 4 2 7 1 10 2 9 1 11 2 13 10 9 15 3 4 2 16 3 10 9 4 13 4 15 1 12 9 13 2
21 15 13 16 15 3 4 7 3 0 4 3 15 13 1 9 1 10 9 4 4 2
26 7 3 4 3 10 9 3 15 15 9 7 15 13 16 15 3 1 10 0 9 3 10 9 4 4 2
10 15 9 13 15 15 3 1 9 4 2
7 10 9 13 10 0 9 2
5 11 13 15 2 2
43 1 15 9 13 9 3 9 3 0 3 8 1 4 2 7 2 15 13 15 0 2 15 4 3 10 9 2 15 13 10 0 9 3 15 3 13 4 4 3 15 4 2 2
22 15 13 1 10 0 9 1 10 9 1 8 1 11 1 15 9 13 3 15 9 4 2
9 10 9 1 9 8 11 13 0 2
40 11 13 15 1 10 9 4 4 1 10 9 1 9 2 15 13 9 7 9 4 4 7 15 1 10 9 1 10 0 2 11 2 3 0 4 4 1 0 9 2
23 2 8 2 1 8 4 10 0 2 6 2 15 4 10 9 3 2 13 9 1 0 9 2
10 13 2 3 3 1 10 0 0 9 2
2 13 2
3 12 9 2
22 16 1 13 2 8 2 16 0 13 1 8 7 15 0 10 0 9 1 15 9 13 2
19 9 8 13 10 9 3 1 4 1 10 0 9 7 9 8 2 11 2 2
7 15 13 3 3 15 3 2
2 3 2
43 2 8 2 2 10 0 9 1 10 9 15 10 9 1 10 9 9 2 13 1 10 9 2 13 1 15 9 2 16 15 0 15 9 1 15 13 2 5 7 15 13 15 2
7 1 10 9 4 12 4 2
5 10 9 13 0 2
22 11 13 0 9 3 1 12 4 4 2 16 0 0 3 1 13 1 12 2 12 2 2
12 3 13 1 15 9 3 9 9 1 0 9 2
27 1 10 9 4 3 10 0 9 11 1 12 1 4 4 3 15 9 1 10 0 9 3 13 1 4 4 2
6 11 4 0 1 9 2
22 3 13 3 10 9 1 10 11 7 1 11 15 15 12 1 12 9 1 15 9 4 2
35 15 13 1 10 9 1 11 9 4 1 13 9 1 10 9 8 8 9 1 10 9 1 10 9 1 10 9 15 1 12 1 10 9 13 2
14 0 4 1 10 9 1 11 7 11 15 12 9 4 2
7 3 3 12 3 1 11 2
14 1 10 0 9 13 3 12 9 15 9 1 10 11 2
20 10 9 3 2 3 1 11 2 1 15 9 3 12 9 3 10 0 9 13 2
28 9 7 9 1 15 8 4 15 3 1 9 0 4 1 10 0 9 1 9 1 10 13 9 1 10 0 9 2
8 10 0 9 3 4 3 0 2
12 10 0 2 2 0 2 9 1 10 9 2 2
7 10 9 7 9 1 12 2
32 10 9 1 10 9 13 9 11 0 15 9 1 12 1 12 9 1 4 7 15 9 2 1 10 9 2 3 1 4 1 12 2
16 0 13 15 10 9 4 4 1 10 9 1 8 1 15 9 2
18 8 13 10 9 1 9 1 8 0 7 13 2 16 0 9 8 4 2
33 1 1 0 4 15 3 3 3 16 3 1 11 15 9 1 10 12 9 13 2 15 10 9 1 15 9 3 1 10 9 13 4 2
5 13 15 3 3 2
8 11 2 11 2 11 2 11 2
16 1 15 0 9 13 15 3 3 15 15 3 1 15 9 4 2
16 15 4 10 0 9 9 2 10 9 2 15 1 15 8 13 2
7 1 10 9 4 15 4 2
11 3 1 10 9 2 15 15 1 9 13 2
11 0 4 10 9 10 9 1 10 0 9 2
11 15 4 3 10 9 9 3 1 9 4 2
28 16 15 1 10 0 9 2 15 0 1 9 4 13 2 10 9 4 2 4 3 1 15 9 10 9 0 4 2
31 10 12 9 1 10 9 13 3 1 11 3 13 7 13 2 1 10 9 4 3 1 4 4 4 1 10 9 1 0 9 2
21 10 0 9 12 10 0 9 15 10 1 8 13 0 9 13 4 2 1 0 9 2
17 1 10 9 1 10 11 9 9 8 7 9 11 3 10 9 3 2
16 5 10 13 9 4 4 1 10 9 3 10 9 1 9 13 2
28 5 8 13 15 9 4 16 10 0 9 1 10 0 9 4 4 1 10 0 9 15 1 12 13 4 4 4 2
15 3 4 15 12 9 3 16 10 0 0 0 9 4 4 2
15 15 9 4 0 4 1 10 9 1 10 9 1 10 9 2
18 10 0 13 9 3 4 1 4 1 10 0 9 11 2 9 2 8 2
24 15 13 15 9 1 10 9 1 10 9 2 10 9 1 10 0 9 15 1 10 9 3 13 2
12 1 15 9 13 1 10 9 3 10 9 4 2
10 15 4 10 9 1 10 9 1 8 2
31 10 9 13 0 10 9 1 10 9 9 7 1 15 9 9 4 16 9 0 1 13 16 15 9 15 0 9 1 13 4 2
14 10 13 9 1 3 12 9 1 10 9 1 12 9 2
9 5 0 9 7 9 1 10 9 2
11 5 0 9 7 9 1 9 1 0 9 2
23 5 10 9 1 9 2 9 7 0 9 13 10 9 4 1 10 9 8 10 9 1 9 2
10 3 13 15 12 9 3 3 9 4 2
8 3 13 15 3 15 3 3 2
9 10 9 1 10 9 13 15 0 2
19 2 10 9 2 15 3 4 4 4 3 15 1 10 9 2 2 13 8 2
20 15 13 3 0 10 9 3 2 16 15 13 3 15 1 15 9 1 4 4 2
14 7 10 12 9 13 3 0 4 16 15 9 0 4 2
15 15 13 3 3 2 16 10 9 1 11 3 4 4 4 2
7 0 13 15 3 9 4 2
27 15 13 15 3 3 2 7 15 13 3 3 10 9 0 16 15 2 9 2 1 10 0 9 3 1 4 2
12 13 15 15 9 3 1 9 9 3 1 13 2
12 1 11 5 3 0 0 5 9 8 13 8 2
14 2 15 0 9 4 3 16 15 3 0 3 13 4 2
9 15 13 3 3 9 9 0 4 2
4 10 9 9 2
7 15 13 10 9 3 4 2
13 15 4 13 15 3 10 0 9 1 9 11 2 2
8 15 13 10 2 0 9 2 2
22 10 9 1 10 0 9 16 3 1 4 13 8 2 12 9 3 12 9 2 3 3 2
5 2 6 2 6 2
32 1 10 0 9 4 3 10 9 4 16 12 9 3 12 13 2 3 0 0 9 2 1 10 11 1 10 9 1 9 4 4 2
13 10 9 1 15 15 1 10 9 13 4 13 3 2
19 10 0 9 2 8 2 15 10 9 9 3 8 15 9 4 4 4 4 2
21 10 9 1 10 11 1 10 9 1 9 1 11 13 1 8 1 10 3 0 9 2
22 8 13 1 10 1 12 1 13 0 9 10 9 1 10 9 1 10 9 1 9 4 2
8 15 13 3 10 9 1 8 2
29 10 9 11 13 2 16 13 2 8 2 15 4 4 1 9 1 10 9 1 9 10 0 9 1 10 0 9 4 2
20 10 9 8 13 8 3 2 15 15 9 13 4 1 15 13 1 10 0 9 2
34 15 13 3 4 16 15 1 10 9 8 9 1 10 11 5 8 11 2 11 2 11 7 11 5 1 10 9 1 10 0 9 4 4 2
51 10 9 1 15 0 8 13 9 11 7 9 11 2 10 9 4 2 3 15 9 2 15 1 0 9 10 9 4 4 1 10 9 1 11 8 15 2 15 1 15 1 10 12 13 9 13 1 10 0 9 2
24 16 1 12 15 9 4 4 2 13 10 9 5 16 15 10 9 13 5 10 9 1 10 9 2
8 3 10 9 4 3 3 13 2
26 16 10 9 10 9 1 15 15 9 9 1 11 13 4 10 9 1 15 13 3 3 1 10 9 4 2
14 11 13 15 9 1 12 9 1 15 7 15 9 11 2
30 10 11 13 1 11 0 9 10 13 7 0 9 4 15 10 13 9 13 16 10 13 9 1 10 9 9 3 1 13 2
11 15 4 10 9 15 8 0 4 13 4 2
34 10 11 13 10 9 1 10 9 1 13 7 0 9 5 7 3 0 10 2 13 9 2 5 16 0 9 1 10 9 3 0 1 4 2
22 10 11 13 3 9 1 15 1 0 9 3 3 4 1 4 1 13 9 8 0 9 2
10 15 13 1 0 9 1 10 13 9 2
19 0 12 9 1 10 9 12 0 9 13 3 10 9 1 15 0 9 3 2
17 7 3 13 3 3 10 9 4 4 16 3 3 0 4 4 4 2
14 10 13 13 9 13 1 15 9 10 3 0 9 4 2
10 7 15 9 4 3 1 12 9 4 2
10 10 0 9 7 10 9 1 15 9 2
12 10 0 9 13 1 15 0 9 4 1 4 2
21 1 0 11 13 10 9 4 2 15 1 15 9 1 3 1 3 1 15 9 13 2
16 2 7 3 10 0 9 11 13 1 9 2 2 13 10 9 2
24 1 9 1 12 7 12 9 13 10 0 9 3 0 0 16 11 9 3 3 3 15 9 4 2
36 10 9 9 1 15 10 9 3 16 1 9 1 4 16 10 9 15 1 9 13 4 4 1 2 0 9 2 1 10 2 11 10 0 9 2 2
17 10 11 13 15 9 4 16 10 9 9 10 3 0 9 1 13 2
9 15 13 7 13 10 0 9 4 2
16 8 2 8 7 8 2 1 11 9 1 9 2 13 10 9 2
26 1 1 15 9 13 16 16 15 8 3 1 9 7 3 1 10 9 4 4 10 9 10 9 13 4 2
9 10 9 13 3 0 3 3 4 2
17 1 15 0 8 4 15 0 16 10 9 16 10 13 9 13 4 2
10 9 8 4 1 9 4 16 9 8 2
26 15 0 8 5 2 1 12 9 1 10 9 1 11 2 2 9 7 9 2 9 2 13 10 9 4 2
2 8 2
18 3 3 1 10 9 1 15 0 9 2 8 9 2 4 15 9 4 2
9 10 9 1 11 13 0 0 4 2
38 15 4 3 0 10 9 1 10 9 3 1 13 2 16 1 12 9 7 9 2 15 3 16 9 13 3 1 4 2 9 7 9 8 10 9 8 13 2
7 1 9 4 10 9 9 2
10 11 2 12 2 8 4 0 0 9 2
2 12 2
12 1 10 9 13 10 9 1 0 9 10 9 2
9 1 12 13 15 10 9 1 12 2
7 9 8 2 9 1 11 2
13 2 10 9 4 3 10 9 1 9 1 15 9 2
19 1 10 13 9 13 15 3 15 8 7 15 13 3 10 13 9 1 4 2
6 15 13 3 1 13 2
15 2 15 13 2 16 0 3 1 10 9 10 9 0 4 2
18 3 13 15 8 10 9 12 9 7 3 13 10 9 3 3 1 15 2
11 15 13 3 1 10 15 13 9 1 11 2
9 11 4 1 9 3 10 0 9 2
13 0 9 13 15 15 0 9 10 0 0 9 4 2
4 15 13 4 2
18 16 3 3 10 0 9 1 10 9 4 4 2 13 3 10 9 3 2
12 10 9 4 4 2 15 13 10 9 8 4 2
11 10 9 1 10 11 13 15 9 9 4 2
20 10 9 13 15 9 15 1 12 9 13 4 2 1 10 9 1 10 9 4 2
9 3 13 15 3 3 10 9 4 2
10 10 9 13 3 10 0 10 9 4 2
22 1 10 0 13 5 16 16 3 9 4 4 5 4 4 15 1 10 9 3 1 4 2
38 10 9 2 15 1 15 9 10 9 13 1 10 0 2 0 9 1 15 9 2 15 13 4 2 16 15 3 0 7 1 9 4 2 4 8 1 11 2
7 8 13 7 9 16 9 2
18 3 4 15 0 9 2 2 8 2 1 8 1 11 1 10 9 4 2
43 1 10 9 8 1 10 0 9 2 15 0 4 4 1 10 9 1 10 9 1 9 2 13 3 10 9 1 9 7 9 1 10 0 9 1 11 10 0 9 0 9 3 2
29 1 12 9 13 10 9 3 12 9 1 9 4 1 0 9 15 0 2 8 2 5 3 9 7 9 5 4 13 2
20 1 12 4 3 12 0 9 4 2 1 10 13 9 13 15 9 3 1 12 2
43 10 12 2 9 2 2 15 8 1 11 2 11 2 8 7 11 13 2 4 4 1 15 0 8 2 15 1 15 1 10 12 9 10 0 13 9 1 2 9 2 13 4 2
24 1 12 13 15 9 1 10 9 1 11 0 4 4 1 10 9 1 8 1 10 12 0 9 2
21 1 10 9 1 15 9 13 1 10 0 11 10 9 1 15 2 9 2 4 4 2
28 0 9 13 4 4 1 0 2 1 10 9 1 10 9 2 9 2 16 3 9 3 1 2 9 2 4 4 2
4 7 15 0 2
29 10 9 2 0 2 8 2 4 1 11 4 1 10 11 1 12 7 13 3 3 0 9 1 10 0 9 7 9 2
33 9 1 10 9 1 9 12 1 10 0 9 2 3 0 1 9 2 9 7 9 1 10 9 4 4 2 13 7 13 0 4 4 2
10 7 16 10 9 3 3 3 1 13 2
18 13 15 9 3 0 3 3 7 4 3 10 13 9 3 0 7 13 2
21 10 0 9 1 9 2 13 15 0 0 4 4 2 7 15 13 15 0 0 4 2
8 1 10 9 4 15 9 0 2
20 15 0 9 1 1 10 9 13 15 1 10 9 1 10 0 9 1 10 9 2
31 15 4 2 7 15 13 15 9 2 15 7 15 10 9 15 1 15 0 9 3 9 13 2 7 10 0 9 16 0 13 2
8 1 15 9 13 15 1 4 2
17 7 10 0 9 4 10 9 2 15 1 15 0 9 8 4 4 2
8 10 9 9 13 10 9 4 2
33 10 0 0 9 13 15 0 2 16 10 0 9 1 0 9 2 1 9 0 9 1 3 13 7 10 0 9 1 9 9 3 1 2
22 3 13 10 9 9 1 10 0 9 1 4 16 10 9 1 13 1 10 0 9 9 2
27 10 9 2 15 0 1 10 9 3 1 10 9 4 4 2 13 15 15 0 7 15 0 9 1 13 9 2
11 3 13 10 9 4 1 10 12 9 8 2
7 1 9 4 12 9 4 2
17 8 13 1 9 12 1 9 12 2 8 1 9 12 1 9 12 2
16 8 13 1 9 12 1 9 12 7 1 9 12 1 9 12 2
15 8 1 9 12 1 9 12 7 1 9 12 1 9 12 2
22 12 0 9 13 4 2 16 15 1 9 1 8 8 5 3 9 5 1 9 4 4 2
21 10 9 13 8 16 10 0 9 10 0 9 11 8 13 1 10 9 1 10 9 2
46 15 13 2 16 9 11 10 0 7 15 0 9 4 1 10 9 2 3 3 15 9 9 8 2 12 2 7 9 8 2 12 2 9 1 12 9 7 1 9 1 10 0 2 9 13 2
12 9 7 8 9 4 15 0 9 1 10 9 2
15 10 1 15 8 13 9 13 10 9 1 10 9 1 8 2
31 1 10 9 1 10 9 13 10 9 4 1 9 1 10 0 9 1 9 2 15 4 9 1 9 2 3 9 0 4 2 2
19 10 9 1 8 13 4 2 16 15 3 10 0 9 1 15 9 4 4 2
18 10 9 13 0 2 7 0 7 0 9 1 10 9 1 10 0 9 2
46 10 0 9 1 10 9 4 8 2 9 1 10 9 9 1 10 0 0 9 1 11 2 15 8 2 0 0 2 2 15 3 10 9 13 2 7 3 1 10 0 7 15 0 9 13 2
12 10 9 4 4 1 9 1 10 9 1 8 2
28 16 15 8 4 1 10 9 1 10 9 13 10 9 1 11 15 3 1 15 9 8 10 9 1 9 7 9 2
13 10 9 1 15 8 2 0 0 0 2 13 8 2
28 10 11 13 13 12 9 1 11 1 12 7 12 1 8 7 12 9 1 11 1 8 2 1 15 9 2 4 2
10 15 9 4 1 15 9 1 12 8 2
12 1 8 13 15 9 1 15 9 7 9 3 2
27 10 9 1 15 8 13 0 1 12 2 0 9 1 10 9 2 16 10 11 0 1 11 10 9 9 13 2
39 10 9 13 3 10 9 3 2 3 3 15 9 13 7 16 10 9 3 3 4 2 4 10 9 3 0 16 10 13 9 1 8 10 9 1 10 9 13 2
24 1 9 4 2 10 15 9 2 1 10 0 9 4 16 15 8 10 11 1 13 1 10 9 2
15 15 4 3 10 0 9 2 3 9 7 9 3 4 4 2
13 15 13 0 3 10 9 7 10 3 1 13 0 2
16 15 4 3 16 8 15 3 3 1 11 0 13 4 8 11 2
12 7 3 3 3 1 10 9 1 11 7 11 2
19 15 13 16 15 9 1 10 9 1 11 7 10 9 1 11 3 0 4 2
34 15 13 16 12 2 11 7 11 2 15 3 3 0 4 16 10 9 9 4 2 7 16 10 0 9 4 2 3 0 15 15 9 0 2
14 11 13 15 0 9 3 0 9 4 0 9 1 4 2
14 15 13 3 15 0 15 9 2 7 3 0 13 9 2
21 10 9 1 15 13 2 16 11 1 15 9 3 13 9 7 9 4 3 1 4 2
8 2 15 13 3 0 1 4 2
9 15 4 3 0 13 7 0 13 2
13 15 4 4 7 4 2 8 1 10 9 9 2 2
25 11 13 15 1 15 9 3 0 0 4 1 15 9 2 15 1 15 8 3 3 10 0 9 13 2
26 10 9 2 15 1 11 1 15 9 4 4 2 13 8 2 16 8 1 12 1 15 1 11 13 4 2
26 10 0 9 4 1 10 9 1 11 7 13 11 10 9 1 4 1 10 0 9 8 10 9 1 11 2
12 16 11 15 9 13 2 13 11 15 0 3 2
11 15 13 3 16 10 9 1 11 0 4 2
25 3 13 4 4 2 16 11 15 4 1 10 9 1 10 9 1 10 9 2 16 15 0 9 13 2
12 10 9 13 1 15 9 2 15 15 8 13 2
12 1 10 9 13 15 1 4 15 1 13 13 2
13 7 10 9 3 10 9 4 4 2 4 15 0 2
12 15 9 15 4 3 0 2 7 0 2 0 2
41 7 15 13 15 1 9 1 10 9 15 0 13 4 2 8 2 10 9 13 4 7 15 13 15 3 2 16 10 3 0 9 16 11 4 2 13 4 1 15 9 2
19 3 15 9 4 9 4 16 10 9 1 10 9 1 10 9 0 1 13 2
26 15 13 1 10 3 13 0 9 2 8 2 4 4 4 16 9 7 9 2 0 9 2 9 7 9 2
36 1 10 9 11 4 10 0 9 3 1 4 1 10 9 16 10 9 1 8 10 9 1 10 9 4 4 2 16 15 3 1 9 1 9 13 2
21 10 0 9 13 10 9 3 10 9 1 4 16 10 9 1 15 9 8 1 13 2
30 9 8 13 1 15 9 0 1 15 13 1 9 7 9 16 1 10 0 9 1 9 1 10 9 1 10 9 1 4 2
6 3 10 9 1 9 2
7 3 3 3 15 0 13 2
19 16 3 15 1 3 4 4 2 13 10 12 9 0 15 0 0 4 4 2
4 7 10 9 2
13 15 13 1 10 9 1 10 9 2 1 10 9 2
3 8 11 2
19 2 15 13 10 9 3 4 2 16 15 9 12 1 10 9 9 4 4 2
23 3 13 16 10 0 9 4 13 1 4 1 12 9 1 9 7 9 1 10 9 16 9 2
9 10 9 13 15 3 3 4 4 2
9 15 13 15 1 15 9 4 2 2
24 10 9 9 13 1 11 1 10 9 16 12 9 7 9 15 9 4 1 15 13 1 10 9 2
7 11 4 10 0 0 9 2
7 15 4 15 16 9 3 2
9 10 9 15 4 1 10 9 8 2
18 11 13 16 13 9 1 10 0 9 2 15 1 12 7 12 9 4 2
42 11 4 15 0 9 2 7 15 13 16 0 9 3 0 1 10 9 1 10 9 2 15 0 9 13 16 11 2 11 2 11 2 11 7 10 12 11 2 11 7 11 2
19 3 13 10 9 2 15 8 4 15 9 1 10 9 1 8 3 1 4 2
34 1 10 9 13 15 3 4 4 2 7 3 4 1 10 9 3 15 13 4 2 7 3 1 8 4 3 3 15 3 16 3 1 13 2
16 10 9 13 1 10 12 9 1 8 2 13 3 3 1 9 2
9 8 10 0 9 13 15 8 4 2
24 8 13 10 9 1 8 12 1 10 9 1 10 0 9 1 10 11 1 10 9 8 10 9 2
32 11 13 10 9 1 8 1 10 9 1 15 9 7 10 9 1 10 9 1 8 1 10 9 1 10 9 11 2 11 7 11 2
27 1 10 9 1 10 9 1 10 11 13 3 4 4 2 16 9 4 4 1 10 9 1 9 1 15 9 2
11 1 10 12 9 13 15 15 0 9 3 2
17 1 8 3 13 10 9 3 4 2 3 3 1 12 9 8 12 2
38 7 1 10 9 8 15 8 1 11 2 3 10 0 9 11 7 9 9 13 4 16 10 9 1 13 2 4 10 9 3 1 10 0 9 15 9 0 2
29 1 15 9 4 0 10 3 0 9 3 0 15 9 8 2 0 9 1 10 0 9 2 8 1 10 9 13 4 2
23 15 13 3 3 3 3 1 4 16 15 2 12 2 1 10 9 3 1 0 9 13 4 2
30 16 10 9 1 10 11 3 3 0 4 4 13 3 0 2 16 10 9 1 15 12 13 9 13 1 9 1 10 9 2
12 3 10 0 9 8 13 1 10 0 9 4 2
17 15 13 3 3 3 16 10 12 9 1 3 3 16 9 4 4 2
40 10 9 15 15 15 13 1 10 0 9 15 11 1 15 8 13 4 2 10 0 9 1 9 13 3 3 3 10 9 10 9 1 10 9 1 15 9 4 4 2
18 1 15 9 3 10 9 1 9 4 4 4 1 10 0 9 13 15 2
8 2 3 13 15 9 1 4 2
23 15 13 1 10 3 0 9 0 12 9 0 2 7 10 0 12 9 13 15 15 4 2 2
12 1 3 4 1 11 3 12 9 1 9 4 2
29 10 12 0 9 4 4 1 15 8 2 15 1 12 1 10 15 9 0 10 15 9 13 2 7 8 10 9 4 2
13 10 9 13 10 9 2 10 9 13 10 0 9 2
33 1 10 13 9 2 15 1 10 9 1 12 9 13 1 10 9 1 10 9 2 4 2 3 0 2 10 0 9 1 10 9 4 2
15 3 13 3 10 2 0 9 2 1 10 0 9 2 8 2
11 2 0 2 9 13 8 0 7 0 9 2
22 0 13 3 3 2 16 9 3 15 16 9 0 4 1 15 9 7 15 9 8 2 2
42 10 9 4 16 9 0 4 7 0 3 16 10 9 15 9 13 1 10 9 2 9 1 9 2 2 15 9 1 10 15 4 4 7 9 1 9 15 4 16 13 9 2
34 10 9 1 15 8 15 12 9 1 10 9 1 9 13 2 4 4 1 12 9 7 15 1 9 1 9 2 13 9 2 1 12 9 2
34 10 9 1 0 9 15 1 9 1 15 9 13 7 1 10 9 9 13 1 10 9 2 16 10 9 2 13 15 10 9 1 12 9 2
27 8 13 15 0 9 3 0 2 1 10 0 7 1 10 9 13 9 15 1 10 11 1 15 9 4 4 2
12 1 12 13 15 3 1 10 15 9 9 4 2
16 15 13 3 1 10 9 1 10 0 7 15 0 13 9 4 2
13 15 4 3 0 1 13 1 15 10 9 3 13 2
29 15 13 10 9 0 4 16 15 3 7 15 13 3 10 3 0 9 3 2 7 15 0 9 1 9 13 1 9 2
33 10 9 13 3 1 10 0 15 15 9 13 7 15 13 3 1 0 9 3 15 3 1 10 9 3 4 2 3 15 15 3 4 2
8 15 15 13 4 8 10 9 2
8 10 9 13 15 15 15 9 2
29 3 13 3 10 9 1 15 9 15 9 13 4 1 10 9 1 15 8 16 10 9 1 11 1 8 3 1 4 2
10 10 9 4 13 2 8 12 1 12 2
11 8 12 1 10 0 9 2 7 3 0 2
17 15 4 3 0 16 10 9 3 1 10 9 1 15 8 4 4 2
21 2 13 2 15 9 13 15 3 15 8 7 15 13 15 1 10 9 1 15 9 2
19 1 9 7 1 9 13 10 0 7 13 9 15 9 1 10 11 1 4 2
31 9 11 13 1 15 1 15 0 9 1 10 0 9 1 9 2 15 15 13 1 9 3 4 4 2 7 15 13 1 9 2
39 16 15 1 10 9 13 1 10 9 1 13 7 3 1 13 2 13 15 1 10 9 3 3 13 2 15 9 4 7 13 10 2 9 2 10 9 3 4 2
14 1 10 9 1 10 9 15 9 1 3 8 12 0 2
30 10 0 9 13 1 10 9 2 1 9 2 1 12 9 1 9 7 1 10 13 9 13 10 9 3 0 4 1 4 2
14 10 9 13 1 10 13 9 1 12 9 1 8 12 2
20 1 10 9 16 9 4 12 9 2 3 12 9 2 9 2 8 12 2 4 2
12 10 9 1 11 1 10 9 4 3 3 0 2
24 10 12 0 0 9 4 3 1 10 0 9 0 1 4 7 9 11 13 3 1 10 0 9 2
23 7 11 2 15 1 10 0 9 8 1 10 0 9 11 13 4 4 2 13 3 10 9 2
19 7 15 13 15 0 2 3 16 15 13 13 15 3 3 15 15 3 4 2
37 0 4 16 1 8 10 0 9 8 9 1 13 7 1 15 3 0 3 4 8 12 9 13 1 4 2 0 15 16 10 0 9 2 12 9 2 2
34 15 13 10 9 4 16 15 10 9 1 10 9 1 10 0 9 1 11 1 10 11 16 15 1 11 8 1 12 4 4 2 4 4 2
27 9 1 11 13 3 3 16 3 1 10 9 1 11 15 9 1 11 2 1 10 9 2 1 10 11 4 2
14 3 13 9 15 9 10 9 1 10 13 9 1 4 2
12 1 13 9 4 10 3 3 13 9 0 4 2
17 10 9 7 10 9 1 10 0 9 13 1 10 0 9 9 4 2
24 3 10 0 9 13 10 9 1 4 2 16 15 13 16 10 9 8 4 2 13 15 10 9 2
6 1 8 13 10 9 2
15 2 16 8 1 10 9 4 4 2 13 15 3 10 9 2
5 15 4 4 2 2
17 10 9 15 1 10 9 3 13 4 13 1 10 13 9 1 4 2
23 1 11 13 15 10 9 1 0 9 2 7 3 3 13 3 0 3 3 10 0 0 9 2
33 1 15 12 9 9 13 10 0 0 0 9 3 1 10 9 2 15 9 13 4 8 10 9 2 16 10 9 1 10 9 4 4 2
18 1 11 2 11 7 3 1 11 13 15 1 10 13 9 0 15 4 2
8 7 3 4 3 9 1 4 2
27 3 13 3 1 10 3 3 0 13 9 1 11 5 7 3 3 3 5 10 9 16 15 0 8 1 4 2
4 0 7 0 2
9 7 13 15 15 1 10 0 4 2
34 15 0 4 2 1 15 9 2 10 9 9 5 16 15 3 9 2 9 2 9 2 9 2 9 2 0 8 7 15 2 9 2 4 2
31 10 9 9 1 7 1 11 1 15 9 13 15 1 10 0 9 1 10 9 8 2 15 3 1 9 1 8 1 11 13 2
53 16 15 3 0 7 0 3 0 0 0 9 4 11 3 3 2 10 11 1 10 9 2 4 2 7 3 2 10 9 2 16 15 15 0 7 0 9 15 13 4 1 10 9 1 11 0 9 1 15 9 1 12 2
21 15 13 3 12 9 4 2 12 9 0 4 7 1 10 9 4 1 10 0 9 2
25 0 0 9 13 15 9 2 15 3 0 4 4 1 10 9 1 10 9 7 10 9 1 10 9 2
31 8 4 10 1 10 0 9 13 0 9 2 1 15 10 9 1 10 9 7 10 2 0 9 1 10 9 2 3 0 4 2
20 15 13 3 10 3 0 0 9 1 15 13 1 10 9 15 1 10 9 13 2
13 3 13 1 11 3 0 3 15 9 16 1 11 2
26 10 9 13 11 7 10 11 3 16 9 1 0 9 7 10 0 13 9 2 15 9 7 0 9 13 2
11 10 0 9 1 10 9 4 3 8 0 2
7 1 8 13 11 3 3 2
24 15 13 3 12 9 1 15 4 5 3 8 5 7 13 3 3 3 10 9 0 9 3 1 2
34 1 10 9 2 7 10 9 2 1 10 9 13 15 1 10 9 1 10 9 10 9 8 2 15 3 9 4 1 10 0 13 0 9 2
30 1 10 13 9 13 10 9 1 13 9 9 4 16 9 1 13 1 10 9 3 10 9 15 9 13 1 9 15 13 2
6 8 13 15 9 4 2
7 10 1 10 0 8 0 2
9 15 9 13 8 3 0 15 4 2
17 10 9 13 3 3 3 16 10 9 15 3 4 4 1 15 9 2
16 15 4 1 15 9 10 9 1 10 0 9 2 3 13 15 2
31 10 0 9 13 10 9 1 8 2 16 3 1 4 10 9 1 10 0 9 3 0 1 15 1 4 2 15 9 4 4 2
34 16 1 15 3 0 13 13 4 4 4 2 13 15 4 4 9 12 1 10 9 1 10 0 9 3 3 1 4 2 3 10 9 8 2
12 16 9 1 13 13 10 9 1 15 9 3 2
23 10 9 13 16 10 9 3 0 9 9 1 11 4 16 9 1 8 1 11 1 13 4 2
18 1 15 9 13 15 3 16 10 0 9 7 10 0 9 1 0 4 2
24 2 10 0 9 13 10 9 1 10 9 7 13 9 15 1 10 0 9 1 11 1 4 2 2
20 3 4 10 9 4 1 8 7 8 1 10 9 2 16 2 8 2 13 4 2
10 15 9 13 15 3 3 1 11 4 2
25 9 1 10 9 13 15 1 15 0 0 9 1 10 9 4 1 10 9 1 10 9 7 10 9 2
17 12 9 13 10 9 4 1 9 11 3 8 9 10 9 4 4 2
11 3 13 10 9 1 10 9 11 4 4 2
12 1 9 8 13 10 9 10 9 3 0 3 2
28 2 16 15 4 4 10 9 1 15 9 8 8 1 4 2 3 4 15 15 15 10 9 1 10 9 0 13 2
40 16 15 3 4 4 1 9 16 9 11 7 9 11 16 0 9 1 13 2 3 13 15 10 0 9 9 16 15 3 1 10 0 9 1 10 9 3 13 2 2
28 9 11 10 9 1 11 2 13 10 9 1 9 11 4 10 9 1 10 0 9 1 10 9 3 0 1 4 2
22 8 2 9 1 10 9 1 8 2 8 2 2 4 4 1 9 1 10 9 1 11 2
17 10 9 1 9 2 8 2 13 10 9 3 1 11 1 8 4 2
19 0 4 15 2 16 3 4 4 2 4 1 10 9 1 10 0 0 9 2
17 9 8 13 10 9 4 2 16 15 1 15 9 15 9 3 4 2
23 8 13 1 11 3 10 9 8 2 15 10 9 15 13 4 1 15 9 1 10 0 9 2
20 15 9 13 3 3 2 1 10 9 2 2 3 1 9 1 0 9 4 4 2
31 3 13 1 9 12 2 9 2 7 9 12 2 0 9 2 1 10 9 1 9 10 9 1 0 9 1 10 9 4 4 2
7 10 9 13 10 0 9 2
4 10 0 9 2
16 15 13 15 3 1 10 9 3 1 15 8 7 8 1 9 2
28 10 9 16 0 9 4 3 1 13 9 1 15 9 13 2 3 8 0 9 1 10 9 1 15 9 1 9 2
18 4 4 10 9 1 9 3 1 4 16 10 9 13 7 10 9 13 2
9 12 9 13 1 4 8 0 9 2
30 0 13 10 13 9 1 10 9 1 4 4 16 10 0 9 1 13 4 7 16 1 13 16 13 9 10 0 9 4 2
15 11 13 5 16 15 0 9 3 1 13 5 4 4 4 2
23 10 9 1 9 1 9 13 11 1 11 1 9 9 4 1 10 9 1 10 9 1 9 2
19 3 13 10 0 9 1 9 4 4 1 15 1 10 9 13 7 13 9 2
15 1 10 9 1 15 9 13 10 0 9 3 10 9 4 2
21 9 11 13 3 16 15 15 0 4 4 16 10 0 0 9 1 12 9 1 9 2
5 3 4 11 15 2
10 3 13 15 15 15 10 9 13 4 2
40 7 11 13 3 5 1 15 1 10 0 0 9 13 15 3 3 15 9 1 0 9 1 4 5 7 15 13 3 1 9 10 9 10 1 9 13 0 9 4 2
4 2 8 2 2
4 13 15 9 2
12 15 13 3 2 13 3 10 0 9 7 13 2
14 11 4 1 10 9 1 15 9 1 11 1 8 4 2
4 2 8 2 2
4 15 4 4 2
11 1 10 9 1 10 9 4 15 15 9 2
18 3 13 3 3 15 9 8 4 2 3 10 9 13 1 10 9 13 2
22 10 9 1 10 2 13 2 9 4 0 3 4 7 3 13 9 1 9 1 10 9 2
15 8 3 4 3 4 1 10 0 9 1 10 0 0 9 2
17 3 13 10 9 1 10 9 15 3 13 9 1 4 1 12 9 2
4 11 1 11 2
54 10 9 1 9 1 10 9 1 10 0 9 13 1 9 1 9 11 2 9 2 7 9 8 2 9 2 4 10 9 1 15 3 15 9 3 1 4 16 10 9 3 3 0 3 1 13 8 11 7 10 9 0 9 2
21 15 13 3 4 16 10 0 0 9 4 4 1 10 9 1 10 9 7 10 9 2
23 16 10 9 3 0 4 4 2 13 10 9 15 11 1 15 1 9 13 4 1 12 9 2
14 15 9 13 3 1 10 9 2 8 2 3 15 9 2
37 10 9 1 10 11 13 0 1 15 8 2 16 15 1 10 0 9 9 13 4 1 10 11 9 1 10 9 3 15 1 12 1 10 9 13 4 2
18 1 10 15 9 4 15 3 3 0 2 7 3 13 15 0 1 9 2
21 15 13 9 8 1 15 9 1 10 9 1 10 11 9 2 16 12 13 4 4 2
55 7 10 1 11 0 13 9 1 15 3 13 2 4 4 2 15 1 9 1 13 5 16 3 1 9 4 1 4 5 13 10 0 9 7 9 3 0 15 0 3 16 10 2 1 9 1 3 0 2 0 7 3 13 11 2
21 1 15 9 13 3 3 15 15 10 9 1 9 1 0 9 1 15 9 1 9 2
16 15 13 3 15 4 16 10 9 10 9 3 3 4 4 4 2
23 9 8 13 3 1 10 1 11 13 9 4 16 10 9 1 10 13 0 9 4 4 4 2
24 10 0 9 1 12 7 0 9 13 2 3 13 15 2 3 4 4 1 9 1 15 13 9 2
44 10 9 11 13 1 4 16 10 0 0 9 1 10 9 2 3 10 0 0 9 1 10 0 9 13 4 2 3 4 9 1 4 1 9 1 9 11 16 10 11 3 1 4 2
34 3 13 10 0 9 1 9 13 2 4 8 1 10 9 1 10 9 15 1 10 9 13 7 10 0 9 15 3 1 10 9 4 4 2
16 7 3 10 9 1 10 0 9 2 10 9 1 9 7 9 2
10 10 9 1 11 4 13 7 3 13 2
17 10 9 1 9 7 9 2 10 9 1 10 0 9 2 4 13 2
13 7 3 15 9 13 16 10 9 15 9 13 4 2
16 9 15 13 1 10 9 1 10 0 9 13 1 15 10 9 2
17 10 11 13 3 10 9 16 15 1 10 0 9 1 12 13 4 2
22 2 15 13 4 15 15 0 1 4 4 16 10 9 1 15 3 3 3 13 4 2 2
33 15 4 15 1 10 9 1 10 9 1 8 15 1 11 10 9 8 13 4 2 15 4 4 1 10 11 11 11 8 10 0 9 2
21 10 9 2 15 0 1 11 4 4 2 13 10 9 3 15 1 10 9 4 4 2
23 3 1 10 0 9 13 11 10 9 3 1 10 0 13 9 11 7 13 15 3 3 3 2
15 15 13 3 3 1 10 9 16 10 13 9 3 1 4 2
15 8 13 15 10 9 1 8 9 2 12 9 1 9 2 2
49 10 1 15 15 1 10 12 9 2 1 10 9 13 0 9 2 12 9 1 9 2 13 15 3 3 4 2 16 10 9 1 10 9 1 10 1 10 9 10 9 13 3 1 4 1 10 0 9 2
22 15 1 10 10 9 1 10 13 9 4 2 16 9 11 15 0 13 1 4 1 11 2
35 10 9 13 15 0 9 1 10 9 2 1 8 2 1 9 16 11 1 12 1 12 9 7 11 1 12 1 12 9 1 10 9 1 13 2
11 8 13 10 0 0 9 1 10 0 11 2
20 11 13 10 9 3 1 12 7 11 13 10 11 3 3 10 9 1 15 9 2
2 12 2
25 15 0 9 2 16 9 0 9 1 11 10 0 9 13 4 2 13 1 15 9 10 0 0 9 2
12 3 3 13 3 12 9 13 7 0 1 11 2
24 10 9 4 10 0 9 0 9 2 1 0 9 15 0 4 10 9 1 10 0 9 1 4 2
13 15 13 10 9 1 15 9 3 9 1 10 9 2
29 1 0 9 13 3 15 8 2 3 8 15 0 9 3 13 7 8 13 1 10 3 0 9 11 2 8 7 8 2
33 3 13 8 10 9 1 9 11 8 16 15 13 16 10 0 9 3 8 4 4 16 1 12 1 12 9 13 16 10 9 13 4 2
32 10 9 16 0 15 15 9 13 8 10 9 15 9 4 4 16 15 3 0 4 16 12 9 2 13 10 9 11 10 0 9 2
15 3 3 3 10 9 1 10 0 2 2 13 15 15 3 2
23 11 7 11 13 15 4 1 10 1 11 13 9 1 9 2 11 2 2 3 13 15 8 2
22 1 15 9 2 15 1 12 1 0 9 4 4 2 4 3 4 11 2 11 7 11 2
9 9 4 13 1 10 9 1 11 2
13 1 10 9 12 9 3 13 11 3 12 9 4 2
31 0 1 10 9 4 3 16 10 9 11 2 15 16 10 0 9 1 11 4 4 1 12 9 4 4 7 15 0 8 13 2
26 0 0 4 8 2 15 1 10 9 2 15 13 12 9 1 11 4 2 10 13 9 4 1 4 4 2
7 15 4 10 9 4 9 2
22 7 11 2 15 15 3 0 13 4 1 15 9 7 1 10 9 1 10 9 13 3 2
15 3 13 3 9 8 1 10 0 9 3 10 11 13 4 2
12 3 1 11 2 3 10 11 11 15 8 13 2
8 1 11 13 9 7 9 4 2
15 10 9 15 0 0 4 2 13 3 3 4 3 1 4 2
19 7 0 13 15 3 10 9 8 3 10 0 9 3 2 3 3 2 13 2
19 10 0 4 15 2 3 0 10 9 4 2 8 0 10 9 10 9 4 2
17 10 1 12 0 0 9 8 4 1 15 8 10 0 9 10 9 2
21 8 4 15 9 7 9 8 2 15 1 15 13 8 11 8 7 11 8 13 4 2
20 7 11 13 10 9 7 11 2 3 9 1 10 9 1 11 13 8 11 4 2
10 15 13 4 15 13 9 3 1 13 2
34 0 4 15 1 15 0 9 1 9 1 11 1 11 11 2 10 3 0 16 0 9 2 15 15 3 3 15 13 2 7 1 11 11 2
14 15 13 16 10 8 13 9 3 0 4 1 10 9 2
33 10 9 1 10 3 13 9 4 16 10 9 11 0 10 9 13 4 5 0 1 11 2 7 3 8 10 9 1 9 1 15 9 2
15 8 13 3 1 4 16 11 15 9 1 15 0 9 4 2
15 15 13 15 8 2 11 2 1 15 9 8 1 15 9 2
25 10 13 9 2 3 10 11 2 13 15 3 3 1 10 9 2 1 10 9 2 8 1 10 9 2
25 1 10 9 4 15 3 3 0 2 1 15 9 3 2 9 3 1 13 1 15 13 1 0 9 2
19 13 3 9 3 2 3 13 15 0 10 9 4 1 10 9 1 10 9 2
16 1 0 15 9 4 10 9 16 11 3 0 16 9 13 4 2
7 15 13 15 9 4 4 2
27 11 13 1 10 9 12 2 8 10 0 8 7 8 2 4 1 10 0 9 16 9 10 0 9 1 4 2
30 1 10 9 1 11 1 10 0 9 2 3 1 10 9 2 16 15 13 7 13 2 13 9 7 9 8 10 0 9 2
9 10 9 1 9 4 10 0 9 2
21 15 1 10 10 9 1 10 10 9 15 10 9 13 8 1 10 9 7 1 15 2
18 2 9 2 9 7 9 13 15 3 2 9 4 4 1 9 7 9 2
6 15 4 1 15 0 2
7 7 15 9 13 4 0 2
18 15 9 4 4 7 0 1 9 1 10 0 9 4 15 16 9 4 2
20 15 13 3 1 15 15 2 3 1 10 13 9 2 7 10 9 4 3 15 2
19 3 8 1 10 2 0 2 9 13 15 8 10 9 4 1 8 1 11 2
31 13 4 10 15 3 0 9 2 7 15 4 4 1 10 13 9 1 10 9 12 2 15 1 9 8 0 4 4 7 4 2
29 3 1 10 0 9 1 15 9 13 10 9 1 10 9 15 9 16 3 15 0 9 2 3 9 2 1 13 4 2
12 0 9 4 3 1 15 9 3 1 11 4 2
17 15 9 2 15 3 15 9 13 2 13 10 9 3 1 10 9 2
40 16 15 0 2 0 9 4 4 5 3 16 3 0 9 3 13 2 16 3 10 9 4 4 1 10 9 1 9 3 5 3 4 10 9 0 10 9 3 4 2
13 10 13 9 2 9 3 4 1 12 9 0 4 2
24 10 9 9 15 1 10 9 4 4 13 10 9 1 10 9 3 15 10 1 9 13 9 13 2
14 1 0 11 13 10 9 3 1 10 0 9 10 9 2
46 15 13 15 9 7 1 0 7 1 9 2 16 15 13 4 1 10 9 1 0 9 7 10 0 9 1 0 9 7 0 9 3 10 13 0 9 2 1 10 13 9 2 9 2 13 2
22 15 4 4 1 10 9 1 8 7 3 13 10 9 1 15 3 2 15 15 16 8 2
11 10 9 4 4 1 15 10 9 9 13 2
39 15 13 15 3 2 16 15 13 4 4 16 3 1 15 9 9 1 10 13 11 15 9 4 4 5 3 13 15 9 1 10 9 15 3 15 0 9 4 2
26 1 8 11 4 8 10 0 9 1 10 8 9 11 15 1 10 0 9 4 4 2 11 2 11 2 2
12 3 3 16 0 9 15 1 10 9 13 4 2
30 15 4 10 9 1 8 2 15 16 15 1 10 0 9 1 11 10 9 1 10 9 13 4 4 7 3 15 3 13 2
40 15 4 10 9 2 1 11 2 1 10 9 2 10 9 15 1 10 9 9 13 2 3 3 1 15 9 3 3 1 15 9 2 3 1 10 9 2 10 9 2
37 1 10 9 11 7 11 13 10 11 8 10 9 4 4 16 1 15 0 0 8 1 4 2 7 3 3 10 9 3 0 9 1 15 9 1 4 2
27 15 13 3 3 3 0 15 9 15 4 4 1 10 9 1 10 9 15 13 1 10 9 1 10 13 9 2
16 8 13 3 15 15 9 1 4 1 10 9 1 10 13 9 2
38 1 10 9 11 2 1 10 9 1 11 2 4 12 9 13 4 7 13 12 15 4 1 15 10 9 11 13 2 9 2 15 1 12 1 12 13 4 2
9 1 10 9 4 10 9 3 4 2
28 10 9 1 10 9 4 1 10 0 9 10 9 8 2 15 9 13 4 4 1 12 9 15 9 13 4 4 2
6 15 9 4 3 4 2
13 12 9 9 13 15 9 1 11 2 15 15 13 2
14 8 13 1 12 1 11 2 8 4 3 3 12 9 2
5 15 4 0 9 2
25 15 4 4 1 9 2 9 2 9 2 9 2 9 2 9 2 9 2 8 7 9 1 10 9 2
21 11 4 1 10 9 4 16 10 9 1 11 7 8 2 13 1 4 1 9 2 2
24 1 11 13 15 10 0 9 1 12 9 1 15 9 15 11 1 10 0 9 1 11 0 13 2
27 10 9 13 16 2 8 15 9 1 9 11 2 10 0 9 15 0 9 4 16 9 1 15 1 9 11 2
22 15 13 15 0 8 4 15 1 9 13 9 1 4 15 15 0 13 1 10 0 9 2
16 11 13 3 1 15 9 3 3 15 9 4 16 11 7 11 2
36 15 13 3 3 8 4 2 3 8 2 16 10 0 9 4 16 3 3 3 10 9 4 15 1 10 1 15 13 9 2 9 1 10 9 13 2
16 1 10 9 1 10 9 13 10 9 15 1 10 9 3 4 2
19 15 4 3 1 10 9 10 0 9 16 10 9 1 13 1 15 0 9 2
25 1 9 2 15 3 0 1 15 13 16 9 7 9 2 13 11 7 11 15 9 1 0 9 4 2
24 2 15 4 0 16 2 3 2 13 9 1 10 9 1 10 9 1 9 1 0 9 4 4 2
39 8 13 4 4 1 10 0 3 0 13 9 7 1 9 1 10 9 1 10 9 10 9 1 10 9 1 10 9 1 4 16 3 10 9 1 13 4 2 2
7 2 8 2 9 12 2 2
24 2 10 9 1 9 1 10 0 9 13 10 9 4 16 1 4 1 10 0 9 1 15 9 2
18 6 2 10 9 2 3 10 0 2 0 9 2 13 3 3 0 3 2
39 1 10 9 1 15 8 13 15 15 8 1 11 2 0 13 2 4 7 10 11 1 11 2 0 13 2 2 7 3 11 9 1 10 9 1 8 16 9 2
18 3 8 4 15 9 4 1 15 0 13 2 8 2 1 8 7 8 2
12 9 13 1 10 9 1 11 2 15 1 11 2
18 15 13 3 0 2 7 3 3 15 0 2 1 9 3 15 0 4 2
18 10 9 1 15 4 1 0 9 4 2 15 4 3 3 0 1 4 2
22 1 12 1 12 1 10 9 13 12 9 1 12 7 12 9 1 10 9 1 10 9 2
25 2 1 15 13 3 15 1 8 1 11 1 11 0 2 10 15 13 1 8 2 13 1 11 2 2
27 0 13 11 3 15 9 2 16 11 2 15 10 9 1 15 9 10 2 1 10 0 9 0 9 2 13 2
28 10 0 0 9 1 9 7 9 2 11 2 13 11 16 15 9 4 16 11 10 9 1 12 9 4 4 4 2
48 1 11 13 15 0 8 2 16 10 9 1 10 9 1 10 9 1 10 0 13 9 1 15 4 13 2 10 9 1 12 9 9 7 13 15 1 10 9 1 10 9 3 3 12 9 1 4 2
18 10 9 4 1 8 7 15 1 12 4 7 10 9 13 1 12 9 2
7 0 13 13 15 3 3 2
20 5 2 15 13 10 9 7 9 16 1 10 15 9 1 10 0 9 1 4 2
6 5 15 13 0 9 2
15 5 15 13 10 9 1 15 13 1 10 9 1 15 9 2
12 5 15 13 10 0 9 2 0 9 2 9 3
20 15 13 3 3 2 15 13 0 16 9 8 2 15 9 13 2 15 13 4 2
12 5 15 13 9 1 10 9 1 15 0 9 2
16 10 9 2 15 1 10 0 9 9 13 4 2 13 9 4 2
12 3 3 10 9 0 4 2 15 9 3 8 2
24 1 10 9 13 10 9 3 3 3 0 2 7 15 4 1 15 9 1 10 9 1 10 9 2
42 1 12 2 16 10 9 1 8 2 10 0 9 1 11 1 3 12 12 9 2 1 10 9 1 9 4 4 2 4 3 15 4 16 1 10 0 9 7 9 1 13 2
20 1 9 1 9 13 15 1 10 0 9 8 4 1 10 0 9 1 10 9 2
16 10 1 15 8 13 9 9 1 12 9 4 3 3 3 8 2
29 11 13 3 1 12 7 15 9 3 1 9 2 3 1 10 0 9 7 10 0 9 2 10 9 1 10 9 4 2
10 3 13 3 10 0 0 9 4 4 2
2 3 2
45 1 15 9 13 1 3 0 9 10 9 2 10 9 13 10 9 1 10 9 2 13 10 9 3 2 9 1 10 9 1 2 15 8 4 4 2 3 1 10 9 1 10 9 1 2
27 15 15 1 15 13 7 13 9 13 7 1 15 0 13 1 10 0 9 13 2 13 15 9 0 4 4 2
36 10 9 4 3 3 15 0 3 2 7 15 13 3 1 4 3 1 10 9 10 9 2 0 3 0 7 0 2 1 9 1 4 7 1 4 2
14 6 2 15 13 3 3 3 3 9 1 15 3 4 2
13 15 9 13 10 9 1 15 0 9 8 4 4 2
10 3 8 2 9 4 15 1 9 0 2
20 10 11 13 10 0 9 1 10 9 8 2 13 1 10 9 1 9 7 9 2
12 15 4 1 15 0 16 1 15 9 1 13 2
33 10 9 7 9 5 16 1 10 9 1 13 5 13 15 3 3 1 0 9 3 7 13 3 1 10 13 9 1 9 1 10 0 2
9 15 0 9 1 10 9 4 4 2
5 4 4 3 3 2
16 10 9 1 12 13 1 15 0 9 8 1 10 0 9 4 2
11 12 10 9 13 1 10 9 1 10 9 2
23 15 4 15 0 2 7 15 13 15 4 16 15 13 1 15 9 1 10 9 15 9 4 2
5 3 13 15 3 2
18 1 10 9 1 10 9 1 10 9 7 3 3 3 1 10 15 9 2
24 1 10 9 12 13 15 10 0 9 4 2 16 10 9 1 10 9 3 15 0 9 13 4 2
16 10 0 9 4 9 13 9 2 16 15 9 4 4 2 4 2
5 10 0 9 4 2
10 9 12 2 0 9 8 2 9 8 2
13 0 9 8 2 3 12 9 2 15 13 3 8 2
13 0 9 8 2 3 12 9 2 15 13 3 8 2
22 3 1 10 13 9 1 8 4 1 10 9 1 15 9 3 3 12 9 9 1 4 2
1 2
10 3 13 12 9 9 4 1 10 9 2
10 16 15 12 13 11 2 11 7 11 2
7 15 12 13 3 9 4 2
15 10 0 9 4 11 2 1 10 9 10 9 1 10 11 2
11 11 13 1 9 1 9 3 15 9 4 2
38 1 10 9 1 10 9 1 9 7 9 4 10 9 1 11 3 4 1 1 10 9 16 10 12 9 15 3 13 4 15 1 15 0 4 1 10 9 2
22 3 1 9 2 3 10 9 3 15 9 1 4 13 2 13 3 10 0 9 4 4 2
18 9 1 10 0 9 4 3 0 9 2 16 8 10 9 1 8 13 2
39 1 9 1 10 9 1 15 9 2 3 15 10 0 9 1 10 9 7 10 0 9 13 2 7 1 10 0 9 2 4 10 9 3 8 1 10 9 4 2
19 10 9 13 3 1 11 4 11 15 13 9 1 10 9 1 9 4 4 2
29 16 15 9 1 11 10 0 9 1 13 13 15 1 15 10 9 1 15 9 3 2 3 15 0 15 9 13 4 2
30 10 0 9 1 11 4 10 9 7 3 4 1 10 0 3 0 0 9 10 0 9 0 1 11 1 11 7 11 4 2
52 16 3 3 15 0 9 0 4 13 10 9 1 0 9 3 4 4 16 16 15 9 1 10 9 7 9 0 9 13 4 2 3 13 10 9 11 1 0 9 7 9 8 9 1 10 9 11 2 9 2 4 2
15 0 9 4 0 0 1 10 0 1 3 1 9 0 9 2
17 10 9 1 10 9 13 4 4 16 0 0 9 7 9 0 13 2
21 10 9 4 10 0 9 15 1 10 9 4 4 7 10 0 15 4 4 1 12 2
24 10 9 16 10 11 10 9 1 11 4 4 4 4 1 10 9 1 3 1 10 9 1 11 2
20 10 0 9 13 3 4 16 12 0 9 1 11 4 4 7 10 15 4 4 2
18 10 9 13 2 3 15 9 2 0 4 4 16 0 9 3 1 13 2
19 16 10 9 1 15 8 13 2 4 10 9 1 10 9 15 3 1 4 2
21 15 13 1 10 0 9 1 9 7 11 2 1 11 2 11 2 4 1 0 9 2
21 9 3 13 4 3 10 9 1 10 11 2 15 9 13 1 10 9 1 10 11 2
32 12 9 2 9 8 2 12 2 7 9 8 2 12 2 2 4 3 1 10 9 1 10 11 1 11 4 1 10 3 0 9 2
20 8 10 9 4 9 1 10 9 4 1 12 0 9 2 15 8 7 15 8 2
40 1 10 9 13 3 10 11 1 12 1 15 9 1 12 9 1 10 11 4 16 15 9 1 4 15 4 4 1 8 7 1 8 2 10 9 1 10 9 2 2
18 10 9 13 3 13 9 4 1 8 7 1 15 8 7 1 10 9 2
24 10 9 1 10 9 4 1 10 9 4 2 7 9 1 9 11 13 1 3 1 15 9 4 2
34 9 11 2 9 2 13 3 8 0 9 1 10 9 11 1 15 8 4 2 16 9 4 4 1 10 0 9 1 10 9 1 0 9 2
13 10 9 13 3 4 10 9 15 9 8 4 4 2
16 15 13 3 2 16 1 15 13 1 15 9 9 4 4 4 2
30 10 9 11 13 1 10 9 1 15 9 4 1 2 10 0 13 2 9 3 10 9 1 15 8 1 11 4 4 4 2
33 7 3 0 15 9 3 13 4 1 10 0 9 8 0 9 2 15 13 3 3 1 15 9 1 10 9 2 10 9 2 10 9 2
23 3 13 10 9 0 4 2 16 16 15 3 15 3 3 13 7 3 10 9 3 8 13 2
10 9 8 4 0 13 1 10 11 4 2
12 3 13 10 9 16 11 3 1 9 4 4 2
6 13 3 3 3 3 2
11 10 0 9 13 3 10 0 9 3 4 2
14 2 1 10 9 13 10 0 9 2 8 2 3 2 2
2 8 2
24 2 3 4 0 15 9 1 4 1 10 9 0 9 1 10 9 1 15 9 1 9 7 9 2
11 3 4 15 9 1 4 1 15 12 9 2
25 7 16 15 3 3 13 2 13 15 3 3 0 4 4 2 7 3 13 15 3 1 15 1 2 2
10 2 10 9 13 11 0 9 4 2 2
36 1 11 4 8 1 10 9 10 9 8 1 10 0 0 9 8 8 4 2 10 9 15 10 0 9 13 1 10 9 1 11 2 1 0 9 2
9 10 15 9 13 1 9 3 4 2
16 10 9 4 1 10 9 3 0 4 16 15 0 7 0 9 2
24 10 9 4 4 1 15 9 8 2 1 15 8 1 10 9 2 8 2 1 15 8 3 13 2
9 2 10 9 1 10 9 4 13 2
40 15 13 1 10 9 1 10 11 2 10 9 11 1 11 2 2 1 0 9 2 2 4 0 10 0 9 1 15 13 1 10 0 9 1 10 11 2 15 8 2
20 15 9 4 0 13 1 10 0 9 7 10 9 1 10 0 9 1 10 11 2
27 10 9 13 1 3 1 11 10 9 4 2 3 10 9 1 10 11 2 8 7 10 10 9 0 13 4 2
34 7 15 13 3 16 10 9 1 11 15 0 4 4 7 16 15 3 3 1 11 0 1 10 9 4 4 16 1 10 0 9 1 11 2
16 0 4 0 10 9 1 10 9 1 10 0 9 8 7 8 2
27 10 0 13 15 1 10 0 9 3 4 16 10 9 1 10 0 9 7 3 1 11 4 15 9 3 0 2
18 1 11 4 4 16 9 1 10 9 4 4 1 10 9 1 10 9 2
13 1 10 9 13 10 9 16 15 10 9 4 4 2
15 9 11 13 3 1 10 9 11 4 16 10 9 1 4 2
14 0 13 15 1 4 16 10 9 0 7 0 4 4 2
25 10 1 10 9 13 9 1 9 2 10 9 1 10 0 0 9 1 11 2 13 3 1 8 0 2
44 1 10 1 15 0 9 2 3 1 10 0 9 1 10 13 9 16 3 15 13 7 9 1 10 9 4 2 13 3 10 9 2 3 0 2 9 1 10 9 11 1 11 4 2
13 15 13 2 1 13 9 2 10 9 1 10 9 2
7 0 4 15 1 11 4 2
24 10 9 13 3 1 4 1 10 9 3 10 9 1 10 9 11 4 4 2 7 15 13 3 2
27 1 15 8 7 10 0 9 1 10 9 13 10 9 11 10 0 9 4 15 13 16 15 9 3 0 4 2
16 15 9 13 15 1 10 1 11 1 9 4 9 1 10 9 2
21 10 9 1 10 0 9 4 10 0 0 9 1 9 15 15 11 13 9 1 4 2
12 15 4 1 15 9 1 10 9 3 3 4 2
37 3 4 10 9 1 10 9 10 9 9 3 1 4 2 0 9 1 11 2 11 2 11 7 11 2 9 3 3 10 9 10 9 2 9 2 13 2
23 3 13 4 3 10 9 1 8 7 8 2 10 12 0 9 1 8 15 15 3 0 13 2
35 3 2 9 2 7 10 0 2 11 2 13 1 15 15 9 15 15 0 9 1 7 0 0 8 13 16 10 0 9 15 3 3 0 13 2
31 7 3 4 13 4 13 3 1 9 4 1 10 9 10 0 9 2 15 15 3 3 3 13 4 1 10 9 1 10 9 2
26 15 13 8 3 10 9 4 1 12 1 15 9 2 1 10 0 0 9 1 10 9 1 8 1 11 2
26 11 13 3 4 4 2 16 15 1 10 9 15 9 3 4 16 1 15 9 1 10 9 3 4 4 2
56 3 10 9 15 1 10 2 9 2 1 9 7 9 1 11 2 1 10 9 1 9 2 9 7 9 1 11 7 1 10 9 1 9 7 9 1 8 15 9 0 15 9 10 9 3 0 4 4 4 16 16 15 15 13 4 2
10 3 4 10 9 1 0 9 1 4 2
13 3 10 9 13 1 10 0 9 7 10 0 9 2
17 15 13 3 10 9 4 4 2 1 15 10 9 1 11 1 13 2
26 3 13 0 9 1 10 9 2 15 15 2 1 12 9 1 11 1 4 4 2 13 4 3 1 4 2
31 10 0 9 2 13 1 10 9 1 10 9 1 10 9 2 13 9 1 11 10 0 9 3 1 10 1 11 13 0 9 2
23 11 2 1 10 0 9 7 12 9 1 9 2 13 10 9 15 11 10 9 1 12 13 2
17 8 10 0 9 1 12 9 13 10 13 0 9 10 9 0 4 2
37 10 9 8 2 11 2 13 9 11 2 9 2 4 2 16 10 9 1 9 10 0 9 11 4 4 12 9 9 1 9 1 9 1 11 1 4 2
14 3 4 15 9 3 3 1 11 4 3 10 9 11 2
27 15 13 3 3 2 16 11 3 9 3 4 1 9 1 10 0 9 15 1 9 1 10 11 13 4 4 2
20 3 4 10 0 9 1 11 4 1 9 1 0 1 9 1 10 9 1 11 2
34 16 3 15 9 4 4 13 15 9 1 10 9 1 10 0 9 1 12 9 4 4 1 9 2 15 3 0 9 13 16 11 0 13 2
38 10 9 1 10 9 4 1 13 1 10 9 0 9 1 10 0 9 1 11 2 16 15 13 1 10 9 7 15 13 1 9 1 10 9 1 10 9 2
17 3 13 1 11 10 9 1 10 9 2 9 8 2 10 9 3 2
12 10 9 3 15 15 13 2 4 3 3 13 2
16 15 13 15 8 10 9 1 9 2 15 10 9 1 9 13 2
45 1 15 9 4 3 4 16 8 10 0 9 1 10 9 0 1 10 2 9 2 1 10 9 0 4 7 16 3 3 4 4 4 1 9 2 15 10 9 1 15 15 9 0 13 2
15 3 13 3 10 13 0 9 7 3 10 9 15 15 4 2
18 9 1 10 9 1 10 9 1 10 9 3 2 7 15 13 10 9 2
20 16 10 9 1 9 3 13 4 16 10 0 9 1 10 9 13 4 3 0 2
24 3 13 11 2 10 9 1 10 0 9 2 16 3 3 10 9 1 13 1 12 0 9 4 2
18 10 9 11 9 1 10 11 2 13 10 0 9 1 10 9 10 9 2
28 10 9 11 13 15 9 1 15 8 1 10 9 1 10 9 1 9 2 8 10 9 1 10 11 1 10 9 2
25 10 9 11 13 16 15 9 1 15 9 9 2 13 16 3 12 2 4 1 10 9 1 10 9 2
18 4 3 15 4 2 3 13 9 3 3 3 2 13 1 3 13 9 2
4 3 13 15 2
13 12 9 0 9 2 3 0 4 4 2 7 9 2
38 13 15 3 3 15 10 9 1 10 9 4 4 2 3 13 15 1 12 9 1 15 9 15 3 1 4 2 7 15 4 7 4 10 9 1 10 9 2
18 10 0 9 4 15 0 8 2 10 0 9 2 13 1 8 1 11 2
38 13 1 10 3 13 9 1 10 9 1 10 9 1 11 7 15 8 8 10 9 2 8 2 2 13 10 13 9 15 3 3 10 9 3 3 4 4 2
29 10 9 13 0 10 9 10 9 1 10 9 1 9 2 9 7 9 1 9 7 9 1 10 9 16 0 3 4 2
7 10 9 13 10 9 0 2
9 15 13 0 9 7 3 0 9 2
23 11 9 1 9 7 2 1 15 9 10 9 1 9 2 13 3 10 0 9 1 10 9 2
45 1 10 13 9 1 10 9 13 10 9 1 10 0 9 1 9 8 9 1 9 9 7 15 9 2 15 1 10 10 0 9 3 11 10 9 13 2 13 13 1 1 9 13 9 2
23 1 12 1 12 13 10 9 9 15 1 9 1 10 9 1 9 13 2 1 12 1 12 2
19 2 11 13 0 12 12 9 2 11 3 12 12 5 3 13 11 9 2 2
7 1 12 4 15 9 12 2
7 8 10 9 1 15 9 2
20 8 13 1 10 9 1 0 9 7 3 0 9 10 9 1 10 9 1 4 2
41 15 13 0 10 9 9 2 16 9 1 9 1 9 2 9 1 10 9 1 15 9 2 9 1 0 9 3 1 0 9 2 7 9 1 10 9 1 9 1 9 2
28 10 9 1 8 2 9 1 10 9 10 9 2 16 10 9 1 0 7 0 9 1 4 13 10 0 9 4 2
13 1 10 0 9 1 12 9 13 8 15 9 4 2
27 16 9 1 15 9 13 15 3 2 16 3 1 10 13 9 10 9 1 13 2 13 7 9 4 4 2 2
14 10 0 9 11 13 4 4 1 10 9 8 1 11 2
17 10 9 13 1 12 1 11 4 4 2 16 11 15 12 9 4 2
18 10 9 4 2 16 11 12 9 1 10 9 1 12 12 9 13 4 2
19 15 9 13 9 0 3 1 12 1 10 11 2 8 2 11 2 1 4 2
10 2 15 13 15 15 9 1 13 2 2
13 3 13 12 9 3 1 15 9 1 15 4 4 2
17 15 9 13 15 0 3 4 1 10 9 7 1 15 13 1 9 2
7 15 1 15 9 13 4 2
20 7 13 16 3 10 0 9 3 4 2 3 13 15 0 9 1 10 0 9 2
17 1 10 11 13 9 1 10 9 1 9 1 10 9 7 0 9 2
15 1 10 9 1 9 7 9 13 0 7 0 9 10 9 2
15 10 9 4 1 0 0 13 2 7 4 1 15 9 4 2
17 3 13 9 1 10 0 9 1 10 9 1 10 0 9 4 4 2
7 1 0 9 13 15 3 2
9 15 13 1 0 9 15 0 9 2
33 2 15 3 0 1 15 1 4 13 3 9 13 1 10 9 16 15 1 13 9 4 5 4 16 15 15 9 8 3 3 0 13 2
15 1 10 9 4 15 10 9 7 15 4 0 1 9 4 2
29 2 10 13 9 13 3 3 10 0 9 1 10 0 9 2 15 0 9 13 0 0 9 2 15 9 2 15 9 2
14 1 10 9 4 8 15 9 1 10 16 12 9 0 2
16 15 4 8 2 9 1 8 15 1 0 3 16 9 9 13 2
11 15 4 8 2 15 1 11 3 13 9 2
7 3 13 15 10 0 9 2
57 3 4 15 3 3 0 7 1 15 9 15 8 1 15 1 15 13 13 15 3 4 3 11 10 9 1 10 0 9 7 10 0 13 9 1 0 9 4 4 1 10 0 9 1 10 9 12 2 15 0 7 0 1 10 9 13 2
19 2 10 0 9 13 9 1 9 2 3 15 15 0 0 9 13 4 2 2
13 15 13 3 8 2 9 1 15 8 1 10 9 2
15 15 13 15 0 16 15 8 15 3 1 13 9 4 4 2
20 1 10 9 1 12 13 10 9 1 9 7 9 10 9 0 16 1 0 9 2
14 15 13 2 3 10 9 2 3 1 9 1 0 9 2
35 10 9 11 4 3 8 16 9 4 4 4 1 10 9 1 10 0 9 1 10 13 0 9 7 10 9 3 10 9 1 15 9 13 4 2
19 10 9 15 15 8 1 12 13 4 3 13 7 0 0 16 15 1 12 2
10 10 9 13 8 2 3 12 2 12 2
20 10 9 4 8 2 12 2 12 2 3 1 9 4 4 8 2 12 2 12 2
10 1 9 4 0 8 2 12 2 12 2
26 16 0 2 4 10 0 9 1 12 2 12 2 9 4 2 3 12 9 1 9 7 12 9 1 9 2
33 15 9 4 10 0 11 1 8 2 15 11 4 4 1 10 0 9 1 11 7 1 9 1 10 9 1 9 4 4 1 10 9 2
20 10 9 13 15 9 1 10 9 1 11 4 7 4 1 8 1 10 9 4 2
16 2 15 4 3 3 0 2 2 13 10 9 1 11 9 11 2
8 10 9 13 1 12 1 4 2
21 2 16 15 1 15 1 10 9 13 4 2 13 15 0 2 2 4 10 9 2 2
11 10 0 9 1 15 2 8 2 2 8 2
22 2 15 13 1 11 0 3 15 9 16 1 15 9 1 9 3 7 9 1 13 4 2
5 15 4 13 2 2
34 10 12 9 13 11 16 9 3 1 13 1 10 0 9 1 10 9 2 16 10 0 0 9 9 8 12 9 3 10 9 1 11 4 2
16 1 15 13 3 9 2 16 8 2 15 9 1 15 11 4 2
14 16 3 3 0 10 9 13 2 4 10 9 9 4 2
20 9 1 0 9 13 10 0 9 3 2 9 1 10 9 9 1 10 0 9 2
8 3 13 15 3 1 15 9 2
30 0 2 1 11 3 16 15 1 15 0 13 2 4 10 9 1 10 9 1 0 9 4 2 15 0 1 10 9 13 2
15 10 0 9 1 10 9 4 3 10 9 0 4 16 0 2
18 11 13 3 15 10 9 3 4 16 10 0 9 7 9 1 4 2 2
25 15 8 9 7 9 2 15 10 9 13 1 15 12 9 7 9 2 4 3 3 1 15 9 0 2
13 0 7 0 13 10 0 9 15 9 16 15 9 2
31 13 4 16 10 9 10 9 2 10 9 1 10 9 8 10 1 10 9 13 9 7 10 1 10 9 0 9 1 10 9 2
37 10 9 2 15 3 1 10 0 9 1 10 9 1 10 11 4 4 7 1 10 0 9 11 1 10 9 13 2 4 1 10 9 4 1 15 8 2
8 10 9 4 4 1 10 11 2
10 15 13 8 4 15 9 0 1 4 2
23 10 0 9 2 15 1 15 9 1 9 4 4 2 10 0 9 8 2 13 1 10 9 2
44 2 15 1 10 9 1 10 9 13 15 1 10 13 9 1 9 2 10 9 2 10 0 9 2 10 9 7 10 9 1 0 9 2 13 9 1 10 9 7 10 9 2 3 2
13 15 9 13 15 3 15 7 15 0 1 4 2 2
4 9 0 9 2
43 10 9 2 15 15 1 10 0 9 3 13 9 13 2 10 9 8 2 15 9 2 8 2 5 3 1 10 0 1 9 1 8 13 5 4 3 1 10 0 0 9 4 2
22 3 4 3 10 9 4 1 15 13 1 10 9 2 2 10 9 1 9 7 9 2 2
32 10 9 13 0 2 16 10 9 1 10 11 4 4 2 16 15 9 10 9 4 4 1 0 9 2 15 15 3 13 4 2 2
8 15 13 3 16 10 8 9 2
17 16 11 0 1 13 13 10 11 15 12 9 4 2 3 15 13 2
25 1 10 0 9 4 10 9 2 13 1 10 1 10 0 9 13 9 0 9 1 10 9 1 4 2
15 10 9 2 15 8 2 4 12 9 3 4 1 15 8 2
17 1 10 15 9 2 15 1 10 9 4 4 2 13 3 12 4 2
16 3 4 12 9 4 2 3 3 15 3 10 0 9 0 4 2
6 10 9 4 12 9 2
3 9 12 2
19 9 1 10 9 4 3 3 16 9 7 10 9 15 0 13 1 10 9 2
25 1 12 9 13 11 15 3 7 13 1 10 9 1 9 2 3 15 10 9 13 2 16 15 4 2
16 12 9 0 13 15 1 15 9 1 11 2 3 1 10 9 2
11 10 12 9 13 15 3 1 10 0 9 2
12 10 9 1 11 4 10 0 9 3 0 4 2
20 10 9 4 8 1 12 2 16 15 1 9 13 4 2 3 0 1 10 9 2
15 10 0 9 4 1 10 0 9 7 10 9 1 11 4 2
64 10 0 9 1 9 1 13 0 9 2 9 1 12 9 9 1 15 9 2 1 11 7 10 0 2 15 13 9 1 11 1 10 9 15 1 10 0 9 1 8 9 11 13 13 1 10 9 2 13 2 10 9 4 4 2 15 3 1 11 15 9 13 4 2
6 9 9 2 9 0 2
26 9 7 9 13 3 1 9 1 2 15 7 15 2 11 1 0 9 2 0 2 2 1 12 9 13 2
2 12 2
16 10 9 11 13 16 9 2 12 9 2 9 13 7 9 13 2
8 9 13 1 9 1 9 9 2
21 9 13 9 3 2 9 13 9 7 13 1 9 5 9 13 7 13 10 9 3 2
28 16 10 9 15 3 0 13 7 9 15 9 1 9 10 9 1 4 2 13 10 9 12 13 9 5 12 9 2
12 8 13 1 10 9 1 12 10 0 9 4 2
36 10 9 2 15 1 11 0 9 4 4 7 11 2 11 2 11 2 11 2 11 7 15 8 13 2 13 10 9 1 8 2 3 12 2 12 2
9 1 9 4 15 8 2 12 2 2
18 1 10 9 1 8 2 12 2 12 13 15 8 2 12 2 9 4 2
23 16 10 9 1 8 10 0 9 4 1 13 9 1 10 0 9 2 13 9 8 3 0 2
23 7 16 15 8 13 4 1 9 1 9 9 2 9 7 9 1 10 9 2 13 15 8 2
3 9 12 2
19 12 9 3 13 15 9 2 1 15 9 2 3 10 9 1 10 9 9 2
16 10 9 1 10 9 16 1 4 4 3 0 16 10 9 15 2
6 3 15 9 4 4 2
39 10 9 4 16 15 1 10 9 1 10 9 1 9 4 7 1 10 9 1 10 9 4 4 2 16 15 15 9 13 2 7 16 15 1 10 9 4 4 2
8 10 9 13 3 1 12 4 2
16 16 10 9 1 15 9 3 4 4 4 2 13 15 10 0 2
11 10 9 1 15 13 4 1 15 10 9 2
52 15 13 3 10 9 3 2 3 10 9 1 10 15 9 10 9 4 4 1 8 7 15 1 10 15 9 0 4 4 1 10 0 9 2 15 0 1 15 9 0 4 7 1 15 9 3 15 9 13 4 4 2
25 2 15 13 3 1 10 9 3 3 3 0 1 2 2 13 10 9 2 16 3 0 9 4 4 2
17 2 15 4 3 0 2 16 3 15 0 9 13 2 16 15 13 2
2 12 2
4 13 3 3 2
19 16 10 9 10 9 7 10 9 13 13 10 9 3 3 3 10 9 4 2
20 10 0 9 15 13 4 1 10 9 1 10 9 1 10 9 3 10 9 13 2
16 13 1 15 13 1 10 9 13 15 10 9 15 9 7 13 2
15 2 10 0 12 9 13 3 7 10 9 13 15 4 2 2
50 10 9 1 10 0 11 13 3 1 12 10 9 8 2 12 2 0 2 4 2 15 3 4 4 2 1 12 10 0 9 8 8 1 4 4 2 16 15 3 1 8 1 15 13 4 2 9 8 2 2
22 8 10 9 4 3 3 3 10 0 9 8 2 12 2 2 7 15 1 15 9 4 2
13 10 9 4 3 4 1 10 9 9 1 0 11 2
9 10 9 2 3 8 3 0 4 2
11 8 4 10 0 9 1 10 9 1 11 2
13 1 15 9 13 15 0 4 15 9 15 13 4 2
3 9 12 2
21 1 10 9 12 13 15 3 1 8 2 15 9 3 15 1 15 9 4 1 4 2
31 16 15 1 13 15 10 9 0 9 4 2 1 10 11 13 3 12 3 2 2 15 15 1 15 9 7 0 9 3 4 2
20 11 13 1 15 9 7 9 3 15 1 11 13 7 13 12 9 10 9 4 2
17 10 9 1 15 0 9 9 3 1 12 1 10 9 1 10 11 2
14 10 9 4 15 9 2 16 11 2 1 12 9 4 2
11 0 13 15 1 15 9 4 1 9 12 2
24 1 9 1 8 2 7 15 4 3 15 1 11 2 10 0 9 15 1 4 1 15 0 9 2
21 10 0 9 1 11 13 1 10 9 1 10 9 7 4 10 9 3 3 1 9 2
19 11 4 3 10 0 15 15 0 1 10 0 9 1 15 9 13 9 13 2
30 8 2 15 9 15 13 7 1 15 9 1 11 3 13 2 13 1 15 9 1 8 10 9 10 9 3 3 1 4 2
2 12 2
20 10 9 8 13 1 11 10 0 9 1 10 12 9 9 1 10 9 1 12 2
22 10 0 9 13 1 10 9 1 12 8 10 9 8 2 11 13 3 0 1 10 9 2
21 3 10 9 8 2 15 1 12 9 4 7 10 0 9 8 2 12 2 4 0 2
28 11 13 3 3 10 12 9 9 1 12 1 10 9 8 2 15 12 13 4 7 10 12 9 0 9 1 12 2
20 16 10 9 1 8 10 9 1 8 0 4 13 2 4 10 9 0 3 4 2
34 15 8 13 10 9 1 12 9 1 12 2 7 3 4 3 3 9 2 15 1 10 13 9 1 0 9 4 13 4 2 9 3 4 2
20 15 13 3 15 3 2 16 10 9 1 10 9 10 9 1 10 13 9 4 2
26 8 10 9 2 15 9 13 1 12 0 9 2 4 10 9 1 10 11 8 16 15 0 15 8 4 2
51 10 11 13 10 9 16 0 9 1 4 1 10 0 9 2 3 4 13 4 1 1 13 1 15 9 10 9 11 7 11 1 0 9 4 4 4 1 0 9 7 9 7 15 10 9 1 10 9 4 4 2
15 16 1 0 9 1 13 13 10 11 9 4 1 10 9 2
3 9 12 2
21 3 13 10 9 4 15 2 3 16 13 15 1 10 0 9 2 13 1 0 9 2
24 7 3 4 10 9 1 11 2 1 10 0 9 1 11 2 1 15 11 7 11 2 3 0 2
24 10 0 9 2 15 1 10 9 1 10 11 13 2 4 3 10 0 1 13 9 1 10 9 2
2 3 2
6 15 0 1 15 9 2
17 3 13 10 9 2 16 8 15 1 9 13 11 0 3 4 4 2
16 2 15 13 15 9 1 9 2 3 15 13 11 15 9 4 2
16 16 15 15 3 13 4 2 13 15 10 15 9 3 8 4 2
9 7 3 13 15 15 9 3 2 2
35 15 4 15 0 9 1 10 9 1 8 1 10 3 13 9 1 10 9 1 10 0 9 1 9 7 9 1 11 1 10 0 9 1 11 2
2 12 2
23 15 13 0 4 16 15 0 13 1 10 9 2 15 15 9 1 10 9 1 15 9 13 2
13 15 13 15 4 3 15 4 16 10 9 3 4 2
19 15 1 9 7 9 1 10 0 7 9 1 0 9 13 10 0 9 4 2
5 0 13 3 3 2
6 9 3 4 3 15 2
8 7 3 13 15 10 11 3 2
3 8 2 2
25 16 8 1 12 1 9 1 10 9 13 4 2 4 15 9 1 9 2 7 10 9 1 10 9 2
14 8 13 3 0 9 4 8 10 1 15 13 0 9 2
8 15 9 4 15 9 3 4 2
3 9 12 2
13 10 9 4 3 4 1 10 9 1 3 0 9 2
14 15 13 9 11 8 9 1 10 0 8 2 11 2 2
17 3 12 9 0 13 15 1 10 9 16 15 0 9 3 1 4 2
27 10 9 1 11 1 12 2 16 11 1 10 9 4 4 16 4 1 4 2 4 3 3 1 10 13 9 2
9 11 4 3 1 15 0 9 0 2
48 4 15 1 12 3 10 9 15 1 11 2 3 10 9 15 13 4 2 11 1 10 9 13 2 1 12 2 1 10 0 9 1 10 9 2 13 10 9 3 3 1 10 9 1 10 0 9 2
14 1 10 9 13 10 9 1 10 9 1 10 9 3 2
18 7 8 9 13 10 9 13 9 2 10 0 9 15 3 15 9 4 2
23 16 0 3 10 0 9 0 4 2 13 15 8 2 16 8 3 10 0 9 13 4 4 2
18 10 9 4 3 12 9 0 16 10 9 7 3 10 9 13 0 9 2
2 12 2
22 2 10 0 9 2 9 1 10 9 15 15 3 13 13 3 16 15 3 4 4 2 2
40 15 13 10 9 8 2 9 1 11 8 1 10 9 2 8 1 11 2 15 8 1 4 13 16 10 9 1 9 2 9 7 9 1 9 7 15 3 9 13 2
14 15 9 13 1 10 9 3 12 9 15 4 13 4 2
8 15 4 10 0 2 9 2 2
16 10 9 8 13 11 0 0 3 1 15 8 1 8 4 4 2
33 1 9 1 10 0 9 4 15 9 1 3 12 15 9 0 4 2 16 10 13 9 1 10 9 3 0 2 12 2 0 4 4 2
30 10 9 1 11 13 3 1 4 4 1 15 8 1 10 0 9 2 3 10 9 1 15 9 3 1 10 0 9 13 2
26 11 4 4 16 8 2 12 2 1 10 9 2 15 1 12 9 1 11 13 2 4 4 4 7 3 2
27 11 0 9 1 9 1 15 9 5 7 3 0 9 1 10 12 9 4 0 4 1 10 9 1 10 9 2
8 1 11 13 15 3 1 9 2
18 1 9 13 10 9 1 10 0 9 7 9 1 3 12 7 12 9 2
12 15 13 3 15 9 7 13 3 15 9 3 2
52 0 9 4 3 1 10 0 9 3 10 9 2 16 10 9 1 11 4 4 2 16 10 13 9 1 15 9 1 10 9 11 3 12 12 9 1 9 4 2 15 4 1 11 10 9 1 3 10 16 12 9 2
16 8 13 10 0 9 1 12 2 15 4 12 9 15 16 11 2
6 3 8 4 3 0 2
35 10 0 9 8 1 11 7 15 0 0 9 8 1 11 13 1 10 0 9 0 1 12 0 1 10 9 1 8 1 11 8 1 4 4 2
10 3 4 9 8 1 10 9 0 4 2
10 10 9 13 2 16 10 9 0 4 2
20 3 1 10 9 2 15 12 9 13 4 2 13 15 16 10 9 11 4 4 2
10 15 0 8 13 10 9 3 0 13 2
33 1 10 9 11 7 1 15 2 0 2 9 13 10 9 10 9 1 10 13 9 1 10 9 1 10 11 13 11 1 10 0 9 2
21 10 9 2 10 0 9 2 13 1 9 2 16 15 10 0 9 1 15 9 13 2
12 10 9 1 10 9 13 3 4 1 10 9 2
18 16 15 13 1 10 9 13 9 11 7 9 11 15 1 10 9 4 2
12 15 13 3 3 3 2 3 15 3 4 4 2
15 15 13 15 3 1 2 9 2 2 10 9 1 10 9 2
12 1 15 9 13 3 3 9 4 1 0 2 2
51 10 9 2 15 1 11 3 10 9 1 12 9 13 5 3 10 9 13 8 10 9 2 10 15 13 5 13 3 10 9 1 10 9 1 9 1 0 2 0 2 7 3 15 15 3 13 4 5 9 9 2
28 15 10 9 1 9 1 9 2 9 7 9 1 13 9 13 4 2 16 15 8 13 4 2 4 3 3 0 2
23 3 3 15 9 2 15 8 1 11 1 11 2 9 1 9 13 2 4 15 10 0 9 2
15 1 15 9 13 15 9 2 9 2 9 2 0 9 3 2
12 15 1 10 9 4 3 4 7 1 9 4 2
35 2 15 13 10 15 0 9 9 16 1 10 9 13 7 3 13 15 3 2 1 10 0 9 1 2 15 9 3 4 4 2 13 15 0 2
26 3 4 3 3 9 4 16 15 9 0 1 4 7 15 1 4 4 15 3 1 15 0 9 4 4 2
49 15 4 3 0 9 1 11 2 1 13 9 7 9 5 15 0 3 0 5 1 10 0 13 9 2 3 10 9 11 1 9 1 4 4 2 7 1 10 0 9 2 9 2 1 0 9 1 9 2
20 0 10 0 9 9 1 10 0 9 8 2 15 3 10 9 8 13 1 9 2
30 11 13 0 1 10 9 2 1 10 9 1 10 16 12 9 1 9 15 1 3 3 3 0 9 1 9 13 4 4 2
16 15 13 10 9 1 11 1 11 1 12 9 7 12 9 4 2
10 10 0 9 13 3 3 12 9 0 2
7 10 9 4 1 11 4 2
13 1 10 9 1 11 13 10 9 3 15 13 4 2
5 3 13 10 9 2
46 10 9 1 10 0 9 2 1 13 13 15 10 9 1 10 9 4 7 9 15 15 3 13 1 4 13 16 15 9 8 4 2 13 1 10 13 9 3 4 1 11 2 11 7 11 2
22 3 4 10 9 0 16 1 10 0 9 10 0 9 13 2 3 15 3 15 3 13 2
17 1 11 4 0 16 15 10 9 3 13 1 15 13 1 0 9 2
22 9 11 13 10 0 9 11 4 15 1 9 1 9 0 3 3 1 4 16 1 11 2
25 15 13 1 10 9 15 10 9 1 10 0 9 3 1 10 0 9 1 11 1 10 9 13 4 2
16 10 9 1 11 4 16 15 1 11 13 9 3 8 1 13 2
9 1 11 13 8 1 9 12 4 2
15 1 10 9 9 13 8 2 9 2 1 10 9 4 4 2
9 8 13 3 1 10 9 1 12 2
65 2 3 4 3 4 1 10 0 9 3 9 3 1 10 0 9 10 9 1 13 7 13 9 7 1 10 9 13 4 2 7 16 9 4 4 2 16 10 9 9 3 0 13 4 4 7 3 16 10 0 9 8 15 10 13 2 0 7 0 9 13 4 4 2 2
26 3 12 9 1 10 12 1 12 7 12 1 11 7 11 0 9 2 13 9 15 15 1 11 0 4 2
21 15 4 10 0 9 16 10 9 1 10 0 0 9 3 10 9 1 10 9 4 2
24 13 10 9 2 15 15 13 2 3 3 3 4 2 3 13 15 1 10 0 9 1 15 4 2
20 1 9 13 15 15 9 4 2 7 3 13 15 0 3 3 15 3 4 2 2
14 15 12 9 13 1 12 9 9 15 1 11 4 0 2
36 12 9 1 10 9 13 1 11 7 11 2 12 9 1 11 2 12 9 1 15 9 7 12 9 1 2 15 9 2 2 3 11 7 15 8 2
33 15 13 1 15 9 1 15 13 1 10 9 4 4 16 10 0 7 0 9 15 1 15 15 9 1 4 4 2 3 10 9 11 2
28 15 13 3 16 10 9 1 0 9 1 10 9 3 3 4 16 10 9 0 4 3 1 15 9 3 1 4 2
21 15 9 4 0 16 10 9 15 3 13 4 7 15 1 10 0 9 13 4 4 2
33 1 15 1 10 0 9 1 10 2 9 2 2 15 15 1 9 13 4 4 2 13 10 9 1 9 1 10 9 7 1 10 9 2
20 7 11 0 9 2 3 15 9 13 7 13 2 4 10 0 9 1 10 9 2
20 10 9 1 11 13 1 9 1 3 12 12 9 3 2 15 15 4 13 4 2
30 7 1 10 0 9 3 10 0 9 1 10 16 12 12 2 16 1 10 0 12 9 1 12 3 15 12 9 4 4 2
33 0 9 13 15 3 7 1 15 0 9 3 4 4 16 9 1 10 0 9 7 3 1 3 10 16 12 9 0 9 1 10 9 2
18 7 9 2 3 15 0 3 3 3 13 4 2 4 15 3 3 0 2
24 15 13 3 16 11 15 1 15 0 0 15 0 9 10 0 9 1 10 9 4 1 4 4 2
39 3 13 10 13 9 1 10 11 1 10 9 1 10 9 1 9 4 1 10 9 1 10 0 9 2 16 1 15 9 10 9 1 11 7 11 13 4 4 2
21 10 9 4 3 4 1 15 9 16 15 1 10 0 9 10 9 7 9 4 4 2
32 1 11 13 15 3 3 3 16 15 0 13 2 9 11 1 9 11 7 3 11 1 9 11 2 3 1 11 1 11 4 4 2
14 10 11 1 11 13 3 3 10 9 1 10 9 4 2
9 9 4 8 9 1 10 13 9 2
13 1 15 13 8 2 8 8 7 8 1 15 9 2
23 16 15 3 13 4 13 10 11 7 10 11 1 11 1 10 13 9 4 1 10 9 8 2
28 1 9 4 4 10 9 1 12 9 8 1 15 9 1 4 1 13 1 10 9 1 10 11 8 10 9 8 2
32 8 10 9 16 10 9 3 1 10 9 1 10 9 1 4 13 15 3 10 3 0 0 9 4 4 15 11 9 3 13 4 2
11 15 13 3 16 15 3 10 9 4 2 2
26 1 15 9 4 4 16 9 11 10 0 0 9 1 10 15 9 1 9 1 11 9 3 4 4 4 2
30 7 16 15 3 2 8 10 0 9 2 10 3 1 10 9 15 0 9 0 1 10 0 9 10 9 13 4 4 4 2
16 15 9 1 9 3 4 3 1 4 1 11 0 9 0 9 2
4 15 13 4 2
60 15 9 1 9 13 15 3 3 1 10 0 9 2 16 3 3 3 0 0 2 7 3 13 15 1 15 13 1 0 0 9 2 10 0 9 2 2 16 3 0 1 13 16 10 9 1 10 9 1 10 9 2 0 9 2 4 1 4 2 2
17 7 15 9 1 9 13 3 10 9 1 0 0 9 2 10 0 2
36 1 10 9 8 1 10 9 1 11 0 4 10 13 9 4 2 15 10 9 13 4 4 16 1 10 11 10 9 11 10 0 9 8 4 4 2
6 10 0 9 13 4 2
34 2 10 15 0 9 4 11 4 2 1 15 10 0 9 8 2 0 1 10 0 9 2 3 10 0 9 1 10 0 9 13 4 2 2
39 9 11 2 15 13 13 4 16 15 3 3 13 9 15 15 9 4 13 2 13 15 3 3 7 1 15 0 9 7 0 9 2 13 15 11 3 15 9 2
14 2 13 15 16 1 10 9 12 10 9 4 4 2 2
22 16 13 11 16 1 10 9 1 10 9 2 15 15 13 1 10 9 4 3 3 0 2
24 3 13 9 11 1 9 10 13 11 4 7 13 8 10 1 11 13 9 3 3 1 10 9 2
39 9 8 2 15 1 15 0 13 3 1 11 2 13 10 9 1 10 9 1 10 9 16 10 9 11 15 9 4 7 16 10 9 2 15 3 3 4 2 2
31 3 13 8 3 1 13 16 15 1 10 11 10 9 1 9 1 11 4 4 16 15 9 10 0 0 9 9 13 4 4 2
14 10 11 4 3 10 9 13 1 10 9 8 1 8 2
11 9 8 1 11 13 7 13 15 3 4 2
22 8 13 1 12 10 13 9 1 15 9 4 7 3 3 10 9 4 1 10 9 9 2
12 10 9 1 10 9 13 15 13 1 10 9 2
9 7 13 1 10 9 4 11 15 2
14 2 15 13 10 0 9 2 15 3 10 9 13 4 2
5 15 13 7 13 2
14 13 15 9 1 11 2 15 13 0 3 15 0 4 2
13 10 9 4 0 1 7 0 1 15 15 9 4 2
12 3 12 9 1 9 13 8 10 13 9 4 2
18 11 13 10 0 9 1 10 9 1 9 1 11 1 10 9 1 8 2
14 11 13 1 10 0 9 10 9 1 12 1 11 4 2
17 11 13 1 11 10 9 2 7 1 10 9 1 11 4 15 12 2
16 1 10 9 13 11 3 1 9 1 11 2 12 2 7 11 2
13 3 4 10 9 1 15 9 1 15 9 0 4 2
18 8 13 16 15 10 13 9 1 9 0 4 4 4 3 1 4 4 2
15 10 9 13 9 3 1 4 16 15 10 9 3 1 13 2
8 2 4 10 9 3 3 4 2
10 1 10 9 15 13 13 15 0 9 2
21 2 15 13 10 9 1 4 2 16 15 3 15 9 4 16 15 3 1 9 4 2
20 9 11 13 1 11 4 16 15 9 1 10 11 3 1 13 4 1 10 9 2
17 15 4 2 13 15 2 15 9 2 16 15 3 3 15 13 4 2
18 15 4 10 0 0 9 1 0 9 15 10 0 9 1 10 11 13 2
20 15 13 3 10 9 1 0 0 9 1 10 11 2 3 9 1 10 0 9 2
8 3 13 15 1 11 7 11 2
10 10 9 1 8 13 3 0 9 4 2
28 16 15 8 11 10 0 9 4 4 2 13 10 9 3 1 10 0 9 1 10 9 1 10 0 9 0 3 2
11 10 9 13 3 1 3 12 9 1 3 2
25 15 13 16 16 15 3 10 0 9 13 1 10 9 1 9 2 0 9 2 15 3 9 4 4 2
27 1 10 0 9 1 10 9 13 10 9 0 9 3 2 3 10 9 13 4 1 10 9 1 0 12 9 2
20 9 8 2 12 2 1 10 9 11 13 3 3 3 1 10 9 1 15 8 2
35 7 15 13 10 9 1 15 9 2 7 15 1 15 3 13 2 7 0 9 2 16 15 3 12 9 3 13 4 2 4 1 11 1 4 2
4 1 10 9 2
36 15 4 15 0 2 0 2 8 2 2 15 15 1 12 13 7 1 12 1 9 13 1 9 11 1 10 0 11 1 10 9 1 10 0 9 2
12 15 13 3 15 9 3 0 8 4 1 4 2
15 15 13 15 10 9 1 10 9 2 15 15 13 4 4 2
21 11 7 15 4 8 2 16 15 15 9 16 9 1 10 9 1 13 9 4 4 2
9 15 13 15 9 0 0 1 4 2
8 1 15 0 9 13 8 3 2
36 10 9 11 13 0 0 16 10 9 1 8 10 9 0 0 4 2 1 15 9 15 0 16 10 9 1 11 2 3 8 15 9 3 13 4 2
28 2 3 15 2 11 2 1 10 9 1 10 9 13 2 4 15 15 0 15 15 15 4 4 15 9 1 13 2
17 0 4 15 13 16 10 9 1 13 2 7 10 9 3 4 0 2
10 15 13 3 3 9 1 0 9 4 2
12 15 13 1 10 9 2 2 3 10 9 11 2
9 3 9 13 10 9 1 10 9 2
22 10 9 13 1 0 9 1 3 2 7 10 0 0 9 4 0 1 10 9 1 4 2
20 3 13 15 10 9 1 10 9 4 2 3 0 4 4 0 0 9 1 4 2
9 10 9 2 8 2 13 3 4 2
22 10 9 2 3 9 1 10 9 1 9 9 10 9 2 4 3 1 9 7 1 9 2
16 10 9 4 1 10 9 1 8 1 10 13 9 4 1 11 2
23 2 15 4 16 3 8 16 10 9 11 13 7 3 4 15 0 1 15 1 10 9 4 2
12 10 9 13 1 10 9 1 9 11 1 11 2
7 15 13 15 9 9 3 2
11 2 15 13 15 3 2 2 13 15 3 2
11 15 9 4 2 13 15 10 0 9 2 2
9 3 13 10 11 3 3 10 9 2
27 16 11 7 11 12 9 10 0 9 1 11 13 4 2 4 15 3 4 1 10 9 2 13 1 15 8 2
20 15 13 3 9 1 10 2 9 2 2 9 2 15 10 9 13 8 1 4 2
19 12 9 3 13 1 10 9 2 16 12 1 12 1 15 9 0 13 4 2
23 16 15 1 10 9 13 2 4 15 1 15 9 4 7 4 15 4 1 10 9 0 9 2
21 15 4 10 0 9 2 7 8 13 3 4 16 15 1 10 0 2 0 9 4 2
37 10 9 13 15 3 16 1 15 9 3 15 9 3 1 4 7 15 13 3 15 9 2 10 9 8 2 15 9 4 2 2 3 13 10 9 11 2
30 7 1 10 9 13 15 3 3 9 7 9 1 8 2 15 15 0 9 4 2 3 3 15 9 13 7 0 13 4 2
12 15 4 15 3 3 16 10 0 9 1 13 2
42 10 0 9 1 9 13 3 1 10 0 9 1 12 2 9 2 2 10 0 9 8 7 10 0 9 8 2 12 9 9 4 1 15 13 1 10 9 9 7 0 9 2
29 10 9 4 4 1 10 9 1 10 11 2 15 1 15 9 2 1 10 9 2 0 4 9 1 15 9 1 4 2
15 11 13 10 9 2 16 15 15 9 4 16 0 1 4 2
8 11 13 3 15 8 4 4 2
15 10 9 15 3 3 2 7 15 4 3 15 0 1 4 2
53 13 1 10 9 16 11 1 11 13 4 2 13 10 9 10 9 1 10 9 3 3 3 3 16 13 9 7 4 15 1 10 9 3 1 4 2 16 3 15 9 1 10 9 4 16 15 15 11 1 10 9 13 2
12 8 4 10 9 1 10 0 11 9 1 11 2
31 15 9 13 1 10 16 13 9 4 2 7 1 10 9 13 15 9 10 9 1 10 9 1 10 0 9 1 10 0 11 2
40 8 1 11 4 1 8 2 3 15 10 0 9 1 15 8 1 12 9 1 8 13 7 3 8 10 9 8 13 2 3 3 10 3 13 9 1 10 0 9 2
12 10 9 1 8 13 15 7 13 10 9 9 2
12 2 15 13 9 2 13 9 8 15 0 3 2
23 2 11 13 9 2 2 13 8 7 10 9 1 15 0 9 4 1 15 9 1 0 9 2
14 0 3 7 1 11 10 0 9 16 15 1 4 4 2
14 3 10 9 3 15 15 3 0 1 10 9 4 4 2
17 15 13 15 1 15 9 4 1 15 11 2 10 0 9 2 13 2
12 2 16 11 15 13 13 15 1 15 9 2 2
8 15 13 11 4 8 1 11 2
34 2 10 9 4 10 0 9 2 2 13 10 9 1 8 2 15 15 3 13 4 2 7 15 13 1 11 15 9 11 3 1 15 9 2
22 15 13 3 3 7 10 9 1 10 0 9 13 3 1 10 9 1 10 9 1 4 2
35 8 2 1 8 7 8 9 1 10 0 9 2 12 9 2 13 10 0 12 9 4 16 15 3 1 10 9 1 15 9 1 10 9 4 2
16 15 8 13 12 1 10 9 3 1 10 9 0 1 13 4 2
21 15 4 3 3 0 1 10 9 2 1 12 9 2 2 16 15 15 9 4 4 2
12 10 9 15 3 3 10 9 13 4 4 8 2
33 2 15 13 15 9 3 3 16 15 4 13 2 3 0 9 13 15 10 9 2 2 13 8 2 9 1 10 3 0 11 0 9 2
28 7 1 15 9 13 13 15 15 0 0 2 7 3 13 15 9 2 10 15 9 1 3 0 9 16 10 15 2
24 15 9 4 10 9 1 8 1 10 11 4 7 1 10 9 4 10 0 9 7 10 9 4 2
20 12 9 13 4 15 9 7 10 9 15 1 10 0 9 4 4 16 15 8 2
11 15 9 4 3 3 3 0 16 0 9 2
28 3 13 3 1 11 12 9 15 15 9 9 1 10 0 9 1 12 9 5 15 9 1 13 9 5 13 4 2
28 1 10 9 13 10 9 10 9 3 1 10 9 15 0 8 13 7 16 15 1 10 9 4 2 3 3 13 2
42 10 9 1 11 4 4 1 8 2 15 1 11 1 10 0 9 2 0 4 7 10 0 9 1 8 1 11 2 10 0 1 8 1 11 7 10 0 1 8 1 11 2
11 10 9 4 0 0 2 3 12 12 9 2
17 10 9 2 15 3 10 9 1 11 1 9 1 10 9 3 13 2
21 10 9 13 3 12 9 1 11 2 15 3 3 10 9 1 12 9 13 1 4 2
7 2 10 9 13 0 0 2
7 15 13 15 15 9 2 2
54 15 4 10 0 9 1 9 8 2 15 1 15 0 9 1 11 1 10 0 9 1 10 0 1 10 0 9 13 2 7 3 1 10 9 9 10 0 9 13 1 10 0 9 1 10 0 11 1 10 9 11 3 9 2
19 13 7 13 1 9 9 7 9 2 13 15 3 3 0 10 9 8 4 2
3 3 9 2
39 0 4 15 15 10 0 9 1 9 2 3 15 13 1 10 0 9 2 7 3 15 0 7 13 4 2 13 15 3 3 15 3 1 4 2 1 15 9 2
7 0 0 13 8 3 13 2
7 13 9 8 2 8 2 2
21 13 9 13 8 1 12 2 8 2 7 8 1 12 2 8 2 2 1 0 9 2
19 1 10 9 13 15 10 0 9 4 2 3 15 0 1 15 0 3 13 2
19 3 13 11 3 0 9 7 10 9 13 3 7 3 3 3 1 12 9 2
15 10 9 13 15 0 1 10 11 1 10 9 1 10 9 2
26 15 13 8 1 15 2 8 3 1 11 7 11 2 3 10 0 9 3 3 0 4 2 10 0 9 2
34 2 15 4 2 9 2 1 15 0 9 3 2 13 1 15 0 0 9 2 0 1 10 9 2 10 0 9 3 15 15 13 2 2 2
14 11 2 2 8 2 8 2 5 12 9 2 12 9 2
47 15 13 15 3 4 1 15 0 2 1 10 9 13 9 2 13 9 2 0 2 0 13 9 2 9 0 3 1 10 9 2 7 15 1 10 9 10 9 13 2 10 9 3 1 15 13 2
18 8 13 15 9 1 3 12 9 2 15 15 1 9 1 0 11 13 2
26 3 4 3 3 12 4 2 16 3 15 9 3 1 11 7 1 10 9 1 11 1 10 9 13 4 2
14 3 13 0 9 1 4 2 7 15 4 10 9 3 2
9 1 8 13 1 9 12 9 3 2
8 7 10 9 4 0 1 0 2
31 13 0 3 4 8 2 15 16 11 10 9 9 13 1 11 7 10 9 1 10 9 2 1 11 7 10 9 1 10 9 2
8 13 11 15 8 3 4 4 2
33 1 10 9 1 15 13 2 0 13 8 2 1 8 2 4 1 15 0 13 10 9 1 11 4 1 10 9 0 0 9 8 8 2
21 15 13 8 7 8 16 15 9 7 13 3 1 10 9 1 8 3 1 9 3 2
10 11 4 0 1 10 0 9 13 4 2
35 13 15 1 15 9 1 9 11 10 0 9 1 15 4 8 15 8 2 15 13 10 9 16 15 3 4 16 15 3 8 11 15 3 4 2
23 15 13 3 2 11 2 1 11 4 7 13 0 15 9 4 15 8 1 10 9 13 4 2
17 15 9 13 15 0 2 3 1 9 2 1 15 9 3 4 4 2
18 10 13 9 7 10 9 15 13 1 13 9 4 15 15 0 13 4 2
12 0 4 1 10 9 11 12 9 0 1 12 2
19 3 1 10 0 9 0 1 10 9 15 7 10 9 15 15 9 13 4 2
9 15 13 16 16 9 15 3 0 2
32 15 13 10 9 3 1 10 9 3 7 15 13 0 1 10 9 1 10 9 15 3 1 11 1 15 9 8 4 13 4 4 2
34 10 0 9 8 2 15 9 1 10 0 11 13 7 15 0 9 1 10 3 1 10 9 13 0 9 11 13 13 1 11 0 9 4 2
19 16 15 15 9 3 13 4 15 15 3 4 1 4 1 10 0 9 8 2
23 10 9 8 2 15 10 13 9 10 9 1 15 1 11 13 4 2 13 1 10 0 9 2
7 10 12 9 4 0 9 2
23 10 9 7 10 13 9 1 8 2 7 10 0 0 9 1 10 9 10 9 12 1 11 2
14 3 13 15 9 3 15 3 15 9 1 11 11 4 2
13 10 3 13 9 1 0 9 2 16 15 9 8 2
17 10 11 1 11 13 15 2 16 9 2 1 13 9 4 1 8 2
19 8 13 15 0 9 3 4 2 3 3 1 8 3 2 8 2 4 4 2
10 0 4 15 3 2 3 4 15 3 2
30 10 9 4 3 0 13 1 4 2 3 3 10 9 1 15 8 1 10 0 9 12 9 0 4 16 1 15 9 12 2
19 15 13 4 4 16 10 9 1 15 8 10 9 1 3 10 11 4 4 2
31 7 10 9 8 1 10 9 1 11 7 11 13 10 3 0 9 1 4 2 16 10 9 0 1 0 13 9 13 4 4 2
13 1 15 8 2 0 1 11 2 13 10 0 9 2
9 1 10 9 2 11 11 2 13 2
19 15 13 3 9 0 7 10 9 13 2 1 11 2 3 9 1 9 4 2
49 10 9 1 10 0 9 11 7 8 2 10 9 7 9 8 13 1 15 1 15 9 10 9 4 15 0 9 2 15 0 1 10 0 9 13 2 1 4 7 3 10 2 0 9 2 3 1 4 2
57 11 13 3 3 0 1 10 9 2 4 4 1 10 15 9 2 13 13 1 10 9 2 13 3 1 10 13 9 15 13 2 13 10 9 1 3 7 13 15 1 10 9 1 3 2 3 10 9 1 10 9 1 10 13 9 13 2
14 1 12 4 10 9 1 15 0 9 4 1 10 11 2
5 10 9 4 13 2
28 9 8 2 12 2 1 11 2 15 10 0 9 1 9 1 10 9 8 1 8 13 2 4 3 0 4 4 2
38 10 9 2 10 9 3 10 9 1 10 9 0 13 2 4 1 11 15 16 15 13 4 4 16 10 9 10 9 1 13 1 9 1 10 9 1 4 2
19 10 9 4 3 0 4 2 16 1 10 9 10 9 1 10 9 0 4 2
20 1 11 12 9 2 1 11 12 9 2 1 11 12 9 7 1 11 12 9 2
16 3 13 15 16 10 9 10 9 1 15 9 1 15 9 4 2
17 10 9 13 15 4 1 10 9 2 15 9 13 4 1 10 9 2
16 1 10 9 4 10 9 1 10 9 3 4 2 7 0 4 2
17 10 9 13 16 1 10 9 1 10 15 9 0 9 13 4 4 2
11 3 13 15 10 0 9 1 15 9 3 2
21 10 9 13 1 10 9 8 7 10 9 4 4 1 10 11 1 11 1 12 9 2
6 0 4 15 10 9 2
33 13 16 10 9 15 9 4 4 4 13 10 9 10 9 1 15 9 0 1 10 9 1 10 9 2 3 15 3 0 1 9 13 2
11 1 10 13 9 13 15 9 1 10 9 2
6 9 13 3 3 3 2
12 10 9 1 10 11 1 11 13 1 8 0 2
34 1 15 9 1 9 13 1 4 2 3 10 9 15 1 9 10 0 9 4 2 3 3 3 4 4 2 3 10 11 1 15 9 4 2
18 15 13 10 9 1 10 9 2 3 1 9 1 15 9 2 3 3 2
18 7 15 13 15 0 10 9 1 15 0 9 2 16 15 1 15 13 2
6 10 9 3 13 15 2
16 2 1 12 2 16 10 9 9 4 2 4 3 3 15 4 2
3 12 9 2
46 9 8 1 8 13 9 8 1 11 7 9 8 9 1 10 9 1 8 4 1 10 9 1 4 4 2 16 10 9 1 11 1 10 0 9 15 9 1 13 16 1 10 0 9 2 2
32 2 10 9 13 3 1 10 9 2 2 13 9 8 3 1 10 9 1 10 9 1 10 9 8 9 2 1 10 0 9 13 2
8 15 4 3 8 1 10 11 2
14 3 4 10 9 2 3 15 0 13 1 10 0 9 2
30 15 13 10 11 1 10 11 2 16 10 11 9 11 10 9 13 2 3 4 4 1 0 7 13 9 1 10 0 11 2
4 10 11 13 2
17 2 15 13 10 9 3 2 16 3 4 4 1 10 9 1 9 2
41 15 0 9 1 10 9 1 3 4 10 0 9 1 10 11 11 2 10 9 1 0 9 2 3 13 1 8 7 8 2 3 8 10 9 1 10 0 9 0 13 2
32 10 9 2 3 8 2 10 13 9 1 8 2 15 13 16 11 15 0 9 7 9 4 10 9 4 4 4 2 0 0 2 2
12 10 0 15 15 3 13 4 4 10 9 15 2
25 1 15 9 4 15 9 3 3 3 1 4 2 7 10 9 1 11 4 3 15 15 15 0 13 2
8 8 2 9 1 10 9 13 2
22 16 10 9 3 3 1 10 9 11 4 4 2 4 10 9 11 3 3 1 10 9 2
5 1 10 9 13 2
23 2 2 13 1 9 1 4 4 16 15 9 1 10 9 3 1 15 3 10 0 9 4 2
10 3 13 15 9 3 3 4 4 2 2
17 10 9 13 3 1 10 0 9 1 10 9 2 3 1 10 9 2
10 10 9 13 15 3 8 8 3 3 2
28 15 13 0 2 16 15 10 9 2 15 10 9 1 13 7 15 10 0 9 10 9 1 9 15 9 4 4 2
26 10 9 8 2 9 2 13 2 16 3 9 4 4 4 16 9 1 4 1 10 0 9 1 10 9 2
32 16 10 9 13 1 10 9 2 13 1 15 3 1 10 0 9 4 4 2 2 3 13 3 3 3 3 10 0 9 3 2 2
13 1 11 13 10 9 3 10 9 1 15 9 4 2
11 2 1 8 13 15 4 4 1 15 9 2
8 7 10 9 4 3 0 9 2
29 3 2 10 9 13 1 10 9 1 10 9 0 9 4 1 10 9 1 10 9 2 15 0 13 4 1 10 9 2
45 4 3 3 10 9 2 16 3 10 0 9 1 10 9 4 13 4 2 0 4 3 3 10 9 3 4 1 10 9 2 10 1 9 13 9 13 3 15 15 1 10 9 3 2 2
13 15 4 3 0 16 8 1 11 1 11 13 4 2
32 10 9 4 3 0 9 8 2 7 10 0 9 3 11 13 2 8 1 11 2 13 10 9 3 0 16 11 3 3 13 4 2
24 3 13 10 9 15 9 3 4 2 16 9 1 11 3 1 11 13 16 10 9 3 1 13 2
9 15 13 0 9 1 9 1 4 2
28 10 9 1 11 13 3 1 12 1 10 9 1 10 11 10 0 9 4 1 10 9 8 2 12 2 1 11 2
6 10 9 9 1 9 2
13 9 4 15 1 9 4 1 15 9 1 10 9 2
5 3 4 15 0 2
21 0 4 10 9 8 2 16 15 1 10 9 13 2 0 4 7 1 10 9 4 2
10 15 13 3 10 0 9 3 4 4 2
9 3 3 4 15 0 13 9 4 2
22 12 9 2 8 1 11 7 8 1 11 2 15 9 0 13 4 1 10 9 1 11 2
32 10 1 10 9 11 13 9 13 15 9 2 16 15 1 10 9 1 11 13 2 3 8 1 11 15 3 13 7 10 9 13 2
31 16 10 0 9 8 1 11 11 1 10 9 11 1 11 15 9 13 1 10 0 9 8 2 3 1 11 2 13 10 9 2
44 1 9 13 3 15 0 2 16 2 8 10 10 9 2 15 9 15 13 2 13 2 1 15 10 9 16 15 1 15 9 15 13 1 10 0 9 2 9 13 2 3 15 13 2
16 15 3 13 10 9 15 15 0 9 0 1 4 7 1 4 2
29 3 0 4 15 9 1 0 9 1 10 9 13 7 15 3 9 4 4 1 10 9 7 9 2 8 2 1 13 2
46 10 9 1 10 0 9 13 10 0 12 9 8 4 10 13 9 8 1 4 16 1 0 9 9 1 13 1 0 9 1 10 9 7 10 9 1 10 0 9 1 10 0 9 7 9 2
2 11 2
28 1 10 13 9 5 8 0 5 4 10 9 4 1 10 9 3 15 15 15 3 0 1 3 13 2 13 4 2
12 9 7 4 2 9 7 9 2 13 7 0 2
25 10 9 15 10 9 3 13 4 2 4 10 9 1 9 1 10 9 1 10 9 1 10 0 9 2
17 10 9 1 10 9 4 1 10 0 9 1 12 9 0 0 4 2
7 3 13 10 9 8 9 2
32 10 9 4 0 2 7 3 4 0 4 2 16 10 9 3 0 16 12 9 4 4 7 16 15 3 15 0 9 3 4 4 2
10 3 4 8 0 4 1 3 15 9 2
5 11 13 0 0 2
17 15 13 15 15 9 3 0 4 4 2 7 3 4 15 3 0 2
8 3 4 3 15 9 3 2 2
7 2 3 4 15 10 9 2
29 11 8 2 3 15 13 16 9 15 16 15 1 15 0 4 2 13 2 16 3 1 8 3 3 10 9 4 4 2
13 2 15 13 3 3 15 9 4 2 2 3 11 2
11 2 7 3 4 1 15 15 3 15 4 2
7 11 13 15 10 0 9 2
25 10 9 4 0 3 0 15 0 2 7 13 3 15 9 16 10 0 0 9 1 0 9 1 4 2
14 10 0 9 8 2 11 2 11 7 11 13 3 0 2
15 11 13 0 8 7 3 1 10 0 9 13 10 9 8 2
7 11 13 0 1 10 9 2
27 10 13 9 4 1 8 0 4 7 1 10 0 0 9 13 15 10 9 0 1 10 0 9 2 12 2 2
15 9 11 7 11 13 10 12 9 10 0 7 0 9 3 2
7 9 13 15 3 3 3 2
18 16 11 3 1 10 12 9 3 4 13 15 1 4 1 15 0 9 2
19 3 4 10 9 10 3 1 13 9 2 3 10 9 1 11 3 4 4 2
15 10 9 13 1 10 0 9 10 9 1 11 2 12 2 2
18 1 10 9 13 11 10 9 3 0 0 1 10 0 9 2 12 2 2
28 9 8 1 11 13 3 3 3 4 16 8 2 11 1 10 9 1 8 9 13 2 9 1 8 4 4 4 2
14 2 8 2 15 15 9 15 13 4 2 4 3 4 2
6 15 4 3 3 13 2
22 0 13 15 2 16 15 11 13 2 10 9 0 16 1 13 7 15 13 15 4 2 2
9 10 9 13 3 1 10 9 3 2
22 1 10 0 9 13 15 0 8 1 8 3 10 9 1 10 0 13 9 1 11 4 2
10 15 4 10 9 15 1 10 9 4 2
26 3 1 10 0 9 13 15 9 10 9 7 13 15 1 0 9 1 8 7 11 1 10 9 1 4 2
7 10 9 8 13 3 3 2
27 3 13 8 15 1 10 9 1 0 9 7 10 9 13 3 0 3 1 10 9 7 15 13 10 0 9 2
16 1 10 9 1 9 8 1 11 4 15 9 10 0 9 4 2
14 11 4 10 9 11 8 4 8 0 9 1 10 9 2
21 15 9 1 8 4 3 4 1 8 2 15 0 3 1 8 10 9 1 11 13 2
23 9 8 1 15 8 2 15 10 9 1 11 0 1 10 9 1 11 13 2 13 1 9 2
19 2 11 13 10 9 1 10 9 1 15 9 1 9 1 9 1 10 9 2
35 1 10 9 13 8 2 9 1 15 8 2 16 0 13 3 4 4 1 10 0 9 2 7 1 10 9 9 2 10 9 9 1 10 9 2
15 15 13 2 16 10 9 15 9 3 4 1 10 0 9 2
2 0 2
26 2 10 9 9 2 2 3 8 2 2 4 0 15 0 16 15 7 13 3 1 4 1 10 9 2 2
5 15 13 3 3 2
23 2 1 0 13 2 9 7 8 2 10 9 13 9 2 9 2 4 1 15 9 15 9 2
43 1 0 0 9 2 16 3 1 10 9 3 4 4 4 2 15 13 15 9 3 9 3 1 3 10 0 9 2 4 15 0 4 1 10 9 2 15 3 12 9 3 13 2
19 15 4 8 4 15 2 1 15 15 3 13 9 0 2 9 3 1 4 2
19 0 9 13 3 3 0 9 1 9 2 16 15 8 15 3 0 4 4 2
29 3 13 15 10 0 9 1 10 9 2 15 9 13 1 10 9 2 15 15 1 10 9 1 15 9 1 12 13 2
16 1 15 9 13 15 10 0 9 9 3 2 3 10 1 11 2
25 16 15 15 9 1 10 15 9 7 9 1 9 1 9 13 2 13 3 10 0 9 1 15 9 2
18 1 11 13 3 15 9 7 9 1 3 12 9 1 10 9 1 9 2
9 15 8 4 1 15 10 9 4 2
20 15 13 15 13 1 10 9 2 16 15 9 1 10 0 2 0 9 2 13 2
19 1 12 9 13 10 9 2 8 10 9 13 1 9 2 15 13 8 4 2
17 3 4 10 9 2 3 11 2 1 0 9 4 7 4 1 0 2
31 3 13 8 10 11 10 9 1 10 9 7 10 9 1 7 10 11 7 1 15 8 4 4 4 2 15 15 8 13 4 2
11 3 13 3 9 2 16 1 10 9 8 2
33 10 9 1 10 0 9 11 13 8 4 2 16 3 10 15 9 4 16 1 10 9 1 11 7 11 2 15 3 0 8 4 4 2
32 8 2 0 9 1 8 2 13 11 1 11 10 9 1 11 5 9 1 11 1 10 9 1 15 8 1 9 5 7 8 4 2
7 11 13 11 1 11 3 2
26 10 0 9 1 11 7 11 2 12 1 10 0 9 2 13 4 4 1 10 3 3 1 13 0 9 2
14 10 0 9 2 12 2 13 8 4 1 10 9 11 2
4 13 15 4 2
10 15 4 4 1 15 9 11 7 11 2
35 1 12 9 9 1 10 0 9 1 9 1 10 11 2 13 15 8 11 7 11 10 9 1 10 9 4 2 15 3 1 15 9 4 4 2
25 8 7 8 13 1 10 9 1 4 4 1 10 9 7 9 7 10 9 15 1 15 9 4 4 2
31 10 9 13 1 12 9 4 4 1 12 9 2 1 15 10 9 1 9 1 10 9 0 1 12 9 4 4 1 10 9 2
36 15 13 3 3 3 4 2 16 15 8 1 11 3 3 10 9 4 4 1 10 9 16 0 9 1 10 9 8 7 1 10 9 11 1 4 2
22 9 4 8 2 16 11 1 10 9 1 12 9 10 9 1 8 1 9 4 4 4 2
22 1 11 13 15 15 9 0 4 4 1 8 1 9 2 3 1 10 9 1 12 9 2
14 1 10 9 4 3 10 13 12 9 13 0 8 4 2
14 10 9 1 15 9 13 1 12 1 12 1 3 12 2
14 3 13 1 15 9 3 0 9 2 3 1 10 9 2
23 15 9 8 10 0 9 1 15 9 2 15 1 10 9 11 4 4 2 13 3 0 9 2
7 3 13 15 3 3 4 2
15 1 10 3 0 9 13 3 15 9 2 3 10 0 9 2
12 10 0 12 9 4 0 1 15 0 1 12 2
14 3 1 10 0 9 13 0 9 2 3 1 0 9 2
18 1 15 8 4 3 0 9 4 1 10 9 1 10 0 9 1 11 2
35 3 9 11 2 11 2 2 8 2 11 2 7 11 2 11 2 13 10 0 9 1 10 9 3 2 3 15 9 10 9 2 9 2 13 2
21 9 11 13 3 3 16 15 3 10 9 4 16 3 0 4 4 1 10 0 9 2
22 15 13 3 9 4 1 10 9 1 9 7 10 9 1 11 7 15 13 15 9 4 2
32 15 13 10 9 1 8 7 10 9 2 15 1 11 0 2 2 2 0 9 1 12 3 15 10 9 3 13 2 0 0 4 2
21 1 8 13 10 9 3 1 4 4 11 0 5 15 13 1 10 9 1 10 9 2
21 8 2 16 15 9 11 2 0 0 13 2 13 10 15 9 1 10 9 16 11 2
7 15 13 1 10 9 2 2
9 15 13 3 3 1 15 3 4 2
16 1 15 9 13 10 0 9 8 15 1 4 16 15 3 4 2
14 15 9 4 15 1 10 0 9 8 1 10 9 4 2
8 10 9 13 3 1 15 9 2
16 1 10 9 1 10 0 9 13 10 9 3 10 16 12 9 2
17 10 9 13 16 10 9 1 0 9 1 9 1 15 9 4 4 2
29 1 10 0 9 1 10 9 2 8 2 1 8 1 10 15 9 13 10 11 15 1 10 0 9 4 1 10 9 2
33 10 0 9 4 15 10 0 9 1 2 8 2 1 9 1 13 9 1 10 9 0 0 9 2 15 9 4 10 9 2 8 2 2
17 7 3 13 10 11 0 15 16 2 9 2 7 2 9 4 2 2
5 2 15 13 2 2
2 11 2
16 15 13 0 9 1 10 9 1 10 0 9 1 10 0 9 2
8 1 8 1 8 4 4 3 2
3 10 0 2
11 15 13 8 9 15 10 0 9 13 4 2
35 7 10 9 1 15 9 2 8 2 16 10 9 1 10 9 2 8 1 11 2 13 16 10 9 1 10 9 0 15 3 0 13 4 4 2
10 2 11 7 11 13 0 15 1 9 2
17 10 9 1 11 13 1 15 1 0 9 4 1 10 9 1 11 2
16 16 10 9 1 10 9 1 10 9 1 4 13 15 13 0 2
31 11 7 11 13 3 0 9 3 2 0 11 2 11 7 11 2 7 15 13 3 3 1 4 1 3 15 1 9 4 4 2
11 1 11 4 10 0 9 2 8 2 4 2
11 2 15 13 12 9 16 10 9 1 4 2
15 9 8 13 1 10 0 9 2 3 1 9 11 1 11 2
15 15 13 1 0 9 2 7 10 9 1 15 0 9 13 2
12 15 0 9 1 9 7 9 1 10 0 9 2
44 3 13 15 10 13 9 2 7 10 9 13 2 3 1 9 1 10 0 0 9 1 9 0 13 8 1 10 0 11 2 1 10 9 9 2 3 8 9 15 3 4 13 4 2
40 10 9 11 13 10 9 3 2 10 9 15 10 9 1 10 0 9 1 10 9 1 9 7 9 13 4 2 3 1 4 4 1 9 16 10 9 15 9 13 2
31 2 16 10 9 1 10 15 9 13 2 3 13 9 7 9 15 1 0 9 1 10 9 3 4 4 2 2 3 13 15 2
30 0 1 9 2 1 0 9 2 9 1 9 2 0 1 9 2 13 16 9 1 8 7 11 7 3 10 9 1 9 2
32 15 9 4 0 2 1 10 9 1 10 9 8 1 9 2 9 7 9 2 1 11 2 8 1 11 7 10 9 11 1 11 2
11 2 8 2 13 11 1 9 1 10 11 2
12 15 2 9 1 9 2 4 3 3 0 9 2
8 1 0 13 15 15 8 4 2
14 1 11 13 15 9 15 1 10 9 1 15 9 4 2
31 8 4 10 9 3 1 10 0 9 4 2 7 15 13 3 10 0 9 2 16 10 0 9 3 3 0 9 1 15 13 2
19 10 0 0 0 9 2 1 0 9 13 3 3 10 13 9 1 9 4 2
32 10 9 13 10 9 4 2 7 10 9 13 15 3 0 4 16 10 9 1 13 1 10 0 13 13 9 1 10 9 1 9 2
20 15 9 13 15 2 1 0 9 2 4 7 3 13 15 12 9 3 4 2 2
23 10 9 8 1 10 11 1 10 11 13 2 3 15 9 2 1 4 2 7 15 15 2 2
34 9 11 13 10 11 4 10 9 3 3 0 1 4 4 2 16 10 11 1 15 9 1 15 9 1 2 10 0 0 9 2 13 4 2
11 15 13 10 9 1 10 9 0 3 4 2
30 15 13 9 1 10 9 15 13 1 10 2 13 9 2 2 15 13 1 10 9 7 10 9 1 10 9 15 13 4 2
19 7 3 9 7 9 1 10 9 7 12 9 3 0 13 2 4 15 0 2
12 7 1 0 13 15 3 15 9 15 4 2 2
27 15 13 10 0 9 0 0 13 1 10 0 9 2 2 8 2 2 16 1 10 9 13 9 1 2 8 2
12 3 13 15 0 1 10 0 9 3 9 2 2
20 10 0 9 1 11 13 16 15 3 1 15 9 2 15 0 4 2 4 4 2
15 15 13 15 3 0 7 13 15 9 4 10 9 1 4 2
19 2 7 2 16 10 0 9 1 12 9 4 4 2 3 13 15 3 3 2
14 10 9 4 3 0 2 15 13 0 3 15 15 4 2
9 15 13 3 3 0 0 4 2 2
20 1 11 13 10 9 1 10 9 1 9 4 16 10 9 1 10 9 1 4 2
10 15 9 4 3 3 9 1 15 8 2
3 9 8 2
12 15 13 3 3 15 9 1 15 9 3 4 2
9 10 11 13 3 10 9 4 4 2
13 3 13 15 10 9 3 16 10 9 1 4 4 2
16 7 10 9 13 4 4 2 16 10 9 3 0 4 1 9 2
10 9 9 1 10 0 9 11 8 11 2
38 10 1 15 9 13 9 1 12 9 2 1 10 9 13 1 10 9 1 12 9 2 13 3 1 10 0 9 1 10 3 3 0 9 1 10 0 9 2
28 16 10 9 4 4 7 10 9 4 13 15 12 13 1 10 9 1 10 9 7 10 0 9 1 10 13 9 2
52 10 9 1 10 9 2 9 8 2 0 9 1 10 0 0 9 1 11 2 13 3 1 0 9 10 9 4 7 1 11 13 10 9 1 9 2 16 0 3 1 13 3 15 9 10 9 1 10 9 4 4 2
36 3 13 3 0 9 4 1 8 2 12 2 2 15 1 10 0 9 1 15 8 2 10 3 0 9 7 0 9 1 10 11 8 7 9 8 2
21 10 9 13 1 10 9 1 0 9 1 11 7 13 1 10 9 1 12 9 4 2
29 2 15 13 15 3 1 15 13 7 13 3 3 15 9 1 15 9 1 15 9 7 16 15 15 3 3 13 4 2
3 15 13 2
23 2 16 15 13 10 9 3 1 4 2 3 10 9 1 10 13 9 2 3 13 15 3 2
9 7 3 16 15 1 10 9 4 2
16 15 13 10 9 4 1 11 15 1 15 1 15 9 13 2 2
5 8 13 3 0 2
10 2 1 0 9 13 15 3 15 4 2
9 9 13 3 1 15 9 0 4 2
11 9 7 9 1 10 9 4 3 1 4 2
19 11 13 15 9 1 10 9 8 1 11 4 1 10 0 9 11 1 11 2
35 10 9 2 15 15 9 13 1 10 0 9 1 10 9 11 2 13 1 10 9 1 3 12 9 0 0 12 12 9 9 1 3 0 9 2
14 15 13 0 2 6 2 2 16 15 0 3 0 4 2
24 10 11 4 0 10 9 1 10 9 3 1 4 16 1 10 9 1 9 7 9 15 9 13 2
17 10 0 9 1 10 9 4 3 2 16 10 9 1 10 0 13 2
9 3 15 0 3 4 10 0 9 2
23 10 0 13 7 9 13 0 4 4 2 16 15 1 0 9 15 3 3 3 4 4 4 2
14 15 2 15 3 4 4 4 2 13 15 1 9 4 2
25 10 0 9 13 2 16 10 9 4 4 7 13 0 15 2 9 2 16 15 3 4 4 2 4 2
17 2 15 13 10 9 4 1 10 0 9 7 1 10 0 0 9 2
11 15 4 4 1 10 9 7 3 9 3 2
26 7 15 4 3 2 16 15 3 13 16 16 11 3 0 4 2 15 1 15 9 3 0 0 3 4 2
32 7 15 13 1 15 4 2 1 15 9 7 9 2 7 1 15 15 9 2 16 11 15 4 2 16 15 15 13 4 7 4 2
15 15 13 15 10 9 4 16 15 10 9 13 6 7 6 2
28 0 9 1 11 13 1 0 9 4 1 4 1 0 9 1 10 9 1 0 9 7 10 3 0 13 9 8 2
24 1 10 0 9 9 15 9 13 10 9 9 4 7 4 2 9 4 7 4 7 4 1 9 2
28 8 13 3 3 2 16 10 9 5 1 10 9 4 3 10 16 12 0 9 4 5 0 9 0 9 4 4 2
28 10 0 9 13 1 10 9 10 9 1 15 9 1 10 9 2 3 15 3 13 4 2 3 13 10 9 0 2
18 10 9 2 15 10 9 13 1 4 2 13 0 1 10 9 4 4 2
13 10 9 4 10 0 1 11 3 10 9 13 4 2
24 1 11 0 9 4 12 0 9 5 1 15 12 9 5 1 0 9 4 7 4 8 0 13 2
31 15 13 9 13 9 4 1 13 9 2 15 13 9 9 2 1 10 9 3 0 9 13 15 16 1 0 9 3 4 4 2
24 3 13 15 9 2 3 0 9 10 9 13 2 7 3 1 10 9 13 15 0 7 13 3 2
25 10 13 0 9 2 0 9 15 1 10 9 4 4 2 9 2 15 3 3 0 4 16 10 9 2
15 1 10 0 0 9 9 10 0 9 1 9 1 15 9 2
9 15 15 13 13 15 15 10 9 2
35 10 13 9 1 9 4 10 10 9 0 4 2 3 12 9 1 0 12 9 15 4 13 1 10 9 1 15 8 1 10 0 9 1 11 2
22 1 9 1 10 9 1 0 9 13 15 9 12 9 7 15 9 4 1 10 0 9 2
29 1 10 9 1 10 0 9 5 15 9 13 3 0 4 4 5 4 12 9 1 10 0 9 0 1 10 0 9 2
7 15 9 1 3 0 9 2
21 1 11 4 11 10 9 4 1 15 13 1 0 9 2 15 4 4 1 15 13 2
18 10 9 10 0 11 1 10 9 11 1 11 2 13 9 1 10 9 2
16 10 9 13 16 10 9 1 10 9 1 10 9 11 9 13 2
21 10 9 13 9 1 4 1 10 9 0 9 1 15 13 2 15 1 10 9 13 2
33 10 0 9 7 9 13 4 16 15 4 1 10 9 1 15 11 8 1 15 9 13 4 4 1 10 9 1 10 11 1 13 9 2
18 10 11 13 13 9 1 11 3 16 1 13 1 10 9 1 10 9 2
9 15 4 3 0 1 15 9 3 2
17 10 0 9 7 9 7 10 11 4 0 9 1 9 1 10 9 2
13 10 9 1 11 13 10 9 8 12 9 4 4 2
18 10 9 1 10 9 7 10 9 13 15 1 15 0 0 9 1 9 2
7 3 13 3 0 9 0 2
19 1 10 9 3 4 10 0 0 9 1 10 0 9 0 16 3 0 4 2
29 15 13 1 9 2 15 1 10 9 3 0 4 2 13 1 10 0 9 3 9 1 0 9 1 10 0 9 4 2
48 1 10 13 9 13 10 9 1 9 8 1 10 9 1 15 8 1 10 0 9 1 10 16 12 9 10 0 9 4 7 3 1 10 9 1 10 9 15 9 4 7 10 9 2 8 2 4 2
30 1 10 9 13 10 9 10 9 1 12 9 2 3 3 10 0 2 9 2 9 7 0 2 7 1 10 0 8 3 2
28 2 15 13 15 9 1 10 9 4 2 2 3 13 10 9 2 2 7 15 4 10 0 9 15 15 0 13 2
24 4 4 3 10 9 1 4 1 15 0 8 2 15 3 13 4 1 10 0 9 1 10 9 2
26 8 10 0 9 15 10 9 1 15 9 13 2 13 10 9 1 10 9 2 15 0 2 11 2 4 2
14 15 8 13 2 8 10 9 2 10 9 4 2 0 2
4 9 1 9 2
10 15 9 13 13 1 10 9 0 9 2
20 10 9 13 3 1 10 0 9 1 9 15 10 0 9 1 11 0 9 9 2
11 8 12 13 10 9 10 9 1 12 9 2
38 1 12 7 1 12 13 10 0 9 1 10 9 9 4 2 0 1 10 9 1 10 9 1 9 2 7 3 13 1 9 3 3 16 9 9 0 4 2
23 3 4 10 9 1 9 1 12 9 4 1 3 8 2 16 10 9 9 1 12 4 4 2
24 1 10 0 9 1 9 13 3 10 9 7 1 0 1 10 9 10 9 3 3 1 10 9 2
7 9 13 3 10 9 9 2
15 9 7 9 2 15 3 0 4 4 2 13 3 0 3 2
18 12 1 9 13 9 1 12 9 9 13 7 12 9 0 9 9 13 2
22 1 10 9 1 9 13 1 11 7 9 10 9 9 3 2 15 1 10 9 4 4 2
21 15 13 0 10 0 9 1 1 10 9 13 9 2 15 0 1 10 9 4 4 2
13 9 2 15 1 10 9 13 4 4 2 4 8 2
43 2 0 0 9 2 2 2 9 2 9 2 9 7 9 2 2 2 10 9 2 2 2 9 2 2 2 9 2 2 2 0 9 2 2 7 2 10 9 1 10 9 2 2
40 10 9 2 10 9 2 2 7 2 10 9 2 13 8 4 1 9 2 15 15 9 1 10 9 1 15 8 7 1 10 9 1 10 9 1 12 13 4 4 2
12 10 0 9 1 15 8 4 0 16 10 9 2
7 15 9 4 0 1 4 2
19 1 9 1 10 9 10 9 1 11 13 10 9 1 11 15 0 8 4 2
30 10 9 13 0 16 15 3 1 10 0 9 1 10 0 11 13 9 1 10 11 1 11 1 11 10 13 9 4 4 2
23 10 9 1 0 9 2 9 7 15 9 15 1 10 9 4 4 2 4 1 11 3 4 2
20 12 9 9 2 12 9 2 1 10 12 9 13 1 9 1 15 9 7 9 2
8 10 9 1 12 9 13 8 2
6 8 4 15 0 8 2
17 10 9 13 3 10 9 2 3 15 11 1 11 1 10 9 13 2
13 8 3 2 10 9 2 4 1 3 1 8 4 2
21 3 13 11 9 1 10 9 1 10 0 9 11 7 11 2 15 9 15 9 13 2
17 11 13 0 3 1 10 9 11 2 10 3 0 1 10 0 9 2
29 8 2 10 0 9 15 10 9 1 15 9 13 2 4 1 10 9 1 15 9 4 3 15 1 9 3 4 4 2
20 15 4 3 10 3 0 9 4 2 15 10 0 9 1 10 9 3 0 13 2
42 3 13 15 1 12 1 15 0 15 9 0 9 1 9 7 13 1 15 15 13 9 1 0 9 2 9 7 9 1 9 2 9 7 9 9 16 10 0 9 1 11 2
28 15 8 2 15 15 0 13 1 9 1 10 9 7 1 10 9 1 10 9 7 10 9 2 4 13 1 11 2
13 1 15 13 10 9 1 9 2 0 13 2 13 2
30 10 9 15 13 16 1 10 11 1 11 1 4 4 1 15 4 7 3 13 10 9 1 13 0 1 11 1 4 4 2
22 1 10 9 4 1 15 8 4 16 10 0 9 1 10 9 1 10 13 9 4 4 2
15 3 13 15 10 9 1 10 9 1 10 9 7 10 11 2
8 10 9 8 13 3 15 13 2
39 15 4 3 10 9 1 10 9 16 1 10 9 10 9 1 4 1 10 0 9 7 11 7 10 9 16 1 11 7 11 10 9 1 4 13 3 1 15 2
17 12 9 3 13 15 1 10 0 9 10 9 3 1 10 9 11 2
32 15 4 3 0 2 13 10 9 11 2 9 2 7 11 2 9 2 16 0 9 10 9 1 15 13 1 8 8 13 4 4 2
15 3 13 10 9 10 9 8 1 8 2 9 1 15 8 2
8 10 9 11 13 3 9 3 2
31 1 10 0 9 13 8 10 0 9 1 10 9 7 10 9 1 9 1 8 4 2 13 10 9 1 15 9 1 10 9 2
8 0 0 1 10 0 0 9 2
18 1 2 11 2 4 3 10 0 0 9 4 1 10 9 1 10 9 2
16 3 0 7 1 15 0 9 2 16 15 3 10 0 9 13 2
26 4 4 3 10 9 1 10 0 9 1 10 0 9 8 2 15 0 13 1 10 1 15 9 13 11 2
12 7 3 10 9 1 11 7 11 1 10 9 2
10 12 2 4 10 0 9 1 11 2 2
23 10 9 1 10 9 0 13 1 15 0 0 13 3 8 1 10 9 1 10 9 1 11 2
17 15 9 1 9 2 9 2 9 7 11 4 3 1 0 9 4 2
44 16 10 0 13 9 4 10 9 7 9 0 10 9 1 4 7 1 0 15 0 9 13 0 9 1 15 9 1 10 0 9 4 4 4 2 1 10 3 0 9 1 11 9 2
20 15 13 10 9 16 10 0 9 1 10 9 4 1 10 15 9 1 10 9 2
25 10 13 9 9 7 0 9 4 15 0 16 10 9 9 2 7 1 10 0 9 0 1 15 8 2
25 10 12 0 9 15 11 9 11 5 10 3 0 9 1 8 1 15 8 5 8 13 2 4 0 2
19 1 15 9 4 1 8 10 9 1 10 9 1 10 9 0 9 0 4 2
23 10 9 13 3 1 10 9 3 3 2 3 1 0 9 15 9 1 4 2 3 13 15 2
50 10 11 13 3 4 10 0 9 8 2 11 2 2 16 9 1 15 0 13 7 16 9 1 15 7 15 0 9 2 2 1 10 0 9 8 2 8 2 8 7 8 16 0 9 1 11 3 1 4 2
13 10 9 2 15 1 2 9 2 8 0 4 4 2
12 2 3 4 3 4 16 3 12 9 4 4 2
7 3 13 3 3 3 12 2
11 7 3 4 3 3 3 10 9 4 2 2
25 10 9 13 1 8 2 8 2 8 2 8 2 8 7 8 13 1 10 13 9 12 0 9 4 2
21 15 13 1 10 9 1 9 12 8 4 4 15 9 3 1 4 7 1 4 4 2
18 10 9 13 3 8 10 9 2 1 9 1 10 1 15 2 9 2 2
16 8 13 10 9 3 10 9 4 2 3 10 9 1 9 13 2
20 9 1 10 9 1 10 9 2 15 4 4 1 15 8 2 13 9 1 8 2
57 3 13 10 9 1 9 4 3 9 11 2 0 9 2 7 9 11 2 9 2 1 15 9 1 10 9 1 0 9 1 15 9 0 4 1 4 1 10 0 13 9 2 16 10 0 9 4 4 1 4 1 11 7 1 10 11 2
15 1 10 3 13 9 13 10 11 1 12 9 4 4 4 2
21 10 9 1 11 13 0 12 9 0 4 2 1 0 3 10 0 9 1 12 9 2
12 0 16 10 9 1 11 13 11 15 3 4 2
13 2 15 13 3 15 3 2 7 15 13 3 0 2
15 15 13 15 4 1 15 0 9 16 8 7 8 3 2 2
12 1 8 13 11 12 9 3 8 1 10 11 2
9 1 15 9 13 15 10 0 9 2
23 15 13 3 1 9 8 13 4 1 9 12 7 15 15 9 4 10 9 10 13 9 4 2
4 15 13 0 2
16 2 15 4 10 0 9 3 3 15 15 9 4 4 1 9 2
15 3 15 0 4 3 16 8 13 1 15 1 11 4 4 2
20 2 15 13 1 10 9 9 1 15 9 0 0 7 0 0 2 2 13 15 2
21 15 13 3 3 3 7 3 1 10 9 1 10 9 13 15 3 1 15 0 9 2
24 10 9 13 15 1 15 9 1 10 11 3 4 2 4 1 10 0 9 1 10 13 9 4 2
31 10 11 12 15 9 0 16 9 1 4 1 15 0 9 8 2 15 10 9 8 1 10 9 1 12 2 0 2 13 4 2
34 8 2 0 9 1 10 11 2 13 15 1 10 9 1 10 9 8 8 10 9 1 15 9 3 1 10 9 1 10 9 11 4 4 2
22 2 10 9 11 4 15 0 9 1 0 9 9 2 2 3 10 9 11 1 15 9 2
26 10 9 1 10 0 9 1 10 13 9 13 10 9 1 15 3 4 4 1 3 12 1 12 12 9 2
27 15 13 10 0 7 0 9 1 4 2 7 3 10 16 12 9 13 4 1 10 9 1 10 9 1 11 2
11 15 4 3 4 7 1 10 9 4 4 2
29 10 0 9 1 9 7 9 13 1 10 0 9 1 10 9 7 10 9 1 10 9 15 9 1 10 0 9 4 2
11 10 9 1 0 9 13 4 1 13 9 2
26 10 0 0 0 9 2 15 1 10 11 1 10 11 1 11 2 4 1 10 0 0 9 1 11 4 2
26 3 10 9 1 10 0 9 4 3 1 9 1 10 0 0 9 2 3 3 3 10 16 12 9 13 2
44 3 13 1 10 0 9 1 10 9 4 4 16 10 9 8 0 4 4 4 7 3 10 0 9 1 11 2 3 3 1 0 9 1 15 9 1 10 9 2 1 10 9 4 2
25 10 9 13 1 10 0 9 10 0 9 4 2 15 13 1 10 9 1 0 9 1 0 12 9 2
16 2 10 13 7 3 8 13 9 1 10 9 1 10 9 2 2
32 15 13 10 9 8 2 12 2 2 9 1 10 0 1 10 9 13 9 8 2 1 10 9 1 9 8 16 1 9 1 4 2
14 2 1 15 9 13 15 15 1 15 15 1 15 9 2
9 3 13 15 1 10 9 1 15 2
21 1 10 0 9 2 15 15 3 1 8 13 4 2 13 15 9 1 15 13 9 2
30 10 9 13 1 10 9 15 11 1 12 9 1 12 1 12 9 0 9 13 7 12 9 1 10 9 1 10 9 13 2
16 10 9 4 8 9 4 1 10 0 9 1 10 9 1 11 2
24 10 15 9 4 1 9 4 7 13 10 9 4 2 15 15 1 15 9 3 1 10 9 13 2
6 15 13 15 13 3 2
11 15 13 15 3 3 15 10 9 2 6 2
10 7 9 13 15 3 8 9 1 15 2
8 1 15 3 13 15 9 3 2
29 15 9 2 2 11 13 12 9 7 12 9 1 10 12 7 12 9 2 2 13 3 1 10 9 7 10 9 9 2
16 15 13 15 3 0 3 4 2 7 3 13 15 15 15 4 2
9 7 16 15 13 4 15 3 3 2
13 2 11 7 3 10 9 0 9 13 10 9 3 2
17 10 11 13 10 0 7 0 9 1 10 9 0 4 1 10 0 2
9 1 12 7 12 9 10 0 9 2
23 15 13 10 0 9 3 2 16 2 3 9 8 2 2 15 3 3 1 15 9 4 2 2
3 15 13 2
24 2 15 4 15 0 15 3 1 13 16 15 1 10 9 3 4 4 3 8 10 9 0 4 2
4 1 15 9 2
18 16 10 0 9 1 15 9 10 9 13 2 13 10 11 0 15 9 2
32 10 0 9 13 3 1 10 9 9 3 4 2 16 15 1 10 9 1 11 7 11 10 9 1 10 9 1 15 9 4 4 2
23 15 13 1 10 9 1 12 2 13 8 2 12 1 12 9 0 2 3 15 9 13 4 2
14 10 9 13 10 9 1 8 1 10 9 1 8 4 2
14 15 13 1 10 9 1 10 0 9 2 2 13 15 2
27 15 13 15 1 11 1 10 9 4 4 7 13 15 3 2 13 1 10 9 2 1 10 9 1 15 9 2
26 3 13 3 3 11 7 11 10 9 2 7 3 11 7 11 13 3 12 1 12 12 9 3 10 9 2
24 3 13 3 10 9 1 12 9 1 9 3 3 15 8 4 2 15 15 3 0 3 15 13 2
8 11 13 3 13 1 11 3 2
11 1 10 16 12 9 13 15 15 9 4 2
13 3 13 8 1 10 9 1 8 10 0 9 4 2
25 1 15 13 10 9 3 3 0 9 1 15 7 13 1 10 9 3 15 2 0 9 2 4 4 2
23 9 8 13 3 1 10 9 3 16 15 3 1 15 8 4 4 15 1 15 13 1 13 2
14 15 13 3 4 1 1 10 13 0 9 1 10 9 2
18 8 13 0 4 16 3 0 4 4 4 1 10 0 9 1 10 9 2
9 2 15 13 10 9 7 10 9 2
38 11 9 4 3 3 3 16 1 15 1 0 9 13 9 1 11 2 15 1 15 9 16 10 0 11 10 9 1 15 11 3 13 2 10 9 1 4 2
53 11 2 10 0 9 2 10 0 2 15 3 13 16 10 0 9 1 10 0 12 9 1 11 9 2 13 8 15 3 1 9 15 9 4 3 10 9 4 2 7 13 1 0 2 0 9 15 9 1 10 9 3 2
8 0 9 2 9 13 15 3 2
13 13 1 10 9 8 4 13 1 10 9 1 11 2
13 10 9 2 8 10 9 2 7 10 0 0 9 2
10 3 13 1 10 9 2 8 10 9 2
12 2 3 4 4 1 10 9 2 2 13 15 2
24 2 3 13 16 10 9 3 15 0 4 4 2 16 15 3 1 10 0 9 13 4 7 4 2
10 10 9 4 9 2 9 2 9 2 2
12 1 11 13 15 9 0 9 4 1 0 9 2
10 1 12 4 15 3 0 4 16 9 2
12 9 1 15 0 9 2 0 1 9 7 9 2
9 8 13 3 10 9 3 4 4 2
10 7 15 13 15 0 9 3 0 4 2
13 15 4 2 16 15 15 13 2 3 1 10 9 2
12 2 15 13 15 9 3 1 15 9 7 9 2
16 15 13 15 3 1 15 1 13 4 7 15 13 3 3 9 2
9 8 4 0 1 15 15 4 13 2
23 15 13 4 16 15 3 1 10 9 3 15 4 4 15 15 1 10 9 3 3 13 4 2
23 15 9 13 3 1 0 9 10 0 9 1 15 9 1 10 9 16 15 16 9 0 13 2
6 10 9 1 10 9 2
16 15 13 10 0 9 4 4 16 10 9 3 8 1 13 4 2
21 7 3 4 10 9 3 3 4 2 8 2 2 3 1 10 0 0 9 1 8 2
25 0 7 13 9 13 1 10 9 0 4 4 2 13 15 15 10 9 8 13 2 16 15 9 4 2
30 1 9 13 11 15 12 1 15 2 9 2 2 7 0 13 3 11 2 11 2 11 2 11 2 11 7 11 9 4 2
12 8 4 10 9 1 3 10 9 9 7 12 2
17 10 3 0 9 15 11 1 15 13 9 13 4 2 4 10 9 2
19 10 9 9 3 13 10 0 9 16 9 1 10 0 9 1 11 7 11 2
21 15 13 10 9 1 13 1 13 16 15 10 9 4 7 9 0 1 10 9 13 2
19 7 1 10 0 9 16 3 3 1 9 9 4 16 10 9 3 1 13 2
15 15 9 13 8 4 16 15 3 3 1 15 9 0 4 2
9 12 9 3 15 15 13 0 4 2
7 10 9 4 3 3 15 2
16 10 9 4 3 3 3 1 16 15 9 3 0 0 1 4 2
7 10 9 1 10 9 4 2
3 0 9 2
6 9 7 10 9 9 2
3 0 9 2
4 12 9 9 2
3 0 9 2
4 10 9 9 2
3 0 9 2
8 0 9 7 9 1 10 9 2
14 15 16 9 13 3 1 0 9 10 9 3 1 4 2
4 1 10 9 2
3 0 9 2
3 1 9 2
12 12 0 9 9 2 10 9 9 0 7 9 2
3 1 9 2
30 12 9 9 2 10 9 9 0 2 9 1 10 0 9 1 10 9 1 10 0 9 7 12 9 9 1 10 0 9 2
11 11 9 8 1 10 9 9 1 10 9 2
19 15 9 4 4 1 10 9 1 10 9 1 10 9 8 2 9 1 11 2
11 10 9 11 13 0 4 1 9 7 9 2
19 15 4 3 1 10 9 4 16 13 1 10 9 2 8 13 2 0 4 2
19 15 13 3 3 3 15 9 0 4 2 1 15 9 13 10 9 3 4 2
9 3 13 15 15 15 9 3 3 2
22 15 9 1 10 9 16 9 1 10 9 11 1 0 2 1 15 13 9 0 2 9 2
22 15 4 3 13 4 2 3 16 1 10 0 9 3 4 4 3 15 0 1 4 4 2
26 10 9 2 13 1 10 9 8 2 9 11 2 9 11 7 8 2 4 1 10 9 4 16 10 9 2
26 1 3 1 10 9 1 10 9 2 1 12 2 4 3 9 1 15 0 13 1 10 3 3 0 9 2
11 7 3 4 3 3 8 10 9 1 4 2
11 3 4 12 9 1 10 9 1 8 4 2
20 10 9 11 7 10 9 11 13 3 4 16 12 1 10 12 9 0 1 4 2
29 10 9 1 11 2 11 2 11 2 11 7 11 13 10 9 2 16 10 9 13 2 3 1 10 9 1 12 9 2
26 0 13 10 12 9 15 15 1 10 13 9 4 7 15 16 9 1 10 9 10 9 4 1 10 9 2
41 10 9 1 15 9 2 15 1 10 3 12 9 0 9 12 9 13 4 2 4 11 2 11 2 8 7 11 2 15 0 9 8 4 4 1 9 1 8 12 9 2
39 3 13 4 12 9 1 10 9 2 10 0 9 8 2 12 2 7 8 2 12 2 2 0 1 10 9 11 2 8 1 10 9 3 10 0 0 9 13 2
23 10 9 1 10 9 2 11 1 11 2 13 1 10 11 1 10 9 11 7 13 15 9 2
20 15 13 1 10 11 8 1 10 9 13 1 10 9 11 13 1 11 1 11 2
24 15 4 10 3 0 0 9 2 3 11 0 9 13 7 1 10 11 1 11 4 4 1 9 2
7 15 13 3 10 9 3 2
19 10 0 9 13 3 10 13 9 2 15 3 10 9 1 10 9 13 4 2
8 10 0 9 4 3 9 4 2
39 1 12 9 1 7 12 9 2 10 9 11 7 8 2 13 10 9 10 9 1 10 9 1 11 2 10 9 1 8 7 15 1 10 9 1 9 1 4 2
26 3 13 10 9 0 1 10 9 16 1 15 9 2 13 1 10 11 7 10 11 2 10 9 1 4 2
11 8 4 10 9 15 1 10 11 4 4 2
13 0 1 9 2 7 1 15 9 1 9 1 8 2
8 15 13 10 9 1 9 4 2
23 1 12 4 15 8 1 8 2 16 9 1 15 8 1 11 7 1 10 11 2 0 9 2
17 15 13 10 0 9 1 8 8 1 11 7 13 1 11 7 11 2
10 16 9 13 11 11 1 12 0 4 2
20 3 13 12 9 1 12 9 1 11 2 3 3 12 3 3 1 9 4 4 2
24 9 11 13 1 0 9 7 1 9 9 1 10 9 7 1 10 9 1 0 9 10 9 4 2
19 10 9 13 3 4 0 0 1 4 1 15 13 1 0 9 1 0 9 2
20 10 9 4 0 4 7 13 15 9 7 1 9 7 1 0 9 1 9 4 2
10 15 8 13 9 1 10 9 1 11 2
11 3 13 10 9 1 8 2 8 2 4 2
17 2 10 0 9 1 11 4 15 0 8 4 2 2 3 13 15 2
7 10 9 13 0 15 9 2
35 3 13 10 9 1 3 9 2 3 11 10 9 1 10 9 1 11 15 3 10 10 9 1 10 9 13 2 13 2 1 3 10 9 3 2
10 15 8 13 13 9 1 8 4 4 2
17 16 1 12 4 10 9 4 1 10 9 15 1 11 1 11 13 2
26 1 10 9 16 10 9 4 1 15 8 7 10 11 1 11 13 10 9 3 10 0 9 1 10 9 2
13 15 8 13 4 1 15 0 2 8 2 1 9 2
21 2 8 2 2 10 9 1 10 2 0 9 1 10 9 11 13 1 12 9 3 2
27 10 0 13 1 10 9 9 1 0 9 2 11 2 11 2 8 7 8 2 15 3 1 11 15 0 4 2
29 3 3 10 9 1 9 8 1 10 9 11 7 10 9 1 15 0 0 2 8 2 2 15 10 9 1 11 13 2
12 10 9 1 10 9 4 3 13 1 10 0 2
36 15 9 13 15 4 16 10 13 9 1 10 9 1 10 9 1 15 8 0 1 15 9 2 3 16 15 9 1 11 3 0 13 4 13 4 2
21 2 15 4 11 2 6 2 2 13 15 1 0 0 2 2 9 11 2 6 2 2
26 1 11 4 15 15 3 3 0 2 16 10 9 15 3 0 4 4 1 9 1 9 2 9 7 9 2
26 10 9 1 10 0 9 13 3 10 9 1 9 1 8 4 4 7 1 15 9 13 15 0 9 4 2
17 15 0 9 4 16 15 10 9 1 15 9 1 8 13 4 4 2
25 15 9 13 9 1 15 9 1 9 1 10 9 1 10 9 16 11 7 11 15 1 10 9 4 2
14 11 13 15 10 9 1 9 1 10 9 1 4 4 2
21 3 13 15 1 4 4 15 9 1 10 9 0 2 8 1 12 2 3 1 4 2
28 9 4 3 1 10 0 9 4 7 10 3 13 9 2 10 9 1 3 0 9 9 2 4 1 10 9 4 2
30 9 12 13 10 9 1 12 9 1 10 9 2 9 12 1 12 9 2 9 12 1 12 9 7 9 12 1 10 9 2
31 10 9 13 16 1 10 0 13 9 2 15 0 1 10 9 12 7 12 13 2 10 9 0 4 4 16 0 9 1 13 2
13 15 4 1 10 9 10 9 1 10 9 1 11 2
12 15 4 15 3 2 10 11 1 10 0 9 2
36 11 9 2 9 7 9 8 7 10 15 2 8 2 9 2 2 8 2 9 2 7 8 2 9 2 2 13 0 4 15 3 1 15 4 4 2
41 13 16 10 9 13 15 3 10 9 3 2 15 3 13 1 9 1 10 13 9 8 2 8 2 8 7 8 2 7 0 15 9 1 15 9 7 9 1 15 9 2
20 10 2 9 2 1 15 15 4 3 0 0 7 4 0 3 3 1 15 9 2
21 1 10 0 9 13 10 0 9 11 1 10 9 1 1 15 12 7 12 12 9 2
25 0 7 0 1 10 9 4 10 9 11 7 8 2 15 12 9 13 1 1 15 12 7 12 12 2
18 10 0 9 1 10 0 9 8 2 11 2 13 15 3 0 9 4 2
15 15 9 4 1 12 4 1 10 9 1 12 1 12 12 2
21 1 10 9 3 1 10 9 1 15 0 8 4 10 0 9 11 1 9 8 4 2
20 1 10 9 1 10 0 9 11 2 15 1 9 11 1 9 4 2 4 4 2
9 15 13 1 0 9 1 10 11 2
15 8 2 12 9 3 2 7 3 3 10 0 9 1 9 2
26 3 13 9 3 4 4 2 16 12 9 10 9 4 4 1 10 9 15 10 9 10 0 9 0 13 2
34 11 13 1 10 9 1 15 9 2 7 3 3 4 15 15 0 16 15 10 0 15 9 4 16 15 0 9 15 15 3 8 13 4 2
20 10 9 13 11 3 2 7 15 4 3 11 1 13 7 15 13 15 15 3 2
19 10 9 13 7 0 13 3 10 9 1 15 3 0 1 11 8 4 4 2
13 10 9 13 15 0 10 2 0 9 2 1 4 2
17 8 10 9 13 10 9 15 9 1 10 0 9 1 10 13 9 2
34 2 15 13 15 4 1 15 0 0 0 7 0 9 1 9 7 9 2 15 15 0 9 1 11 7 1 10 9 1 10 0 9 13 2
12 9 15 9 3 10 9 1 10 9 13 2 2
23 1 10 9 1 10 11 13 10 11 4 16 10 11 16 9 1 10 0 0 9 4 4 2
21 5 10 0 9 2 3 16 0 0 2 0 7 0 9 1 10 13 9 1 4 2
15 15 4 13 2 10 0 9 2 15 4 15 3 1 4 2
17 5 9 1 10 9 1 15 9 7 9 1 10 1 11 13 9 2
8 5 0 9 1 10 0 9 2
16 5 9 1 0 9 1 11 2 1 10 11 2 1 15 8 2
4 1 0 9 2
25 8 4 3 0 1 15 9 1 10 0 9 1 9 1 8 7 3 1 8 1 10 2 11 2 2
13 3 15 2 0 13 2 1 9 4 10 0 9 2
16 15 2 8 2 7 10 2 11 2 13 15 15 1 13 3 2
42 7 15 4 1 10 9 13 10 3 0 9 1 10 0 0 9 2 3 1 9 13 9 1 10 0 9 1 15 13 5 15 13 15 3 3 5 1 10 9 4 4 2
2 11 2
22 2 7 15 13 8 1 10 9 3 2 13 15 4 8 9 15 3 1 8 4 2 2
10 7 15 13 15 0 2 15 13 13 2
18 9 1 10 11 2 10 9 1 10 11 13 3 3 1 10 15 9 2
41 16 10 9 1 10 9 4 4 4 3 3 15 0 0 9 1 10 9 4 2 7 1 10 12 9 15 0 9 1 10 11 4 4 2 13 10 9 12 9 3 2
7 10 9 11 13 15 3 2
19 3 10 9 1 11 2 1 3 13 2 4 2 16 0 1 9 2 4 2
10 3 1 12 13 10 9 10 9 3 2
27 1 11 4 1 10 13 9 10 0 9 4 2 15 4 3 3 3 10 9 16 15 13 4 4 4 2 2
2 8 2
2 11 2
2 8 2
2 11 2
17 2 6 2 1 10 9 16 15 4 10 13 9 0 1 10 9 2
2 8 2
2 11 2
9 10 9 1 8 4 3 15 0 2
26 15 13 15 0 4 16 10 9 1 0 9 2 10 9 2 3 15 3 15 9 1 10 9 13 4 2
19 15 9 3 2 16 15 9 1 10 9 1 10 9 2 9 11 2 13 2
53 3 13 10 9 3 10 0 9 3 1 2 10 0 7 0 9 2 7 13 15 10 9 3 1 15 1 2 10 9 1 4 16 15 9 1 10 13 9 3 1 4 1 15 9 1 10 9 1 3 10 9 2 2
15 0 1 10 0 2 13 9 1 13 10 0 9 15 4 2
31 1 10 9 4 10 9 1 8 3 3 10 9 2 15 9 3 3 9 2 15 13 9 3 3 9 1 10 13 9 2 2
14 15 0 8 13 3 10 0 9 4 4 1 10 11 2
17 10 9 4 10 9 1 9 1 9 7 9 8 10 9 1 9 2
40 10 0 9 2 15 15 15 9 3 1 10 0 9 13 1 10 0 9 1 11 2 13 10 9 9 1 10 9 2 15 15 13 1 10 0 9 1 12 13 2
14 1 15 9 1 10 9 1 11 13 15 10 9 8 2
16 15 13 1 15 8 7 13 16 9 8 11 2 8 7 11 2
11 15 4 10 0 9 1 10 0 9 8 2
20 1 12 13 8 15 8 7 1 12 4 15 4 1 9 1 10 9 1 8 2
25 10 0 11 4 10 9 9 2 13 1 8 2 8 2 8 2 8 2 8 8 2 8 7 8 2
25 15 13 3 10 9 1 10 9 1 12 2 7 15 13 3 16 15 3 1 10 0 9 4 4 2
44 3 13 15 3 1 10 0 9 2 15 3 3 10 0 9 4 4 1 10 5 10 0 9 5 3 0 9 2 3 11 3 3 13 4 16 15 10 9 0 4 3 1 4 2
17 3 4 15 3 2 16 10 9 13 1 10 9 1 12 1 11 2
25 1 12 13 3 10 9 1 11 2 15 1 10 0 10 9 13 1 2 8 2 2 3 10 9 2
23 7 15 9 13 3 3 1 10 9 1 10 0 9 15 0 10 9 13 1 10 0 9 2
19 8 10 9 1 9 7 9 13 10 11 3 10 9 4 1 9 7 9 2
49 2 10 0 9 15 15 3 13 4 4 10 9 1 12 0 9 1 10 0 9 8 2 15 1 10 9 9 12 7 9 12 13 4 4 7 10 9 1 10 9 1 10 9 1 12 9 1 8 2
19 10 0 9 13 1 15 13 1 15 9 2 16 15 3 9 13 4 4 2
12 15 4 1 15 9 10 9 1 11 0 9 2
11 10 9 13 3 1 10 9 1 15 8 2
13 10 9 4 11 2 10 9 4 3 10 0 9 2
7 16 1 10 0 1 13 2
14 15 4 10 9 1 11 9 7 10 9 1 15 8 2
15 11 15 13 10 9 2 7 10 8 13 9 13 15 3 2
6 15 8 13 15 13 2
21 15 13 9 3 2 15 15 13 9 0 13 16 15 10 15 9 0 1 15 13 2
11 9 7 9 3 13 3 13 1 10 9 2
9 11 13 15 13 3 7 13 3 2
25 10 9 1 15 8 13 15 13 9 2 16 9 8 1 12 9 1 10 9 3 1 9 13 4 2
26 7 3 13 11 2 1 10 0 9 1 10 9 2 0 1 9 3 1 13 3 3 10 9 1 4 2
20 11 2 15 13 1 10 0 9 1 10 9 9 12 2 13 15 3 3 4 2
16 10 9 3 4 0 3 3 1 4 16 3 10 9 1 13 2
22 11 3 2 8 9 1 9 7 0 9 2 13 8 11 3 1 10 0 9 1 11 2
14 10 0 9 8 13 10 9 1 11 1 10 9 4 2
16 10 9 1 11 1 11 4 0 4 7 10 9 13 3 3 2
15 11 13 10 9 3 4 2 7 15 0 4 3 3 0 2
6 15 13 3 15 3 2
9 9 8 13 1 10 9 10 9 2
20 11 2 1 10 9 2 13 1 10 9 1 15 9 3 3 15 8 4 4 2
2 11 2
6 15 13 3 0 9 2
8 15 13 15 10 0 9 4 2
9 15 4 3 1 10 9 1 9 2
14 10 9 8 13 9 10 9 10 0 9 15 15 13 2
9 15 13 3 3 3 10 13 9 2
10 15 9 13 13 15 1 15 9 0 2
18 2 3 13 0 3 4 4 4 16 10 9 3 1 12 9 4 4 2
17 8 2 1 15 10 0 13 0 9 2 13 13 1 11 2 11 2
16 0 9 13 15 3 3 1 11 1 15 0 13 1 10 9 2
18 1 15 9 1 10 9 1 15 8 2 13 15 0 1 15 0 9 2
11 2 15 13 15 3 4 1 15 12 9 2
9 15 13 15 0 1 10 13 9 2
5 15 13 1 9 2
29 11 13 15 9 3 3 0 16 16 15 10 9 0 0 13 7 15 10 9 13 3 1 15 9 15 3 1 4 2
10 10 9 9 4 3 1 3 12 4 2
21 0 9 1 10 9 4 10 5 8 1 10 15 0 9 5 13 9 16 10 9 2
31 10 9 2 10 0 9 1 10 9 2 13 0 9 1 0 12 2 12 2 12 2 9 3 7 13 3 15 12 12 9 2
32 1 0 9 3 4 3 4 10 9 15 10 9 13 4 1 10 0 9 2 10 0 11 2 2 15 0 0 4 16 1 12 2
24 10 0 9 4 8 1 0 9 8 2 15 1 0 9 1 15 9 2 8 2 4 13 4 2
18 16 15 9 9 13 1 15 9 1 15 9 1 4 2 4 3 0 2
12 15 13 1 15 15 9 3 1 4 4 2 2
7 10 9 13 3 15 9 2
24 15 13 8 10 9 9 2 10 0 0 9 8 4 4 1 9 1 2 0 9 1 9 2 2
12 15 9 13 9 4 1 10 9 1 10 9 2
21 15 9 4 15 2 8 2 2 16 10 9 15 1 10 9 2 8 2 13 4 2
7 15 4 3 10 0 9 2
9 8 3 1 10 9 13 1 4 2
6 8 13 10 0 9 2
14 15 13 4 16 15 1 15 9 9 3 0 9 4 2
13 10 0 9 1 10 9 13 15 3 3 1 4 2
8 7 15 4 15 0 3 3 2
4 5 7 3 2
7 16 13 1 10 0 9 2
13 7 9 0 13 3 15 9 16 3 8 1 4 2
23 1 11 4 15 0 3 2 16 15 1 10 9 13 4 2 1 10 9 7 9 1 13 2
12 15 4 1 10 9 7 10 0 9 4 2 2
29 3 13 10 9 1 10 9 7 0 9 3 3 3 4 2 15 13 16 10 9 0 10 9 1 10 0 9 4 2
5 2 15 13 3 2
17 8 13 3 15 8 2 10 9 1 12 9 1 0 9 2 4 2
12 11 13 10 9 3 1 12 9 7 12 9 2
36 1 10 9 2 3 10 9 11 7 11 0 13 4 2 4 10 9 1 10 9 4 1 8 2 11 2 11 2 11 2 11 2 11 7 11 2
13 1 15 9 13 8 15 1 10 9 3 10 0 2
2 11 2
10 10 9 11 4 0 1 11 7 11 2
13 10 0 9 13 7 1 0 7 9 10 0 9 2
8 10 0 0 9 4 3 4 2
16 10 9 15 3 15 3 13 2 13 15 15 9 8 1 4 2
9 3 4 3 9 1 15 0 4 2
23 15 13 0 0 4 16 1 10 9 1 8 12 9 2 0 0 9 7 9 2 1 4 2
17 10 0 9 0 12 9 2 13 3 8 4 4 2 3 13 15 2
13 3 13 15 15 13 16 1 4 1 10 9 3 2
22 2 3 1 15 9 2 2 3 10 9 2 2 13 11 15 0 9 16 9 4 2 2
22 1 9 13 10 9 3 9 4 4 7 9 1 9 16 9 2 7 1 15 0 9 2
18 2 15 13 16 15 0 4 4 1 10 9 15 15 8 9 13 4 2
4 1 0 9 2
24 8 13 1 10 9 4 2 16 15 1 15 8 2 16 8 2 10 11 1 11 13 4 4 2
16 15 9 2 13 10 9 3 2 13 10 9 1 0 12 9 2
6 3 4 15 3 4 2
20 7 3 1 12 9 4 10 9 1 3 1 0 4 1 0 9 7 9 3 2
18 10 9 1 10 9 13 15 9 15 15 4 4 1 10 3 0 9 2
23 10 9 1 10 9 1 10 0 9 4 4 2 7 10 9 1 10 9 4 10 0 9 2
17 10 0 9 13 3 1 12 2 12 2 12 1 0 12 12 9 2
15 10 13 9 13 1 12 2 12 2 12 1 0 12 12 2
20 1 10 13 9 4 10 9 10 9 0 15 3 0 3 16 1 12 13 4 2
37 3 13 15 1 10 9 3 15 13 9 16 15 9 2 15 9 2 15 9 7 15 9 2 16 3 0 10 9 9 3 1 4 13 4 2 8 2
23 15 1 8 2 0 9 2 4 7 1 8 2 0 9 2 2 13 8 2 0 9 2 2
45 11 13 15 16 2 10 9 2 15 3 0 13 7 13 2 1 15 15 15 1 10 15 1 4 4 2 7 15 3 15 0 1 15 0 13 7 0 1 10 15 2 3 13 2 2
17 15 9 1 15 8 13 8 1 9 4 1 10 0 7 13 9 2
21 9 12 1 10 9 13 16 1 9 1 9 1 0 9 10 0 9 4 4 4 2
7 10 0 9 13 4 4 2
59 10 9 13 10 9 1 10 9 7 10 3 13 9 1 10 9 1 10 9 2 13 1 10 9 0 9 3 1 10 11 2 8 1 15 9 15 5 1 9 1 10 9 1 10 9 5 9 1 10 3 1 10 0 9 13 9 4 4 2
7 10 0 9 13 0 4 2
20 1 10 9 1 10 1 9 15 9 13 11 3 3 0 9 8 3 15 9 2
5 15 0 13 15 2
7 2 1 11 13 15 4 2
15 15 4 10 15 9 7 15 13 3 1 12 9 4 2 2
5 3 13 15 8 2
13 1 10 0 9 13 15 1 15 0 9 8 2 2
42 10 9 1 12 1 10 1 9 0 0 9 13 11 3 3 15 4 2 16 9 13 1 10 15 9 15 9 15 3 1 4 1 15 0 12 1 10 0 9 1 9 2
11 1 10 11 4 12 10 9 1 13 9 2
12 10 9 13 1 12 9 1 3 12 12 9 2
50 10 0 9 4 12 9 0 7 13 12 2 12 2 12 9 2 16 10 9 0 13 2 1 12 9 2 13 10 9 0 12 9 0 3 1 12 2 12 2 12 3 4 4 12 2 12 2 12 9 2
16 10 9 4 16 0 4 1 8 2 12 2 1 9 1 8 2
17 3 16 15 10 9 15 13 4 4 2 7 10 9 13 0 4 2
15 7 9 2 9 7 9 4 3 3 10 13 2 0 9 2
27 13 15 3 1 10 9 1 10 9 2 0 1 9 7 1 10 9 10 9 1 10 9 3 3 1 4 2
17 0 13 1 11 1 10 9 1 15 0 1 9 13 9 4 4 2
17 10 9 8 2 12 2 0 9 1 11 2 3 0 1 10 9 2
33 15 0 9 1 9 7 10 9 1 10 13 9 1 11 1 15 8 2 10 9 1 11 2 10 9 1 11 2 10 9 1 8 2
26 7 0 3 13 12 9 8 10 9 1 10 1 9 7 9 13 9 15 15 8 13 2 1 10 9 2
6 7 11 13 13 9 2
6 10 9 4 13 4 2
6 10 9 13 9 4 2
7 10 9 11 4 3 4 2
2 9 2
4 4 15 13 2
2 9 2
2 6 2
13 2 15 4 0 15 3 1 10 9 15 1 4 2
38 7 1 10 9 16 8 3 1 10 9 1 10 9 10 9 4 2 4 10 9 2 1 10 9 1 10 0 9 3 2 4 1 9 15 0 0 4 2
11 15 0 13 8 1 10 9 1 10 0 2
15 3 10 0 15 9 13 13 15 10 0 9 1 10 0 2
33 1 10 9 1 10 9 1 11 13 10 9 1 10 3 3 10 9 13 9 2 8 2 16 10 9 9 1 10 9 4 4 4 2
25 4 4 16 3 3 3 9 4 4 1 0 9 7 15 1 10 9 1 9 7 9 7 10 9 2
14 3 15 0 2 0 8 13 15 1 3 12 9 0 2
5 15 13 1 8 2
10 16 10 9 13 15 15 1 11 0 2
11 3 13 11 1 10 0 9 10 0 9 2
18 10 0 9 1 11 4 0 1 10 9 1 11 2 3 11 13 4 2
16 3 13 15 10 9 1 9 3 0 2 3 1 15 12 9 2
20 15 4 3 3 8 15 0 1 9 1 4 2 3 9 8 13 9 13 4 2
18 15 9 13 3 1 9 7 9 2 15 15 1 9 3 0 0 13 2
7 1 9 13 15 15 4 2
7 15 13 1 10 0 9 2
22 1 10 9 10 9 13 15 9 4 1 9 1 9 1 0 7 9 7 0 9 4 2
14 15 9 3 13 15 10 0 9 8 10 13 9 9 2
23 16 15 1 15 8 3 0 13 1 4 2 13 10 9 1 10 0 9 1 15 9 3 2
28 10 8 13 9 4 4 7 10 9 16 10 9 1 11 10 9 4 2 13 10 9 1 10 9 10 9 3 2
19 7 13 9 11 9 8 1 10 9 1 2 0 16 15 3 3 4 4 2
19 16 10 9 1 13 13 15 9 1 15 0 9 2 9 7 0 9 4 2
21 3 3 4 3 1 11 10 9 1 0 7 0 9 1 10 9 10 9 1 4 2
24 10 10 9 7 9 13 10 9 1 15 3 0 9 1 15 9 3 3 1 0 7 0 9 2
22 3 13 15 16 10 0 9 1 10 9 7 1 10 9 15 15 0 1 15 9 13 2
15 3 15 0 0 4 10 9 1 8 2 11 2 8 2 2
36 10 9 13 10 9 3 9 1 10 9 1 9 4 4 2 10 9 13 10 9 1 10 9 2 2 15 13 3 10 0 2 13 2 13 9 2
20 16 10 9 3 7 3 0 13 5 15 0 9 4 5 13 15 0 10 9 2
16 10 9 1 10 9 7 10 0 9 1 10 9 1 10 9 2
24 9 11 2 11 11 2 13 0 1 10 9 10 9 1 10 0 13 9 8 2 3 1 4 2
31 16 3 15 0 9 13 1 10 9 1 10 9 1 10 9 2 13 10 9 11 1 10 11 2 3 13 15 13 9 4 2
14 7 2 13 15 3 4 2 15 9 13 15 3 3 2
17 1 10 9 13 3 3 10 9 8 3 10 9 3 1 4 13 2
15 11 13 3 1 9 2 16 15 10 9 1 15 9 13 2
3 11 3 2
9 2 15 13 15 9 2 13 11 2
17 7 16 15 1 10 0 9 13 2 13 15 3 1 10 0 9 2
12 7 3 13 15 3 10 9 16 1 4 2 2
12 1 10 0 9 13 11 1 11 15 9 3 2
18 15 13 9 1 11 2 1 10 13 9 13 2 4 3 10 9 3 2
18 7 1 11 13 10 13 2 0 2 1 11 3 1 10 9 4 4 2
13 16 15 3 13 13 15 1 15 9 3 4 4 2
12 15 13 1 9 2 16 10 9 15 0 4 2
7 9 2 9 2 11 2 2
10 15 4 0 0 5 3 3 10 9 2
18 16 15 15 1 10 9 3 10 9 13 4 2 3 13 15 15 4 2
7 3 13 15 3 0 4 2
8 7 3 13 15 3 4 2 2
22 11 4 3 3 0 1 15 12 1 10 9 2 16 13 15 3 10 9 3 3 4 2
11 2 1 10 9 4 10 9 1 3 4 2
26 9 11 13 15 9 7 13 10 9 1 10 0 9 2 1 15 9 8 9 11 0 13 2 12 2 2
48 3 4 10 9 1 9 4 16 16 10 9 3 13 9 3 13 1 4 2 16 8 10 9 1 11 1 10 9 13 2 7 11 13 3 15 9 10 9 1 10 0 9 1 10 9 1 4 2
18 15 13 10 9 3 4 7 1 12 9 13 11 1 10 0 9 3 2
7 7 8 2 0 7 0 2
12 8 2 10 0 9 1 8 2 13 16 9 2
15 2 15 13 3 10 9 4 1 10 9 16 15 4 4 2
5 3 3 1 11 2
16 16 15 13 13 15 3 10 9 16 15 3 3 15 3 4 2
6 7 15 4 9 2 2
17 11 13 1 15 9 1 10 13 12 9 12 9 4 4 1 11 2
16 10 3 0 9 2 3 16 13 11 10 15 0 9 16 11 2
21 3 1 10 0 9 13 11 15 10 0 9 4 1 10 3 3 13 9 1 11 2
9 1 10 9 13 3 9 1 11 2
19 8 7 11 13 3 1 9 2 15 1 3 1 15 0 9 13 1 11 2
28 1 10 9 1 11 13 3 3 9 8 1 10 0 9 1 10 9 9 4 1 10 0 9 1 10 0 9 2
11 2 0 16 15 1 10 0 9 4 4 2
3 11 13 2
23 7 9 8 1 10 0 9 13 0 16 15 10 9 4 1 10 9 3 11 15 9 13 2
18 2 15 13 3 3 10 9 16 15 0 4 16 15 10 9 8 4 2
21 0 4 3 9 4 2 7 16 15 3 13 4 4 3 0 15 10 13 4 2 2
33 10 9 13 1 9 1 10 9 4 2 16 10 9 1 8 4 4 2 16 10 9 13 7 1 10 9 9 13 3 1 4 2 2
16 10 9 13 15 1 10 0 7 0 9 3 3 1 9 4 2
17 15 9 3 16 1 15 1 4 7 15 13 9 7 9 1 4 2
4 15 4 13 2
13 1 12 13 10 9 3 2 16 8 12 9 4 2
15 10 9 2 3 9 1 10 9 3 3 1 9 13 4 2
13 15 13 0 9 16 15 4 4 16 3 4 4 2
22 15 0 8 5 1 12 9 10 9 1 15 13 1 12 9 5 13 3 10 15 9 2
3 9 4 2
15 8 13 1 15 2 16 15 13 1 9 15 10 9 4 2
24 10 9 15 1 10 11 13 2 15 4 3 15 12 2 13 12 9 1 10 9 0 1 9 2
18 13 15 1 10 9 3 13 15 12 9 0 2 1 10 9 12 9 2
18 15 15 9 3 1 10 0 9 13 4 13 10 9 1 15 9 8 2
5 7 8 13 15 2
19 10 9 11 13 15 9 1 10 9 4 3 12 9 1 10 9 4 4 2
21 1 10 9 1 10 11 4 3 12 0 4 15 1 9 1 9 7 9 4 4 2
8 15 13 3 3 10 9 4 2
15 15 13 3 1 15 4 15 9 1 10 0 9 1 4 2
15 15 12 1 15 9 4 0 3 1 15 9 1 0 4 2
8 3 4 15 9 7 9 4 2
12 10 9 7 9 13 15 10 9 3 3 4 2
33 10 0 9 1 10 9 1 10 9 8 2 0 11 2 13 3 4 1 10 9 1 9 7 9 1 10 11 2 1 15 10 9 2
20 10 9 13 16 10 9 15 9 1 10 9 13 16 10 0 9 8 1 13 2
31 10 9 2 15 0 8 2 7 10 9 2 15 0 8 2 12 1 11 0 2 13 4 16 10 9 1 10 9 15 4 2
4 7 3 8 2
9 15 9 4 1 15 0 0 4 2
32 7 10 9 15 3 1 8 1 8 13 2 15 13 3 3 15 8 1 15 0 9 2 15 13 3 4 10 0 12 9 3 2
14 3 13 15 15 2 7 15 4 0 13 10 0 9 2
6 9 13 15 3 2 2
20 3 13 3 10 9 3 8 4 2 2 3 8 2 0 0 1 10 0 9 2
12 10 12 0 9 13 8 3 0 3 3 3 2
19 15 13 10 9 2 16 15 3 3 10 3 0 9 3 4 2 1 11 2
24 1 9 1 15 9 13 15 1 10 0 9 3 1 11 3 15 10 9 1 10 9 13 4 2
16 10 15 9 1 10 0 9 4 10 0 9 1 9 1 9 2
8 2 3 4 0 15 4 2 2
22 1 11 4 15 3 3 0 16 3 1 10 13 12 9 10 9 4 4 1 0 9 2
21 2 15 13 3 15 0 9 2 15 0 9 2 3 13 10 0 9 4 4 2 2
29 1 12 13 11 2 3 11 3 8 13 2 10 0 9 1 10 9 3 2 3 10 0 9 1 2 11 2 13 2
11 0 13 16 9 4 15 9 10 0 9 2
18 3 13 3 11 1 10 9 1 11 2 3 10 0 2 11 2 13 2
12 15 13 10 9 11 15 9 16 9 10 9 2
16 8 13 2 16 15 13 1 10 13 9 15 9 1 9 4 2
12 8 2 9 1 10 0 9 2 13 8 9 2
7 9 1 0 2 0 9 2
7 10 9 13 15 9 3 2
4 15 4 9 2
51 2 10 0 9 15 10 9 13 1 10 9 1 15 15 3 13 4 13 3 1 10 9 2 7 10 0 9 15 1 0 9 4 2 4 3 10 9 1 9 2 2 13 10 9 8 2 9 1 15 8 2
31 2 0 2 2 13 9 8 2 12 2 2 0 9 1 8 2 2 13 10 0 9 3 9 1 10 9 1 15 9 2 2
26 10 13 9 4 3 2 16 15 9 15 1 10 9 1 9 4 4 1 10 9 1 10 0 9 13 2
17 15 4 0 16 10 3 13 9 3 3 1 0 9 1 13 13 2
7 10 13 9 4 3 4 2
13 3 3 1 10 9 2 7 15 13 12 13 9 2
24 10 9 1 10 9 2 15 13 1 10 15 13 9 3 10 9 0 9 2 4 3 0 13 2
12 10 9 1 10 1 12 13 9 13 3 3 2
33 1 10 9 1 10 0 9 13 10 0 9 8 2 15 1 10 9 1 15 9 9 13 1 10 9 2 1 1 15 9 0 9 2
30 15 13 16 1 10 13 9 2 3 10 9 15 3 13 13 1 10 15 0 9 2 10 9 1 10 11 3 4 4 2
13 10 9 1 10 9 13 1 8 0 4 4 4 2
12 3 13 10 9 1 3 12 12 9 0 4 2
61 16 10 9 1 10 9 3 13 2 13 10 9 1 10 13 12 9 9 4 1 10 0 9 1 10 9 1 10 0 9 1 9 2 15 8 10 0 9 1 10 9 1 10 0 9 2 3 12 9 1 10 9 2 16 11 1 13 4 1 4 2
17 10 0 9 11 13 10 9 1 10 9 1 15 8 1 11 4 2
11 9 4 4 1 10 9 1 10 13 9 2
18 3 10 9 13 11 0 9 0 9 8 10 9 1 11 7 1 11 2
12 2 15 13 15 0 16 10 0 9 1 4 2
14 10 9 1 15 0 0 9 1 9 13 3 4 4 2
16 1 11 1 11 7 2 8 2 1 11 13 3 0 12 9 2
8 10 9 13 3 12 12 9 2
41 3 4 1 15 9 10 0 9 4 1 10 9 2 3 3 16 10 9 1 11 3 3 15 9 4 1 4 2 7 13 9 2 3 10 9 0 1 10 9 13 2
16 2 0 2 2 2 9 2 7 2 9 2 4 10 9 9 2
13 1 15 0 9 16 8 13 10 9 12 1 8 2
21 11 2 0 16 9 7 3 3 16 9 2 13 1 11 10 9 1 10 9 0 2
40 7 1 10 11 13 15 1 10 16 12 9 7 1 9 15 1 9 13 4 4 2 13 15 9 1 10 9 15 1 10 9 1 9 13 3 16 3 1 4 2
50 10 9 13 15 2 15 9 15 1 15 0 9 4 13 2 16 1 10 9 0 9 3 15 13 1 10 9 13 1 9 2 9 7 9 2 2 13 2 1 0 9 2 10 0 9 4 4 7 4 2
9 0 13 13 9 7 4 15 9 2
14 3 13 3 3 2 16 12 15 9 9 1 9 13 2
14 0 13 13 13 10 9 3 7 13 15 0 3 4 2
23 3 15 0 2 0 13 2 15 3 9 3 15 9 13 2 13 10 9 3 1 15 4 2
11 7 3 13 10 0 9 0 1 0 9 2
8 0 13 2 9 2 0 9 2
11 15 9 13 1 9 1 0 9 4 4 2
20 1 15 4 10 9 3 0 2 16 15 0 4 4 7 1 10 13 9 13 2
14 16 15 12 13 13 3 3 12 9 1 0 9 13 2
26 10 9 9 13 0 1 9 2 1 10 9 1 10 9 13 3 1 10 9 1 0 3 10 15 9 2
19 9 1 0 9 2 13 13 7 15 9 2 1 15 12 2 0 3 0 2
3 9 3 2
29 3 13 15 9 15 0 10 0 9 13 2 3 3 0 16 3 9 13 15 15 0 13 16 1 10 9 1 4 2
25 2 1 10 9 2 2 13 9 0 3 2 2 13 15 3 0 9 13 1 10 9 1 10 9 2
16 16 10 9 13 3 10 0 9 10 0 9 4 1 15 9 2
7 15 0 9 8 13 4 2
2 9 2
16 13 7 13 7 3 10 9 0 1 15 13 16 16 1 13 2
5 3 4 10 9 2
30 9 13 3 3 1 16 15 10 9 1 15 9 4 2 16 3 0 15 9 4 16 1 15 9 0 15 9 1 4 2
22 15 4 0 3 0 10 0 9 1 13 2 16 10 9 1 10 0 3 3 0 4 2
24 1 0 9 13 9 12 9 2 9 13 1 12 9 2 12 9 7 9 13 3 12 9 3 2
24 9 13 2 0 2 1 10 0 9 3 2 15 9 1 10 9 13 4 7 10 9 4 0 2
7 11 13 3 0 0 9 2
23 13 4 15 3 15 1 10 9 8 15 1 10 1 15 9 13 9 1 10 9 3 4 2
28 3 13 8 2 15 10 9 1 10 9 13 2 9 4 4 1 10 9 16 15 10 9 3 1 15 9 4 2
14 8 13 15 15 1 10 13 9 1 0 9 7 9 2
11 15 13 15 9 3 3 0 7 0 0 2
18 1 10 0 9 1 10 9 1 11 13 13 8 2 12 2 15 0 2
61 11 2 0 3 3 0 2 1 10 9 15 13 11 1 10 0 9 1 10 9 13 2 13 15 15 9 3 0 10 9 1 10 0 9 2 9 2 9 7 3 9 8 16 1 9 1 13 16 15 0 15 1 13 4 4 1 10 15 8 9 2
7 2 15 4 15 0 9 2
25 8 10 0 11 7 10 9 8 2 11 2 4 1 12 8 12 10 9 4 8 10 0 9 12 2
20 16 2 9 2 4 10 9 2 8 2 4 2 3 9 4 4 1 3 8 2
8 8 2 8 2 8 7 8 2
11 15 4 9 1 9 1 10 0 0 9 2
23 15 15 1 10 9 1 8 1 9 13 13 10 9 0 2 7 15 4 3 1 9 0 2
20 0 16 15 9 3 4 10 9 2 15 3 10 9 13 7 15 9 9 13 2
52 10 0 9 1 10 9 1 9 2 10 9 8 2 13 10 9 1 10 9 1 10 0 0 0 9 1 11 10 2 0 0 9 2 2 15 3 0 13 7 3 10 9 13 16 1 15 9 16 9 7 9 2
28 10 9 11 13 10 9 1 10 9 3 1 13 1 10 9 9 1 11 2 15 3 4 4 1 12 1 9 2
9 10 9 4 16 15 0 0 4 2
36 3 13 15 10 9 1 10 0 9 16 1 15 9 3 3 1 15 9 7 1 10 9 1 9 7 9 4 4 4 4 15 15 4 4 4 2
32 15 13 4 0 7 1 10 9 16 15 1 4 4 1 10 9 15 13 1 9 1 4 3 0 9 1 9 7 0 9 4 2
16 1 10 9 13 8 16 9 1 10 9 0 4 8 10 9 2
20 10 9 1 9 7 9 13 10 0 9 1 4 1 10 0 13 9 7 9 2
12 10 0 9 3 13 1 15 9 4 4 4 2
14 15 0 9 13 15 1 10 9 4 16 9 1 9 2
16 10 9 13 15 0 9 4 4 1 15 1 0 9 13 4 2
4 15 9 4 2
10 13 3 10 0 9 1 10 9 4 2
9 4 10 9 0 10 9 1 4 2
13 15 13 15 1 10 9 3 0 13 13 4 2 2
11 10 0 9 1 8 7 8 13 1 12 2
10 10 9 13 16 9 1 10 0 9 2
9 3 13 8 10 9 4 7 4 2
19 13 9 4 12 9 1 10 0 9 7 12 9 1 10 9 1 15 8 2
16 15 0 9 4 4 1 15 1 12 9 2 15 16 9 13 2
14 1 11 4 15 8 2 16 11 10 0 9 4 4 2
32 11 13 15 3 1 10 0 9 11 3 4 1 10 0 9 1 10 11 16 1 10 0 9 1 9 12 11 1 12 1 13 2
9 10 9 1 10 0 9 4 13 2
25 1 10 9 16 10 9 1 8 1 10 0 9 3 1 10 0 9 1 4 2 13 15 10 9 2
17 8 2 10 9 1 10 9 8 2 13 3 1 10 9 1 8 2
2 12 2
23 1 10 9 1 15 12 9 1 10 9 4 15 3 1 10 0 9 0 10 9 1 13 2
43 8 15 9 1 0 9 16 10 9 1 9 11 1 11 1 10 9 1 4 4 2 4 11 3 3 3 4 9 11 7 11 0 9 8 1 9 1 10 9 11 1 4 2
23 10 9 1 9 13 15 3 10 9 1 10 9 1 10 9 1 9 1 10 9 1 4 2
8 3 4 3 10 0 9 4 2
17 9 11 13 15 2 16 10 0 9 1 15 8 3 4 4 4 2
14 3 13 8 3 4 16 10 9 9 0 1 11 4 2
20 15 4 3 11 9 10 9 1 13 2 15 10 9 11 7 15 9 13 4 2
31 16 15 9 13 4 1 10 0 9 2 13 10 11 10 9 4 16 1 10 0 9 1 10 9 1 4 2 13 10 9 2
26 3 13 15 0 9 1 8 1 10 9 16 10 0 9 1 15 1 8 13 8 3 3 3 4 4 2
18 10 9 1 11 13 3 10 9 1 0 12 9 0 1 9 1 8 2
16 3 1 10 9 1 10 9 1 11 1 8 13 10 0 9 2
29 2 3 8 8 13 0 9 8 1 8 2 10 9 11 7 1 0 7 0 9 2 1 7 0 1 10 9 11 2
41 10 9 1 10 9 2 10 9 8 2 13 3 3 16 10 9 12 1 10 3 12 9 4 2 1 15 12 3 15 13 4 3 0 1 10 9 13 1 4 4 2
15 1 15 12 4 3 12 0 16 12 9 1 10 9 4 2
24 1 10 0 12 9 2 15 4 4 2 13 3 12 2 15 0 16 12 9 1 15 8 13 2
20 10 9 1 10 9 1 8 2 1 11 2 4 10 0 9 1 12 9 4 2
7 10 9 4 15 16 13 2
11 8 4 3 0 4 2 16 15 9 13 2
16 10 9 4 8 10 9 1 10 3 13 9 1 11 16 9 2
5 10 9 4 4 2
23 1 15 9 13 10 9 10 0 9 1 10 9 1 10 9 8 7 8 10 3 0 9 2
14 10 9 1 12 4 4 1 12 12 9 1 12 12 2
15 10 9 1 10 9 8 13 3 3 3 12 1 12 9 2
11 10 9 1 11 4 1 15 9 3 4 2
11 10 9 11 13 3 3 3 0 16 8 2
13 10 0 9 13 8 0 3 3 3 1 15 9 2
32 10 9 1 10 11 4 3 3 4 16 1 10 9 1 11 12 9 1 13 9 1 15 13 1 9 12 0 1 10 0 13 2
9 1 10 9 8 11 13 15 8 2
9 9 11 4 3 3 10 9 3 2
20 15 13 16 15 8 10 13 9 4 1 10 0 9 1 15 8 2 13 15 2
17 1 10 9 13 3 15 9 12 1 12 9 7 9 1 15 8 2
23 16 15 1 10 0 9 2 15 8 8 13 2 13 3 15 1 10 0 9 0 10 4 2
21 11 13 16 3 10 9 4 16 3 1 4 16 10 11 10 9 3 0 4 4 2
13 10 9 13 16 10 11 3 4 1 9 1 11 2
21 10 11 13 1 10 9 1 10 9 7 10 0 9 3 3 15 9 2 3 11 2
30 10 9 13 1 0 9 1 10 9 2 7 3 10 9 4 4 4 2 16 10 9 13 0 1 10 11 3 1 4 2
24 10 9 9 16 3 3 3 0 13 16 15 1 15 9 7 3 11 12 9 3 3 9 4 2
22 10 0 13 10 9 3 2 16 15 0 1 15 9 0 0 4 16 1 10 9 3 2
4 15 13 3 2
9 15 13 10 9 0 7 0 3 2
8 15 9 13 3 1 10 9 2
17 0 2 10 11 4 8 3 1 10 9 2 15 15 16 9 13 2
14 15 9 2 11 2 13 15 1 10 9 3 0 0 2
33 10 9 1 11 1 8 16 9 13 10 0 9 2 12 2 1 10 9 1 12 9 2 8 2 1 10 0 0 9 1 15 8 2
17 10 9 1 11 2 12 2 7 11 2 12 2 4 0 7 0 2
43 1 10 15 9 13 15 3 3 16 3 1 4 2 15 1 10 0 9 10 9 4 4 2 3 13 15 0 13 1 10 0 12 9 10 9 1 12 2 12 7 15 9 2
19 15 13 3 3 4 1 8 2 15 15 9 10 9 3 1 11 4 13 2
30 9 1 10 9 1 11 13 15 10 9 1 10 0 9 1 11 2 3 10 9 1 10 9 0 4 2 10 9 11 2
9 15 13 3 9 4 2 13 15 2
26 16 10 0 9 3 4 4 2 13 3 9 3 2 15 3 3 3 0 2 3 3 3 3 0 4 2
5 7 11 13 15 2
21 10 9 4 3 4 15 3 0 3 1 4 1 10 9 1 0 9 1 10 9 2
17 16 10 9 3 10 0 9 3 13 3 13 15 3 0 9 4 2
31 0 13 10 9 11 15 1 10 9 1 10 0 9 11 2 16 10 0 9 1 11 3 1 10 11 9 4 4 1 11 2
11 2 15 13 0 3 2 15 0 13 2 2
15 15 8 13 3 1 0 9 12 9 0 10 0 9 4 2
26 10 9 1 11 4 1 8 12 3 0 4 8 10 9 7 9 1 10 0 9 1 10 11 1 11 2
15 1 10 9 8 4 9 3 10 9 0 0 1 15 9 2
12 10 3 13 9 13 1 9 1 3 12 9 2
39 10 11 13 1 15 9 15 13 9 1 9 2 15 1 10 0 9 3 3 9 8 4 4 16 1 9 1 10 0 9 7 8 1 11 2 1 4 4 2
18 0 4 4 10 9 1 10 9 1 11 1 10 9 11 3 1 4 2
10 15 4 10 9 1 10 0 15 9 2
16 10 13 9 4 10 9 1 10 11 1 10 0 9 11 4 2
21 7 10 0 9 13 3 3 1 10 11 9 3 10 9 13 3 15 1 9 4 2
26 16 9 1 10 0 9 13 9 1 4 1 15 9 2 0 2 1 10 9 15 15 13 1 10 11 2
18 7 16 15 3 0 4 4 16 9 1 13 1 0 9 13 9 3 2
16 2 16 15 13 13 13 15 16 15 1 10 9 4 4 2 2
33 16 15 15 15 9 3 13 1 4 1 15 8 13 1 10 0 9 9 12 2 13 15 15 3 4 8 9 15 11 1 4 4 2
12 3 2 15 13 15 9 10 0 9 1 4 2
25 15 4 15 9 16 3 3 3 10 9 1 11 1 2 13 2 2 7 10 0 9 1 12 9 2
17 10 0 9 4 3 1 10 9 1 15 9 3 3 1 3 4 2
7 15 4 0 16 3 2 2
2 9 2
14 11 13 15 3 3 2 16 15 10 0 9 8 4 2
23 2 16 15 10 9 13 4 2 1 15 12 0 9 1 11 2 13 15 10 9 1 11 2
13 1 15 0 9 13 15 3 3 3 1 15 9 2
6 3 13 15 3 4 2
9 3 13 15 1 15 9 3 3 2
20 3 13 0 2 0 9 4 2 15 10 9 13 7 3 13 15 1 10 9 2
4 1 9 13 2
25 1 10 0 11 13 10 0 9 9 15 1 10 9 1 15 9 0 4 1 10 9 1 15 9 2
29 2 15 8 13 4 10 0 9 1 15 9 1 4 16 3 10 0 9 1 4 2 2 3 10 9 1 10 9 2
20 3 10 9 15 13 10 9 8 7 10 9 13 1 15 9 3 15 9 4 2
11 10 0 9 13 3 10 0 9 1 15 2
30 10 0 9 13 1 10 0 9 7 1 13 9 10 9 1 10 9 3 4 7 10 2 9 2 10 2 9 2 4 2
13 11 13 1 10 0 9 10 9 1 15 13 4 2
14 3 13 10 3 0 9 1 9 2 9 7 0 9 2
13 0 10 9 1 9 7 9 13 15 9 3 0 2
22 15 13 3 1 15 8 2 15 3 1 15 8 4 4 2 11 12 7 12 11 2 2
35 10 0 9 1 10 0 9 2 11 2 13 3 15 9 10 9 4 16 10 0 9 13 4 1 10 9 7 10 9 1 10 9 1 11 2
20 1 10 11 11 9 13 10 9 2 16 11 1 0 9 1 10 11 4 4 2
32 11 13 1 10 9 10 0 9 1 10 9 3 2 15 3 1 9 4 1 10 9 1 10 11 2 15 11 10 9 13 4 2
17 1 11 4 15 3 1 10 9 4 2 16 15 9 3 4 4 2
13 10 9 13 15 3 1 10 9 1 10 13 9 2
35 15 2 8 2 13 15 0 16 2 10 0 9 2 0 1 15 9 2 2 15 1 10 9 2 15 9 13 15 9 1 9 1 13 2 2
25 10 13 9 4 3 0 3 15 8 10 9 0 1 4 2 7 3 3 16 13 9 0 1 4 2
33 10 15 9 2 11 2 13 3 10 9 9 2 7 13 1 10 9 3 13 0 1 4 2 16 3 15 9 10 15 13 9 13 2
11 3 10 0 9 1 10 11 4 3 0 2
20 3 1 10 9 1 10 11 7 10 9 1 11 4 10 9 1 9 3 0 2
41 1 9 4 4 16 10 9 3 0 12 9 1 0 9 13 2 16 10 9 9 1 10 15 9 1 10 9 2 16 11 4 4 2 0 3 12 1 0 9 13 2
13 10 9 13 1 10 9 1 12 8 12 0 3 2
12 10 9 0 9 1 15 9 13 1 12 12 2
7 1 12 4 15 9 12 2
22 8 15 9 13 1 12 5 13 1 10 9 1 12 9 1 10 9 5 12 9 8 2
15 13 1 12 2 12 0 2 13 15 10 9 1 12 9 2
19 3 3 10 9 13 3 10 13 9 0 1 10 3 0 13 9 1 11 2
10 15 9 4 1 15 8 1 15 8 2
19 10 9 1 10 9 1 12 13 4 4 1 10 0 9 1 10 0 9 2
7 9 13 1 10 9 3 2
56 10 9 1 11 13 7 15 9 3 13 13 2 3 0 0 15 0 0 9 4 16 15 3 1 10 0 9 1 15 8 13 2 10 9 2 3 10 9 3 1 9 13 7 15 3 0 4 16 15 0 1 10 9 4 4 2
8 7 3 13 15 11 0 4 2
17 10 9 13 9 1 9 1 10 9 7 0 0 9 1 10 9 2
31 9 8 13 4 1 10 0 9 1 0 3 1 13 9 7 9 2 7 15 3 1 10 9 13 2 4 1 10 9 13 2
22 10 9 1 15 8 13 0 9 8 8 2 7 4 1 10 9 0 0 1 15 9 2
13 1 10 9 13 8 1 1 15 9 1 9 11 2
14 15 13 1 9 4 9 2 3 4 15 0 3 2 2
9 13 0 10 0 9 1 10 9 2
16 10 9 4 0 3 10 9 16 10 0 0 0 2 0 9 2
32 15 9 9 4 13 3 3 4 4 16 15 8 5 15 13 0 16 15 8 3 15 3 1 13 4 5 12 9 9 4 4 2
11 16 3 12 9 4 4 7 12 0 9 2
22 8 2 15 1 10 9 1 10 9 2 4 0 8 1 15 8 15 0 13 1 4 2
12 10 9 1 10 9 4 4 8 10 0 9 2
3 4 4 2
27 10 9 1 10 9 1 8 2 15 0 9 7 10 9 1 10 9 1 10 9 7 10 9 1 10 9 2
13 10 9 2 8 2 4 1 10 0 4 1 12 2
4 9 11 13 2
21 2 10 0 4 1 10 0 9 4 1 10 9 1 10 9 1 10 0 12 9 2
16 10 8 13 9 13 3 1 10 9 1 11 12 0 9 4 2
52 0 13 13 15 1 15 13 9 1 9 3 3 16 15 1 15 0 9 7 1 10 15 1 10 9 13 9 15 4 3 15 10 0 9 1 10 9 13 1 4 4 16 10 0 9 15 13 4 1 10 9 2
28 15 1 10 9 4 1 9 7 9 1 10 9 4 2 10 15 4 3 1 9 4 7 13 3 1 9 4 2
30 10 9 4 4 1 10 0 9 1 8 2 15 1 10 9 10 9 3 15 9 4 7 1 10 9 1 10 9 13 2
29 1 11 13 3 2 15 15 13 13 2 3 10 9 11 8 0 10 9 1 12 0 9 8 4 4 1 10 9 2
11 15 3 1 9 13 9 4 9 3 4 2
16 10 9 4 3 0 1 10 9 9 4 2 3 13 10 9 2
8 0 13 11 10 9 1 9 2
19 10 9 4 3 3 4 7 4 3 4 2 7 15 4 3 3 0 4 2
49 10 9 1 10 9 13 4 2 16 10 9 15 4 4 3 10 15 9 1 10 9 2 16 10 9 4 2 1 4 2 8 10 9 7 16 15 0 10 9 13 8 16 10 9 1 10 0 9 2
17 3 1 10 0 13 10 0 9 15 0 1 10 9 3 4 4 2
18 2 15 13 3 10 9 1 8 7 15 13 1 9 15 9 1 9 2
23 16 1 13 4 15 11 2 15 15 1 10 2 0 2 0 7 0 9 2 8 13 4 2
35 12 0 9 3 10 0 9 1 10 0 9 2 4 2 3 16 1 11 10 9 13 16 11 1 15 8 1 13 2 1 15 9 4 4 2
18 15 13 10 9 4 15 15 1 15 9 1 11 13 1 15 1 11 2
10 7 15 13 2 0 13 2 1 4 2
21 10 12 9 2 10 0 2 10 0 7 10 0 2 13 12 9 4 1 0 9 2
21 1 10 9 1 9 1 10 0 11 13 8 10 0 9 1 8 10 0 9 4 2
7 10 9 4 1 15 4 2
8 10 0 9 8 13 10 9 2
18 10 9 1 10 9 4 15 16 0 1 15 16 15 8 4 13 4 2
22 10 9 2 16 12 9 13 2 13 10 0 9 7 10 0 9 13 10 9 8 4 2
27 12 9 4 3 8 4 1 10 9 1 10 9 7 10 9 1 10 1 0 9 13 9 1 10 9 11 2
37 1 9 1 15 13 1 15 9 1 10 9 1 11 13 11 1 15 9 2 2 11 11 11 2 15 9 1 15 13 1 10 9 1 10 11 3 2
7 10 9 13 1 10 9 2
7 10 0 9 4 0 13 2
8 10 9 1 10 9 4 0 2
12 1 10 9 13 7 10 9 7 10 9 8 2
7 3 4 15 9 13 4 2
26 10 0 9 13 3 15 9 4 1 10 9 1 9 11 1 10 9 7 10 9 1 11 1 10 9 2
12 3 13 10 0 9 15 1 15 9 4 4 2
35 1 10 9 1 10 9 4 4 2 16 10 9 15 3 1 11 4 4 10 9 1 10 9 1 11 3 4 4 2 16 12 9 0 4 2
27 10 0 9 13 3 1 12 9 1 9 0 1 15 1 10 11 2 15 16 10 9 1 10 13 9 13 2
12 10 9 13 1 0 2 13 9 1 9 4 2
16 3 4 3 10 2 8 0 9 3 4 1 10 9 1 9 2
37 0 0 9 2 1 3 12 2 13 7 13 1 10 11 13 3 1 12 9 9 10 0 9 4 1 10 9 15 13 1 10 12 7 12 12 9 2
13 9 8 2 3 13 2 13 15 12 9 1 9 2
27 3 1 11 16 3 10 9 7 10 9 3 3 3 13 2 3 3 3 9 11 16 3 10 9 4 4 2
21 1 10 9 13 15 3 0 1 10 9 7 13 15 0 15 0 9 1 10 9 2
16 3 4 3 9 1 9 4 2 15 3 3 3 13 4 4 2
5 10 0 9 3 2
12 15 9 13 1 11 12 1 9 1 15 9 2
5 2 8 8 2 2
28 1 15 9 4 3 1 15 13 10 13 9 8 4 2 13 1 15 0 9 10 9 2 9 7 2 9 2 2
7 9 1 10 9 1 8 2
53 15 13 8 9 1 10 9 10 0 9 1 10 1 11 13 11 2 15 9 1 10 9 1 10 0 9 5 3 13 10 9 15 16 9 1 10 9 4 4 2 5 7 15 9 1 8 0 0 9 1 10 9 2
16 10 0 9 4 10 13 9 3 3 4 1 10 0 0 9 2
21 15 4 0 3 3 0 2 16 10 10 9 0 13 4 2 3 4 15 3 0 2
25 16 9 3 1 9 13 15 0 13 0 3 9 2 16 10 9 1 0 13 1 10 0 9 2 2
25 1 10 9 13 3 3 10 9 3 10 9 0 8 13 7 3 10 9 3 10 9 3 0 4 2
34 15 13 3 15 0 9 10 9 4 1 0 9 10 9 1 13 1 10 0 9 1 15 8 2 3 1 15 0 9 9 4 13 4 2
11 10 9 1 8 4 10 0 13 9 4 2
35 7 15 2 15 9 13 1 10 0 9 1 15 2 8 2 2 13 16 15 15 0 9 3 1 9 7 9 16 1 9 7 9 4 4 2
42 15 13 15 10 0 9 4 8 2 7 15 13 16 11 3 1 10 9 1 11 7 11 4 8 2 9 13 15 3 1 15 9 2 3 16 13 15 3 1 15 9 2
4 6 2 9 2
26 7 3 15 8 1 10 9 15 11 13 4 7 15 10 15 1 15 15 11 10 9 10 9 13 4 2
21 10 9 13 12 9 9 1 10 9 1 12 2 3 11 2 11 2 11 7 11 2
16 10 0 9 2 15 13 15 3 16 15 10 0 9 13 4 2
13 11 13 3 3 3 9 1 10 0 9 1 8 2
38 1 15 13 2 16 8 2 10 9 1 12 13 9 1 15 0 9 2 3 15 8 2 8 2 8 2 8 2 8 2 8 7 8 1 15 13 4 2
28 1 15 3 3 13 9 11 13 3 10 9 16 3 15 1 4 4 2 16 13 15 11 15 3 3 3 3 2
2 9 2
13 8 2 8 2 8 2 3 2 8 2 8 2 2
9 8 2 9 1 10 9 13 0 2
24 2 3 13 10 9 4 1 10 9 15 15 3 1 12 13 7 13 15 3 3 15 9 4 2
15 15 13 1 10 9 1 10 9 9 15 0 0 4 2 2
13 0 13 15 10 9 1 11 2 15 15 0 13 2
17 15 9 1 15 3 1 8 9 13 1 11 13 15 2 0 2 2
16 2 1 15 9 13 15 1 15 9 3 15 3 0 4 2 2
22 8 8 2 11 2 2 8 2 11 2 2 8 2 11 2 7 10 9 8 7 8 2
8 8 13 3 3 10 0 9 2
57 10 9 13 15 9 15 3 5 9 13 3 1 15 0 1 10 0 9 13 1 10 9 5 7 10 9 8 2 9 1 10 9 7 9 1 10 9 2 15 15 15 13 2 13 4 2 16 3 1 0 3 10 9 9 4 13 2
7 10 9 4 3 3 0 2
20 12 9 13 15 3 3 4 7 12 1 15 13 1 9 1 10 9 4 4 2
11 10 9 13 3 1 9 10 13 9 4 2
21 10 9 13 1 10 9 3 7 1 12 4 1 10 13 9 10 13 9 3 4 2
11 1 10 9 1 10 9 13 15 3 8 2
15 3 13 9 4 1 11 2 11 2 11 2 11 7 11 2
11 10 9 4 1 12 9 1 10 9 4 2
7 10 0 9 4 0 9 2
15 3 13 15 15 0 16 0 9 1 10 9 4 1 4 2
28 7 0 13 15 16 15 3 3 10 9 4 4 4 16 3 10 9 16 9 10 9 1 10 9 13 4 4 2
10 15 13 15 1 10 0 9 4 4 2
3 13 15 2
6 1 10 0 9 3 2
14 2 10 9 3 1 10 9 1 11 4 3 3 0 2
11 16 3 3 3 10 9 3 0 0 4 2
12 10 9 4 3 0 15 16 15 3 4 4 2
13 15 10 9 13 4 2 13 10 9 1 8 4 2
18 15 13 15 9 2 3 2 7 15 4 1 15 15 15 16 9 2 2
27 9 1 10 9 1 10 9 2 7 1 9 7 1 9 2 4 3 1 10 0 0 9 1 11 3 4 2
42 16 11 13 4 10 11 3 1 4 2 7 3 3 1 11 4 4 2 13 15 10 13 9 4 1 10 9 2 15 3 13 4 4 10 0 0 0 9 3 1 4 2
18 15 1 10 1 10 9 13 9 4 3 0 1 0 9 8 10 9 2
20 15 1 10 0 9 3 11 1 4 13 4 10 3 0 4 1 10 0 9 2
22 1 10 9 1 9 1 10 11 4 9 3 10 3 12 9 0 0 9 1 3 4 2
17 10 9 13 1 10 0 9 1 13 9 3 1 10 9 13 9 2
8 0 9 13 15 3 3 4 2
18 1 10 9 4 0 9 4 7 3 0 9 13 15 10 15 9 4 2
12 3 13 12 9 2 15 1 12 9 1 3 2
25 16 10 9 13 2 13 15 1 11 7 11 3 1 13 9 1 10 0 9 1 15 9 4 4 2
6 15 9 4 15 4 2
11 2 15 4 10 0 9 1 8 13 9 2
3 15 9 2
13 3 13 3 9 3 2 8 2 13 9 2 2 2
5 11 4 15 9 2
10 2 1 11 13 15 0 7 0 4 2
20 15 4 0 1 15 12 7 13 1 10 9 0 7 1 13 9 4 4 2 2
16 1 15 1 8 13 3 3 3 10 0 0 9 2 1 8 2
14 15 4 10 9 15 15 1 9 13 2 2 3 8 2
20 9 1 15 9 4 1 10 11 4 16 15 1 10 9 16 10 9 1 4 2
27 16 10 0 9 1 10 9 3 3 3 0 4 2 13 8 10 9 1 10 11 1 9 3 1 4 4 2
9 3 4 3 10 9 1 0 8 2
11 2 10 9 13 1 8 3 1 10 9 2
10 10 9 4 4 1 11 16 0 9 2
20 1 10 9 1 10 0 9 13 15 3 15 4 16 16 15 15 12 9 13 2
23 10 9 13 3 3 1 9 13 9 2 3 9 1 11 2 4 15 15 9 3 1 4 2
42 15 4 3 4 1 10 9 1 10 11 2 8 2 1 10 9 2 3 11 13 3 10 0 9 1 10 11 1 4 7 15 1 4 4 15 8 1 10 11 13 4 2
9 10 9 13 10 9 1 9 4 2
22 15 13 15 1 9 11 1 13 4 1 15 9 1 10 11 1 10 9 1 15 9 2
18 10 9 13 15 1 15 9 1 10 9 13 1 10 9 1 10 9 2
25 10 9 4 3 0 10 9 1 4 4 16 13 9 1 0 9 1 0 9 1 9 4 4 4 2
11 7 1 9 4 10 9 1 10 0 9 2
16 8 9 2 15 3 15 12 9 13 1 10 0 9 4 4 2
29 16 15 11 0 9 4 7 15 9 13 2 15 13 15 9 3 3 4 16 15 13 1 10 3 0 9 1 9 2
10 15 0 2 3 13 8 4 1 11 2
38 10 9 2 0 4 1 10 0 9 1 15 9 1 10 9 1 12 2 4 1 10 9 1 9 4 16 15 15 9 13 1 15 13 1 10 0 9 2
6 10 9 13 15 3 2
8 2 9 13 3 1 9 2 2
18 11 2 11 2 13 16 1 10 9 1 15 9 10 9 3 4 4 2
29 15 13 16 10 11 2 10 11 7 15 8 9 4 4 16 1 10 0 9 10 9 3 10 0 9 1 13 4 2
28 10 13 9 13 1 10 9 1 10 9 10 9 1 12 9 1 10 0 9 2 16 15 0 4 16 12 9 2
13 1 10 9 4 3 1 11 10 0 9 8 4 2
25 8 2 0 1 12 1 11 2 13 10 0 12 9 1 11 2 3 15 9 10 3 0 9 13 2
16 11 13 15 9 15 1 10 9 2 16 1 15 9 4 4 2
20 0 13 15 1 11 2 3 15 10 1 10 0 9 4 1 10 11 8 8 2
29 15 13 3 0 2 13 15 9 3 1 11 2 13 9 2 13 3 1 10 9 1 10 9 1 10 11 1 11 2
40 8 13 1 8 3 16 9 2 9 7 9 3 3 13 4 16 4 4 16 10 9 1 9 4 4 4 1 10 15 9 2 15 3 10 0 9 13 4 4 2
18 3 13 3 9 1 10 0 9 1 10 9 11 1 4 3 13 8 2
17 0 13 15 1 0 4 15 9 1 10 13 9 2 11 2 4 2
22 10 9 1 10 9 1 10 0 9 2 8 2 13 16 10 9 11 1 11 4 4 2
8 15 13 3 12 4 4 4 2
14 10 9 11 13 3 1 4 3 11 1 15 9 4 2
13 10 0 9 1 11 8 4 3 3 4 1 11 2
9 15 13 3 1 15 9 9 4 2
26 15 1 10 9 1 10 9 4 10 9 15 4 4 1 8 3 0 0 9 8 10 9 1 10 11 2
25 10 0 9 1 9 2 11 2 1 8 13 8 12 0 3 1 10 11 7 15 0 9 4 4 2
20 15 13 3 3 15 9 3 4 16 10 9 10 0 9 1 10 9 13 4 2
22 1 10 9 1 10 11 4 10 0 9 8 7 8 2 8 1 12 1 12 9 4 2
26 1 10 9 1 3 0 9 13 3 3 10 9 7 10 9 1 13 3 3 3 1 10 9 4 4 2
9 1 8 4 3 0 10 0 9 2
38 1 10 9 1 9 8 13 10 9 1 10 9 1 11 2 15 1 10 9 1 10 0 9 15 0 9 13 4 7 15 3 3 1 10 9 13 4 2
15 2 15 13 0 4 2 16 15 13 4 2 2 13 8 2
22 2 1 15 4 15 0 15 1 9 2 3 16 15 3 1 10 9 3 13 13 4 2
10 15 9 2 6 2 15 4 3 15 2
7 15 4 15 3 0 2 2
25 16 15 9 3 3 4 4 1 1 3 5 16 10 9 1 13 10 9 1 15 8 5 4 0 2
29 15 13 2 15 10 9 3 13 4 2 4 3 10 0 9 1 10 9 1 10 9 2 15 0 1 9 4 4 2
12 13 3 16 11 3 3 1 15 9 4 4 2
10 6 2 3 13 9 1 10 9 0 2
18 9 8 7 8 2 10 0 9 1 10 9 2 9 1 10 0 9 2
21 7 3 1 13 11 9 8 15 15 1 9 7 9 1 15 9 3 7 3 13 2
37 15 13 10 0 9 1 15 12 1 9 13 9 1 10 0 7 0 9 2 3 15 10 15 9 1 10 15 13 4 2 7 15 4 3 4 2 2
10 9 13 15 0 1 0 7 0 9 2
23 7 15 13 15 3 4 16 8 1 15 13 1 10 9 7 9 1 9 15 9 4 4 2
25 10 15 9 4 3 15 10 9 1 10 9 15 15 10 13 9 9 7 9 13 4 16 10 15 2
34 0 0 9 2 1 13 9 2 9 0 1 10 9 7 10 0 9 1 0 9 1 10 9 2 15 1 15 9 1 10 9 4 4 2
23 11 7 11 13 1 15 9 0 3 10 0 0 9 1 1 10 9 0 0 9 7 9 2
15 1 15 9 1 10 11 4 15 4 1 10 0 9 0 2
34 1 10 9 13 2 13 10 9 9 1 3 12 15 9 15 1 9 1 8 7 11 1 11 4 4 2 16 10 9 8 1 13 2 2
20 0 13 15 1 13 9 1 15 8 1 10 11 3 15 10 0 0 0 13 2
7 3 4 3 15 9 4 2
32 15 0 9 15 15 13 8 1 10 0 9 13 4 2 13 9 1 10 0 9 1 10 0 9 1 11 1 10 11 4 4 2
25 3 13 0 15 9 1 8 2 15 3 10 9 13 4 1 10 9 1 10 9 1 11 1 11 2
13 7 1 9 4 15 0 11 1 11 0 1 13 2
14 15 13 16 15 15 9 1 15 9 15 9 4 4 2
32 10 9 13 3 13 9 3 3 16 1 0 9 10 9 4 4 1 15 13 2 3 16 10 9 3 16 2 8 2 4 4 2
28 1 10 9 1 10 0 9 13 10 9 1 10 9 3 4 4 16 15 3 3 3 4 16 12 9 4 4 2
12 15 13 3 15 16 10 0 9 0 9 13 2
9 15 9 4 0 2 3 10 9 2
29 10 0 0 9 13 8 15 0 9 2 15 1 10 0 0 9 4 4 2 1 12 3 1 10 9 3 1 4 2
19 9 2 0 1 15 9 2 13 3 3 3 1 10 0 9 4 4 4 2
29 10 9 1 10 0 9 4 3 1 10 9 1 10 9 1 9 7 9 1 11 4 1 10 9 2 10 9 11 2
8 11 9 4 3 3 15 0 2
50 3 13 1 10 15 9 10 9 1 10 0 9 11 16 10 0 9 15 10 2 9 2 4 4 16 15 4 4 9 1 4 4 2 7 1 10 15 9 10 0 9 16 3 3 15 0 9 4 4 2
13 1 10 1 11 13 9 4 15 9 0 0 4 2
26 16 13 7 13 2 13 11 2 16 15 0 8 2 3 1 8 9 15 9 7 3 15 9 1 15 2
24 7 3 2 11 2 4 15 1 15 1 11 1 9 7 15 13 15 3 3 3 10 9 9 2
40 15 13 15 3 0 15 9 2 7 16 15 3 13 4 16 15 3 12 9 10 11 4 4 7 3 0 3 4 0 10 9 1 4 2 4 15 15 3 4 2
24 15 4 3 3 3 8 4 1 10 9 2 8 2 1 8 2 15 8 15 9 3 3 13 2
13 1 15 13 1 15 9 15 0 8 1 11 0 2
32 8 2 10 9 1 8 15 15 3 15 9 1 15 9 13 2 13 15 3 0 16 11 3 10 0 0 9 1 0 9 4 2
15 1 11 7 11 3 4 10 0 9 3 10 9 3 4 2
10 10 9 4 3 0 4 16 15 13 2
12 10 13 9 13 3 3 15 9 3 3 4 2
17 9 8 16 3 3 0 3 1 4 1 15 15 0 8 4 4 2
13 15 13 3 3 3 16 10 9 1 9 1 4 2
9 10 9 3 4 4 1 10 9 2
18 10 0 9 2 10 9 2 0 9 2 9 1 13 2 9 1 9 2
18 10 0 9 13 3 3 4 2 15 13 4 16 15 15 0 13 4 2
32 1 10 9 2 8 2 4 15 3 1 10 9 4 1 10 0 9 8 7 10 9 4 8 10 9 1 4 1 10 0 9 2
34 15 13 1 15 13 5 10 9 1 1 10 9 9 12 9 2 16 3 15 3 2 5 13 15 4 1 10 9 5 3 15 13 7 2
7 1 15 9 10 9 13 2
29 10 15 9 4 10 0 9 1 10 0 9 2 15 3 15 0 9 13 7 1 10 9 4 4 1 10 0 9 2
21 15 9 13 3 3 1 13 9 7 0 4 3 3 9 3 4 2 1 15 3 2
23 1 10 0 9 13 3 10 0 9 15 3 3 4 2 1 10 9 1 0 9 1 9 2
19 13 0 9 1 10 9 3 2 1 7 3 2 1 10 9 13 15 3 2
36 8 1 11 13 1 10 9 1 9 11 0 9 1 10 9 1 10 11 1 0 9 3 1 4 1 10 9 1 10 9 9 7 9 1 9 2
12 1 11 4 12 1 10 12 9 1 9 4 2
24 3 4 9 4 1 10 9 16 1 0 9 1 4 1 9 1 10 9 1 10 9 1 9 2
2 9 2
16 15 13 10 9 4 1 8 12 2 10 9 13 12 9 4 2
15 15 4 8 2 9 1 10 9 8 2 15 15 13 4 2
22 1 10 0 13 9 2 3 10 9 8 4 1 4 2 13 10 0 9 9 15 0 2
20 1 16 9 10 9 1 9 2 2 9 2 2 15 13 1 9 1 10 9 2
5 15 4 10 9 2
21 10 9 3 15 15 13 2 4 3 10 9 7 10 9 1 10 12 9 0 9 2
26 3 1 8 4 10 9 1 11 4 16 10 9 0 10 0 9 1 10 11 1 11 4 2 4 2 2
44 1 15 13 1 10 9 13 10 12 0 1 9 13 1 12 1 12 9 15 10 0 9 1 10 9 1 0 9 13 4 2 15 9 1 10 1 12 9 7 10 9 13 9 2
18 10 9 4 1 10 9 4 4 7 13 15 4 4 10 9 1 4 2
26 16 9 8 13 3 10 9 8 0 9 4 8 10 2 0 9 2 2 13 1 12 1 10 9 11 2
19 15 13 10 0 7 0 9 1 10 9 1 10 9 1 0 1 15 9 2
38 1 15 9 13 2 1 15 9 2 3 4 4 4 10 9 1 10 9 8 1 11 2 10 9 1 12 9 1 9 7 1 9 2 9 7 10 9 2
48 0 13 8 3 9 4 2 7 0 13 3 16 3 1 12 7 12 10 0 9 1 10 11 4 4 2 3 10 0 9 15 3 0 2 7 3 16 15 15 1 13 2 10 13 9 13 4 2
8 10 9 4 3 8 10 0 2
23 15 9 13 15 13 16 15 3 1 10 0 9 4 4 1 15 15 3 15 1 4 13 2
6 10 9 13 15 9 2
8 3 13 15 3 15 0 9 2
32 9 16 15 2 1 15 10 0 1 15 9 1 15 13 4 1 9 4 4 2 13 15 1 10 9 16 15 3 16 9 13 2
18 10 0 9 2 7 3 4 10 11 3 3 2 15 10 11 13 4 2
16 10 9 2 3 13 16 8 10 9 1 10 11 3 13 4 2
38 0 15 3 10 9 2 10 9 1 8 13 10 0 9 4 2 10 9 13 15 1 9 4 4 2 7 10 11 13 3 15 0 9 4 4 7 4 2
11 15 13 0 3 10 9 1 10 9 4 2
8 9 8 13 10 0 9 11 2
37 1 12 4 1 10 11 10 9 4 1 10 0 9 2 16 15 15 1 10 9 1 11 13 2 9 7 13 9 1 15 9 3 1 10 9 2 2
18 15 13 15 9 1 10 9 2 16 15 1 10 11 10 9 4 4 2
40 3 15 7 3 3 10 9 2 13 15 9 4 2 7 15 4 10 0 0 2 0 9 2 15 1 12 9 10 0 9 13 4 1 10 9 1 10 0 9 2
13 15 0 9 2 2 8 2 2 4 10 13 9 2
10 15 13 1 0 9 3 1 10 15 2
17 3 13 11 15 16 10 0 9 0 15 9 1 10 9 1 4 2
6 7 15 4 15 2 2
13 10 9 13 3 1 10 9 1 10 0 9 4 2
21 3 11 3 13 2 10 9 13 3 1 10 9 1 10 9 1 10 9 1 11 2
17 11 11 13 10 9 4 7 10 9 13 0 4 10 9 1 4 2
48 15 0 4 1 15 9 1 10 11 4 1 15 9 3 0 9 16 9 2 8 10 9 1 10 9 11 2 3 10 9 9 0 4 4 2 16 3 10 9 1 10 9 1 9 0 4 4 2
5 1 11 13 15 2
18 9 13 3 3 9 3 4 2 16 10 9 1 10 11 3 4 4 2
15 10 13 9 13 1 10 0 9 1 13 9 4 4 4 2
32 10 11 2 15 15 3 9 3 13 1 9 1 11 2 13 1 15 9 10 9 1 9 7 9 1 9 16 9 1 11 13 2
27 3 13 10 11 9 11 1 10 3 1 12 1 15 8 13 9 10 9 1 13 9 1 11 3 1 4 2
31 9 11 13 10 11 4 15 2 1 0 9 1 4 16 9 0 4 4 2 16 15 15 9 1 9 3 13 0 13 4 2
42 3 13 10 9 1 10 13 9 15 13 1 10 9 16 9 11 3 3 4 4 4 4 1 4 16 15 9 1 8 4 4 2 16 3 1 13 15 15 0 8 4 2
9 10 9 1 13 1 15 0 13 2
20 11 7 11 13 10 9 8 1 10 9 4 16 15 2 8 2 3 1 13 2
16 15 13 10 9 3 1 10 9 4 1 0 9 1 0 9 2
31 10 9 3 4 10 9 1 10 9 16 10 9 1 11 2 0 9 11 1 10 9 13 2 3 3 1 4 1 10 9 2
27 15 13 1 9 3 16 15 9 1 10 11 1 15 0 9 4 4 7 16 15 9 1 10 11 4 4 2
10 3 4 11 0 1 15 0 9 11 2
14 1 15 9 13 10 0 9 3 3 3 15 9 4 2
16 16 15 15 0 13 2 13 15 3 0 1 10 0 9 3 2
21 8 2 15 15 1 15 11 1 10 0 9 13 4 2 4 3 3 3 1 4 2
17 8 4 15 3 3 4 16 10 9 13 1 10 9 1 12 9 2
36 15 4 15 9 2 7 10 15 9 4 3 0 1 10 9 2 15 0 1 0 9 13 7 16 15 3 0 4 3 1 10 0 9 13 4 2
23 3 16 3 3 9 4 4 1 12 9 2 12 7 12 9 7 16 12 9 10 9 4 2
5 15 4 15 4 2
31 8 2 10 11 2 8 2 8 2 8 2 8 2 8 2 8 2 8 2 8 2 8 2 8 2 8 2 8 7 8 2
10 10 0 9 13 1 10 9 1 11 2
21 15 13 0 2 16 8 2 9 1 10 9 2 8 2 2 3 10 11 4 4 2
26 1 10 11 13 10 9 1 12 9 4 2 3 10 9 13 4 2 15 4 4 1 10 9 1 8 2
20 1 15 11 1 12 9 13 15 15 9 1 10 9 1 9 8 7 9 8 2
19 11 7 11 13 3 3 10 9 1 11 4 2 11 7 11 4 3 3 2
5 3 12 9 15 2
13 10 9 8 13 13 3 1 10 9 1 10 11 2
18 15 13 15 10 9 8 0 3 1 10 9 3 3 10 9 1 4 2
8 10 9 13 1 10 11 4 2
8 7 15 13 15 0 4 4 2
34 10 9 1 10 12 9 13 9 11 13 1 10 9 1 11 4 10 0 9 16 13 9 3 1 4 1 10 0 9 1 10 9 11 2
17 11 7 11 4 1 10 9 0 7 0 3 13 1 11 7 11 2
6 11 0 9 4 4 2
25 10 9 2 12 2 9 1 11 13 15 15 3 3 4 4 7 13 1 10 9 12 9 0 4 2
6 10 9 4 9 0 2
12 3 4 15 9 3 4 1 10 0 0 9 2
19 9 7 15 9 4 0 0 4 7 1 10 9 13 15 3 3 15 3 2
14 10 9 1 15 9 13 3 3 1 10 0 0 9 2
6 10 9 4 3 0 2
9 7 15 13 0 9 3 4 4 2
10 8 13 1 12 7 12 11 1 11 2
15 8 1 8 1 11 7 10 13 9 1 10 11 1 11 2
29 1 10 9 13 9 1 10 9 2 11 2 7 1 10 9 2 8 2 2 15 1 11 3 10 0 9 13 4 2
26 15 13 15 4 4 2 15 10 9 13 4 1 15 13 1 10 0 0 9 1 9 2 9 7 9 2
10 1 15 8 4 3 10 0 9 0 2
24 15 13 1 12 9 3 10 16 12 9 4 2 3 1 12 11 2 11 1 10 0 11 2 2
28 3 13 12 0 4 2 13 15 3 4 2 15 13 15 3 1 10 9 1 2 1 10 9 1 3 4 4 2
6 15 13 15 3 3 2
8 0 13 15 0 1 10 9 2
4 15 4 0 2
15 1 11 13 15 3 1 15 9 2 7 15 4 3 3 2
12 1 11 13 3 3 3 10 0 0 9 4 2
6 15 13 10 9 4 2
5 10 0 0 9 2
11 2 15 13 15 0 0 2 2 13 11 2
48 1 10 9 1 11 4 3 15 1 15 9 1 9 1 4 2 8 3 3 0 7 1 10 9 1 9 2 9 2 9 2 9 7 9 2 9 15 15 3 13 16 3 10 9 16 1 13 2
10 3 13 1 15 9 3 0 9 3 2
27 1 15 0 9 4 15 3 15 0 2 13 0 9 2 9 2 9 7 9 7 13 15 9 3 3 3 2
13 1 15 8 13 1 15 9 2 10 8 13 9 2
12 3 4 10 0 9 1 10 9 15 0 9 2
16 10 9 7 9 1 10 9 4 3 0 7 0 1 9 13 2
30 7 15 15 1 11 2 9 7 9 13 2 13 3 10 0 9 7 10 0 9 1 10 9 1 10 0 9 10 9 2
31 3 13 15 15 0 9 2 13 1 10 9 1 8 1 8 4 8 10 9 1 9 7 9 1 10 0 9 13 4 4 2
45 15 4 3 0 2 3 2 0 9 2 1 15 9 2 15 3 1 9 1 10 9 1 10 9 1 9 4 4 2 4 1 4 1 12 7 12 9 1 1 10 9 0 13 9 2
37 1 15 13 1 3 12 9 11 13 3 0 3 10 9 1 9 2 3 13 10 9 3 3 12 7 12 9 15 4 2 16 3 15 9 3 13 2
14 2 3 13 3 0 16 3 10 9 1 15 9 13 2
13 3 3 4 10 9 1 15 9 3 3 0 3 2
10 10 9 1 15 9 13 0 9 4 2
15 1 11 13 10 9 15 1 1 11 7 11 15 9 13 2
11 11 12 2 11 12 2 11 12 9 9 2
27 3 9 11 7 9 8 2 12 8 2 15 4 4 1 15 13 1 10 9 13 1 10 9 11 10 9 2
11 10 9 13 7 15 0 13 8 10 9 2
49 9 8 13 3 15 9 4 16 10 9 0 9 2 15 0 13 4 4 2 16 10 9 1 9 11 3 3 0 4 4 1 10 9 16 10 11 15 13 2 16 13 16 10 9 11 3 0 13 2
14 13 9 13 1 3 10 9 1 15 8 1 11 13 2
13 1 9 13 9 1 10 9 8 1 10 11 3 2
11 10 9 1 10 11 4 0 1 15 9 2
23 1 11 7 11 13 10 9 0 12 12 9 1 9 4 2 1 11 7 11 0 12 12 2
12 15 13 3 3 3 3 4 16 15 1 4 2
13 15 13 1 9 16 10 9 1 15 9 13 4 2
28 1 10 9 1 15 8 2 11 2 4 12 9 3 3 4 16 1 10 11 7 11 9 1 10 11 13 4 2
26 15 9 3 4 15 4 1 10 9 1 10 9 2 3 10 9 10 9 4 8 10 9 1 10 9 2
12 1 10 9 4 15 12 9 1 10 9 4 2
14 1 10 12 9 1 11 13 3 3 15 0 7 0 2
22 10 13 9 2 7 11 2 13 10 9 9 3 4 1 10 9 1 9 1 10 9 2
39 8 13 10 9 11 16 15 15 1 10 9 4 1 10 9 2 10 9 15 15 9 3 1 10 9 13 1 9 1 13 7 15 10 9 1 10 9 13 2
15 7 16 10 9 10 9 13 2 4 15 0 3 3 13 2
6 0 13 3 9 0 2
31 3 13 9 15 1 10 9 4 16 15 15 1 15 9 13 7 16 15 3 15 15 9 0 13 4 2 4 15 9 0 2
19 3 15 1 3 13 2 4 10 9 2 7 15 4 3 10 0 9 2 2
15 9 11 13 10 9 1 10 0 9 8 1 10 0 9 2
37 15 4 10 0 9 3 4 2 3 13 15 3 1 15 8 2 1 15 9 1 10 9 15 10 9 3 1 10 9 1 10 9 1 8 4 4 2
35 10 9 1 8 1 11 13 8 1 9 4 2 7 15 15 3 0 1 10 9 1 8 2 9 1 10 11 1 15 8 2 1 15 9 2
16 15 13 1 10 9 7 13 15 16 15 15 1 10 9 13 2
17 16 15 9 4 2 13 15 1 10 9 11 10 9 4 1 8 2
11 15 13 0 16 15 1 10 0 9 13 2
16 1 12 4 3 12 9 7 3 13 3 12 1 15 9 3 2
23 15 13 15 0 9 2 7 15 9 1 10 9 10 9 15 3 1 10 9 4 4 2 2
8 11 4 0 1 15 0 9 2
23 10 9 1 11 13 3 0 4 7 1 15 9 13 15 15 10 9 13 9 3 13 4 2
10 10 9 1 10 9 13 10 0 9 2
39 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 9 7 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 3 2
25 11 2 11 7 11 13 3 1 15 9 2 10 9 4 3 0 1 11 2 3 15 4 15 9 2
5 10 9 4 0 2
15 15 13 3 3 1 10 9 1 10 9 1 10 9 4 2
13 1 11 2 11 2 11 2 11 2 11 2 8 2
13 3 4 11 1 10 11 3 8 2 0 3 8 2
5 12 9 1 11 2
21 15 4 3 1 8 2 9 2 9 1 10 9 7 1 10 0 9 2 3 4 2
16 0 3 2 7 0 2 1 10 13 9 15 10 9 13 4 2
29 3 4 10 9 3 15 16 11 3 1 4 2 8 4 1 9 11 4 16 3 1 0 9 10 9 1 13 4 2
16 10 2 9 2 1 11 13 16 10 9 1 10 9 2 7 2
26 7 3 2 1 15 0 9 1 11 1 7 1 10 9 1 0 9 1 1 10 9 13 10 9 3 2
23 1 1 10 0 9 2 16 11 1 9 15 0 0 9 1 10 9 3 1 10 9 13 2
18 10 0 9 1 15 0 9 4 0 10 9 1 12 2 11 0 2 2
12 1 10 9 13 10 13 9 10 0 4 4 2
35 10 0 9 4 15 1 8 12 7 12 9 1 15 3 8 0 0 3 2 1 4 16 15 1 15 0 9 1 15 0 9 3 0 4 2
22 10 9 1 11 13 15 15 1 15 9 2 16 10 9 3 0 1 15 9 4 4 2
22 1 10 0 9 13 10 9 8 3 1 11 1 10 0 9 1 10 9 15 9 8 2
13 9 8 13 1 10 9 15 1 10 9 1 4 2
35 10 9 1 10 9 4 1 15 0 8 1 8 0 4 2 15 1 10 0 9 0 4 4 2 7 10 9 1 10 0 9 4 3 13 2
18 1 10 0 9 13 10 9 3 0 0 4 16 8 3 9 13 4 2
17 2 3 4 0 4 1 10 9 2 15 15 0 1 15 9 13 2
15 8 3 3 0 9 4 3 4 7 11 13 3 10 9 2
13 8 13 1 11 1 10 12 9 1 12 1 11 2
11 10 0 9 13 1 10 0 9 10 9 2
14 10 9 1 11 4 1 10 12 9 1 11 3 0 2
7 11 7 8 4 3 4 2
27 1 15 9 4 12 9 1 10 0 0 9 3 9 3 4 10 9 2 8 2 1 10 11 3 1 4 2
31 12 9 1 10 0 9 2 15 3 10 9 3 10 9 13 4 7 9 1 2 11 2 1 10 9 13 4 2 4 4 2
6 15 4 9 3 4 2
19 8 1 11 13 9 10 9 10 9 4 16 15 1 8 10 9 4 4 2
30 16 9 7 9 13 10 9 4 1 10 0 9 1 12 1 12 9 11 7 10 0 9 3 15 3 10 9 13 4 2
18 15 13 3 2 13 1 15 9 7 13 15 9 1 15 1 10 9 2
15 3 4 15 3 0 3 4 15 1 10 9 3 3 0 2
18 1 11 13 15 9 3 2 10 11 4 10 0 9 2 3 1 15 2
25 16 10 9 13 3 10 9 3 3 10 9 1 15 9 1 10 16 12 9 1 3 12 9 13 2
33 3 13 15 10 9 1 15 9 4 4 7 15 4 3 15 4 2 16 3 3 3 9 13 3 15 8 1 10 9 9 13 2 2
32 2 15 13 4 4 15 10 9 4 3 15 3 3 3 13 16 15 3 3 0 1 9 13 9 1 15 9 0 1 4 2 2
21 1 0 9 4 15 9 3 3 0 15 1 4 16 1 10 0 9 8 1 13 2
33 2 16 15 0 13 3 13 15 1 10 9 4 16 10 9 4 4 1 9 15 15 0 4 16 15 13 1 3 12 0 9 2 2
31 15 13 9 2 8 11 11 2 9 1 10 0 9 1 10 13 7 0 13 0 9 2 11 2 9 1 10 11 1 11 2
21 15 9 5 9 3 8 5 4 3 0 4 2 3 8 10 0 9 1 10 9 2
18 15 13 3 1 10 0 0 9 1 10 9 1 15 9 2 9 2 2
16 2 3 2 13 2 1 11 7 1 11 13 15 15 3 4 2
52 3 9 8 1 11 7 2 0 2 1 11 15 1 0 9 15 9 8 13 4 1 10 9 1 8 7 15 3 0 13 13 1 10 9 8 7 2 1 10 9 3 1 15 10 9 3 1 15 9 1 8 2
23 3 13 15 9 1 10 1 9 11 13 9 16 9 16 15 0 15 1 10 0 9 4 2
24 10 9 13 9 1 15 8 16 9 2 7 15 15 11 3 0 13 2 13 15 3 0 8 2
41 2 10 9 9 2 15 3 3 13 2 4 15 1 10 9 15 10 9 11 1 4 13 16 15 9 0 9 10 9 13 1 10 9 15 10 9 13 1 10 9 2
31 10 0 9 13 4 2 15 9 2 1 4 1 10 9 1 10 11 7 8 12 9 13 15 3 1 0 9 1 10 9 2
10 1 0 9 13 4 9 10 0 9 2
20 7 9 7 9 13 9 0 2 13 15 1 10 9 1 15 13 3 8 4 2
26 10 9 13 10 9 1 9 7 9 15 2 4 2 2 16 10 9 10 9 7 10 0 9 13 4 2
14 10 0 4 2 16 8 3 1 10 9 8 13 4 2
17 3 13 10 9 7 10 9 16 10 9 2 16 10 9 2 8 2
11 15 13 16 15 15 4 3 0 1 4 2
18 15 13 15 3 15 3 7 13 10 9 8 1 10 9 3 3 4 2
11 15 8 13 1 15 0 9 3 3 8 2
14 10 3 0 0 9 13 15 7 0 7 0 3 3 2
12 15 13 15 3 0 4 1 10 0 0 9 2
16 2 10 9 4 0 0 1 10 9 15 13 4 1 10 9 2
5 15 13 3 15 2
29 11 4 10 9 7 3 13 3 2 16 11 13 4 4 1 10 9 2 15 10 9 13 1 10 9 1 15 9 2
28 16 11 3 10 0 9 4 2 4 15 3 0 2 16 10 9 13 4 4 1 9 10 9 1 10 9 13 2
24 10 9 1 10 9 2 15 10 9 1 10 9 13 16 15 9 1 13 4 4 3 0 8 2
24 10 13 9 1 10 11 1 15 8 1 11 13 3 1 3 12 15 9 0 1 15 9 4 2
7 15 13 3 15 16 8 2
42 15 13 3 0 7 3 10 9 11 2 9 1 10 11 2 13 15 10 9 1 10 9 1 10 9 1 13 9 15 13 4 15 15 9 3 1 10 9 4 1 4 2
10 10 9 11 13 3 10 9 0 4 2
24 1 10 0 9 1 10 11 1 8 13 15 1 12 7 12 3 4 1 10 9 2 8 2 2
19 1 15 9 4 10 9 1 10 9 8 1 10 9 1 10 0 9 4 2
23 1 10 9 2 8 2 13 10 11 15 9 10 9 1 10 9 1 9 7 9 1 11 2
12 10 9 10 9 8 13 3 10 0 9 4 2
11 15 9 2 10 9 8 2 13 10 9 2
41 15 3 15 15 13 4 1 10 11 2 13 8 16 10 9 1 10 9 11 4 2 7 16 15 1 9 1 15 9 4 4 16 15 9 1 9 7 11 1 13 2
30 15 4 3 10 11 2 8 1 11 2 3 12 9 13 4 4 2 4 1 9 1 4 1 10 11 2 8 1 11 2
43 2 10 9 4 0 16 0 15 8 1 4 1 10 0 9 2 2 3 8 1 11 1 10 9 1 2 8 2 2 15 15 3 1 10 1 11 13 9 1 15 8 13 2
21 15 13 15 3 2 7 15 13 15 3 4 2 16 15 13 3 10 9 3 4 2
5 10 9 13 9 2
22 15 13 1 10 9 15 9 7 13 1 10 9 3 10 9 15 1 15 13 4 4 2
9 3 13 15 15 1 10 9 3 2
6 10 9 13 15 3 2
14 9 8 4 3 12 9 1 9 2 1 12 3 8 2
35 1 10 1 10 0 12 9 1 12 13 9 9 4 4 12 2 12 2 0 9 2 3 9 2 7 1 10 9 13 9 12 2 12 2 2
36 13 1 9 13 10 9 13 9 1 10 0 12 9 1 12 1 12 2 12 2 9 2 12 2 12 2 2 9 7 12 2 12 2 0 9 2
22 8 10 9 8 4 1 10 9 1 11 15 0 0 8 4 2 15 3 10 9 13 2
9 10 9 8 1 11 4 0 0 2
31 10 0 9 13 11 1 10 0 13 11 1 10 13 0 9 1 8 2 11 2 7 10 15 0 4 11 1 8 2 11 2
25 0 9 8 1 10 9 8 2 15 8 2 4 3 0 13 1 10 9 1 15 8 1 9 4 2
10 6 2 3 13 15 15 9 3 3 2
19 10 0 9 4 1 11 1 8 1 11 15 3 10 0 4 1 15 9 2
30 10 0 0 9 4 1 10 0 9 4 1 9 1 9 3 16 1 9 7 9 3 4 4 1 9 8 1 10 9 2
14 10 0 9 3 13 8 4 4 2 3 12 9 0 2
17 10 9 13 10 9 1 12 9 7 4 9 1 15 8 1 11 2
21 1 15 9 2 9 11 2 4 15 3 0 2 16 3 15 9 13 3 1 4 2
13 10 9 13 8 3 8 4 1 9 15 3 4 2
36 3 13 15 0 9 15 1 10 9 7 16 15 13 15 3 13 1 10 9 4 4 2 3 3 15 9 1 4 1 10 0 9 1 0 9 2
15 3 13 3 15 9 15 3 8 9 3 13 15 1 4 2
12 3 4 10 9 4 16 10 9 15 1 13 2
14 13 13 11 3 10 15 9 1 15 9 9 4 16 2
26 6 2 15 9 4 0 3 0 2 7 15 13 3 10 0 9 1 15 10 9 0 9 3 0 13 2
28 2 13 15 3 10 9 2 2 7 2 11 3 10 9 1 2 7 2 15 13 15 9 1 10 0 9 2 2
13 11 13 15 3 15 3 1 15 9 3 1 4 2
17 15 13 16 15 15 0 4 4 2 10 13 9 4 3 1 4 2
14 15 8 13 1 12 12 9 10 9 4 16 1 12 2
20 3 4 4 1 10 0 9 1 3 2 15 4 4 8 9 1 9 10 9 2
21 15 10 9 13 1 4 10 9 1 10 9 0 1 9 3 1 4 1 10 9 2
14 1 9 4 4 2 16 3 3 10 9 4 4 4 2
13 10 9 1 9 10 9 4 0 1 15 9 4 2
18 10 11 7 10 11 4 1 10 9 1 10 10 9 10 3 0 9 2
25 15 4 4 1 10 9 3 10 9 2 4 3 3 9 15 15 0 13 2 1 12 9 4 4 2
8 7 15 9 13 15 0 0 2
21 1 10 9 13 2 16 12 9 1 15 13 10 11 0 13 7 12 9 10 11 2
11 10 11 13 1 10 0 9 1 12 9 2
31 10 9 1 10 0 11 2 9 11 2 13 3 1 10 9 1 12 9 2 15 1 10 9 8 7 15 1 10 9 11 2
41 10 9 1 10 0 9 8 1 11 2 3 13 2 1 10 9 2 13 15 9 11 1 10 9 2 16 15 1 12 15 9 5 13 1 10 9 5 1 9 13 2
12 1 15 0 9 1 10 11 4 10 9 4 2
44 16 15 15 9 13 2 13 15 3 3 4 16 15 3 1 12 15 12 9 0 4 16 10 9 8 15 9 13 1 15 13 1 10 0 9 15 15 1 15 9 3 13 2 2
18 15 13 3 1 9 11 1 11 10 9 1 10 11 1 15 8 8 2
21 10 11 7 10 11 4 10 0 9 1 15 9 7 3 10 0 9 1 10 11 2
29 15 13 3 3 3 1 4 2 3 16 13 10 15 9 5 15 13 3 15 5 3 10 0 9 1 15 4 2 2
13 13 10 9 1 15 9 8 9 4 1 15 9 2
9 15 13 2 8 2 3 3 0 2
24 2 10 9 1 11 4 1 15 10 9 3 4 16 3 1 4 2 7 15 4 3 0 4 2
13 15 13 12 9 0 1 10 0 9 1 11 4 2
9 15 4 15 3 3 1 15 9 2
37 8 1 11 3 2 10 0 9 1 10 0 9 2 15 3 1 10 3 0 9 13 16 1 10 0 1 9 9 1 12 9 12 9 9 1 13 2
27 2 15 13 15 0 4 1 10 9 2 2 13 2 8 2 2 7 15 13 15 0 16 3 1 4 2 2
24 16 3 13 13 11 1 10 12 9 0 9 1 12 9 15 15 1 9 13 1 8 7 8 2
29 15 8 1 11 4 0 7 3 13 10 9 1 11 10 9 1 9 7 15 9 8 1 9 1 9 3 3 4 2
23 10 11 2 15 1 12 1 10 9 1 9 4 4 2 13 1 12 1 10 0 9 0 2
24 1 10 9 11 4 15 3 10 9 1 10 9 2 10 0 9 2 10 9 7 10 0 9 2
24 10 9 9 1 10 9 2 10 9 9 2 10 9 1 10 9 7 10 0 9 8 1 11 2
14 15 8 1 10 9 13 2 15 13 15 15 16 0 2
10 3 13 15 15 12 9 15 0 13 2
20 0 2 1 10 0 9 2 15 3 8 3 10 0 9 1 9 3 13 4 2
9 10 9 3 15 13 2 13 8 2
8 15 13 1 12 9 10 9 2
8 3 13 10 9 1 12 9 2
21 15 4 10 3 13 9 8 8 1 13 1 10 9 1 12 9 2 12 9 2 2
37 15 13 3 8 2 10 9 1 10 0 9 1 15 8 2 15 1 15 9 1 15 8 15 9 4 4 1 4 16 15 15 9 3 1 10 9 2
14 2 15 13 3 8 1 15 9 2 2 3 13 15 2
24 15 13 3 1 10 9 1 10 9 1 9 1 10 15 9 13 2 3 0 2 13 15 3 2
16 15 13 0 10 9 2 13 8 2 7 13 8 15 1 11 2
11 15 13 10 9 1 11 16 10 9 9 2
10 15 13 3 1 15 9 1 15 9 2
26 3 13 15 15 0 1 10 9 4 2 10 9 13 1 9 3 10 9 2 7 13 3 10 9 9 2
10 15 13 1 15 1 10 9 8 4 2
24 8 2 8 1 10 9 1 11 2 13 1 10 9 1 9 9 4 1 10 9 1 10 11 2
19 15 13 15 1 9 1 10 9 1 12 4 1 10 0 9 1 9 11 2
30 15 13 15 9 1 10 9 2 16 9 9 4 4 2 15 1 15 9 4 4 2 3 15 0 4 4 1 15 9 2
16 1 10 1 10 9 13 9 13 3 12 9 1 10 0 9 2
30 11 13 10 12 12 9 0 9 1 10 11 4 1 9 1 3 2 3 4 1 9 1 10 9 1 8 1 11 4 2
31 9 2 15 1 10 9 13 16 15 9 9 0 4 4 3 0 16 1 1 11 13 9 15 1 4 2 3 10 0 9 2
22 1 15 9 2 15 13 1 9 2 13 15 3 1 12 9 1 13 9 4 4 4 2
9 16 15 3 15 9 0 9 4 2
31 10 0 9 8 4 1 10 9 1 10 9 1 15 9 4 2 16 15 1 12 0 13 4 10 9 1 8 3 1 4 2
20 10 9 2 15 3 3 0 4 4 2 4 1 10 9 1 9 1 10 9 2
21 3 13 3 15 9 4 1 10 9 7 1 10 9 1 10 9 8 9 4 4 2
16 10 11 13 3 10 9 1 15 9 16 10 0 9 1 4 2
11 10 9 1 8 4 4 1 10 9 8 2
34 8 2 9 1 8 9 16 8 2 8 7 8 1 15 9 12 9 1 10 0 9 4 4 2 4 3 10 9 1 11 0 9 8 2
23 15 13 10 9 1 10 9 7 9 16 10 9 3 1 13 1 10 0 9 1 15 9 2
7 15 4 1 10 9 4 2
18 1 10 15 9 1 10 9 13 1 12 9 0 12 9 7 9 3 2
25 10 9 1 10 9 2 8 2 13 1 10 10 0 9 7 15 9 10 9 1 10 9 4 4 2
40 10 9 8 13 12 9 3 8 1 15 4 1 10 9 0 9 2 13 1 10 9 1 11 2 13 16 9 1 15 2 8 2 1 10 9 1 11 1 11 2
5 3 4 9 4 2
6 10 9 4 15 4 2
10 15 13 3 0 3 3 9 3 4 2
6 9 1 8 1 11 2
2 8 2
7 8 7 10 0 9 8 2
19 10 9 2 15 1 8 13 2 4 4 1 10 3 13 9 8 7 8 2
20 10 0 13 10 9 3 16 9 1 15 13 1 8 7 8 1 10 0 11 2
15 15 13 15 9 1 11 7 13 15 11 2 13 1 11 2
16 1 15 9 1 10 13 9 13 8 15 13 1 12 0 9 2
7 15 13 15 9 1 8 2
15 10 9 1 15 8 2 11 2 7 10 9 1 9 11 2
38 15 8 13 1 15 9 16 10 11 15 3 8 4 4 1 2 0 9 3 0 9 10 9 4 4 2 7 15 1 0 9 3 4 1 4 4 2 2
18 1 8 13 10 0 9 3 4 4 16 3 10 9 13 1 0 9 2
9 7 1 10 9 13 8 15 3 2
8 3 3 13 8 15 0 9 2
15 7 16 15 1 15 9 13 2 13 10 9 3 0 3 2
17 7 1 10 9 13 15 5 1 9 2 13 11 0 4 5 8 2
17 15 9 0 13 10 9 1 10 9 7 13 11 3 10 9 3 2
11 8 8 11 2 12 2 1 15 0 9 2
13 2 15 13 15 0 16 11 3 15 9 4 4 2
14 3 4 15 3 3 7 13 15 15 9 1 15 9 2
25 10 9 15 1 10 3 0 13 9 8 10 0 9 1 10 9 13 2 13 15 3 3 1 4 2
10 0 9 13 1 11 10 0 13 9 2
17 10 9 15 8 13 1 15 0 13 13 1 0 9 1 9 8 2
6 11 4 3 1 4 2
29 13 8 3 10 9 4 16 8 10 9 13 2 16 11 10 9 1 15 9 1 10 9 13 4 4 2 12 2 2
16 8 13 3 1 4 1 10 13 9 1 10 9 1 15 9 2
15 2 3 3 10 0 9 4 10 9 1 15 13 0 9 2
17 10 9 2 3 11 1 9 0 1 11 4 4 2 4 0 4 2
14 15 13 0 1 15 9 1 2 2 13 11 1 13 2
27 2 7 16 15 8 7 15 8 4 4 1 10 9 16 10 3 0 0 9 3 1 13 2 13 15 3 2
20 10 9 13 15 12 9 3 1 11 16 1 12 10 9 9 13 1 10 9 2
13 11 13 10 0 9 4 16 15 13 9 1 4 2
45 13 2 13 15 15 7 13 3 3 2 3 13 10 15 0 9 3 8 2 8 2 2 9 1 10 9 9 2 3 0 9 2 3 1 10 0 9 1 10 0 9 3 4 4 2
27 15 13 3 3 10 0 9 1 4 15 10 0 3 1 10 9 1 15 9 1 10 0 13 9 13 4 2
10 16 10 0 9 13 2 13 15 4 2
7 8 2 3 13 15 3 2
6 13 9 4 10 9 2
7 13 15 15 3 3 4 2
6 15 9 1 3 2 2
10 3 13 10 9 15 3 9 1 8 2
17 2 13 15 2 13 9 13 15 3 0 12 9 9 1 10 9 2
14 15 13 4 4 16 10 15 9 15 8 4 1 15 2
16 9 13 10 9 16 15 0 1 10 9 4 7 15 9 4 2
8 15 13 15 4 7 15 15 2
17 15 13 3 0 3 15 3 3 2 7 15 13 15 3 0 2 2
19 1 15 9 10 0 9 10 10 9 13 2 4 3 3 3 0 8 4 2
11 11 4 1 12 1 9 13 9 3 4 2
3 11 3 2
30 7 16 15 1 11 7 10 11 3 3 10 9 0 4 4 3 8 3 10 9 1 10 9 1 11 7 1 11 4 2
11 15 13 3 10 9 12 9 3 4 4 2
17 10 9 13 3 10 9 3 2 15 1 15 10 0 9 13 4 2
18 1 10 0 9 13 9 8 15 1 10 1 10 9 13 11 0 0 2
19 8 13 16 10 9 3 8 1 15 9 1 10 1 15 0 9 4 4 2
32 10 9 1 10 9 13 0 1 10 9 1 13 13 4 2 7 16 15 9 3 3 0 13 13 10 9 1 12 9 4 4 2
14 11 13 1 8 4 4 10 9 1 1 10 9 4 2
9 16 15 13 4 2 4 0 0 2
13 15 0 9 2 2 15 13 9 4 1 10 11 2
3 1 9 2
6 10 9 4 3 0 2
16 13 13 15 10 9 8 1 15 15 1 10 0 0 9 13 2
16 15 13 15 15 0 1 4 1 10 9 15 1 15 8 4 2
13 15 13 3 3 15 16 3 3 3 15 9 4 2
10 3 13 10 9 8 4 1 0 9 2
15 8 2 11 4 10 9 2 16 3 0 9 7 9 13 2
10 10 9 13 3 3 3 3 0 4 2
11 15 9 0 7 10 0 9 10 13 9 2
24 7 3 13 15 3 1 10 0 9 1 15 8 2 1 10 0 0 9 2 1 12 0 9 2
11 10 9 4 0 2 15 4 0 7 0 2
6 15 4 1 15 13 2
15 15 13 1 10 9 1 10 9 1 15 0 9 1 12 2
8 15 9 13 15 3 3 4 2
10 10 9 1 9 1 9 4 15 9 2
16 15 13 15 9 3 3 2 16 10 9 3 3 1 4 4 2
7 1 9 2 1 10 9 2
14 10 9 4 0 16 15 9 10 9 1 10 9 13 2
35 7 3 13 10 9 15 10 0 9 13 3 0 2 0 2 3 16 15 0 9 1 9 0 13 4 2 3 10 9 15 3 0 13 4 2
3 8 3 2
7 7 3 2 9 1 9 2
19 9 4 0 2 15 13 0 2 15 4 3 0 4 7 3 3 0 4 2
16 10 9 7 10 9 1 8 1 10 9 1 11 4 3 4 2
19 10 9 2 3 3 10 9 1 15 9 2 4 1 0 12 12 9 4 2
21 10 9 4 1 12 4 1 10 9 11 2 10 9 1 12 9 1 10 9 8 2
20 10 9 0 13 3 15 3 1 10 9 15 13 4 2 15 4 4 7 4 2
8 9 11 2 4 1 0 9 2
19 15 13 3 0 3 4 12 9 1 10 9 8 1 15 8 1 4 4 2
12 1 15 13 2 13 9 13 15 1 9 4 2
15 15 13 15 0 7 3 13 15 3 3 3 0 16 0 2
11 9 8 13 10 9 1 12 9 1 13 2
25 1 15 9 9 4 10 9 0 4 15 2 13 2 9 1 10 11 1 10 0 9 3 1 4 2
10 1 10 9 13 2 16 15 9 13 2
6 11 7 11 13 3 2
32 15 13 1 15 9 3 1 15 9 1 10 9 3 9 1 0 9 15 3 13 1 15 9 2 11 2 4 4 16 10 9 2
3 8 13 2
40 2 0 13 15 3 3 2 16 3 13 1 10 9 7 13 1 10 9 3 15 9 4 1 15 13 1 10 0 9 7 10 0 4 1 15 0 7 0 9 2
37 10 0 9 13 10 13 9 12 9 4 2 15 13 0 10 0 9 1 11 2 11 2 11 2 11 7 11 1 9 12 9 1 9 1 4 4 2
9 15 9 13 0 12 9 9 4 2
29 10 9 13 10 9 4 2 16 9 10 9 8 4 4 16 15 1 10 9 1 10 0 9 13 9 3 1 4 2
17 15 13 3 1 4 16 15 15 13 3 4 4 1 15 13 3 2
6 15 13 15 1 8 2
17 2 15 0 9 4 1 15 10 9 1 0 9 7 10 0 9 2
11 15 15 0 13 4 10 9 1 10 9 2
14 0 13 10 9 0 9 2 3 16 15 3 13 4 2
15 15 13 15 0 7 0 16 10 9 16 10 2 11 2 2
8 15 4 0 1 15 0 9 2
29 15 8 2 11 2 7 8 13 1 10 0 9 4 16 3 1 10 9 1 15 15 9 4 7 3 3 4 4 2
36 10 9 1 10 12 9 13 15 3 1 10 0 9 1 10 9 2 7 1 10 9 1 15 2 3 9 13 7 1 11 13 9 8 10 11 2
10 9 13 16 10 9 10 9 4 4 2
36 10 0 9 1 10 9 9 1 10 11 13 9 13 15 9 3 4 4 16 10 9 1 9 2 12 2 15 10 9 1 4 4 1 10 9 2
12 3 13 15 10 13 9 3 0 10 9 4 2
20 10 9 2 1 10 9 1 10 9 2 4 1 4 1 8 1 12 1 12 2
16 10 9 4 8 1 10 9 1 9 2 8 2 1 11 4 2
18 10 9 1 15 8 1 11 2 8 2 13 15 12 9 13 9 4 2
14 15 13 16 15 13 1 8 15 1 13 4 1 9 2
17 2 13 1 10 0 9 13 15 15 1 10 9 1 10 9 2 2
18 10 9 1 10 9 7 9 13 1 10 0 13 9 1 9 11 9 2
24 1 10 9 13 10 11 16 10 9 1 13 1 0 9 10 0 9 4 1 10 9 1 9 2
13 10 9 13 15 8 1 9 2 10 9 1 4 2
21 10 11 13 11 1 12 9 1 11 10 0 9 4 1 10 9 1 10 0 9 2
42 1 9 1 10 0 9 1 9 1 10 9 10 9 13 10 9 1 9 1 11 15 9 4 1 15 9 16 1 15 1 9 1 13 7 9 1 13 1 9 7 9 2
21 1 8 9 11 1 1 11 2 13 15 2 13 15 3 1 10 9 10 9 4 2
11 10 0 9 4 1 15 9 10 9 4 2
27 9 11 15 10 9 1 11 13 2 13 0 1 10 9 1 10 1 10 0 0 9 1 9 7 0 9 2
15 10 9 1 10 9 1 9 1 10 11 1 12 9 3 2
20 10 9 1 12 9 2 15 10 0 9 3 0 4 2 13 3 0 1 3 2
14 10 9 13 5 13 10 0 9 5 10 9 8 4 2
16 16 0 4 11 0 1 10 9 1 10 9 12 12 9 4 2
12 1 10 9 4 10 9 1 10 0 9 4 2
11 1 10 0 0 9 13 11 1 10 9 2
29 10 0 9 2 16 9 0 9 4 4 2 4 10 9 16 10 9 1 15 9 3 8 1 3 4 1 8 13 2
16 11 13 10 9 1 8 1 8 7 11 13 12 9 1 12 2
9 1 10 9 13 15 15 12 9 2
24 15 9 4 15 9 1 4 1 10 9 2 16 3 0 4 4 1 10 9 1 9 7 9 2
18 10 9 4 3 13 2 10 9 13 1 10 9 3 16 10 9 4 2
35 1 15 9 13 0 1 10 9 10 9 3 2 16 12 9 13 2 16 15 4 4 4 1 10 9 1 10 9 11 2 10 0 13 9 2
8 10 9 13 15 1 0 9 2
15 10 9 13 0 7 0 0 15 1 10 0 9 1 13 2
10 10 9 4 4 1 10 0 13 9 2
6 1 3 4 15 0 2
19 7 3 13 10 15 9 1 3 15 10 9 13 7 1 10 9 13 4 2
8 15 13 10 9 1 0 9 2
22 9 7 15 9 1 10 9 13 3 3 2 13 10 9 0 7 13 15 10 9 3 2
17 0 13 15 15 15 4 4 16 10 0 9 13 2 13 2 13 2
10 1 10 12 9 4 3 9 11 13 2
19 3 8 13 15 16 1 15 16 0 10 9 3 0 3 13 4 1 4 2
18 10 9 1 10 9 1 10 9 13 1 11 2 11 7 11 0 0 2
11 1 10 9 13 10 9 0 1 10 9 2
21 8 9 1 13 13 10 9 3 1 10 9 1 10 9 7 10 9 1 10 9 2
19 3 10 9 1 10 0 11 13 1 10 9 3 7 13 10 9 0 3 2
16 15 9 13 10 0 9 2 13 1 10 9 1 10 0 9 2
24 10 0 9 4 4 7 0 4 1 10 0 2 9 2 2 3 10 0 7 0 9 4 4 2
38 1 15 9 13 15 10 0 0 9 4 2 15 16 9 13 4 4 1 10 0 0 9 1 15 9 2 3 15 13 4 4 15 15 9 7 9 13 2
11 10 13 9 4 13 7 9 1 10 9 2
17 10 9 1 10 9 13 15 1 15 9 3 9 4 1 15 9 2
14 16 15 10 9 1 9 4 1 13 2 4 3 0 2
13 1 11 13 15 15 4 1 10 12 7 12 9 2
15 3 13 3 10 9 1 8 1 9 7 15 4 0 4 2
25 10 9 13 2 16 1 10 9 10 9 4 4 2 16 10 9 1 10 9 1 10 9 4 4 2
8 10 9 4 3 10 0 9 2
6 7 10 9 4 0 2
21 2 10 9 13 2 2 3 11 2 2 8 10 9 2 16 15 10 9 13 4 2
12 15 9 13 3 1 10 9 3 4 4 2 2
18 13 3 2 16 8 3 1 8 1 9 4 7 3 8 1 11 4 2
14 1 10 9 13 3 3 7 3 10 0 9 4 4 2
27 1 8 4 12 0 9 5 1 9 1 10 0 9 5 4 2 3 0 9 0 1 10 9 13 4 4 2
25 10 9 4 1 4 1 0 9 7 1 12 9 13 10 9 1 8 2 8 7 8 0 9 4 2
24 9 13 1 11 1 10 9 10 0 9 3 0 2 1 10 9 4 8 15 9 3 0 13 2
34 12 1 10 9 13 0 1 0 9 2 12 13 1 10 9 15 8 4 4 7 12 4 1 10 9 4 16 8 10 9 3 1 13 2
11 1 10 11 2 4 15 8 2 9 2 2
19 12 9 1 15 8 7 1 11 2 11 7 8 13 1 8 1 8 4 2
7 10 9 9 13 4 4 2
13 1 10 9 1 8 13 8 9 7 9 1 9 2
21 7 15 15 8 10 9 16 15 8 12 9 3 16 0 10 9 8 1 9 4 2
11 3 13 3 3 12 9 1 15 9 4 2
14 9 11 13 1 12 5 11 0 9 5 10 0 9 2
13 10 9 1 9 2 9 8 12 2 9 8 12 2
8 1 3 0 2 1 3 0 2
10 10 0 13 16 10 0 1 10 9 2
37 10 9 2 1 10 0 9 2 7 3 1 10 0 9 1 10 0 9 1 8 7 10 9 2 15 3 1 10 0 9 4 4 1 10 0 9 2
28 1 10 9 4 3 12 9 0 4 2 7 10 9 13 3 1 12 2 16 10 9 13 10 0 9 1 4 2
22 13 1 10 9 9 13 2 8 2 15 0 13 9 1 15 7 15 0 7 0 9 2
11 0 13 15 9 15 15 1 15 9 0 2
20 7 1 10 9 7 1 10 9 4 3 1 10 9 1 10 9 0 9 4 2
17 1 0 9 13 3 3 10 9 1 4 1 12 15 13 0 9 2
20 9 1 9 13 9 4 4 2 3 16 15 13 1 10 9 3 10 9 13 2
21 15 13 10 9 0 7 11 3 1 10 9 2 16 15 3 1 15 8 13 4 2
23 1 10 9 13 15 9 3 9 4 2 16 15 3 13 1 10 9 3 15 9 4 4 2
16 10 12 9 13 3 16 9 1 0 7 9 15 9 4 4 2
11 1 15 9 4 15 15 9 3 8 4 2
16 10 0 9 1 15 8 1 10 11 1 11 4 8 0 4 2
14 8 2 9 1 10 9 1 8 2 13 10 9 4 2
11 10 9 4 1 10 9 1 15 9 8 2
24 10 9 1 15 8 1 11 4 3 0 4 1 10 9 15 1 9 1 10 0 9 4 4 2
13 15 13 3 2 1 10 0 0 9 10 0 9 2
3 8 13 2
15 2 10 0 3 13 15 9 1 10 0 9 1 10 9 2
8 15 13 15 1 13 1 13 2
13 15 13 15 0 9 1 10 0 0 9 8 4 2
24 15 13 15 9 3 0 1 4 2 16 15 9 13 1 4 1 10 1 10 9 13 9 2 2
15 3 15 13 1 8 13 1 10 0 9 13 9 10 9 2
4 15 9 13 2
17 3 1 15 1 11 2 15 3 3 4 4 1 10 0 13 9 2
19 1 11 13 10 0 9 5 3 0 15 3 13 4 5 0 3 10 9 2
17 10 0 9 4 3 0 0 1 4 2 3 3 3 0 9 13 2
30 15 4 3 4 1 15 13 9 2 3 15 3 15 0 13 7 10 15 0 9 1 10 15 1 15 0 13 9 13 2
11 15 4 10 13 9 0 0 1 10 9 2
25 3 13 16 1 0 9 1 10 9 1 9 1 11 15 0 1 4 4 16 10 9 0 4 4 2
18 9 1 13 9 13 1 9 2 16 10 9 1 10 7 15 9 4 2
17 1 10 9 4 10 9 3 0 0 2 3 10 9 0 15 13 2
17 0 9 1 13 9 13 0 10 9 2 16 10 9 3 0 4 2
13 3 4 1 10 9 2 8 2 3 0 9 4 2
23 0 9 4 3 3 2 16 3 10 9 1 9 3 11 10 0 9 3 4 3 1 4 2
6 7 10 9 13 3 2
30 1 10 9 1 8 4 3 3 10 0 0 9 1 4 2 13 1 10 9 1 15 15 1 15 9 10 9 13 4 2
26 10 0 9 4 3 16 15 9 15 9 1 11 13 2 16 10 9 10 9 4 1 9 7 0 9 2
16 16 15 3 1 13 1 9 4 1 4 2 13 3 10 9 2
4 10 13 9 2
23 10 9 13 16 3 1 13 2 0 0 4 2 15 4 13 2 7 13 15 3 3 0 2
13 3 13 15 13 3 16 9 2 7 15 4 0 2
13 16 1 13 4 15 3 0 2 4 10 9 4 2
10 3 13 15 9 3 16 1 15 13 2
19 1 15 9 3 1 13 4 2 4 15 3 0 1 3 2 7 13 15 2
3 10 9 2
10 9 0 9 13 10 9 1 10 9 2
5 3 13 12 9 2
13 10 0 1 10 12 9 13 9 4 4 1 9 2
15 8 1 12 13 10 9 1 10 9 10 9 3 1 4 2
17 1 15 9 13 15 10 0 9 7 15 9 4 7 10 9 1 2
5 2 13 15 0 2
7 15 13 3 15 0 9 2
9 15 13 10 9 3 3 3 3 2
33 7 16 11 1 11 13 10 9 1 4 2 4 0 0 2 8 10 9 15 1 10 9 1 15 9 3 10 0 9 13 4 4 2
21 15 9 4 3 3 10 9 0 3 1 13 2 3 3 13 16 15 15 9 4 2
14 7 10 9 2 15 15 9 8 8 13 2 13 4 2
7 15 13 1 15 0 2 2
11 3 13 3 1 8 10 9 1 9 3 2
14 10 0 9 4 15 3 0 2 3 1 10 9 3 2
34 13 15 0 9 3 2 3 13 3 9 1 8 8 7 12 9 1 8 1 15 1 4 2 8 16 10 9 1 12 3 1 15 3 2
6 8 2 8 2 11 2
10 3 10 0 9 2 15 3 0 4 2
14 1 10 0 9 4 3 3 10 9 1 10 9 0 2
10 9 8 13 10 9 1 15 13 8 2
9 11 13 3 1 3 3 10 9 2
23 15 13 16 10 9 15 9 4 16 1 4 1 10 9 1 10 13 9 1 10 0 9 2
24 2 10 9 4 0 15 1 4 2 13 15 2 2 7 1 15 9 13 10 9 3 15 3 2
10 15 4 3 9 16 10 9 8 4 2
15 8 1 10 9 2 7 3 13 15 10 9 3 4 2 2
29 10 9 13 10 9 10 9 3 1 4 2 7 10 15 9 3 1 4 15 9 13 4 1 10 9 7 10 9 2
21 3 13 1 10 9 10 0 9 4 1 4 7 10 9 1 10 9 4 1 4 2
19 15 9 3 13 10 9 10 9 3 1 4 8 9 1 9 1 10 9 2
13 0 13 15 1 10 9 3 9 4 4 1 4 2
26 15 9 13 4 4 10 0 9 2 16 1 10 0 9 1 10 9 1 10 0 9 13 4 4 4 2
15 1 15 9 13 15 15 3 1 10 9 1 10 0 9 2
9 15 4 4 1 10 9 1 11 2
13 10 9 8 7 11 4 1 12 1 11 8 4 2
35 15 13 3 10 9 2 16 10 0 9 1 10 9 7 9 2 3 15 3 10 0 9 13 2 10 9 8 10 9 1 15 9 4 4 2
14 1 10 9 13 10 9 1 10 0 9 3 3 8 2
22 9 8 13 1 15 9 1 15 1 10 9 2 10 9 0 1 3 4 1 10 9 2
12 2 10 9 13 13 1 10 9 1 10 9 2
19 10 9 1 15 8 13 1 10 0 0 9 1 9 2 2 3 10 9 2
16 15 13 0 16 1 10 9 10 9 1 10 9 1 4 4 2
21 16 3 3 15 1 4 13 1 11 4 15 3 3 1 15 9 10 9 3 4 2
10 0 13 15 3 0 2 0 13 3 2
11 9 11 13 15 0 2 9 2 1 4 2
27 2 15 4 0 0 1 15 2 2 13 10 9 11 2 16 15 0 4 13 15 0 0 3 4 4 2 2
37 1 10 9 8 2 9 2 7 11 2 9 2 2 13 15 9 3 1 10 0 9 2 2 3 13 15 3 1 9 1 10 9 8 2 11 2 2
20 1 10 9 13 9 11 0 15 9 1 4 16 9 11 0 1 15 9 13 2
46 10 0 9 1 10 0 9 9 13 15 9 5 16 3 1 13 16 3 3 0 9 4 5 12 9 9 4 1 10 9 1 12 9 2 12 7 12 9 2 16 10 9 0 0 0 2
26 15 9 13 10 9 2 15 0 0 15 9 4 2 1 15 15 9 4 7 15 3 10 9 3 4 2
28 15 13 3 3 3 3 2 7 1 10 0 9 1 10 13 9 4 15 0 3 1 4 2 9 3 1 4 2
19 10 0 9 1 10 9 13 15 16 10 9 3 1 10 9 15 4 4 2
18 3 12 15 10 9 1 10 9 2 12 9 2 15 2 16 9 13 2
27 15 7 15 9 4 3 8 4 1 10 9 1 10 9 1 10 11 2 3 3 15 13 1 11 0 4 2
22 8 9 1 10 9 10 9 8 13 3 10 9 8 2 10 9 1 10 9 2 8 2
38 13 9 11 4 3 1 2 8 2 1 11 10 0 9 1 9 4 1 15 9 2 15 16 0 9 13 10 9 1 15 9 1 0 12 9 1 9 2
16 15 4 3 1 10 9 2 15 1 10 9 1 11 13 4 2
34 12 9 4 1 10 9 1 12 1 10 9 1 10 0 9 1 9 1 9 4 1 10 9 2 15 3 1 10 9 8 9 13 4 2
34 1 15 9 13 3 3 10 0 9 4 4 2 7 13 10 9 3 4 3 10 9 1 12 1 10 0 9 1 10 9 11 4 4 2
19 1 10 0 9 1 15 9 13 15 0 10 9 1 10 9 7 10 9 2
34 15 13 15 3 4 2 16 10 9 0 1 9 4 7 16 3 4 10 9 1 10 12 13 9 1 10 9 2 15 0 0 4 4 2
7 15 4 0 10 0 9 2
17 3 13 10 9 15 16 10 0 9 1 10 9 1 10 13 9 2
5 10 9 7 9 2
16 3 4 9 11 3 3 4 16 15 10 0 9 1 11 13 2
38 16 15 1 10 9 1 11 2 3 1 10 9 2 1 10 9 1 12 9 13 4 2 13 10 9 10 0 9 16 3 1 10 9 10 9 4 4 2
9 3 13 0 9 1 10 9 4 2
11 1 15 9 4 9 11 4 1 10 9 2
10 11 7 8 4 12 9 1 10 9 2
6 2 13 8 0 2 2
10 8 15 1 9 7 9 3 13 8 2
22 10 0 9 13 1 0 9 1 10 9 7 13 15 10 9 4 16 10 9 1 13 2
26 8 8 2 15 11 13 4 2 13 11 0 1 10 9 1 10 0 9 2 15 3 3 10 9 13 2
10 2 15 13 15 9 2 2 13 11 2
3 3 8 2
12 2 15 13 10 9 0 1 15 4 4 2 2
43 10 12 9 1 10 0 0 9 2 15 9 2 15 9 10 9 8 7 10 0 9 9 1 10 0 9 11 4 3 1 9 1 9 1 10 0 9 1 10 9 11 4 2
13 1 15 9 13 15 4 1 9 1 10 0 9 2
19 13 1 9 7 9 13 15 1 10 9 1 11 15 9 1 10 9 0 2
16 15 4 10 0 9 11 4 1 15 8 1 11 2 8 2 2
27 8 10 0 9 8 13 12 0 9 5 10 11 2 10 11 7 15 8 5 10 9 1 10 9 4 4 2
15 1 0 7 0 9 4 10 0 9 0 3 10 9 4 2
30 15 9 13 15 8 3 1 12 3 2 3 1 4 10 0 9 1 9 1 0 9 3 1 4 8 10 0 0 9 2
35 10 0 9 1 0 9 1 11 2 8 2 13 4 0 1 4 1 10 9 10 9 3 1 4 3 4 4 3 9 1 10 9 1 4 2
25 1 15 13 10 9 2 9 7 9 2 7 10 9 3 1 4 2 4 15 3 4 1 10 9 2
24 15 13 3 12 9 0 1 4 2 15 1 10 9 1 10 9 1 9 1 10 9 9 13 2
18 10 0 4 2 16 10 9 1 15 9 1 10 9 1 9 4 4 2
15 15 13 3 10 9 3 16 15 1 9 1 9 1 13 2
10 10 9 1 9 13 1 10 9 4 2
28 3 4 3 3 4 16 15 1 15 9 3 4 4 2 6 2 15 4 3 0 3 15 1 9 3 1 4 2
25 1 11 2 12 2 12 7 12 2 7 1 9 2 12 2 12 7 12 2 1 12 7 12 9 2
28 8 4 4 16 15 9 1 9 4 1 0 11 2 15 13 10 9 4 2 3 10 15 9 4 3 3 4 2
16 15 4 3 3 1 10 9 4 3 0 1 10 9 4 4 2
13 15 4 0 0 2 7 10 9 9 13 1 4 2
13 15 13 15 3 2 7 15 13 3 10 9 3 2
22 9 7 9 13 8 10 9 9 2 9 12 7 12 2 3 1 15 9 10 9 4 2
13 15 4 10 9 1 10 9 3 15 3 1 13 2
16 11 13 16 10 9 1 10 9 1 9 7 9 8 3 4 2
22 15 13 0 16 15 10 9 1 10 9 1 10 9 0 4 16 10 9 1 10 9 2
7 10 0 9 9 1 11 2
27 3 13 15 13 3 1 10 9 1 10 9 9 1 4 4 1 10 9 1 15 8 2 15 15 8 13 2
2 6 2
27 10 9 7 3 10 9 2 4 3 0 7 8 8 2 15 3 13 4 16 15 15 4 16 10 0 9 2
8 3 15 3 3 13 1 4 2
28 13 15 3 3 1 8 15 15 3 3 1 9 7 9 9 4 5 0 9 1 9 5 4 1 15 10 9 2
12 15 13 10 13 9 3 7 3 10 9 3 2
15 15 13 9 2 7 15 4 1 10 9 1 11 15 9 2
3 10 9 2
7 15 13 0 1 15 9 2
15 3 3 1 10 9 2 7 1 15 9 3 1 10 9 2
44 15 9 16 15 15 0 13 9 1 10 9 13 2 13 8 1 10 9 1 8 1 11 2 3 15 10 9 1 10 0 11 2 10 9 1 10 12 9 3 13 11 2 13 2
11 3 13 15 10 0 9 1 7 1 9 2
15 10 9 1 10 11 13 3 1 10 0 9 1 9 4 2
5 12 9 15 9 2
9 15 13 1 8 4 16 15 9 2
17 10 9 13 2 16 11 10 9 1 10 9 13 9 3 4 4 2
24 10 0 9 2 1 0 13 9 2 4 1 0 9 0 0 2 13 13 1 10 9 0 9 2
2 11 2
14 2 15 13 15 4 16 15 1 0 9 7 9 13 2
19 1 10 0 9 4 15 3 0 0 1 0 2 10 9 2 1 13 2 2
15 9 1 0 15 9 13 9 15 12 9 1 9 13 4 2
23 15 13 3 10 9 8 7 15 0 9 8 2 15 15 1 15 9 1 8 3 13 4 2
8 15 13 3 3 1 15 9 2
13 10 9 5 8 2 8 5 13 15 15 4 4 2
6 15 4 0 8 4 2
15 4 15 8 0 15 16 1 10 0 9 1 9 1 13 2
26 2 16 15 15 3 4 2 13 15 3 3 2 2 13 11 3 2 2 13 15 3 3 15 8 2 2
23 3 3 13 4 4 16 10 0 9 4 4 1 10 9 3 10 0 9 3 10 9 4 2
25 1 15 9 2 9 7 0 9 13 1 10 13 9 10 0 9 4 4 2 15 0 9 13 4 2
47 3 13 1 10 9 8 8 3 1 15 8 1 10 11 1 10 9 1 10 13 0 9 8 5 10 9 0 1 10 9 1 8 7 11 3 3 10 0 9 1 9 1 10 9 4 4 2
23 10 9 1 2 8 2 4 15 10 9 2 15 15 13 2 15 10 0 9 8 13 4 2
9 3 3 10 13 9 1 15 9 2
18 10 12 0 9 4 0 1 10 13 9 1 10 9 1 10 0 11 2
23 3 1 10 9 2 15 1 10 9 9 1 10 9 1 10 9 4 2 13 10 9 9 2
18 10 0 9 4 10 9 1 15 9 1 10 9 1 15 9 3 3 2
8 15 9 4 1 10 9 4 2
11 10 9 1 9 7 9 4 3 0 0 2
16 9 11 13 3 3 15 9 1 15 13 1 15 9 0 4 2
8 3 13 10 9 1 10 11 2
18 15 13 2 16 15 3 0 4 4 2 16 10 0 9 4 13 4 2
11 3 4 10 9 1 0 9 3 3 0 2
11 13 1 10 0 9 2 13 3 10 9 2
21 3 13 10 0 7 0 9 11 3 3 10 0 9 1 10 0 7 0 9 11 2
2 8 2
8 11 13 0 1 10 0 9 2
19 15 13 0 3 1 10 0 9 1 3 2 7 15 9 4 3 3 4 2
45 15 13 15 3 10 0 9 1 11 4 1 15 13 1 10 0 9 2 15 10 0 9 13 4 4 16 3 1 13 15 9 1 10 9 13 4 1 4 7 3 15 4 1 4 2
39 8 2 15 1 8 7 8 15 1 10 10 9 1 15 9 4 15 0 0 13 4 1 10 9 2 13 1 10 9 3 3 9 4 15 15 9 1 4 2
3 15 13 2
25 2 15 13 15 3 3 4 4 2 15 13 3 1 15 9 2 7 15 13 15 3 3 1 9 2
16 15 13 15 0 0 16 9 2 7 3 10 15 9 1 4 2
20 1 9 1 10 9 7 15 8 4 3 3 10 9 4 3 9 0 3 13 2
26 1 10 9 4 4 2 16 9 3 0 13 1 9 1 9 2 3 9 2 9 7 3 9 4 4 2
6 9 1 15 9 4 2
20 3 3 13 10 0 9 16 10 9 1 9 13 2 16 15 4 4 1 11 2
25 0 1 9 2 0 0 2 3 15 15 13 10 9 7 10 9 2 0 0 1 13 2 0 0 2
17 1 15 13 13 3 0 9 7 12 4 7 0 16 1 9 0 2
8 15 4 3 0 0 1 11 2
14 10 0 9 13 1 9 3 7 13 3 1 10 9 2
8 1 10 15 9 4 15 4 2
7 3 13 12 9 1 8 2
6 2 11 13 3 2 2
15 11 13 15 0 1 10 0 9 15 1 15 9 13 4 2
4 2 8 2 2
4 0 9 3 2
11 3 4 15 15 9 15 3 0 1 4 2
9 3 13 15 0 8 1 13 9 2
26 11 13 1 10 0 9 1 10 9 1 11 1 11 10 9 3 2 15 15 13 15 9 9 1 4 2
36 15 9 4 3 4 1 8 1 11 2 15 1 11 13 4 1 8 2 7 15 15 3 13 4 1 8 2 15 1 10 9 10 0 9 13 2
9 1 11 13 11 3 3 3 4 2
14 15 13 13 1 11 13 1 10 9 9 8 8 4 2
15 7 16 15 13 4 13 0 1 15 13 1 10 9 3 2
10 10 9 1 11 4 15 16 0 9 2
17 0 1 10 9 13 11 2 11 2 8 7 11 15 3 9 3 2
26 15 13 15 4 16 10 9 1 15 3 0 4 4 16 15 1 10 11 1 12 9 1 10 9 13 2
5 15 13 3 4 2
11 15 4 13 1 10 0 9 7 10 9 2
5 2 13 15 3 2
8 3 4 15 9 3 4 2 2
9 3 10 15 9 13 3 3 3 2
20 1 10 11 4 15 3 15 9 7 10 9 15 9 13 4 4 16 10 9 2
18 2 10 9 4 3 2 16 3 0 10 9 13 15 10 0 9 13 2
17 7 15 13 15 15 9 4 1 10 9 1 10 9 1 9 2 2
14 10 0 9 13 10 0 0 9 4 1 9 7 9 2
36 10 9 1 11 1 11 4 10 0 9 2 3 16 4 15 15 3 0 16 3 9 4 1 10 0 9 1 10 13 0 9 1 10 13 9 2
25 15 9 13 3 1 10 9 1 4 1 10 9 15 8 9 0 4 4 1 15 0 13 1 11 2
26 10 0 11 13 8 10 9 8 1 12 1 9 11 1 10 12 9 3 2 10 9 1 10 9 2 2
9 15 15 13 16 3 0 9 13 2
15 15 9 13 3 1 10 9 4 4 1 10 3 0 9 2
30 0 9 13 0 12 9 7 9 10 9 1 10 9 16 4 1 4 1 10 9 1 10 9 7 16 0 9 1 13 2
11 1 10 9 8 1 10 11 13 4 4 2
25 10 9 13 12 9 0 4 7 13 15 11 1 10 12 9 1 12 9 8 1 10 9 1 8 2
25 10 2 0 2 9 1 11 13 1 15 13 1 10 9 1 12 9 3 10 9 1 12 9 4 2
18 15 4 3 1 11 0 4 2 7 1 10 9 1 11 2 15 8 2
9 1 10 9 4 10 9 10 9 2
33 1 10 0 9 1 10 0 1 10 9 4 10 9 10 13 9 3 0 4 2 7 3 3 0 4 16 12 3 10 9 4 4 2
52 16 15 15 9 8 13 1 11 2 15 4 3 3 3 0 1 10 0 9 7 1 10 0 0 9 2 7 0 1 15 8 5 16 10 0 9 1 13 2 13 10 9 1 10 9 15 1 3 13 9 3 2
8 15 13 16 15 15 13 4 2
8 2 1 15 4 15 15 9 2
2 8 2
16 15 9 13 3 3 9 3 4 2 16 11 9 4 4 2 2
17 1 0 9 13 8 2 9 1 11 1 8 2 9 7 10 9 2
28 10 0 9 2 15 1 10 9 15 8 13 2 4 15 1 10 10 9 15 3 7 0 13 4 1 15 9 2
13 15 9 13 15 3 10 0 9 1 10 0 9 2
15 10 9 8 4 1 12 1 12 9 1 10 0 9 4 2
12 1 10 9 13 15 12 9 1 10 9 8 2
2 11 2
34 2 1 10 0 9 7 9 1 11 1 15 9 2 3 15 0 7 0 15 9 13 2 4 15 9 1 10 0 9 0 1 10 9 2
16 10 9 4 1 10 9 1 9 11 16 0 9 4 7 4 2
36 15 15 15 1 10 0 9 1 15 9 13 2 13 3 3 4 16 15 3 8 1 12 9 0 0 4 7 10 9 1 10 9 3 4 4 2
8 2 10 9 13 15 0 3 2
34 15 13 16 8 10 0 9 4 2 16 10 0 9 1 15 1 10 15 0 9 13 4 1 4 16 10 15 9 15 0 1 11 13 2
19 9 11 13 15 0 3 3 15 3 3 7 4 16 9 1 9 12 4 2
12 9 11 13 3 1 10 0 9 15 9 4 2
18 10 9 13 3 12 9 1 12 2 16 16 15 13 1 15 9 13 2
28 16 0 4 10 9 1 10 9 4 1 10 9 1 11 7 10 9 16 10 9 15 9 1 9 4 4 4 2
15 11 9 13 0 3 1 10 3 13 9 1 10 0 9 2
11 15 4 1 4 1 10 0 9 1 8 2
15 15 13 0 16 10 9 3 3 3 3 0 3 1 4 2
33 15 13 4 16 10 9 13 4 7 16 10 9 3 0 4 2 7 15 13 3 4 2 16 15 15 9 0 4 16 15 15 9 2
17 3 11 15 3 10 9 1 10 9 13 1 15 9 1 10 9 2
20 15 13 16 15 13 1 10 9 15 10 9 0 4 7 1 2 0 9 2 2
15 15 3 2 1 15 15 9 7 9 2 13 3 15 3 2
25 16 10 13 0 9 0 9 1 11 13 4 16 9 1 13 2 4 10 9 0 1 10 9 4 2
23 1 10 9 4 10 9 4 10 9 1 4 2 1 15 9 15 15 9 9 8 4 4 2
20 16 3 15 1 9 1 10 9 13 4 4 2 13 15 10 13 9 4 4 2
17 9 3 10 9 5 0 5 4 4 2 13 15 9 0 3 4 2
5 15 4 15 13 2
9 13 4 1 10 9 1 10 9 2
9 15 4 8 10 9 1 10 9 2
7 10 9 13 0 12 9 2
15 12 9 3 4 15 9 3 12 9 13 15 3 3 3 2
36 1 10 9 1 2 8 2 2 10 9 1 15 8 2 4 8 2 0 1 11 2 8 15 0 9 1 10 9 8 0 2 8 0 9 4 2
7 9 11 13 10 9 0 2
8 2 10 0 4 10 9 0 2
10 10 9 1 10 9 9 13 15 9 2
14 9 13 3 1 9 2 7 3 4 15 0 3 1 2
14 15 9 4 1 10 0 9 7 9 3 0 0 4 2
32 15 13 2 16 10 9 1 10 9 1 10 9 0 16 10 9 1 15 2 8 2 4 4 2 7 3 1 9 4 1 4 2
21 1 15 9 13 2 16 10 0 10 9 1 10 9 13 4 16 10 9 1 13 2
15 15 13 9 13 1 10 9 2 3 10 9 10 9 13 2
30 10 0 9 8 4 0 4 1 10 9 13 9 1 9 1 10 9 8 3 1 4 2 16 10 9 0 15 9 13 2
28 8 4 13 11 1 8 1 10 9 4 16 15 1 10 9 8 1 10 9 13 16 10 9 8 0 1 13 2
33 2 3 1 10 9 3 15 15 13 2 11 1 11 2 4 1 9 2 15 15 9 0 3 0 13 2 10 3 0 9 4 2 2
16 10 9 13 3 15 9 7 13 10 0 9 1 15 13 3 2
31 1 10 0 9 4 3 9 4 1 9 2 9 1 9 7 9 2 9 2 0 9 2 9 2 0 9 2 9 7 9 2
38 1 9 1 15 13 1 15 9 2 13 10 9 1 10 11 10 0 0 9 8 4 4 3 15 15 9 7 10 10 15 9 1 10 11 8 4 4 2
19 1 10 9 1 10 9 13 10 9 8 10 9 7 10 0 9 1 8 2
22 15 13 2 15 15 1 15 9 1 10 9 10 13 9 4 7 10 9 1 0 9 2
14 10 0 9 2 1 10 9 1 9 4 3 10 9 2
15 1 0 9 4 9 2 9 7 9 3 15 1 15 13 2
16 3 4 0 9 1 10 13 2 9 2 2 3 10 0 9 2
24 1 15 4 15 0 2 7 9 16 9 1 10 0 9 1 13 16 3 9 3 3 1 13 2
50 10 0 9 2 15 3 15 9 10 9 13 1 10 9 1 12 9 2 15 1 15 9 1 15 8 3 0 4 4 7 0 4 1 3 0 9 2 13 8 15 9 5 15 9 15 9 13 5 4 2
11 9 4 15 15 0 2 13 8 4 4 2
10 1 10 9 4 10 9 12 9 0 2
10 0 9 13 10 0 9 3 3 4 2
15 1 10 9 11 13 10 12 0 9 0 9 1 15 9 2
36 12 9 3 4 10 9 11 1 10 9 4 7 15 13 15 3 1 15 9 8 7 10 0 9 8 1 4 16 15 3 4 7 15 4 4 2
19 10 9 13 11 9 2 9 7 12 9 4 2 7 15 0 9 4 13 2
23 8 13 10 13 9 4 2 7 3 13 15 10 9 4 4 2 3 11 13 9 4 13 2
21 2 15 15 15 15 9 3 0 3 4 2 13 4 2 16 15 15 3 4 4 2
29 1 15 13 15 15 10 9 2 15 15 3 4 4 10 9 1 10 0 7 13 9 1 10 9 3 1 4 2 2
22 3 13 1 10 3 0 9 1 15 9 3 3 1 4 2 16 15 0 0 4 4 2
28 8 1 10 3 0 9 2 15 1 15 9 13 2 8 1 10 0 9 2 15 15 10 13 9 13 4 4 2
14 10 0 9 13 9 0 0 9 7 9 1 10 9 2
30 10 0 13 9 2 15 8 0 1 10 11 13 4 2 7 16 10 9 10 0 9 0 13 4 2 13 0 3 3 2
28 10 9 8 13 15 1 10 9 2 15 11 0 1 15 9 13 7 3 10 9 1 10 9 13 9 4 4 2
33 8 7 8 13 2 1 15 13 1 15 8 1 8 2 10 0 9 3 2 3 9 1 15 8 7 11 0 1 15 9 13 4 2
8 10 13 9 13 15 0 9 2
22 0 9 7 10 3 0 9 13 10 9 1 10 0 9 1 11 1 11 12 9 4 2
14 15 4 3 10 0 9 2 7 15 13 10 0 9 2
40 1 10 9 2 16 3 15 9 3 13 2 13 15 4 4 2 13 1 10 0 9 11 8 11 10 9 0 9 0 16 3 10 0 11 15 1 15 13 4 2
28 1 10 0 9 4 3 1 10 0 9 1 10 9 1 11 1 10 9 1 3 12 9 8 8 10 9 4 2
29 10 9 4 10 0 9 2 15 3 9 13 1 10 9 1 15 9 2 3 15 10 0 9 3 10 9 13 4 2
17 15 9 4 3 0 1 10 9 15 3 10 9 3 3 0 4 2
23 10 0 9 4 15 4 2 16 1 10 9 1 10 9 13 9 7 13 9 2 13 2 2
10 7 15 13 3 15 0 9 1 11 2
10 15 13 2 16 10 9 4 1 12 2
17 15 4 3 3 12 2 7 3 13 15 0 10 0 9 1 15 2
4 10 0 9 2
31 1 10 9 1 0 9 2 15 3 0 13 1 9 1 10 0 9 1 4 5 7 3 15 5 13 15 15 9 9 4 2
17 1 10 9 4 15 0 2 7 15 13 15 9 15 3 15 4 2
19 10 9 2 15 12 9 3 1 9 4 4 2 13 1 10 9 3 3 2
35 1 10 9 10 9 4 3 0 9 7 9 1 10 9 4 2 15 4 13 2 16 15 3 3 13 4 1 10 13 9 1 10 0 9 2
34 3 4 15 1 10 9 12 0 4 10 9 9 1 10 9 1 13 2 16 15 3 0 0 4 2 10 9 1 10 9 15 1 13 2
13 3 13 8 10 9 1 15 9 1 9 3 4 2
8 3 13 3 0 9 1 9 2
26 8 8 2 10 9 15 1 11 7 9 3 10 9 13 4 2 4 10 9 15 0 1 15 8 4 2
20 0 2 16 15 12 9 0 4 16 1 10 9 15 15 1 10 9 4 4 2
21 3 13 11 2 3 1 10 0 9 2 7 9 11 2 10 9 2 0 10 9 2
41 10 0 9 5 0 11 5 13 3 8 9 7 15 4 3 3 11 2 15 1 10 0 9 2 16 10 9 1 10 0 9 1 13 2 13 7 1 10 9 13 2
19 15 4 3 1 11 0 8 4 2 3 9 8 15 13 3 10 9 13 2
19 3 13 11 10 0 0 11 1 10 12 9 7 8 3 1 10 13 9 2
32 16 10 9 1 8 1 10 0 11 15 9 4 13 9 1 10 9 1 11 3 15 1 10 0 9 1 11 15 0 9 13 2
42 10 9 13 3 3 4 2 7 16 10 0 11 10 0 9 3 1 10 9 13 13 9 8 16 15 15 3 3 3 3 1 10 0 9 5 3 12 9 5 4 4 2
21 10 9 4 3 0 7 1 10 0 9 4 15 1 10 9 1 12 9 10 9 2
20 3 9 15 3 13 16 8 7 8 12 13 9 1 9 8 13 4 2 12 2
15 15 13 15 3 1 10 9 4 4 4 15 15 15 13 2
27 10 0 9 1 15 9 4 10 2 9 2 1 10 13 9 7 9 2 3 10 9 15 15 9 13 4 2
28 10 9 4 3 13 1 10 9 1 11 2 7 15 16 10 9 1 8 13 15 9 3 3 2 2 12 2 2
14 1 15 13 1 10 9 1 8 4 15 3 10 9 2
34 16 15 9 2 0 1 10 9 7 9 8 2 1 10 0 9 2 3 13 1 10 9 2 4 10 9 1 15 9 3 3 0 4 2
24 10 0 9 1 15 9 4 3 15 1 10 0 11 7 10 9 10 9 2 8 2 11 2 2
23 10 9 13 1 10 9 1 10 0 9 1 10 0 9 11 2 3 1 10 13 9 11 2
15 1 10 0 9 13 11 3 1 12 0 9 10 0 9 2
26 1 10 0 9 3 13 10 9 1 15 0 9 0 3 2 7 3 13 11 1 12 1 10 0 9 2
27 8 13 8 0 7 13 3 1 10 0 9 1 11 1 8 2 10 9 15 3 1 15 0 9 4 4 2
9 1 8 4 10 13 9 0 4 2
32 12 9 3 13 15 10 0 9 1 2 8 2 2 7 16 15 1 15 0 9 3 3 4 1 4 13 15 0 4 7 4 2
24 0 7 0 9 2 13 11 2 7 10 9 2 7 15 0 9 2 1 10 9 1 10 9 2
26 3 3 10 9 1 15 8 1 8 7 11 16 8 9 4 4 4 10 9 1 0 9 3 0 4 2
14 1 10 11 4 3 9 3 15 0 9 3 1 4 2
23 2 15 4 1 10 9 0 1 9 1 11 7 3 8 11 13 15 15 15 1 4 2 2
21 3 4 11 3 1 11 4 7 10 9 13 9 1 10 9 1 8 2 12 2 2
15 10 11 9 1 9 2 12 2 13 12 9 3 1 8 2
43 15 4 3 10 0 9 1 11 2 10 9 1 10 9 2 10 9 1 11 16 10 9 1 10 9 3 4 13 4 7 10 0 9 2 8 2 2 3 13 1 10 9 2
2 9 2
20 8 2 15 4 13 15 9 1 10 9 8 1 4 2 8 15 0 9 2 2
7 15 4 3 9 7 9 2
9 13 7 13 0 9 1 15 9 2
24 11 13 9 7 0 0 9 2 1 10 9 2 1 9 16 16 10 9 3 10 9 3 4 2
20 9 1 9 2 9 2 9 7 0 9 2 15 9 3 3 13 1 15 9 2
30 15 0 9 4 15 1 10 0 9 1 15 9 2 13 9 12 9 2 1 15 13 9 2 1 15 15 15 3 13 2
30 1 11 2 2 8 2 2 0 8 4 12 7 13 3 0 9 2 16 15 13 1 10 0 9 8 2 3 12 2 2
38 10 9 13 10 9 10 9 4 4 16 1 10 9 1 11 1 10 9 1 13 1 10 9 1 10 9 15 11 1 10 0 9 1 15 12 9 13 2
24 10 9 1 10 9 3 10 9 1 10 9 13 4 2 13 1 10 9 1 0 9 4 4 2
30 1 9 12 1 10 9 13 10 9 1 15 13 1 10 9 4 4 1 9 1 10 9 2 15 3 1 13 9 13 2
24 8 13 16 10 0 9 1 10 0 9 3 0 4 2 7 16 15 1 0 9 0 0 4 2
14 10 0 9 13 1 15 9 10 15 0 9 1 4 2
40 1 8 12 9 4 10 9 4 2 1 15 15 13 4 4 1 10 0 0 9 2 15 13 4 10 9 1 9 1 4 2 7 0 1 10 0 9 13 4 2
15 3 13 1 10 9 9 4 4 3 1 10 0 9 9 2
39 15 9 4 9 1 1 10 9 7 8 13 15 15 9 1 0 9 7 3 0 2 16 10 9 3 3 1 4 13 2 3 10 9 3 1 10 9 13 2
17 3 13 15 8 3 9 3 4 4 13 9 1 10 9 1 11 2
7 10 9 4 10 0 9 2
9 7 15 13 3 3 9 4 4 2
9 10 9 13 4 3 8 15 9 2
26 1 15 10 9 1 15 8 13 10 9 4 4 4 15 15 0 9 1 0 9 1 10 9 4 4 2
25 15 13 3 3 1 9 1 4 16 1 13 16 15 9 1 9 10 9 1 10 9 3 8 4 2
14 15 9 13 3 0 8 4 1 10 0 2 13 9 2
13 7 3 4 15 15 9 3 3 3 9 1 4 2
21 10 13 9 4 3 1 10 0 7 0 9 1 11 11 4 2 8 1 13 9 2
55 8 7 11 4 3 3 3 3 9 15 3 3 13 2 7 10 9 1 11 1 10 9 11 2 11 11 1 10 0 9 11 2 1 9 11 1 10 3 0 9 11 7 1 10 0 11 1 10 15 13 11 13 0 9 2
23 10 0 9 1 10 9 9 2 15 1 11 1 8 4 4 2 4 3 0 16 4 4 2
35 0 13 15 10 9 15 3 3 1 4 2 16 10 9 1 8 3 3 3 4 2 16 15 15 8 1 15 9 3 3 8 13 4 4 2
3 3 8 2
14 3 3 13 10 9 1 10 0 9 3 15 1 4 2
24 10 9 1 10 0 9 13 3 0 9 1 4 2 7 10 9 1 10 9 4 3 3 0 2
13 8 4 1 8 3 8 0 16 10 9 1 3 2
6 11 4 0 1 8 2
10 11 13 8 4 1 10 9 1 8 2
29 3 13 10 1 15 12 9 13 9 3 1 10 9 1 10 9 3 15 9 4 4 2 3 1 9 1 15 9 2
48 15 9 2 15 12 9 0 4 4 3 4 4 2 13 16 10 9 15 3 0 4 16 10 13 9 15 0 4 1 15 13 1 10 0 9 1 9 2 8 7 3 0 0 4 1 4 4 2
15 10 0 9 4 16 15 9 1 10 3 0 9 13 4 2
12 15 4 1 4 1 10 9 1 9 1 9 2
33 9 7 9 1 11 13 10 9 4 1 0 9 1 10 9 1 10 9 1 10 9 15 3 10 0 9 1 10 0 9 0 13 2
20 1 10 0 2 0 9 2 1 10 9 4 0 12 9 1 13 9 13 4 2
15 8 4 10 9 1 10 9 15 3 13 4 4 2 4 2
17 10 9 1 11 2 3 10 9 9 13 4 4 2 13 3 3 2
31 15 13 15 3 16 8 10 0 9 7 10 0 9 1 9 4 4 2 7 10 11 4 4 2 1 15 1 15 9 3 2
24 0 13 15 1 10 9 2 15 1 10 9 4 4 2 10 9 1 0 7 0 9 1 4 2
31 15 9 13 15 1 10 13 9 1 9 1 10 11 2 16 15 1 15 13 1 9 1 10 9 1 10 9 13 4 4 2
24 3 13 15 10 9 11 3 2 15 0 1 10 9 3 13 4 4 15 1 10 9 1 4 2
24 15 13 10 9 10 9 2 3 15 15 13 16 15 1 4 4 4 1 10 9 1 10 9 2
11 11 13 3 3 3 0 10 9 4 4 2
31 15 9 3 4 10 9 1 10 9 1 10 9 1 10 0 9 1 11 15 16 12 9 1 9 13 16 1 11 1 4 2
28 15 13 3 9 4 1 9 2 9 1 9 7 9 1 9 2 2 3 1 15 9 10 0 9 4 13 4 2
14 3 13 10 9 13 1 3 10 0 9 0 9 13 2
35 10 3 13 9 13 10 0 12 9 10 9 4 16 0 3 1 13 1 15 15 9 1 10 8 12 9 15 1 15 9 7 9 4 4 2
30 10 0 9 1 10 9 13 8 1 11 15 15 1 15 9 3 0 4 7 13 16 15 10 0 9 9 3 4 4 2
15 3 12 9 1 15 13 13 15 1 10 0 9 4 4 2
5 9 1 10 9 2
12 2 1 0 9 4 1 11 3 3 9 2 2
27 0 9 13 3 10 10 9 1 11 2 3 1 10 9 1 10 0 9 15 9 4 4 1 10 0 9 2
15 12 9 1 10 0 9 13 3 1 10 9 1 4 4 2
7 3 11 4 0 15 0 2
7 10 9 13 8 0 4 2
9 3 13 12 9 3 1 10 9 2
22 10 9 3 15 15 4 4 7 3 8 10 9 15 10 9 13 1 10 15 4 0 2
18 9 8 13 15 0 4 10 9 1 10 9 1 0 0 9 1 4 2
24 3 13 15 10 0 9 4 2 3 0 1 10 0 7 13 15 10 9 15 4 1 0 9 2
8 10 9 1 10 9 4 0 2
29 8 1 11 13 10 9 10 1 10 9 1 0 9 13 9 1 10 0 9 3 1 9 1 10 0 9 1 4 2
12 2 10 9 13 10 0 0 9 1 10 9 2
33 15 13 1 10 0 9 3 2 16 15 13 13 4 2 16 10 9 1 10 0 9 10 0 9 1 10 9 4 2 2 13 15 2
15 15 13 0 9 13 1 12 9 1 10 0 9 15 9 2
43 9 16 11 2 11 2 15 12 1 8 1 11 13 2 7 11 2 11 2 13 1 9 13 1 10 13 9 2 7 1 10 9 13 3 8 2 11 7 11 2 0 9 2
16 11 7 11 2 13 1 10 0 9 2 13 3 15 9 3 2
6 10 0 9 13 15 2
4 11 13 0 2
18 10 0 9 13 15 3 3 3 0 1 3 16 10 9 0 4 4 2
31 11 13 11 3 1 4 2 3 15 9 1 11 15 9 8 9 13 9 12 9 1 15 9 1 11 13 4 2 15 8 2
37 13 9 4 1 10 0 9 7 9 1 10 9 2 10 9 1 11 4 2 2 10 0 9 2 2 16 10 0 9 8 15 2 9 11 2 13 2
22 0 1 15 9 7 9 13 3 10 9 1 9 2 13 1 10 9 1 11 16 9 2
11 2 15 13 15 3 4 1 15 0 9 2
20 15 13 10 0 9 1 10 9 15 15 16 10 0 0 9 1 10 11 2 2
18 15 13 15 0 16 10 9 4 4 7 1 10 0 15 9 4 4 2
37 1 10 9 1 11 7 11 7 10 0 9 13 3 0 9 9 1 10 9 1 12 9 2 3 1 10 9 1 3 10 9 10 0 9 4 4 2
26 1 0 9 13 10 9 10 9 4 4 2 3 10 9 3 13 4 2 16 10 9 15 0 13 4 2
44 10 9 1 10 0 9 1 9 2 11 2 8 2 13 3 1 15 9 1 10 0 9 1 10 11 1 11 2 16 10 9 1 10 9 1 15 15 9 10 0 9 4 4 2
26 10 0 9 1 9 1 9 7 9 4 0 0 3 7 1 9 13 3 3 3 0 16 12 9 3 2
14 8 13 0 16 11 3 3 4 1 10 9 1 9 2
15 2 3 10 9 16 15 9 10 0 9 4 2 4 0 2
19 10 9 1 10 9 4 0 1 15 1 10 11 7 15 9 13 15 9 2
10 10 9 13 3 9 4 1 15 9 2
18 10 9 1 10 0 9 1 10 9 4 3 3 1 15 9 3 4 2
10 15 4 1 10 11 10 0 9 2 2
20 1 10 9 1 9 8 2 9 2 13 3 10 9 8 2 0 2 1 4 2
10 15 4 1 0 9 1 15 9 4 2
9 15 13 3 0 9 1 15 9 2
4 15 13 0 2
9 15 4 3 1 3 0 3 4 2
9 15 13 0 1 16 15 3 4 2
7 15 4 3 1 9 11 2
10 13 15 1 10 9 1 15 16 15 2
12 15 2 1 2 3 3 2 13 15 1 4 2
5 12 4 10 9 2
13 11 2 13 15 3 9 7 9 2 11 2 11 2
5 0 9 13 3 2
6 15 13 1 10 9 2
7 9 8 13 1 10 9 2
10 9 8 7 9 8 13 1 10 9 2
8 9 8 13 0 1 10 9 2
10 9 8 13 0 9 3 1 10 9 2
8 9 8 13 1 10 9 4 2
8 9 8 13 1 10 9 4 2
9 9 8 13 1 10 9 4 4 2
11 9 8 13 0 1 10 9 4 4 4 2
11 10 9 13 1 10 9 3 1 10 9 2
9 10 9 13 9 1 10 9 11 2
4 10 9 13 2
6 10 9 13 1 9 2
9 11 13 10 0 9 3 4 4 2
10 15 13 3 3 15 9 1 4 4 2
7 11 13 10 0 9 4 2
6 11 13 10 0 9 2
6 11 4 1 9 4 2
4 11 4 3 2
6 11 13 10 9 4 2
6 11 13 1 10 9 2
4 11 4 9 2
8 11 13 3 3 9 4 4 2
4 11 4 9 2
5 11 13 9 4 2
5 11 4 9 4 2
7 15 9 4 15 0 9 2
8 11 13 0 4 4 4 4 2
7 15 4 15 10 9 0 2
9 15 13 15 0 15 1 13 4 2
11 10 9 13 1 10 0 9 1 10 9 2
8 15 9 13 0 1 10 9 2
8 10 0 9 13 3 3 9 2
5 15 4 3 13 2
6 15 4 3 0 4 2
6 15 4 3 0 0 2
9 10 9 4 3 1 3 15 0 2
9 15 4 11 7 15 4 3 0 2
6 15 4 10 0 9 2
8 15 4 10 0 9 1 4 2
5 11 13 10 9 2
6 11 13 10 9 4 2
6 11 13 10 9 4 2
8 15 9 4 3 1 15 4 2
9 15 9 13 3 1 15 4 4 2
9 11 13 15 9 0 4 4 4 2
15 2 15 13 15 9 4 2 16 10 0 9 1 13 4 2
9 15 13 3 15 9 1 4 4 2
6 15 13 15 9 0 2
7 6 2 9 2 15 13 2
5 15 13 10 9 2
7 15 13 3 1 10 9 2
5 9 13 10 9 2
6 9 13 3 1 9 2
5 15 13 10 9 2
7 15 13 3 9 3 3 2
6 13 15 15 8 4 2
5 13 15 3 4 2
6 15 13 15 9 4 2
7 15 13 3 1 4 4 2
5 15 13 10 9 2
4 15 13 0 2
6 15 13 15 9 8 2
5 15 9 13 8 2
8 15 13 10 9 1 10 9 2
7 10 9 13 1 10 9 2
6 15 13 15 9 4 2
4 10 9 13 2
8 6 2 15 13 15 3 3 2
10 10 0 9 13 10 9 1 10 0 2
4 15 9 13 2
5 15 13 10 9 2
4 10 9 13 2
6 10 9 13 10 9 2
6 10 9 13 3 15 2
5 15 13 10 9 2
5 10 9 13 0 2
5 15 13 10 9 2
4 10 9 13 2
8 15 0 9 13 15 1 9 2
6 15 0 9 13 9 2
6 13 15 9 3 0 2
7 9 13 8 0 16 9 2
7 15 0 9 13 3 3 2
8 15 9 13 3 12 9 4 2
9 13 15 15 9 3 15 9 4 2
5 15 13 15 0 2
6 15 13 15 9 0 2
6 15 13 15 9 0 2
8 15 13 10 9 1 15 9 2
10 11 13 1 9 10 9 1 10 9 2
9 15 13 15 9 1 15 9 4 2
4 15 9 9 2
12 15 13 2 15 13 3 4 2 15 0 9 2
7 15 13 10 0 9 4 2
6 15 4 10 9 4 2
6 15 13 15 10 9 2
6 13 15 10 9 4 2
7 15 13 3 10 9 4 2
9 15 13 10 9 1 0 12 9 2
13 2 15 13 3 3 3 1 4 2 2 13 15 2
8 15 13 10 0 9 7 13 2
6 10 9 13 10 9 2
13 2 13 3 3 2 6 9 2 2 13 10 9 2
13 2 15 13 15 3 3 4 2 2 13 11 3 2
8 15 4 3 3 1 15 4 2
10 3 4 1 15 9 3 15 9 4 2
5 10 9 13 0 2
6 10 9 13 3 0 2
10 9 16 10 9 13 11 1 10 9 2
9 15 13 3 3 9 1 15 9 2
4 15 13 15 2
5 0 9 13 0 2
6 13 13 0 16 9 2
5 15 9 13 0 2
6 15 9 13 3 0 2
7 15 13 3 15 9 0 2
9 15 13 15 3 15 1 15 9 2
7 15 13 15 1 15 9 2
7 15 13 15 1 15 9 2
6 15 9 13 15 3 2
7 11 13 15 1 10 9 2
7 11 13 15 1 10 9 2
8 10 9 13 15 1 10 9 2
8 10 9 13 15 1 10 9 2
4 11 13 15 2
7 11 13 15 9 1 9 2
4 11 13 15 2
5 10 9 13 15 2
9 10 9 13 10 9 1 10 9 2
5 10 9 13 15 2
7 15 13 15 1 10 9 2
10 10 9 13 15 9 1 10 0 9 2
9 10 9 13 15 1 0 9 3 2
10 10 9 13 10 9 1 0 9 4 2
11 15 13 15 3 3 0 16 15 3 4 2
8 15 9 13 15 3 0 4 2
11 15 13 15 3 3 0 16 15 3 4 2
7 15 13 15 1 10 9 2
4 11 13 15 2
7 15 13 15 3 16 9 2
9 15 13 15 3 1 10 9 4 2
9 15 13 15 3 1 10 9 4 2
7 15 13 15 15 3 4 2
7 15 13 15 15 3 4 2
4 11 13 15 2
4 11 13 15 2
4 11 13 15 2
5 11 13 10 9 2
9 15 13 15 3 16 9 0 4 2
7 15 13 10 0 9 4 2
8 15 9 13 15 15 0 4 2
6 15 13 10 9 4 2
12 15 13 15 3 1 10 0 9 1 10 9 2
6 15 9 13 15 4 2
9 15 13 15 3 1 10 9 3 2
8 15 4 3 4 1 10 9 2
12 16 10 9 15 13 2 13 15 3 3 4 2
7 10 9 13 10 9 3 2
11 1 15 9 13 15 15 3 10 9 4 2
7 3 13 15 15 9 4 2
9 15 13 15 3 4 1 15 9 2
6 13 15 15 3 4 2
4 15 9 3 2
5 15 9 9 0 2
5 15 13 3 0 2
8 15 13 15 0 1 15 9 2
14 15 13 0 16 15 1 15 9 3 3 0 9 13 2
7 15 13 0 1 15 9 2
6 15 13 0 1 9 2
3 15 9 2
4 15 9 13 2
4 15 9 13 2
4 15 13 0 2
7 10 9 13 1 10 9 2
14 15 13 3 3 4 2 15 13 3 0 1 15 12 2
18 15 9 4 3 0 16 1 13 2 7 1 15 12 13 15 3 0 2
5 15 13 1 9 2
6 10 9 1 9 13 2
8 15 9 3 3 2 15 0 2
7 10 9 13 1 10 9 2
6 15 13 3 3 0 2
7 15 9 13 1 10 9 2
6 15 9 1 9 11 2
15 10 9 13 8 2 1 0 9 13 2 4 1 10 9 2
6 15 13 15 9 0 2
8 9 4 15 3 3 3 0 2
10 15 0 9 13 0 3 10 0 9 2
7 13 11 1 10 9 3 2
10 13 10 9 3 3 4 1 9 12 2
15 16 10 9 3 3 13 4 2 3 13 15 10 9 4 2
11 9 13 0 3 15 9 16 3 1 4 2
4 13 10 9 2
4 0 15 13 2
5 15 13 15 0 2
5 10 9 13 15 2
4 11 0 15 2
4 15 4 3 2
5 15 13 1 4 2
4 11 3 3 2
4 13 3 3 2
5 4 3 3 0 2
3 13 12 2
6 13 15 3 3 4 2
7 4 7 0 1 9 4 2
3 13 3 2
4 0 3 3 2
10 3 13 13 15 3 15 0 9 4 2
5 15 4 11 0 2
5 3 13 13 15 2
5 15 13 10 9 2
3 10 13 9
5 15 13 10 9 2
3 10 13 9
5 9 0 1 4 2
3 8 12 2
6 15 13 3 1 9 2
6 13 15 7 13 15 2
6 13 15 10 9 3 2
5 13 15 2 9 2
5 13 15 2 9 2
5 15 4 3 4 2
8 7 3 4 15 0 3 4 2
11 15 4 10 9 4 10 9 0 1 13 2
6 10 9 4 3 4 2
7 11 4 4 1 15 9 2
9 3 4 15 3 15 15 9 4 2
7 4 15 9 3 3 4 2
10 15 9 13 3 0 9 3 3 4 2
7 10 9 4 15 0 4 2
8 15 0 9 13 15 3 4 2
8 15 4 3 3 10 9 4 2
5 10 9 4 4 2
6 10 9 4 0 4 2
8 15 4 15 3 3 0 4 2
6 10 9 4 0 4 2
8 1 10 9 4 15 3 4 2
5 4 15 3 4 2
10 9 12 13 10 11 0 4 1 4 2
7 15 4 3 4 1 13 2
12 15 4 4 15 3 3 10 9 0 3 13 2
8 15 4 3 3 15 0 4 2
10 15 4 4 16 15 3 0 3 13 2
7 15 13 15 9 0 4 2
7 15 4 8 4 8 9 2
13 3 0 15 9 13 15 3 0 1 10 9 4 2
5 15 13 3 4 2
7 10 9 13 12 9 4 2
6 15 13 10 9 4 2
8 15 13 10 9 1 9 4 2
5 15 13 0 4 2
6 15 13 13 9 4 2
6 15 13 0 0 4 2
16 15 13 3 9 15 9 10 4 2 7 0 13 15 3 4 2
8 15 13 15 3 0 3 4 2
7 15 13 15 3 4 4 2
7 15 4 1 0 9 4 2
6 15 4 10 9 4 2
6 15 9 4 0 4 2
8 15 9 4 15 10 9 4 2
7 15 4 10 15 9 4 2
6 15 4 15 9 4 2
7 10 9 4 10 9 4 2
7 15 4 15 3 3 4 2
8 10 9 4 0 10 9 4 2
10 15 4 15 13 3 3 4 1 4 2
6 15 13 15 3 4 2
5 15 4 3 4 2
6 10 9 13 15 4 2
4 15 4 4 2
7 3 13 15 10 9 4 2
6 10 9 4 3 4 2
6 10 9 13 15 4 2
6 15 4 1 11 4 2
6 15 13 10 9 4 2
5 10 9 4 4 2
7 15 13 15 9 4 4 2
6 15 4 3 0 4 2
8 3 0 13 15 3 3 4 2
8 15 4 1 11 1 11 4 2
10 15 4 1 10 9 1 10 9 4 2
12 10 9 4 3 10 9 4 7 3 0 4 2
7 15 4 10 9 3 4 2
7 15 13 1 10 9 4 2
9 10 9 13 8 3 1 11 4 2
16 15 13 3 3 12 9 4 7 4 2 1 15 3 4 4 2
6 4 15 3 0 4 2
11 15 4 3 0 0 4 1 10 0 9 2
13 4 15 9 3 3 1 10 9 1 15 9 4 2
9 10 9 4 3 10 9 0 4 2
9 10 9 4 4 2 15 13 1 9
10 15 9 13 3 10 0 9 3 4 2
6 15 4 15 9 4 2
11 15 13 3 3 15 9 1 10 9 4 2
13 15 13 3 3 4 15 9 1 15 9 1 4 2
13 15 13 3 3 15 9 1 15 9 4 1 4 2
10 15 4 10 9 1 15 0 0 4 2
18 11 2 3 13 15 15 9 4 2 11 2 1 10 9 1 15 13 2
17 15 13 15 3 4 3 13 15 4 2 7 15 4 15 9 4 2
10 1 15 15 9 4 15 15 8 4 2
10 16 15 15 0 4 15 15 3 4 2
11 15 4 15 1 10 9 1 15 9 4 2
8 10 9 13 15 9 0 4 2
7 11 13 10 9 0 4 2
7 15 13 10 0 9 4 2
10 15 13 10 9 10 0 9 0 4 2
5 15 13 8 4 2
7 15 13 15 9 3 4 2
7 15 13 15 9 0 4 2
9 11 13 10 0 9 1 9 4 2
10 11 13 10 0 9 1 9 4 4 2
9 9 2 15 13 15 3 0 4 2
7 15 13 3 0 4 4 2
6 15 13 10 9 4 2
7 15 13 10 9 4 4 2
9 8 13 15 3 4 2 7 0 2
11 8 13 15 3 4 1 4 2 7 0 2
10 15 15 10 0 9 1 10 9 4 2
11 15 15 10 0 9 1 10 9 4 4 2
9 9 4 3 1 15 13 9 4 2
6 9 4 3 4 4 2
6 10 9 4 3 4 2
7 15 4 3 4 1 4 2
10 11 4 3 15 1 9 4 4 4 2
10 11 13 3 15 1 9 4 4 4 2
9 3 4 15 3 3 4 4 4 2
9 3 13 15 3 3 4 4 4 2
10 15 13 3 0 16 10 9 4 4 2
10 15 4 3 0 16 10 9 4 4 2
9 1 10 9 13 15 3 4 4 2
9 1 10 9 4 15 3 4 4 2
11 16 9 13 15 1 10 0 9 4 4 2
11 16 9 4 15 1 10 0 9 4 4 2
7 10 9 13 4 1 4 2
7 10 9 4 4 1 4 2
8 10 9 13 3 4 1 4 2
8 10 9 4 3 4 1 4 2
10 15 13 3 3 3 3 3 4 4 2
10 15 4 3 3 3 3 3 4 4 2
12 15 13 10 9 3 15 3 0 4 4 4 2
16 15 13 3 1 9 4 4 4 2 7 15 13 3 1 15 2
7 15 13 0 4 1 4 2
9 15 13 3 3 0 4 1 4 2
9 15 4 3 3 0 4 1 4 2
9 15 13 3 3 0 4 1 4 2
8 10 9 13 3 15 9 4 2
13 10 9 13 15 3 3 4 1 10 1 13 9 2
23 1 10 3 0 3 1 4 9 1 10 0 9 1 10 9 13 0 1 15 9 4 4 2
2 13 2
8 11 15 13 1 10 9 13 2
4 15 3 13 2
3 3 13 2
4 9 5 11 2
4 1 9 13 2
7 15 13 10 9 1 4 2
5 11 10 9 13 2
4 15 15 13 2
5 7 15 9 13 2
8 7 15 3 1 10 9 13 2
9 10 9 13 10 9 3 3 0 2
7 9 4 15 9 8 4 2
5 9 13 1 13 2
10 2 11 13 15 2 11 3 1 4 2
5 16 15 0 1 13
13 1 3 0 1 13 9 13 10 9 1 10 9 2
8 15 4 10 0 1 13 9 2
4 13 10 9 2
4 11 0 15 2
11 15 13 3 4 2 15 9 15 15 13 2
12 3 15 3 4 2 15 13 3 9 3 4 2
17 15 13 15 9 4 2 15 4 15 3 1 4 2 15 4 3 2
10 15 13 15 1 15 0 9 0 4 2
5 0 11 9 4 2
5 15 13 15 0 2
7 0 15 9 1 9 4 2
13 3 15 3 13 4 2 15 13 3 9 3 4 2
5 15 4 1 4 2
5 15 9 13 4 2
15 10 9 13 1 10 9 1 12 9 16 4 15 10 9 2
6 15 13 15 8 8 2
4 15 9 11 2
4 15 9 13 2
7 3 0 0 15 11 0 2
6 15 4 8 0 4 2
10 8 15 13 0 3 13 15 9 4 2
4 11 13 15 2
4 13 15 4 2
6 13 15 10 9 0 2
6 13 15 3 3 0 2
15 13 15 1 15 15 4 7 15 13 15 4 15 15 4 2
12 13 15 9 3 7 15 13 15 3 3 3 2
7 13 1 16 15 13 4 2
10 4 15 1 15 0 7 15 13 9 2
7 4 3 3 9 1 10 9
7 13 3 3 3 0 4 2
6 4 3 15 0 4 2
5 13 10 9 0 2
7 13 10 9 0 2 15 2
3 13 12 2
7 6 2 13 3 15 4 2
4 13 3 3 2
6 13 3 3 2 15 2
3 13 0 2
11 13 3 15 3 1 10 9 1 10 9 2
7 0 0 2 13 10 9 2
9 13 10 9 3 7 13 10 9 2
13 13 10 9 3 7 13 10 9 12 9 3 4 2
9 13 1 9 10 9 1 10 9 2
3 13 15 2
5 13 15 3 4 2
4 13 11 3 2
4 15 4 13 2
7 9 13 13 10 9 3 2
10 1 0 9 9 13 13 10 9 3 2
8 8 13 13 15 3 3 3 2
12 15 3 1 10 9 4 13 10 9 10 9 2
8 13 10 9 4 15 9 4 2
1 13
5 15 4 3 13 2
4 15 13 13 2
4 15 13 13 2
5 11 13 13 3 2
6 13 13 10 9 3 2
9 15 13 15 9 3 3 13 4 2
5 3 13 13 15 2
10 3 13 13 15 1 9 3 1 4 2
5 15 13 0 4 2
10 13 15 9 13 15 3 1 9 4 2
8 0 0 13 16 10 9 13 2
6 3 13 2 3 13 2
6 11 13 2 3 13 2
2 6 2
4 13 2 9 2
1 13
2 13 9
3 10 13 9
7 15 9 4 3 9 13 2
5 15 4 13 4 2
9 3 13 13 15 1 10 9 3 2
6 11 13 15 0 13 2
13 15 13 15 3 4 16 15 9 3 9 0 4 2
13 15 13 15 3 4 16 15 9 3 9 13 4 2
13 15 13 15 3 4 16 15 9 1 12 4 4 2
13 15 13 15 3 4 16 15 9 1 12 4 4 2
6 15 9 13 3 4 2
6 15 13 10 9 4 2
8 13 13 15 1 10 9 3 2
6 11 13 15 0 13 2
7 3 13 13 15 3 3 2
11 11 13 7 9 13 13 10 9 1 9 2
11 1 15 13 7 13 13 15 15 0 4 2
6 10 9 4 0 9 2
9 10 9 13 1 10 9 4 4 2
8 15 9 13 4 2 4 2 2
4 11 13 9 2
6 11 13 1 10 11 2
17 3 10 9 1 15 9 13 10 9 15 9 3 4 1 10 11 2
5 15 13 3 4 2
9 3 13 15 11 1 10 9 3 2
6 15 13 3 3 4 2
9 16 15 15 4 2 13 15 15 2
4 13 15 3 2
5 4 15 3 4 2
7 15 13 15 4 1 4 2
9 9 2 10 9 13 0 1 3 2
11 15 13 1 9 11 2 0 13 2 11 2
9 3 3 1 10 9 2 15 13 2
7 13 15 3 3 1 9 2
4 3 13 9 2
7 9 13 8 0 1 15 2
8 15 13 10 9 1 15 9 2
7 15 13 8 1 12 3 2
6 15 9 13 1 9 2
8 9 2 11 13 3 10 9 2
5 15 13 2 9 2
10 15 13 1 0 9 11 1 10 9 2
10 15 13 3 3 12 9 1 15 9 2
7 15 9 13 1 10 9 2
8 1 12 4 8 1 11 4 2
20 3 1 12 13 10 9 2 15 4 3 0 2 15 13 2 15 13 15 3 2
26 3 13 15 1 10 11 11 3 2 15 13 2 15 13 15 3 3 2 15 13 2 15 13 11 4 2
14 3 4 15 3 0 2 16 15 1 15 13 2 2 2
6 15 4 1 0 3 2
9 3 13 10 0 1 0 0 9 2
7 10 9 13 1 8 3 2
24 10 9 13 1 8 4 2 10 9 7 15 9 13 1 10 9 4 4 1 10 9 2 2 2
11 3 13 9 2 9 2 7 15 9 13 2
8 15 13 1 10 13 9 3 2
9 13 9 13 15 3 1 15 8 2
8 3 13 10 0 9 0 9 2
7 15 13 15 9 3 0 2
16 16 10 9 1 13 13 10 9 3 10 0 9 1 10 9 2
14 15 4 1 4 16 10 9 10 1 1 13 9 4 2
14 15 15 0 13 2 13 3 16 15 10 0 9 13 2
8 3 4 15 16 15 15 13 2
15 15 13 16 15 10 9 4 2 1 15 9 13 15 4 2
16 15 13 16 15 1 15 9 9 4 2 1 15 9 13 15 2
10 15 13 3 1 13 1 0 9 4 2
18 15 13 1 10 9 4 4 2 6 2 15 9 1 13 1 0 9 2
10 15 13 3 4 2 10 9 4 0 2
12 6 2 15 9 7 3 4 15 15 9 4 2
9 15 13 8 3 7 13 15 9 2
13 11 13 0 10 9 4 2 16 15 3 0 13 2
8 11 4 0 7 13 10 9 2
7 0 9 13 9 3 4 2
6 0 9 13 9 3 2
11 10 9 4 3 2 11 13 15 0 4 2
11 10 9 4 3 0 16 11 15 15 13 2
14 15 13 0 15 4 2 3 13 15 3 15 0 9 2
15 15 13 0 15 2 15 4 3 3 15 0 1 10 9 2
16 15 13 3 15 9 4 2 15 13 3 16 15 15 9 4 2
12 6 2 15 13 15 9 2 15 13 10 9 2
7 3 13 15 3 1 9 2
12 3 13 15 3 10 9 4 2 1 15 9 2
12 15 13 0 9 9 4 2 15 4 3 4 2
14 15 4 4 1 10 9 2 15 13 3 1 10 9 2
9 15 4 12 9 4 1 10 9 2
7 15 13 3 1 9 4 2
6 15 13 3 1 9 2
8 16 15 9 13 10 9 4 2
7 16 15 9 13 10 9 2
14 3 4 3 0 3 2 3 15 9 13 10 9 4 2
5 15 13 3 4 2
4 15 13 3 2
15 16 15 1 8 13 2 4 10 9 3 0 3 0 3 2
13 15 13 3 1 15 9 4 7 4 3 3 4 2
10 16 15 13 13 15 9 3 3 4 2
10 11 13 15 0 9 1 15 9 4 2
10 11 13 15 0 9 3 1 15 9 2
16 15 4 10 0 9 3 1 10 9 4 7 15 13 15 4 2
16 15 4 10 0 9 3 3 1 10 9 7 15 13 15 4 2
10 15 9 13 3 1 10 9 1 4 2
10 15 9 13 3 3 1 10 9 3 2
9 15 9 13 3 1 10 9 3 2
10 15 13 1 0 9 11 1 10 9 2
11 15 13 1 0 9 11 1 10 9 4 2
10 15 13 3 3 12 9 1 15 9 2
11 15 13 3 3 12 9 1 15 9 4 2
7 15 9 13 1 10 9 2
8 15 9 13 1 10 0 4 2
11 15 13 1 9 11 2 0 13 2 11 2
15 15 13 3 1 15 9 2 16 15 1 9 1 11 4 2
9 13 9 13 15 4 1 15 8 2
9 3 13 10 0 9 0 9 4 2
8 15 13 15 9 3 0 4 2
17 16 10 9 1 13 13 10 9 3 10 0 9 4 1 10 9 2
15 15 4 1 4 16 10 9 10 1 1 13 9 4 4 2
15 15 15 0 13 2 13 3 4 16 15 10 0 9 13 2
10 3 13 10 0 1 0 0 9 4 2
7 10 9 13 1 8 4 2
13 1 12 13 10 9 10 9 1 10 9 4 4 2
12 1 12 13 10 9 10 9 1 10 9 4 2
11 3 1 15 9 13 10 9 3 4 4 2
10 3 1 15 9 4 10 9 3 4 2
15 13 3 1 15 13 1 15 9 16 15 15 9 13 4 2
14 13 3 1 15 13 1 15 9 16 15 15 9 13 2
11 15 13 3 3 1 15 15 9 13 4 2
10 11 13 15 9 3 13 1 15 3 2
10 11 4 15 9 3 13 1 15 4 2
7 10 9 13 0 1 9 2
8 10 9 4 0 1 9 4 2
36 3 4 15 1 10 9 4 2 3 4 3 10 9 2 0 16 15 15 0 3 4 2 15 4 0 0 1 10 9 2 3 13 3 15 0 2
11 2 2 2 2 2 3 13 3 15 4 2
11 2 2 2 2 2 7 3 13 15 15 2
21 9 13 2 1 10 0 9 2 15 9 2 9 7 9 1 10 9 1 12 9 2
9 3 13 3 10 9 16 8 4 2
14 3 13 3 15 4 15 15 9 1 10 9 4 13 2
45 0 9 13 8 1 10 9 8 2 8 0 2 16 3 1 10 9 3 10 9 1 9 1 9 10 9 13 2 10 9 11 13 15 8 7 13 3 16 10 13 9 3 0 4 2
10 16 15 9 13 2 13 15 1 9 2
9 15 4 0 16 15 1 15 4 2
11 15 13 15 11 16 10 9 9 9 4 2
10 15 13 15 16 10 9 9 9 4 2
10 15 13 15 11 16 10 9 9 4 2
9 15 13 15 16 10 9 9 4 2
20 15 13 15 3 3 0 16 15 4 4 2 15 13 3 0 1 15 9 4 2
13 9 4 0 9 11 4 2 9 13 15 3 4 2
15 15 4 3 4 2 13 1 12 9 4 16 10 9 13 2
18 10 9 1 10 0 9 1 11 13 1 10 0 9 11 3 4 4 2
8 1 9 2 3 1 0 9 2
13 11 13 16 15 9 8 10 0 0 9 1 11 2
19 1 9 1 10 9 1 9 11 13 11 10 0 9 11 1 10 0 9 2
18 16 10 9 3 4 4 2 4 15 3 0 16 10 9 11 0 13 2
9 3 8 13 3 3 9 3 3 2
11 9 13 1 15 9 15 3 2 13 11 2
12 1 10 0 9 13 0 10 0 9 4 4 2
13 15 13 10 9 1 10 0 11 7 0 9 11 2
20 2 15 13 10 9 0 1 9 2 2 13 11 1 10 9 1 10 0 9 2
16 10 0 9 11 4 0 16 15 1 10 9 1 11 4 4 2
34 0 9 13 16 10 0 9 1 10 9 11 2 10 0 9 1 11 2 0 1 15 9 3 4 4 7 1 10 0 9 9 4 4 2
13 1 11 15 4 10 9 1 10 9 15 11 13 2
31 2 15 13 16 11 7 11 3 0 15 0 9 4 4 1 10 9 1 10 9 1 0 9 2 2 13 10 0 9 11 2
21 2 7 16 11 15 9 13 1 10 9 1 15 2 3 13 15 3 9 3 2 2
22 10 0 9 11 13 16 9 11 3 4 1 10 9 1 10 9 1 10 0 0 9 2
23 9 13 16 10 9 0 9 4 4 1 10 13 0 9 16 10 9 1 10 9 1 4 2
10 10 9 13 4 16 11 10 9 4 2
17 15 13 3 9 1 10 9 4 1 3 0 9 1 11 7 11 2
15 10 9 4 16 10 0 9 1 3 1 13 1 0 9 2
17 10 0 9 1 11 13 1 10 9 1 10 0 9 1 10 11 2
16 15 9 1 10 9 1 10 11 13 0 3 0 10 9 4 2
19 10 0 9 13 15 9 16 10 9 1 11 10 9 1 0 9 4 4 2
18 15 13 3 16 10 9 1 10 9 0 4 1 10 2 0 2 9 2
10 2 15 4 10 9 1 10 9 2 2
15 8 12 9 7 9 4 13 9 1 0 9 1 11 4 2
20 3 3 1 9 2 7 1 9 13 12 9 16 2 3 13 10 0 9 11 2
12 10 0 9 13 3 1 9 7 9 10 9 2
37 10 9 13 0 12 12 13 7 15 0 12 0 9 5 7 3 7 3 13 3 10 0 9 1 12 12 9 1 4 2 3 12 9 1 10 9 2
16 1 15 9 4 15 9 4 1 9 2 9 2 9 7 9 2
19 1 9 4 4 15 15 3 1 10 0 9 1 1 3 0 9 9 4 2
28 10 15 9 4 1 13 9 4 1 0 0 2 15 0 4 1 0 9 7 10 9 15 10 0 9 15 13 2
12 11 4 10 0 9 1 9 1 11 7 11 2
27 1 10 12 9 0 0 9 13 1 0 9 10 13 9 2 7 9 13 15 3 3 1 9 1 15 8 2
19 12 9 1 10 9 13 1 11 15 9 1 11 7 3 0 1 10 9 2
15 10 9 1 13 9 15 9 1 10 0 9 1 10 9 2
20 3 0 13 3 9 1 9 1 15 13 1 9 1 3 3 10 9 7 15 2
12 11 13 10 13 12 9 10 16 12 9 4 2
13 15 12 8 13 13 3 1 10 9 1 15 9 2
25 10 0 9 1 15 9 13 8 8 10 0 9 13 3 1 10 9 3 0 9 1 10 9 4 2
17 2 10 15 9 15 15 13 4 2 4 15 1 10 9 3 3 2
10 15 13 2 15 13 15 15 1 9 2
12 7 10 13 9 13 15 15 3 3 4 2 2
14 7 9 13 3 10 0 9 16 9 10 9 1 4 2
16 3 13 10 9 1 10 0 9 10 9 0 16 11 1 11 2
18 8 13 10 9 1 10 9 7 13 3 1 10 9 1 15 13 9 2
13 3 1 9 7 9 8 13 10 9 1 10 9 2
12 2 9 7 9 13 8 15 2 2 13 8 2
5 8 4 0 4 2
8 15 13 3 0 1 15 4 2
24 12 9 3 13 15 9 1 10 9 1 8 3 1 11 3 15 10 9 1 15 9 13 4 2
7 1 10 9 13 8 3 2
5 15 13 1 9 2
14 1 9 1 9 13 15 8 15 1 4 1 10 11 2
13 7 3 13 3 0 9 1 10 0 0 9 8 2
12 8 2 2 15 9 13 3 1 0 9 2 2
24 8 2 12 2 13 3 1 10 9 1 10 0 0 9 1 15 1 12 1 15 15 9 13 2
15 15 13 1 11 1 11 1 15 1 15 9 1 13 4 2
36 10 0 9 4 15 0 3 3 5 9 4 0 3 0 7 13 3 3 16 15 3 10 9 1 10 9 13 5 7 15 13 3 15 9 3 2
9 2 15 9 4 0 3 4 2 2
15 10 13 9 13 15 3 16 15 3 4 4 1 10 11 2
10 9 11 13 15 3 3 3 1 4 2
16 1 1 10 9 13 8 9 16 15 0 1 4 1 10 9 2
8 2 15 9 13 15 9 3 2
20 16 9 1 13 13 15 15 4 16 15 3 3 1 10 9 0 1 4 2 2
12 12 9 1 10 9 13 10 9 1 12 9 2
16 16 8 7 15 0 8 4 3 8 1 10 9 1 8 4 2
11 1 0 9 0 10 0 11 10 9 3 2
10 3 10 9 1 15 9 8 4 4 2
10 1 10 9 1 9 13 10 9 3 2
14 15 13 9 1 9 11 15 13 1 4 1 10 9 2
8 2 15 13 2 13 1 15 2
7 15 4 3 10 9 2 2
9 13 1 11 13 15 1 10 9 2
7 11 13 3 2 13 8 2
6 2 15 9 15 3 2
7 15 4 3 10 9 2 2
16 8 13 16 15 10 9 4 2 1 10 9 1 10 9 8 2
6 15 9 13 15 4 2
15 11 7 3 2 3 0 15 4 2 3 0 15 3 4 2
12 2 15 13 16 15 9 1 10 9 0 4 2
7 15 9 13 15 4 2 2
27 10 9 1 10 9 12 1 10 9 2 12 12 12 12 2 4 10 0 9 1 10 9 15 9 1 11 2
13 1 10 9 13 10 0 9 8 0 1 15 8 2
25 1 11 13 10 9 1 10 0 0 9 2 15 1 11 3 0 16 10 9 13 2 10 0 9 2
13 8 1 12 9 13 10 9 10 0 9 1 11 2
20 1 10 9 1 10 9 2 2 15 13 0 0 3 2 10 9 3 1 9 2
9 10 9 13 8 15 8 11 9 2
11 1 11 13 15 3 1 10 9 1 11 2
12 1 10 16 12 9 1 9 4 15 3 0 2
9 10 9 1 15 9 4 15 9 2
6 9 13 15 15 9 2
8 10 0 9 13 10 0 9 2
17 10 9 1 8 13 1 11 12 9 1 10 0 9 1 10 9 2
12 2 0 9 4 15 8 4 2 1 15 9 2
13 15 13 15 8 16 3 3 1 4 1 15 9 2
7 15 13 0 8 1 4 2
7 1 15 9 13 10 9 2
16 15 4 3 3 0 16 15 13 16 15 1 15 4 4 2 2
20 10 0 9 4 0 2 7 0 1 13 9 2 4 1 10 9 1 12 9 2
16 10 9 13 15 3 7 1 0 16 1 0 9 3 1 11 2
20 10 9 13 1 10 9 1 11 10 12 9 2 10 9 13 13 7 13 3 2
31 11 13 3 3 10 2 3 13 2 9 7 1 9 13 15 12 9 1 10 0 9 2 8 7 2 1 10 9 2 11 2
18 9 8 13 3 8 1 10 9 4 3 15 9 1 10 9 4 4 2
20 1 11 13 11 11 11 2 15 3 3 13 1 9 13 1 11 2 12 2 2
16 1 10 15 0 9 2 1 8 2 13 11 7 11 1 15 2
10 10 9 13 3 11 3 2 12 2 2
12 11 4 1 10 9 1 12 9 10 0 9 2
13 11 13 1 12 1 11 2 1 10 9 1 11 2
26 1 11 13 11 3 10 9 15 15 3 0 2 1 12 9 1 12 9 2 1 10 0 9 13 4 2
9 3 13 11 3 1 12 1 11 2
17 1 10 9 13 10 9 3 0 13 4 1 15 8 2 12 2 2
17 9 8 13 3 8 12 9 3 2 3 15 8 1 12 13 4 2
10 10 9 4 0 4 1 10 0 9 2
10 11 13 3 3 10 13 9 1 4 2
31 3 13 10 0 9 10 0 9 3 1 10 12 9 2 1 9 3 1 10 13 0 9 2 15 10 9 1 9 8 13 2
31 15 4 3 3 10 9 1 10 1 10 10 0 0 9 1 11 2 7 3 15 0 13 10 9 13 1 8 10 0 9 2
20 1 10 9 1 10 0 9 4 10 9 1 10 9 4 1 10 0 9 11 2
13 8 4 1 10 0 9 1 15 0 0 9 4 2
8 10 0 9 13 3 3 3 2
16 11 2 9 1 10 9 2 13 15 1 10 9 3 0 4 2
16 10 0 9 4 1 10 0 9 10 0 9 1 10 0 9 2
19 11 13 2 1 10 0 9 2 3 1 10 0 9 1 10 0 9 4 2
26 9 11 13 9 11 1 3 2 12 2 2 1 10 9 1 9 8 15 1 8 3 1 9 4 4 2
13 3 13 10 9 16 15 3 3 1 15 9 4 2
20 10 13 11 13 2 16 3 3 3 1 15 9 2 3 1 10 15 0 9 2
14 1 10 0 9 13 10 9 10 0 13 7 13 9 2
22 8 2 15 1 8 13 2 13 15 4 1 10 9 1 10 0 0 9 2 12 2 2
14 10 0 9 1 0 9 13 3 10 9 9 0 3 2
10 7 10 10 9 13 10 13 11 15 2
25 10 9 13 10 9 3 1 12 9 2 16 1 10 9 3 9 11 1 10 9 2 0 2 13 2
12 15 4 10 0 9 2 15 4 10 0 9 2
12 9 1 9 13 1 0 9 9 1 0 9 2
7 3 13 10 0 9 0 2
12 7 3 13 1 9 1 15 13 9 7 9 2
19 1 8 12 9 13 9 8 3 10 0 9 15 13 1 15 13 1 4 2
12 3 4 10 9 15 7 15 9 11 3 0 2
9 12 1 10 12 9 13 15 9 2
18 3 13 15 3 3 3 1 10 9 7 1 10 0 9 1 10 9 2
11 3 13 15 1 10 0 1 10 0 9 2
3 13 3 2
14 8 2 2 15 13 16 15 1 15 9 0 4 4 2
6 15 13 16 15 4 2
14 1 15 11 13 4 15 0 15 1 15 9 1 13 2
17 16 3 10 0 13 2 4 15 3 0 10 0 3 1 13 2 2
12 8 13 15 0 1 0 9 1 15 0 9 2
7 15 13 1 15 9 4 2
7 2 10 9 13 15 4 2
10 3 13 15 10 9 7 4 15 3 2
6 15 4 3 1 15 2
7 10 9 13 3 4 2 2
22 10 9 4 3 15 10 9 1 8 16 1 10 9 15 15 10 0 9 3 13 4 2
31 10 9 2 15 1 15 13 1 8 7 8 9 13 1 10 0 9 2 13 3 8 15 1 10 0 9 1 10 9 4 2
15 10 9 4 0 2 12 9 1 10 9 11 2 7 9 2
9 0 13 15 8 10 9 3 4 2
15 10 9 2 15 10 0 9 1 10 11 16 0 9 13 2
19 10 9 15 10 9 3 1 10 9 13 4 2 0 16 15 13 1 9 2
14 9 1 10 13 9 3 3 9 15 1 11 4 4 2
8 11 4 10 9 3 9 13 2
17 3 0 4 3 10 9 15 8 1 10 13 9 1 10 11 4 2
17 7 3 13 4 10 9 16 8 13 1 10 9 1 15 9 11 2
18 7 3 0 4 15 16 10 0 9 2 0 9 11 2 1 9 13 2
18 15 13 3 3 1 3 0 9 2 10 9 1 12 9 2 12 13 2
22 1 10 0 0 13 8 15 9 4 2 3 16 11 7 10 9 11 2 15 0 9 2
23 1 10 0 0 9 15 3 10 9 2 3 16 12 15 2 7 0 0 4 16 9 3 2
17 3 13 8 2 1 15 10 0 9 9 2 7 15 12 9 13 2
2 12 2
3 3 9 2
7 7 3 13 4 10 9 2
22 7 16 15 10 9 1 11 3 3 4 4 4 2 4 4 2 7 3 1 15 9 2
41 10 9 13 15 1 11 1 10 9 2 13 15 7 13 3 1 10 9 1 10 9 1 10 9 3 15 15 3 15 1 9 13 1 4 10 9 13 1 10 9 2
9 3 13 15 15 9 3 1 4 2
8 6 2 15 4 15 9 4 2
10 2 1 10 9 13 15 3 3 13 2
11 15 13 3 1 10 9 0 0 3 2 2
35 7 6 2 15 4 13 2 7 3 3 0 2 2 0 9 13 15 3 3 16 15 3 3 13 4 7 3 13 15 1 10 0 3 3 2
11 16 15 3 3 4 2 4 10 9 0 2
15 7 15 13 3 9 1 10 9 2 3 15 0 13 4 2
18 15 4 0 1 11 1 13 2 7 15 4 15 11 3 3 4 2 2
22 10 9 15 3 1 10 9 1 11 1 10 9 4 4 2 4 10 9 1 10 11 2
27 7 1 11 2 3 11 7 1 8 1 10 2 0 2 9 13 15 10 9 10 9 0 13 1 10 9 2
13 2 15 13 11 3 16 10 9 1 15 13 4 2
20 15 4 3 16 15 1 10 9 3 0 13 2 7 15 4 0 3 0 2 2
6 3 9 8 4 0 2
17 2 15 3 13 2 4 10 9 1 15 15 15 15 9 4 4 2
10 15 13 4 16 11 3 0 4 4 2
9 3 13 15 15 3 3 4 2 2
6 9 4 1 15 0 2
13 2 1 10 0 9 1 10 9 13 15 0 4 2
17 16 11 15 4 2 16 8 3 1 9 4 2 13 15 3 4 2
13 15 4 10 0 9 15 15 13 1 12 7 12 2
8 10 12 15 13 1 15 3 2
9 8 13 4 4 16 15 4 4 2
10 11 11 13 15 16 15 10 9 4 2
10 1 15 10 9 13 15 3 4 4 2
12 15 13 15 1 4 2 15 13 15 0 4 2
9 6 2 15 13 15 1 11 4 2
7 3 4 15 9 0 2 2
12 2 10 9 4 3 1 10 9 1 4 2 2
9 8 13 1 15 9 1 10 9 2
18 0 13 15 15 3 1 10 0 9 15 15 11 1 10 11 13 3 2
8 4 7 4 2 13 10 9 2
11 10 0 9 1 10 9 13 1 9 9 2
21 1 10 0 9 1 11 13 10 9 3 3 1 10 9 1 9 1 9 1 4 2
14 1 10 0 7 0 9 13 15 10 13 9 3 4 2
17 1 15 13 1 10 0 9 4 10 9 1 10 9 8 3 4 2
8 10 9 13 8 10 0 9 2
5 10 9 16 8 2
16 12 9 16 15 1 8 15 9 13 4 2 4 15 9 0 2
18 11 13 1 12 7 12 1 9 1 11 3 13 3 15 9 3 4 2
20 15 13 8 15 9 1 9 2 3 15 15 3 0 13 1 10 9 16 9 2
11 2 15 4 3 4 16 15 3 15 4 2
16 15 13 16 8 3 3 4 4 16 15 15 0 4 4 2 2
8 11 13 13 3 10 9 3 2
22 2 11 13 10 0 9 1 15 4 4 2 7 3 13 15 9 3 15 0 4 2 2
11 1 10 9 1 10 11 13 3 15 9 2
17 10 9 13 0 10 9 7 15 9 13 15 15 9 15 9 4 2
10 3 1 10 9 13 15 1 9 4 2
13 10 9 13 15 1 10 11 3 0 1 10 9 2
18 8 2 10 9 1 10 9 1 10 11 2 13 16 3 3 10 9 2
18 15 13 1 10 9 1 12 9 2 1 12 9 2 1 15 3 8 2
17 8 2 2 15 4 10 9 2 3 0 3 2 10 9 9 2 2
25 15 9 2 3 4 15 2 7 10 9 13 9 1 9 1 10 9 4 16 10 9 8 1 13 2
3 15 13 2
26 3 13 8 2 11 2 3 1 10 9 3 2 7 1 10 9 1 11 13 10 9 3 13 4 4 2
10 10 9 13 10 0 9 3 1 9 2
16 9 2 2 15 13 16 10 9 1 15 3 10 0 9 4 2
13 15 13 10 9 0 4 2 7 3 0 15 2 2
14 13 15 13 1 10 0 9 3 3 9 1 15 9 2
16 1 15 13 1 10 9 13 9 3 1 10 9 1 12 9 2
23 11 4 3 3 1 12 9 4 2 7 9 2 11 7 11 13 10 0 1 15 3 4 2
23 10 2 9 2 13 11 2 7 0 9 3 0 9 1 15 1 2 11 2 11 7 8 2
15 3 3 13 11 15 1 10 9 1 8 7 15 13 11 2
15 2 15 13 16 11 1 10 9 1 15 9 4 4 2 2
16 8 13 10 9 1 10 9 0 10 9 10 9 0 1 4 2
7 15 13 10 0 9 3 2
9 3 13 10 9 1 9 7 9 2
16 9 13 15 2 7 3 8 2 8 7 11 13 1 10 9 2
9 8 13 3 16 10 9 4 4 2
12 2 10 9 13 3 4 16 15 4 4 2 2
20 13 4 10 0 9 3 3 1 4 16 15 1 10 0 9 12 9 9 13 2
12 2 15 13 0 16 15 1 15 1 13 2 2
12 13 4 0 2 11 0 2 7 11 4 0 2
14 15 13 1 15 13 3 3 3 9 16 16 1 4 2
14 1 8 2 0 2 13 15 3 10 9 1 10 9 2
11 11 2 2 15 13 0 1 15 9 4 2
21 16 15 13 16 15 1 8 4 2 13 15 16 15 1 15 15 3 0 4 4 2
12 7 1 10 9 1 10 9 13 15 1 9 2
22 1 10 13 12 9 13 15 12 9 4 2 3 15 1 10 9 16 9 1 13 2 2
22 11 13 15 0 4 4 1 10 9 16 9 2 3 0 4 15 4 16 10 13 9 2
6 15 9 13 0 0 2
28 1 10 0 9 3 15 1 10 9 13 5 11 2 11 2 11 7 11 5 13 15 3 0 1 10 9 4 2
11 1 10 9 1 10 9 0 9 13 15 2
25 15 9 13 15 1 10 0 11 2 7 15 9 13 1 15 9 1 10 13 9 3 3 4 4 2
8 9 13 15 3 3 16 9 2
14 10 9 1 10 9 4 0 2 9 13 3 3 0 2
11 2 15 13 15 3 0 1 10 9 4 2
11 1 12 9 13 15 9 1 15 9 2 2
17 3 13 9 8 1 11 16 15 2 7 9 8 2 9 1 13 2
12 10 8 9 11 13 4 15 8 3 1 4 2
12 10 9 13 1 12 8 12 1 11 4 4 2
14 10 0 9 13 15 11 9 1 10 9 1 10 9 2
9 1 11 4 10 9 3 0 4 2
24 1 10 9 1 8 4 11 3 4 10 9 3 1 11 1 4 4 2 8 0 0 1 8 2
31 10 0 9 1 10 9 1 10 9 2 15 3 0 1 11 4 4 2 4 10 9 1 10 9 1 10 0 9 2 8 2
14 15 4 12 4 3 1 11 2 15 1 10 13 9 2
23 10 9 1 11 0 1 11 4 10 0 1 10 9 1 9 15 8 4 4 1 15 8 2
15 1 11 13 9 1 10 9 11 2 11 2 11 7 11 2
14 9 16 10 9 1 11 4 4 4 2 4 3 0 2
13 1 12 13 10 0 9 11 1 10 0 9 11 2
15 1 10 0 9 1 10 11 13 15 10 0 9 1 11 2
13 11 13 15 13 1 10 11 0 1 10 0 9 2
12 2 15 13 9 4 1 9 2 2 13 15 2
23 7 10 13 9 13 15 10 11 2 15 11 1 3 13 2 3 3 10 9 13 1 13 2
19 1 10 9 1 11 4 1 10 9 1 11 2 11 7 11 10 9 4 2
19 15 13 10 0 9 1 10 11 7 15 13 15 9 3 4 4 1 11 2
8 11 13 10 9 3 1 4 2
22 0 16 9 11 11 10 9 10 9 1 4 0 13 4 2 4 11 4 1 15 9 2
12 15 13 2 1 9 2 4 4 1 10 9 2
16 16 15 13 1 15 13 1 10 11 2 13 15 15 3 0 2
15 11 4 3 4 1 10 9 16 10 11 11 11 1 13 2
22 10 9 13 15 9 8 1 8 10 9 4 4 1 10 0 9 16 10 11 1 13 2
22 10 13 9 13 10 11 1 0 9 0 12 13 9 7 9 0 16 15 9 1 13 2
21 0 13 7 9 13 11 9 1 10 9 1 9 11 10 9 1 1 10 0 9 2
18 11 13 2 2 16 10 11 3 13 2 4 15 10 9 1 15 9 2
11 15 13 10 9 4 1 15 9 7 9 2
10 15 4 9 1 10 9 1 10 9 2
17 9 15 15 3 13 1 10 11 2 13 15 3 1 15 13 2 2
13 11 13 10 9 0 16 10 11 11 11 1 13 2
26 15 13 0 1 9 1 15 0 9 1 10 9 15 0 9 1 4 1 10 9 1 10 9 1 11 2
21 11 2 11 2 11 2 11 7 11 13 0 10 9 1 11 1 10 9 1 8 2
5 11 2 11 2 11
6 7 11 4 3 3 2
17 10 9 1 10 11 13 1 10 9 10 9 7 10 9 1 4 2
15 1 10 0 9 4 1 9 4 1 15 13 1 10 9 2
12 10 9 8 13 10 0 9 1 12 12 9 2
26 1 10 9 1 10 9 8 2 3 12 10 9 13 4 4 2 4 10 9 9 7 9 0 8 4 2
6 8 13 10 9 3 2
10 15 13 15 13 16 10 11 3 4 2
16 2 15 4 1 15 10 9 16 3 10 15 11 1 4 4 2
9 10 0 9 4 3 0 1 15 2
12 7 15 16 3 3 3 3 10 0 9 13 2
11 13 3 15 2 4 15 3 3 3 0 2
13 10 9 9 13 4 3 15 10 9 0 13 2 2
18 1 10 9 16 15 0 4 16 10 9 1 11 4 2 13 15 3 2
9 2 15 13 3 3 1 10 9 2
9 15 13 16 15 3 0 4 2 2
11 10 0 11 1 15 9 13 1 10 9 2
12 8 4 0 8 16 15 1 4 1 15 9 2
10 2 15 4 1 10 0 9 4 2 2
19 11 13 10 3 0 9 1 12 9 15 1 9 1 10 0 9 1 11 2
10 10 0 0 9 13 3 2 8 8 2
12 3 13 4 3 0 10 0 9 1 11 4 2
12 7 16 10 9 1 9 7 9 3 4 4 2
13 9 16 1 4 13 10 0 1 15 9 3 3 2
9 15 13 10 9 1 10 9 4 2
15 2 15 4 0 3 9 1 10 9 10 9 1 9 13 2
20 15 16 3 13 15 15 16 10 9 16 3 13 1 10 9 1 4 4 2 2
17 13 9 13 10 0 9 8 1 10 0 9 1 10 0 9 13 2
12 15 4 0 13 2 7 15 4 3 10 9 2
15 15 0 9 7 0 9 2 8 2 4 4 1 0 9 2
12 2 15 0 9 13 15 3 13 1 15 9 2
4 3 3 3 2
5 0 3 3 2 2
14 9 11 13 10 9 1 11 2 1 10 9 1 11 2
8 15 4 10 9 1 0 3 2
11 0 1 8 13 15 10 9 1 9 11 2
10 2 3 13 15 4 15 9 4 2 2
6 3 13 3 1 11 2
10 8 1 12 13 10 0 9 15 8 2
9 0 16 15 0 3 3 0 4 2
12 2 15 13 16 15 15 15 15 3 4 4 2
5 15 4 3 0 2
20 3 4 15 0 1 15 1 10 9 15 15 3 3 4 4 1 15 9 2 2
21 16 8 1 11 15 0 9 1 10 9 13 2 13 11 10 9 16 1 10 9 2
23 15 13 15 8 16 3 3 1 4 1 15 12 13 8 7 10 9 15 3 1 15 13 2
6 3 4 9 3 9 2
14 2 3 13 4 15 0 15 0 4 16 15 0 4 2
4 15 4 12 2
7 8 2 8 9 13 15 2
22 15 4 3 12 9 7 3 13 15 3 10 9 1 10 9 1 15 9 1 4 4 2
10 3 4 10 9 1 10 9 8 2 2
14 2 15 4 10 0 9 1 9 2 0 1 10 9 2
6 9 7 9 13 8 2
22 15 13 4 10 9 1 10 9 1 10 9 1 4 2 10 9 15 1 15 9 13 2
7 15 4 0 1 10 0 2
17 10 0 15 13 10 0 9 1 15 0 3 9 0 1 4 2 2
14 2 3 16 15 13 1 13 2 13 15 9 0 9 2
8 0 13 15 15 3 0 4 2
6 8 16 15 4 4 2
9 3 3 13 15 16 15 0 4 2
11 15 13 15 9 1 15 15 9 4 2 2
9 2 0 13 15 3 3 3 13 2
12 9 13 4 7 13 2 3 13 15 15 3 2
7 15 4 3 1 15 12 2
16 7 15 13 3 3 15 15 3 1 15 9 3 4 4 4 2
9 10 9 7 10 9 7 10 9 2
11 1 10 0 9 13 15 1 15 9 2 2
13 3 4 15 3 3 3 10 0 1 10 0 9 2
21 15 9 4 0 1 15 9 2 2 0 2 3 13 10 9 15 3 3 4 2 2
18 0 1 9 13 15 0 10 9 3 1 15 9 3 10 9 1 11 2
30 10 9 11 13 1 9 2 16 9 2 15 1 15 9 2 11 13 1 10 9 7 11 2 6 15 13 3 3 3 2
9 3 16 11 9 1 3 2 8 2
11 10 9 1 12 13 3 15 9 1 8 2
10 2 15 13 1 12 9 1 10 9 2
8 3 16 10 9 1 15 9 2
26 15 13 16 15 3 10 0 9 4 1 15 15 9 13 2 7 1 15 10 9 1 10 9 13 2 2
15 11 9 4 1 15 9 4 2 10 9 13 0 15 9 2
12 1 11 4 15 9 10 0 9 3 0 9 2
19 10 9 4 0 2 13 10 9 1 10 0 0 9 1 8 2 11 2 2
19 15 1 9 4 2 13 1 9 2 13 15 1 10 9 15 9 1 11 2
10 7 10 9 0 13 10 9 3 3 2
21 10 9 9 13 10 9 3 2 10 9 4 1 9 1 12 9 1 15 9 4 2
9 10 9 4 10 9 2 15 9 2
2 9 2
23 2 16 13 15 9 4 2 2 13 1 9 10 9 10 9 1 1 15 9 1 15 8 2
21 16 15 0 4 2 13 1 4 2 7 10 9 1 10 0 9 4 13 2 8 2
16 10 9 9 13 3 15 8 1 9 1 15 9 2 0 13 2
23 1 11 8 13 13 9 1 9 4 2 7 3 10 11 13 10 0 9 16 3 1 4 2
25 8 2 10 9 1 8 2 13 3 2 1 9 0 4 3 2 1 12 9 2 1 15 9 4 2
13 10 0 9 11 13 10 9 1 10 9 1 11 2
20 15 13 15 15 9 1 10 9 2 7 15 9 13 15 9 3 4 4 4 2
8 1 11 13 16 3 3 3 2
21 10 9 9 13 10 2 13 0 9 1 9 2 2 8 2 9 2 3 3 4 2
20 16 15 1 2 9 2 3 1 2 9 2 13 2 13 3 1 15 0 9 2
5 7 15 13 3 2
9 10 9 0 15 9 15 0 9 2
32 10 9 2 10 0 9 13 1 10 0 0 9 1 11 2 12 2 2 13 10 9 4 2 7 9 4 3 0 9 16 9 2
21 3 13 10 9 15 3 3 1 10 9 9 3 13 3 10 0 9 1 10 9 2
26 1 10 0 9 8 2 12 2 13 9 1 15 0 0 2 6 2 1 10 0 9 10 9 1 3 2
5 9 4 3 9 2
13 9 16 1 11 1 4 1 9 9 1 0 9 2
31 0 9 13 10 9 1 11 2 8 2 15 4 1 10 0 9 2 7 1 10 0 2 11 13 4 2 10 9 4 4 2
8 0 13 11 10 9 1 4 2
13 15 13 10 9 1 10 9 1 15 3 1 4 2
10 0 13 10 9 15 13 1 9 4 2
28 10 9 8 4 10 0 9 1 10 9 15 15 1 4 13 1 15 9 2 10 15 4 3 7 3 3 9 2
42 0 9 13 10 9 2 0 9 15 1 0 13 2 9 13 10 9 2 13 11 2 3 1 10 3 0 7 0 9 4 9 0 2 3 0 7 15 13 1 10 9 2
41 1 10 9 4 10 9 1 15 15 0 9 13 7 13 16 15 15 16 10 0 9 2 16 15 3 10 9 13 0 10 9 3 16 10 9 3 10 9 4 4 2
15 11 13 3 15 15 4 2 15 13 3 0 15 9 3 2
7 15 13 8 3 9 3 2
18 15 4 1 15 9 0 3 2 3 15 4 4 1 9 1 10 9 2
14 8 12 9 13 3 4 15 9 1 4 4 16 11 2
27 10 9 13 3 1 0 9 1 0 16 11 7 11 15 1 15 9 1 9 3 3 1 15 9 13 4 2
31 10 13 9 11 2 15 1 10 13 9 1 10 9 2 13 15 13 0 1 0 9 4 2 7 13 3 3 0 9 3 2
16 1 15 13 0 9 10 9 15 9 13 2 9 13 16 3 2
11 1 11 13 12 0 2 3 1 10 9 2
28 13 16 15 3 15 15 1 15 9 4 16 10 9 1 9 1 9 2 13 11 3 1 11 2 2 4 0 2
14 3 13 15 9 4 16 15 15 9 13 1 10 9 2
29 0 9 4 15 3 1 11 7 13 10 9 2 15 13 3 1 0 9 7 0 9 2 3 1 13 0 9 2 2
24 3 13 11 10 0 9 8 2 10 9 3 2 10 9 2 6 13 2 4 1 15 3 0 2
14 1 15 9 13 11 1 11 13 15 3 1 10 9 2
19 9 13 10 9 4 1 10 0 9 16 0 9 15 3 1 10 9 13 2
23 3 13 15 3 2 7 15 9 0 13 15 1 15 15 2 10 9 2 15 15 0 13 2
14 3 13 15 9 1 11 2 9 2 3 3 10 9 2
12 3 13 10 9 1 10 9 1 10 9 0 2
13 15 13 15 1 10 9 15 0 4 3 1 4 2
15 16 15 1 10 0 9 1 0 13 2 13 10 9 8 2
37 2 16 9 9 13 16 11 9 4 7 16 15 3 3 4 4 2 4 15 9 0 1 4 2 9 13 1 0 9 3 0 10 0 9 4 2 2
16 3 3 13 9 1 10 9 0 9 10 9 16 15 0 13 2
16 13 15 15 3 4 2 3 4 15 10 13 9 8 1 9 2
22 10 0 0 9 1 10 0 9 8 4 9 1 11 1 15 13 1 10 9 8 4 2
23 10 9 13 1 12 9 9 1 10 9 1 4 16 15 1 3 13 7 1 15 9 13 2
8 0 3 13 15 1 15 9 2
9 10 9 13 15 13 3 1 4 2
24 10 9 13 1 10 9 1 11 1 11 10 0 9 4 8 9 1 10 0 9 1 15 9 2
16 1 10 9 1 10 9 1 11 13 1 12 10 0 0 8 2
23 10 9 1 10 9 13 16 10 13 9 7 10 9 1 10 9 10 9 1 15 4 4 2
16 10 0 9 1 11 1 10 11 13 15 9 3 12 9 4 2
20 10 9 13 1 8 2 3 10 11 15 9 1 9 1 9 1 9 7 9 2
13 1 10 9 4 8 9 4 1 15 12 12 9 2
21 12 0 0 9 13 13 1 15 9 1 0 9 4 4 1 10 9 1 10 9 2
41 10 9 1 10 9 1 9 13 11 4 16 10 0 0 9 11 1 11 7 15 8 1 11 10 9 4 4 3 0 13 4 4 7 10 9 1 10 9 4 4 2
21 10 9 1 10 9 0 13 9 3 1 10 9 1 9 8 2 9 1 9 11 2
23 1 10 9 1 9 4 10 9 3 10 9 13 4 4 10 0 9 1 10 15 0 9 2
20 2 15 13 10 9 1 15 13 2 7 3 15 9 7 10 9 1 9 2 2
36 1 10 9 1 10 9 1 10 9 13 9 11 0 1 4 4 1 3 10 9 1 15 9 10 0 9 4 1 3 1 13 1 15 0 9 2
16 3 13 15 16 12 1 10 12 9 1 15 2 9 3 8 2
25 12 9 1 12 7 12 9 1 11 7 11 4 11 1 10 9 1 11 1 15 9 1 9 4 2
12 10 12 9 13 15 1 10 9 1 10 9 2
18 10 9 13 16 10 9 1 10 9 7 15 9 10 9 0 4 4 2
24 10 9 1 10 1 10 9 13 1 10 9 12 9 0 1 10 9 4 7 13 10 9 3 2
20 9 13 3 4 1 4 2 7 1 9 1 10 9 4 10 9 1 4 4 2
7 10 0 9 13 10 9 2
33 1 10 9 1 10 11 1 11 1 8 2 15 9 10 9 2 12 2 7 10 9 2 12 2 1 15 8 2 11 2 8 4 2
20 12 15 0 1 10 9 1 1 9 12 9 4 3 13 2 1 15 9 0 2
16 1 10 9 1 11 13 10 9 1 10 9 1 10 9 13 2
16 10 13 9 2 15 13 2 7 10 9 4 1 10 9 4 2
16 1 9 1 10 9 1 8 1 11 4 11 12 9 13 4 2
20 15 13 1 10 9 9 7 9 15 1 10 9 1 10 9 1 10 9 13 2
10 1 10 9 13 10 9 1 0 9 2
8 10 9 13 3 1 10 9 2
18 15 4 1 10 9 1 10 9 4 2 15 13 9 1 9 7 9 2
11 10 9 4 1 10 11 7 10 9 4 2
7 15 13 3 0 1 9 2
21 10 0 9 13 1 10 9 1 11 1 11 10 9 4 1 10 9 9 1 11 2
18 10 0 1 10 3 13 9 0 9 2 3 9 4 4 2 4 4 2
16 10 9 1 12 9 1 10 9 13 8 10 9 15 9 4 2
18 12 9 1 11 4 1 10 9 1 11 1 11 4 1 10 0 9 2
13 1 10 9 1 10 9 13 15 13 1 10 9 2
15 10 9 7 9 8 4 1 10 9 1 11 1 11 4 2
21 8 13 3 16 9 7 13 1 10 9 11 1 10 11 2 3 1 15 9 8 2
12 8 4 12 9 4 2 3 13 10 9 3 2
15 1 10 9 12 7 12 13 11 9 1 10 0 0 9 2
12 1 10 0 11 13 15 3 16 10 0 9 2
27 1 15 9 11 4 11 1 0 9 8 4 2 0 9 7 9 1 10 9 11 1 15 8 2 11 2 2
12 11 13 9 9 10 9 1 10 11 1 11 2
12 1 15 9 13 15 1 0 9 9 16 9 2
12 9 2 1 9 9 2 13 1 10 0 9 2
8 15 9 13 15 13 3 4 2
15 8 4 1 12 10 0 9 11 1 10 9 1 11 9 2
14 0 4 1 8 9 8 1 10 9 1 9 7 9 2
6 3 4 15 9 11 2
11 1 15 9 4 15 8 10 9 8 4 2
13 15 4 1 15 9 1 10 0 9 1 10 11 2
15 0 4 10 9 1 8 2 15 13 1 10 9 4 4 2
15 10 0 9 8 4 11 1 0 9 4 1 15 9 11 2
10 11 4 15 1 10 9 1 15 8 2
7 15 13 3 9 1 9 2
17 11 13 10 9 7 4 1 12 4 16 9 1 15 8 1 11 2
8 3 10 0 9 13 15 9 2
19 11 2 0 2 8 2 1 9 1 15 9 2 13 15 16 12 12 9 2
16 15 13 15 1 10 9 2 1 8 1 8 2 9 7 9 2
9 7 15 4 10 9 3 15 13 2
15 8 4 0 1 12 1 11 2 11 2 1 10 0 9 2
15 15 4 4 1 9 7 9 8 7 13 16 9 3 9 2
8 15 0 13 13 15 3 0 2
47 9 1 2 8 2 2 12 2 13 15 10 16 12 9 1 15 9 2 3 2 11 2 2 12 2 2 2 8 2 2 12 2 2 2 8 2 2 12 2 7 2 8 2 2 12 2 2
11 15 13 3 9 1 12 9 1 15 9 2
16 11 2 15 13 1 10 0 9 2 4 9 3 13 16 9 2
12 15 13 3 1 9 16 2 8 2 1 8 2
10 3 13 15 8 3 1 8 7 8 2
24 10 0 9 11 13 8 2 11 2 1 10 9 11 1 12 12 9 2 3 12 12 9 2 2
17 8 2 11 2 13 2 13 7 13 9 1 9 1 15 0 9 2
13 1 10 0 9 1 10 9 1 13 9 0 9 2
16 15 8 13 0 12 12 9 1 12 9 7 13 1 12 9 2
16 9 2 9 3 13 16 8 7 11 2 4 9 1 0 9 2
12 15 8 13 3 3 1 10 9 1 10 9 2
17 10 0 9 3 8 9 7 9 4 11 7 11 0 4 1 9 2
24 15 8 10 9 7 9 1 10 9 1 11 2 10 9 1 10 9 15 10 9 1 9 13 2
17 11 13 16 11 12 9 13 1 10 0 9 1 10 9 4 4 2
6 11 4 15 3 0 2
11 15 13 1 13 1 0 9 1 10 9 2
9 10 9 3 4 2 13 11 3 2
17 7 11 16 11 13 10 2 9 2 1 15 9 2 3 10 9 2
30 9 8 1 10 0 0 9 8 2 11 2 13 10 9 1 15 9 1 11 16 10 13 9 1 10 12 9 1 4 2
6 15 8 13 10 9 2
8 15 13 3 0 4 1 11 2
14 8 1 10 9 13 10 9 10 0 9 1 10 9 2
24 11 13 9 3 16 15 9 15 4 1 4 1 11 16 15 15 9 13 16 15 8 0 13 2
19 11 11 13 3 16 1 15 13 1 15 9 10 9 1 10 9 4 4 2
15 9 1 0 3 10 9 4 8 3 10 9 0 1 4 2
19 1 10 9 11 7 11 3 4 3 15 4 2 3 9 8 1 11 3 2
17 10 9 13 1 10 9 4 1 10 9 1 9 11 2 9 2 2
23 1 8 4 10 9 1 10 9 2 3 15 9 4 4 2 10 9 15 10 9 13 4 2
20 8 13 0 1 10 0 9 3 9 1 15 8 4 4 7 10 9 1 11 2
12 15 13 12 1 12 9 1 9 2 13 15 2
32 9 4 4 1 8 10 9 1 10 11 7 11 1 11 2 10 11 1 10 11 1 11 7 10 11 1 10 9 8 7 11 2
15 1 8 4 3 9 16 10 11 1 11 7 8 1 4 2
10 1 8 4 10 9 4 1 9 11 2
15 1 12 9 13 3 1 10 0 9 11 0 1 9 4 2
14 15 13 1 15 9 1 10 9 2 15 12 9 13 2
6 0 13 9 13 13 2
13 10 9 13 1 2 10 9 1 10 9 9 2 2
11 1 11 4 1 11 15 2 8 2 4 2
28 3 12 9 7 9 1 11 7 9 1 11 7 11 13 3 1 10 0 9 1 10 9 7 1 10 0 9 2
25 10 0 9 8 2 15 9 10 9 1 0 9 13 2 13 16 15 15 9 4 3 9 1 4 2
15 1 10 0 9 8 13 15 16 2 10 9 3 4 2 2
22 11 2 15 1 12 7 12 1 9 13 2 13 10 9 1 10 9 1 10 0 9 2
13 10 9 1 10 0 0 9 8 4 1 9 4 2
19 15 13 16 15 1 10 0 9 1 11 4 4 1 10 9 1 10 9 2
12 11 4 11 1 11 4 7 3 4 1 11 2
15 1 11 4 3 10 9 1 10 9 7 0 9 3 4 2
7 3 4 10 0 9 4 2
17 9 13 9 1 10 9 1 10 9 1 11 1 15 13 1 11 2
20 3 4 3 4 8 10 9 11 2 1 10 9 11 15 1 0 9 4 4 2
16 10 0 9 11 13 11 12 9 7 9 4 15 0 4 4 2
16 10 9 4 10 9 1 10 9 16 11 7 9 0 9 9 2
21 3 13 0 9 12 9 4 1 10 9 1 10 15 9 0 0 9 2 10 11 2
13 15 13 13 9 1 9 2 15 1 15 0 9 2
15 10 16 12 9 4 1 10 9 1 15 8 4 1 9 2
15 10 9 13 12 9 3 1 9 1 10 9 1 10 9 2
23 1 10 9 11 4 1 12 10 0 9 2 3 3 1 15 9 9 1 9 8 4 4 2
8 12 9 4 1 9 11 4 2
18 0 9 13 1 11 3 12 9 4 15 1 10 9 13 13 4 4 2
13 9 13 10 0 9 1 9 1 15 0 8 4 2
8 3 4 0 9 7 9 4 2
29 10 9 1 15 8 9 10 9 1 10 9 1 15 12 9 7 9 15 13 1 10 0 0 9 1 12 7 12 2
19 16 15 10 9 13 2 13 10 0 9 8 11 2 3 2 10 9 4 2
19 15 13 1 15 8 1 15 9 10 9 9 1 10 9 3 10 9 3 2
15 10 1 9 1 13 9 1 15 8 13 3 9 1 9 2
9 15 13 10 13 9 3 12 9 2
20 10 9 2 9 2 13 7 16 10 9 1 4 16 2 16 0 2 1 4 2
18 10 9 13 3 16 10 0 11 3 0 8 4 1 10 9 1 4 2
7 2 15 13 3 9 1 2
8 10 0 9 8 4 3 4 2
28 15 13 3 15 9 0 2 16 15 4 4 16 15 8 2 11 2 9 12 3 13 4 1 15 13 1 9 2
28 1 15 13 1 10 0 9 4 3 10 0 9 4 1 10 0 9 2 3 1 10 9 10 0 9 4 4 2
27 15 4 10 0 9 1 10 9 15 1 8 12 4 4 2 7 3 9 1 10 0 9 10 0 9 4 2
33 10 11 13 15 3 3 3 4 2 1 15 0 9 2 8 2 16 15 9 1 9 1 10 0 9 7 9 1 0 9 4 4 2
27 2 15 4 0 16 3 1 4 2 2 13 11 3 2 2 7 3 16 15 10 9 3 1 15 13 2 2
25 1 15 8 13 10 9 12 9 16 11 1 13 3 1 4 13 15 1 13 2 3 13 3 9 2
26 15 9 13 16 11 3 4 16 10 11 1 15 9 3 1 9 4 1 4 16 10 9 3 0 13 2
28 3 13 15 10 9 1 15 15 9 2 15 8 2 1 13 1 4 16 15 15 3 0 15 4 1 10 11 2
41 7 8 2 15 13 1 10 9 2 13 16 10 11 15 3 4 4 2 7 13 15 8 1 10 0 9 3 1 4 7 1 10 2 0 7 0 9 2 1 4 2
29 11 9 13 3 1 10 9 1 10 0 9 2 3 0 9 3 1 0 9 13 16 0 9 1 0 9 1 13 2
16 1 10 0 9 1 10 9 2 1 11 2 4 11 9 3 2
16 1 10 9 13 10 9 0 4 1 13 9 1 9 7 9 2
13 0 9 13 3 10 0 9 1 10 0 11 4 2
26 10 9 4 10 9 1 10 9 11 1 10 1 11 13 0 9 11 1 10 0 1 11 13 9 9 2
20 1 10 0 9 13 10 0 7 12 0 9 13 2 1 15 1 11 13 11 2
23 11 13 0 3 1 10 9 1 10 9 1 11 2 10 9 9 16 11 0 9 3 13 2
17 10 0 9 3 13 3 0 2 10 0 9 8 4 1 9 4 2
6 12 9 13 15 9 2
20 10 0 9 4 9 1 10 9 16 11 1 4 4 1 10 9 1 10 9 2
21 9 11 13 3 16 2 9 1 9 4 2 2 7 1 11 4 3 15 9 4 2
28 1 10 0 0 9 1 10 0 9 1 11 1 11 2 13 10 0 9 11 13 9 4 2 7 13 15 9 2
10 10 0 9 11 13 3 3 3 3 2
16 2 8 4 15 13 1 9 15 10 11 3 1 10 9 13 2
12 11 4 3 3 3 13 16 3 1 4 2 2
17 8 5 8 13 3 16 0 9 10 9 1 15 8 1 9 4 2
14 15 13 10 9 1 12 9 1 12 9 7 12 9 2
15 10 0 0 9 13 10 0 9 2 9 13 2 1 15 2
7 8 13 15 0 9 4 2
12 1 10 9 1 12 9 13 15 8 1 12 2
23 10 9 4 0 4 2 16 8 7 8 1 12 9 1 12 9 1 10 0 9 4 4 2
12 9 8 4 0 4 1 10 11 11 1 11 2
11 1 0 9 13 10 0 9 10 0 9 2
11 1 10 0 9 13 10 0 9 16 0 2
11 8 1 11 13 2 3 2 15 9 3 2
15 10 0 9 13 1 11 10 0 9 1 10 0 9 4 2
11 1 10 9 13 10 9 1 12 1 11 2
12 11 2 16 11 1 12 13 2 13 10 9 2
5 11 4 1 11 2
15 11 13 10 9 16 0 3 7 13 15 3 1 10 11 2
19 8 13 1 10 11 13 1 11 1 10 12 9 0 9 3 9 1 8 2
24 10 0 9 13 15 3 4 1 15 9 2 7 1 10 9 13 9 8 3 1 15 9 4 2
15 10 0 9 13 10 9 1 15 9 3 3 1 15 12 2
18 10 0 9 13 10 9 1 15 8 2 10 11 11 11 2 13 4 2
9 15 8 4 1 12 9 9 4 2
17 10 9 13 3 3 10 0 9 7 13 11 3 1 3 12 9 2
16 8 13 15 13 9 1 10 9 16 10 9 1 15 8 4 2
7 10 9 13 1 15 8 2
13 15 13 15 9 11 7 8 1 10 15 12 9 2
4 8 4 0 2
21 10 0 0 9 1 15 9 1 8 7 8 13 1 11 1 10 0 9 1 11 2
14 10 9 13 1 15 8 7 15 12 16 10 12 9 2
14 1 12 1 12 4 10 9 1 10 0 9 0 8 2
15 11 4 16 11 8 1 12 1 12 9 1 15 12 9 2
19 8 8 4 10 0 9 1 10 0 9 4 1 10 9 1 15 8 9 2
21 9 2 11 7 11 13 1 12 9 16 0 1 10 0 9 1 11 2 12 2 2
21 0 13 11 10 9 1 12 9 2 1 10 9 1 10 11 1 11 2 12 2 2
8 8 4 10 0 0 9 13 2
13 10 0 9 13 1 10 9 1 11 10 9 8 2
15 11 11 13 10 12 9 1 12 9 3 2 9 12 2 2
24 10 9 11 2 11 2 7 11 2 11 2 13 10 9 3 4 1 10 9 1 10 0 9 2
21 12 9 3 4 10 9 1 12 9 2 3 0 1 11 2 1 0 9 4 4 2
6 11 4 10 9 4 2
27 10 0 0 9 2 1 11 7 3 3 11 2 13 9 11 1 10 9 4 1 10 0 9 2 9 2 2
11 10 9 1 10 9 4 1 10 13 9 2
21 10 2 0 9 2 13 1 9 9 4 1 12 1 12 13 7 13 9 7 9 2
16 11 7 11 13 0 12 9 2 7 4 3 0 1 10 9 2
20 10 0 7 0 9 4 10 0 7 0 9 16 11 0 1 10 9 1 4 2
20 11 13 3 9 3 10 9 1 15 8 7 3 10 0 9 1 8 7 8 2
9 1 11 13 16 9 15 9 9 2
18 8 7 8 2 9 1 8 2 13 1 8 15 8 2 11 2 3 2
7 7 3 3 10 9 11 2
29 10 0 9 8 13 16 8 2 10 9 1 10 11 2 15 1 10 9 1 11 4 4 3 1 11 1 4 4 2
9 10 9 13 3 1 10 9 4 2
17 0 13 10 9 1 10 9 3 1 4 1 10 9 1 15 8 2
19 1 11 13 1 16 10 9 1 11 13 2 16 10 13 9 7 9 13 2
50 10 0 9 8 7 8 2 15 1 12 9 8 12 13 1 11 7 3 1 10 9 4 1 10 0 9 2 13 15 1 10 11 1 11 3 3 8 10 9 1 10 0 9 7 10 9 0 1 4 2
28 9 8 2 11 7 9 8 13 1 15 8 0 1 15 15 9 3 3 1 10 9 1 9 7 10 0 9 2
16 15 9 1 10 0 13 9 1 11 7 10 9 1 0 9 2
9 1 11 7 3 11 4 15 3 2
21 3 13 8 2 10 9 3 10 0 9 8 4 4 2 10 0 1 10 9 4 2
15 10 0 9 13 1 15 8 1 11 1 9 2 9 9 2
26 15 9 1 11 10 0 9 1 9 11 2 12 2 2 7 13 16 9 1 10 9 1 11 2 12 2
10 11 13 1 10 9 1 12 1 12 2
12 11 7 11 3 11 1 10 0 9 1 15 2
6 11 13 10 0 9 2
5 13 9 4 8 2
9 15 13 9 8 1 12 9 3 2
7 10 0 9 13 1 9 2
8 15 13 10 9 1 10 9 2
13 10 9 1 10 9 9 4 13 2 10 9 13 2
15 7 10 9 13 4 2 1 1 10 11 1 11 1 11 2
8 11 13 10 9 1 15 9 2
23 2 15 13 2 2 3 11 2 2 3 15 9 13 2 1 10 11 1 12 9 1 11 2
14 7 15 13 3 4 16 15 3 1 10 9 4 4 2
7 15 13 3 1 10 9 2
15 3 1 15 9 3 15 15 15 9 7 15 3 13 2 2
19 13 13 11 1 10 9 0 8 7 3 13 4 11 1 12 9 0 8 2
30 8 2 12 1 12 2 2 8 2 12 1 12 2 2 11 2 12 1 12 2 13 3 1 15 9 12 1 15 9 2
16 10 9 13 1 12 1 10 0 9 10 0 9 1 10 9 2
30 8 2 10 0 0 9 1 10 9 7 13 1 15 8 2 13 10 9 11 1 10 9 1 10 9 8 3 1 4 2
17 10 9 13 2 10 9 13 10 0 9 1 10 9 1 10 9 2
19 9 11 15 1 9 9 4 4 1 11 2 15 11 1 10 9 13 4 2
13 10 9 13 15 0 9 1 10 9 10 9 3 2
24 11 13 3 10 9 0 4 1 11 0 12 0 1 13 2 3 11 16 0 9 10 9 13 2
12 10 9 13 3 3 1 10 0 9 1 4 2
14 9 7 11 13 8 7 11 1 10 9 2 12 2 2
27 1 10 0 9 13 8 10 9 1 15 0 9 9 2 12 1 11 2 3 11 8 3 13 2 12 2 2
11 2 15 4 9 2 2 13 9 11 0 2
3 2 11 2
5 13 7 13 2 2
11 10 9 13 12 9 7 9 3 12 9 2
7 2 16 2 2 13 11 2
6 2 15 3 0 4 2
5 15 13 15 3 2
8 10 9 13 1 15 9 4 2
10 15 13 15 9 4 1 10 9 2 2
10 10 9 0 13 10 9 1 11 0 2
5 10 0 1 11 2
12 10 9 13 10 0 9 1 11 1 12 9 2
18 10 0 9 13 1 10 0 9 1 11 3 11 11 11 13 1 12 2
15 11 13 16 10 9 11 2 11 2 11 7 11 1 11 2
20 15 13 3 12 9 1 10 0 9 7 13 10 9 1 12 8 11 0 9 2
9 10 9 13 11 3 1 0 9 2
4 11 4 0 2
16 13 13 3 9 3 1 12 0 0 9 1 10 9 1 13 2
14 1 15 15 8 13 15 10 9 3 1 10 0 9 2
11 15 13 10 9 4 7 13 10 9 4 2
5 10 9 13 0 2
10 10 9 13 3 3 10 9 3 4 2
24 7 10 0 9 1 10 9 4 1 8 1 15 13 8 0 1 15 8 7 15 13 15 4 2
13 1 12 0 13 9 13 15 0 8 1 10 11 2
14 10 9 13 10 0 9 1 10 0 9 3 1 4 2
9 10 0 9 9 13 4 9 4 2
8 10 9 13 3 1 9 0 2
25 2 16 15 3 0 4 2 13 15 0 2 7 3 13 3 10 0 3 4 2 2 13 15 13 2
16 2 15 13 2 16 15 10 9 4 2 13 15 10 9 2 2
9 7 8 1 12 9 4 15 0 2
3 3 0 2
13 1 10 0 9 13 10 9 1 10 9 0 8 2
13 10 9 13 1 0 1 15 2 1 12 9 3 2
6 0 4 10 9 0 2
13 1 15 9 13 15 10 0 9 1 10 0 9 2
31 2 15 13 3 3 2 7 15 13 3 10 0 9 1 15 9 7 13 1 10 9 10 9 4 1 11 2 10 9 12 2
9 10 9 12 4 1 15 0 2 2
18 10 9 1 10 9 13 16 13 1 10 0 9 11 2 11 7 11 2
7 15 13 3 15 0 9 2
16 3 11 2 10 9 1 0 9 2 13 1 15 1 10 9 2
22 15 13 1 9 1 10 9 2 7 13 3 10 9 10 0 0 1 10 9 0 4 2
14 11 13 3 10 9 3 1 11 2 16 10 9 13 2
9 15 13 15 9 16 15 0 9 2
29 2 7 15 13 1 15 9 12 9 2 3 4 10 9 1 11 1 10 9 12 9 2 2 13 9 11 15 0 2
3 11 13 2
16 15 13 10 9 2 3 16 0 9 2 7 4 3 3 0 2
10 11 13 3 13 9 3 1 15 8 2
20 10 0 9 13 1 9 1 10 9 10 9 4 16 10 9 15 9 4 4 2
16 15 9 13 1 9 1 4 4 7 4 4 1 8 12 9 2
23 16 15 9 3 4 4 2 13 10 9 1 12 9 7 0 15 0 9 1 15 8 12 2
30 16 9 1 11 7 11 15 9 1 15 13 0 0 13 5 11 13 3 5 4 15 1 11 3 0 10 9 1 13 2
11 3 4 10 9 1 9 1 15 9 13 2
27 11 13 1 11 3 16 10 12 9 1 12 2 3 10 13 11 2 15 15 9 4 1 4 1 13 9 2
7 10 9 4 4 1 11 2
20 13 10 9 3 1 10 9 1 10 9 4 4 2 3 13 10 9 1 11 2
10 10 9 13 10 0 9 1 15 8 2
18 1 10 9 1 10 9 1 11 13 10 0 9 15 15 9 1 11 2
9 15 4 12 1 11 1 10 9 2
7 10 9 4 15 0 9 2
23 10 1 11 3 0 9 2 1 12 8 7 0 9 1 15 8 2 4 1 12 9 0 2
19 1 15 0 12 2 8 11 7 11 2 4 10 9 1 12 12 9 4 2
9 11 13 3 3 12 0 9 3 2
14 8 4 10 0 9 1 10 9 2 8 10 0 9 2
9 1 11 13 10 9 10 0 9 2
22 0 9 1 15 8 1 11 13 10 9 3 1 10 0 9 3 1 10 0 9 11 2
18 10 9 13 3 1 10 0 9 1 11 2 7 10 9 4 3 3 2
