2432 17
12 13 3 15 13 16 15 0 13 9 7 9 2
20 10 3 9 3 1 15 13 0 2 7 3 0 3 3 13 1 10 0 9 2
5 13 15 10 9 2
8 3 15 3 10 9 0 13 2
7 3 15 3 10 9 13 2
28 15 3 13 1 15 15 0 3 15 13 2 16 10 9 13 2 16 15 0 13 2 0 13 2 13 0 13 2
6 3 15 13 10 9 2
31 3 0 3 3 13 2 13 7 10 0 9 7 0 0 10 0 13 2 3 13 1 10 9 13 2 13 15 7 10 9 2
22 3 3 13 13 2 3 3 13 10 9 2 7 3 13 3 0 13 7 13 10 13 2
34 9 3 13 13 2 13 2 3 0 13 10 9 3 0 13 3 3 13 7 1 15 13 2 3 3 13 10 9 9 1 10 13 13 2
25 13 3 13 16 2 16 13 15 0 3 15 13 13 2 15 9 9 13 3 15 13 7 9 13 2
13 16 3 3 10 9 13 2 15 13 10 15 0 2
8 15 3 13 10 1 15 13 2
20 16 3 10 0 10 13 13 2 0 13 2 16 0 9 13 0 13 10 9 2
52 16 3 15 13 2 3 0 10 1 10 9 13 2 7 3 10 0 13 7 10 0 13 2 7 13 0 0 9 13 10 9 2 16 13 1 10 15 10 9 3 15 13 7 0 9 10 13 1 10 9 13 2
28 3 3 3 13 13 10 9 7 3 0 15 0 13 7 0 3 13 10 10 9 9 16 10 1 10 0 9 2
26 15 13 13 15 3 10 9 13 2 7 0 0 13 16 9 10 3 13 10 0 13 1 15 3 13 2
27 13 3 15 13 7 13 2 3 13 10 9 9 0 9 13 2 16 15 0 0 7 3 0 0 0 13 2
21 15 16 15 13 13 2 16 0 1 15 13 13 2 3 3 13 9 0 10 9 2
22 3 16 3 9 13 3 0 13 0 15 13 2 1 10 10 9 9 0 10 0 13 2
19 16 3 1 10 15 13 13 3 10 15 9 2 1 10 9 13 15 13 2
22 15 3 13 9 10 15 13 13 10 1 10 9 13 2 16 0 15 10 13 13 13 2
25 15 3 13 2 16 3 13 10 13 7 13 1 9 16 13 1 10 9 7 16 13 13 2 13 2
35 16 3 0 13 0 13 15 13 2 13 13 16 13 15 13 7 10 9 3 13 2 7 16 3 3 10 13 13 0 10 0 9 13 13 2
26 15 0 15 13 2 16 13 16 3 3 3 15 13 2 3 15 3 13 2 10 7 15 9 0 13 2
13 1 3 10 0 10 15 13 3 3 15 9 13 2
7 13 3 15 1 15 13 2
41 16 3 3 10 13 13 13 10 0 15 9 7 10 10 9 9 2 13 15 3 10 0 13 2 16 13 10 13 0 1 15 13 7 10 9 15 0 0 0 13 2
58 15 3 9 3 13 1 9 10 9 2 10 3 0 10 0 13 2 0 13 13 1 10 0 9 13 2 13 7 1 9 2 0 9 13 2 13 10 15 9 2 7 13 3 3 13 0 13 0 13 2 16 3 0 13 0 13 13 2
9 13 3 1 9 2 16 3 13 2
22 3 0 15 13 15 1 15 13 13 2 15 3 15 15 13 13 15 10 15 15 13 2
9 1 9 3 13 10 9 9 13 2
18 10 3 13 10 9 0 3 13 15 0 13 2 13 7 13 9 13 2
17 10 3 9 15 3 13 3 2 16 3 3 13 13 10 9 13 2
9 13 3 15 9 13 9 15 13 2
17 3 0 3 9 9 13 10 9 2 1 9 9 13 10 0 13 2
26 9 3 0 13 13 10 15 9 2 13 15 3 3 9 15 7 3 9 15 1 10 9 13 10 15 2
102 3 15 13 7 3 0 3 0 7 0 13 3 10 13 15 13 7 10 13 13 2 7 15 13 0 13 10 9 2 9 13 10 15 9 10 10 9 9 2 15 0 13 13 2 16 13 3 0 9 10 9 10 15 13 10 15 13 2 7 15 9 13 9 2 15 13 3 9 9 13 2 1 3 10 9 13 13 2 9 3 10 10 9 0 13 2 3 7 1 10 0 1 10 9 13 16 1 10 9 1 15 2
14 1 15 3 15 7 10 13 13 13 13 15 13 15 2
29 3 3 13 13 16 3 13 13 10 3 9 15 13 9 1 10 9 13 2 15 7 3 1 10 9 10 15 13 2
30 15 3 13 0 13 2 16 10 3 9 15 13 3 3 3 13 2 0 7 13 13 3 10 9 0 1 10 9 13 2
13 13 3 13 16 9 15 0 13 1 10 9 13 2
26 3 3 3 0 13 0 13 16 15 3 13 13 3 10 3 10 9 9 0 13 2 15 7 15 13 2
19 10 3 0 9 13 10 3 0 13 2 10 7 9 3 10 13 13 13 2
11 3 3 0 10 9 0 13 10 9 13 2
33 3 3 0 9 7 3 15 0 13 1 10 10 9 9 13 2 7 13 16 3 15 0 13 2 16 10 9 0 10 0 0 13 2
51 3 15 3 0 10 15 9 2 15 3 3 13 13 0 13 3 10 0 15 13 13 10 9 2 13 3 3 15 3 13 10 9 2 13 3 3 15 3 13 10 9 2 13 7 3 10 13 13 10 0 2
53 3 3 3 2 16 3 13 2 1 10 9 3 0 3 13 13 10 9 2 16 7 15 13 13 7 0 13 9 2 3 10 0 13 1 10 9 13 2 3 0 15 13 3 0 13 2 7 0 15 0 15 13 2
20 3 3 0 13 16 9 9 3 15 10 15 13 2 9 7 10 9 0 13 2
14 15 3 3 13 10 0 3 13 2 9 15 0 13 2
28 16 3 13 15 13 2 15 0 13 15 13 2 7 13 1 15 13 9 9 2 0 16 0 9 10 9 13 2
43 3 3 0 13 1 15 13 2 16 13 13 3 9 13 7 9 13 3 13 9 13 13 2 7 9 15 13 3 9 7 0 9 13 9 13 3 16 10 9 13 10 15 2
109 3 16 15 15 3 10 13 1 10 9 13 2 3 1 10 13 10 0 13 2 3 10 9 13 13 2 3 0 13 2 7 10 0 13 2 15 0 13 10 15 9 0 13 2 7 13 16 9 3 10 9 15 7 10 9 1 9 9 9 10 0 9 3 0 13 2 10 7 9 15 10 0 15 9 13 2 16 3 13 13 0 0 15 13 10 9 13 2 7 3 9 3 9 7 9 15 1 0 13 10 9 10 13 7 10 9 15 13 2
7 3 3 13 7 13 0 2
17 3 3 13 2 16 1 3 10 0 13 2 1 7 10 0 13 2
35 0 3 9 1 15 15 0 13 10 9 2 15 15 2 16 3 15 0 13 2 16 13 2 13 2 16 7 0 13 1 10 0 9 13 2
32 3 3 3 3 3 13 1 10 9 15 13 0 15 13 2 0 13 3 9 3 13 0 3 10 0 0 7 1 10 15 13 2
46 3 3 15 1 15 0 13 2 7 0 3 9 13 3 10 15 7 10 15 0 2 15 10 3 13 13 3 13 2 0 7 9 13 2 7 1 10 0 15 3 13 1 10 0 13 2
43 15 3 3 16 13 0 13 2 13 7 16 10 3 15 10 13 13 2 16 3 3 3 13 13 10 15 9 2 15 7 15 13 2 16 3 0 9 13 10 15 13 0 2
32 15 3 3 10 13 7 10 13 13 0 3 15 13 2 13 16 0 3 13 10 9 2 0 7 9 10 0 9 13 10 9 2
12 13 3 15 10 9 3 10 9 7 10 9 2
7 3 15 13 13 10 0 2
54 15 3 3 0 9 7 0 9 15 1 10 9 13 2 16 13 10 3 9 1 10 10 9 9 13 7 13 10 9 15 15 3 13 13 2 10 7 9 7 10 0 13 1 10 9 10 1 15 13 2 16 3 3 2
50 13 3 15 2 16 0 13 2 13 3 9 2 16 13 10 9 9 13 10 9 2 13 3 10 9 2 16 13 9 1 10 9 0 13 10 15 9 2 13 7 10 9 13 15 1 10 10 9 9 2
39 3 3 15 15 13 2 7 1 3 10 9 13 15 1 0 13 7 1 10 9 13 2 16 7 15 13 1 10 13 9 13 2 13 13 1 15 15 13 2
38 16 3 0 13 13 13 2 13 13 16 13 10 0 13 2 7 3 15 15 3 15 13 13 2 16 15 13 10 13 1 0 15 15 7 10 9 13 2
43 13 3 13 1 10 9 3 13 10 9 7 10 9 13 0 13 2 7 1 15 10 9 3 3 9 3 9 7 15 15 0 15 13 2 1 15 9 13 10 9 15 13 2
21 15 3 3 3 0 13 9 13 2 7 9 0 13 15 13 2 13 10 0 13 2
19 15 3 13 10 15 9 13 10 9 13 2 15 16 13 1 10 0 13 2
6 3 15 13 10 9 2
12 1 3 15 13 1 10 9 15 10 9 13 2
6 3 15 13 10 9 2
9 1 15 13 13 1 3 13 13 2
6 3 15 13 10 9 2
6 3 15 13 10 9 2
6 3 15 13 10 9 2
45 16 3 10 1 15 13 10 9 13 13 10 1 0 10 9 9 2 3 9 13 10 13 0 1 10 9 7 9 10 0 9 1 10 0 0 13 10 9 9 10 10 13 9 9 2
65 15 3 3 13 0 7 0 9 15 3 3 13 13 3 7 0 9 9 13 3 0 10 1 10 9 3 0 0 7 0 9 1 0 9 13 10 9 2 15 0 3 13 13 2 15 7 3 3 0 1 15 10 0 9 7 9 15 0 3 15 13 0 10 9 2
42 16 3 13 0 7 0 10 1 10 0 9 9 13 3 3 3 0 2 16 10 0 10 13 9 2 1 15 10 9 10 0 13 9 2 13 7 13 1 10 9 9 2
10 13 3 10 10 9 0 7 9 15 2
10 9 1 0 9 0 9 13 7 9 2
21 3 3 13 13 10 10 9 9 2 3 0 1 10 9 2 7 3 1 15 13 2
21 9 0 13 9 1 10 10 9 9 2 16 3 13 2 3 9 0 13 15 0 2
27 9 10 3 9 13 1 10 1 10 9 9 7 1 10 9 9 2 15 0 3 3 13 9 10 13 9 2
15 1 3 15 13 10 10 9 9 2 13 10 10 9 9 2
21 3 3 15 0 13 3 9 7 9 13 9 2 10 0 9 3 13 10 9 0 2
26 9 3 3 3 9 7 9 3 13 3 13 2 10 7 9 10 0 9 10 0 9 3 13 3 13 2
33 9 3 3 3 0 9 2 3 7 0 13 10 9 9 15 2 0 3 10 13 0 2 0 7 3 10 13 9 13 10 15 9 2
18 3 3 3 1 10 0 7 0 13 13 10 13 10 10 0 9 9 2
64 13 3 10 9 15 10 3 9 9 0 3 7 0 2 10 7 9 1 3 10 9 10 13 0 9 2 15 0 13 1 9 1 9 9 2 9 3 9 2 9 7 9 2 1 7 10 10 9 13 10 1 0 9 2 15 9 7 9 10 9 13 1 15 2
12 15 3 13 0 10 0 10 1 9 0 9 2
39 1 3 3 10 1 15 9 3 9 13 13 10 10 9 9 1 10 3 1 10 9 2 3 3 7 10 9 15 3 7 3 1 10 9 13 0 10 13 2
36 1 3 0 10 9 3 0 13 13 10 9 2 13 7 10 0 7 0 9 10 3 1 10 9 7 10 0 7 1 0 13 9 10 9 0 2
13 3 3 10 9 10 15 9 1 0 13 10 9 2
48 10 3 13 9 13 9 9 7 13 10 0 7 0 9 15 13 1 10 10 0 9 2 3 3 3 0 13 1 10 9 10 9 13 7 13 1 9 1 3 10 9 7 10 1 10 9 9 2
41 16 3 3 15 13 0 7 0 10 9 10 1 10 10 0 9 13 2 3 15 3 9 13 1 10 3 10 13 1 0 9 7 9 13 13 10 0 7 0 9 2
116 16 3 3 10 9 7 10 9 9 0 13 10 0 10 9 10 13 9 7 10 9 15 2 9 13 13 13 0 7 10 3 9 1 10 9 2 16 15 13 1 0 10 10 9 9 3 13 7 13 0 9 7 0 9 7 9 13 9 1 0 13 10 9 2 1 15 3 10 9 7 10 9 10 1 9 13 0 0 2 7 1 0 10 9 7 10 1 15 9 0 13 10 13 16 3 3 0 9 13 1 3 10 9 13 7 1 10 9 13 10 10 0 9 7 9 2
32 3 3 10 13 15 7 13 1 10 9 10 9 3 15 13 2 1 7 15 3 10 15 10 1 15 13 10 10 3 9 9 2
11 0 3 3 0 15 1 0 10 9 13 2
5 15 13 3 13 2
45 3 3 3 15 13 10 13 1 10 1 9 9 3 13 10 0 0 15 13 2 16 3 16 15 0 7 0 9 13 13 10 9 13 13 3 9 13 10 9 0 10 9 7 9 2
48 16 3 15 3 3 13 7 0 3 13 10 9 10 3 9 7 10 10 9 9 3 3 13 10 0 15 2 3 3 13 0 15 13 16 3 3 0 15 10 9 13 3 7 0 10 13 13 2
18 9 3 3 13 1 9 10 0 0 2 9 7 7 9 0 13 0 2
18 3 3 0 15 0 13 10 1 9 9 1 10 10 0 9 7 9 2
13 13 3 0 9 10 9 10 0 9 1 9 9 2
23 15 3 13 0 3 10 1 15 9 13 2 13 7 1 10 0 7 0 1 10 12 9 2
24 3 3 0 3 13 3 7 3 13 10 1 10 9 7 0 9 1 15 13 13 13 1 9 2
12 0 3 10 9 0 13 10 1 9 10 9 2
25 3 0 0 10 10 9 9 3 2 16 3 10 9 9 13 0 10 10 0 9 9 13 7 9 2
22 16 3 10 1 15 13 13 9 2 3 3 3 0 10 0 9 9 13 1 10 13 2
66 9 3 3 13 1 3 10 1 9 9 9 0 2 1 7 10 1 9 9 0 2 1 15 9 3 10 1 9 13 9 1 9 10 9 13 7 0 9 10 1 10 9 9 9 13 10 1 10 9 9 13 9 2 9 7 1 9 13 0 10 9 13 1 10 9 2
31 1 15 13 9 9 7 9 13 9 3 13 3 3 10 9 0 7 13 0 9 10 9 13 1 10 3 9 1 10 0 2
41 13 3 0 0 10 9 1 3 10 9 7 10 1 10 9 9 1 15 13 9 2 3 9 2 3 7 9 10 1 3 10 9 7 10 9 13 10 10 9 9 2
103 1 3 0 9 9 1 10 1 10 9 9 9 7 10 1 15 9 13 9 2 0 0 9 10 10 9 9 10 3 1 9 13 7 13 1 10 9 2 9 9 3 7 9 1 15 13 2 10 7 1 10 9 9 0 9 3 13 2 3 0 1 10 0 9 10 9 13 2 3 16 1 0 2 1 7 10 0 16 1 0 3 7 13 15 13 2 9 13 0 10 1 10 9 9 1 10 1 10 9 7 9 9 2
26 13 3 3 0 0 7 13 10 10 9 13 1 15 1 9 1 15 13 13 10 3 13 10 9 9 2
14 0 3 15 13 7 0 0 10 1 10 9 13 9 2
7 13 3 15 9 7 9 2
35 9 3 3 3 0 0 9 10 3 13 9 9 1 9 13 7 3 1 10 9 7 10 0 9 10 9 13 1 10 13 9 3 13 13 2
28 13 3 15 10 3 9 7 10 9 10 13 2 16 3 10 9 13 1 0 10 10 9 9 0 2 3 13 2
12 10 3 0 9 7 10 9 1 15 13 13 2
17 0 3 7 3 0 9 7 9 0 13 1 9 13 9 10 9 2
30 9 3 2 1 0 9 9 1 9 13 2 0 13 10 9 15 2 13 7 3 9 13 13 9 3 7 9 1 9 2
24 10 3 13 9 3 0 13 10 9 7 10 15 9 2 13 0 10 9 2 15 13 9 0 2
19 3 10 3 13 2 10 7 13 10 9 10 0 9 10 9 13 10 9 2
9 10 3 9 3 3 13 10 13 2
13 3 3 13 3 13 15 1 10 13 10 13 9 2
16 16 3 1 15 13 2 13 15 13 10 9 2 16 3 13 2
26 13 3 10 3 0 1 0 10 9 13 2 3 13 1 10 13 10 13 2 9 7 13 0 16 0 2
43 15 13 1 10 9 2 10 9 13 1 10 9 7 13 0 1 10 1 15 9 13 2 13 1 10 1 15 9 2 1 0 0 3 13 2 13 1 10 0 10 15 9 2
11 10 3 9 7 10 9 3 10 9 13 2
32 16 3 13 10 13 9 2 13 10 10 9 13 1 10 9 2 1 9 1 10 9 15 3 13 1 10 9 1 0 0 9 2
48 10 3 13 10 9 3 13 1 10 9 1 0 0 7 9 13 10 13 3 13 3 7 3 10 9 2 16 10 9 2 16 3 13 1 10 10 9 9 2 3 0 3 13 9 15 13 9 2
19 15 1 10 0 9 3 0 13 10 3 13 0 13 9 7 1 10 9 2
74 13 3 10 9 2 16 13 10 9 7 10 9 1 10 9 2 15 1 15 13 7 13 3 15 2 10 7 9 13 3 10 9 7 10 9 0 13 10 0 9 2 13 3 7 1 10 9 3 2 13 9 1 15 2 13 0 9 13 1 10 9 15 2 16 15 13 13 1 10 9 1 10 9 2
26 13 3 10 9 10 13 7 13 10 0 0 9 13 7 0 13 9 16 1 10 0 10 10 9 13 2
17 1 3 10 10 15 9 9 3 15 13 1 10 9 1 10 9 2
30 13 3 10 13 3 7 13 0 10 0 7 0 10 9 2 13 1 15 9 0 0 2 3 3 10 1 10 9 13 2
31 9 3 13 15 0 7 10 9 0 13 9 10 3 10 0 13 9 2 15 7 13 1 10 9 9 1 0 13 10 0 2
16 9 3 0 3 9 13 1 10 13 0 13 10 9 10 9 2
42 10 3 0 0 10 0 9 1 10 0 13 9 2 16 9 13 2 3 9 13 13 10 10 0 13 3 0 1 10 9 2 7 3 10 9 9 2 0 13 10 9 2
69 3 9 13 3 15 15 2 13 3 10 9 3 0 10 1 10 9 2 7 3 10 9 9 0 9 13 2 3 7 10 9 0 0 13 10 1 10 0 7 0 9 2 13 2 16 9 3 13 2 16 3 0 7 0 9 15 13 2 9 0 13 7 9 10 10 9 9 13 2
18 16 3 3 1 15 13 10 9 2 3 13 9 10 9 2 0 13 2
22 13 3 13 15 10 9 13 1 0 9 10 9 13 1 10 0 3 13 10 0 9 2
17 13 3 10 1 10 9 10 10 9 9 13 10 1 10 9 13 2
40 10 3 0 13 3 1 10 13 9 7 13 0 9 2 1 7 10 3 13 1 10 3 13 10 9 3 1 0 0 9 0 7 0 13 10 9 2 13 13 2
25 13 3 10 9 1 10 9 2 13 10 0 10 0 9 9 9 13 2 13 13 7 13 1 9 2
22 10 3 9 10 3 10 9 9 3 13 10 9 13 2 10 3 13 2 10 7 13 2
10 10 3 9 13 7 15 10 9 13 2
19 9 3 10 3 9 15 13 2 13 15 3 2 3 7 3 13 10 9 2
23 15 3 10 3 0 9 1 9 13 2 10 7 0 9 1 10 9 13 3 13 10 9 2
31 1 3 10 9 0 9 13 3 13 10 13 1 10 10 0 10 10 9 13 3 13 1 10 9 2 13 1 10 9 9 2
15 3 1 15 13 1 10 9 13 10 9 1 10 13 9 2
20 13 3 1 0 9 1 10 0 9 13 13 3 15 10 9 10 1 10 9 2
17 10 3 9 10 9 9 9 7 3 13 10 9 13 1 10 9 2
45 13 3 3 3 13 10 0 7 13 3 3 0 2 3 7 0 13 10 9 15 2 10 3 9 10 0 13 7 10 9 2 10 3 0 13 1 0 2 13 13 10 9 10 9 2
15 15 3 13 15 2 9 13 13 13 7 0 13 10 9 2
20 13 3 10 9 13 1 9 2 3 1 10 9 13 15 3 10 10 9 9 2
18 1 0 3 9 13 13 10 0 7 13 10 0 16 1 10 9 0 2
12 9 3 3 13 10 0 13 3 1 10 9 2
20 10 3 9 13 15 1 10 0 9 2 13 10 9 13 1 9 1 10 9 2
23 10 3 1 9 9 13 9 10 9 10 13 7 13 0 13 3 13 2 7 13 10 9 2
17 13 3 10 9 1 9 13 10 9 2 1 10 9 10 9 13 2
20 13 3 10 0 0 3 15 13 2 10 7 0 13 13 3 1 10 13 9 2
30 13 3 10 9 0 7 13 10 9 2 0 13 3 13 10 3 10 9 7 10 10 13 15 9 2 15 13 10 0 2
10 10 3 0 13 15 13 13 10 9 2
52 10 3 3 0 9 1 10 9 9 1 9 0 3 1 15 7 1 15 13 10 9 2 15 0 13 9 13 10 0 9 2 1 15 13 10 9 2 13 3 10 9 10 15 9 13 1 10 1 10 9 9 2
48 10 3 3 7 3 13 15 10 9 9 10 1 10 0 13 9 7 3 3 7 3 13 10 1 10 9 10 3 13 13 9 2 9 13 13 13 10 13 3 10 0 15 10 3 9 3 13 2
19 3 3 13 13 3 1 10 3 2 16 3 13 10 9 1 10 0 9 2
33 15 3 13 1 10 13 9 15 2 1 15 13 3 13 1 15 0 3 3 7 3 13 1 15 13 10 9 2 1 15 13 3 2
8 15 3 3 1 9 3 13 2
17 15 13 0 1 10 9 10 13 9 7 9 1 10 1 9 9 2
32 15 13 1 10 15 9 10 0 9 9 1 10 9 7 15 10 9 10 9 2 1 7 10 13 10 1 10 1 9 9 9 2
29 15 3 1 10 15 9 1 10 9 10 0 13 13 9 2 1 15 3 10 9 13 10 0 9 7 10 0 9 2
21 3 3 13 1 15 13 2 13 7 3 13 1 10 9 10 13 1 15 13 9 2
23 3 1 0 13 1 10 0 10 13 13 13 10 9 10 9 10 10 0 9 9 7 9 2
37 15 3 10 9 0 13 10 9 2 15 3 13 3 13 10 3 13 0 2 10 7 13 1 10 0 9 0 7 0 1 10 13 13 13 10 9 2
16 0 7 0 13 13 1 10 0 13 9 9 7 9 1 9 2
27 7 3 0 15 9 13 9 3 9 0 3 0 9 3 0 9 7 9 0 10 1 10 13 9 13 0 2
25 15 3 10 9 1 15 10 9 3 0 3 13 10 9 2 0 3 10 9 2 0 7 10 9 2
26 3 3 10 13 3 13 10 0 10 9 9 7 9 3 3 1 10 13 9 16 1 15 0 10 9 2
18 0 3 3 13 10 9 3 13 2 13 1 10 9 7 10 9 15 2
9 13 3 15 13 15 0 10 13 2
31 1 3 10 9 7 10 0 9 9 3 0 13 10 9 13 3 2 3 2 3 2 10 7 9 0 2 9 7 3 15 2
15 1 3 3 10 0 9 10 15 9 3 3 3 15 13 2
21 3 3 0 13 13 10 0 9 7 9 7 13 10 0 10 0 7 13 10 0 2
49 16 3 10 10 9 9 13 15 2 13 13 0 10 15 7 3 3 13 7 13 10 0 9 10 0 2 16 10 9 13 15 2 3 7 13 7 13 3 10 0 2 16 10 10 9 9 15 13 2
23 16 3 9 10 9 13 13 10 0 2 3 1 9 13 10 9 10 13 15 0 13 9 2
36 3 3 10 0 13 7 10 0 13 0 2 7 3 10 15 13 2 3 7 13 0 2 16 10 1 9 13 3 13 3 0 7 13 3 13 2
17 13 3 10 13 15 10 13 0 10 13 9 7 9 1 10 9 2
14 16 3 13 0 10 3 1 15 13 13 1 15 13 2
38 10 3 9 13 3 10 9 7 10 0 9 13 13 10 9 13 10 3 9 7 10 9 2 13 7 10 9 1 9 1 10 9 3 13 1 10 9 2
46 15 3 13 10 3 9 13 1 10 13 9 3 1 13 10 13 16 3 0 3 10 9 7 10 9 13 13 9 1 10 9 2 7 3 10 9 0 13 10 13 1 10 10 9 9 2
19 15 3 2 16 15 13 2 10 0 13 9 0 7 9 3 13 10 3 2
21 15 3 13 7 13 13 2 15 13 3 3 13 10 9 7 9 13 10 9 13 2
7 15 3 13 15 3 13 2
16 3 9 3 10 9 13 10 0 0 7 10 1 10 13 9 2
6 13 3 15 3 0 2
38 3 3 13 10 9 7 9 10 0 2 7 10 9 13 10 9 1 9 2 16 3 15 13 2 7 10 9 2 1 9 13 10 10 9 7 9 9 2
25 9 3 3 1 0 3 15 10 9 13 15 13 2 3 3 3 9 2 16 1 0 13 10 9 2
34 15 3 16 10 13 13 9 1 10 9 2 13 1 10 9 13 13 3 10 3 9 1 0 9 13 1 9 10 13 1 10 13 9 2
37 13 3 1 10 9 1 10 9 10 1 10 9 7 10 9 9 2 13 0 9 9 7 9 9 10 3 9 0 13 7 10 9 0 1 10 9 2
18 13 3 1 9 10 0 9 9 0 1 10 0 2 10 1 9 13 2
10 15 0 1 0 0 2 9 7 0 2
18 15 13 1 3 10 9 10 0 13 9 13 10 9 1 7 10 9 2
37 10 3 9 13 10 9 7 9 10 9 2 3 7 10 9 7 10 9 10 0 9 2 1 0 13 15 0 13 10 10 9 7 10 10 9 9 2
11 10 3 9 13 2 3 3 1 10 9 2
25 13 3 10 9 13 16 3 13 10 0 1 10 3 1 10 1 15 13 9 0 9 13 10 0 2
17 3 13 10 9 0 1 0 10 9 15 13 9 3 13 10 9 2
34 13 3 9 1 15 10 3 0 1 9 13 10 9 9 2 9 7 13 9 15 12 2 0 3 9 3 16 0 7 0 13 10 9 2
35 10 3 9 9 13 15 1 10 9 9 7 13 3 15 1 10 13 10 9 3 13 10 9 10 1 15 9 2 13 7 13 1 10 9 2
23 0 3 3 0 15 13 7 0 9 13 10 0 9 1 3 10 1 9 7 10 3 9 2
56 13 3 10 9 1 10 9 2 3 13 10 9 7 13 10 1 9 9 2 0 3 0 13 13 10 9 10 9 2 7 0 0 9 2 13 3 3 13 10 9 15 13 10 9 2 3 7 3 13 3 13 10 9 10 0 2
39 10 3 9 13 10 3 9 0 15 13 2 10 7 9 0 13 1 10 1 10 9 13 0 13 9 2 1 15 13 13 10 0 7 13 10 1 10 9 2
25 3 3 13 1 10 0 9 0 3 9 7 9 2 3 7 0 15 9 2 0 1 10 9 13 2
37 13 3 10 10 9 9 0 13 1 10 9 7 0 3 10 15 9 1 15 13 10 3 9 7 10 9 2 9 13 13 15 10 9 1 10 9 2
14 10 3 9 10 3 1 10 9 13 9 10 9 13 2
18 10 3 1 15 13 9 9 7 9 9 13 1 10 9 1 10 9 2
18 13 3 10 10 9 9 7 10 1 10 9 9 13 0 13 10 9 2
20 3 3 10 3 15 9 10 9 13 2 13 7 0 10 9 1 15 9 13 2
14 3 13 1 0 9 1 10 9 13 1 9 10 9 2
22 13 3 10 10 9 9 2 7 13 0 9 2 13 0 10 13 10 9 1 10 13 2
16 10 3 9 13 10 0 13 1 10 9 2 13 13 10 13 2
19 13 3 15 3 10 3 1 10 10 9 9 13 2 10 7 1 10 9 2
15 3 10 10 9 9 3 3 7 3 3 13 10 9 9 2
18 10 3 9 1 15 9 13 10 13 10 9 7 13 10 3 1 9 2
22 3 3 3 0 13 10 0 13 3 0 3 10 0 13 2 3 7 0 10 0 13 2
27 9 3 13 10 0 0 3 13 10 9 2 10 3 15 13 2 10 7 0 13 7 13 13 1 10 9 2
21 1 3 15 13 10 3 9 0 13 1 10 9 2 10 7 9 0 13 10 9 2
43 16 3 3 13 10 9 16 1 9 2 13 10 9 10 9 1 0 9 10 9 10 3 9 1 10 1 10 9 9 13 2 0 7 13 1 10 1 9 13 9 10 9 2
51 10 3 1 10 9 1 0 10 9 10 9 13 7 10 3 1 15 9 13 1 10 1 10 13 1 10 9 9 2 10 7 1 15 13 2 9 13 10 3 9 7 10 13 7 13 13 1 10 13 9 2
20 10 3 1 10 9 7 10 9 9 9 13 2 13 10 0 10 9 1 9 2
25 0 3 3 3 9 1 10 15 13 2 15 0 9 13 13 1 15 1 10 1 15 10 9 13 2
23 10 3 1 10 9 10 13 9 7 9 13 10 9 13 1 10 9 1 9 10 0 9 2
13 1 15 13 10 9 1 0 13 7 13 10 9 2
19 1 3 15 13 10 9 7 9 10 9 16 3 13 1 10 13 10 9 2
24 15 3 3 9 3 13 2 16 3 0 9 7 9 13 9 10 0 7 0 15 13 10 9 2
87 1 3 15 13 10 13 9 10 3 9 1 3 10 9 7 10 9 3 13 1 10 0 13 1 15 9 2 10 7 0 9 13 0 1 9 13 2 13 10 3 9 1 0 10 9 13 7 10 0 9 0 13 1 9 1 10 9 2 13 10 0 9 13 3 13 10 9 10 0 13 7 13 10 9 15 13 2 7 3 13 13 2 16 3 15 13 2
15 10 3 9 13 1 10 9 2 16 13 10 1 10 9 2
23 0 3 1 9 13 13 10 0 7 0 3 15 13 2 10 7 0 16 1 10 9 13 2
25 13 3 15 13 10 1 10 9 10 9 2 13 10 9 10 13 9 2 3 0 9 13 10 0 2
18 3 0 3 9 13 1 10 13 2 15 0 13 16 13 1 0 9 2
54 10 3 9 13 7 13 3 1 10 9 1 10 9 7 13 16 10 9 10 9 3 13 2 0 3 7 1 10 0 13 1 10 9 2 13 13 10 10 9 9 2 3 0 1 15 13 3 10 9 1 10 13 9 2
14 3 13 0 10 9 1 10 1 9 10 9 13 15 2
17 1 0 3 9 13 10 9 9 13 10 13 0 10 9 10 9 2
20 15 3 13 1 10 9 7 10 0 9 10 13 13 0 13 10 10 9 9 2
16 13 3 9 0 10 3 0 13 15 2 15 7 1 9 13 2
13 10 3 9 10 3 0 13 9 7 10 9 0 2
51 13 3 10 9 2 3 1 10 1 10 9 9 7 1 10 9 0 10 9 15 13 2 13 9 10 9 7 13 13 0 9 1 9 1 10 13 9 2 13 1 9 9 1 10 9 2 13 10 0 9 2
15 13 3 9 9 13 10 9 13 10 0 13 3 10 9 2
28 10 3 9 10 9 13 13 10 13 7 10 9 10 10 1 10 9 1 0 13 1 15 0 13 1 10 9 2
23 15 3 3 15 13 2 13 13 10 9 7 0 3 9 2 0 7 3 0 13 9 0 2
13 15 3 3 1 10 0 9 13 1 9 15 13 2
12 10 3 9 3 10 9 13 13 15 10 9 2
39 1 3 10 3 9 2 13 15 3 10 9 2 0 3 9 13 10 0 10 9 2 13 10 0 9 2 3 7 0 13 10 0 2 13 10 10 9 9 2
48 3 13 3 7 3 1 0 10 9 9 13 10 9 1 10 13 9 2 3 7 10 3 9 13 3 1 10 0 9 2 10 7 9 1 9 0 13 2 13 1 10 13 10 9 1 10 9 2
37 3 3 15 10 9 3 0 15 13 13 9 1 0 10 13 9 1 10 3 15 13 10 9 2 3 3 3 7 1 0 9 0 13 1 9 9 2
32 10 3 9 1 9 0 13 10 1 10 9 9 1 10 15 3 10 1 10 9 13 0 9 2 0 15 13 15 10 9 9 2
15 1 15 3 3 13 15 3 10 0 7 0 10 9 9 2
48 3 3 0 0 9 13 2 7 3 9 3 7 9 3 13 10 9 2 3 3 0 1 9 13 3 3 13 16 3 16 13 10 9 2 3 13 9 13 10 1 9 13 10 1 9 9 0 2
21 9 3 3 15 13 1 10 9 10 3 1 15 13 7 1 10 0 15 10 9 2
50 16 3 10 0 13 13 1 10 9 10 9 2 3 0 0 15 13 9 2 7 3 3 0 9 7 9 3 9 2 7 1 9 7 9 3 7 9 7 9 13 9 7 9 1 15 3 13 10 9 2
60 1 15 3 9 10 9 1 10 9 13 15 2 7 0 9 0 1 10 9 13 2 16 13 13 10 9 0 2 15 9 13 3 1 15 13 10 10 0 9 9 2 16 16 3 15 13 13 2 0 16 1 10 9 1 9 3 13 10 9 2
31 3 3 3 15 3 0 13 10 9 2 13 1 10 10 9 9 2 10 7 10 9 13 13 1 10 9 13 10 9 15 2
54 13 1 10 9 1 10 9 10 9 10 15 13 9 10 1 15 10 9 9 2 0 7 1 15 13 10 9 2 3 0 13 1 15 13 10 9 7 3 13 13 15 13 13 3 7 13 10 9 1 10 10 9 9 2
30 13 3 15 2 1 10 13 10 9 13 7 0 9 1 0 10 9 1 9 13 13 1 10 9 1 10 9 10 9 2
50 10 3 1 10 0 9 13 10 9 9 9 0 9 0 2 13 10 9 2 16 13 10 9 2 0 16 1 10 9 2 15 13 1 9 0 13 1 10 9 2 13 10 13 1 10 9 13 10 9 2
27 13 3 15 9 3 1 10 10 9 9 2 13 10 9 0 10 13 13 10 13 9 7 13 1 10 9 2
23 10 3 10 9 9 9 2 13 1 10 9 10 13 13 9 10 9 13 2 9 0 13 2
12 15 13 9 1 10 9 13 10 1 10 9 2
28 9 3 13 10 3 9 1 9 13 1 10 9 2 10 7 9 0 13 7 13 13 15 9 13 15 10 0 2
19 10 3 9 10 3 9 7 10 9 10 0 0 13 3 1 10 9 13 2
28 1 3 0 3 9 2 3 0 13 7 0 10 1 10 9 9 2 1 0 0 9 1 10 0 9 3 13 2
30 13 3 10 10 9 9 13 1 10 9 3 13 2 13 13 10 3 9 7 10 0 9 10 0 2 13 0 9 13 2
35 13 3 1 10 10 9 9 13 10 0 1 9 7 9 13 10 9 7 10 3 0 13 10 9 2 15 7 1 10 13 3 7 3 13 2
21 9 1 9 0 13 2 9 3 9 9 2 1 7 10 9 0 9 13 10 9 2
28 15 15 3 1 10 9 9 13 2 13 7 15 9 0 9 13 2 9 3 9 9 2 10 7 9 0 9 2
21 10 3 9 10 9 13 0 7 13 1 10 9 1 10 0 3 10 9 0 9 2
26 1 3 10 9 0 13 0 0 9 13 2 13 9 1 10 9 2 16 10 0 13 0 10 0 9 2
45 1 3 15 10 9 13 9 2 15 1 10 9 10 9 13 10 9 1 10 1 10 9 9 13 1 10 9 10 0 9 3 3 1 9 2 3 7 13 10 1 10 9 13 9 2
39 16 3 10 9 10 9 13 10 9 3 13 10 9 2 16 3 0 13 15 2 3 13 2 16 7 1 3 2 1 0 10 9 1 0 0 13 10 9 2
32 15 10 3 13 10 1 9 9 13 10 10 9 9 2 10 7 13 10 1 10 9 13 9 1 10 9 13 10 9 10 9 2
11 15 3 3 15 13 9 9 13 1 9 2
27 10 3 9 9 16 0 13 10 9 10 10 0 9 13 2 13 10 0 9 10 9 15 13 1 10 9 2
40 13 3 10 9 1 9 7 9 13 9 0 7 0 2 13 10 9 10 9 2 7 0 13 0 10 0 2 3 9 13 10 9 2 7 3 1 9 0 0 2
26 1 3 10 13 13 13 10 9 1 10 0 9 2 1 0 3 13 10 9 2 13 10 10 9 9 2
13 3 3 3 3 13 10 0 13 10 0 13 3 2
8 0 3 9 13 10 9 13 2
21 3 3 0 3 10 0 13 9 0 13 2 1 15 13 0 3 10 10 9 9 2
11 9 3 3 7 3 0 1 10 9 13 2
33 10 3 0 9 10 9 13 3 10 9 16 1 9 2 1 7 10 13 13 10 13 1 10 13 9 13 7 13 10 10 9 9 2
21 13 3 10 13 2 10 3 1 9 2 10 7 1 9 13 3 13 13 10 9 2
18 10 3 9 3 13 10 1 9 9 2 3 13 10 9 1 10 9 2
28 3 3 3 13 10 9 10 3 9 13 9 3 15 3 13 1 7 10 1 10 9 9 9 9 1 9 13 2
69 1 3 10 9 9 2 10 10 9 9 10 13 1 10 0 9 2 13 1 9 2 13 1 10 0 9 13 10 0 1 10 9 1 10 1 10 9 9 2 7 13 13 15 1 15 10 0 1 10 9 7 10 9 10 9 2 13 15 3 13 1 0 10 9 3 1 0 13 2
34 1 3 15 10 9 10 3 9 13 10 13 9 13 1 10 9 2 3 3 0 7 3 1 9 13 2 13 9 7 15 10 0 9 2
28 9 3 3 0 3 1 10 9 13 1 9 1 15 9 7 0 13 10 9 2 3 13 1 10 13 9 13 2
14 9 3 3 10 9 13 7 10 1 9 9 3 13 2
42 10 3 1 10 9 9 10 9 1 3 10 3 9 15 0 13 9 2 3 7 13 10 13 9 9 9 7 9 9 13 1 10 9 1 10 10 10 9 9 3 13 2
12 10 3 9 13 10 9 1 0 10 9 13 2
19 10 3 9 9 0 0 1 15 13 2 3 13 9 7 13 10 9 13 2
8 1 3 15 13 9 13 13 2
41 10 3 3 9 9 9 10 9 10 9 1 9 13 7 13 3 13 10 10 9 9 2 13 10 0 9 13 10 13 2 0 13 1 10 15 2 13 0 9 13 2
27 10 3 9 13 10 0 10 3 3 13 2 10 3 13 2 10 7 0 0 13 10 15 2 13 15 13 2
17 3 13 10 3 15 13 2 10 7 10 9 9 1 0 0 13 2
25 3 9 3 15 3 10 9 13 7 13 13 3 10 9 2 10 7 0 10 9 13 1 0 13 2
18 13 3 1 9 13 10 0 7 0 3 0 9 13 2 0 7 13 2
12 10 3 0 10 9 13 1 10 9 13 9 2
26 1 3 15 10 9 0 13 0 13 10 9 2 13 0 1 10 13 0 9 7 10 1 9 13 9 2
25 10 3 0 9 1 10 1 15 9 15 13 0 9 2 7 1 0 3 10 13 9 13 10 9 2
24 3 13 2 16 13 2 1 10 13 0 13 9 3 0 7 0 0 9 0 7 13 1 9 2
28 3 13 13 9 13 10 9 2 13 7 10 9 13 1 9 1 10 3 10 0 9 1 15 15 13 10 9 2
19 9 3 0 7 0 9 0 13 9 13 2 3 7 1 9 10 0 13 2
35 13 3 10 3 9 9 1 10 9 13 7 10 9 3 13 2 16 10 9 3 1 9 2 7 1 15 15 7 10 0 9 10 9 13 2
7 10 3 9 0 15 13 2
33 13 3 16 0 13 10 9 7 0 10 1 10 9 9 0 10 3 1 15 13 2 3 0 3 13 13 2 7 13 7 13 13 2
25 13 3 10 3 1 10 13 2 10 7 1 10 13 2 0 13 10 13 9 1 10 0 13 9 2
22 3 13 1 10 0 9 10 0 9 13 10 0 9 2 15 13 13 2 1 9 9 2
8 10 3 9 0 0 13 9 2
14 0 3 3 13 9 7 0 9 7 10 9 1 9 2
9 10 3 0 3 0 0 3 13 2
11 9 3 13 1 10 1 10 0 9 9 2
16 10 3 9 10 3 0 3 10 0 13 1 10 1 9 9 2
15 10 3 3 9 15 13 1 0 9 1 10 10 9 9 2
42 1 15 3 0 3 15 13 7 13 1 10 9 2 7 3 13 13 10 10 9 9 7 10 10 9 0 9 7 9 2 13 1 3 10 10 9 7 10 10 9 9 2
26 10 3 9 13 16 10 3 9 13 13 0 2 10 7 0 13 2 3 13 13 10 9 0 7 0 2
24 10 3 3 0 0 13 2 1 15 13 10 9 9 9 7 9 9 2 0 1 9 0 13 2
33 15 3 0 0 1 0 9 13 10 3 10 0 2 10 7 10 0 9 13 2 3 1 0 9 0 10 9 0 10 3 13 9 2
13 10 3 9 3 13 10 9 10 9 1 15 13 2
10 15 13 13 0 10 0 9 10 9 2
17 1 3 15 13 10 0 2 9 13 1 15 10 10 0 9 9 2
27 15 3 3 13 10 0 9 2 10 9 13 2 1 0 13 9 2 16 13 1 0 10 9 10 1 15 2
46 3 13 0 1 10 13 9 2 10 3 0 13 9 10 9 9 2 15 10 3 1 10 9 9 13 0 2 10 3 1 10 9 0 2 10 7 0 0 7 0 2 3 7 3 0 2
47 10 3 10 9 9 1 10 0 9 13 10 0 1 9 7 13 15 16 13 3 10 9 1 9 13 10 9 2 13 7 1 10 0 9 13 7 10 9 2 3 15 13 13 1 10 9 2
20 3 3 0 13 10 13 1 10 13 10 13 1 10 13 2 3 13 7 3 2
45 13 3 10 10 0 9 10 9 7 1 15 13 10 3 9 9 10 15 9 1 0 13 9 2 1 10 9 13 10 0 9 2 3 13 10 0 2 0 13 0 10 9 10 0 2
16 10 3 0 0 10 0 9 13 2 1 0 13 1 10 9 2
29 13 3 10 9 10 3 0 9 2 13 9 7 9 10 3 13 1 10 9 2 9 10 1 10 9 13 10 9 2
13 10 3 0 13 10 9 9 10 1 10 9 13 2
17 15 3 1 0 10 9 13 10 9 13 0 9 1 10 9 0 2
24 10 3 9 13 1 0 13 10 9 7 13 10 9 1 0 2 10 3 9 10 9 13 15 2
33 0 3 10 1 10 9 9 1 9 13 1 9 1 10 13 10 10 9 9 2 15 3 13 1 9 2 10 7 9 3 13 3 2
35 10 3 3 0 7 0 9 13 10 13 2 10 7 0 7 10 0 9 13 2 10 3 13 10 0 9 2 10 7 9 13 7 13 15 2
30 16 3 10 0 7 0 9 0 10 15 13 13 9 10 9 2 9 13 1 10 9 9 13 0 3 7 13 10 13 2
62 9 3 13 0 2 10 3 13 13 7 3 3 13 3 7 13 0 13 10 9 2 10 7 13 1 10 9 7 13 10 9 10 3 13 2 3 3 7 10 13 0 10 9 1 9 10 13 13 10 9 2 3 0 0 13 10 9 10 9 10 9 2
10 10 3 3 1 15 9 15 13 9 2
38 1 3 10 15 9 10 3 0 9 13 9 2 10 13 1 9 1 10 0 9 2 10 7 9 13 13 10 10 9 9 7 0 9 13 7 9 15 2
26 10 3 1 10 9 13 10 9 13 1 9 1 10 13 9 7 13 0 10 9 13 10 13 10 0 2
11 10 3 13 10 9 13 7 13 10 0 2
18 13 3 9 9 10 0 9 2 7 0 9 13 0 13 10 9 15 2
19 10 3 0 0 10 9 13 1 10 1 9 9 0 13 13 3 10 9 2
23 3 9 3 10 1 9 1 0 13 1 10 9 2 15 13 16 13 0 0 10 10 13 2
11 9 3 13 10 1 10 9 1 9 13 2
9 10 3 3 9 13 10 0 9 2
25 10 3 9 13 10 1 10 9 7 10 0 9 1 9 13 15 2 13 10 0 9 10 0 9 2
26 13 3 7 13 15 10 1 10 9 2 3 13 10 9 2 3 3 3 13 2 3 13 1 10 9 2
31 10 3 9 2 10 3 1 9 15 13 2 10 7 1 9 13 2 13 7 3 1 10 13 13 2 13 0 13 10 9 2
43 1 3 10 15 9 10 3 9 13 3 7 13 13 1 10 9 10 0 9 1 10 10 9 0 9 2 10 7 9 1 0 13 10 0 7 10 9 13 0 13 10 13 2
8 0 3 13 3 10 13 9 2
35 3 0 3 13 15 3 3 2 16 3 13 10 9 10 9 13 3 15 1 10 9 13 2 1 7 10 9 1 10 9 3 13 3 13 2
26 3 3 13 7 13 10 9 10 9 0 3 13 0 9 10 0 2 0 7 15 1 10 9 13 13 2
22 10 3 3 1 9 9 0 13 10 9 2 10 7 9 10 0 9 13 1 10 9 2
15 13 3 15 3 0 7 9 9 2 10 7 9 1 0 2
19 9 3 10 3 9 0 15 10 0 13 0 2 10 7 9 0 7 9 2
32 1 3 15 3 10 9 13 7 10 0 9 13 2 3 7 10 13 10 9 9 13 10 9 13 13 10 9 3 1 10 9 2
53 13 3 10 0 13 9 1 10 9 10 9 13 2 15 1 0 10 1 10 9 9 13 13 0 16 1 10 9 2 3 13 10 13 3 9 7 0 13 10 9 13 1 10 9 2 16 1 10 9 13 9 13 2
32 13 3 10 9 3 7 13 2 3 7 9 7 9 13 10 9 13 1 10 13 15 2 3 13 3 15 13 10 13 10 9 2
42 10 3 13 1 10 1 10 9 9 10 9 13 7 13 10 0 1 10 13 9 13 3 13 10 9 1 15 10 9 2 13 10 0 7 0 9 10 13 10 9 9 2
33 13 3 10 9 3 13 7 13 10 9 2 10 3 13 10 9 13 2 13 7 10 9 7 1 9 13 10 3 9 7 10 9 2
58 10 3 9 13 10 9 7 9 13 10 9 7 9 2 3 7 9 1 10 9 13 10 13 3 1 10 13 2 13 7 1 10 13 15 13 13 7 3 13 10 9 2 1 3 15 0 10 9 1 9 13 13 1 10 13 10 9 2
20 15 3 3 13 2 0 3 9 3 13 13 2 0 7 9 10 9 0 13 2
10 9 3 0 10 0 1 10 9 13 2
34 1 3 15 10 9 13 1 10 9 10 13 16 13 10 3 9 10 9 13 13 9 10 13 2 10 7 0 13 1 10 9 10 9 2
19 10 3 3 9 13 2 13 9 0 7 0 0 7 0 2 9 7 0 2
22 10 3 9 13 10 9 7 10 10 0 9 7 13 1 10 9 3 13 1 10 9 2
13 10 3 13 9 0 7 0 0 13 1 10 9 2
16 3 13 9 0 13 1 10 1 10 9 3 13 13 10 13 2
13 13 3 15 13 10 9 7 3 13 15 3 13 2
22 10 3 9 1 15 9 13 2 10 3 0 10 9 1 9 13 2 10 7 13 13 2
16 13 3 1 9 9 0 2 13 15 13 1 9 9 7 9 2
17 10 3 9 10 3 9 13 13 7 10 0 13 13 13 10 9 2
18 3 13 9 0 3 10 0 2 0 7 10 15 9 2 1 15 13 2
39 0 13 3 10 0 9 1 10 9 7 10 9 2 13 7 10 0 9 7 13 15 15 1 9 0 7 0 2 13 13 10 0 15 13 13 13 1 15 2
6 15 3 3 13 13 2
48 13 3 10 10 9 9 3 16 10 0 7 0 10 10 0 9 13 1 10 9 2 3 13 16 15 13 1 10 9 13 2 13 7 10 0 9 1 10 9 13 1 0 10 9 1 10 9 2
13 10 3 3 9 7 10 9 10 9 13 0 3 2
17 10 3 0 3 3 7 3 13 10 3 0 9 13 13 7 13 2
22 16 3 13 7 13 1 10 1 0 9 13 13 2 1 15 0 3 1 10 9 13 2
20 10 3 3 9 1 10 9 2 16 0 10 0 13 2 1 9 13 10 9 2
26 10 3 9 10 0 0 13 9 7 10 9 13 2 1 7 15 0 13 10 9 3 10 9 3 13 2
33 13 3 10 13 9 9 0 2 0 13 1 10 13 9 2 3 7 13 3 1 3 10 9 7 10 3 15 9 2 13 1 15 2
37 10 3 9 0 3 0 1 9 2 3 7 1 9 13 2 3 1 10 10 0 9 2 7 1 10 10 13 9 2 1 0 9 13 1 0 9 2
23 1 3 10 13 3 10 10 9 9 13 15 3 0 2 0 7 10 9 13 0 10 9 2
44 10 3 9 13 10 9 3 1 9 7 1 9 13 7 13 0 3 13 10 9 2 13 7 16 13 10 13 9 1 10 9 13 10 9 10 9 13 2 13 10 9 1 9 2
10 10 3 3 13 13 15 10 0 9 2
26 10 3 13 15 15 13 10 13 10 9 1 10 13 15 10 13 16 3 13 13 13 10 9 10 9 2
26 10 3 3 9 3 3 13 10 0 2 10 2 15 3 13 2 0 13 13 15 1 9 7 9 13 2
32 10 3 9 13 16 3 13 15 0 15 3 13 0 10 3 9 2 3 0 13 10 13 13 2 7 3 13 10 9 10 9 2
51 10 3 9 10 9 13 10 13 1 10 9 10 9 2 3 3 13 10 10 9 9 2 3 3 3 13 7 3 16 0 13 13 7 0 9 7 9 13 13 1 15 15 0 7 0 10 1 15 9 13 2
26 0 3 1 10 9 10 10 9 9 13 1 10 9 7 10 9 2 13 10 13 13 7 9 15 13 2
47 10 3 13 1 10 9 13 10 13 10 9 3 1 15 3 13 2 7 16 13 15 7 13 10 0 10 9 1 3 10 9 3 9 7 9 3 15 3 10 9 13 13 7 10 0 13 2
14 10 3 9 13 10 13 7 13 15 3 10 9 13 2
22 13 3 3 3 1 15 10 1 10 9 13 9 10 9 7 9 15 9 1 10 0 2
56 16 3 13 1 10 9 10 9 1 9 13 7 15 3 13 10 9 1 9 7 13 1 9 13 2 15 13 9 1 10 10 0 9 9 16 1 9 13 10 0 7 13 3 0 13 10 0 2 13 15 3 13 0 13 9 2
27 15 3 13 10 9 13 10 9 13 3 10 9 2 13 15 10 13 10 9 1 0 9 13 13 10 9 2
24 15 3 13 0 3 1 0 7 0 2 9 3 0 2 10 7 10 9 9 0 3 10 0 2
40 10 3 9 13 10 9 10 3 9 13 1 10 0 9 7 10 9 13 1 10 0 10 9 2 1 0 3 15 13 13 2 10 3 3 0 13 13 10 0 2
14 13 3 10 3 0 9 13 3 0 9 13 10 0 2
19 3 3 1 9 10 3 13 10 9 13 3 7 15 0 13 1 10 13 2
25 10 3 0 3 13 1 10 9 2 13 1 9 7 1 9 10 9 13 13 15 13 13 10 0 2
32 10 3 13 10 9 2 10 3 9 13 1 0 1 0 10 9 1 9 13 2 10 7 9 10 9 1 9 0 15 1 13 2
22 10 3 0 10 3 1 10 0 9 13 2 10 7 0 3 10 9 0 10 9 13 2
10 10 3 9 13 13 10 0 13 3 2
37 10 3 0 9 0 3 16 3 2 0 7 13 10 3 1 10 9 9 3 13 13 2 10 7 1 10 9 2 0 13 10 1 15 2 3 13 2
30 16 3 0 1 10 15 9 3 3 7 1 9 0 13 1 10 13 9 2 13 1 9 2 13 10 9 10 15 9 2
54 1 3 10 10 9 10 3 1 10 9 13 13 7 13 10 10 0 9 2 10 7 9 1 0 10 9 13 7 13 10 0 2 3 3 3 10 10 9 9 1 10 1 15 9 13 10 9 7 13 13 1 10 0 2
19 10 3 3 9 10 9 3 1 0 10 9 13 1 10 0 13 10 9 2
31 10 3 0 10 13 1 10 0 9 2 3 3 13 10 10 9 9 2 3 7 13 10 0 13 1 10 0 9 10 9 2
12 13 3 15 13 7 13 15 16 1 10 9 2
41 10 3 1 10 9 13 10 3 0 13 1 10 9 10 9 13 7 13 3 1 9 9 13 2 10 3 3 0 9 10 9 1 10 9 10 13 1 15 0 13 2
87 16 3 10 3 10 0 13 9 13 3 1 10 9 13 1 15 13 13 2 10 7 1 0 10 9 1 10 3 13 7 1 9 13 10 9 1 0 7 13 13 10 10 9 9 13 2 3 3 3 13 10 3 0 10 9 13 1 10 0 9 10 9 2 10 3 0 13 1 10 9 10 9 1 15 10 10 9 9 2 3 7 15 0 1 9 13 2
37 13 3 0 10 9 2 3 15 10 3 1 10 9 7 10 9 13 2 0 7 3 10 1 9 10 9 13 1 0 0 13 1 15 15 0 13 2
51 10 3 3 1 10 9 0 13 1 0 10 1 10 0 10 9 13 2 10 7 9 13 3 1 0 10 1 10 9 10 13 1 13 10 9 2 10 7 0 9 13 1 9 10 9 7 10 1 15 13 2
14 10 3 3 9 10 9 10 13 13 1 10 9 3 2
22 10 3 9 10 0 13 7 10 9 3 1 10 0 13 13 0 10 13 1 10 9 2
17 1 15 9 0 15 3 3 13 13 1 9 10 10 9 9 13 2
22 3 3 10 13 10 9 2 7 3 1 10 9 2 0 13 0 3 1 10 9 9 2
22 10 3 0 0 3 13 9 7 9 10 13 1 9 15 13 13 15 1 10 15 9 2
33 9 3 9 7 0 9 10 3 0 9 7 0 13 13 13 2 10 7 3 13 3 9 7 10 13 9 10 9 1 10 0 13 2
12 15 3 15 13 1 10 10 13 10 9 9 2
32 3 10 3 3 3 0 2 16 1 0 9 7 9 13 10 9 2 10 7 3 0 2 16 1 9 13 13 1 15 10 0 2
17 1 15 13 0 9 0 1 0 9 10 1 10 0 9 13 9 2
16 0 3 15 1 9 1 0 9 7 9 9 0 13 10 0 2
8 15 3 3 15 1 15 13 2
27 9 3 2 1 9 0 15 13 2 9 9 3 13 1 3 10 1 10 9 9 7 1 10 1 15 9 2
22 9 3 15 9 7 9 13 10 9 9 1 3 0 9 13 3 2 3 7 3 13 2
17 10 3 0 7 0 9 0 3 10 9 2 0 7 10 9 13 2
33 15 10 3 0 1 3 10 9 7 10 10 0 9 0 3 3 13 1 0 9 13 2 10 7 0 3 1 0 15 13 7 13 2
20 13 3 3 0 1 10 9 10 9 9 2 15 13 13 0 13 10 13 9 2
29 9 3 2 13 15 1 9 10 1 9 13 2 3 13 1 10 13 10 9 7 10 9 13 10 1 10 9 13 2
19 10 3 9 1 15 13 13 10 9 2 13 0 13 10 1 10 9 13 2
16 1 3 10 9 7 9 10 9 3 13 13 9 13 10 9 2
29 13 3 15 13 10 9 10 9 7 13 3 1 10 9 13 10 9 2 10 3 13 9 2 10 7 1 9 13 2
13 0 3 13 9 0 13 7 13 10 9 10 0 2
21 10 3 9 10 0 13 13 0 7 0 9 7 9 13 9 9 7 9 9 13 2
12 10 3 13 13 1 10 9 16 1 10 9 2
23 13 3 1 10 9 10 10 9 9 2 15 3 1 9 3 3 13 9 13 0 0 0 2
16 10 3 1 9 13 9 13 1 10 9 13 3 1 10 9 2
29 13 3 10 9 3 7 13 10 10 9 9 0 13 9 7 0 9 16 3 3 13 3 13 1 10 9 10 13 2
43 10 3 0 7 9 1 10 0 9 0 0 13 13 9 2 10 7 0 10 3 0 13 2 10 7 1 10 9 1 10 9 7 10 9 13 0 13 9 10 0 7 9 2
13 15 3 0 9 1 9 9 1 9 3 13 13 2
14 15 10 9 3 3 1 10 9 16 1 10 9 0 2
11 1 3 13 10 9 10 9 7 9 9 2
23 15 13 10 13 13 3 0 2 13 15 10 1 10 9 9 10 10 13 9 9 13 13 2
15 3 15 3 0 9 1 0 13 9 3 10 15 9 13 2
33 1 3 3 10 9 1 9 7 10 15 9 13 10 9 10 3 0 13 1 10 1 0 9 13 10 9 2 3 7 3 3 13 2
17 1 3 10 9 7 1 10 13 16 13 7 13 2 0 9 13 2
34 15 3 3 7 3 15 3 13 7 13 13 2 16 3 3 13 10 15 9 7 9 2 1 15 13 13 15 0 9 13 0 7 0 2
45 10 3 9 2 13 10 13 9 10 10 9 9 7 13 1 3 9 0 15 13 1 10 13 9 2 1 7 9 1 10 13 10 9 9 2 13 0 1 3 10 0 7 0 9 2
31 3 10 3 9 3 13 1 10 9 2 13 15 10 3 13 7 10 1 10 9 13 9 2 1 7 15 9 0 7 0 2
14 15 3 13 0 13 9 7 15 10 1 10 9 13 2
22 10 3 9 13 1 10 9 3 10 3 9 7 10 9 13 7 0 13 13 10 0 2
17 9 3 10 1 10 9 13 13 10 1 9 3 3 13 10 13 2
16 3 13 3 3 13 2 3 13 1 9 0 7 0 13 9 2
13 13 3 1 0 9 9 7 15 13 13 10 9 2
23 3 3 10 1 9 9 13 2 7 13 3 10 9 2 10 3 13 9 9 13 1 9 2
8 10 3 9 13 15 13 13 2
10 13 3 1 10 9 13 3 0 9 2
25 1 15 15 0 13 13 1 10 10 9 9 2 10 13 3 9 2 3 3 7 13 10 0 9 2
21 1 15 13 1 0 9 1 10 9 2 13 9 7 13 10 9 1 0 13 9 2
24 3 3 3 3 3 1 15 9 13 10 9 2 13 1 10 9 0 10 9 3 13 10 9 2
8 15 13 9 0 13 10 0 2
12 13 3 10 9 7 13 10 9 13 1 9 2
27 3 3 13 3 3 1 9 10 9 1 10 9 3 13 9 15 10 9 16 0 10 0 7 0 9 13 2
14 1 3 10 13 9 13 3 0 13 10 10 9 9 2
19 10 3 3 9 3 13 13 10 9 2 1 7 10 0 9 0 13 9 2
6 3 15 13 3 3 2
81 10 3 9 2 13 9 1 10 1 10 9 9 16 10 9 10 3 9 15 13 7 10 0 13 10 9 2 3 13 0 10 9 16 1 0 9 10 1 10 13 9 3 3 1 10 0 9 2 3 3 1 10 0 13 10 0 1 0 7 0 9 3 13 3 13 10 9 7 1 10 0 3 13 9 2 13 10 10 9 9 2
18 9 3 0 7 9 13 1 0 10 9 2 13 10 0 7 0 9 2
21 3 3 13 10 9 10 1 10 0 9 9 7 9 3 13 1 9 13 10 9 2
18 3 13 9 9 9 7 9 9 13 0 9 3 13 7 13 9 3 2
72 10 3 13 10 9 9 2 13 13 10 9 1 10 13 9 2 13 10 3 9 10 9 1 10 0 9 1 10 9 13 2 10 7 9 1 10 9 13 10 0 9 13 10 9 2 13 13 10 10 0 9 13 10 9 2 13 1 10 9 10 9 13 7 13 1 10 9 10 9 10 9 2
22 10 3 9 2 13 15 13 2 7 13 13 10 9 15 2 13 10 9 1 10 9 2
24 15 13 9 2 16 3 13 13 10 9 2 3 13 0 10 9 13 1 10 9 1 10 9 2
27 13 3 10 9 15 1 10 9 2 13 1 10 13 9 10 9 2 16 15 13 13 10 1 10 9 9 2
27 16 3 10 9 13 10 9 7 10 9 2 10 3 3 10 0 13 13 2 16 0 15 13 10 9 13 2
51 13 3 13 15 13 2 15 3 10 0 1 10 9 7 9 13 2 13 2 16 13 10 9 1 15 2 13 10 9 3 2 16 7 13 2 13 1 10 9 7 3 1 15 13 13 1 10 13 10 9 2
19 10 3 1 10 9 0 13 13 10 9 7 13 1 1 10 0 10 9 2
25 15 3 10 9 13 1 10 1 10 0 9 10 0 13 9 13 2 0 3 7 0 13 10 13 2
29 1 3 10 15 0 13 10 9 13 10 10 9 9 1 10 9 7 13 1 15 13 10 9 0 13 1 10 13 2
9 13 3 15 3 13 1 10 9 2
10 10 3 13 10 9 13 10 9 3 2
31 3 13 1 0 1 9 13 10 0 0 13 7 13 9 13 10 0 0 7 0 3 15 13 2 10 7 0 13 13 3 2
22 9 3 1 0 3 9 13 0 2 10 7 0 10 9 13 1 10 9 13 13 0 2
21 15 3 13 3 0 13 13 10 9 9 10 3 13 10 0 9 7 13 10 9 2
32 10 3 9 0 13 1 10 9 2 0 13 3 3 1 10 10 0 13 10 9 13 2 16 1 10 10 0 13 10 9 13 2
33 3 3 3 13 1 15 1 10 1 9 9 1 10 1 9 7 0 9 10 9 1 10 9 13 2 13 1 9 9 13 10 9 2
17 13 3 10 0 1 10 9 13 10 9 0 9 16 1 10 9 2
7 9 3 13 10 9 0 2
29 13 3 1 10 9 2 3 7 10 0 3 9 15 13 2 13 13 2 16 13 15 3 13 10 9 1 10 9 2
21 3 3 1 3 0 10 9 3 10 9 10 13 13 7 10 0 13 9 10 9 2
35 3 3 15 0 13 1 10 13 13 3 13 7 0 13 1 10 13 9 1 10 0 9 13 15 2 0 7 10 0 9 13 9 1 9 2
26 16 3 3 10 13 10 9 0 10 13 13 2 13 1 9 13 1 9 10 9 7 9 15 10 13 2
13 15 3 3 10 3 9 13 0 2 15 7 0 2
62 10 3 9 10 9 13 3 0 2 10 7 9 10 9 0 9 13 9 2 15 10 3 1 9 13 2 1 7 10 0 9 13 9 13 2 10 7 1 10 9 13 13 3 10 9 10 1 9 9 2 13 7 10 9 3 0 0 2 13 7 9 2
45 1 3 15 9 0 13 10 9 2 1 15 3 13 10 9 13 10 9 2 9 3 3 13 7 1 9 0 7 9 1 9 2 1 15 13 1 10 9 9 0 13 9 7 9 2
35 15 3 13 1 0 9 10 9 7 10 1 10 9 9 3 9 7 9 13 13 13 9 1 10 0 13 10 9 9 16 1 10 0 9 2
59 13 3 0 7 0 10 9 2 7 10 9 10 3 13 1 0 9 2 10 7 13 2 3 3 7 10 9 13 3 3 3 1 10 9 2 13 0 9 7 9 1 10 13 2 3 13 1 10 9 1 10 0 9 0 10 0 1 0 2
29 3 3 3 10 3 9 15 9 15 13 10 9 2 7 10 3 13 2 10 7 13 3 10 13 9 13 10 0 2
49 3 3 1 0 9 13 7 10 9 13 2 16 3 13 9 13 2 0 1 0 10 9 7 0 9 3 13 3 1 9 7 3 2 16 0 3 13 0 1 10 0 9 10 13 13 1 10 9 2
40 10 3 0 9 10 3 10 9 1 10 3 9 0 13 10 9 2 1 15 9 13 13 15 10 10 9 0 2 7 3 0 13 10 9 13 10 9 10 9 2
34 10 3 13 3 13 10 13 10 9 7 13 1 9 2 0 9 7 9 13 2 16 13 10 1 15 9 7 3 13 10 13 10 9 2
48 13 3 3 10 9 2 3 1 15 13 1 3 10 9 9 10 9 10 9 10 13 1 9 1 10 13 1 10 9 1 15 9 2 1 7 10 0 0 9 1 10 1 15 9 15 7 9 2
27 10 3 13 10 9 3 13 2 3 7 13 10 13 0 9 1 10 9 2 3 13 15 13 1 10 13 2
19 9 3 3 1 10 13 9 1 0 13 13 10 9 2 13 1 10 0 2
35 9 3 0 9 13 1 10 9 3 0 10 9 7 10 9 2 7 3 10 9 7 10 9 2 3 7 9 0 13 10 3 13 10 0 2
65 10 3 1 10 9 15 3 15 13 2 13 7 10 1 10 9 9 2 13 9 0 9 7 13 10 13 9 10 9 10 1 15 13 9 2 15 13 9 3 9 9 7 7 0 9 0 2 13 1 9 2 13 3 13 2 13 7 1 9 10 9 13 10 13 2
35 13 3 0 7 0 9 2 13 0 10 9 7 13 1 0 10 9 10 9 13 10 9 2 13 13 7 1 9 0 10 9 1 10 9 2
34 10 3 1 10 9 9 13 1 10 9 0 3 3 13 10 13 2 3 7 1 10 0 10 9 0 13 1 9 7 9 13 10 13 2
17 9 3 3 7 3 13 7 13 1 10 9 1 9 13 10 9 2
36 10 3 1 10 9 0 3 3 13 1 10 10 9 9 0 2 3 0 9 7 9 13 2 16 1 10 3 13 10 9 13 10 9 10 9 2
63 13 3 10 9 10 13 1 0 7 13 9 13 1 3 10 9 10 9 10 1 0 13 7 10 1 0 13 9 15 7 9 1 9 2 3 13 7 13 3 13 2 7 13 15 2 3 3 13 7 13 10 9 13 2 13 13 1 9 7 13 10 13 2
40 1 3 0 3 13 10 13 15 13 10 13 1 10 9 0 9 3 10 9 7 10 9 10 9 13 7 13 10 9 1 0 10 13 1 10 9 0 13 9 2
17 10 3 13 2 13 10 9 1 10 9 1 0 9 13 10 9 2
26 10 3 9 1 10 13 10 13 3 3 7 3 13 2 7 3 13 1 10 13 7 13 10 0 3 2
14 0 3 1 0 9 13 15 13 9 0 1 10 9 2
18 10 3 3 1 10 9 13 3 0 0 2 10 7 3 3 0 15 2
41 0 3 13 10 9 1 9 13 10 9 3 1 10 15 9 2 15 0 13 10 9 2 16 3 1 0 9 1 9 7 1 9 3 0 13 1 10 13 10 9 2
16 3 3 3 10 3 9 7 10 9 13 13 1 0 10 9 2
40 10 3 3 1 15 13 2 9 3 9 7 9 13 2 3 3 7 3 3 13 13 10 9 16 10 9 1 10 0 13 9 2 3 13 13 10 10 0 9 2
32 10 3 10 9 9 13 1 3 10 9 0 13 2 15 7 1 15 13 2 3 13 13 10 9 2 13 10 15 13 10 9 2
21 10 3 9 1 15 13 10 0 13 10 9 2 9 13 10 9 7 0 13 3 2
27 10 3 3 9 1 10 9 0 13 3 3 1 10 9 13 10 0 1 10 9 1 9 10 10 9 9 2
25 1 3 10 9 10 9 7 10 9 10 1 10 9 9 3 0 13 9 10 9 1 10 9 15 2
26 10 3 10 9 3 3 13 2 3 3 13 3 1 10 10 9 10 9 1 10 1 10 9 9 13 2
8 10 3 13 10 0 9 13 2
32 3 13 1 15 10 1 10 9 13 9 2 10 1 9 9 13 3 9 0 1 0 9 0 10 0 13 7 13 10 9 13 2
31 10 3 9 10 9 1 0 10 9 2 1 0 13 0 0 10 9 13 2 13 13 1 10 9 7 9 10 13 13 9 2
53 10 3 0 1 10 0 10 9 13 3 13 10 0 10 3 9 7 10 13 16 3 0 0 13 10 9 13 7 10 9 2 0 13 13 10 9 10 0 2 7 3 0 13 13 13 10 9 2 16 13 10 0 2
22 15 3 13 1 15 13 1 10 9 10 9 2 13 13 0 9 0 10 10 0 9 2
33 3 10 0 3 3 13 0 15 0 9 13 2 10 3 9 3 10 13 13 2 10 3 13 0 13 2 10 7 9 13 10 0 2
19 0 3 13 1 10 9 15 10 1 10 0 1 10 9 3 13 10 9 2
33 13 3 7 13 3 3 1 10 1 10 9 9 13 10 1 10 9 9 1 9 3 16 10 1 10 9 13 9 10 9 13 0 2
15 1 15 9 3 13 0 1 9 10 1 10 9 9 13 2
17 10 3 10 0 9 13 3 0 13 10 13 10 9 10 0 13 2
14 1 15 10 9 13 10 13 13 10 9 10 9 13 2
78 1 3 3 10 0 9 10 9 15 13 1 10 9 10 9 7 1 10 15 13 10 13 13 7 13 10 3 2 7 1 3 10 9 7 10 10 9 9 10 13 3 1 10 9 13 7 13 2 1 7 0 9 13 9 13 9 1 0 9 2 1 15 9 13 9 13 7 10 0 0 13 2 13 10 9 10 9 2
19 15 10 9 13 7 9 13 0 0 10 13 2 3 7 10 0 2 13 2
12 10 3 1 9 13 9 1 15 3 13 3 2
14 13 3 1 9 15 10 9 13 2 13 10 9 13 2
8 10 3 3 0 13 3 13 2
14 10 3 10 9 9 13 2 9 13 13 13 10 0 2
19 13 3 10 0 1 3 10 9 7 1 10 9 10 9 13 10 0 0 2
29 10 3 9 2 13 3 0 10 9 3 13 7 13 15 10 1 10 9 2 3 13 10 13 7 13 1 10 9 2
49 10 3 13 10 3 9 3 13 2 10 7 13 7 13 10 10 0 9 13 2 13 0 9 9 13 0 9 7 9 1 0 10 10 9 9 16 3 10 9 13 7 10 13 15 9 10 9 13 2
23 1 0 9 13 15 10 0 0 10 9 10 9 1 10 10 9 9 13 10 9 10 9 2
24 10 3 13 7 3 13 0 10 1 10 9 13 2 13 10 9 1 0 9 13 9 10 9 2
53 16 3 3 10 3 9 1 10 9 3 13 1 10 3 13 2 10 7 10 9 9 13 1 0 10 9 7 9 2 10 3 9 10 9 0 13 13 7 0 2 10 7 9 7 9 10 9 1 9 0 7 0 2
52 0 3 9 13 10 13 10 13 16 3 13 7 13 13 10 13 2 7 13 1 10 1 15 13 9 7 10 9 2 3 7 10 10 9 9 2 3 0 13 7 13 2 3 13 13 1 0 10 10 9 9 2
25 0 3 0 13 13 10 9 1 10 0 1 10 13 9 2 15 0 9 1 10 13 13 10 9 2
26 10 3 9 0 13 13 10 9 10 9 16 3 10 9 10 9 7 10 9 10 9 1 10 9 13 2
14 15 3 13 10 3 3 1 10 9 13 13 10 9 2
22 13 3 7 9 13 9 10 9 2 3 7 10 0 9 9 13 10 9 13 10 9 2
15 10 3 1 10 9 10 13 13 9 3 13 3 10 9 2
32 15 1 10 9 13 7 0 13 1 10 9 2 13 10 9 10 9 10 9 9 9 13 9 13 13 1 10 9 0 10 9 2
12 15 3 13 13 1 0 9 2 13 10 0 2
12 3 10 3 9 0 13 2 0 13 10 9 2
22 1 3 10 9 10 0 1 10 9 9 13 2 13 9 10 3 0 13 1 10 0 2
29 0 3 1 15 13 7 13 10 9 10 0 13 0 9 9 13 7 0 13 1 10 3 13 15 1 0 13 9 2
20 3 3 10 3 9 13 1 10 9 2 10 7 1 10 9 0 13 1 9 2
34 3 3 15 13 1 10 9 7 13 13 7 3 13 2 13 7 13 10 9 13 1 9 13 7 13 1 10 15 9 13 15 1 9 2
26 13 3 10 13 1 9 0 13 10 9 2 1 0 10 9 1 0 9 10 9 13 10 10 0 9 2
61 9 3 10 10 9 9 13 10 3 0 1 10 15 9 3 13 7 13 10 9 7 1 10 13 13 2 10 7 0 9 10 3 1 3 10 9 13 10 3 1 0 10 9 2 10 7 13 1 10 9 2 0 13 13 7 13 10 9 3 3 2
36 3 3 10 3 1 10 9 10 7 1 10 9 1 10 9 13 2 3 0 9 13 1 10 9 0 2 7 3 10 9 13 10 9 15 13 2
19 3 3 3 3 10 13 13 10 9 1 0 10 9 3 13 0 10 0 2
31 10 3 9 0 13 3 3 3 1 0 10 9 2 3 7 13 1 0 10 9 1 10 9 13 10 0 10 0 9 9 2
50 3 3 3 10 13 3 10 13 13 15 13 13 1 10 9 2 13 7 0 1 9 13 1 10 9 10 3 9 13 10 9 1 9 2 13 1 10 9 10 9 1 10 13 10 1 10 9 13 9 2
15 1 15 13 0 10 9 13 1 0 10 9 13 10 9 2
16 16 3 3 15 13 2 13 10 9 1 0 10 9 13 15 2
21 10 3 3 0 0 13 10 9 2 3 3 0 10 0 1 10 0 9 9 13 2
16 3 3 3 13 10 9 1 10 0 9 1 0 13 10 9 2
35 10 3 3 13 0 13 1 10 9 10 9 7 10 10 9 9 2 10 7 9 0 13 15 2 16 13 10 9 1 10 1 10 9 9 2
19 16 3 13 15 1 10 0 2 3 13 3 1 10 13 1 10 13 9 2
25 3 13 15 10 0 2 3 13 1 10 0 7 1 9 2 1 10 9 1 10 9 13 10 9 2
8 10 3 3 9 0 15 13 2
41 10 3 3 13 3 13 1 3 0 13 2 1 10 9 13 10 9 2 3 7 10 13 1 10 1 9 9 3 10 0 13 13 1 9 7 1 10 9 13 13 2
40 13 3 3 1 10 0 9 7 3 13 10 3 1 0 13 2 15 1 10 13 13 0 2 3 13 1 3 10 9 10 9 2 3 3 7 10 9 10 9 2
25 3 3 13 10 13 1 9 13 1 10 13 1 10 9 7 3 0 13 9 10 13 13 10 13 2
29 10 3 0 9 2 13 0 7 0 2 13 10 9 7 10 9 2 0 3 10 9 10 9 1 10 9 13 13 2
52 13 3 10 9 0 9 3 13 1 10 9 2 16 1 15 7 1 10 0 9 7 9 13 2 9 7 1 10 9 13 7 13 0 2 16 3 7 3 10 9 13 7 10 1 15 3 0 9 13 10 9 2
11 3 3 1 15 0 9 7 9 13 13 2
27 3 3 10 3 9 2 3 15 13 2 1 10 1 10 0 9 15 13 10 13 2 7 13 10 3 9 2
37 3 3 13 10 1 10 9 9 2 9 0 13 3 10 0 15 13 9 9 2 10 3 9 13 10 10 9 13 7 10 0 9 7 9 10 9 2
9 1 3 3 0 15 13 0 9 2
41 10 3 9 13 1 10 9 7 13 10 13 10 9 1 3 10 9 7 10 0 9 13 1 9 1 10 9 2 13 0 0 9 7 10 9 3 1 0 9 0 2
24 3 3 13 10 9 10 0 0 7 15 10 0 9 13 2 13 13 10 9 10 1 10 9 2
26 15 3 1 10 9 13 2 10 3 1 9 13 1 10 9 13 7 1 10 1 10 0 0 9 13 2
62 1 3 10 0 9 9 3 9 10 1 10 9 13 7 10 0 9 13 1 10 9 2 9 7 10 13 13 0 9 13 1 15 13 15 0 13 2 13 3 13 10 13 1 10 9 10 0 9 2 15 3 16 0 13 13 2 10 3 0 9 13 2
31 13 3 10 9 7 13 10 9 1 10 0 7 10 3 13 10 7 13 10 9 2 0 13 13 9 1 10 10 9 9 2
32 13 3 15 1 10 9 7 13 9 2 13 9 10 10 9 13 7 13 3 10 9 13 10 13 2 13 10 1 10 9 0 2
20 10 3 9 2 10 0 3 15 13 2 3 1 0 7 1 10 13 13 9 2
35 10 3 10 9 9 0 10 9 10 3 13 10 7 13 2 1 15 0 1 10 9 13 16 1 9 13 2 13 13 10 1 10 9 13 2
27 13 3 10 9 9 0 9 13 0 7 13 2 13 13 2 13 13 1 10 13 10 9 1 10 13 9 2
19 3 3 3 10 1 10 9 13 9 13 10 13 13 9 10 9 10 0 2
34 10 3 13 3 3 15 0 13 1 9 2 13 1 0 9 10 1 15 13 2 0 3 2 9 7 13 7 9 13 1 10 9 0 2
22 3 13 10 9 7 10 3 9 7 10 0 10 1 10 9 13 13 10 9 10 0 2
27 10 3 9 13 10 3 0 13 13 15 2 13 10 3 9 13 1 10 9 13 2 10 7 9 3 13 2
40 3 13 3 10 9 2 7 0 13 3 2 7 10 9 0 13 7 0 9 2 0 10 10 9 13 9 13 13 1 0 9 2 1 15 13 13 10 9 15 2
34 10 3 1 10 9 13 9 2 16 10 1 10 9 13 2 13 10 9 13 10 9 3 1 10 9 2 15 13 10 1 10 13 13 2
31 10 3 10 9 9 2 13 10 9 15 3 10 9 10 0 2 13 13 1 9 2 13 15 3 0 13 10 0 9 13 2
62 10 3 9 13 1 0 10 9 10 10 9 7 10 9 10 9 2 3 13 13 7 13 3 0 13 1 10 3 13 10 0 2 13 1 9 0 7 1 0 9 0 13 2 13 0 13 15 2 15 13 13 3 16 10 0 0 10 0 9 0 13 2
46 13 3 9 7 9 13 1 10 9 0 2 10 3 10 9 9 1 3 10 10 9 7 10 10 9 9 13 10 13 7 13 10 13 13 10 9 13 10 9 7 13 10 9 10 9 2
52 13 3 3 2 15 3 0 13 7 3 13 10 9 1 0 13 2 10 7 10 9 9 2 10 9 13 7 10 9 1 9 13 0 2 3 13 16 3 10 9 15 13 0 2 7 0 15 3 7 3 13 2
14 9 3 10 3 9 13 2 10 7 9 3 3 13 2
27 10 3 3 9 3 13 10 1 10 9 2 7 10 3 13 1 9 3 2 10 7 13 15 1 10 0 2
30 10 3 9 13 1 10 9 1 10 9 7 0 13 2 13 1 10 13 15 7 13 10 13 2 13 13 10 13 9 2
23 3 3 0 15 13 9 2 13 13 10 9 7 13 10 3 10 9 9 7 10 9 0 2
45 10 3 9 13 3 9 1 9 10 9 1 10 1 10 9 13 9 1 9 7 9 2 3 7 0 7 13 1 10 9 2 9 7 1 0 13 10 1 10 9 9 1 10 9 2
36 0 3 1 0 3 10 9 2 13 0 2 13 10 10 9 10 0 9 2 15 3 0 13 10 3 9 7 10 0 9 10 1 10 9 9 2
18 10 3 9 1 0 10 9 13 2 3 0 13 7 0 3 10 9 2
41 1 3 3 10 9 13 9 2 3 3 7 10 1 9 9 13 3 0 10 9 7 3 3 10 10 9 2 13 3 3 10 9 3 7 10 0 9 9 15 13 2
20 10 3 9 1 15 9 13 15 9 10 9 13 2 15 10 1 10 9 13 2
10 15 13 10 0 9 13 13 10 9 2
7 9 3 13 0 10 9 2
13 13 3 9 0 13 1 10 13 9 1 9 0 2
38 0 3 10 9 10 3 9 3 13 10 0 9 2 1 15 10 13 9 0 13 7 0 2 1 3 10 0 9 3 13 2 0 7 9 1 9 0 2
28 13 3 9 0 1 3 10 1 9 9 7 10 1 10 9 13 2 10 7 1 15 13 0 7 0 13 9 2
23 13 3 1 15 3 9 2 15 3 3 9 2 3 3 9 0 13 9 1 10 13 9 2
23 13 3 3 9 0 1 10 1 9 7 9 9 1 10 9 2 1 15 9 9 0 13 2
44 0 3 3 3 13 1 9 10 0 10 9 13 1 10 9 9 2 0 7 1 9 13 15 9 1 10 9 9 1 3 0 9 0 7 0 9 13 1 9 3 1 0 9 2
14 1 15 3 0 3 1 10 9 10 1 9 13 9 2
45 10 3 3 9 7 10 9 2 1 15 1 0 9 13 1 15 9 2 9 2 9 2 9 2 3 3 10 13 13 13 2 10 7 13 0 3 7 0 3 1 10 9 13 9 2
21 1 3 10 0 9 1 15 7 10 9 10 9 3 3 15 1 9 13 10 13 2
27 3 3 10 1 9 9 3 10 1 10 9 7 10 13 9 9 7 10 1 0 7 0 13 9 15 13 2
13 9 3 3 0 13 1 0 9 3 0 3 13 2
27 10 3 3 9 0 13 0 2 10 3 1 10 9 3 0 1 10 9 2 10 7 9 10 9 0 3 2
20 15 0 13 3 10 10 3 1 9 9 0 13 1 9 2 0 7 13 15 2
16 15 3 0 3 13 13 1 10 9 2 10 1 9 9 13 2
20 10 3 3 13 3 1 10 0 0 13 1 10 15 9 7 3 1 9 13 2
27 3 3 3 16 0 9 10 9 13 0 0 1 10 13 9 7 10 13 9 1 0 9 7 9 0 13 2
40 10 3 9 2 10 9 10 9 13 1 3 10 9 7 1 10 9 2 16 13 2 13 10 9 10 9 2 15 13 1 10 3 9 7 10 1 10 9 13 2
47 1 15 13 3 3 13 7 13 13 10 10 9 13 10 9 2 3 7 10 9 13 2 10 3 0 3 13 7 10 9 3 3 15 13 2 16 3 10 9 1 0 9 7 0 9 13 2
55 3 3 3 3 3 0 3 0 10 0 9 7 9 13 1 15 2 0 3 9 9 13 2 0 7 9 7 9 9 13 2 9 3 2 16 9 13 2 13 7 13 2 7 3 3 0 7 0 0 9 0 13 10 9 2
27 0 3 16 15 15 13 2 3 0 9 3 1 0 10 9 13 2 1 0 9 13 13 10 9 10 9 2
14 10 3 3 1 10 9 7 10 0 9 0 13 9 2
12 10 3 9 13 15 0 10 13 10 0 9 2
40 15 3 3 3 13 10 9 1 10 9 2 0 7 10 9 13 13 10 9 2 16 3 3 3 13 15 3 15 13 2 7 3 15 13 13 10 0 15 13 2
84 3 3 9 13 2 3 9 3 3 0 10 1 9 9 3 13 1 3 10 9 7 1 10 13 1 0 10 0 9 13 10 9 2 3 13 3 13 15 9 1 10 9 3 3 1 10 9 10 10 9 9 2 13 10 0 13 10 1 10 0 9 9 2 13 1 10 9 0 2 16 3 13 10 9 2 3 3 3 9 13 10 9 13 2
5 15 3 9 13 2
24 10 3 3 0 13 10 9 13 10 1 10 9 9 2 10 7 0 13 10 1 10 9 9 2
29 3 3 0 13 0 10 9 2 1 15 13 7 10 1 10 9 9 10 9 13 10 1 9 9 9 13 10 0 2
8 13 3 10 9 10 13 9 2
12 9 3 3 3 13 1 10 9 1 10 0 2
19 3 3 3 1 10 10 13 9 1 10 0 9 7 9 13 1 10 9 2
29 1 3 10 10 9 9 1 9 3 0 7 0 13 13 9 13 2 1 15 10 9 13 2 1 9 10 9 13 2
33 15 3 3 13 10 1 10 9 9 10 3 1 10 9 9 13 7 10 1 10 9 9 2 0 13 1 10 0 10 10 9 0 2
94 13 3 1 10 1 10 9 9 9 7 15 1 10 9 13 2 3 3 15 13 10 0 13 2 3 7 13 10 9 10 9 9 7 13 10 1 9 9 16 3 13 1 10 1 9 9 9 10 0 13 2 3 0 7 0 13 13 10 9 2 7 1 0 9 9 7 9 13 10 9 3 10 9 10 7 0 10 1 10 9 9 13 9 13 1 10 13 1 3 0 9 10 9 2
47 10 3 9 2 1 10 9 13 15 10 13 9 10 9 7 3 13 10 9 2 3 13 10 9 2 7 13 9 7 10 0 0 13 10 9 2 13 15 13 10 1 10 9 9 10 9 2
10 13 3 3 9 1 10 0 9 9 2
45 15 13 7 13 1 10 9 13 9 13 10 0 13 13 1 10 9 3 10 3 9 13 7 13 10 9 2 13 7 9 1 10 0 10 0 7 9 1 15 2 3 13 10 0 2
35 10 3 9 13 10 9 10 1 10 9 7 13 10 9 15 2 13 1 10 0 9 10 0 9 13 1 10 9 9 10 1 10 9 13 2
18 3 13 10 13 10 9 10 9 13 10 9 3 13 1 10 3 9 2
48 1 3 10 0 2 3 10 9 13 2 13 10 3 0 0 9 13 7 0 2 15 7 0 13 10 9 1 9 10 9 2 0 7 0 13 10 9 2 10 3 0 13 15 13 13 10 13 2
8 3 13 3 13 10 13 9 2
11 13 3 10 10 0 9 13 13 1 9 2
22 10 3 9 3 13 10 9 10 9 2 3 1 0 13 9 0 13 10 0 10 9 2
24 10 3 9 13 10 9 15 13 10 9 2 13 10 9 7 13 1 9 15 0 13 10 0 2
25 10 3 0 9 10 0 13 9 10 1 10 9 13 9 2 3 10 9 0 10 9 3 0 13 2
19 9 3 3 10 3 9 13 7 10 9 0 1 10 1 10 9 0 13 2
23 10 3 9 13 13 15 10 9 13 2 10 7 9 1 9 9 0 1 10 0 9 13 2
8 1 3 10 9 0 15 13 2
34 10 3 3 9 13 3 13 1 10 9 2 10 3 9 3 13 0 7 1 9 13 2 10 7 0 0 7 0 0 9 7 0 0 2
18 1 3 10 3 3 3 10 9 13 10 9 13 13 13 10 0 9 2
25 3 1 10 13 1 0 9 10 9 13 3 13 2 7 0 3 15 9 13 2 0 7 13 0 2
30 10 3 0 9 13 10 9 7 13 3 13 1 10 9 9 2 3 7 3 1 9 15 1 10 13 9 10 9 13 2
27 10 3 3 10 9 9 13 1 10 9 7 10 9 1 10 10 0 9 7 10 9 9 13 2 0 13 2
14 3 3 0 10 0 13 9 10 13 9 1 10 9 2
26 10 3 9 2 13 15 3 10 9 2 10 3 9 7 10 9 3 0 13 13 2 10 7 9 13 2
19 3 3 13 3 10 1 10 9 9 0 15 13 2 13 10 9 10 0 2
18 13 3 15 7 9 9 0 13 2 0 9 7 0 9 13 3 13 2
12 3 3 13 1 10 9 13 15 1 10 0 2
11 10 3 3 3 13 9 9 0 7 0 2
41 1 3 3 1 10 1 9 13 0 9 1 10 13 2 15 10 0 7 0 13 13 13 2 7 0 10 10 13 1 10 13 9 2 16 3 15 0 9 2 13 2
33 16 3 13 10 9 2 7 10 1 9 15 3 13 1 10 13 10 13 2 3 3 7 3 13 10 13 1 9 7 9 13 9 2
22 10 3 0 0 9 13 10 13 13 10 3 10 13 2 3 3 7 10 10 13 9 2
30 10 3 9 3 13 10 13 1 10 13 10 0 9 13 7 13 3 10 9 2 13 9 13 10 9 0 0 9 13 2
14 15 3 13 1 10 9 2 3 13 10 9 10 9 2
10 3 13 9 0 10 13 1 10 9 2
16 15 3 13 10 3 0 15 3 13 2 0 7 13 10 9 2
29 10 3 3 9 10 9 13 0 2 0 9 13 2 10 7 9 13 9 13 2 0 1 10 9 13 7 10 9 2
37 10 3 3 9 7 9 13 1 9 9 1 15 7 15 13 10 9 2 9 13 0 7 0 3 2 9 15 15 13 9 13 0 3 0 7 0 2
32 1 15 1 10 0 9 7 9 2 16 13 0 2 3 3 10 3 0 16 0 2 3 7 0 13 0 9 9 13 1 15 2
41 16 3 15 13 13 10 9 10 9 9 1 10 9 2 15 10 3 9 1 10 9 7 3 9 7 9 1 15 13 2 3 3 3 13 0 9 13 1 9 13 2
33 3 15 3 13 10 0 2 13 15 3 2 16 13 10 0 7 0 13 9 3 16 3 3 3 13 0 9 7 13 0 9 13 2
23 3 3 3 1 3 0 10 9 3 13 10 9 13 2 16 1 10 9 15 10 9 13 2
13 1 15 3 15 1 0 0 7 10 13 3 0 2
21 10 3 3 9 0 2 3 7 16 9 13 0 1 10 3 1 10 1 15 13 2
15 10 3 3 13 2 10 7 0 7 3 0 13 10 9 2
47 1 1 3 10 13 9 10 3 10 9 0 9 0 13 15 3 13 3 0 10 9 7 3 10 9 2 3 7 10 1 10 0 9 2 10 3 3 9 3 0 0 7 0 1 0 9 2
27 9 3 3 9 7 9 0 0 9 10 3 13 10 9 13 2 9 3 1 9 9 10 1 15 13 9 2
13 1 3 10 9 0 0 15 7 0 0 13 13 2
30 1 15 1 10 3 0 1 10 9 2 7 3 1 10 13 3 3 13 10 9 2 0 13 10 0 13 9 10 13 2
43 16 3 0 13 10 13 9 13 10 1 10 9 9 1 10 9 10 9 2 3 15 3 13 10 9 2 10 7 1 10 9 9 9 13 1 10 13 10 9 1 10 9 2
46 13 3 10 13 3 13 1 9 13 15 7 9 13 10 9 2 13 9 13 10 9 1 10 10 13 7 13 10 13 10 9 13 13 1 10 9 1 10 0 3 16 10 3 13 13 2
15 10 3 3 9 13 0 10 9 3 13 10 1 10 9 2
55 13 3 0 9 3 3 7 1 9 2 10 3 0 13 10 9 7 10 13 9 13 10 9 2 16 3 13 3 10 1 10 9 15 2 13 7 10 13 2 13 0 1 0 9 10 13 9 2 13 1 10 13 0 0 2
91 3 3 13 1 10 9 7 13 3 13 10 9 2 16 3 10 0 9 13 2 3 0 13 10 9 1 10 9 2 13 10 9 16 3 1 9 13 2 3 15 3 9 0 7 3 9 13 2 10 3 3 13 10 3 2 10 7 13 3 13 1 15 2 7 10 0 9 15 0 9 13 1 10 9 2 15 13 1 0 9 3 13 10 9 13 10 9 1 15 13 2
35 10 3 0 13 1 10 9 7 1 0 9 13 9 7 9 2 15 0 13 0 9 7 3 16 13 0 3 0 0 13 9 2 13 3 2
28 3 3 13 2 15 3 15 13 10 13 15 10 9 1 10 0 7 13 0 10 13 15 13 13 13 10 9 2
30 0 3 13 10 9 2 15 10 9 1 10 0 10 9 13 15 13 2 0 13 9 7 0 9 10 13 1 15 9 2
73 3 1 10 13 0 1 10 9 2 7 13 9 10 13 9 1 10 9 3 10 9 3 0 10 9 7 10 9 13 2 7 3 13 10 9 10 9 7 10 3 9 10 9 13 13 9 0 10 1 0 13 9 2 3 9 7 9 13 7 9 0 13 2 3 3 1 9 2 3 7 3 0 2
21 16 3 3 3 0 7 0 13 2 13 9 3 9 7 10 13 9 0 10 9 2
50 9 3 3 13 0 7 0 9 2 1 3 10 3 3 13 13 7 0 13 10 13 3 13 2 13 1 0 9 10 9 2 1 7 10 13 9 3 9 7 9 13 3 13 7 13 10 13 3 13 2
30 3 3 0 0 13 9 13 10 0 9 2 16 3 1 9 7 9 13 1 15 2 7 13 10 0 7 0 13 9 2
8 15 3 3 13 13 1 15 2
8 10 3 0 9 15 13 9 2
16 3 3 13 13 0 3 0 13 7 0 0 13 1 15 9 2
10 10 3 3 9 13 10 0 9 0 2
11 0 13 1 10 9 13 10 9 7 9 2
8 15 13 3 3 13 10 9 2
38 1 3 10 15 13 3 10 9 3 10 3 13 9 10 13 9 1 9 1 15 7 13 15 10 9 3 13 3 15 2 10 7 15 15 13 15 13 2
25 9 3 3 13 3 10 9 2 13 3 10 1 9 9 2 13 7 1 10 9 13 1 10 9 2
21 3 13 13 3 3 0 7 0 9 10 9 1 10 13 9 2 0 13 10 0 2
16 10 3 9 3 1 9 13 10 15 9 2 16 13 15 9 2
40 0 3 3 13 2 1 0 9 13 0 9 0 2 13 0 9 0 9 1 10 0 9 2 15 7 0 3 2 13 10 9 7 10 9 7 1 15 10 9 2
77 0 13 9 13 0 3 15 13 1 10 13 2 0 7 15 13 1 10 13 2 3 3 7 3 13 10 9 0 13 2 13 13 10 9 15 2 7 10 3 10 0 9 13 0 13 2 16 15 13 7 13 10 9 2 10 7 10 9 3 0 13 9 2 13 13 0 15 2 15 3 3 15 13 16 1 9 2
60 13 3 0 10 1 0 9 1 10 0 13 2 16 3 13 3 7 13 10 9 7 9 10 9 2 13 7 7 13 1 10 13 15 1 9 1 10 0 9 9 3 0 9 13 3 3 1 15 1 10 9 2 7 3 10 0 9 15 3 2
21 3 1 10 13 10 1 10 9 15 10 9 3 13 7 10 13 9 13 10 0 2
24 13 3 3 15 2 3 10 13 9 1 0 9 10 0 13 1 10 9 9 13 15 13 13 2
24 3 3 3 15 0 7 0 13 2 1 0 13 10 9 1 10 0 9 7 0 1 15 13 2
22 3 3 3 0 10 0 13 10 9 2 13 13 1 10 13 9 10 1 9 13 9 2
35 1 3 3 9 10 9 2 1 15 13 1 10 9 2 3 13 2 13 3 0 1 15 13 10 3 13 1 15 10 7 9 3 13 13 2
30 1 3 9 3 13 3 2 15 13 3 1 9 9 2 13 7 15 9 10 13 1 3 10 15 7 3 1 10 9 2
7 3 13 15 1 10 13 2
17 10 3 0 13 1 10 13 2 13 15 0 13 10 1 9 9 2
17 9 3 13 1 10 13 10 13 10 13 2 1 9 13 10 9 2
32 15 13 16 13 15 10 9 13 2 7 1 10 9 9 13 13 2 0 13 3 13 7 13 2 13 13 10 9 10 1 9 2
40 3 13 10 9 13 16 1 10 9 13 10 0 9 1 10 9 13 3 10 1 15 9 1 15 10 9 7 13 1 10 1 15 9 0 13 10 1 10 9 2
36 0 3 13 10 0 10 0 9 7 13 0 9 1 10 10 9 10 3 9 13 10 7 9 10 3 9 7 10 9 13 2 13 3 1 9 2
30 16 3 15 0 13 13 2 3 0 15 13 16 10 13 0 13 7 13 13 10 1 10 9 2 3 13 10 9 13 2
17 3 0 3 10 0 9 1 10 9 3 10 9 7 10 9 13 2
12 3 3 15 13 2 16 13 1 10 9 13 2
21 3 16 15 13 13 13 2 3 13 3 3 7 3 16 15 13 13 10 3 13 2
17 3 15 3 13 13 1 0 10 9 2 13 15 9 9 7 9 2
33 3 3 3 10 9 3 13 10 9 2 13 7 13 13 15 7 13 3 2 13 10 9 13 10 9 15 2 9 10 9 13 13 2
37 10 3 1 15 13 16 3 10 13 9 9 13 13 10 3 0 1 10 13 10 0 10 9 2 1 7 15 13 10 3 9 7 10 1 15 9 2
52 10 3 1 10 9 7 10 9 13 0 3 3 13 10 9 2 16 0 15 13 7 0 2 13 10 10 9 9 7 10 3 9 10 9 1 10 9 13 2 10 7 9 7 10 1 15 13 3 1 9 13 2
21 3 10 0 13 3 3 1 10 9 2 9 0 7 1 10 0 10 9 9 13 2
18 10 3 3 1 10 9 7 0 13 9 1 15 7 15 13 10 9 2
32 10 3 1 10 9 13 10 13 3 3 13 9 1 10 1 10 9 9 2 13 1 10 9 7 13 15 13 7 13 10 9 2
73 9 3 10 3 1 0 9 3 13 1 10 1 10 9 9 2 10 3 0 9 7 9 13 1 10 1 10 9 9 2 3 7 13 13 0 9 2 3 0 3 15 3 0 13 3 2 7 3 1 15 13 0 10 13 13 2 3 1 0 9 7 9 13 2 16 1 10 9 15 10 9 13 2
19 13 3 1 10 1 9 9 3 13 13 10 9 9 0 13 7 9 13 2
5 13 3 15 0 2
8 0 3 13 9 9 7 0 2
24 1 3 15 3 9 9 2 3 0 9 2 3 9 9 1 15 13 2 3 3 0 9 13 2
17 3 3 3 9 9 7 0 7 0 10 13 3 9 3 0 13 2
17 3 3 3 3 13 0 13 9 0 7 0 9 0 9 7 9 2
13 3 0 3 15 15 10 0 7 0 0 13 0 2
90 1 3 10 13 9 0 9 13 13 3 13 10 1 10 9 9 2 13 3 10 0 0 10 9 10 0 2 0 7 10 9 10 9 16 3 13 2 9 3 10 0 7 9 3 0 1 15 10 13 13 2 13 7 7 13 10 3 9 3 10 3 7 3 10 9 13 2 7 10 15 3 13 0 9 7 9 2 10 7 1 10 9 0 13 2 15 9 13 9 2
16 3 10 3 9 3 0 9 1 10 9 2 7 9 0 13 2
40 10 3 9 10 10 1 10 9 13 13 10 0 9 7 9 1 10 9 2 3 13 1 9 1 15 15 13 10 13 15 2 13 10 9 13 3 1 10 9 2
38 3 0 13 9 10 1 10 9 7 9 16 3 0 13 10 13 10 9 10 0 1 10 9 2 15 13 1 10 9 2 7 3 1 10 0 13 9 2
20 3 3 13 1 10 13 0 2 3 7 3 1 10 13 13 3 10 3 13 2
43 3 3 3 3 1 0 0 13 10 9 2 13 10 9 9 1 10 13 15 3 0 15 10 1 10 9 10 9 13 2 13 3 0 2 13 7 10 1 10 9 10 9 2
8 13 3 7 13 10 0 9 2
29 10 3 9 0 3 1 9 13 2 13 7 13 10 9 2 10 3 10 9 10 7 15 3 9 13 1 10 0 2
16 10 3 13 9 15 10 9 10 9 3 0 7 0 9 13 2
27 0 3 1 3 10 1 10 9 13 9 3 3 10 10 9 13 9 2 1 7 0 1 10 9 10 9 2
42 1 15 0 3 13 10 0 7 13 1 10 9 10 9 0 13 0 10 9 2 7 3 3 9 2 3 7 3 3 13 1 10 9 1 9 7 9 0 13 10 3 2
9 9 3 1 3 10 9 3 13 2
9 3 3 13 1 0 10 9 0 2
8 13 3 1 10 9 0 13 2
14 3 3 10 9 3 13 7 10 0 9 3 7 3 2
7 13 3 3 0 0 9 2
17 3 1 15 13 9 9 0 3 13 3 16 13 13 3 10 13 2
31 13 3 1 10 9 10 9 3 10 9 7 3 0 10 1 10 9 9 7 13 1 10 9 13 13 1 10 10 0 9 2
24 10 3 9 13 1 10 9 2 3 13 10 9 7 10 9 10 0 13 0 13 1 10 9 2
30 3 0 3 15 13 13 1 10 9 2 10 7 13 9 1 0 9 0 7 9 13 2 13 10 1 0 10 9 9 2
58 10 3 9 13 9 7 9 13 2 15 16 3 13 13 10 9 1 0 9 7 0 13 15 2 13 3 3 9 13 10 9 7 13 10 0 2 10 3 9 13 7 3 10 9 2 15 7 13 1 10 9 13 1 10 10 9 9 2
25 13 3 10 9 0 7 10 10 13 9 2 15 9 1 10 15 13 1 10 9 13 10 0 0 2
55 3 0 3 1 0 10 9 3 13 3 2 7 3 1 0 9 1 10 13 9 13 15 10 0 2 13 9 3 3 1 9 1 10 13 3 7 1 9 2 3 3 13 3 15 10 0 2 0 13 15 3 7 3 13 2
57 3 10 9 13 15 3 13 10 9 2 9 10 13 9 3 13 2 7 15 13 1 10 13 9 9 2 13 0 3 9 3 10 13 10 0 7 10 13 1 10 0 2 1 7 15 0 9 7 0 2 16 10 0 1 0 13 2
38 15 1 10 0 3 9 13 10 0 10 9 13 3 10 9 10 0 2 13 3 10 10 9 9 2 13 7 0 10 13 9 7 10 1 10 9 9 2
12 10 3 13 13 1 15 1 10 9 0 0 2
92 10 0 10 13 10 9 10 13 10 9 1 10 9 13 0 7 0 13 9 1 10 9 2 13 10 1 10 9 0 10 1 10 13 9 3 13 9 9 13 2 1 7 15 10 13 9 9 13 1 0 9 3 10 1 10 9 10 1 10 9 9 7 1 10 9 10 9 0 1 10 0 13 2 0 7 13 1 15 9 2 3 0 13 10 9 3 2 9 1 15 13 2
26 1 15 13 10 9 3 0 9 10 9 13 2 7 3 10 1 0 13 13 3 3 13 13 10 0 2
21 1 15 13 9 3 0 9 7 9 9 13 1 10 13 1 10 9 13 0 15 2
45 10 13 9 1 10 1 9 9 13 1 0 9 9 13 10 9 7 0 13 10 1 0 10 9 9 2 13 0 10 9 10 1 10 9 7 13 1 15 10 9 13 10 13 9 2
19 13 3 10 9 2 9 13 13 0 1 10 9 10 13 9 13 10 9 2
31 0 3 10 9 13 3 10 1 10 9 7 10 0 2 10 3 9 13 1 10 9 2 13 10 9 1 10 10 9 13 2
25 16 3 1 0 13 15 2 13 1 0 10 9 13 2 9 13 3 13 15 0 7 13 10 0 2
28 10 3 9 13 3 10 9 0 13 10 9 2 1 3 15 10 9 7 10 0 2 0 7 10 0 10 9 2
13 13 3 0 13 10 0 2 13 13 0 10 15 2
13 3 10 3 1 10 9 13 9 13 10 9 13 2
18 10 3 1 10 9 1 9 13 1 9 13 13 1 10 10 0 9 2
16 0 10 3 10 3 13 13 13 7 13 15 3 7 10 0 2
15 10 3 0 13 2 1 9 10 9 13 15 7 10 9 2
16 13 3 3 1 0 10 9 7 10 0 2 13 7 1 0 2
51 9 3 13 10 9 10 13 9 2 13 1 9 10 0 7 10 3 1 10 9 9 1 9 13 2 13 7 13 1 10 9 10 1 15 0 2 10 7 0 9 13 10 3 13 2 0 7 1 9 13 2
18 10 3 9 0 15 9 13 7 9 2 1 0 15 13 10 13 9 2
26 1 3 10 9 0 3 1 10 9 7 10 9 13 2 13 13 15 7 3 13 10 1 10 9 9 2
37 10 3 9 13 1 10 9 1 0 10 9 10 0 1 0 13 2 10 9 13 10 9 2 13 1 10 13 3 10 1 9 9 2 13 1 0 2
20 10 3 0 9 15 10 1 9 9 13 1 10 9 1 10 1 10 9 9 2
29 10 3 9 13 1 0 9 3 9 13 2 13 10 1 10 9 7 9 9 1 10 9 0 13 10 1 10 9 2
37 13 3 10 9 10 3 10 9 9 0 7 1 9 2 10 3 10 9 1 9 2 10 7 1 10 9 1 9 2 0 15 9 13 13 7 0 2
45 1 3 10 9 0 9 2 15 13 3 9 10 0 9 2 13 7 3 0 9 0 2 0 3 3 3 13 1 10 9 0 13 9 2 3 7 3 13 1 10 9 10 9 9 2
23 3 3 13 13 0 9 1 9 0 7 9 2 13 1 10 9 13 1 15 9 1 0 2
11 3 13 10 9 3 13 2 13 10 9 2
20 10 3 9 13 10 9 7 13 15 10 9 2 1 9 13 13 13 10 9 2
28 13 3 3 7 13 10 10 9 9 2 13 10 9 10 9 7 10 9 10 1 15 13 0 3 1 10 9 2
12 10 3 10 3 13 2 10 7 13 10 9 2
9 3 3 13 7 13 1 10 9 2
18 10 3 13 1 9 13 0 3 9 13 2 3 7 13 9 13 0 2
49 9 3 15 13 3 13 3 1 3 10 1 10 9 9 7 10 1 10 9 9 10 9 2 16 3 0 13 9 15 13 10 9 2 7 3 10 9 13 13 1 9 2 13 15 10 1 9 9 2
32 13 3 10 9 2 10 3 9 13 10 1 15 13 13 9 2 13 1 0 2 10 7 9 13 15 10 9 0 13 10 0 2
19 10 3 1 10 9 13 1 15 10 9 7 13 1 10 9 13 10 9 2
23 13 3 9 0 13 10 1 10 9 2 3 3 10 9 13 2 0 7 10 9 13 9 2
21 10 3 3 9 7 9 13 2 10 7 0 13 3 1 0 2 13 7 1 0 2
42 13 3 10 9 2 9 10 3 13 10 0 1 15 13 9 13 7 13 10 1 10 0 9 2 10 7 3 13 13 13 13 2 3 3 10 3 9 15 13 10 13 2
21 1 3 15 13 15 13 9 0 1 15 2 3 2 7 13 15 2 0 13 9 2
29 1 3 10 0 9 10 10 9 10 9 13 10 0 2 13 10 1 10 9 7 9 2 13 10 1 10 9 9 2
19 3 10 3 3 1 15 13 9 9 13 1 10 9 1 10 15 9 13 2
49 3 3 10 9 9 13 1 9 9 2 3 3 0 10 9 13 10 9 7 13 1 15 2 13 9 9 10 13 2 3 15 3 13 2 1 7 15 13 13 9 0 10 1 10 9 9 13 13 2
27 3 10 0 3 13 10 9 1 15 13 3 10 9 2 16 3 13 1 10 9 13 1 15 1 10 9 2
18 10 3 0 3 0 1 15 13 9 3 0 13 13 13 1 10 13 2
56 9 3 7 9 2 1 7 15 9 10 9 13 10 9 9 1 10 0 7 13 16 10 0 9 13 13 1 10 13 9 10 3 9 7 10 10 0 9 2 13 3 3 13 15 10 1 9 1 9 13 10 9 1 10 9 2
7 13 3 15 13 10 0 2
15 13 3 15 0 13 2 3 13 1 10 1 10 9 9 2
39 10 3 9 13 10 3 9 7 10 1 15 0 2 15 13 1 10 9 2 16 3 13 2 13 3 2 3 13 15 1 10 9 10 9 1 10 15 9 2
25 13 3 10 9 0 10 9 0 3 13 3 13 10 1 10 9 10 10 9 13 9 1 10 0 2
39 1 3 15 13 13 16 13 10 1 10 9 13 3 1 10 0 2 0 7 13 10 0 9 2 9 0 7 9 0 13 13 2 15 13 0 15 13 0 2
24 3 3 15 13 15 13 0 0 2 3 1 10 1 10 9 13 2 0 10 1 10 9 13 2
21 1 15 9 10 9 13 0 13 9 13 10 15 9 10 0 13 10 1 9 9 2
26 3 13 15 13 2 15 13 2 10 15 13 10 9 2 15 3 3 15 10 0 7 0 13 1 9 2
11 10 3 0 15 13 9 7 0 13 13 2
22 15 3 13 13 10 3 9 7 10 1 15 13 7 10 0 13 0 10 9 13 13 2
15 0 3 13 15 1 10 9 1 10 0 10 9 15 13 2
7 3 3 13 13 13 3 2
15 0 3 3 10 0 13 10 9 1 10 9 10 13 9 2
12 3 13 15 3 10 9 2 15 3 13 13 2
44 0 3 13 1 0 9 3 7 13 0 13 10 9 1 10 13 1 10 9 1 15 9 2 3 3 10 13 15 13 0 2 3 3 3 0 2 0 7 1 10 0 9 13 2
23 16 3 3 13 16 10 9 13 2 7 15 1 10 13 13 13 2 0 3 13 10 13 2
11 3 15 3 3 1 9 13 13 10 13 2
20 10 3 1 10 9 13 2 13 1 0 2 13 1 10 9 10 1 10 9 2
38 3 13 0 1 10 9 0 3 13 10 9 2 13 10 9 1 10 9 2 15 0 9 0 1 0 9 13 13 3 9 15 2 13 7 1 10 13 2
10 16 3 10 9 13 2 13 10 0 2
13 13 3 7 10 9 13 3 13 13 1 0 9 2
38 10 3 9 10 9 15 13 13 3 15 13 2 13 7 7 0 13 10 9 1 3 9 7 10 0 10 9 9 9 13 2 13 13 7 13 10 13 2
12 1 3 10 13 9 13 1 10 10 9 9 2
29 10 3 3 13 2 13 7 10 13 3 9 13 1 15 7 9 2 3 10 0 9 13 10 13 15 3 9 13 2
18 1 3 10 0 13 7 13 15 2 15 3 3 13 9 2 13 13 2
7 15 3 3 13 3 13 2
38 3 1 15 13 3 3 15 13 13 16 3 0 10 9 10 9 7 15 10 1 15 13 9 7 9 13 13 7 3 0 13 2 0 7 3 10 9 2
24 1 3 3 10 9 2 16 3 9 10 15 13 15 2 1 0 3 15 13 0 13 10 9 2
23 16 3 3 13 2 1 10 1 15 9 13 10 0 3 13 9 2 16 3 13 10 13 2
20 10 3 9 3 0 3 13 9 7 9 16 15 0 9 7 0 13 10 9 2
23 15 16 3 9 0 13 7 9 2 9 7 9 13 10 13 0 7 0 13 1 10 13 2
25 16 3 13 2 13 10 9 3 13 15 10 13 7 0 0 3 13 2 1 0 13 10 0 9 2
8 9 3 13 13 10 0 9 2
34 10 3 9 0 3 7 0 9 0 9 0 7 9 1 9 0 2 0 7 3 0 2 0 7 10 0 10 3 10 13 9 7 9 2
21 15 3 3 13 3 1 3 10 9 10 0 2 3 7 3 1 10 9 15 13 2
25 9 3 13 10 10 0 9 10 3 9 1 15 13 2 13 13 3 10 9 0 13 9 10 0 2
36 10 3 0 15 3 13 2 10 3 1 9 9 13 2 10 7 9 1 15 13 13 10 9 2 0 13 9 0 2 16 13 10 0 3 13 2
23 13 3 10 9 0 9 13 3 1 10 9 2 13 15 0 7 0 1 15 9 10 9 2
38 10 3 3 9 13 1 15 13 1 15 1 15 16 3 0 10 1 10 0 13 9 2 7 3 1 15 0 0 9 13 10 0 1 10 1 15 9 2
25 15 3 3 13 10 9 10 3 9 10 9 13 13 2 10 7 0 13 2 15 3 10 9 13 2
37 1 3 15 3 10 13 9 1 10 1 15 13 9 2 1 15 13 10 0 9 1 3 10 9 7 10 0 0 2 13 13 1 9 3 1 9 2
26 10 3 1 10 9 2 16 3 13 2 13 13 2 0 15 3 3 9 13 10 9 0 1 10 9 2
33 3 3 1 10 0 1 10 9 9 7 1 10 9 3 15 3 10 0 9 7 9 13 2 1 7 10 9 0 9 13 7 9 2
30 10 3 3 13 15 1 15 2 13 1 0 2 7 10 9 15 13 0 13 1 10 9 2 10 7 9 13 10 9 2
11 10 3 3 9 3 13 13 10 13 13 2
19 15 3 13 10 3 1 10 9 7 9 13 10 13 13 13 0 10 9 2
7 9 3 13 9 10 9 2
34 15 3 13 10 9 1 10 9 2 16 10 9 10 9 13 13 13 1 10 1 10 9 15 13 9 1 10 13 10 9 9 1 15 2
34 3 9 13 15 3 7 9 13 10 9 2 13 10 9 10 1 10 9 7 9 2 0 15 13 9 1 3 15 7 15 9 10 9 2
11 10 3 3 1 10 0 9 1 15 13 2
13 10 3 9 13 3 13 13 1 10 9 9 9 2
60 9 3 3 3 3 1 10 13 9 0 13 9 1 0 10 13 1 15 2 3 7 3 3 13 2 13 13 15 3 1 10 1 9 9 7 1 10 9 9 10 13 9 2 16 3 3 13 10 13 3 13 10 13 2 3 3 7 3 13 2
22 3 3 13 10 15 13 7 0 15 13 9 2 1 15 3 1 10 13 13 0 13 2
15 3 3 3 3 9 13 10 1 10 9 0 9 15 13 2
14 1 9 3 3 13 0 9 1 0 1 0 0 9 2
31 10 9 10 13 1 9 1 9 7 13 10 0 13 1 15 2 7 3 13 15 1 10 9 1 10 0 2 13 10 9 2
28 1 3 15 13 7 13 1 9 0 1 15 13 16 3 10 9 13 10 13 1 15 0 1 10 1 9 9 2
14 1 3 0 10 9 1 0 10 13 3 7 3 13 2
20 3 3 1 3 10 9 13 10 0 13 3 10 13 2 1 7 10 0 13 2
26 1 3 15 10 3 1 10 9 0 2 1 0 9 1 10 9 13 2 13 15 1 10 9 3 13 2
16 10 3 9 13 15 2 3 13 2 13 10 1 10 9 0 2
14 9 3 3 10 1 10 13 0 13 9 13 10 9 2
14 10 3 1 10 9 7 9 3 0 13 13 16 13 2
20 1 0 3 15 10 1 10 9 9 13 10 0 16 13 9 15 13 10 9 2
44 1 3 0 9 13 10 3 0 10 0 7 9 2 10 0 1 0 2 1 15 13 3 9 10 9 13 10 1 15 13 2 13 3 13 1 10 0 7 13 10 1 10 9 2
25 10 3 3 0 9 13 2 13 10 9 7 10 1 10 9 9 2 10 7 0 7 0 13 13 2
22 1 0 9 13 10 3 9 7 9 15 15 13 10 0 2 1 7 10 9 3 13 2
27 3 3 13 2 16 13 2 13 1 0 10 9 0 13 9 9 0 7 0 9 9 7 9 0 7 0 2
47 0 3 3 15 1 10 1 9 9 13 7 13 16 0 9 3 13 2 0 7 1 10 0 9 10 3 1 9 0 13 13 2 10 7 3 7 3 3 3 1 9 3 7 3 13 13 2
10 15 0 13 9 2 0 13 10 9 2
32 1 3 3 10 9 3 13 13 2 0 10 9 7 10 9 10 13 13 2 1 7 9 3 13 13 9 2 13 15 10 13 2
20 13 3 3 10 1 10 9 9 1 10 10 13 9 0 13 13 1 15 0 2
59 16 3 13 3 3 10 0 2 9 0 13 2 13 3 10 0 10 9 2 13 7 1 10 9 15 2 3 0 10 9 1 10 9 1 10 0 10 9 13 2 13 10 1 10 9 3 9 7 9 13 15 10 0 7 13 1 9 9 2
17 13 3 9 7 13 9 1 9 13 2 13 0 2 1 10 9 2
7 1 15 9 9 13 0 2
13 13 3 15 3 9 13 10 13 13 1 10 9 2
21 10 3 3 1 10 9 7 9 7 10 0 10 0 9 0 10 9 13 10 9 2
55 10 3 9 2 16 10 9 13 10 9 2 13 15 13 1 10 10 9 13 2 7 1 0 10 9 13 1 10 9 2 13 15 9 10 3 9 7 10 0 9 0 13 2 0 13 10 0 2 1 10 9 10 9 13 2
17 15 13 1 10 9 10 9 1 10 3 13 9 0 13 10 9 2
21 13 3 10 13 10 3 9 3 9 13 0 1 10 0 2 3 13 3 10 9 2
14 15 3 1 9 7 1 9 10 9 13 7 10 9 2
17 1 3 3 10 1 9 9 13 9 2 1 7 10 3 15 9 2
15 1 3 15 13 1 10 9 10 1 10 9 0 13 3 2
51 15 3 3 3 1 10 10 9 9 13 7 13 3 15 3 13 2 15 7 13 13 7 13 0 10 9 10 0 1 10 10 9 9 2 10 9 16 3 1 9 0 3 13 9 1 9 10 1 15 9 2
18 10 3 9 3 3 13 10 9 10 1 10 9 1 10 9 10 9 2
14 3 3 13 3 3 13 1 10 9 1 10 3 9 2
21 3 13 1 10 9 7 13 1 10 0 9 13 1 10 9 10 9 7 10 9 2
14 10 3 9 0 10 9 15 13 3 7 3 13 3 2
12 3 3 13 10 9 1 9 13 3 10 9 2
10 3 3 13 10 13 10 1 10 9 2
69 3 3 0 3 10 0 13 7 1 15 10 0 3 13 9 9 2 3 7 13 2 1 7 15 10 0 10 1 10 9 13 2 0 0 13 15 2 13 1 10 9 2 13 0 10 10 9 1 0 9 13 10 9 1 10 13 9 7 13 15 13 2 13 1 10 13 10 9 2
29 3 0 15 13 13 3 0 10 0 1 10 9 2 13 7 10 9 1 10 9 2 3 3 13 13 1 10 0 2
16 16 3 0 13 10 1 10 9 0 2 13 13 15 1 0 2
40 13 3 10 9 1 10 9 2 10 3 0 10 9 1 0 10 9 13 2 10 3 1 0 9 13 1 3 0 13 15 2 10 7 9 0 13 10 0 9 2
15 10 3 3 0 9 10 9 1 10 9 3 13 10 9 2
18 3 3 1 0 10 9 0 13 9 10 9 7 10 15 0 13 3 2
20 3 3 3 13 15 3 9 15 7 9 3 13 15 9 13 7 9 13 9 2
33 10 3 3 0 9 1 0 13 9 9 0 13 10 9 16 3 0 13 3 10 9 10 9 2 7 3 10 0 10 9 13 3 2
20 10 3 9 2 13 10 0 10 9 1 10 9 0 9 13 10 1 10 9 2
31 9 3 3 9 7 9 3 9 13 10 0 1 10 9 9 2 15 15 13 9 13 2 0 15 10 15 9 7 9 13 2
23 9 3 1 10 9 0 1 10 1 10 9 13 0 1 15 13 13 13 1 10 13 9 2
53 10 3 3 13 10 13 9 2 1 0 9 3 13 1 10 13 1 10 3 13 10 1 9 9 2 13 10 9 3 0 13 10 9 2 7 3 0 9 7 0 13 10 9 1 15 3 1 10 13 13 10 9 2
5 15 3 3 13 2
7 9 0 10 0 13 9 2
31 13 3 9 13 0 10 9 13 2 9 9 9 2 15 9 3 0 7 9 13 2 9 3 1 12 9 3 1 12 13 2
21 1 15 3 15 13 9 9 2 9 9 9 2 15 0 13 12 9 1 10 9 2
14 1 3 10 9 10 13 9 9 13 2 9 9 9 2
18 7 15 3 13 13 9 3 7 10 9 9 9 2 9 3 7 9 2
37 15 3 3 10 9 13 10 10 9 9 2 10 3 9 0 1 10 9 10 9 13 10 9 10 9 13 2 16 3 10 10 9 9 10 9 13 2
12 9 3 9 13 13 9 13 16 10 13 9 2
34 16 3 9 13 0 2 13 9 15 9 0 2 15 13 9 13 9 2 1 15 15 13 0 3 13 10 9 2 3 10 9 15 13 2
11 1 15 9 10 1 9 7 9 13 9 2
19 13 3 15 9 12 10 9 10 9 13 10 9 2 10 13 16 13 0 2
11 15 3 10 13 15 10 9 9 13 13 2
33 13 3 7 9 7 9 9 0 9 2 9 3 7 9 9 7 9 2 9 3 7 9 9 2 9 3 7 9 9 9 9 9 2
28 10 3 10 9 9 1 9 1 9 13 9 13 9 2 15 15 9 13 1 15 15 1 9 1 10 9 13 2
10 1 3 3 9 15 9 13 9 9 2
18 15 3 13 15 13 2 16 3 13 9 13 16 1 10 9 15 13 2
18 13 3 9 7 10 9 9 2 7 13 1 10 9 13 1 10 9 2
14 0 3 10 9 13 7 10 9 15 7 10 9 13 2
7 9 3 1 9 13 9 2
10 13 3 15 1 9 9 9 13 13 2
15 15 3 13 9 1 9 9 13 9 2 16 9 13 13 2
12 13 3 9 1 9 7 13 10 9 13 9 2
39 13 3 9 9 2 13 1 0 9 1 10 3 13 2 7 15 13 0 13 13 2 16 13 9 13 9 1 10 13 1 15 13 9 2 15 9 9 13 2
5 15 13 13 15 2
19 10 3 9 9 9 3 13 9 15 1 9 13 2 13 10 1 9 9 2
27 9 3 13 9 1 10 9 0 1 9 13 2 16 1 9 13 13 0 9 2 1 15 13 3 9 13 2
5 11 3 13 10 11
5 11 3 13 10 11
5 11 3 13 10 11
15 11 3 13 10 11 10 9 11 1 15 13 11 10 13 11
22 6 10 9 1 9 13 7 13 9 7 13 10 9 15 11 15 13 13 1 15 10 9
6 3 3 13 1 10 9
12 13 3 15 6 9 9 13 1 9 10 11 13
21 13 13 10 9 7 10 9 15 7 13 1 9 11 13 3 10 13 10 9 10 9
15 13 3 15 16 13 10 9 1 10 9 0 13 9 10 11
11 15 9 13 1 15 13 7 15 13 1 15
9 7 13 9 12 7 12 9 0 13
4 13 15 10 11
9 13 3 16 11 13 13 1 10 11
8 15 3 3 13 10 9 13 15
8 7 13 10 9 15 13 15 13
11 13 7 13 16 10 9 15 0 1 10 9
12 15 3 3 13 10 9 15 8 0 13 10 9
18 13 3 15 16 13 12 10 9 15 7 3 0 10 9 15 13 1 11
9 7 1 10 9 16 9 13 10 9
15 7 10 13 15 13 7 10 9 15 13 13 15 7 10 9
7 3 3 10 0 10 15 13
3 6 13 15
4 13 10 9 15
4 13 10 9 15
7 13 10 9 10 9 3 13
5 10 3 3 13 15
21 9 13 0 1 10 9 15 10 9 7 3 13 13 10 9 1 10 9 10 9 15
15 15 3 15 3 13 16 13 15 10 9 3 3 15 13 15
7 10 3 0 9 9 0 13
22 15 3 15 13 15 10 9 0 7 13 15 13 9 0 15 13 15 10 9 1 10 9
7 7 13 10 9 13 15 13
5 13 3 10 9 13
7 0 3 13 13 15 13 0
10 9 13 15 0 13 7 13 10 9 15
4 15 0 13 0
10 16 13 15 13 15 1 10 9 10 9
2 13 9
11 13 13 15 10 9 7 13 1 10 9 15
4 15 3 13 13
9 15 3 13 9 9 0 1 9 0
10 7 13 10 9 0 1 0 10 9 0
6 7 13 15 10 11 13
17 13 3 10 9 13 1 15 16 13 13 7 13 3 9 3 13 9
10 13 3 3 1 10 9 10 13 9 11
14 1 15 3 3 9 7 9 13 13 15 1 15 0 13
5 13 3 1 10 9
4 6 3 13 15
12 13 3 3 10 13 7 9 7 9 13 1 11
4 15 13 10 13
4 9 1 0 13
11 10 3 0 1 10 9 10 9 0 15 13
10 13 10 9 10 9 13 7 13 7 13
19 1 11 13 16 16 1 11 13 10 9 10 13 1 15 13 3 1 10 3
11 10 3 9 15 13 7 13 13 9 7 13
8 7 13 3 13 1 10 9 15
11 13 3 10 9 9 13 1 15 16 15 13
6 1 0 15 9 13 15
7 1 3 10 9 10 9 13
30 3 3 13 11 1 10 9 10 9 12 9 7 12 9 3 13 10 9 10 9 1 10 9 10 9 12 9 7 12 9
8 3 13 7 10 9 0 10 0
20 7 13 1 15 9 0 16 15 1 9 13 13 7 15 10 9 1 10 9 13
6 1 15 1 9 13 15
13 15 3 0 10 9 16 13 7 10 9 15 16 13
13 13 10 9 10 9 9 13 0 9 1 10 9 15
19 0 13 10 9 10 9 9 15 13 9 13 1 9 9 12 16 15 13 0
10 10 3 0 9 0 13 10 9 10 9
15 0 13 10 9 10 9 9 13 1 10 9 15 13 9 13
3 13 0 15
9 7 10 9 15 3 15 1 15 13
5 13 3 10 11 15
14 7 13 13 0 9 7 13 1 15 7 13 10 0 15
4 13 15 3 15
10 13 3 10 9 13 7 13 13 13 13
10 3 13 10 11 1 11 9 7 9 13
7 9 3 13 1 15 11 13
11 15 9 15 3 13 10 9 15 10 0 13
13 1 3 10 9 13 9 0 9 9 9 9 9 9
4 15 3 13 13
6 6 9 0 15 10 9
5 7 13 15 10 9
4 7 13 15 13
10 7 10 12 9 10 12 7 15 9 13
2 13 15
9 7 13 15 10 11 13 13 15 13
14 15 3 13 9 16 10 9 0 13 10 3 9 15 13
14 16 13 13 3 12 9 15 12 7 11 12 7 11 12
6 7 13 15 10 9 13
11 7 13 15 10 9 15 7 3 13 15 13
1 6
9 15 3 0 13 1 10 9 10 9
17 16 3 10 9 15 7 10 9 15 13 15 13 15 7 13 1 15
14 16 3 13 10 9 15 13 13 15 1 15 7 15 0
11 9 3 13 1 15 10 9 15 7 13 15
20 13 3 10 9 0 13 12 10 9 15 15 13 15 12 9 7 13 15 13 13
20 3 3 10 9 15 10 0 13 15 16 3 13 0 10 9 15 1 10 9 15
8 15 3 10 9 13 9 3 13
8 9 15 0 13 16 13 9 0
3 15 0 13
4 15 3 13 13
19 0 3 13 10 9 10 9 9 9 15 13 3 3 13 9 1 10 9 15
2 13 15
4 9 3 13 15
18 3 13 15 10 9 10 9 11 1 10 9 15 13 7 13 15 1 15
2 13 15
21 7 16 13 1 11 7 13 1 11 1 10 9 10 9 3 11 13 12 9 13 15
12 0 3 13 9 1 10 9 7 13 1 10 9
6 15 3 15 13 9 9
9 3 3 1 15 9 13 1 10 9
7 7 15 15 13 10 9 0
2 3 13
6 13 3 10 0 13 3
8 10 3 9 7 10 9 13 15
19 1 0 13 15 16 13 1 15 10 9 10 9 7 13 9 13 10 9 15
4 6 1 10 9
3 7 13 15
6 3 3 13 1 9 9
1 9
9 1 10 9 3 15 10 12 13 9
7 9 15 9 0 1 10 9
2 13 15
8 7 9 3 13 15 1 10 9
10 15 3 3 13 1 10 9 10 9 13
7 0 13 13 7 0 3 13
8 7 15 13 10 9 10 9 15
9 3 3 15 13 1 3 16 3 13
6 7 13 10 11 13 15
5 15 3 0 9 9
18 13 3 3 9 0 15 3 13 1 9 9 1 10 3 7 3 3 13
7 10 3 9 15 3 3 13
16 1 0 7 15 13 0 16 15 3 13 9 10 9 10 9 13
8 13 3 10 9 13 15 7 13
20 13 3 15 13 13 10 9 7 10 0 13 1 15 1 10 9 7 13 10 9
15 10 3 10 12 13 13 13 9 7 13 10 9 10 9 15
7 13 3 10 10 12 9 13
10 7 13 13 13 10 9 15 1 10 9
9 3 13 10 9 7 10 9 10 9
12 1 15 13 12 0 10 9 15 10 0 15 13
4 3 13 15 13
25 10 3 11 13 1 11 1 9 11 10 0 13 15 9 13 9 9 0 7 13 1 10 9 15 13
3 6 13 15
3 7 13 15
4 3 15 13 9
10 13 3 15 13 10 11 9 7 13 13
8 7 13 13 1 10 9 10 9
10 9 16 0 13 13 1 15 10 9 0
6 13 3 15 10 9 13
5 15 3 13 0 13
8 13 10 9 15 1 10 9 15
21 10 3 11 13 15 3 1 10 9 10 9 7 13 3 13 1 10 9 13 10 9
19 13 15 1 10 9 10 13 16 15 13 16 15 13 10 11 10 9 10 9
4 15 3 13 13
4 3 13 15 13
2 15 13
6 15 13 10 9 10 0
10 15 13 13 15 11 7 11 10 13 11
7 15 3 13 11 10 13 11
6 7 13 15 10 9 13
7 0 13 16 13 10 9 15
2 15 13
11 1 3 10 0 9 13 10 11 9 0 13
32 7 13 10 9 10 11 13 15 9 0 7 13 15 1 10 0 15 9 15 13 1 10 9 7 13 9 0 10 9 10 9 13
1 13
7 13 3 16 11 10 13 13
1 13
8 15 3 13 10 9 13 3 13
5 9 13 1 10 0
19 7 13 1 0 10 9 13 11 1 11 10 11 7 13 1 10 11 1 11
3 13 3 9
4 9 0 1 9
14 7 3 0 3 13 13 7 13 1 0 9 7 3 13
1 13
10 7 13 10 11 10 9 15 13 10 0
2 15 13
20 7 13 13 15 1 10 9 15 7 0 9 7 9 13 10 11 7 10 9 15
5 7 13 15 10 11
1 13
16 7 13 10 9 15 16 9 13 15 1 10 9 16 3 13 15
4 7 13 1 9
26 7 3 13 15 1 10 9 10 0 13 10 9 15 13 16 3 0 10 0 13 7 3 10 9 15 13
8 7 13 10 1 15 3 13 13
20 7 15 13 1 10 0 3 3 13 9 0 7 3 13 1 10 3 13 9 9
3 7 13 15
8 7 13 0 7 16 13 1 0
13 3 3 13 10 9 3 13 10 9 16 13 10 9
4 3 3 13 9
8 13 10 9 10 0 1 10 9
27 7 13 10 9 10 0 13 1 10 9 7 13 10 9 1 10 9 1 10 9 3 12 7 13 1 10 9
21 7 13 10 11 1 10 9 1 10 3 3 13 9 0 1 15 7 13 1 10 9
7 13 10 9 13 15 7 13
10 10 3 11 13 10 9 13 13 10 9
5 8 8 15 13 13
10 3 0 0 7 15 10 9 10 13 0
7 13 3 10 11 10 11 16
2 15 13
3 7 13 15
3 7 13 15
31 7 13 10 12 9 7 10 12 9 13 1 10 9 13 7 13 10 9 7 13 10 9 16 13 15 7 10 12 9 13 15
6 15 3 15 13 7 13
30 7 3 3 13 1 9 7 1 9 7 1 9 1 10 9 13 10 13 7 13 15 16 7 3 10 9 10 9 15 13
11 3 13 10 9 10 9 16 10 9 15 13
8 10 3 9 13 0 9 10 9
17 7 13 1 10 9 15 13 10 9 13 1 10 9 7 10 9 13
18 1 0 10 9 3 0 9 13 7 3 13 15 13 13 10 9 13 15
8 7 13 10 9 13 1 10 9
6 7 13 10 9 15 13
4 7 13 13 15
1 12
5 3 1 10 9 13
8 15 3 13 9 9 10 9 15
11 7 13 9 13 15 7 13 9 1 10 9
8 7 3 13 1 10 9 10 9
5 15 3 13 15 13
13 7 3 7 1 9 15 13 7 1 9 16 13 15
6 7 13 7 0 13 13
4 7 13 1 11
4 13 15 10 11
5 15 3 13 13 15
3 7 13 15
15 15 3 3 13 10 9 10 9 3 9 3 3 13 1 15
2 3 13
8 15 3 13 1 10 9 13 13
5 13 15 10 11 13
13 7 13 3 10 12 13 15 13 10 13 15 13 16
14 13 13 10 9 15 15 13 7 10 9 15 15 13 13
2 13 15
5 10 3 11 13 15
7 7 15 10 3 13 13 15
14 7 13 15 3 3 13 10 9 13 1 11 1 10 12
6 15 3 13 15 9 9
3 13 9 9
15 13 15 12 9 7 13 15 7 13 15 1 15 9 0 13
5 7 13 10 11 13
10 13 7 13 10 9 7 13 10 9 15
14 3 3 13 1 9 9 7 1 9 10 9 10 9 13
1 9
6 7 10 12 3 13 9
2 0 13
5 7 13 15 10 9
14 13 1 0 15 16 3 13 10 0 15 9 10 9 15
7 15 3 1 10 13 15 13
19 13 15 1 9 7 1 9 13 7 1 9 7 9 13 1 15 1 9 15
6 13 3 16 3 13 9
19 7 3 13 10 9 7 13 10 0 1 10 12 9 1 9 9 1 9 9
7 3 13 3 3 10 9 13
21 7 13 15 1 11 1 10 9 11 10 0 13 15 13 9 13 9 9 9 0 0
13 3 3 10 0 13 1 15 7 3 13 13 3 13
9 7 13 12 10 9 15 7 13 15
2 3 15
5 7 13 15 10 11
20 7 13 0 13 1 10 9 7 13 16 16 0 13 13 1 15 10 9 7 13
6 7 13 13 15 3 13
28 7 3 3 15 13 13 11 10 11 12 10 12 7 1 15 9 1 9 7 9 1 10 9 7 10 9 7 0
5 7 16 13 10 9
14 15 13 10 9 0 10 0 7 1 12 9 15 0 13
8 10 3 9 13 10 9 15 13
4 15 3 13 13
6 7 13 15 10 9 0
9 13 3 16 1 9 13 15 10 9
20 10 3 11 13 13 10 0 10 9 13 15 10 11 7 13 10 11 13 16 13
5 7 13 15 13 9
2 15 13
1 13
37 7 3 0 13 16 13 9 15 13 9 13 11 10 1 11 0 9 15 3 0 13 13 10 9 10 9 13 13 1 10 11 7 13 10 9 10 11
4 13 3 0 3
3 3 0 13
7 1 0 9 13 7 3 13
5 7 9 13 1 15
17 15 13 11 10 13 1 10 9 7 13 13 1 15 7 13 15 0
7 7 13 1 15 10 9 13
7 3 13 0 16 9 3 13
17 7 13 16 13 10 9 10 11 10 11 13 10 9 1 10 9 15
5 13 9 1 9 15
7 7 3 9 9 13 1 15
36 13 3 3 11 1 10 11 1 9 11 1 10 11 1 9 11 15 13 11 1 10 13 15 1 9 7 9 11 13 1 11 10 13 15 13 0
11 9 1 0 9 7 1 9 9 1 9 9
6 9 9 3 12 9 9
9 7 13 11 9 9 11 1 9 11
11 7 13 15 13 7 13 1 15 10 9 15
50 1 9 3 0 10 9 11 9 13 11 11 10 11 7 13 10 11 11 11 3 10 9 15 13 10 0 7 0 9 7 11 10 11 13 1 9 11 7 11 13 9 9 1 11 10 11 9 1 10 9
6 7 3 13 13 1 15
8 0 15 13 1 9 0 7 9
12 7 3 13 15 1 10 9 0 7 13 15 13
1 13
10 7 15 13 1 10 9 15 13 1 15
4 7 13 1 15
14 7 13 1 11 9 10 11 7 13 13 15 1 10 9
10 7 13 9 1 15 7 13 1 15 13
6 15 13 10 9 10 9
9 13 3 11 11 13 10 9 11 13
7 7 13 10 9 13 15 13
18 7 6 9 13 1 9 9 15 13 13 7 13 15 13 7 13 1 15
15 16 3 13 16 10 9 10 9 9 13 1 10 9 13 9
10 7 13 9 0 11 15 1 10 9 15
15 3 13 10 9 10 9 1 15 10 9 1 15 13 13 13
4 10 0 0 13
16 13 3 10 9 7 10 9 16 1 10 9 13 16 13 13 15
7 13 1 0 10 9 7 13
5 3 13 10 13 15
11 7 16 13 1 15 13 13 15 15 9 13
6 15 3 9 13 13 15
15 3 3 13 9 0 13 9 0 7 3 9 0 13 9 0
3 7 3 13
10 3 3 0 13 16 1 10 9 15 13
11 7 13 1 10 9 10 13 13 10 9 13
20 13 13 11 15 13 7 13 16 0 13 0 13 0 13 0 13 0 13 0 13
3 6 13 15
11 0 13 9 10 1 9 13 7 13 15 13
52 7 6 9 15 13 1 10 9 0 7 13 16 13 1 10 9 10 9 13 9 9 7 13 3 1 10 9 15 13 10 9 13 13 10 9 15 7 10 9 10 9 15 13 7 13 10 9 15 7 13 10 9
3 13 11 13
11 0 3 1 15 13 3 13 13 15 10 9
5 13 3 1 10 9
13 7 0 13 1 10 9 10 0 7 13 13 9 0
12 10 9 15 7 10 9 15 13 3 13 15 13
3 9 9 13
10 15 15 7 15 11 9 10 9 10 0
3 7 13 15
12 7 13 1 0 10 9 13 15 13 15 10 11
7 9 10 9 13 15 7 13
4 3 13 10 9
8 15 3 13 10 9 15 13 13
6 13 3 10 12 13 15
24 13 3 10 12 9 7 10 12 9 13 1 10 9 13 15 7 13 7 13 10 9 13 10 9
33 15 3 13 15 13 15 13 0 13 16 13 10 9 10 9 0 13 7 13 1 10 0 7 9 7 9 7 13 7 10 0 9 13
12 7 13 11 7 11 7 11 13 1 10 9 13
2 15 13
5 13 3 10 9 15
12 15 3 13 0 10 9 1 10 9 15 15 13
12 7 3 13 15 16 10 9 15 13 13 1 11
6 13 3 1 15 10 11
5 15 1 10 9 13
16 1 15 3 3 9 13 7 3 13 15 13 1 10 9 15 13
8 10 3 15 13 13 10 13 15
9 6 10 9 3 3 13 9 1 15
2 3 13
14 1 9 3 9 15 13 1 10 9 0 7 13 15 13
12 13 3 1 10 13 15 7 15 13 1 9 15
6 7 3 13 15 1 9
4 7 15 15 13
8 13 3 10 9 13 13 10 0
6 1 0 15 9 13 15
10 0 10 9 10 13 15 7 9 15 13
11 3 13 1 10 9 11 7 6 0 11 3
6 13 3 10 9 1 15
6 9 0 13 3 15 13
3 6 13 15
12 7 15 15 13 9 1 10 9 10 9 13 15
6 13 3 9 1 15 13
1 13
14 13 10 9 16 7 13 7 13 15 3 13 9 7 9
8 0 3 15 10 9 10 9 13
10 0 10 9 0 15 13 10 9 13 13
57 16 3 13 10 9 0 1 10 9 15 13 10 9 15 13 7 13 13 10 9 7 10 9 13 3 7 13 7 13 13 10 9 10 9 0 1 9 15 3 13 7 1 9 15 3 13 7 13 15 7 10 9 15 1 10 0 13
21 13 3 15 1 0 10 9 13 15 1 10 0 15 10 9 11 13 1 10 9 15
5 13 3 1 10 9
9 13 3 15 10 11 13 7 13 15
2 13 3
5 15 3 13 1 15
5 3 13 15 3 13
17 3 13 15 3 7 3 7 10 13 13 16 3 13 9 13 1 11
6 7 13 13 15 7 13
5 13 16 3 0 13
3 7 0 13
10 13 3 15 9 0 7 13 13 1 15
9 16 3 3 10 9 13 1 15 13
22 13 15 16 3 9 1 10 9 13 1 12 0 13 3 1 12 0 15 3 9 13 9
22 7 1 3 0 9 13 0 10 0 9 13 1 9 3 7 3 13 10 9 15 13 3
7 13 15 3 12 10 0 15
19 7 16 13 13 10 9 13 9 7 9 7 13 12 10 9 13 15 13 0
2 13 13
3 15 3 13
13 7 16 1 10 0 0 3 13 10 15 15 13 15
12 1 3 10 9 10 9 13 7 15 1 15 13
26 9 11 13 15 7 13 11 16 13 10 9 10 9 15 9 7 13 10 9 15 16 13 1 10 9 0
2 13 15
17 3 16 3 10 9 13 1 15 7 3 13 1 15 13 13 13 15
18 13 15 13 7 13 13 15 16 13 7 13 7 1 0 13 7 13 15
15 13 3 1 10 9 3 13 10 9 10 9 13 15 7 13
12 0 3 13 15 0 13 7 13 1 10 9 0
16 15 3 9 13 11 1 11 13 9 7 9 1 9 7 13 0
4 10 3 0 13
6 1 3 0 13 1 15
5 10 9 13 0 13
6 13 3 10 9 13 15
6 15 0 3 3 12 9
9 10 0 1 9 0 1 10 9 13
15 13 3 1 10 13 15 1 11 0 15 13 1 10 9 13
4 15 15 13 13
7 7 15 13 9 7 13 0
7 13 3 1 15 10 11 16
25 7 13 1 10 13 15 13 10 9 7 13 13 15 10 9 0 15 13 10 9 16 13 15 15 13
10 9 6 10 9 15 15 13 13 1 9
3 7 13 15
10 7 15 10 9 1 10 9 13 1 15
7 7 13 10 9 15 9 9
7 15 3 13 1 15 13 16
15 7 9 13 1 10 9 9 16 1 10 9 10 9 13 15
9 13 3 15 10 9 13 1 15 13
10 9 15 13 10 13 0 13 1 9 9
3 13 15 9
7 7 10 0 13 9 13 0
6 13 10 9 10 9 15
12 0 3 1 10 9 15 0 10 9 15 13 13
4 3 13 1 15
17 15 3 13 15 9 7 9 15 3 13 13 7 13 0 10 13 15
15 7 3 13 10 9 10 9 13 1 9 1 9 7 9 0
11 13 3 1 15 10 13 1 9 15 10 9
11 7 13 7 13 9 10 13 15 1 9 15
12 3 13 10 9 3 10 9 1 10 9 15 13
4 15 3 13 15
11 15 3 13 1 15 16 3 13 10 9 15
1 15
11 7 13 13 1 10 9 1 10 9 10 9
18 7 13 1 10 9 13 1 10 9 13 13 15 1 10 9 7 13 15
3 13 1 0
5 3 0 1 15 13
4 13 3 10 11
7 0 3 13 1 10 9 15
20 15 3 13 13 16 13 10 9 13 1 0 10 11 7 13 1 10 11 1 3
14 11 3 13 10 9 7 10 9 7 10 9 13 1 15
9 3 3 10 11 13 13 13 10 11
12 13 3 10 1 9 7 9 13 1 9 15 13
3 7 10 9
5 13 3 10 9 13
7 13 3 10 0 13 15 13
26 0 13 10 11 13 10 9 10 11 7 13 13 15 9 7 13 15 1 9 0 3 3 13 15 3 13
14 0 3 13 15 7 13 10 9 1 10 9 13 1 15
9 10 3 9 15 13 10 3 13 15
11 15 3 13 16 15 13 10 13 13 10 11
12 7 13 1 10 9 3 13 7 15 13 3 13
16 7 15 13 10 1 10 9 7 3 13 15 1 10 9 10 9
5 7 13 1 15 13
17 1 9 13 10 9 7 10 9 13 1 10 9 7 9 13 10 9
4 9 15 13 3
2 3 13
9 13 10 9 9 3 13 11 10 9
11 13 10 9 10 9 10 13 10 9 10 9
5 13 10 9 10 9
17 13 11 10 9 11 11 12 1 10 12 10 13 1 11 7 13 15
12 13 3 10 11 1 11 1 10 9 11 7 11
3 3 15 13
6 13 10 9 15 10 9
12 15 9 0 10 0 9 13 7 3 13 10 0
7 13 3 10 0 7 13 15
8 15 3 13 15 13 1 10 9
12 3 13 1 10 9 10 9 15 0 13 7 13
4 3 13 0 13
16 10 3 13 3 13 16 3 13 1 10 9 10 0 9 10 9
19 9 15 13 1 15 1 10 11 15 15 13 13 0 13 7 15 13 1 15
18 13 3 1 9 10 11 13 11 1 10 9 15 13 11 11 10 9 15
5 13 11 7 13 15
13 9 13 15 0 10 9 16 3 13 7 13 3 13
4 13 15 10 9
12 9 10 9 7 10 13 1 9 7 9 13 13
9 6 13 9 15 13 15 15 15 13
15 15 9 13 16 13 10 9 10 13 15 7 13 15 10 9
12 16 3 13 1 15 10 9 13 15 13 1 15
4 10 9 15 13
16 13 3 1 10 11 1 10 0 9 10 13 3 11 12 9 13
6 13 10 9 15 7 13
3 13 7 13
26 1 0 3 13 15 10 0 13 16 3 0 13 10 9 7 7 9 0 13 10 9 0 15 13 10 9
24 6 6 13 15 16 13 9 7 3 13 3 10 0 13 10 9 10 9 10 9 7 10 13 13
14 15 3 3 1 9 10 9 13 7 0 13 16 15 13
17 9 1 9 3 13 7 13 15 16 3 13 10 9 10 9 1 15
11 13 9 3 15 13 12 9 0 7 12 9
9 10 3 9 13 15 13 9 13 16
18 13 3 13 15 1 10 9 7 3 13 10 9 1 10 9 1 15 13
7 0 3 10 9 13 10 9
5 13 3 15 10 11
36 15 15 13 15 10 9 1 15 13 7 10 13 1 15 3 3 13 3 16 13 1 10 9 3 16 13 10 9 10 15 7 10 9 10 13 15
22 15 13 13 1 15 16 3 10 9 10 13 15 13 15 7 15 13 15 1 10 0 9
17 0 13 10 9 10 1 10 9 13 16 15 1 15 13 7 3 13
3 0 15 13
6 13 3 10 11 10 12
10 0 3 13 15 13 12 13 1 10 12
6 10 9 10 15 3 13
9 7 9 13 1 15 0 1 10 9
20 16 15 13 10 9 15 13 13 1 10 9 3 1 9 13 7 15 1 15 13
6 12 9 13 7 15 13
9 10 3 11 3 13 15 13 3 13
13 0 3 13 1 10 9 15 13 13 10 13 1 15
14 15 3 13 1 15 13 15 7 15 13 1 15 10 9
17 3 10 9 15 13 10 9 16 3 13 0 1 15 7 13 15 13
4 15 3 15 13
3 15 3 13
6 10 9 15 3 13 0
5 3 13 10 9 15
5 3 13 15 16 13
7 0 15 13 0 13 1 15
6 10 9 13 1 10 9
16 3 3 13 15 13 9 15 10 9 15 13 15 13 1 10 9
8 1 15 10 9 10 15 3 13
6 13 10 0 7 13 15
8 11 13 7 10 9 7 15 13
4 15 3 13 15
8 11 3 13 7 13 1 10 9
6 3 3 13 15 10 9
16 13 3 9 1 15 9 10 9 13 10 11 7 13 15 10 9
10 15 15 13 1 15 16 13 15 10 9
4 15 1 15 13
5 3 0 13 3 13
4 15 9 13 0
9 1 9 15 13 0 7 15 13 15
3 7 13 15
13 15 15 13 9 13 7 9 7 3 13 15 10 9
11 3 15 9 13 15 3 13 1 10 9 0
2 15 13
5 13 15 7 3 13
4 13 15 10 0
18 7 13 3 1 10 11 1 10 9 3 13 11 10 0 13 7 13 3
13 13 3 10 11 10 11 7 10 9 15 7 10 11
7 0 13 7 1 0 13 15
4 13 15 10 11
16 15 13 16 15 13 10 11 10 9 10 9 10 1 10 9 13
2 13 15
3 13 10 9
13 7 1 10 9 10 13 13 16 13 16 15 15 13
21 16 13 15 3 15 13 1 15 7 13 10 0 7 13 15 7 10 9 7 10 9
19 10 3 11 1 12 9 10 9 13 1 11 3 13 11 15 13 1 0 11
7 10 0 3 3 13 1 15
8 13 11 7 11 7 13 10 11
7 9 13 15 1 10 9 0
6 3 9 13 10 9 0
12 16 10 9 13 13 1 10 9 16 9 9 13
5 11 3 13 7 13
34 1 3 10 9 10 9 13 10 11 16 13 15 10 9 16 13 1 10 9 0 1 10 9 13 10 0 10 1 10 9 1 9 13 15
9 3 3 13 15 10 9 1 10 9
4 3 15 0 13
10 0 13 11 13 10 9 7 13 7 13
10 13 3 10 9 13 7 13 11 11 11
17 16 10 9 13 1 15 3 10 9 13 15 1 15 7 3 13 15
3 13 3 0
9 1 10 9 10 9 15 9 0 13
7 7 3 13 15 7 13 15
10 10 3 9 1 15 13 13 10 9 15
11 15 13 15 16 1 15 13 7 1 15 13
5 13 16 15 13 15
20 15 9 1 15 3 13 9 13 15 7 15 10 9 13 13 15 16 9 0 13
9 3 13 15 10 9 7 15 13 15
6 0 13 15 16 13 15
9 3 3 9 3 13 1 10 9 15
13 7 13 9 16 15 10 13 15 13 9 13 10 9
7 16 3 13 13 15 1 15
18 15 13 0 15 13 15 0 7 3 13 15 7 3 0 7 13 15 7
5 0 1 9 13 15
3 13 15 11
24 13 15 10 9 16 10 9 13 15 3 13 15 9 15 9 16 15 15 13 15 13 15 9 0
14 7 10 15 15 15 13 7 10 15 15 7 13 1 15
13 3 15 13 1 10 9 7 15 13 15 1 10 9
18 13 3 7 11 10 13 15 10 9 16 3 13 11 3 1 10 9 15
4 3 3 15 13
6 13 3 9 10 9 11
19 15 3 13 1 9 7 1 10 9 3 15 10 0 13 7 1 0 13 15
7 13 3 11 11 13 7 13
3 13 3 3
13 16 10 9 10 11 13 15 13 13 15 9 13 13
10 10 9 10 15 3 13 1 10 9 0
3 15 13 9
5 13 10 9 10 0
4 13 15 10 11
4 9 13 3 0
6 3 13 9 3 3 9
4 9 13 10 0
24 13 3 1 10 9 10 11 10 9 15 7 10 9 10 9 15 11 10 10 11 7 11 10 9
6 16 3 13 10 9 13
4 13 1 15 13
12 13 10 9 1 10 9 7 3 13 3 13 15
29 16 3 13 13 1 10 9 7 13 12 9 1 0 13 12 1 10 9 7 12 1 10 9 3 13 10 9 10 11
14 13 1 10 9 15 7 9 15 7 9 15 7 9 15
3 13 9 0
2 9 15
13 1 0 13 15 3 11 10 9 1 10 9 10 11
4 13 3 15 11
7 10 3 0 9 10 9 13
13 13 11 7 13 10 9 7 13 15 7 10 9 3
2 13 15
6 9 15 13 10 13 15
29 10 3 0 9 13 1 15 6 11 15 13 10 11 13 7 7 13 1 15 9 13 10 9 1 9 0 15 13 13
21 7 16 13 13 1 10 9 13 15 7 6 9 12 13 15 1 9 0 15 3 13
20 0 3 3 13 9 1 9 10 9 7 0 13 13 0 7 13 15 10 9 15
19 7 13 3 1 10 9 9 3 13 9 0 7 13 0 10 9 3 13 13
8 0 3 13 13 16 9 13 13
6 16 13 9 9 10 0
7 13 15 9 1 10 9 15
29 3 15 3 10 13 13 1 10 15 7 13 0 0 7 10 9 7 10 9 13 7 13 15 15 3 3 15 9 13
6 9 7 9 3 13 15
29 15 3 10 0 7 0 13 7 13 9 9 13 15 10 3 9 10 9 13 15 10 9 13 1 0 15 15 9 13
17 7 15 3 10 9 1 11 7 10 3 15 13 3 13 10 9 0
50 9 10 9 7 0 16 15 3 13 1 9 9 0 1 15 0 13 0 13 15 15 7 15 10 9 11 16 1 10 9 11 11 10 0 15 15 13 15 10 9 13 1 0 1 0 0 13 1 15 0
9 10 3 11 7 11 13 13 1 15
37 13 3 1 9 1 10 9 0 1 10 0 9 15 11 15 13 11 7 7 11 11 1 9 7 9 11 13 15 10 9 15 7 10 9 15 13 13
4 13 3 10 11
8 7 13 3 0 1 10 9 11
5 13 3 13 13 16
9 9 13 15 3 13 1 10 9 0
11 9 9 13 15 1 10 9 0 15 13 13
15 15 3 3 13 13 1 9 10 9 16 13 1 10 9 13
14 11 3 0 9 7 9 13 9 7 9 0 1 10 9
4 3 0 3 13
5 7 13 15 9 9
13 10 7 13 9 13 15 13 7 13 15 1 9 13
13 15 10 9 10 9 15 10 9 11 7 11 7 11
11 9 15 13 10 9 1 10 9 15 3 15
64 10 9 10 9 13 10 9 15 1 10 0 3 13 10 13 10 11 13 15 1 10 9 15 13 15 3 13 13 10 9 15 1 11 1 10 9 10 9 15 13 10 9 1 9 10 9 15 1 10 9 11 15 13 9 1 10 9 7 13 13 9 10 9 11
8 15 10 9 3 13 10 9 15
7 9 3 13 15 10 9 0
20 13 3 10 9 10 13 1 10 11 3 1 10 13 15 7 13 10 9 15 13
29 13 3 10 1 11 9 16 13 10 11 10 9 10 9 13 1 15 11 7 11 15 13 13 1 15 16 13 9 0
20 7 6 9 9 9 9 11 9 9 15 13 1 15 10 9 15 13 13 1 11
19 3 9 1 9 13 7 3 9 1 10 13 15 0 3 3 13 10 9 15
4 15 13 15 13
3 15 13 9
1 11
20 13 16 9 9 13 15 0 10 13 10 9 15 1 9 7 7 9 9 7 11
10 16 3 13 9 0 13 10 0 13 15
13 13 3 10 9 13 15 1 11 7 13 15 1 11
6 13 3 15 9 13 15
13 7 3 13 9 1 11 7 13 11 15 15 13 11
7 7 9 3 1 0 1 15
3 15 3 13
8 7 13 15 13 7 13 13 0
10 13 3 1 11 7 13 11 15 13 11
30 11 10 1 11 16 13 15 10 9 9 0 7 9 15 13 13 7 13 15 10 13 1 10 9 16 10 9 13 1 15
19 3 10 9 13 13 15 10 3 13 0 15 10 9 10 0 13 3 3 15
23 13 1 11 7 13 11 10 13 11 15 13 9 1 15 1 15 13 15 7 15 10 9 15
6 7 13 9 9 1 15
4 15 13 1 11
11 7 6 9 9 13 7 9 13 1 10 9
4 13 3 9 13
5 15 3 13 3 13
21 11 3 13 15 7 3 13 13 10 9 13 13 7 13 1 10 11 1 10 11 13
12 13 3 15 10 9 7 13 13 10 9 10 0
53 10 9 10 9 0 11 13 10 9 15 7 10 9 13 1 10 9 1 9 11 7 1 9 0 13 15 1 15 7 3 0 9 13 15 1 10 0 7 13 9 12 1 9 11 13 10 9 15 3 9 12 7 12
32 10 3 13 1 11 7 10 9 15 0 13 7 10 9 10 9 10 1 15 9 13 13 13 7 15 9 9 13 13 11 13 15
5 3 3 1 0 13
14 10 3 13 9 3 15 10 9 13 13 10 9 10 9
12 15 3 13 10 9 10 9 1 15 13 1 11
18 0 13 10 11 13 15 13 15 7 13 16 13 9 10 13 13 0 9
13 15 1 10 13 9 13 15 10 9 13 10 9 15
17 7 3 13 1 11 3 13 13 10 9 10 9 1 10 9 15 13
14 11 13 3 0 10 9 13 13 1 9 9 10 9 15
46 16 13 16 15 1 15 13 13 15 9 13 10 9 15 15 3 13 13 15 13 3 13 9 13 1 15 1 10 0 15 11 7 11 9 13 10 9 15 1 10 9 10 9 15 11 11
8 1 3 15 9 13 1 11 11
9 13 3 0 10 9 15 16 9 13
25 13 3 1 11 13 1 11 10 3 13 1 0 9 7 3 1 11 15 13 0 10 9 11 9 9
6 0 3 13 1 0 9
11 3 3 9 13 0 16 13 10 9 10 9
14 7 13 15 10 9 10 9 1 15 10 1 10 9 15
14 3 13 3 15 13 11 7 15 9 1 10 9 13 16
24 10 3 13 10 11 13 1 11 7 13 9 1 10 11 7 10 11 16 3 0 13 1 15 13
8 13 3 15 13 1 10 9 15
8 1 15 3 13 7 13 7 13
9 1 0 13 1 10 11 13 1 11
20 7 13 3 13 1 9 15 9 11 11 13 10 9 15 10 9 13 13 10 9
6 7 13 15 1 10 9
24 0 13 13 10 9 10 9 7 13 10 9 13 7 13 3 10 1 10 11 13 0 10 9 11
18 13 3 1 10 9 13 1 9 12 13 7 13 10 1 10 9 10 9
27 7 13 10 9 1 15 1 15 13 10 9 10 0 13 0 13 1 15 16 0 7 13 13 1 10 9 0
40 9 13 16 1 0 10 9 10 9 15 13 7 13 7 13 16 3 0 11 7 3 15 10 11 10 11 0 13 13 0 9 13 16 3 13 9 10 1 9 13
10 1 3 10 9 13 11 13 15 10 0
11 16 3 15 1 0 13 1 10 0 9 13
6 13 7 10 9 1 9
12 16 3 13 15 1 10 11 13 15 13 1 11
34 7 3 6 13 15 10 9 13 1 11 10 1 15 13 15 3 13 1 16 10 9 10 0 1 9 13 15 13 16 9 7 9 15 13
19 13 3 10 9 13 3 9 12 15 10 11 13 1 10 9 3 13 1 11
6 3 13 10 11 7 13
6 15 3 13 13 10 9
19 1 3 10 13 9 15 13 13 13 15 10 7 0 7 9 7 0 7 9
19 3 13 10 9 13 15 7 13 13 9 12 7 13 15 13 7 15 13 13
22 3 3 15 13 10 0 10 1 0 10 9 13 7 13 1 10 0 10 12 9 10 9
34 15 13 9 0 13 1 11 10 11 13 3 1 10 9 0 1 10 9 11 13 1 9 10 0 9 9 13 10 9 3 15 15 13 3
9 10 3 1 15 13 10 3 9 13
8 13 16 15 1 9 3 13 15
6 13 3 10 9 13 15
31 10 3 3 13 13 10 0 10 15 13 1 10 0 13 15 7 13 13 10 9 7 15 10 9 7 13 10 11 13 1 15
6 3 13 9 16 13 9
7 3 3 9 13 15 7 9
11 15 3 1 10 13 15 0 13 10 13 15
5 15 3 3 13 15
17 10 3 3 9 1 10 13 15 13 10 11 13 1 9 1 10 11
7 3 3 0 15 13 13 15
12 10 11 3 13 10 0 9 13 13 10 11 13
15 9 3 13 15 11 10 9 7 11 13 1 11 13 10 11
6 13 3 0 10 9 13
6 11 3 1 10 11 13
5 15 3 13 1 11
4 10 3 9 13
3 10 3 11
15 7 3 13 10 9 9 0 13 1 10 11 13 15 1 15
19 9 3 15 13 13 11 13 3 0 13 10 9 15 13 9 13 13 10 9
15 9 15 13 13 7 6 13 15 10 9 15 10 13 1 15
12 3 13 10 9 10 9 10 9 7 13 15 13
8 16 3 9 13 10 9 3 13
9 10 7 0 13 3 10 13 9 15
28 0 3 13 3 10 0 10 1 10 9 13 9 13 7 13 15 3 0 9 13 15 7 13 13 10 1 10 9
10 1 0 3 10 9 13 15 13 7 13
41 9 3 15 13 10 9 15 13 1 10 9 15 1 10 9 10 9 15 16 3 9 15 13 3 1 10 9 15 13 16 3 3 13 1 10 9 10 9 13 1 15
27 13 3 9 9 1 9 1 15 9 7 9 9 10 10 9 1 9 13 16 10 0 10 9 0 13 1 15
23 15 10 9 10 9 13 16 10 10 0 13 0 9 13 3 0 15 13 7 3 13 10 13
16 9 7 9 1 15 9 9 10 13 10 0 0 7 0 7 9
5 10 13 3 13 13
23 7 10 1 10 0 0 7 9 9 1 9 3 9 15 10 9 3 1 9 7 1 10 9
13 16 3 13 1 10 9 15 7 13 1 10 13 15
2 15 3
24 13 3 16 15 10 9 13 10 1 10 9 13 16 15 9 13 7 0 13 15 10 9 10 9
3 1 15 9
8 16 3 11 1 9 13 13 9
3 3 3 13
5 9 0 9 13 15
21 10 3 9 3 13 16 10 9 10 9 13 1 10 9 15 1 9 0 10 13 15
7 9 3 3 13 3 13 9
7 9 3 13 16 13 10 9
21 3 13 16 15 13 15 9 1 9 9 13 15 13 7 9 1 9 7 9 1 9
13 10 3 9 10 9 9 0 1 11 11 10 9 15
3 10 9 9
6 10 3 0 15 13 9
11 10 3 13 13 15 10 3 13 10 0 3
8 15 3 3 9 10 1 11 11
15 15 3 3 13 1 9 7 1 9 16 9 9 13 1 15
11 0 10 9 13 10 9 15 16 13 9 9
5 15 3 13 1 0
4 13 3 9 9
5 9 3 10 9 0
4 10 11 3 13
10 6 9 3 15 15 13 10 13 10 9
6 11 3 13 1 10 11
5 13 10 9 10 9
5 15 13 1 10 9
8 3 0 10 9 10 13 10 0
4 3 11 3 13
7 3 13 10 9 10 9 15
12 16 3 9 3 1 9 16 10 9 3 13 9
4 3 13 16 13
12 16 3 13 3 15 10 9 13 7 10 9 15
9 1 3 15 9 9 16 13 10 9
7 1 3 10 9 0 1 15
6 16 10 13 1 10 9
3 10 9 13
3 13 1 13
2 15 13
6 10 3 13 15 9 13
6 1 0 3 3 9 13
7 10 9 10 3 0 3 13
10 10 3 13 10 9 13 3 1 9 9
10 16 7 3 13 16 7 13 10 9 13
4 3 3 15 13
8 3 1 9 13 10 9 10 9
3 7 3 13
2 7 3
14 3 3 13 13 3 3 13 11 16 3 1 0 9 13
11 13 3 16 13 1 15 1 9 9 11 13
7 13 9 10 0 15 1 9
15 13 15 9 10 0 15 7 9 7 9 7 9 10 0 15
16 0 10 9 1 15 13 1 9 10 9 15 11 11 10 9 15
20 13 16 15 15 13 3 3 11 7 11 16 3 15 13 16 1 10 15 9 13
5 3 9 10 9 0
46 7 15 1 9 7 1 9 7 1 9 0 13 1 15 7 10 9 15 7 10 9 15 3 1 0 9 9 7 1 9 9 7 9 16 10 9 15 3 13 1 9 9 7 1 9 9
16 15 3 13 9 0 10 9 3 3 10 9 10 9 10 1 15
16 7 15 9 3 13 13 15 3 0 7 3 0 3 0 1 11
2 15 13
3 15 15 13
3 15 3 11
29 0 3 9 13 1 15 7 11 1 15 16 1 15 13 10 3 1 15 13 16 3 12 1 10 12 13 1 10 0
4 15 0 1 11
9 3 9 10 9 13 15 9 1 3
2 15 13
8 13 15 1 10 9 3 13 9
11 7 16 1 15 13 10 9 0 13 9 0
9 10 9 10 9 7 10 9 10 9
3 13 10 9
7 3 3 3 10 9 10 9
6 0 3 13 13 3 13
7 1 3 9 13 15 10 9
2 9 13
15 13 3 0 0 13 1 10 13 9 16 0 9 10 3 13
5 9 10 9 13 13
3 10 9 13
11 13 3 16 10 9 15 0 9 13 10 0
10 10 3 9 15 10 9 15 13 1 9
4 3 13 9 13
9 3 13 3 0 16 3 13 1 15
12 0 3 13 1 15 15 15 13 16 10 0 13
7 15 3 3 13 3 3 3
2 3 13
4 16 0 15 13
8 15 10 15 13 7 10 10 0
7 9 15 13 3 3 15 11
13 9 3 3 3 13 13 10 9 9 7 9 9 13
21 7 10 9 0 13 15 16 9 3 16 13 9 15 13 9 3 16 13 9 15 13
3 15 13 15
22 3 15 3 13 10 9 7 13 10 9 10 9 3 0 13 10 9 7 10 9 10 9
14 13 16 16 9 13 1 10 9 10 0 3 3 13 13
10 7 3 10 9 3 13 12 9 7 0
30 7 0 3 10 13 9 10 9 0 13 0 13 7 15 13 0 13 10 9 0 9 0 13 7 10 0 15 9 0 13
3 3 15 9
3 13 10 9
2 15 13
6 16 13 0 13 3 0
3 13 10 9
27 3 3 9 16 13 1 15 9 13 15 15 13 16 3 15 13 7 1 9 7 1 9 7 1 9 7 9
19 7 1 9 13 12 9 10 9 15 13 16 3 0 13 3 12 9 1 9
4 15 3 13 9
10 9 3 12 7 12 13 7 10 0 13
14 16 15 13 9 13 7 0 13 15 13 15 16 9 13
19 15 3 13 10 0 10 9 15 3 13 0 13 9 16 13 10 9 10 9
7 3 3 10 13 1 11 13
5 0 0 13 10 9
3 3 3 13
3 13 1 9
6 10 0 11 1 9 13
12 15 3 13 1 0 1 9 9 1 10 0 9
24 3 9 15 0 0 13 0 13 1 10 9 10 9 3 13 16 10 9 15 3 13 0 1 9
7 13 3 1 11 1 10 9
1 13
14 13 15 1 9 0 11 7 11 1 10 1 9 15 9
44 0 10 9 3 9 10 9 15 11 11 10 9 10 9 3 9 15 9 10 13 15 1 15 10 9 15 1 10 13 15 13 10 1 15 9 1 10 9 15 13 0 1 10 9
12 3 16 13 15 10 9 7 0 13 10 9 15
6 15 3 15 13 3 15
9 7 3 1 9 1 9 1 11 13
15 16 3 10 9 10 9 9 0 3 13 10 9 10 9 9
21 15 3 15 13 9 10 9 9 13 10 15 9 13 1 9 1 9 3 1 9 9
5 10 3 9 1 15
15 10 3 13 15 1 15 0 9 10 13 15 10 9 10 9
4 16 3 13 9
59 15 1 15 13 9 16 3 13 10 9 7 1 15 13 15 3 9 9 1 9 0 1 9 1 9 1 9 1 9 1 9 1 9 1 9 1 9 1 9 1 9 1 9 1 9 1 9 1 9 0 1 9 0 1 9 9 1 9 9
6 7 15 9 9 1 9
2 13 15
16 7 3 13 15 1 11 15 13 9 10 9 15 7 1 15 13
8 1 15 13 15 0 13 10 9
27 7 3 1 15 13 9 7 9 7 9 7 15 9 7 10 1 15 1 15 9 3 3 1 0 10 9 13
11 10 10 0 3 13 7 10 10 0 3 13
22 13 3 10 9 15 15 1 15 13 9 16 11 13 1 3 7 10 15 9 13 10 0
4 10 1 9 13
10 1 3 3 15 13 1 10 9 10 11
7 13 3 15 13 10 3 9
20 15 3 13 3 13 16 13 10 9 10 13 9 16 1 15 13 13 3 3 15
8 16 0 13 1 9 3 15 13
2 3 15
41 9 3 9 9 9 9 9 1 9 9 1 9 9 1 9 9 1 9 9 1 9 9 1 9 9 7 9 1 9 3 1 9 7 9 1 9 3 1 9 7 9
27 13 9 1 11 1 9 12 7 1 9 3 13 7 1 10 9 3 13 10 9 13 13 10 0 1 0 9
17 15 3 13 15 13 1 10 0 9 3 3 16 0 15 3 13 15
10 3 15 15 13 1 15 1 15 13 15
9 1 9 12 9 7 12 13 15 9
26 13 3 1 10 9 3 13 15 0 15 3 16 15 0 13 7 16 15 10 0 13 15 3 3 0 13
10 7 10 9 10 9 7 9 13 1 15
9 16 15 15 13 1 15 13 9 13
11 15 3 13 15 6 1 10 9 16 3 13
10 7 3 11 10 1 15 9 13 13 13
4 13 3 3 15
3 0 13 3
16 16 3 1 9 15 13 1 10 9 0 16 10 0 1 9 13
8 10 3 11 1 9 13 10 9
12 3 10 9 9 15 13 1 11 16 1 9 13
24 1 15 9 10 9 0 13 15 13 9 9 15 13 7 1 9 13 7 9 1 10 9 10 9
7 13 15 16 3 13 1 15
26 9 15 15 3 13 16 15 13 11 1 15 13 3 13 1 15 3 7 13 10 9 15 16 13 1 15
9 3 9 3 13 9 9 7 10 0
2 13 3
14 0 3 10 9 1 9 10 9 7 1 10 9 13 15
15 10 3 9 10 9 13 9 9 9 9 9 9 9 9 9
11 13 3 10 13 10 9 10 13 1 15 0
17 15 13 13 1 9 0 13 15 13 0 16 10 9 10 11 3 13
130 0 10 9 7 9 10 9 15 11 11 10 13 15 1 15 9 0 1 10 0 1 11 3 13 15 1 15 1 9 9 13 15 0 7 0 1 15 1 9 13 15 1 9 1 11 11 1 15 1 10 9 10 9 15 1 9 9 10 9 15 15 13 15 1 10 13 1 15 13 10 9 1 10 9 15 10 9 10 9 1 10 9 10 9 15 15 13 1 15 1 15 9 7 9 13 15 10 9 10 9 15 1 10 9 15 15 13 1 15 1 9 10 9 10 9 13 10 15 1 10 11 10 1 10 9 7 10 1 10 9
5 7 0 3 1 15
2 3 13
7 10 9 3 13 1 9 15
24 0 3 13 13 16 15 9 7 0 7 9 15 13 9 3 13 9 1 10 9 10 11 7 9
8 10 3 15 13 1 10 9 13
12 3 13 10 9 13 10 15 9 3 10 15 9
23 13 10 9 15 7 10 9 15 13 9 0 1 9 16 3 15 13 7 13 0 1 10 9
39 16 3 3 15 13 10 1 15 15 13 15 13 15 11 10 0 9 7 0 9 1 9 15 13 1 15 1 0 0 16 13 10 1 15 7 13 10 9 15
7 15 3 7 1 9 7 9
40 3 3 10 9 15 13 7 13 15 10 9 10 1 15 9 16 1 10 9 11 15 9 13 0 7 0 7 0 7 15 9 13 16 9 11 11 1 9 9 9
12 0 3 3 13 13 16 3 13 10 1 15 3
3 13 10 9
22 10 3 3 13 10 3 3 13 1 9 13 1 10 9 10 3 9 10 9 1 11 11
24 0 0 13 15 15 1 10 9 13 15 1 3 11 7 10 0 0 15 15 10 9 1 9 9
8 7 10 9 10 9 13 1 15
13 3 3 1 11 7 3 7 3 1 10 9 15 13
7 3 3 10 1 10 9 9
25 3 3 13 10 11 11 10 9 1 15 13 13 7 13 1 15 7 13 10 9 3 13 13 1 9
21 15 13 9 3 13 9 1 9 7 9 7 9 9 3 1 9 15 1 9 10 9
9 3 7 10 11 13 15 3 3 15
7 10 9 13 10 9 1 15
15 10 9 15 3 1 9 9 13 13 3 13 15 12 0 13
3 7 13 11
46 0 3 1 15 13 15 9 13 1 15 7 3 13 1 10 9 1 10 9 13 9 13 7 0 7 13 10 9 15 1 10 9 15 13 1 10 0 11 10 13 15 1 10 9 10 13
67 15 3 9 13 9 10 9 10 9 10 13 1 10 11 1 11 11 16 10 15 13 3 15 1 10 0 9 3 3 0 1 10 0 10 7 10 9 13 11 7 10 9 7 15 13 7 9 3 13 7 15 9 0 13 15 10 9 13 16 13 1 10 13 15 10 9 3
9 1 3 10 9 3 9 13 13 15
7 3 13 15 1 10 9 0
31 3 3 13 15 10 9 1 9 7 1 9 9 1 10 9 15 11 11 10 13 1 15 16 7 13 7 13 3 1 15 13
2 3 13
7 0 10 13 15 15 3 13
47 13 3 15 9 1 10 9 10 9 15 11 11 7 15 9 1 15 1 10 3 3 13 15 1 10 9 7 13 7 1 9 7 1 9 7 1 9 3 1 15 3 16 13 10 9 10 9
17 3 3 9 13 7 13 10 9 15 13 7 1 9 7 1 9 15
17 7 3 16 13 1 15 0 13 15 16 16 15 3 13 13 7 13
20 0 10 9 7 15 9 0 16 11 11 13 1 10 9 0 13 15 0 13 15
17 1 15 13 15 9 7 9 9 13 3 13 9 9 1 9 7 9
3 0 10 9
12 9 13 12 9 9 9 3 13 7 10 0 9
7 10 3 0 7 0 9 13
2 0 13
5 10 3 13 13 13
14 10 3 13 0 0 9 13 3 10 13 1 9 7 9
20 9 3 15 10 0 13 10 9 15 15 13 13 1 10 9 7 15 13 9 0
4 10 9 1 15
11 10 0 9 13 1 9 0 10 13 1 15
3 13 15 13
5 13 3 15 3 13
20 16 3 15 13 15 1 0 13 9 1 9 13 0 10 9 1 15 9 0 13
5 7 3 13 1 0
3 13 3 3
6 13 3 15 0 1 9
24 13 15 10 9 1 15 9 0 7 13 1 10 9 15 10 0 15 10 9 1 10 9 10 9
12 9 7 9 1 9 9 7 11 11 10 9 15
3 9 13 13
3 15 15 13
4 3 3 13 13
26 3 0 1 11 9 13 13 15 10 13 1 10 9 3 13 0 13 3 9 9 3 3 3 9 11 11
7 6 9 15 15 13 1 9
5 13 9 7 13 9
23 16 3 10 1 9 13 9 13 0 7 15 9 7 9 13 0 9 3 15 13 0 13 9
25 10 3 0 15 1 9 13 13 11 1 10 9 10 9 9 7 9 13 16 9 9 1 15 13 9
24 3 13 1 15 10 9 13 16 0 13 7 0 9 10 1 10 9 1 10 13 10 9 10 9
7 3 13 10 9 0 7 13
9 7 3 15 10 13 1 11 1 11
7 13 3 3 1 10 0 3
31 13 3 10 9 10 9 7 0 7 0 1 15 9 0 7 13 1 9 9 7 9 9 7 7 9 7 0 9 7 9 9
35 3 13 10 10 9 10 9 9 1 10 9 13 3 3 9 13 9 1 0 9 7 9 1 9 9 9 9 7 9 9 7 0 7 9 0
15 9 3 1 10 0 13 7 15 15 9 9 1 9 10 9
25 7 0 3 0 13 16 1 10 9 11 13 9 0 15 3 1 9 9 0 13 7 1 9 9 0
28 0 13 9 15 13 1 0 10 9 10 9 1 10 9 10 0 9 7 10 9 10 0 15 13 10 9 3 9
2 13 9
12 13 3 3 3 10 0 9 9 10 7 0 0
12 9 3 1 0 0 16 3 13 16 13 10 13
29 9 3 13 10 9 10 13 0 3 0 10 9 10 9 1 9 10 0 9 15 13 1 10 0 3 13 10 13 13
8 3 3 9 0 3 9 1 9
26 13 3 10 0 9 1 15 13 0 9 13 9 0 3 9 7 7 9 13 0 3 9 10 3 13 13
27 9 0 9 11 1 11 13 10 9 1 15 13 13 0 13 1 10 9 15 10 9 7 1 15 13 3 13
27 3 3 1 12 13 7 0 13 3 10 9 10 9 10 9 7 3 10 9 10 1 10 9 10 9 10 0
16 9 11 13 0 10 9 11 13 7 13 1 10 9 10 9 15
4 7 15 3 13
7 13 9 1 9 10 0 15
17 3 1 9 13 1 10 9 13 7 13 10 9 15 15 3 9 13
5 13 16 13 10 13
6 13 3 1 9 15 13
4 13 3 0 15
10 13 3 9 9 7 3 0 9 13 15
5 15 3 13 10 0
8 10 3 9 0 10 3 13 9
2 3 13
11 3 0 9 13 9 15 13 16 0 9 13
11 3 13 0 10 9 3 13 7 0 0 0
13 13 7 3 13 16 3 13 16 1 10 9 15 13
8 13 3 10 9 7 13 1 15
11 12 13 10 9 7 9 10 13 13 7 13
4 13 3 10 0
3 3 13 15
17 1 15 3 9 15 3 13 7 10 9 7 10 9 7 0 15 9
11 13 3 15 10 9 7 13 1 15 16 13
9 0 3 13 10 9 10 13 1 15
3 15 3 13
12 0 3 9 16 1 9 9 13 15 9 13 3
6 15 3 13 1 9 13
2 6 6
7 10 9 10 1 11 9 13
8 7 10 9 10 1 11 9 13
37 13 3 13 3 10 9 10 11 7 13 10 9 15 7 3 13 10 9 15 1 10 9 11 10 9 15 10 0 15 15 13 1 15 3 10 11 13
12 13 15 10 9 16 9 13 16 13 7 0 13
4 13 15 10 9
8 7 10 9 10 1 11 9 13
25 10 13 13 15 13 1 15 1 10 9 15 3 3 15 13 7 13 1 10 9 15 1 10 9 15
29 7 10 9 10 0 0 9 7 10 0 9 0 9 7 10 0 9 13 10 9 3 9 7 10 0 9 0 9 13
37 7 13 1 0 10 9 7 10 12 9 7 1 0 10 0 9 13 3 13 13 9 12 7 9 12 15 13 10 12 9 10 9 13 1 15 10 9
12 7 16 13 10 9 10 0 13 10 0 9 13
63 7 13 16 13 10 9 10 0 7 9 0 13 7 10 9 0 13 3 9 0 7 10 9 0 13 3 9 7 10 9 10 9 13 1 10 9 3 9 13 10 9 15 1 9 0 13 7 10 9 13 3 9 13 7 15 9 7 9 1 10 9 15 13
33 7 15 9 13 7 13 1 10 9 13 9 0 7 13 15 9 0 16 13 10 9 10 0 15 1 10 9 10 0 10 1 10 9
26 7 13 10 0 10 9 9 7 13 10 0 10 9 10 1 10 9 10 13 9 7 10 0 10 9 13
20 7 1 10 9 13 9 1 10 9 7 13 15 9 3 13 9 10 9 10 9
7 6 13 3 12 9 1 0
72 7 10 0 10 9 15 3 13 1 10 9 0 7 13 1 10 9 10 9 15 16 3 13 10 9 7 10 9 10 0 7 10 0 7 10 0 7 10 0 7 10 0 15 7 13 13 7 13 7 13 7 3 13 1 10 9 15 7 1 10 9 15 7 1 10 9 15 7 1 10 9 15
3 7 13 15
23 7 3 13 10 9 15 10 9 10 13 1 10 9 13 1 15 9 7 13 15 7 13 15
7 6 10 9 10 0 13 0
24 7 15 13 15 1 10 9 10 9 7 1 10 9 10 9 15 7 3 13 10 9 15 1 9
21 7 10 9 15 13 13 0 9 7 10 9 15 3 9 7 10 9 15 3 9 9
10 16 15 1 9 13 13 15 1 9 13
8 10 13 9 13 10 9 10 9
19 0 13 1 10 9 9 10 9 7 10 9 7 1 10 9 15 3 13 9
16 3 10 9 10 0 13 10 13 10 9 10 9 7 10 9 11
17 7 13 10 13 1 10 9 10 9 15 1 10 9 7 13 10 9
10 0 7 0 10 9 15 10 9 10 9
12 6 9 10 9 10 9 0 7 0 10 9 15
1 6
8 7 15 9 13 7 9 3 13
5 7 13 15 10 9
11 10 0 3 13 7 3 13 0 15 13 13
6 7 13 1 0 9 13
11 13 9 7 9 3 13 7 9 3 3 13
34 7 15 9 7 15 10 1 9 13 7 9 7 15 10 9 13 1 3 13 7 13 13 10 9 10 9 15 13 15 0 10 9 10 0
23 1 3 0 9 15 3 3 13 10 9 13 13 10 11 1 11 13 13 10 9 10 9 11
23 15 3 13 0 13 15 11 10 9 16 3 13 15 9 7 13 13 13 15 1 0 9 13
9 1 3 10 11 3 13 9 3 9
15 0 10 11 9 0 15 15 13 15 3 13 9 1 9 9
41 1 0 9 13 13 10 9 1 9 1 9 7 10 11 13 7 11 13 3 1 12 7 7 12 9 9 9 12 7 7 12 9 1 9 13 10 9 1 11 10 11
9 1 3 9 13 13 3 10 9 9
6 13 3 1 10 9 9
8 3 3 3 3 15 13 9 13
11 13 3 10 9 7 13 1 10 1 11 9
19 0 3 10 11 0 9 15 15 13 1 11 13 9 1 11 10 11 11 9
27 0 3 11 7 10 11 0 13 7 9 0 7 1 10 11 13 11 7 10 1 11 13 13 1 11 7 13
13 10 3 9 10 0 13 16 9 3 13 9 10 9
12 16 13 3 10 9 9 13 13 9 11 9 11
24 11 3 16 15 0 13 3 13 9 1 11 13 9 13 11 7 7 0 9 15 3 10 9 13
12 1 3 10 1 0 7 7 11 9 11 3 13
5 13 3 13 15 13
36 13 3 15 15 0 1 10 9 15 3 11 13 10 9 13 1 11 15 3 11 10 0 13 11 16 15 13 0 1 10 11 13 0 13 10 9
58 13 3 0 7 13 11 9 13 1 11 13 9 15 7 10 15 1 10 11 9 15 0 10 9 13 13 3 15 15 13 7 3 3 11 9 0 15 0 9 13 13 13 9 12 1 9 9 13 16 3 3 15 10 9 13 13 15 13
9 11 3 15 13 7 10 13 13 13
3 15 3 13
15 0 3 3 13 13 10 9 10 9 10 3 0 10 9 15
17 1 3 10 0 9 0 3 13 13 15 3 15 13 0 3 3 13
19 10 3 3 0 0 0 3 12 13 10 0 0 0 3 10 0 7 0 0
24 15 3 3 15 0 13 13 7 3 13 3 10 9 0 1 15 10 9 0 6 9 0 13 13
3 13 3 11
14 6 9 9 9 0 13 15 1 10 9 15 10 9 13
15 13 3 0 10 9 13 10 10 11 9 13 15 13 10 9
5 1 3 9 0 13
4 3 3 1 9
9 0 7 3 15 13 7 3 9 13
5 13 3 10 11 9
10 11 3 3 13 3 9 13 10 15 9
16 16 3 3 13 1 10 9 10 0 13 10 0 10 9 13 0
36 13 3 10 11 0 13 1 11 3 0 7 3 15 9 12 9 0 0 7 0 15 10 3 0 13 1 0 13 1 10 9 10 3 0 1 0
16 3 3 3 10 15 9 10 1 10 9 13 10 11 7 10 9
35 16 3 13 10 9 13 10 11 13 7 10 9 3 7 13 13 10 11 9 13 3 1 11 11 13 13 15 10 9 1 9 12 9 0 9
15 0 3 13 10 13 13 10 0 10 3 0 10 3 0 9
16 13 7 16 10 13 9 9 13 1 0 10 9 0 13 1 9
11 13 3 9 7 10 9 10 0 13 13 0
18 13 3 10 9 10 11 13 11 16 13 15 10 9 13 9 1 10 9
16 16 3 13 1 10 11 15 13 1 10 9 3 3 13 1 15
6 13 10 9 1 9 13
21 11 10 9 0 9 13 1 11 1 10 9 16 13 1 10 9 3 10 11 13 0
37 15 3 1 7 9 0 7 9 3 0 9 3 7 13 3 7 13 7 3 15 3 13 9 13 7 13 9 0 13 13 1 11 1 15 10 9 9
21 13 3 10 9 15 15 13 9 7 13 15 13 0 7 9 13 10 9 10 9 13
13 0 3 10 9 11 13 1 11 7 9 13 7 9
19 15 3 13 1 11 7 13 10 15 9 1 10 9 13 1 3 13 10 9
6 11 3 15 13 13 9
13 3 3 9 3 1 0 13 13 1 3 10 0 9
20 9 3 13 7 3 13 10 9 1 9 7 3 15 13 7 3 13 13 15 15
14 10 3 13 15 13 0 11 7 10 9 7 11 10 0
10 3 16 3 13 3 10 9 3 0 13
14 9 3 0 13 7 13 15 0 9 15 13 13 9 13
17 13 3 10 0 7 13 1 9 15 13 13 10 9 3 13 11 13
12 13 3 15 13 10 0 9 13 1 10 11 9
8 9 3 13 15 0 13 10 9
7 13 3 7 15 0 13 0
29 1 3 0 13 10 9 16 3 13 3 10 0 13 9 0 13 13 15 9 13 11 1 0 10 9 15 15 13 9
13 13 15 9 15 3 0 13 10 3 15 0 0 3
18 10 3 9 0 10 0 16 13 13 10 9 1 9 7 7 0 13 9
17 16 3 3 15 13 0 13 7 7 13 1 0 9 1 3 13 11
9 3 15 13 3 13 3 10 9 13
16 1 3 3 15 10 9 10 9 13 1 3 15 10 9 10 9
3 15 3 13
9 11 3 13 15 15 15 0 13 13
25 13 3 11 16 3 1 10 9 10 11 13 10 11 9 7 3 1 0 11 3 0 3 13 13 9
7 13 3 3 10 11 0 9
5 15 3 13 10 9
14 12 3 9 0 0 13 1 10 7 0 9 7 10 0
27 9 3 9 3 0 13 3 9 1 3 16 10 0 9 13 0 3 9 15 15 13 9 9 7 9 13 13
19 10 3 0 10 9 13 15 16 3 3 13 9 10 3 0 13 13 10 9
33 0 13 10 3 11 1 9 12 7 12 0 1 15 9 13 13 7 3 0 1 10 9 13 10 0 13 9 0 7 13 10 9 13
24 3 3 13 15 13 9 10 11 13 0 1 15 9 7 13 7 13 16 15 0 13 9 15 13
14 10 3 15 0 13 9 1 10 11 9 3 3 10 9
6 0 3 1 10 9 13
33 0 13 0 3 13 0 10 9 7 0 7 13 1 9 10 1 10 11 7 0 13 3 0 13 10 7 0 7 10 0 7 10 9
7 0 3 13 13 1 10 0
27 3 3 13 7 10 9 1 0 15 13 7 13 1 15 10 13 1 10 0 9 3 13 15 13 11 10 9
20 3 3 10 11 0 13 3 9 0 9 3 10 15 0 15 13 9 13 10 9
5 13 3 1 15 13
17 9 3 10 9 13 15 13 11 1 10 9 9 1 3 10 0 11
27 13 3 1 9 0 15 1 15 3 10 9 10 9 13 10 3 9 15 15 3 13 10 11 13 15 10 9
16 13 3 13 9 7 7 9 13 3 3 7 9 13 0 1 11
3 13 3 13
13 13 3 1 10 11 13 13 0 13 10 9 10 9
22 12 3 0 10 9 13 13 11 9 9 0 1 9 3 3 3 13 10 13 1 10 11
8 6 9 15 0 0 13 1 9
5 10 3 3 11 13
7 11 3 3 10 0 13 9
5 0 3 13 13 0
13 0 3 13 7 13 10 0 10 9 13 1 10 9
8 7 3 1 15 15 0 13 13
25 3 3 3 13 1 10 9 0 13 13 9 7 15 13 9 13 7 7 9 15 13 1 9 13 9
5 9 3 15 3 13
23 10 3 9 13 10 9 0 16 3 13 10 9 13 15 10 9 13 9 16 13 11 9 13
37 13 3 10 9 10 9 7 9 13 3 9 10 9 10 0 13 1 10 9 13 15 1 9 13 10 9 11 13 9 15 13 7 15 15 0 13 13
12 3 7 13 13 6 9 13 15 13 0 13 9
37 1 3 0 10 7 9 7 10 9 7 10 9 10 11 15 10 9 13 1 15 0 13 7 13 3 13 10 9 9 1 3 9 7 7 9 3 0
20 15 3 13 11 3 1 10 0 10 9 13 9 13 10 9 15 10 9 11 13
11 15 3 10 15 9 13 3 13 7 10 9
18 7 1 0 13 9 10 9 13 13 13 16 15 1 9 13 15 9 0
8 1 3 10 13 15 13 10 9
19 7 3 3 10 0 9 13 10 15 13 0 13 7 1 10 9 10 0 9
35 13 3 3 0 10 9 13 3 3 0 10 3 12 9 1 7 0 10 9 15 13 7 10 0 9 15 10 15 9 1 12 9 0 9 13
8 13 3 3 10 9 9 9 13
21 9 3 16 13 0 13 1 10 9 9 7 13 0 7 13 1 11 10 15 1 0
14 9 3 3 7 0 1 10 0 13 0 3 1 15 0
9 13 3 1 10 15 9 13 10 9
17 7 3 13 10 9 3 15 10 0 9 13 3 3 10 3 13 9
9 13 3 3 0 12 10 1 10 9
15 0 3 3 7 0 3 3 9 10 10 9 13 13 0 15
18 0 1 10 15 9 13 10 11 10 9 16 9 13 9 7 7 9 13
4 0 13 15 9
14 11 3 13 0 13 9 1 15 13 13 13 13 1 11
10 13 3 1 11 13 1 15 11 13 0
8 6 9 0 3 3 10 9 13
8 13 3 10 9 1 10 11 9
27 13 3 0 11 13 9 10 9 9 3 0 13 9 15 10 9 9 11 0 9 13 10 10 11 10 9 13
25 0 3 10 9 0 10 9 3 3 15 13 16 10 3 0 15 13 11 13 10 15 9 13 3 13
35 10 3 9 16 15 9 10 9 10 11 13 3 13 13 13 13 16 15 3 9 13 10 3 15 9 13 0 1 1 0 10 9 13 1 11
26 3 3 0 15 10 13 10 9 1 15 10 9 13 13 13 0 7 0 7 0 3 9 7 9 7 9
24 10 3 15 9 1 0 1 9 3 13 11 3 3 10 13 7 9 13 0 1 15 15 0 13
18 11 3 13 11 13 9 1 9 7 0 7 0 3 13 7 9 7 9
19 13 3 1 11 11 0 9 0 15 9 3 7 9 13 3 9 13 10 9
24 16 3 3 15 11 13 15 3 13 15 3 7 13 9 7 3 3 13 1 10 0 10 0 9
15 3 3 10 0 9 1 10 9 13 0 10 9 13 15 13
20 0 10 1 11 9 0 7 13 9 11 7 9 13 0 9 13 15 9 13 11
6 10 3 3 15 0 13
9 13 3 0 1 10 11 9 10 9
12 13 3 3 0 0 13 3 0 1 0 10 9
37 13 3 10 10 0 15 3 3 0 13 10 9 0 13 7 1 10 9 7 13 1 10 9 3 3 1 11 10 0 1 10 0 9 3 13 10 0
7 15 3 13 1 0 0 13
37 0 3 10 11 9 13 0 0 15 15 1 10 9 0 13 0 3 9 13 3 3 15 13 0 16 3 3 1 10 15 9 10 1 10 11 13 13
6 0 3 3 1 0 13
15 1 10 3 0 9 10 9 9 15 13 0 9 0 10 9
9 0 3 3 10 9 0 15 13 13
19 10 3 9 9 13 1 10 9 13 9 10 0 9 0 13 13 13 10 9
13 10 3 9 9 13 0 13 9 0 0 9 12 0
9 16 3 0 15 15 13 1 12 13
9 10 3 0 15 3 12 9 9 13
17 1 0 3 9 13 13 7 9 7 9 7 9 7 9 7 15 15
13 15 3 3 13 0 10 0 0 13 15 13 10 13
5 9 3 15 1 9
6 9 3 15 3 13 0
14 16 3 10 11 7 0 10 9 13 13 9 1 15 13
12 10 3 11 9 13 1 15 3 13 10 0 9
20 10 3 3 9 0 10 0 3 0 9 13 10 9 1 15 10 11 13 9 13
7 6 9 9 13 13 15 13
17 13 3 7 13 10 9 0 11 10 9 13 0 10 13 9 13 0
15 10 0 3 13 0 16 13 10 13 13 3 10 9 10 11
16 16 3 13 10 11 9 13 13 9 13 1 10 9 10 9 0
24 15 3 10 0 13 3 1 9 7 13 16 16 15 0 13 13 3 3 15 13 10 9 1 9
8 11 3 9 15 0 13 13 9
23 10 7 3 0 10 0 9 3 3 13 7 3 3 0 11 13 13 10 15 12 13 12 9
13 15 3 3 1 9 7 9 7 9 9 10 15 13
8 9 3 9 15 13 0 3 15
4 0 3 13 13
15 7 10 7 0 13 9 0 7 9 0 13 1 9 10 9
21 13 3 1 10 9 7 13 15 13 13 0 10 11 9 0 10 9 15 9 13 11
7 13 3 10 0 1 9 9
16 13 3 10 0 7 10 9 13 9 10 9 0 15 9 13 11
9 10 3 11 15 3 3 9 15 13
6 0 3 0 3 13 13
16 0 3 15 10 0 1 9 0 11 13 0 9 13 10 11 13
18 10 3 11 13 0 10 11 9 1 11 13 15 0 9 0 13 11 13
16 9 3 3 9 0 7 0 13 7 10 3 15 0 9 13 0
12 0 3 13 9 13 10 1 9 9 1 0 9
7 9 3 13 10 1 9 9
11 10 3 9 15 0 1 13 10 11 13 0
19 9 3 0 13 9 13 15 10 9 9 9 0 0 13 1 0 15 3 13
6 13 3 3 0 9 13
14 7 10 3 9 10 1 13 10 9 10 3 9 10 3
3 0 3 13
26 13 3 3 15 15 9 0 13 15 10 3 9 13 0 9 3 13 0 9 7 13 7 10 3 13 0
23 1 3 11 1 12 9 0 9 0 9 9 7 9 7 9 0 0 3 3 3 1 10 0
15 10 3 9 9 9 0 9 15 13 15 15 1 9 13 13
10 10 3 9 0 15 1 10 0 9 13
7 7 1 0 15 13 13 0
6 13 3 9 7 9 0
12 9 3 0 1 9 13 1 9 13 7 0 0
59 7 3 10 9 10 0 7 10 9 1 0 13 7 10 9 7 7 9 7 9 7 7 9 10 10 9 13 7 10 0 7 10 0 10 1 10 9 10 9 13 3 3 13 3 1 9 7 10 0 9 7 9 0 7 15 9 0 9 0
9 15 3 15 0 15 1 10 9 13
9 15 3 13 3 12 9 1 10 9
3 13 3 15
11 10 3 3 9 9 9 13 0 9 3 13
8 1 9 3 1 9 13 10 0
7 0 3 10 9 13 10 11
9 10 3 9 0 13 9 15 13 13
14 1 3 3 11 10 11 0 7 7 0 9 13 1 0
22 16 3 13 10 11 13 11 10 9 1 10 11 15 9 7 15 9 10 3 13 13 9
9 1 3 10 13 15 7 13 13 0
8 10 3 3 0 9 13 0 9
6 13 3 9 15 0 13
8 13 3 15 1 11 13 15 9
9 16 3 13 10 9 0 10 11 13
6 15 3 3 0 0 13
19 10 3 9 13 13 10 9 7 10 1 9 9 13 13 9 10 3 9 13
11 10 3 0 9 13 10 9 9 16 13 13
23 10 3 9 10 13 0 1 10 11 16 13 13 13 1 9 10 11 11 9 9 7 7 9
10 15 3 16 13 13 3 0 13 10 9
7 13 3 0 13 10 9 0
28 9 3 13 0 10 1 11 13 3 3 0 13 0 7 3 13 13 7 3 3 1 10 3 9 13 16 13 9
5 9 3 0 13 13
6 11 15 15 13 0 1
3 13 3 11
39 0 3 1 10 0 9 10 11 0 7 15 3 3 3 13 7 3 3 10 11 13 9 1 3 0 1 12 9 9 13 1 10 3 9 16 15 15 0 13
9 1 11 13 9 10 0 1 10 9
13 10 3 11 15 11 3 13 9 11 3 10 9 9
11 13 3 11 9 11 13 10 9 1 10 11
11 13 3 3 0 13 10 11 7 13 10 11
37 16 3 15 3 13 13 9 10 9 0 13 15 7 0 10 11 13 0 10 0 7 13 10 9 3 9 10 9 10 0 13 13 1 10 9 3 13
9 9 3 13 0 13 9 13 1 9
37 16 3 10 9 13 10 1 10 9 10 1 11 15 11 10 9 13 0 13 9 13 10 9 7 3 15 7 13 10 9 13 7 10 0 3 13 15
7 3 3 3 15 10 0 13
3 0 3 13
14 9 3 3 0 13 10 3 13 9 13 10 3 11 0
23 9 3 15 15 13 9 13 10 1 9 9 3 3 11 10 9 9 0 0 7 0 9 0
16 15 16 13 15 9 1 10 11 13 9 13 1 7 9 7 0
6 11 3 3 9 0 13
12 3 3 1 9 10 0 13 9 1 9 9 0
14 0 3 0 9 13 1 9 0 1 15 0 11 9 13
9 6 9 0 13 15 1 0 9 13
9 10 3 11 13 9 13 1 10 11
16 9 7 3 13 0 7 9 0 1 13 7 10 9 0 7 0
15 13 3 10 11 1 10 11 13 1 10 11 13 9 3 0
9 13 3 10 9 0 13 10 0 9
6 11 15 13 9 1 9
19 10 3 3 9 10 11 9 7 10 0 3 13 15 13 10 11 9 13 15
6 13 3 15 9 1 15
20 11 3 13 1 10 9 1 0 10 13 13 0 13 10 9 13 1 10 0 9
10 11 13 3 3 0 3 13 9 13 0
9 13 3 1 11 13 16 13 10 11
19 0 10 9 10 9 13 10 0 7 1 11 9 7 0 13 3 1 9 12
11 13 11 10 0 13 15 9 1 10 9 9
9 3 13 3 13 9 13 1 10 9
11 0 3 10 0 10 0 13 13 15 9 12
5 0 3 3 13 13
32 11 7 3 9 0 13 1 11 7 10 9 1 9 11 13 7 11 9 10 0 10 11 9 7 1 10 0 13 13 9 10 11
10 0 10 9 1 11 13 0 3 3 13
8 10 3 9 13 10 0 10 9
11 3 3 3 15 13 0 7 7 0 7 9
9 15 3 15 13 9 10 9 13 13
11 13 3 10 0 3 9 13 10 9 7 9
10 9 3 3 3 1 10 9 3 12 13
11 10 3 9 13 15 7 7 0 13 15 9
14 1 9 3 15 15 13 7 10 1 0 9 13 3 13
5 7 0 3 3 13
40 9 7 3 13 10 11 10 0 7 0 13 1 9 13 13 9 1 11 13 1 10 9 9 12 9 10 0 11 9 13 13 10 1 9 9 7 15 13 15 13
6 10 3 3 15 9 13
5 9 3 15 13 11
3 13 3 11
16 13 3 0 1 10 11 7 13 1 10 9 10 11 13 10 9
4 15 3 3 13
19 13 3 0 1 12 9 7 13 10 9 3 9 15 10 9 10 9 11 13
25 11 3 13 10 13 7 9 13 16 15 13 11 10 0 10 9 13 3 3 15 9 13 1 10 9
7 13 3 1 9 11 13 13
5 3 3 3 3 13
5 10 3 3 15 13
26 9 3 15 1 10 0 9 13 7 9 1 15 10 13 15 9 0 13 0 13 1 0 13 11 15 13
13 9 3 13 15 1 9 15 13 13 15 3 9 13
20 9 7 3 13 1 10 11 7 10 9 9 13 1 10 11 13 1 10 11 3
24 3 3 13 1 10 9 10 0 10 9 13 10 9 10 0 10 3 0 0 1 10 0 9 13
12 9 3 7 9 0 13 13 9 7 7 9 13
20 13 3 10 9 10 9 1 10 11 9 3 10 9 9 13 13 10 9 10 9
23 13 3 10 9 13 1 0 7 9 13 7 9 11 15 13 1 10 0 9 1 10 11 13
12 13 3 15 0 13 13 0 7 7 10 0 9
20 11 3 3 0 13 10 13 10 1 11 13 9 13 1 10 11 13 11 10 0
9 3 3 1 0 13 13 1 10 11
12 10 3 11 13 15 13 13 13 10 9 10 9
24 15 3 13 15 16 9 11 13 9 3 13 1 10 11 13 9 3 1 10 11 7 0 1 13
13 7 3 9 3 13 9 13 13 10 11 1 10 11
11 15 3 3 1 10 11 7 10 0 11 13
12 10 3 9 10 9 13 9 0 1 10 15 13
9 7 15 7 13 7 15 15 0 13
49 13 3 0 10 13 1 10 9 10 9 10 0 3 3 1 11 10 11 0 15 0 13 9 10 11 13 10 9 13 15 13 10 9 9 10 0 3 13 13 3 3 9 0 1 10 9 13 10 9
27 7 15 10 0 10 0 13 1 0 10 9 1 9 13 3 3 9 0 13 7 13 0 10 9 1 10 9
6 0 3 3 0 13 9
6 9 3 15 11 0 13
15 11 3 13 1 9 0 15 3 13 10 9 7 9 0 13
34 13 3 0 10 11 9 11 3 13 0 10 0 13 10 0 13 16 0 13 0 3 9 1 15 13 13 13 10 3 11 13 13 0 9
12 10 3 3 1 11 13 9 13 11 11 9 9
8 1 3 10 9 13 11 0 13
18 16 13 10 9 10 9 1 10 11 10 0 9 15 3 13 9 1 0
14 16 3 13 15 10 9 3 0 13 10 9 13 10 9
12 10 3 1 0 0 10 9 0 13 13 1 9
17 0 3 10 9 13 9 1 0 1 11 13 10 9 1 10 9 13
16 3 3 13 1 11 13 10 9 16 13 15 3 15 10 9 13
8 16 3 3 15 9 9 13 13
11 13 7 10 11 7 10 9 15 13 10 9
43 0 7 13 13 7 10 9 13 15 1 9 15 13 10 9 10 12 9 1 3 0 13 9 13 0 15 1 9 13 13 1 0 10 9 3 3 7 1 15 3 13 1 11
22 3 1 9 13 15 3 0 13 13 10 0 9 0 3 3 10 9 0 3 9 13 13
12 11 3 7 10 0 13 1 11 9 9 9 13
51 1 3 3 10 1 11 10 0 9 10 3 12 9 13 1 3 10 1 0 11 0 3 0 0 3 3 16 10 3 0 13 9 0 13 1 7 10 9 7 10 9 9 0 12 9 16 3 10 0 13 12
15 10 7 3 0 9 13 9 7 7 9 11 7 3 3 9
11 3 3 13 6 9 10 9 3 13 0 0
12 3 3 15 13 15 13 3 7 0 7 0 13
9 3 3 0 13 1 11 3 13 15
6 13 3 0 13 10 9
13 10 3 0 13 9 1 11 13 1 10 9 10 0
14 0 3 13 10 9 13 1 10 0 10 9 13 3 0
17 16 3 13 9 12 9 3 13 15 7 9 13 7 13 0 10 9
11 11 13 1 11 7 13 9 12 9 3 13
12 7 3 3 13 1 10 9 10 9 9 13 13
11 13 3 3 15 1 9 9 13 11 10 11
21 0 0 3 9 11 3 9 13 1 15 3 10 9 10 1 11 13 9 13 9 13
11 15 3 13 10 9 13 13 3 15 15 13
4 13 3 3 9
9 15 15 3 13 10 9 13 10 0
5 13 3 1 0 11
16 7 3 1 10 9 0 13 7 15 9 13 11 10 9 7 11
22 15 3 13 7 15 13 7 9 13 13 1 11 10 9 13 16 1 11 13 10 9 13
7 1 11 3 13 13 9 11
11 16 3 15 13 9 13 1 10 9 10 9
9 1 3 0 13 10 9 13 1 11
11 7 3 15 1 0 13 10 9 10 0 13
12 1 12 3 3 10 0 3 0 13 10 11 13
6 13 3 13 15 10 9
10 3 15 0 13 3 1 15 10 11 13
12 1 7 0 3 0 13 16 0 13 13 9 13
7 6 0 13 3 15 13 0
16 13 3 15 10 9 16 9 10 9 13 10 11 13 0 10 9
11 3 0 7 13 1 9 15 3 3 13 13
6 0 3 3 13 1 9
27 1 0 3 3 9 15 13 15 13 3 0 3 13 13 7 13 13 0 1 10 9 3 15 0 13 10 9
11 0 3 3 13 13 13 12 9 13 0 13
13 13 3 13 13 11 7 11 13 15 1 9 10 9
12 0 3 13 3 13 10 0 13 9 13 15 0
6 13 3 11 0 3 13
18 10 3 0 11 7 10 11 7 11 10 11 9 10 9 0 13 10 9
22 3 3 10 0 9 10 0 9 13 13 11 13 7 10 9 13 0 13 1 10 15 0
12 13 3 3 0 9 3 0 13 13 1 10 9
6 15 3 13 3 13 0
17 0 3 13 1 10 11 10 9 13 0 13 7 1 9 10 0 13
19 7 3 3 13 15 0 10 0 10 9 7 9 1 15 10 0 0 3 13
8 0 3 13 0 13 1 10 9
25 10 3 0 9 13 3 10 9 15 3 3 13 13 0 3 13 9 10 9 13 15 3 7 11 13
11 3 3 13 10 0 1 10 11 13 0 15
9 10 3 9 0 13 0 7 7 9
12 0 3 13 10 9 13 9 13 3 1 10 9
8 7 15 3 13 10 9 3 13
3 13 3 9
10 0 3 13 10 9 13 3 13 10 9
12 0 3 1 10 15 9 13 12 15 15 9 13
10 15 3 13 10 13 3 13 3 13 0
33 1 3 11 11 10 0 9 9 11 11 3 10 10 9 13 0 7 13 0 3 9 15 15 13 10 0 9 0 10 1 11 9 13
18 16 3 1 9 13 10 9 9 13 1 7 9 7 10 13 1 10 0
8 6 9 11 13 3 3 10 9
23 0 7 3 13 11 7 11 1 3 11 11 7 0 7 11 0 1 10 11 11 13 10 9
18 0 13 1 9 11 13 16 1 0 13 11 13 15 3 15 13 0 13
7 0 3 3 0 10 11 13
15 13 3 3 10 15 9 7 7 10 9 1 9 1 10 11
13 7 3 3 13 7 10 9 10 9 13 7 0 13
27 13 3 11 1 11 7 11 10 9 15 9 13 0 1 10 9 16 13 15 13 9 1 10 9 9 3 13
10 7 15 13 7 10 13 0 7 0 13
14 0 13 3 0 9 9 13 7 13 0 10 11 9 13
14 0 7 3 13 13 7 10 7 9 7 10 9 9 13
27 13 3 13 3 3 9 7 15 13 9 7 15 3 13 3 0 7 0 0 7 3 3 9 7 7 9 13
26 13 3 3 13 7 15 9 9 15 7 9 15 9 13 15 15 0 7 13 13 1 9 0 15 13 13
38 7 3 0 3 13 9 16 9 3 7 9 7 9 7 7 0 0 7 9 0 7 0 13 9 15 7 9 13 13 13 9 13 9 3 13 9 3 13
17 15 13 13 0 9 7 13 7 9 13 10 9 7 15 3 3 9
21 7 3 3 11 10 11 9 16 13 10 0 9 10 9 7 13 13 3 10 9 9
11 13 10 13 9 16 13 10 9 7 13 13
7 9 3 13 13 0 9 13
19 7 16 3 3 15 13 13 9 10 9 13 10 15 9 1 3 15 3 15
7 10 3 0 15 10 9 13
11 15 3 9 13 15 3 0 13 13 15 0
18 11 3 0 13 10 9 3 7 13 1 10 9 7 13 9 1 11 13
5 11 3 0 15 13
15 7 7 1 10 3 7 1 10 3 3 13 13 10 0 13
27 13 3 11 13 1 0 0 9 1 10 9 13 15 10 9 13 13 13 7 1 15 9 13 7 15 15 9
5 15 3 1 0 13
16 9 3 0 7 9 3 0 1 9 10 0 1 9 10 0 11
15 10 3 9 9 1 7 10 0 9 13 7 3 3 1 0
20 13 3 10 9 13 13 16 0 13 15 15 13 9 7 7 9 1 10 11 3
3 15 3 13
6 11 3 13 10 13 13
36 3 1 0 9 0 3 0 1 11 10 11 9 0 11 9 9 13 11 9 13 1 9 13 15 3 1 10 11 10 9 1 11 13 9 0 13
17 10 7 3 9 13 0 13 7 10 13 10 9 10 11 13 10 9
34 13 3 0 9 13 9 3 13 7 10 9 9 13 13 3 7 10 9 9 13 3 7 3 16 3 13 10 9 10 9 13 7 10 9
12 10 3 12 13 1 15 7 13 15 13 13 3
20 13 3 0 3 10 0 7 7 10 9 1 3 0 0 9 0 9 3 3 13
6 13 3 3 1 11 11
15 1 3 10 9 13 3 12 9 7 3 10 0 9 13 3
11 7 13 3 1 9 3 15 3 9 9 0
25 16 15 10 9 10 9 3 0 3 13 13 3 10 0 9 3 13 15 13 1 10 11 7 13 3
4 15 3 13 13
16 7 3 3 3 15 13 13 10 9 0 1 0 9 13 9 13
3 13 3 3
8 1 9 3 7 3 9 13 9
18 1 9 3 13 3 10 0 9 16 3 13 10 3 1 9 15 9 13
9 3 3 13 13 10 9 15 9 13
12 3 3 10 7 9 10 0 7 10 9 10 0
49 3 3 13 10 9 10 0 13 7 0 9 3 13 3 10 9 10 9 7 13 0 10 9 13 1 15 3 10 9 0 10 9 13 13 1 9 11 7 9 0 7 0 9 13 16 15 13 1 11
13 15 3 3 0 13 9 1 9 3 13 13 10 0
29 1 3 10 9 13 9 13 9 0 1 3 10 9 9 0 0 9 0 9 0 1 3 10 9 9 1 3 9 9
9 0 3 0 10 9 13 7 3 0
18 0 3 1 3 10 9 3 10 0 13 13 9 3 0 0 7 9 0
6 13 3 13 11 10 11
7 9 3 9 3 13 13 13
7 9 3 0 13 1 0 0
8 10 3 0 0 1 9 9 13
12 9 3 1 3 10 9 13 9 0 9 3 0
4 13 3 3 9
16 9 3 1 3 10 9 9 0 0 13 9 3 0 0 7 9
7 9 3 7 9 13 15 9
12 9 3 15 1 10 0 9 9 7 7 9 13
5 0 0 13 1 9
11 0 3 13 3 3 1 10 0 7 0 3
4 13 3 15 0
4 0 3 3 13
6 0 3 10 0 0 13
5 9 3 12 13 9
6 0 3 9 7 9 0
16 9 3 7 9 7 9 7 0 9 0 13 1 10 9 13 12
13 3 3 13 0 7 13 1 9 1 9 12 0 13
27 3 3 3 15 13 3 16 15 9 7 10 0 10 1 9 13 9 13 3 0 13 15 13 13 3 13 0
30 16 3 0 0 12 9 10 9 10 15 0 13 15 3 3 13 12 13 0 7 3 3 13 3 10 9 10 1 15 13
13 13 3 9 10 15 9 15 13 9 9 12 3 13
17 3 3 3 0 1 3 12 13 0 13 0 9 0 3 0 9 0
15 11 3 1 9 7 13 7 3 13 9 15 7 3 15 13
20 1 3 0 10 9 0 10 1 10 9 7 10 9 13 1 10 9 1 10 11
9 13 3 10 0 10 9 3 0 9
20 9 3 15 3 9 0 13 15 15 13 7 13 10 1 15 3 13 0 0 9
20 12 3 9 13 10 9 0 13 0 1 15 9 7 7 9 9 10 0 13 13
13 13 3 3 1 9 10 1 10 0 13 1 10 11
8 7 3 15 13 1 10 0 13
22 13 3 0 9 13 1 10 11 16 11 13 9 1 11 0 3 3 13 13 1 10 11
12 9 3 11 3 13 13 7 15 13 9 11 0
12 1 11 9 10 1 11 13 13 9 9 9 13
12 15 3 13 9 0 1 11 15 13 9 1 11
11 0 3 9 0 10 9 10 0 10 0 13
28 16 3 15 3 15 13 15 3 3 13 13 10 3 13 10 11 13 0 0 3 3 0 13 16 13 15 10 11
12 16 3 15 9 10 1 9 13 10 0 15 13
9 15 3 13 0 3 3 0 13 0
17 13 3 10 11 10 15 9 13 3 16 10 9 1 10 9 13 13
16 3 3 3 0 3 13 13 10 11 10 9 13 1 11 10 9
19 13 3 11 9 7 0 3 9 13 7 0 3 0 7 0 0 3 15 13
39 3 3 13 13 10 9 7 1 11 7 11 9 10 0 13 10 9 13 3 0 10 9 3 13 13 3 10 9 13 13 3 10 9 13 0 13 15 10 11
15 13 0 0 1 11 10 9 13 16 15 0 13 13 10 11
5 1 3 13 9 9
16 10 3 9 1 0 13 1 11 13 1 9 0 9 13 10 9
21 0 13 10 1 11 9 9 7 13 13 1 10 11 1 10 11 7 13 3 1 11
13 10 3 3 1 11 9 1 10 11 13 3 0 9
7 1 0 3 13 13 10 9
29 10 3 0 11 9 13 1 11 9 13 9 10 0 13 12 3 11 3 13 13 9 12 0 0 7 7 0 7 0
8 10 3 3 12 10 9 3 13
19 13 3 1 0 10 9 1 0 10 0 9 9 7 7 9 7 9 12 9
24 0 3 10 1 0 10 11 9 13 13 1 7 10 9 10 13 7 10 0 9 7 15 13 0
5 0 3 10 9 3
22 10 3 3 0 15 13 13 10 9 0 3 3 0 13 7 9 13 11 13 1 9 11
27 10 3 9 10 0 1 10 9 10 0 13 0 9 1 15 10 9 10 0 13 13 15 10 13 1 10 9
7 10 11 1 9 0 9 13
18 10 3 1 11 9 13 3 15 0 15 13 11 3 0 13 3 3 3
16 1 3 10 9 0 13 9 0 3 3 0 3 3 3 3 0
4 9 3 0 13
14 0 3 1 11 13 1 3 9 9 7 12 7 0 12
10 13 3 1 10 0 11 0 10 9 13
12 15 3 10 3 13 15 1 10 9 10 9 13
14 13 3 15 13 11 0 0 13 13 10 13 1 10 0
15 3 3 1 9 7 7 0 9 10 1 9 13 7 9 0
6 13 3 10 9 1 9
18 1 0 10 9 10 9 13 9 13 3 13 1 10 9 13 1 10 9
17 10 3 11 0 13 3 11 1 0 9 15 15 1 10 3 9 13
9 10 3 9 0 13 3 10 0 9
9 13 3 3 13 10 9 3 1 9
8 15 3 3 3 13 10 9 13
9 3 3 15 9 13 9 7 9 3
8 13 3 15 11 1 9 9 13
10 0 3 3 13 15 1 10 9 7 13
14 10 3 11 11 3 10 9 13 9 11 3 10 11 9
12 0 3 7 0 0 9 13 11 10 0 13 9
13 10 3 10 9 11 11 10 11 13 1 9 10 13
8 10 3 3 1 11 9 3 13
2 0 3
8 1 0 10 9 13 13 10 0
8 10 7 13 13 7 10 0 13
5 9 3 13 1 15
27 13 0 16 9 13 1 10 11 0 7 3 3 1 10 9 10 1 11 13 3 3 15 13 15 0 0 13
40 16 3 3 13 1 10 11 3 13 13 10 0 16 3 3 15 3 15 13 11 3 9 11 3 9 11 13 13 0 10 9 13 13 3 13 15 9 1 10 9
