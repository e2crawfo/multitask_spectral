3557 11
6 9 9 1 11 1 9
10 11 3 13 9 9 1 9 0 9 2
9 3 1 9 2 13 16 0 9 2
19 11 13 9 2 13 15 9 15 9 2 7 9 1 9 13 9 0 9 2
27 16 1 11 2 9 13 16 4 0 9 15 15 13 1 9 0 7 3 0 2 15 13 0 9 1 9 2
19 13 16 15 9 7 9 13 13 0 9 1 9 16 0 14 13 3 15 2
32 7 13 14 0 9 2 1 9 16 9 1 0 9 13 13 16 9 2 7 3 7 3 2 13 1 9 16 13 9 1 9 2
7 11 11 4 12 15 9 2
32 2 15 4 9 13 1 9 11 2 2 16 14 15 2 1 9 12 9 2 16 3 4 13 9 3 15 4 15 0 9 13 2
19 13 4 15 16 4 1 9 13 3 15 9 2 7 15 15 4 13 2 2
41 1 15 4 11 0 12 9 2 2 4 13 15 9 2 7 3 4 15 15 9 3 14 13 2 1 9 16 4 0 9 13 15 9 2 2 13 4 11 1 11 2
19 1 15 9 2 9 4 0 3 1 9 16 1 9 16 15 13 1 9 2
20 15 4 0 2 0 9 15 4 13 0 9 13 4 9 11 16 13 15 9 2
39 1 15 2 0 9 15 4 0 13 4 9 9 2 7 3 3 15 0 2 16 15 4 11 2 13 1 0 9 2 15 13 1 0 9 1 9 1 9 2
14 11 11 2 0 9 1 9 11 2 0 4 9 15 2
11 2 9 3 2 13 16 4 9 3 0 2
30 9 0 9 3 14 13 7 15 13 1 9 9 2 9 16 9 2 13 15 2 4 4 3 9 2 7 9 15 13 2
25 1 9 4 14 9 0 9 4 3 0 2 16 14 9 15 4 13 2 2 13 4 11 1 11 2
28 3 1 12 9 9 0 1 9 1 9 2 7 15 0 9 14 13 2 13 4 9 0 7 0 9 0 9 2
24 11 13 16 4 15 3 2 7 16 4 15 9 1 9 13 3 12 7 3 9 1 15 9 2
15 11 11 2 0 9 9 1 0 9 2 13 15 1 15 2
35 2 0 9 4 9 1 0 9 2 1 9 16 15 9 2 9 2 13 1 0 9 2 9 9 7 9 1 9 2 2 13 4 1 11 2
22 3 4 7 9 0 9 2 2 1 15 9 2 9 4 13 13 0 9 7 9 2 2
34 11 13 3 4 2 1 15 9 2 9 2 4 0 2 2 2 1 9 1 0 9 2 2 7 16 4 9 13 1 0 9 1 9 2
24 13 1 9 1 0 9 11 11 2 3 4 3 4 2 3 12 9 1 9 15 4 3 0 2
23 3 15 9 13 2 3 1 2 12 15 2 7 12 9 0 9 4 0 2 2 13 11 2
11 11 13 3 4 0 9 13 1 0 9 2
9 2 3 4 0 9 9 0 9 2
10 9 4 13 13 9 15 13 0 9 2
5 3 4 9 0 2
20 3 4 1 9 15 15 7 3 13 2 2 14 13 2 9 1 9 1 9 2
26 11 4 0 9 1 15 9 0 9 16 15 13 9 9 1 9 13 9 9 2 2 13 4 1 11 2
29 0 9 0 4 3 9 9 11 1 0 11 2 15 4 13 9 9 11 11 16 13 1 9 0 7 0 9 9 2
6 8 4 0 12 9 2
7 9 0 9 13 9 1 11
24 15 13 16 4 9 11 11 9 1 9 9 2 16 0 13 3 9 1 15 0 9 13 3 2
30 0 9 7 0 9 0 9 11 11 2 15 4 3 13 0 9 2 13 4 13 9 2 13 9 1 15 0 0 9 2
54 11 2 0 9 0 9 8 2 12 9 7 0 9 2 0 4 1 0 9 1 11 12 9 1 12 9 9 1 9 9 2 0 9 2 9 9 7 9 9 2 12 9 13 4 0 9 1 9 1 12 1 12 9 2
18 9 8 7 12 9 0 4 3 15 4 13 9 7 13 9 1 9 2
43 2 9 4 16 4 9 0 1 15 9 2 15 4 0 9 2 0 7 16 9 14 13 0 9 1 9 9 1 0 9 2 2 13 4 1 11 9 0 9 11 11 11 2
43 0 9 2 7 3 0 9 8 11 2 13 16 15 9 2 1 9 2 0 9 2 2 13 9 1 9 7 3 0 0 9 1 11 2 15 4 13 15 9 7 13 9 2
20 2 0 0 9 13 4 1 0 9 15 0 9 7 15 9 15 4 1 15 2
45 15 9 2 7 3 15 15 7 13 2 4 4 13 8 11 7 11 11 2 16 9 9 1 9 2 9 2 11 11 2 2 13 4 0 9 8 11 7 9 0 0 9 11 11 2
25 9 4 13 16 4 8 11 0 3 16 4 15 9 9 2 7 16 4 11 0 1 0 0 9 2
45 2 15 4 0 9 1 9 7 9 15 13 1 0 9 2 7 15 9 13 3 1 0 9 0 9 7 9 9 16 3 13 15 9 2 2 13 4 9 0 11 11 11 1 11 2
37 9 4 13 12 9 15 4 13 16 4 11 13 13 12 9 9 9 2 7 16 4 13 12 9 9 1 9 2 16 15 4 9 9 1 0 9 2
27 11 4 13 1 15 12 9 2 15 13 7 1 11 7 0 0 9 2 15 4 9 13 1 9 8 11 2
23 1 9 9 0 9 8 8 11 11 2 3 13 15 15 4 9 13 7 13 9 8 11 2
16 11 4 13 16 4 8 13 9 0 9 11 1 9 9 9 2
21 2 0 4 16 4 2 0 9 2 13 15 9 1 0 9 2 2 13 4 11 2
24 15 0 2 16 15 4 0 9 11 11 2 13 16 14 13 9 15 13 9 0 1 9 9 2
10 2 13 14 16 15 9 13 7 14 2
26 9 9 1 11 0 4 7 0 2 7 9 1 8 11 15 4 13 1 9 3 3 13 1 15 9 2
22 15 2 2 2 4 13 0 9 1 9 7 13 0 9 2 0 4 0 1 0 9 2
16 1 15 4 9 0 9 9 2 2 2 13 4 11 1 11 2
9 9 9 11 11 13 9 1 15 9
18 9 9 11 11 11 13 4 9 0 0 9 2 3 0 9 1 9 2
35 9 9 11 7 11 2 11 2 11 11 13 4 1 9 2 12 9 2 9 1 9 9 0 9 2 11 2 7 0 9 1 0 9 9 2
18 11 2 0 9 0 9 2 12 4 1 0 9 1 9 11 7 11 2
40 2 13 9 9 2 11 2 7 13 1 15 9 13 1 0 9 1 0 9 1 9 2 2 13 4 11 9 1 15 4 13 16 13 9 1 0 9 1 9 2
39 16 1 11 4 4 9 2 0 13 16 0 0 9 13 1 15 9 1 9 9 11 11 2 15 4 13 9 0 9 0 9 11 11 1 0 0 9 11 2
26 9 9 11 11 0 9 4 4 9 9 2 16 4 11 13 9 11 2 9 7 9 9 15 9 11 2
14 2 4 4 3 16 13 1 9 7 16 13 12 9 2
9 15 13 2 2 2 13 9 11 2
24 1 0 4 4 0 9 1 0 9 2 2 13 4 11 9 1 11 1 9 1 11 12 9 2
17 11 4 13 0 9 1 0 9 1 11 1 0 0 9 12 9 2
13 0 4 15 4 3 9 15 9 9 9 1 9 2
45 0 9 9 13 4 16 4 0 9 1 9 1 9 1 9 0 9 2 11 2 4 0 2 7 0 9 13 15 4 7 9 0 9 2 16 7 9 15 4 13 9 11 1 9 2
15 2 11 7 11 13 4 11 3 15 1 9 0 0 9 2
22 15 9 3 4 9 9 9 2 2 13 4 1 11 9 1 0 9 1 11 11 11 2
6 9 1 11 13 3 2
7 0 0 9 13 4 9 2
6 2 9 13 9 9 2
26 15 4 15 0 9 7 15 9 1 9 4 9 15 2 2 13 4 1 11 11 11 2 0 9 11 2
18 11 11 2 9 11 2 13 16 4 0 9 13 13 1 0 9 9 2
36 2 15 4 13 13 9 9 11 7 9 0 9 1 9 16 4 11 2 3 1 0 9 9 2 0 1 0 9 2 2 13 4 11 1 11 2
25 3 3 9 1 0 0 9 2 9 4 13 9 7 13 11 1 0 9 2 1 9 1 0 9 2
17 2 15 3 4 13 12 9 2 7 15 13 1 9 2 1 11 2
20 15 4 4 15 9 16 13 1 15 2 2 13 4 1 11 11 11 1 11 2
10 2 9 4 0 9 16 15 4 11 2
13 16 4 9 13 15 9 2 0 4 16 15 13 2
17 1 15 15 3 3 13 2 2 13 4 9 11 11 11 1 11 2
10 0 9 11 13 4 15 1 9 7 9
13 1 3 12 9 1 9 2 11 3 13 0 9 2
20 0 9 11 2 0 0 9 11 11 2 13 4 16 4 13 9 9 9 11 2
12 3 2 3 4 15 13 2 13 13 3 9 2
9 11 13 9 1 0 9 0 9 2
9 9 4 4 1 9 3 12 9 2
9 2 12 1 0 0 9 4 0 2
32 0 9 9 9 0 4 1 9 7 9 2 2 13 4 11 9 1 9 2 12 9 2 3 4 9 13 9 9 1 12 9 2
9 15 0 9 4 4 9 0 9 2
25 1 0 9 0 4 16 15 9 13 13 2 7 13 16 0 9 13 9 2 7 14 3 0 9 2
16 2 13 13 16 0 9 2 15 4 13 12 9 2 4 0 2
27 3 15 13 1 0 9 15 13 14 3 1 0 9 2 7 7 1 0 0 9 2 2 13 4 11 9 2
21 9 1 9 7 9 11 11 13 4 16 4 0 9 11 13 4 0 9 7 9 2
13 2 13 16 4 15 9 13 1 9 1 0 9 2
29 3 2 15 4 0 7 0 9 2 7 0 9 13 13 16 9 13 1 9 0 9 2 2 13 4 11 1 11 2
19 9 4 12 9 13 13 9 2 7 4 13 13 9 15 4 13 9 9 2
32 9 13 1 9 16 9 1 0 9 2 15 13 9 9 1 9 2 13 12 9 2 16 4 9 0 9 13 13 1 9 9 2
18 1 9 12 9 2 3 4 9 13 15 9 7 13 0 9 1 9 2
12 1 9 12 9 2 15 4 15 13 0 9 2
11 0 9 4 13 16 4 9 11 4 9 2
17 2 0 15 4 9 16 3 13 9 2 16 15 13 3 16 9 2
9 7 13 16 4 15 9 0 9 2
31 9 4 13 13 16 4 11 9 9 7 9 2 7 13 4 9 15 2 7 13 13 0 9 2 2 13 4 11 1 9 2
16 12 1 15 9 4 2 13 4 9 9 11 11 2 9 9 2
16 2 1 9 4 0 9 1 11 7 9 0 9 3 4 0 2
24 13 4 15 13 0 15 9 7 9 1 9 1 9 1 0 9 2 2 13 4 11 1 11 2
4 11 15 13 2
10 2 0 0 9 0 4 1 9 9 2
29 1 15 13 9 2 0 9 2 9 9 2 9 1 9 1 9 7 9 0 9 1 9 7 9 2 2 13 4 2
29 16 15 9 13 1 15 9 1 15 13 14 0 9 13 9 15 9 2 0 15 13 16 4 3 3 14 13 9 2
8 2 11 3 3 4 13 9 2
7 15 4 16 9 1 9 2
26 9 15 14 13 13 1 9 2 15 14 13 1 9 2 2 13 4 1 11 11 11 2 9 1 11 2
26 2 13 0 9 2 13 13 2 9 2 15 9 2 16 4 13 9 2 2 16 3 14 13 9 9 2
7 13 14 9 13 15 9 2
23 13 16 4 2 7 9 13 0 0 9 9 2 2 13 4 0 11 11 1 9 1 11 2
15 2 4 4 1 9 1 9 9 2 13 0 9 1 9 2
12 0 9 7 9 13 4 7 13 2 9 2 2
8 15 15 13 16 4 15 0 2
31 1 3 4 0 2 13 4 3 12 0 9 2 15 4 0 0 9 1 15 9 2 2 13 4 1 11 0 9 11 11 2
9 11 11 2 11 4 13 9 1 11
30 9 1 11 1 11 2 11 7 11 3 4 13 0 9 0 11 2 13 0 9 11 11 1 0 9 1 8 8 8 2
5 0 9 11 11 2
18 8 8 8 2 9 9 2 13 14 9 9 1 9 1 9 9 11 2
11 11 11 2 9 9 11 3 13 0 9 2
33 9 16 15 16 11 16 0 9 11 2 16 7 9 9 3 9 14 13 1 15 9 13 15 9 1 15 4 15 13 1 0 9 2
18 13 16 4 0 9 9 9 9 1 9 11 2 3 13 0 0 9 2
45 16 14 4 0 0 9 0 9 7 0 0 9 1 15 9 2 13 4 4 9 0 2 0 9 2 11 2 15 4 13 3 13 9 3 0 11 2 16 13 0 0 9 1 9 2
15 11 2 16 4 9 13 13 1 11 7 15 9 1 11 2
8 13 14 0 7 15 0 9 2
14 11 2 9 11 3 4 13 15 0 9 1 9 11 2
28 3 3 13 9 16 4 15 2 16 9 9 1 9 1 11 7 11 2 13 0 9 15 9 3 1 15 9 2
28 3 2 3 4 16 4 0 9 7 9 1 15 4 4 0 3 13 1 9 0 1 9 15 0 7 0 9 2
16 16 0 9 2 0 4 13 3 0 9 1 11 7 1 11 2
17 13 14 1 15 13 14 13 3 1 15 2 3 7 1 15 9 2
24 11 2 13 14 16 4 11 13 9 1 11 1 11 7 16 4 15 13 1 0 9 1 9 2
10 3 2 13 14 9 0 9 1 9 2
13 0 9 13 9 1 9 1 9 9 9 1 11 2
15 9 4 13 15 9 1 9 9 1 9 3 9 3 9 2
15 11 2 9 11 13 4 0 9 0 1 9 9 1 11 2
29 13 9 16 4 15 9 1 9 2 16 7 9 0 12 9 9 0 9 2 11 7 11 2 3 13 0 9 9 2
14 0 9 15 13 9 9 11 7 9 15 1 15 13 2
28 15 0 9 9 1 0 7 0 9 2 7 9 1 11 13 15 9 2 0 4 9 9 0 9 7 0 9 2
17 11 2 13 14 9 1 9 1 11 7 11 9 9 11 1 11 2
37 11 2 9 1 9 1 11 7 11 0 4 9 7 7 1 15 9 14 13 1 9 1 9 2 7 1 9 14 4 13 13 9 15 9 1 11 2
13 3 2 11 16 0 9 9 13 16 4 13 9 2
15 15 13 13 15 0 9 1 9 9 2 7 3 0 9 2
12 11 2 15 4 15 13 16 3 4 0 9 2
25 15 7 9 13 0 9 2 16 15 9 13 1 9 9 7 9 1 11 2 11 13 13 15 9 2
12 11 2 3 2 13 15 16 1 15 4 13 2
13 9 11 0 4 7 0 1 9 16 13 9 11 2
13 0 4 9 3 13 1 9 15 9 7 13 9 2
24 9 9 9 1 15 0 7 0 9 7 4 0 2 7 4 1 9 0 9 1 15 9 13 2
12 11 2 13 4 0 9 15 13 9 1 11 2
15 16 4 15 13 7 3 11 13 15 9 15 9 9 9 2
19 11 2 0 9 13 1 0 9 1 11 2 11 2 11 7 11 7 11 2
22 1 15 15 9 3 13 16 0 2 0 9 11 7 13 15 9 9 9 9 3 9 2
32 0 9 13 3 3 16 15 13 1 15 9 2 16 15 4 3 0 3 4 1 15 9 9 7 0 4 15 13 1 15 9 2
22 0 9 11 11 8 11 11 2 3 2 7 11 13 1 9 1 0 9 1 9 11 2
9 11 2 4 14 0 9 1 9 2
22 11 2 3 4 9 1 0 9 1 9 11 2 1 9 13 0 9 7 13 0 9 2
23 3 2 9 4 3 7 3 13 1 0 9 2 16 1 15 1 15 9 14 4 13 13 2
15 11 2 3 4 11 13 1 15 9 1 0 9 1 11 2
6 4 14 0 9 9 2
34 11 2 15 4 9 9 0 0 9 9 12 3 4 13 9 1 9 9 1 9 2 16 7 1 0 7 0 9 9 1 9 0 9 2
9 3 0 2 9 4 1 0 9 2
17 3 15 4 3 15 15 2 1 15 0 9 2 4 13 0 9 2
12 0 4 3 4 15 9 13 1 0 3 9 2
15 11 2 13 14 16 11 1 9 9 13 9 1 9 9 2
28 11 2 9 11 13 7 0 9 7 0 9 2 7 3 4 0 15 0 9 16 13 9 9 9 1 9 12 2
22 11 2 3 4 9 11 13 1 9 9 0 9 9 7 0 9 1 9 2 8 2 2
6 13 14 9 15 9 2
10 11 2 9 15 13 3 4 15 13 2
15 1 0 2 16 15 13 0 9 2 13 15 9 0 9 2
25 13 15 3 4 9 15 4 13 0 9 2 3 9 11 7 9 8 11 11 2 15 1 9 0 2
9 11 2 3 13 1 9 1 9 2
22 15 4 15 9 1 9 9 1 11 7 1 15 4 9 15 2 1 15 9 2 0 2
9 11 2 0 4 9 1 0 9 2
17 0 4 9 3 4 1 15 9 9 3 3 0 7 1 12 9 2
8 1 9 15 13 0 0 9 2
12 0 9 15 13 9 13 9 2 7 14 9 2
11 0 4 0 0 0 9 7 0 0 9 2
5 15 13 4 0 2
3 11 13 9
18 0 9 13 4 1 9 0 9 0 9 2 1 9 9 9 9 11 2
25 9 11 11 11 13 4 1 9 2 12 9 2 0 9 0 9 2 1 9 9 0 9 9 11 2
35 9 1 12 9 13 4 9 0 9 9 7 9 2 8 2 2 7 13 4 15 0 0 0 9 2 11 2 7 9 0 9 2 11 2 2
14 9 15 9 9 11 13 15 3 0 9 1 12 9 2
19 0 9 13 4 0 9 1 9 1 12 9 2 7 15 13 13 12 9 2
60 9 9 2 0 1 9 9 11 1 9 1 11 2 13 15 0 0 0 9 2 8 2 7 9 9 9 9 0 9 1 0 9 1 9 2 8 2 2 13 15 9 9 2 13 0 9 2 9 9 13 1 0 9 0 9 7 13 9 9 2
7 0 4 3 12 9 9 2
15 9 12 9 0 4 9 2 9 7 9 13 0 9 2 2
11 2 9 0 9 2 0 4 1 9 12 2
28 1 9 12 0 4 9 1 15 15 13 0 9 2 16 7 9 2 1 9 9 0 9 1 9 0 9 2 2
28 9 2 1 7 15 13 1 9 1 0 9 0 1 9 9 2 9 9 7 0 9 2 0 4 1 9 12 2
8 15 9 13 15 1 9 9 2
46 9 2 0 9 15 14 13 13 3 16 9 4 0 1 9 7 9 0 0 9 7 1 0 9 2 2 0 4 1 9 12 2 7 0 4 9 2 15 14 13 4 0 0 9 2 2
10 9 12 9 15 13 9 9 0 9 2
23 0 4 9 12 2 15 4 0 9 0 9 0 9 0 1 0 9 2 1 9 0 9 2
16 1 9 12 0 4 9 9 9 0 9 1 9 15 9 11 2
15 0 4 9 12 2 1 15 4 0 9 7 9 9 11 2
24 9 9 9 2 0 1 9 12 2 0 4 7 0 4 9 15 15 13 1 0 9 0 9 2
14 1 9 2 1 9 0 9 0 4 0 9 1 9 2
19 1 3 12 9 15 4 13 9 1 9 9 2 12 4 13 1 15 9 2
35 16 9 9 13 0 9 9 15 4 11 13 1 9 1 9 9 11 2 3 3 12 9 9 13 4 0 3 4 15 9 13 1 9 11 2
22 1 9 9 9 8 8 2 0 9 9 4 1 9 1 9 11 7 3 0 0 9 2
8 11 0 1 9 9 15 13 11
33 11 1 0 12 9 13 13 9 9 15 13 11 2 7 13 13 1 9 9 9 12 2 13 4 9 11 1 9 11 11 1 9 2
30 2 13 4 3 3 9 2 3 2 1 9 9 7 0 9 7 9 1 9 2 2 13 4 9 11 1 9 11 11 2
40 0 12 9 4 4 0 1 0 9 16 13 12 9 11 12 9 2 13 4 0 9 0 9 2 11 2 1 9 2 12 9 2 2 3 11 1 9 0 9 2
47 2 11 13 0 9 1 9 2 7 7 3 9 1 15 2 3 2 1 9 9 7 0 9 7 9 1 9 2 2 13 4 9 11 1 9 11 11 1 9 1 0 9 0 9 11 11 2
19 2 0 4 15 13 1 9 16 4 1 0 0 9 4 3 3 13 2 2
25 11 4 13 16 13 13 9 1 11 1 9 12 2 15 4 15 13 9 9 15 9 1 9 12 2
24 9 4 13 1 9 12 2 1 3 4 0 12 1 12 0 9 2 1 15 4 12 3 0 2
29 11 11 2 9 11 1 11 2 13 4 16 4 15 12 1 12 9 1 15 15 3 13 13 13 1 9 15 9 2
32 1 15 2 15 4 9 13 4 0 12 0 9 7 3 3 15 1 16 15 11 13 0 9 1 9 9 0 9 11 12 9 2
35 2 0 1 0 2 9 1 11 3 13 2 2 13 4 11 2 3 9 3 4 11 13 0 9 1 9 9 1 15 1 0 9 1 9 2
17 9 4 3 13 11 1 9 1 9 11 2 15 4 13 0 9 2
32 1 15 2 11 4 13 16 2 3 16 4 9 1 11 7 11 1 0 9 0 2 13 9 1 9 9 1 9 7 0 9 2
27 11 4 9 1 11 13 3 4 15 9 13 0 9 1 9 0 9 7 4 0 13 0 9 11 1 9 2
15 2 0 4 1 15 7 15 4 7 13 2 2 13 4 2
25 3 2 1 9 1 9 2 11 4 13 3 15 4 4 0 9 7 16 4 4 3 3 0 9 2
40 1 0 9 1 0 9 11 11 2 9 11 11 11 11 13 4 3 4 9 15 9 13 0 9 1 0 9 9 1 12 2 1 9 16 11 13 9 0 9 2
38 11 4 13 16 4 2 1 9 1 11 2 2 3 13 9 11 16 13 0 15 4 1 15 9 3 4 13 9 1 0 9 7 13 9 11 12 2 2
11 9 11 13 11 1 9 9 1 9 1 9
25 1 9 15 13 1 11 1 0 9 11 1 11 2 9 13 9 1 9 9 9 1 9 1 11 2
29 0 9 11 11 11 2 3 2 13 1 0 9 11 11 2 1 9 2 7 9 11 11 1 0 9 11 1 11 2
24 1 9 11 1 9 9 1 9 1 11 0 9 2 9 4 13 3 4 13 13 1 9 9 2
34 1 9 2 12 9 2 2 9 4 13 3 4 15 9 13 9 1 9 9 0 9 1 9 1 11 2 15 4 11 13 9 1 11 2
19 16 4 9 9 13 3 4 11 13 9 1 9 2 9 1 9 13 9 2
13 11 4 13 16 4 15 9 13 15 9 4 0 2
26 9 11 11 13 4 1 9 1 0 9 11 11 8 11 11 2 15 4 13 16 4 9 13 9 11 2
22 15 4 2 3 2 13 16 4 2 15 9 4 0 2 11 3 13 9 9 15 9 2
25 11 4 13 16 4 0 13 9 1 9 1 15 9 2 7 3 15 14 13 13 1 0 9 9 2
8 9 11 11 13 4 0 9 2
24 2 13 4 9 15 4 3 13 0 9 1 9 1 0 7 0 9 0 9 2 2 13 4 2
11 11 4 13 13 15 9 1 0 9 9 2
26 9 0 0 9 11 11 13 4 1 9 0 9 0 9 11 11 3 4 13 13 14 11 13 0 9 2
16 11 4 3 13 1 0 9 7 11 2 2 15 9 11 11 2
16 11 15 1 9 13 1 9 0 0 9 1 9 1 15 9 2
18 15 4 13 3 4 1 9 13 16 3 13 13 14 15 1 0 9 2
24 3 2 9 9 0 4 1 9 3 16 15 13 3 4 0 0 9 1 0 9 13 0 9 2
28 0 9 11 11 11 2 15 15 1 9 13 1 11 7 11 1 11 2 13 4 9 9 11 1 9 1 11 2
20 3 1 11 2 8 4 13 9 1 15 15 11 4 13 9 1 9 1 11 2
27 15 4 13 9 0 9 15 15 13 1 9 1 9 7 13 9 3 4 11 13 9 11 3 1 9 9 2
32 2 15 15 4 0 4 16 13 13 9 15 9 1 9 11 2 3 4 15 13 9 0 12 9 2 2 13 4 9 0 9 2
9 9 11 13 15 1 9 1 0 9
25 9 11 13 4 3 4 9 9 15 15 13 1 9 1 8 9 13 13 0 9 9 1 0 9 2
13 0 9 9 0 9 11 0 4 9 13 12 9 2
20 0 9 1 11 7 11 2 11 2 13 4 3 9 9 1 9 9 0 9 2
20 9 4 2 1 9 2 12 9 2 2 13 3 0 9 1 0 9 1 9 2
17 9 0 9 13 4 3 4 1 9 0 9 7 9 1 0 9 2
26 9 4 13 3 12 9 1 0 9 11 7 11 2 7 4 15 9 13 9 15 15 13 1 9 9 2
14 3 4 0 9 2 0 9 2 9 7 9 0 9 2
15 15 4 4 0 0 9 0 1 0 9 1 9 9 11 2
11 1 9 4 0 0 9 1 11 7 11 2
21 0 9 13 4 9 12 9 0 1 9 2 1 15 4 12 3 0 1 9 9 2
19 9 0 9 13 4 3 13 16 4 12 1 9 0 2 11 11 2 9 2
12 0 0 2 11 11 2 3 4 13 1 11 2
50 9 4 1 9 13 12 9 7 15 9 13 0 9 9 7 0 9 2 0 9 2 0 9 2 0 9 2 9 9 2 0 9 2 9 2 9 1 9 0 9 2 9 7 9 9 15 15 13 9 2
37 0 0 13 15 1 9 11 1 11 7 0 4 1 9 1 0 9 1 11 11 2 15 4 0 9 0 1 12 9 9 1 9 1 9 0 9 2
37 11 11 0 4 1 9 0 9 0 9 2 16 4 11 11 3 0 9 11 11 2 0 9 9 11 1 11 2 15 4 0 9 13 1 0 9 2
16 9 4 0 16 4 9 3 13 0 9 1 0 9 3 11 2
24 9 9 0 9 0 4 1 9 1 0 9 7 9 9 4 7 4 13 1 0 9 7 9 2
6 11 7 11 13 0 9
13 0 9 1 11 7 11 13 13 0 9 12 9 2
36 1 9 1 15 15 13 1 0 9 1 11 7 11 2 9 9 9 11 11 11 11 7 0 9 11 11 13 4 13 0 9 15 13 0 9 2
17 3 15 13 1 9 12 9 0 9 1 11 1 11 1 0 11 2
23 11 4 13 3 4 15 13 1 9 0 0 9 2 15 4 13 7 9 0 9 11 11 2
32 9 0 0 9 11 11 13 4 1 11 1 9 1 12 9 2 3 3 4 9 1 9 9 2 7 3 9 13 9 0 9 2
16 8 2 1 15 4 9 3 9 9 7 9 1 11 7 11 2
38 11 2 14 13 0 9 2 1 9 16 1 15 9 0 9 9 11 14 13 0 9 0 9 2 7 13 9 9 2 3 0 0 9 16 13 0 11 2
11 1 15 4 0 9 13 0 1 0 9 2
9 8 2 4 14 13 9 1 11 2
6 15 15 0 9 13 2
6 11 2 0 4 9 2
7 0 4 4 1 9 9 2
28 0 4 0 9 16 15 13 1 9 0 9 2 15 4 13 4 0 1 0 9 1 9 9 1 0 0 9 2
14 8 2 13 14 13 0 9 0 9 1 11 7 11 2
11 4 14 9 0 9 13 0 9 12 9 2
13 11 2 11 7 11 14 13 0 9 1 0 9 2
20 12 9 9 4 11 7 0 15 15 13 4 11 2 7 9 2 1 0 9 2
12 9 13 0 9 12 9 7 9 13 9 9 2
43 9 12 9 2 11 4 1 11 13 9 1 9 12 9 9 2 7 12 9 3 16 1 12 9 2 7 13 9 1 9 12 9 9 2 7 12 9 3 16 1 12 9 2
15 8 2 15 4 9 0 9 1 11 1 9 1 15 9 2
18 11 2 0 9 13 4 9 9 1 15 15 13 7 13 1 15 9 2
20 8 2 4 14 9 9 1 12 9 4 0 9 2 7 13 14 11 15 13 2
17 11 2 14 13 9 1 9 1 9 15 13 4 0 1 12 9 2
8 11 7 11 13 9 1 9 9
21 0 9 11 7 11 13 4 15 1 11 1 9 9 1 9 9 7 0 9 0 2
38 16 9 1 11 13 13 0 9 1 11 16 9 15 4 13 1 9 9 0 11 2 9 15 4 13 0 1 0 9 7 16 0 9 1 9 9 11 2
30 1 9 9 1 11 2 9 9 0 9 2 11 11 2 13 4 16 9 14 13 2 7 0 7 0 9 9 11 2 2
29 3 9 9 0 9 11 11 3 4 9 1 11 2 0 9 11 1 9 11 2 2 13 4 16 4 15 9 0 2
38 2 11 11 15 4 13 1 0 9 7 1 0 9 0 9 2 2 13 4 11 9 2 3 3 4 11 13 1 9 0 9 7 0 9 9 1 11 2
24 1 9 2 9 11 13 4 13 1 11 1 0 0 9 2 7 4 15 0 9 13 0 9 2
18 3 4 4 0 7 1 0 9 2 1 9 16 11 13 13 0 9 2
27 9 1 11 13 4 13 0 0 9 1 0 9 9 9 1 11 2 16 1 15 9 13 9 1 9 11 2
18 9 1 9 9 2 15 4 0 2 3 13 13 9 1 11 7 11 2
24 15 9 2 15 4 13 13 12 9 2 13 4 9 1 15 4 4 9 11 2 11 7 11 2
25 16 4 11 13 13 9 16 15 15 4 13 9 0 11 2 9 15 4 3 13 1 9 0 9 2
41 2 9 1 9 0 9 11 9 4 9 11 7 9 12 9 9 11 7 9 0 9 1 15 13 9 11 2 2 13 4 1 11 11 11 2 9 0 0 9 11 2
8 9 4 3 3 13 1 9 2
38 9 9 0 9 9 1 11 2 11 11 2 13 4 1 11 16 4 0 15 4 9 0 2 7 16 4 11 2 3 1 9 13 9 11 7 11 2 2
35 1 9 13 14 9 0 9 11 2 11 4 13 16 2 11 3 3 13 15 4 0 9 1 9 1 11 2 7 15 0 9 4 13 2 2
21 3 2 9 9 9 1 11 11 11 13 4 1 11 16 4 15 9 1 0 9 2
27 2 1 9 11 11 9 4 14 0 9 11 7 11 16 15 3 13 9 11 1 11 9 0 9 1 11 2
18 15 4 9 3 0 9 1 9 0 9 9 11 2 2 13 4 11 2
8 9 4 3 13 7 0 11 2
31 11 11 2 12 1 9 11 1 9 11 2 3 14 13 0 9 2 13 4 16 4 9 0 1 0 9 7 13 9 11 2
30 2 3 4 16 11 13 1 11 2 15 13 9 1 11 1 9 1 9 1 0 9 2 2 13 4 11 1 0 9 2
24 3 2 11 11 2 9 11 15 13 1 0 9 2 13 4 3 4 9 13 15 9 1 11 2
30 2 1 9 2 11 13 0 9 16 15 2 1 9 0 9 2 13 9 11 7 9 9 9 0 11 2 2 13 4 2
7 11 13 9 9 9 1 11
11 0 9 13 4 13 0 0 9 8 9 2
49 9 9 15 4 13 13 9 1 9 11 13 15 1 9 2 12 9 2 1 0 9 2 1 15 4 0 9 13 15 9 7 13 9 12 1 9 15 4 13 1 0 9 2 15 4 13 0 9 2
30 11 11 0 4 1 9 9 16 4 13 13 9 11 1 9 7 13 1 9 9 12 9 2 12 9 9 7 12 9 2
9 13 4 1 9 1 9 1 9 2
30 0 9 4 4 9 0 9 12 9 1 9 11 11 2 15 4 4 1 9 1 11 3 16 15 4 15 13 0 9 2
22 15 9 13 4 4 0 0 9 8 9 2 15 4 13 13 9 9 1 9 12 9 2
22 3 4 11 13 9 1 9 15 4 4 1 9 9 2 1 15 4 13 9 0 9 2
50 9 9 2 15 4 0 1 15 4 0 9 1 9 9 11 11 13 1 9 16 4 0 9 1 0 7 0 9 1 9 1 11 4 0 13 1 0 9 1 9 9 2 13 4 9 0 9 1 11 2
10 15 13 16 4 11 13 1 9 11 2
21 9 9 13 4 1 9 9 1 0 9 1 11 2 3 0 9 1 9 9 9 2
16 0 9 0 9 13 4 9 9 3 16 9 2 0 9 2 2
15 9 4 13 11 16 13 9 2 7 4 15 9 3 0 2
34 2 9 13 13 15 1 15 9 2 3 4 13 3 9 1 11 11 2 2 13 4 0 9 0 9 11 11 1 9 0 9 1 9 2
14 2 13 0 9 0 1 9 15 9 2 2 13 4 2
20 9 0 9 0 9 11 11 13 4 1 11 16 4 9 1 11 13 0 9 2
15 9 1 15 9 13 16 1 3 12 9 14 0 0 9 2
8 0 9 11 13 4 9 11 2
22 1 9 1 11 2 9 4 13 16 4 15 9 2 0 7 0 0 9 7 9 2 2
20 9 4 13 0 9 7 0 0 9 16 13 9 1 11 3 4 13 9 9 2
58 1 9 2 9 0 0 9 2 15 13 11 2 0 0 9 2 11 7 11 2 13 4 1 9 9 1 15 13 2 0 15 13 13 9 9 11 16 15 13 1 0 9 2 16 4 15 15 9 13 13 7 13 3 0 0 9 2 2
20 1 9 1 9 2 11 4 13 15 9 2 3 16 4 15 13 1 0 9 2
17 1 9 9 2 9 4 13 9 9 9 0 9 15 4 0 11 2
4 0 9 1 11
12 0 9 13 13 0 9 11 1 9 12 9 2
15 1 3 3 3 1 12 9 11 4 13 9 1 0 11 2
26 15 9 4 1 9 12 9 4 3 12 9 1 9 2 15 4 9 13 0 9 1 9 9 1 11 2
16 12 7 3 9 1 9 9 11 4 3 0 13 12 9 11 2
10 15 4 15 3 13 12 9 12 9 2
26 1 9 9 9 9 2 9 11 11 13 4 9 16 2 0 0 9 1 15 4 0 9 3 0 2 2
23 2 0 7 0 11 0 4 9 1 15 9 2 2 13 4 11 1 9 1 9 0 9 2
22 2 11 4 3 0 16 9 1 0 9 15 13 9 7 0 9 11 2 2 13 4 2
15 0 9 1 11 13 4 12 9 2 1 9 9 9 11 2
15 3 0 9 2 9 4 3 13 11 16 13 1 0 9 2
41 2 11 4 13 13 15 0 9 1 0 9 2 3 1 9 7 0 9 2 7 4 1 9 1 9 13 9 9 1 9 9 2 2 13 15 1 0 9 1 9 2
18 2 9 0 9 1 9 13 4 15 0 9 11 7 0 9 9 2 2
17 16 4 0 0 9 0 1 9 9 2 0 9 4 14 3 0 2
20 9 13 16 13 9 15 15 13 9 11 2 16 7 3 4 0 1 12 9 2
47 11 11 2 0 9 7 0 9 2 13 4 1 11 16 4 15 0 0 9 2 1 9 16 4 0 9 1 9 0 9 3 0 2 13 1 9 9 2 7 13 13 14 3 9 1 9 2
47 2 4 4 9 9 16 15 13 15 4 3 13 9 2 15 4 13 2 3 7 3 2 16 4 13 9 9 11 7 15 4 3 13 4 0 1 0 0 9 2 2 13 4 11 1 11 2
9 2 15 4 9 1 0 0 9 2
23 9 1 11 14 13 15 16 0 2 0 7 0 9 2 16 16 9 0 7 0 9 2 2
7 11 9 9 2 9 9 2
31 3 15 9 9 11 11 11 7 0 9 11 11 11 4 4 9 0 9 15 4 9 9 9 2 9 7 9 1 0 11 2
20 0 0 9 1 9 2 9 1 9 2 4 4 12 9 0 1 0 9 11 2
50 9 15 3 13 11 2 11 7 9 1 9 9 13 4 9 11 2 11 7 11 2 11 2 11 2 11 7 11 7 11 11 2 3 1 9 11 2 11 2 0 9 2 9 7 9 1 3 12 9 2
33 9 9 4 4 0 1 9 9 2 9 7 9 2 9 0 2 0 7 0 9 2 7 9 9 9 2 9 9 7 9 0 9 2
33 9 9 4 13 9 7 9 9 11 7 11 1 9 1 15 9 2 13 9 9 7 13 1 0 9 1 15 15 13 9 0 11 2
14 9 9 4 0 9 11 11 7 0 9 11 11 11 2
32 9 9 13 9 9 9 7 9 0 9 1 15 4 15 13 1 12 0 9 2 9 7 9 2 9 7 0 9 7 0 9 2
16 9 9 15 4 13 9 13 4 9 13 15 9 1 0 9 2
62 3 11 1 2 9 7 9 2 15 4 13 1 9 9 2 11 4 13 9 11 3 13 13 0 9 2 1 0 9 7 9 2 0 9 0 9 7 0 9 7 9 1 9 0 0 9 2 16 4 13 13 2 0 9 15 4 4 0 7 0 2 2
44 9 9 0 9 11 12 9 12 9 2 11 4 0 9 13 15 9 1 9 0 9 1 11 16 0 9 1 9 0 9 9 1 9 7 15 9 9 15 4 0 1 0 9 2
21 1 9 12 9 15 9 0 4 1 9 0 9 11 0 9 0 9 1 0 11 2
54 2 13 16 4 9 1 0 9 2 9 7 9 0 9 15 4 13 13 0 9 2 3 9 2 9 9 2 9 0 9 7 9 0 9 7 9 2 3 3 9 9 1 0 2 0 7 0 9 2 2 13 4 11 2
51 2 9 7 9 1 9 14 4 15 13 13 9 7 9 16 9 1 9 7 9 2 2 13 4 11 3 9 16 4 9 2 13 9 1 0 9 1 15 15 13 9 7 13 15 9 1 9 0 9 2 2
10 0 9 13 0 9 1 9 7 0 9
17 0 9 13 16 0 9 1 3 9 9 4 3 13 1 0 9 2
12 9 9 4 3 15 9 13 0 9 1 9 2
54 9 1 9 0 9 0 9 3 0 9 2 12 9 2 2 15 4 13 0 9 2 13 7 0 9 0 2 9 9 2 15 4 13 0 9 2 1 15 4 1 3 0 0 9 2 12 1 12 9 2 13 0 9 2
52 15 14 4 0 9 1 9 0 9 1 9 2 9 9 9 12 0 9 2 0 0 9 11 7 0 0 9 0 9 0 9 2 9 4 9 1 0 2 9 2 1 12 0 9 1 9 0 0 7 0 9 2
47 9 9 11 11 2 0 9 11 15 15 13 12 1 9 0 9 0 9 11 11 1 9 0 9 2 13 4 9 1 9 2 0 2 2 3 16 4 15 15 9 13 13 7 1 0 9 2
32 1 15 2 0 0 9 2 0 9 1 0 9 0 9 7 9 9 16 13 0 9 2 3 4 13 9 1 0 9 15 13 2
18 2 9 3 4 13 9 2 7 9 1 0 2 9 9 2 2 2 2
26 14 15 2 9 2 13 13 9 1 9 1 0 9 7 9 2 2 13 4 9 11 11 11 12 9 2
57 1 0 0 9 1 0 9 2 15 4 0 1 9 0 9 7 9 7 0 9 15 4 3 3 1 9 2 0 9 0 4 2 0 9 2 1 9 7 12 0 0 9 2 15 4 3 13 0 9 7 0 9 0 1 0 9 2
24 3 2 2 0 2 9 1 9 2 12 9 2 13 4 3 12 0 9 15 4 13 9 11 2
29 0 16 13 15 9 7 9 0 9 9 2 11 11 2 0 9 0 9 1 11 2 13 4 1 2 0 9 2 2
22 2 15 4 0 7 3 0 9 2 13 14 9 3 13 2 2 13 4 11 1 11 2
36 2 3 15 14 13 9 9 2 9 2 2 15 4 9 9 7 9 2 2 13 4 2 7 4 3 13 2 9 1 9 2 15 4 13 9 2
14 3 4 13 0 9 16 4 0 2 0 9 2 0 2
22 11 11 2 0 9 7 9 2 7 9 0 9 0 9 2 14 13 15 7 13 9 2
42 2 3 2 0 9 16 15 13 7 13 0 9 1 15 9 4 16 15 13 9 1 12 9 7 16 15 3 3 13 2 7 16 15 0 9 3 13 16 13 9 2 2
25 8 4 13 16 15 13 3 1 0 9 1 0 9 1 3 15 13 1 11 1 3 1 12 9 2
83 1 9 2 0 9 2 1 0 0 9 2 15 4 1 15 9 13 0 0 9 2 1 0 9 4 9 9 0 1 9 1 0 9 2 9 1 9 9 3 4 15 13 9 0 9 0 1 9 2 0 9 9 15 9 2 9 9 0 1 9 9 2 9 7 9 0 9 2 9 9 7 9 1 9 2 7 9 0 9 1 0 9 2
12 0 9 13 4 15 15 1 9 2 13 11 2
8 0 4 4 0 1 9 9 2
6 9 1 9 1 11 2
26 11 13 13 1 9 1 12 0 9 2 11 2 11 2 11 11 7 11 2 1 9 16 13 9 9 2
21 11 7 11 13 4 1 9 2 12 9 2 9 1 9 1 9 9 1 9 9 2
26 15 9 2 13 9 2 0 4 9 16 11 13 13 0 9 1 9 3 4 9 1 9 9 1 9 2
24 2 9 11 16 4 0 9 1 15 9 4 0 2 2 13 4 1 11 0 0 9 11 11 2
20 9 4 13 0 9 0 9 11 11 7 9 0 0 9 1 9 9 11 11 2
15 9 9 13 4 1 0 7 0 9 15 13 9 7 9 2
15 11 4 3 13 0 9 1 9 1 9 1 11 7 11 2
31 1 0 9 11 11 13 15 16 15 9 13 13 0 2 9 2 2 15 4 13 11 2 11 2 11 11 2 11 7 11 2
14 9 4 13 3 16 4 13 9 9 15 13 1 11 2
12 2 0 9 9 4 4 0 0 9 0 9 2
16 11 2 3 2 13 9 0 9 1 0 7 0 9 1 11 2
21 0 9 1 9 13 9 16 0 9 13 4 0 1 9 2 2 13 15 1 9 2
5 9 4 3 0 2
28 11 4 0 9 13 16 4 2 16 0 9 14 13 0 9 1 9 9 2 0 9 13 3 12 9 9 3 2
48 11 2 4 12 1 0 9 15 13 9 15 9 2 3 15 0 9 15 15 13 1 11 2 11 2 11 7 0 0 9 11 13 12 1 0 9 15 15 13 1 15 9 2 2 13 4 11 2
33 11 4 13 16 4 15 9 1 9 1 9 2 9 2 1 11 2 3 3 15 4 1 0 9 0 16 9 1 2 0 2 9 2
33 2 9 1 11 3 4 13 15 9 7 9 16 15 3 13 1 9 9 2 2 13 11 2 3 16 4 9 13 3 15 13 11 2
11 7 2 11 4 13 11 1 15 9 9 2
11 2 13 3 12 9 15 13 11 7 11 2
9 15 1 15 13 0 9 7 9 2
10 11 13 16 9 9 9 1 0 9 2
39 11 4 13 9 11 2 16 1 9 0 9 2 3 15 13 0 9 9 2 15 15 3 13 1 9 7 13 2 2 13 4 11 2 7 13 0 11 11 2
19 9 4 13 9 9 2 9 9 1 0 9 7 9 0 9 9 15 9 2
13 9 11 1 9 1 9 2 11 0 2 7 9 13
19 9 11 8 11 7 9 0 0 9 11 13 4 15 9 2 7 9 13 2
34 0 9 0 15 1 0 0 9 1 12 9 3 4 3 0 2 13 4 9 11 1 9 1 9 11 8 11 1 9 2 12 9 2 2
36 3 2 9 1 11 7 0 9 7 3 15 13 1 9 2 13 4 2 3 16 12 1 15 9 16 0 9 13 9 1 0 9 1 0 9 2
10 2 13 14 15 16 4 3 1 9 2
4 3 14 2 2
37 11 4 3 0 9 15 9 11 8 11 9 9 2 9 0 0 9 9 7 0 9 1 15 15 2 3 15 13 2 13 2 13 4 15 9 11 2
25 2 3 4 3 3 0 3 16 15 4 4 1 12 9 2 2 13 4 9 1 11 2 13 11 2
35 2 15 14 13 16 4 13 0 9 2 0 9 2 7 4 13 4 0 1 9 2 1 9 7 0 9 9 7 1 9 9 0 9 2 2
16 9 1 0 9 3 0 9 13 4 7 1 9 2 1 11 2
20 9 15 9 13 4 16 4 13 9 9 11 0 9 1 9 11 1 9 9 2
36 1 9 15 4 13 0 9 2 15 4 13 1 9 1 11 2 4 4 7 11 11 2 15 4 0 9 4 13 9 1 9 0 9 3 9 2
41 2 11 4 3 1 11 8 11 13 9 16 15 13 1 9 9 1 0 9 1 0 0 9 2 11 7 11 2 2 13 15 1 9 0 9 2 13 0 8 8 2
37 2 13 4 9 1 0 9 1 0 0 9 2 3 9 7 9 2 9 9 2 16 7 9 1 9 7 9 1 9 9 0 9 1 0 9 2 2
23 0 9 1 15 15 9 13 3 13 4 2 3 0 7 0 2 2 13 4 9 1 11 2
40 9 11 1 9 13 4 9 16 4 0 0 9 1 11 3 13 9 0 9 11 16 13 15 9 9 9 2 3 9 9 2 15 15 3 13 1 9 9 9 2
29 2 13 4 9 9 9 2 3 0 9 7 9 2 7 0 9 9 2 15 4 3 0 2 2 13 4 8 11 2
37 0 9 15 2 1 15 9 2 13 2 3 13 11 2 4 2 9 0 9 1 11 7 11 2 1 0 9 15 4 13 15 12 9 3 15 9 2
23 2 14 13 13 0 9 2 2 13 4 8 11 2 3 1 9 9 9 9 1 15 9 2
5 0 9 11 1 11
28 0 9 0 1 0 9 11 1 11 13 7 9 1 9 9 9 0 9 9 7 9 1 9 9 9 1 11 2
20 0 9 9 9 7 9 9 9 11 1 11 0 4 1 9 2 12 9 2 2
25 1 0 9 0 1 0 9 9 4 1 9 9 9 0 9 9 7 9 1 9 9 9 1 11 2
34 9 0 9 13 4 9 9 1 11 1 0 9 0 0 9 1 0 9 2 15 4 0 1 9 2 12 9 1 16 15 4 4 0 2
19 13 4 15 13 0 9 1 9 15 9 9 7 13 9 0 9 0 9 2
10 9 4 0 1 0 9 1 9 11 2
22 0 9 11 11 13 1 15 16 9 9 9 11 13 1 0 9 2 7 14 9 11 2
26 2 13 9 13 3 7 13 2 0 0 9 4 13 2 2 4 13 2 2 13 4 0 9 11 11 2
13 1 15 2 9 4 13 9 0 9 11 1 11 2
25 9 9 3 4 15 13 13 0 12 9 1 0 0 9 1 9 1 11 2 15 3 13 12 9 2
35 9 11 11 11 13 4 0 9 9 7 13 11 1 0 9 0 0 9 3 4 15 13 9 1 15 9 1 0 7 0 9 0 1 9 2
17 2 9 11 15 4 9 0 3 2 14 3 2 2 13 4 11 2
16 9 9 1 11 2 0 9 11 11 11 13 15 9 9 11 2
35 16 4 11 13 1 9 1 9 1 15 9 7 13 13 0 9 2 1 9 4 15 13 13 9 11 7 0 9 2 15 13 11 7 11 2
28 2 15 9 1 0 9 13 9 1 0 9 1 0 9 9 7 14 13 4 9 15 2 2 13 4 0 9 2
20 2 3 13 1 9 9 2 0 9 9 7 0 9 4 15 15 13 1 9 2
17 14 13 15 0 1 0 9 7 0 9 9 2 2 13 4 11 2
13 9 11 4 3 3 13 9 11 1 9 1 11 2
13 2 16 0 9 11 13 9 2 2 13 4 11 2
25 2 15 9 3 4 4 1 0 9 1 9 1 0 9 7 9 2 16 4 15 9 12 9 2 2
23 9 11 1 9 3 4 13 9 1 9 9 11 1 11 7 11 1 9 11 1 9 9 2
38 1 15 2 12 9 15 15 13 9 1 9 2 11 2 11 7 11 2 0 4 1 9 15 4 3 13 2 16 15 4 0 3 4 13 13 9 11 2
12 9 11 13 16 4 0 0 9 0 9 1 11
28 3 4 9 1 9 0 9 9 1 0 9 11 2 13 4 1 9 0 9 11 2 3 1 0 9 1 9 2
24 9 11 1 0 9 11 11 2 3 2 13 15 1 9 0 11 11 11 11 1 9 0 9 2
38 0 9 11 13 4 1 9 2 12 9 2 9 9 16 2 16 7 0 11 7 0 11 13 9 15 4 15 13 9 11 2 14 13 13 0 9 9 2
36 2 0 9 0 0 9 14 4 4 0 2 2 13 4 9 11 1 0 9 11 11 3 9 9 1 15 9 11 2 11 7 11 3 15 9 2
28 2 15 0 14 4 13 0 9 15 4 15 13 2 16 15 4 15 13 0 12 2 0 9 7 0 9 2 2
28 0 0 9 1 9 11 13 4 1 9 0 9 2 3 4 0 11 1 0 9 13 9 9 15 4 13 11 2
30 16 4 9 0 11 13 0 9 2 3 4 3 0 9 0 9 1 9 0 11 1 9 13 1 11 12 9 12 9 2
32 11 4 13 16 4 1 3 13 1 0 9 2 3 2 0 9 2 15 4 13 9 0 11 7 0 11 1 9 9 0 9 2
34 2 13 0 9 7 1 0 9 2 16 1 9 1 0 9 2 3 7 1 0 9 15 3 13 13 1 0 9 2 2 13 4 11 2
26 1 9 9 2 13 4 2 13 15 9 16 13 0 9 1 9 12 9 2 7 7 0 9 4 0 2
17 16 0 9 13 16 13 9 2 13 9 1 9 9 2 13 4 2
35 2 9 1 9 13 13 2 7 0 9 13 13 9 2 9 7 0 9 0 1 9 9 2 1 0 9 15 13 9 2 2 13 4 11 2
12 9 13 13 2 7 14 3 13 15 9 2 2
51 9 0 11 11 11 13 16 4 9 15 4 0 9 13 0 9 11 11 11 9 0 11 7 11 0 2 3 15 15 4 13 2 3 16 15 4 4 0 2 7 3 16 4 0 2 2 13 4 11 9 2
47 9 0 11 11 11 11 1 9 4 13 16 4 15 9 4 2 0 13 0 9 1 9 9 2 16 16 13 16 4 3 0 13 0 7 0 9 9 9 0 11 2 2 13 4 9 11 2
28 11 4 3 13 9 15 9 9 4 13 1 0 0 9 1 12 9 0 9 7 13 9 15 4 0 0 11 2
22 11 4 13 16 15 2 3 1 9 9 2 13 13 2 3 3 2 1 9 1 9 2
7 0 9 1 0 9 0 9
27 0 9 0 7 0 9 13 4 1 0 12 9 1 3 12 9 2 7 3 3 13 3 9 1 0 9 2
22 3 11 3 4 1 9 3 12 9 2 1 9 1 12 3 15 4 4 1 12 9 2
28 1 12 9 2 3 4 12 0 9 13 0 0 9 1 11 2 3 4 12 9 1 9 11 13 13 0 9 2
19 3 15 1 9 11 13 3 12 9 0 7 0 9 7 15 15 9 13 2
22 1 0 9 11 0 9 2 11 2 2 1 0 12 9 0 4 3 12 9 0 9 2
20 0 9 9 13 4 3 12 9 2 1 11 4 4 3 0 2 3 12 9 2
24 9 13 16 4 2 16 15 13 15 9 2 11 1 9 9 13 13 12 9 0 9 1 9 2
21 9 9 4 3 13 2 1 12 9 9 1 12 9 2 1 12 9 1 12 9 2
13 3 1 0 9 12 9 3 4 13 12 9 9 2
14 9 13 16 0 2 3 16 0 9 2 13 0 9 2
26 3 15 13 3 12 9 0 9 9 1 11 2 16 4 15 15 9 13 13 1 9 2 13 9 9 2
13 15 9 13 4 7 15 9 2 3 9 9 9 2
20 3 13 3 12 9 3 11 2 1 9 1 12 3 15 4 4 1 12 9 2
36 9 15 15 13 9 7 0 9 4 4 0 13 1 9 1 0 9 2 11 2 2 7 1 9 12 9 1 9 4 4 3 1 12 15 9 2
18 16 0 9 11 7 11 13 0 9 2 7 9 9 13 13 15 9 2
9 0 9 1 9 3 4 1 9 2
29 0 1 3 1 9 9 2 1 9 11 11 3 4 13 12 9 9 1 9 2 15 4 11 13 9 1 0 11 2
18 16 4 3 1 9 13 0 9 0 0 9 2 13 0 9 1 9 2
18 15 13 9 3 12 9 1 9 9 1 9 15 4 0 9 1 11 2
28 0 13 16 4 9 9 2 15 3 13 3 1 12 9 0 0 9 2 13 13 12 1 12 9 1 12 9 2
9 3 2 15 11 7 3 4 0 2
13 2 13 13 9 1 0 9 2 1 9 15 9 2
13 3 14 13 9 2 2 13 11 11 2 0 9 2
9 2 3 15 13 1 9 1 9 2
26 16 13 1 9 7 1 9 7 15 9 14 13 2 3 4 15 13 2 2 13 11 11 2 0 9 2
28 15 9 4 0 0 9 0 1 0 9 2 3 9 0 9 1 12 9 11 2 15 4 13 9 1 9 9 2
26 15 4 9 16 4 15 0 0 9 15 4 13 0 9 9 9 1 9 9 15 9 3 13 0 9 2
8 0 0 9 1 11 4 4 0
40 9 2 9 1 9 0 9 7 0 0 9 13 9 16 4 13 13 9 1 9 0 9 0 12 9 2 15 4 13 4 0 1 9 15 9 9 1 0 9 2
23 0 0 0 9 1 9 2 11 2 4 4 0 3 9 11 13 1 9 1 9 15 9 2
21 9 2 15 15 13 1 0 9 0 0 9 2 4 4 0 1 3 12 9 9 2
15 16 14 4 0 0 9 2 11 4 13 13 0 0 9 2
32 16 4 13 9 9 0 12 9 2 9 1 9 0 9 7 0 9 13 4 9 9 11 2 1 9 2 14 13 9 11 2 2
17 2 9 0 12 9 13 15 1 9 15 4 13 12 1 12 9 2
32 14 13 16 9 14 13 13 2 16 9 4 15 13 13 1 9 15 4 15 13 9 11 2 2 13 4 9 9 11 11 11 2
29 9 4 13 9 11 2 15 4 3 13 3 13 9 1 11 0 1 9 9 2 1 9 15 9 2 9 12 2 2
41 0 9 1 9 2 0 9 15 13 3 1 12 0 9 2 13 15 0 9 7 11 7 13 9 0 9 0 9 11 11 2 3 9 1 9 11 7 15 0 9 2
35 3 2 1 3 4 0 9 13 15 0 9 13 9 1 0 9 2 9 4 13 0 9 1 9 9 0 1 15 9 3 16 15 15 13 2
28 1 12 9 0 4 0 9 9 2 9 9 2 0 9 7 0 9 2 15 13 1 0 7 14 1 0 9 2
30 0 9 1 9 2 11 2 13 4 9 1 15 9 2 3 16 15 0 9 13 1 9 16 15 14 4 13 1 9 2
11 9 13 16 4 15 15 3 13 0 9 2
15 0 9 15 15 13 4 9 9 1 0 9 1 0 9 2
21 9 1 15 9 2 1 15 0 9 13 1 9 1 9 2 3 13 1 15 15 2
9 9 4 15 13 9 0 1 9 2
20 3 2 9 11 3 4 15 13 9 0 0 9 2 16 7 9 1 9 9 2
15 11 4 1 9 4 0 16 2 0 9 9 9 11 2 2
18 0 1 0 9 2 9 4 13 9 1 12 9 1 9 0 9 11 2
25 1 12 9 9 4 13 9 0 0 9 2 1 0 9 7 0 0 9 1 12 1 12 9 11 2
38 1 0 9 0 4 9 0 9 2 9 1 3 0 0 9 2 9 2 9 1 3 0 9 2 0 9 2 0 9 7 9 2 9 1 9 1 9 2
22 0 9 4 4 1 3 0 3 0 1 15 0 9 2 3 15 4 4 0 0 9 2
6 0 9 0 9 1 11
18 16 4 0 9 1 9 1 11 2 0 9 9 0 9 13 0 9 2
43 0 9 13 4 16 15 2 1 0 9 12 9 2 9 9 1 9 0 9 1 11 13 1 0 9 1 9 0 0 9 2 0 11 7 0 9 1 0 9 9 0 9 2
13 0 9 9 9 0 9 1 9 9 14 13 0 2
16 9 1 15 4 0 2 7 13 9 9 1 0 7 0 9 2
19 0 4 0 9 9 15 3 13 1 9 7 3 0 9 9 1 9 9 2
16 0 9 14 13 13 9 1 0 7 0 9 7 1 9 9 2
13 0 9 9 7 0 9 3 13 9 1 9 9 2
47 3 2 9 1 0 9 2 9 1 0 9 2 11 1 0 9 7 9 7 11 1 9 0 9 2 11 2 1 9 1 0 9 1 9 2 15 4 1 0 9 15 13 9 9 0 9 2
10 1 12 2 15 13 0 0 9 9 2
32 0 9 13 9 1 9 9 9 0 9 9 0 9 2 9 1 0 9 2 9 9 2 9 0 0 9 1 9 7 0 9 2
24 2 1 12 9 0 4 12 9 1 0 9 15 4 13 9 2 1 9 1 0 7 0 9 2
22 1 12 2 0 4 12 9 0 9 2 16 4 1 0 9 15 9 0 12 0 9 2
29 16 4 15 9 1 9 2 3 4 0 9 1 15 0 9 2 2 13 4 11 11 11 1 9 0 1 0 9 2
35 9 0 7 0 9 11 11 7 11 11 2 7 0 9 1 11 11 11 2 13 4 15 9 15 4 13 13 16 0 9 1 9 0 9 2
9 2 9 4 0 9 9 1 9 2
11 9 15 9 14 4 13 13 9 0 9 2
23 3 2 1 11 2 9 13 9 15 15 9 13 9 9 7 0 9 2 2 13 4 11 2
38 2 1 15 4 9 1 9 0 9 1 9 9 2 9 7 9 2 7 16 4 13 1 0 9 2 13 15 13 9 1 9 9 2 0 7 0 9 2
35 0 0 9 1 0 4 9 2 7 1 0 9 13 4 3 3 3 15 13 13 9 7 3 15 13 9 7 9 9 2 2 13 4 11 2
19 9 0 9 9 0 9 13 4 3 9 16 13 15 9 1 9 0 9 2
10 11 1 0 9 1 9 11 7 0 11
28 16 9 1 11 7 11 13 4 15 9 9 1 11 1 9 1 11 7 0 11 2 11 15 13 1 0 9 2
34 9 11 11 11 13 4 1 9 2 12 9 2 16 15 9 15 9 14 13 13 1 4 15 0 9 1 9 2 3 11 7 0 11 2
20 11 4 13 16 4 11 0 9 2 1 0 0 2 0 2 0 7 0 9 2
29 2 15 15 15 13 9 11 13 13 11 16 9 0 9 2 7 13 16 9 13 15 3 0 2 2 13 4 11 2
18 9 9 11 11 13 4 15 9 2 3 16 4 11 2 0 9 2 2
10 11 15 2 3 2 13 1 0 9 2
34 16 11 13 15 2 0 9 2 2 7 11 13 9 15 13 13 9 1 0 9 2 11 13 9 1 0 9 7 9 15 9 1 11 2
29 2 4 4 3 1 11 16 9 1 11 13 1 15 0 9 1 9 11 2 2 0 4 1 0 9 11 1 9 2
12 2 3 2 11 4 15 13 13 1 0 9 2
26 13 4 13 9 0 9 2 15 4 13 1 9 1 0 9 2 1 15 9 11 13 1 0 9 9 2
22 2 9 9 0 11 7 11 4 2 3 2 13 9 11 1 9 11 2 2 13 11 2
19 0 9 1 11 11 11 13 4 16 4 9 13 2 9 2 1 12 9 2
19 2 0 9 14 13 15 13 9 2 9 7 9 0 9 2 2 13 4 2
14 1 0 9 11 11 2 9 11 7 11 4 3 0 2
12 2 13 9 1 15 4 0 2 2 13 4 2
21 2 11 4 4 1 0 9 1 0 9 2 4 4 0 9 3 1 9 0 9 2
36 9 0 9 1 9 4 0 2 3 7 1 15 15 15 15 14 13 7 15 14 13 2 2 13 4 11 2 9 0 9 1 0 9 7 9 2
22 1 9 2 11 0 11 13 9 11 1 0 9 2 16 7 13 16 4 11 0 9 2
23 11 3 13 9 7 9 11 7 13 9 4 15 9 1 11 2 13 4 0 9 11 11 2
13 9 14 13 4 0 1 9 0 9 2 13 4 2
25 2 3 13 9 2 16 7 15 9 13 2 16 15 13 0 9 2 3 4 0 9 3 0 2 2
12 9 0 9 13 4 0 0 1 9 0 9 2
9 9 11 13 9 9 9 9 1 11
40 9 0 9 11 13 4 15 1 9 16 4 13 9 9 1 11 2 15 4 13 9 9 1 15 9 2 3 9 3 0 9 9 12 9 7 11 4 4 0 2
21 9 1 9 13 1 9 0 9 2 12 9 1 11 2 1 9 2 12 9 2 2
40 11 4 1 9 2 12 9 2 13 16 4 0 13 9 1 0 0 9 0 11 2 1 9 9 9 9 1 9 9 15 4 11 7 11 13 7 12 9 3 2
42 2 11 13 4 0 2 2 2 13 0 9 2 3 9 0 9 7 11 2 0 1 0 7 9 9 9 1 11 2 2 13 4 9 0 9 11 1 0 9 1 11 2
40 9 1 12 9 2 15 4 13 0 9 11 11 2 15 4 9 0 9 0 0 9 11 2 13 15 16 11 7 11 13 13 1 9 7 13 0 9 0 9 2
21 1 15 2 0 9 13 15 13 1 15 0 9 2 7 0 9 1 9 1 9 2
20 9 4 0 0 9 1 9 7 9 1 0 11 7 11 2 0 0 0 9 2
28 0 9 13 15 0 9 1 15 4 11 13 0 9 1 0 11 2 15 15 13 1 11 12 7 13 9 11 2
13 11 4 3 13 2 3 11 7 1 9 0 11 2
46 3 11 2 0 9 0 9 11 11 13 4 16 4 9 0 9 1 0 9 11 7 0 9 1 0 0 9 11 2 0 9 1 9 2 2 2 1 15 4 15 13 16 4 13 2 2
22 9 15 11 13 13 1 0 11 13 4 15 12 9 11 15 15 3 13 1 15 9 2
21 0 9 0 9 11 11 2 0 9 11 2 13 4 16 4 13 9 3 12 9 2
28 0 9 0 9 11 11 2 15 4 1 9 13 9 2 13 4 16 15 13 16 15 11 4 13 0 9 11 2
24 13 4 2 3 2 16 15 0 9 11 13 13 9 0 9 9 2 1 15 11 13 9 9 2
39 9 0 9 11 9 9 13 4 16 4 13 9 9 0 9 1 0 9 9 0 9 9 9 11 2 15 4 15 12 7 12 9 13 1 11 2 1 11 2
17 3 0 9 9 13 4 1 9 9 1 11 1 15 9 1 11 2
20 2 3 2 15 9 13 13 15 9 2 2 13 4 0 9 0 9 11 11 2
14 11 4 2 3 2 13 1 9 11 7 9 1 9 2
15 9 4 4 9 0 9 9 0 9 9 9 11 0 9 2
33 0 0 9 11 11 13 4 9 2 1 9 9 2 2 2 1 9 0 0 9 1 11 2 2 13 4 9 11 1 11 1 9 2
49 1 9 2 9 9 11 2 11 2 11 2 11 7 11 2 7 11 2 15 4 9 11 2 13 4 9 12 9 16 11 13 1 0 9 1 9 1 11 16 4 15 13 0 9 11 1 15 9 2
11 9 2 9 13 16 13 9 11 0 1 9
21 3 1 12 9 11 13 16 4 13 0 2 7 0 15 9 13 7 1 0 9 2
16 1 0 9 1 9 2 0 0 9 13 0 9 1 9 11 2
6 9 13 9 1 11 2
15 1 11 13 9 9 16 9 0 0 9 7 9 0 9 2
29 12 11 13 16 4 9 1 9 0 2 13 15 1 9 9 1 0 9 0 0 9 2 0 1 9 2 12 9 2
14 1 11 12 9 13 16 4 0 1 9 1 0 9 2
18 11 4 0 1 12 2 16 12 9 1 11 13 16 15 15 9 13 2
15 1 11 4 12 9 13 9 15 0 9 1 0 12 9 2
12 0 9 8 8 13 4 12 9 9 1 11 2
14 0 4 0 9 4 1 9 1 11 1 11 1 11 2
20 9 4 13 12 9 3 2 7 13 15 16 4 1 9 9 13 1 12 9 2
20 0 9 11 11 13 4 0 0 9 1 9 11 1 11 1 9 2 12 9 2
18 9 9 0 4 1 12 9 9 2 7 4 4 0 12 0 0 9 2
26 0 9 0 9 4 3 12 9 9 7 12 9 9 2 15 4 13 4 0 0 0 9 15 9 9 2
23 0 9 11 11 7 15 0 9 11 11 13 4 0 0 9 1 9 0 12 9 1 11 2
19 11 4 13 16 13 16 4 9 3 13 9 1 9 11 1 9 0 9 2
12 9 4 13 0 9 1 0 9 1 0 11 2
12 11 4 1 9 1 11 13 9 0 0 9 2
23 0 9 11 11 7 15 9 11 11 13 4 1 9 2 12 9 2 1 11 0 0 9 2
10 13 4 15 1 0 9 0 0 9 2
14 3 1 9 0 4 7 9 9 1 9 0 0 9 2
33 0 0 9 11 7 0 11 13 4 0 9 0 9 1 9 11 1 0 9 0 9 0 11 2 13 4 11 1 9 2 12 9 2
9 0 9 9 0 9 0 4 12 2
14 12 9 13 0 9 1 12 2 7 13 9 7 9 2
22 0 9 9 7 0 9 11 11 13 4 1 9 2 12 9 2 9 1 0 9 9 2
31 9 4 15 13 1 12 9 1 12 9 11 2 7 0 4 1 9 9 0 9 1 9 1 9 2 15 15 13 9 9 2
34 0 9 4 1 9 2 12 9 2 13 0 9 15 15 13 9 9 15 0 9 13 13 1 0 9 7 15 13 0 9 1 0 9 2
21 1 0 9 2 0 9 13 13 1 12 15 9 1 9 2 1 9 1 0 12 2
19 9 1 9 7 0 9 7 9 1 0 9 13 4 15 1 9 1 12 2
21 9 1 9 1 0 9 4 4 0 1 12 1 12 16 4 15 13 9 9 9 2
9 9 4 9 0 9 1 9 9 2
9 0 9 2 2 0 9 2 13 11
22 0 0 9 0 4 1 15 9 1 9 2 7 1 0 4 9 9 13 11 7 11 2
30 11 11 1 11 11 13 1 9 11 11 1 11 1 0 0 9 1 0 0 9 1 11 2 1 9 2 12 9 2 2
12 0 0 9 13 4 11 1 9 12 2 12 2
26 11 11 2 11 11 2 11 11 7 11 11 13 4 12 9 2 16 4 11 11 7 11 11 13 12 2
11 11 11 4 4 0 0 9 1 12 9 2
25 0 9 0 9 11 11 13 4 1 9 1 12 9 15 9 1 11 11 11 1 9 12 2 12 2
21 1 9 1 12 11 2 11 11 13 4 1 11 11 1 0 9 2 12 2 12 2
14 0 9 13 4 1 9 1 11 1 9 12 2 12 2
24 11 11 13 4 12 9 2 16 4 1 12 13 11 11 2 11 11 2 11 11 7 11 11 2
11 1 12 9 13 4 11 11 7 11 11 2
20 0 0 9 11 11 12 4 9 13 1 9 2 7 3 4 12 13 1 9 2
30 1 9 1 9 1 9 2 11 11 11 7 11 11 4 4 0 1 11 11 11 7 11 11 2 1 9 12 2 12 2
15 0 9 2 11 11 7 11 11 2 13 4 1 0 9 2
21 1 9 2 11 11 13 4 1 11 11 11 1 0 9 1 9 1 9 9 9 2
19 1 9 0 9 2 11 11 13 4 1 11 11 11 1 9 1 12 11 2
14 1 9 2 11 11 4 4 0 0 9 1 0 9 2
14 13 4 1 12 9 2 16 4 9 4 11 11 11 2
14 1 9 9 2 11 4 13 1 11 11 12 2 12 2
25 0 9 13 4 1 9 0 0 9 1 9 12 2 12 2 1 9 1 3 9 15 4 13 9 2
26 11 11 2 11 11 2 11 11 7 11 11 13 4 1 12 9 2 11 11 13 4 12 9 1 11 2
10 0 9 13 4 1 11 12 2 12 2
33 11 4 13 0 9 1 15 4 9 9 11 11 1 9 13 1 9 1 9 1 12 11 2 14 3 1 12 9 9 13 12 11 2
7 11 4 13 9 0 9 2
43 1 9 2 11 11 13 4 3 1 12 9 2 16 4 9 11 11 0 1 9 0 9 1 12 9 3 2 3 3 1 12 9 1 12 9 1 9 12 2 12 2 12 2
35 3 9 9 2 9 0 9 11 11 7 11 11 13 4 1 9 1 12 11 7 12 11 2 16 4 9 11 11 13 1 9 1 12 11 2
7 9 7 9 2 11 1 11
21 9 2 9 9 7 9 9 11 2 4 4 15 1 0 9 1 11 15 0 9 2
36 3 1 9 9 1 9 7 9 2 11 11 1 0 9 9 0 9 11 7 11 2 11 11 13 9 9 0 1 15 9 2 9 1 9 2 2
24 9 13 1 9 11 7 9 1 9 9 11 0 1 9 1 9 11 1 9 2 12 9 2 2
19 11 4 12 0 9 13 1 0 9 1 11 2 3 12 9 7 9 9 2
22 9 11 11 11 3 4 13 0 9 2 3 9 1 0 0 9 1 9 11 12 9 2
19 9 11 13 4 9 1 15 9 2 3 4 9 13 13 9 16 13 9 2
46 9 11 11 2 9 0 9 11 11 11 7 9 11 11 4 4 1 12 0 9 15 4 9 11 11 13 1 15 9 1 9 9 2 9 2 9 2 9 2 9 7 9 1 12 9 2
17 11 4 13 0 9 11 11 2 16 4 0 9 0 9 0 9 2
18 0 9 11 7 11 2 11 2 13 4 9 11 11 1 9 0 9 2
12 11 4 3 4 9 9 1 12 1 12 9 2
20 13 11 11 2 15 4 3 15 9 0 1 0 9 9 1 9 1 11 12 2
15 9 9 0 9 11 11 0 4 1 9 0 9 1 11 2
12 9 13 12 9 1 9 0 1 12 0 9 2
7 9 4 13 1 12 9 2
33 9 11 11 13 4 16 4 9 9 0 1 15 9 1 12 9 2 9 1 8 2 4 0 1 9 11 1 11 12 9 12 9 2
16 9 4 13 8 9 8 8 8 2 1 15 11 13 0 9 2
5 0 11 13 0 9
38 3 9 11 7 9 11 0 4 1 9 1 9 1 0 9 1 3 0 9 11 1 11 2 1 0 9 1 3 4 11 13 9 1 11 1 12 9 2
16 0 11 13 9 1 9 11 1 9 2 12 9 2 1 11 2
32 9 11 1 11 13 4 1 9 2 12 9 2 15 0 9 1 9 3 0 9 11 0 11 1 15 4 13 9 1 0 9 2
12 0 4 0 9 0 9 15 13 1 9 11 2
32 2 13 9 1 0 9 0 9 7 15 9 15 4 0 1 9 11 7 11 2 2 13 4 1 11 1 11 9 11 11 11 2
29 11 4 3 13 16 4 2 3 0 0 9 2 1 9 1 9 11 9 1 9 11 1 9 15 9 1 15 9 2
37 2 13 0 9 9 3 2 16 15 4 3 0 9 7 3 4 9 9 2 1 9 16 15 13 2 13 13 11 9 1 15 9 2 13 4 11 2
27 15 4 0 1 15 4 15 9 11 13 1 0 9 2 15 4 13 9 0 9 9 1 11 1 9 11 2
13 12 9 3 3 12 0 0 9 3 4 13 9 2
31 0 9 0 4 2 3 15 13 2 9 9 15 4 13 0 9 1 15 4 11 13 1 9 11 1 9 9 12 2 12 2
21 16 4 13 9 2 13 4 9 11 1 9 7 13 9 11 2 3 15 9 11 2
23 9 11 13 4 1 9 9 1 9 1 9 13 15 16 13 9 2 16 4 9 15 13 2
45 3 9 9 11 7 9 11 13 4 2 3 15 13 2 1 9 1 9 0 1 9 2 15 4 0 1 15 4 0 0 9 13 9 1 0 9 1 9 11 1 15 3 13 11 2
31 3 15 13 12 11 0 4 1 9 9 2 16 2 3 15 13 2 3 12 15 13 4 1 15 4 0 9 13 9 11 2
7 11 4 13 9 12 9 2
31 0 9 1 3 13 13 15 9 2 3 1 3 9 11 7 0 9 2 3 2 9 9 2 9 0 9 1 9 0 9 2
35 2 9 4 3 0 2 16 9 7 9 11 0 4 1 0 9 2 2 13 4 11 9 9 0 0 9 2 11 2 1 9 2 11 11 2
9 11 4 0 0 9 0 12 9 2
27 1 9 2 9 0 9 13 15 1 9 9 3 9 7 9 1 9 0 9 15 4 13 1 9 1 9 2
12 15 4 13 9 7 0 9 16 4 13 0 2
23 12 9 11 7 12 9 11 0 4 1 9 7 0 2 13 15 1 9 0 0 0 9 2
28 11 13 16 4 9 2 15 15 13 1 9 9 11 1 9 9 2 2 4 1 0 9 2 0 1 9 9 2
31 1 9 15 4 3 13 11 0 4 9 9 15 4 13 16 4 1 9 1 11 12 0 9 13 9 15 4 0 1 9 2
9 0 9 13 16 4 0 12 9 2
22 3 12 9 11 7 9 11 0 4 2 3 15 13 2 1 15 4 1 9 4 0 2
15 1 9 9 9 11 11 11 13 4 9 9 9 9 11 2
57 1 9 1 0 9 1 11 11 11 1 9 2 12 9 2 2 11 4 13 1 0 9 0 9 0 9 11 11 1 9 9 11 15 4 13 16 11 13 0 0 9 1 11 7 4 9 12 11 0 0 9 15 4 15 13 13 2
26 11 13 3 13 9 1 9 9 1 11 15 15 2 13 9 11 0 9 9 11 2 2 13 4 11 2
7 11 1 0 9 1 9 11
24 3 1 9 9 1 16 4 15 9 11 13 1 11 2 0 9 13 4 15 13 9 11 11 2
17 3 2 0 9 13 4 1 9 3 4 9 0 9 11 13 9 2
15 9 11 11 13 1 0 9 1 9 0 0 9 1 11 2
32 0 0 0 9 13 4 15 1 9 2 12 9 2 16 4 9 11 11 13 13 0 9 1 9 11 1 11 15 13 12 9 2
22 3 1 9 4 13 0 9 3 4 9 0 9 11 2 11 2 13 9 0 9 2 2
16 11 13 4 0 9 0 9 2 3 16 4 11 13 9 9 2
46 3 2 0 0 0 9 2 3 11 2 13 4 15 1 9 16 4 0 9 13 13 1 9 2 16 15 13 1 9 0 9 1 15 15 11 13 1 9 1 15 9 1 9 1 11 2
18 15 9 1 9 4 1 0 9 1 9 1 11 2 15 4 9 9 2
27 11 4 13 16 4 13 15 9 9 16 4 13 9 9 11 1 9 3 16 15 1 9 14 13 0 9 2
27 11 11 13 15 1 3 12 9 9 15 9 1 11 2 3 15 0 9 11 11 11 13 1 9 12 9 2
41 2 1 0 12 7 12 9 13 4 16 0 9 2 1 0 0 9 2 7 13 15 16 4 15 9 4 0 1 9 2 2 13 4 1 9 9 0 9 11 11 2
29 11 11 2 9 0 0 9 2 0 9 11 2 11 2 2 13 4 16 4 16 0 9 2 11 13 9 1 9 2
39 11 4 0 9 13 1 0 9 16 4 13 9 1 15 1 15 9 2 3 0 9 0 9 7 9 2 7 0 9 1 0 11 2 9 9 1 12 9 2
11 11 3 13 16 11 13 0 0 9 11 2
11 1 9 2 9 15 3 13 13 0 9 2
24 3 1 9 2 15 0 9 2 9 9 11 11 2 13 4 16 11 14 13 3 13 1 11 2
21 13 4 16 4 13 1 9 9 16 13 9 2 3 0 11 1 9 1 0 9 2
29 9 11 1 0 3 4 4 0 9 15 4 11 13 1 9 2 7 1 15 4 13 16 11 13 1 9 0 9 2
23 3 7 1 9 11 2 9 11 3 3 4 4 1 9 13 2 3 16 13 0 0 9 2
28 9 11 11 2 9 11 2 13 4 16 4 2 3 12 9 1 0 9 2 9 1 11 1 2 0 9 2 2
9 3 4 13 16 13 9 0 9 2
37 2 16 15 13 9 1 0 9 7 9 2 15 4 13 9 0 9 3 0 9 15 0 9 2 13 16 13 13 9 12 9 2 2 13 4 9 2
19 15 9 3 13 1 0 9 11 2 1 15 4 15 9 9 9 4 0 2
6 9 13 9 0 0 9
31 9 0 9 7 9 9 11 11 11 3 15 13 2 1 9 0 9 11 11 16 15 9 7 3 12 0 9 13 9 9 2
6 0 9 11 11 11 2
16 0 0 9 11 11 13 4 9 0 9 9 3 9 0 9 2
37 9 13 16 4 9 9 7 9 2 11 2 13 2 9 2 9 15 15 13 9 2 7 16 9 13 2 0 9 2 0 1 9 11 1 0 9 2
22 9 4 13 16 15 12 9 9 2 3 9 11 11 11 2 13 9 9 1 12 9 2
28 9 11 0 4 9 0 9 1 9 1 9 1 11 7 0 9 1 9 2 15 13 9 2 9 7 0 9 2
15 16 15 9 13 2 9 12 9 4 4 0 1 9 9 2
15 12 1 12 9 13 4 0 9 11 11 11 2 0 9 2
8 11 13 15 16 0 0 9 2
12 13 4 0 9 1 0 9 3 12 9 9 2
17 0 9 2 1 9 9 2 13 4 13 9 9 0 9 1 9 2
19 1 9 1 12 9 11 4 13 16 4 9 9 0 9 15 13 0 9 2
15 3 4 13 0 0 9 1 15 15 13 9 7 0 9 2
18 15 9 2 13 4 9 2 13 0 9 11 1 9 11 1 0 9 2
20 11 4 3 13 1 9 9 16 13 9 9 1 9 7 9 1 9 0 9 2
22 3 2 3 1 9 9 2 9 1 0 9 13 4 16 4 9 4 0 1 9 9 2
11 1 9 1 9 11 4 13 15 9 9 2
19 3 4 13 9 9 2 3 16 4 9 16 15 13 9 1 9 9 0 2
7 9 1 0 9 4 0 2
30 3 1 11 2 0 9 9 2 9 11 11 13 4 16 15 9 9 11 1 3 4 0 3 13 1 15 1 0 9 2
31 3 4 9 13 11 1 9 2 13 11 2 15 4 13 16 4 13 16 4 13 0 0 9 7 13 0 9 0 9 11 2
55 2 14 4 11 11 13 9 1 15 4 13 15 9 2 13 4 15 9 1 9 1 11 7 0 9 2 7 14 4 15 13 1 15 9 2 2 13 4 9 3 16 4 11 3 0 13 13 14 1 9 4 0 9 11 2
14 0 0 9 2 11 11 1 11 2 3 15 13 9 2
25 2 0 9 13 4 13 9 1 9 9 7 13 13 9 1 9 15 15 11 13 1 9 0 9 2
8 13 4 13 9 0 9 2 2
10 11 4 1 9 13 9 1 0 9 2
32 2 1 0 0 9 0 9 13 15 1 9 7 13 1 0 9 2 7 14 1 9 2 2 13 4 9 11 1 9 11 11 2
24 2 0 9 14 13 15 13 1 9 9 2 16 15 0 9 14 4 13 13 1 0 9 2 2
12 3 0 9 0 1 0 9 1 0 9 0 9
28 9 9 0 9 0 9 11 11 0 4 1 9 3 1 9 9 1 9 2 1 15 15 13 16 13 0 9 2
25 9 13 1 9 9 7 9 0 9 1 11 1 15 4 9 3 13 12 9 1 9 2 12 9 2
28 9 1 0 9 15 4 13 1 9 13 4 1 9 3 2 12 9 2 1 0 9 0 9 2 3 0 9 2
28 1 9 4 13 3 1 12 9 3 2 3 9 1 9 9 0 9 11 11 1 0 9 3 0 9 1 11 2
28 9 13 16 15 9 13 16 4 9 0 9 9 11 11 2 0 9 2 13 13 9 15 15 13 16 9 9 2
37 2 9 4 1 0 9 15 4 13 1 9 9 9 1 15 15 4 2 3 15 13 2 13 1 9 7 13 13 2 2 13 4 0 9 11 11 2
14 2 13 4 0 9 2 4 4 3 9 7 9 2 2
14 9 9 3 4 0 2 7 9 4 13 9 1 9 2
14 11 2 15 4 0 2 13 16 4 9 4 0 15 2
23 3 0 7 0 9 11 2 13 4 16 4 15 15 15 13 1 9 4 0 1 9 9 2
25 2 13 4 9 2 0 9 7 9 9 9 2 2 13 4 11 9 1 15 9 3 9 1 9 2
37 2 15 4 0 9 4 0 1 9 9 2 2 13 4 2 3 16 15 9 4 13 9 1 9 2 16 13 9 15 9 2 15 9 7 9 2 2
6 3 15 4 13 9 2
41 1 9 0 1 11 2 0 9 1 9 11 11 13 4 1 0 9 2 0 0 9 1 9 2 15 15 13 1 9 0 9 11 7 11 2 16 0 9 0 9 2
14 9 4 3 15 9 13 9 7 3 12 9 15 9 2
16 11 13 16 4 9 9 0 1 9 4 9 16 9 4 0 2
34 3 15 16 2 0 9 2 2 9 11 11 13 4 15 9 0 9 2 3 16 15 9 4 13 0 9 16 13 15 9 7 13 11 2
37 2 1 9 3 15 9 7 15 9 3 13 16 13 9 1 9 2 0 9 13 13 9 9 7 15 9 2 2 13 4 1 9 0 3 1 9 2
17 9 13 0 9 16 4 13 4 14 9 0 1 9 3 7 9 2
6 9 9 2 9 11 2
17 1 9 15 9 9 9 2 11 4 13 15 9 1 0 0 9 2
14 3 2 1 9 9 1 0 9 2 0 4 9 0 2
10 11 8 12 4 9 4 9 0 9 2
25 11 4 13 0 9 1 11 2 3 1 9 16 4 9 11 11 1 9 1 9 1 0 9 12 2
42 3 2 9 4 13 13 9 0 9 12 2 12 1 9 11 1 15 0 9 1 9 2 15 4 9 1 0 9 13 0 9 2 1 9 16 4 1 0 9 13 11 2
30 9 1 11 13 4 9 12 9 2 3 16 4 9 11 11 13 15 3 0 9 1 9 2 15 4 13 0 12 9 2
22 11 4 13 16 15 4 13 1 11 1 9 2 16 4 13 13 15 9 0 9 9 2
27 9 4 13 4 14 15 9 4 3 0 9 7 4 2 9 11 2 2 3 15 0 9 3 13 2 0 2
12 0 0 9 11 11 13 15 0 9 0 11 2
41 11 2 12 2 4 4 9 12 0 9 1 11 2 11 11 2 11 11 7 11 11 2 1 15 4 13 7 1 9 0 2 0 9 2 2 11 2 11 7 11 2
27 13 14 15 9 0 2 13 15 16 4 13 2 9 2 9 1 15 4 0 9 1 0 7 0 0 9 2
30 1 9 2 0 9 15 4 13 0 9 1 0 9 4 4 0 1 9 2 16 7 1 9 11 11 1 0 9 11 2
20 9 0 9 3 4 0 1 9 1 9 2 7 9 4 1 0 9 4 0 2
20 12 1 0 9 0 9 2 0 9 1 9 9 2 13 4 15 9 1 9 2
36 15 15 13 0 9 2 0 2 0 2 9 1 0 0 9 1 9 15 9 13 4 15 0 2 3 16 15 1 0 9 4 13 7 0 9 2
22 1 9 1 15 2 9 4 1 0 9 11 13 4 0 1 9 15 4 13 1 9 2
51 3 16 15 4 9 11 11 1 12 9 13 0 9 1 0 9 2 2 0 2 11 4 3 13 13 0 9 1 9 11 11 11 11 2 15 4 0 9 1 0 9 12 13 13 7 9 15 3 0 9 2
13 0 4 9 13 1 0 9 1 0 9 7 9 2
45 13 15 16 4 9 4 0 9 1 0 7 0 9 2 1 15 4 0 4 0 9 9 15 4 13 1 0 0 9 2 16 7 9 7 9 2 15 4 11 13 1 0 11 11 2
24 1 0 2 9 4 4 3 0 2 7 15 15 1 9 7 9 4 13 13 1 9 1 9 2
5 9 2 9 11 2
22 4 14 13 9 16 15 11 13 15 9 1 0 11 16 0 9 1 9 1 0 9 2
9 11 11 13 15 4 9 1 15 2
31 1 0 9 2 0 9 2 0 9 7 0 9 2 11 13 3 1 13 9 2 16 15 9 16 9 1 9 13 3 0 2
13 11 15 13 13 0 9 7 9 0 9 0 9 2
19 9 14 13 4 0 2 16 4 11 0 0 9 9 16 4 13 15 9 2
25 4 14 9 0 2 13 9 16 4 0 9 1 0 0 9 13 13 1 9 0 9 0 0 9 2
10 9 9 1 11 13 4 13 1 9 9
20 0 8 9 9 2 15 15 13 13 3 15 9 2 0 4 1 9 0 9 2
14 9 13 9 0 9 1 9 2 12 9 2 1 11 2
20 0 9 13 9 0 9 15 13 0 2 13 4 9 1 9 2 12 9 2 2
18 9 4 4 9 0 9 15 4 13 1 9 0 8 9 9 1 11 2
27 9 9 9 11 11 13 4 1 11 16 9 13 13 1 0 9 1 11 2 9 0 9 15 13 9 2 2
14 0 9 9 7 0 0 9 12 13 4 15 8 9 2
27 9 9 11 11 13 4 16 4 9 4 0 1 15 15 4 15 13 13 16 15 9 13 16 15 4 0 2
28 1 9 0 9 2 9 1 3 12 9 13 4 13 9 9 9 0 1 0 9 1 9 15 15 9 13 13 2
19 9 4 3 13 9 1 9 11 2 15 4 13 4 9 9 1 9 9 2
24 0 9 15 0 9 3 4 15 13 13 1 9 9 2 15 4 15 13 16 3 3 13 9 2
40 9 0 9 13 4 16 9 14 13 13 9 9 9 7 13 9 9 1 9 9 1 9 9 2 1 9 9 11 7 11 2 3 4 9 9 13 4 3 0 2
20 2 9 0 9 0 4 13 9 1 0 9 3 4 1 9 9 7 0 9 2
30 13 4 9 9 15 4 9 13 13 2 16 14 4 4 0 7 1 12 0 9 2 2 13 4 9 0 9 11 11 2
5 9 4 15 13 2
33 2 9 1 0 0 0 9 4 16 15 15 9 13 1 0 9 2 16 4 15 13 16 4 9 8 7 0 9 9 0 9 9 2
26 14 13 13 1 15 9 1 9 9 2 15 14 4 4 9 9 2 2 13 4 9 0 9 11 11 2
19 9 9 9 13 4 16 4 2 9 13 1 9 9 2 2 13 4 9 2
42 9 0 9 11 11 13 4 1 9 16 4 4 0 2 0 8 2 1 9 15 13 9 2 3 16 4 1 9 0 12 9 1 15 4 13 13 0 9 1 9 11 2
21 9 4 3 13 16 2 3 2 15 0 9 4 4 0 1 9 11 1 0 9 2
6 13 15 9 9 1 11
22 3 9 9 1 9 9 2 0 9 11 11 13 15 1 9 1 9 7 9 0 9 2
21 0 9 11 11 2 1 9 2 13 9 9 1 11 2 1 9 2 12 9 2 2
5 13 4 13 9 2
31 1 11 4 1 9 2 12 9 2 13 7 0 9 9 1 9 7 9 1 0 9 9 15 4 11 13 1 9 9 12 2
42 9 4 13 1 15 4 0 9 1 9 1 9 13 9 9 1 15 9 9 0 9 13 16 11 13 9 1 9 1 9 9 1 9 3 4 13 9 1 0 0 9 2
14 2 3 4 15 13 2 2 13 15 9 11 1 9 2
11 2 7 12 9 1 11 4 4 3 0 2
11 3 4 13 0 9 7 3 2 12 9 2
19 1 0 12 9 4 15 13 2 1 15 2 13 4 1 9 1 9 2 2
18 3 12 9 13 15 1 9 1 0 9 1 9 2 3 1 0 9 2
20 9 4 13 0 3 15 9 1 15 4 9 9 13 7 13 9 9 0 9 2
10 1 11 2 0 4 3 1 12 9 2
16 3 4 3 1 9 13 0 9 1 9 7 9 1 9 11 2
11 0 4 3 12 9 16 15 4 12 0 2
11 9 4 1 9 9 13 9 7 0 9 2
23 1 9 2 0 12 0 9 0 1 9 2 3 0 0 9 0 9 11 2 13 4 9 2
19 3 2 9 11 11 11 13 4 9 1 9 3 15 15 9 1 0 9 2
30 0 9 1 11 13 15 13 1 3 1 12 9 2 13 4 2 7 0 9 13 4 9 1 0 0 9 15 13 11 2
40 2 16 9 9 12 9 13 16 4 0 9 13 9 2 9 13 13 7 1 15 13 9 9 2 2 13 4 11 1 0 9 1 9 2 7 13 0 9 8 2
18 2 9 4 0 2 16 1 15 4 0 9 2 9 7 9 9 2 2
37 11 4 2 1 9 2 3 13 16 14 13 13 1 9 9 7 13 9 2 3 15 16 4 1 15 13 1 0 2 16 0 2 9 9 0 9 2
43 1 0 9 0 9 2 13 15 16 4 15 9 0 9 11 13 12 2 11 2 15 4 0 9 1 11 7 3 1 0 9 1 12 2 1 9 15 15 13 13 1 9 2
16 1 9 16 13 0 0 9 2 11 4 13 9 7 13 9 2
19 0 0 9 13 4 13 9 2 16 7 0 9 1 0 9 7 0 9 2
10 11 2 11 7 11 11 13 13 1 11
32 9 0 9 11 7 11 11 11 11 13 4 16 15 9 13 1 9 13 1 9 11 1 0 9 3 4 15 13 11 7 11 2
43 11 7 11 11 4 4 0 1 11 7 11 16 1 9 14 13 1 0 0 9 1 0 11 2 11 2 2 13 4 1 9 2 12 9 2 9 0 9 15 9 11 11 2
17 1 9 11 2 11 4 0 9 13 16 12 1 0 9 15 9 2
17 2 13 12 3 0 9 15 13 13 16 15 13 13 11 7 11 2
12 13 1 9 1 0 9 2 2 13 4 11 2
22 1 15 9 2 1 9 9 15 9 9 4 13 2 3 9 0 9 1 9 1 11 2
28 11 4 3 0 1 9 0 9 15 15 13 1 9 7 13 11 9 1 0 9 0 1 9 1 11 0 9 2
51 0 0 9 11 11 7 15 15 9 3 4 1 0 9 2 16 11 4 13 9 1 9 0 0 9 1 11 2 3 9 0 0 9 1 15 4 0 9 0 9 1 15 9 1 9 1 11 12 2 12 2
19 9 0 11 1 9 9 11 11 7 11 9 3 15 3 3 13 1 9 2
30 3 16 0 9 15 13 11 13 3 4 0 1 11 2 11 4 13 16 4 15 13 9 15 9 2 7 14 13 9 2
21 2 13 9 1 15 9 2 2 13 4 11 1 9 9 1 11 2 7 13 11 2
18 2 15 0 0 9 13 4 9 15 9 0 9 1 11 7 0 9 2
22 11 7 11 11 4 9 1 11 7 11 4 9 1 11 7 11 11 2 2 13 4 2
22 1 9 2 0 9 9 11 11 13 4 16 4 9 9 11 1 11 13 4 0 9 2
55 2 13 9 9 2 11 2 11 2 13 9 2 11 2 11 2 15 1 11 11 3 4 1 9 2 7 0 3 13 13 1 0 9 2 2 13 4 11 1 9 1 9 11 2 9 1 9 11 2 7 13 0 9 11 2
38 9 11 1 11 7 11 11 11 11 1 9 4 13 9 9 1 15 15 13 0 9 9 11 7 11 1 15 4 15 13 9 9 0 9 1 0 9 2
24 3 1 9 9 11 1 0 9 2 2 3 2 4 3 13 1 15 9 2 13 4 11 11 2
36 2 9 15 3 3 13 1 9 15 9 13 9 2 7 3 3 3 2 13 0 9 16 4 9 0 9 1 15 15 13 13 2 2 13 4 2
10 9 7 9 2 0 0 0 13 0 9
17 0 7 0 9 1 0 11 4 4 0 1 11 2 11 7 11 2
19 3 1 9 9 1 9 7 9 2 11 11 11 13 4 0 9 0 9 2
24 0 0 0 0 1 11 13 4 12 9 1 9 7 9 2 0 9 1 11 2 11 7 11 2
35 1 9 9 9 9 11 11 2 9 4 13 3 12 0 7 0 0 9 1 9 11 2 11 2 11 7 11 2 16 7 9 0 0 9 2
22 12 1 0 0 9 2 11 11 11 2 13 4 1 9 0 9 0 9 12 2 12 2
24 12 0 9 9 9 0 9 7 0 0 9 13 4 16 15 0 9 1 9 1 9 7 9 2
15 0 0 9 2 11 11 2 13 4 9 1 0 9 11 2
44 9 12 9 1 9 12 1 0 0 9 2 9 0 9 2 11 11 2 0 4 1 9 2 12 9 2 1 15 0 9 11 1 11 7 11 0 9 7 0 9 9 15 9 2
6 9 4 13 9 11 2
25 0 9 11 11 2 13 4 2 3 15 13 2 15 9 1 11 1 9 0 9 2 8 8 2 2
21 11 4 13 0 0 9 1 9 2 1 15 4 1 15 13 7 0 9 11 11 2
17 9 15 15 13 0 0 9 0 4 1 0 9 11 11 1 11 2
33 1 9 1 9 2 9 12 9 2 2 0 4 9 2 9 2 9 2 9 7 9 15 13 1 0 9 2 3 0 9 12 9 2
17 9 4 1 11 4 0 1 12 9 2 7 3 15 13 1 11 2
18 9 9 0 0 9 11 11 0 4 1 9 11 11 1 11 1 11 2
12 9 11 0 9 2 0 4 1 9 0 9 2
5 0 9 1 0 9
12 12 4 0 9 0 9 15 9 13 0 9 2
42 9 9 11 11 1 0 0 9 2 11 2 13 4 12 9 9 1 9 9 11 11 1 9 9 1 15 15 4 11 13 13 15 9 1 11 16 13 9 1 0 9 2
37 2 15 4 9 0 9 15 4 13 1 0 0 9 7 15 4 13 3 16 7 15 2 2 13 4 11 1 15 4 4 0 13 9 1 12 9 2
20 11 4 13 16 4 15 9 4 9 1 15 15 13 9 1 0 9 1 9 2
22 13 4 7 16 9 11 11 11 2 15 15 13 1 9 1 11 2 4 13 15 9 2
13 16 4 11 13 9 9 2 0 4 1 12 9 2
27 9 9 0 9 11 11 13 4 9 11 2 3 16 4 4 2 0 1 0 9 1 15 4 13 9 2 2
28 11 15 4 13 1 0 9 15 4 9 13 0 9 11 11 11 2 3 2 2 15 4 9 13 1 9 2 2
26 0 0 9 13 4 9 1 9 7 13 15 9 2 3 16 4 1 15 9 9 13 1 0 9 9 2
40 11 4 9 2 3 7 0 9 3 2 13 15 9 7 13 15 16 2 9 2 2 16 4 0 2 1 11 2 13 16 4 9 4 0 7 13 8 12 9 2
35 9 0 9 0 0 9 11 2 11 2 11 11 13 4 16 4 9 11 4 0 1 15 15 15 13 2 0 9 9 9 2 1 9 9 2
35 13 4 16 2 16 15 3 13 9 3 15 9 2 3 9 2 3 3 9 2 7 2 3 9 2 3 4 15 15 15 4 1 9 2 2
12 3 2 9 0 9 4 13 9 1 15 9 2
19 13 4 16 4 9 4 0 1 9 0 0 9 7 13 9 9 9 11 2
27 11 11 2 9 0 9 0 9 1 0 11 2 13 4 16 4 11 9 9 2 3 3 13 2 0 9 2
16 2 13 3 0 0 9 7 15 13 1 0 2 2 13 4 2
27 2 9 9 16 9 13 1 9 1 15 9 13 4 16 15 4 13 7 15 9 1 3 2 2 13 4 2
9 0 9 0 9 1 11 0 9 9
19 0 9 2 15 4 15 9 13 1 0 9 2 13 4 15 9 1 9 2
5 0 9 1 11 2
27 0 9 0 9 11 11 7 9 11 11 2 0 9 0 9 2 1 9 4 15 13 1 0 9 0 9 2
15 9 4 0 9 13 0 2 7 0 4 9 13 0 9 2
17 9 15 3 13 11 3 13 9 1 9 12 13 4 9 1 9 2
33 9 13 9 15 15 13 1 9 1 15 4 13 9 1 9 11 9 9 1 0 9 1 12 9 2 3 13 9 15 4 13 9 2
21 13 15 15 9 2 7 13 15 16 11 1 0 9 9 9 3 13 9 1 9 2
18 9 4 1 0 9 1 0 9 13 9 9 16 4 15 13 15 9 2
15 9 4 13 9 1 15 15 13 16 4 15 9 13 9 2
32 2 0 9 13 9 0 9 2 4 9 1 0 9 7 1 0 9 0 9 2 2 13 4 11 2 3 9 0 1 12 9 2
29 11 4 13 9 1 9 15 4 0 13 9 0 9 2 16 7 11 11 2 0 9 15 4 13 16 4 13 9 2
45 3 1 1 15 0 9 0 0 9 7 9 11 11 2 0 4 9 11 11 2 15 15 1 3 4 13 1 0 9 2 13 0 9 1 15 4 13 9 16 15 4 15 9 13 2
24 2 3 13 15 11 1 15 15 4 1 15 0 15 15 9 7 9 15 1 15 13 13 2 2
40 9 8 8 2 11 2 2 0 0 0 9 1 9 9 15 4 2 1 0 2 13 9 1 11 2 13 4 2 9 9 7 9 15 13 0 9 1 9 2 2
36 2 1 15 9 2 11 0 9 13 1 9 7 9 9 0 9 2 15 16 16 4 13 16 9 14 13 3 9 2 2 0 4 1 0 9 2
9 2 0 0 9 13 4 0 9 2
26 0 4 0 9 9 0 9 15 9 2 2 13 4 1 11 11 11 2 9 9 1 0 9 11 11 2
36 2 15 0 9 0 4 1 9 0 9 0 9 2 9 0 9 7 9 1 15 9 15 15 4 3 4 0 15 2 9 2 2 2 13 4 2
20 1 9 11 0 1 9 2 11 13 12 2 9 2 16 15 11 13 12 2 2
8 0 9 2 9 9 13 1 9
22 11 2 11 2 11 7 11 11 13 1 9 9 2 16 11 7 11 13 9 15 9 2
41 9 11 11 11 2 3 2 2 9 11 11 11 11 2 0 1 3 2 2 0 9 11 11 11 2 0 1 3 2 7 9 11 11 11 13 15 1 9 1 11 2
44 0 9 11 7 11 11 11 7 9 11 2 11 7 11 11 2 11 11 2 11 11 7 11 11 2 2 13 4 15 1 11 1 9 2 12 9 2 1 9 1 9 1 11 2
17 1 9 15 4 0 1 9 9 13 15 1 0 9 7 0 9 2
28 9 11 11 11 11 13 4 1 9 2 12 9 2 1 11 11 16 15 9 13 9 7 0 9 11 7 11 2
25 1 9 1 9 9 0 2 11 2 11 11 2 11 4 3 13 9 9 11 1 9 11 7 11 2
22 13 4 16 4 12 0 0 9 13 13 9 16 13 9 0 2 1 9 9 15 9 2
18 3 4 13 9 16 4 12 9 13 9 1 0 9 15 4 3 3 2
35 11 7 11 13 1 9 13 0 0 9 2 13 4 1 9 2 12 9 2 9 9 7 9 11 11 1 9 1 0 9 11 11 1 11 2
27 2 1 9 1 15 9 2 13 9 3 13 13 2 3 1 9 2 2 13 4 11 2 3 0 9 11 2
41 9 9 12 9 1 2 0 9 2 2 3 11 2 11 7 11 2 11 2 11 7 11 2 0 4 1 9 2 12 9 2 1 0 9 11 1 15 4 11 9 2
16 9 4 13 0 9 3 1 0 9 9 1 9 7 0 9 2
14 9 4 3 13 9 1 0 9 1 9 7 0 9 2
28 0 9 11 11 13 4 1 0 9 11 1 9 2 12 9 2 15 0 9 9 11 1 9 1 11 7 11 2
24 1 0 0 9 1 0 9 11 11 2 11 4 13 16 11 13 9 1 9 1 9 1 11 2
31 0 9 11 11 7 15 0 9 11 11 13 4 15 1 9 2 12 9 2 16 4 0 9 0 2 7 16 0 9 13 2
29 11 4 13 9 11 9 11 1 9 1 11 2 3 16 11 13 16 0 9 1 9 13 15 9 9 1 11 3 2
29 0 9 11 11 11 13 4 1 9 2 12 9 2 0 0 9 1 11 2 3 0 9 12 9 1 0 9 11 2
34 1 9 1 0 9 1 11 11 2 11 4 13 16 4 11 7 11 2 12 0 9 9 9 11 2 13 9 13 9 0 9 0 9 2
9 9 7 9 2 8 11 13 11 11
17 9 1 9 13 4 11 11 7 8 11 1 9 3 1 11 11 2
24 3 15 9 2 1 11 0 0 9 2 7 11 11 11 13 9 9 1 9 0 9 1 11 2
32 11 11 2 3 2 13 1 9 11 11 1 9 0 9 11 1 11 11 1 9 2 12 9 2 1 9 9 8 11 8 8 2
32 3 12 9 1 11 11 2 11 2 11 7 11 7 11 13 4 1 9 2 12 9 2 9 8 11 1 9 11 1 9 11 2
17 9 9 2 15 4 0 1 9 9 8 8 2 13 4 12 9 2
19 1 0 4 4 0 9 11 11 2 9 11 11 11 7 0 9 11 11 2
24 11 4 13 0 9 1 0 0 9 1 12 11 2 0 0 9 15 4 0 0 9 1 11 2
20 11 9 4 4 0 1 3 12 9 2 1 11 1 12 7 11 1 12 9 2
18 1 3 12 0 9 1 11 2 11 11 7 11 11 13 4 1 12 2
17 0 0 0 9 0 4 1 9 2 12 9 2 1 11 1 11 2
31 9 1 12 9 13 4 15 1 9 9 7 9 2 9 2 9 2 9 2 9 2 8 8 8 2 9 2 9 7 9 2
24 11 4 3 0 16 0 9 9 2 1 9 1 11 11 1 0 9 11 1 0 9 1 9 2
21 0 0 9 11 0 4 1 9 2 12 9 2 1 9 9 1 9 11 1 11 2
14 9 4 13 3 12 9 0 9 11 1 11 7 11 2
17 1 11 1 11 1 12 9 1 12 9 0 4 0 9 0 9 2
40 3 12 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 7 11 13 4 1 9 2 15 4 3 13 9 1 0 9 7 0 9 11 2
21 0 9 11 11 3 4 1 9 2 12 9 2 0 1 0 0 9 2 11 2 2
28 9 11 11 1 9 3 4 0 1 12 9 0 9 11 1 11 11 2 1 15 4 11 11 13 9 0 9 2
5 11 13 0 9 11
19 0 9 11 11 13 4 9 1 12 9 1 15 4 4 0 0 9 11 2
13 13 14 15 11 13 1 9 16 13 0 9 11 2
15 1 9 2 12 9 2 0 4 9 0 1 0 9 11 2
16 12 9 15 13 0 9 9 0 4 1 9 9 0 12 9 2
15 9 7 9 4 4 0 9 9 2 15 4 13 12 9 2
19 2 9 4 1 9 1 0 0 9 2 2 13 4 0 9 9 11 11 2
22 13 4 9 3 1 9 0 9 2 11 11 2 12 9 1 9 9 11 7 0 9 2
22 13 15 16 4 9 0 9 9 4 0 1 0 12 1 12 9 2 3 1 0 9 2
11 9 2 9 7 9 13 15 1 15 9 2
9 9 15 13 1 0 9 7 9 2
11 0 9 4 4 0 1 9 0 9 9 2
14 12 15 9 13 1 9 12 9 2 0 9 12 9 2
14 9 15 13 1 3 0 9 1 9 7 9 0 9 2
8 15 9 13 15 1 12 9 2
10 9 15 13 1 9 0 9 11 11 2
19 9 1 9 0 9 2 15 4 13 9 1 12 2 13 4 1 3 9 2
27 0 9 9 11 11 4 12 13 0 9 1 9 0 9 2 16 9 15 4 3 0 3 4 13 1 9 2
8 0 4 9 0 1 9 12 2
14 11 11 2 0 0 9 2 4 4 12 1 9 9 2
18 13 4 9 11 11 2 9 0 1 11 2 15 3 13 1 8 11 2
16 0 4 9 0 1 9 11 7 1 15 13 9 1 0 9 2
15 9 4 1 0 0 9 1 12 0 9 2 0 1 9 2
19 3 12 9 9 9 7 9 9 2 15 3 13 12 9 9 2 13 11 2
18 3 4 9 13 3 12 9 9 2 16 9 4 0 1 12 9 9 2
19 9 9 2 15 13 1 0 9 11 2 13 9 1 0 9 7 0 9 2
17 0 9 2 0 0 9 2 13 0 9 1 0 9 1 0 9 2
15 13 7 0 9 2 9 1 9 7 9 1 9 1 11 2
10 3 2 1 0 15 9 13 9 11 2
14 0 4 9 4 0 1 0 9 7 0 9 0 9 2
17 9 9 13 9 0 9 1 11 1 0 9 0 9 2 0 11 2
21 9 1 9 9 4 11 1 0 9 2 7 9 13 9 16 15 3 13 1 9 2
20 0 4 9 0 0 9 15 4 0 3 3 11 2 7 9 4 13 1 9 2
11 9 13 16 4 9 3 0 1 15 9 2
24 2 15 4 9 13 16 4 9 0 9 9 11 2 16 15 14 13 9 11 2 2 13 11 2
23 2 13 15 15 9 9 1 15 9 7 16 9 0 12 9 1 15 9 13 15 9 2 2
10 0 4 9 4 1 9 1 9 12 2
21 9 11 13 4 15 0 2 9 12 2 1 15 4 15 3 13 0 9 7 9 2
23 0 15 11 13 16 4 15 0 9 13 1 9 0 0 9 15 4 3 0 1 0 9 2
16 9 0 9 4 4 9 1 15 4 13 9 1 9 15 9 2
10 11 15 3 13 9 0 9 1 11 2
23 2 0 4 3 0 0 9 11 2 2 13 4 11 11 2 0 0 9 1 9 0 9 2
17 2 15 4 0 9 1 11 7 0 9 1 9 0 0 9 2 2
34 9 15 13 2 0 7 1 9 0 9 2 3 4 13 11 7 0 9 11 2 13 3 1 9 15 15 4 13 1 0 9 15 9 2
20 0 4 9 12 9 2 16 15 4 9 1 9 13 0 9 1 9 0 9 2
33 13 12 9 0 9 2 1 0 12 9 2 2 12 9 2 1 0 12 2 0 1 0 9 11 7 12 9 1 0 7 0 9 2
31 1 15 2 9 13 9 1 11 2 1 0 12 2 2 12 9 9 0 9 7 0 9 11 2 11 2 11 7 0 9 2
23 1 0 4 9 9 1 15 4 15 13 13 3 9 4 0 0 2 16 14 0 0 9 2
26 2 9 9 13 4 0 9 1 9 15 9 2 2 13 9 11 11 2 9 9 1 9 0 9 11 2
8 9 7 9 2 11 13 0 9
12 0 9 11 11 0 4 9 1 9 9 11 2
18 1 0 9 1 9 2 0 9 13 4 1 9 0 9 15 13 11 2
3 11 11 2
24 0 9 11 11 13 4 1 9 2 12 9 2 9 1 0 9 1 9 0 9 1 9 11 2
10 9 4 13 1 9 2 0 9 2 2
18 9 15 13 0 9 2 7 13 9 2 9 2 9 2 9 7 9 2
25 0 0 9 9 0 4 1 9 0 0 9 1 9 9 2 13 4 0 9 1 9 2 12 9 2
19 9 4 0 1 0 9 1 9 9 9 9 2 15 4 9 1 11 2 2
19 0 9 11 11 1 0 11 13 15 1 9 9 1 0 9 15 13 11 2
16 11 4 12 1 12 9 7 12 1 1 12 9 1 12 9 2
20 9 9 4 4 0 1 0 9 11 12 9 2 15 4 9 4 0 1 9 2
27 0 0 0 9 11 9 12 13 4 1 9 2 12 9 2 1 11 11 2 1 11 7 11 2 11 2 2
36 9 13 1 9 2 12 9 2 16 13 4 12 0 0 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
33 1 11 4 15 3 13 0 9 15 4 15 4 0 1 0 9 2 13 4 1 9 2 12 9 2 0 9 9 7 9 11 11 2
16 9 1 9 0 9 9 4 4 0 1 9 2 13 4 9 2
23 0 4 9 9 9 9 0 1 9 9 7 9 9 1 12 9 0 9 1 12 7 12 2
25 11 9 11 11 13 4 1 9 2 12 9 2 0 11 9 1 11 2 11 2 13 4 0 9 2
16 1 9 4 0 11 13 11 11 11 1 12 2 12 2 12 2
20 11 4 9 1 9 13 12 9 2 7 4 3 1 12 9 9 0 9 9 2
27 11 11 2 1 11 7 11 2 4 4 9 0 9 0 9 2 11 2 1 9 2 12 9 2 1 9 2
28 9 4 13 9 12 0 2 0 2 0 7 0 9 2 16 9 4 4 1 9 11 2 15 13 9 1 9 2
8 9 0 9 0 9 0 9 11
24 9 9 11 4 4 0 9 1 0 9 15 0 9 1 12 9 2 13 4 0 9 0 9 2
25 3 9 9 2 11 4 13 16 4 9 9 11 4 0 9 1 15 9 15 0 9 1 12 9 2
23 3 0 9 9 4 4 9 1 9 9 2 16 7 9 1 9 1 9 2 9 7 9 2
17 9 9 7 9 9 1 0 0 9 3 15 13 1 9 0 9 2
48 2 0 9 1 11 13 4 0 9 0 9 15 4 13 1 9 15 13 2 2 13 4 1 9 2 12 9 2 1 11 0 9 0 9 11 11 3 1 9 9 0 9 9 9 11 1 9 2
29 2 9 15 9 13 0 3 7 15 4 4 0 9 15 9 1 12 9 2 2 13 4 0 9 2 11 2 11 2
33 0 9 11 7 11 2 13 4 11 2 2 13 4 0 9 1 9 9 7 9 7 9 9 0 9 11 2 2 1 11 1 11 2
42 11 4 2 13 4 15 2 0 9 13 9 1 9 9 9 9 7 9 1 12 9 15 4 0 1 9 1 11 2 16 7 0 0 9 11 1 9 7 9 1 9 2
15 11 4 13 1 2 0 0 9 2 1 9 1 0 9 2
21 3 9 0 9 1 9 9 11 2 11 15 9 13 9 9 1 9 7 9 9 2
41 11 4 13 16 4 15 9 2 2 15 4 4 0 1 0 9 9 7 9 2 9 9 7 0 7 0 9 2 2 13 4 0 1 0 9 15 4 13 7 11 2
14 11 4 3 13 1 3 12 9 15 15 13 15 9 2
25 15 4 4 0 9 2 9 9 7 9 1 9 7 9 7 9 1 0 9 9 7 9 1 9 2
28 11 4 13 9 0 7 0 9 1 11 7 11 2 11 2 11 2 9 11 7 0 0 9 2 13 4 11 2
33 13 4 16 4 9 4 4 3 12 1 15 9 16 11 2 3 9 9 1 9 0 9 2 9 9 7 9 9 1 0 0 9 2
29 3 9 1 15 4 0 0 0 9 1 11 2 11 4 13 9 9 11 15 9 1 9 0 9 7 9 0 9 2
24 3 4 13 16 4 2 1 9 9 0 1 12 9 2 13 1 9 0 7 0 9 0 9 2
30 16 11 2 9 0 9 9 9 11 15 4 0 1 9 0 0 9 9 2 0 4 1 0 0 9 7 9 9 11 2
21 15 16 11 13 0 0 9 1 15 4 15 9 9 0 9 11 2 11 7 11 2
33 11 4 9 9 11 0 9 13 1 11 2 16 11 4 1 9 11 13 0 0 9 0 9 11 8 11 11 2 0 0 9 11 2
16 0 9 0 9 0 9 12 9 13 4 11 1 9 11 11 2
8 1 11 13 0 2 0 0 9
14 11 7 11 13 3 0 9 16 15 13 9 0 9 2
11 9 13 1 0 9 0 0 9 1 11 2
13 9 1 0 9 12 9 0 4 2 13 0 9 2
37 9 11 13 16 0 9 0 9 2 11 0 9 2 11 2 2 7 15 0 9 1 9 2 0 9 2 11 2 2 13 15 1 12 9 9 9 2
27 9 4 3 13 1 9 2 12 9 2 2 3 3 4 13 0 9 1 0 9 1 9 9 0 0 9 2
19 1 0 12 9 9 4 13 11 2 13 9 7 13 9 1 9 1 9 2
25 3 16 4 9 3 0 2 9 13 1 9 9 11 2 11 2 7 0 2 0 2 0 2 9 2
9 15 4 4 0 15 9 1 11 2
22 9 11 11 0 4 13 15 9 2 3 16 4 1 0 9 9 13 4 3 13 9 2
12 16 7 13 0 9 2 3 13 3 9 15 2
14 12 9 13 4 9 2 16 9 4 1 3 4 0 2
21 11 4 2 3 2 13 9 0 1 0 2 15 13 11 2 7 0 2 11 2 2
22 1 0 9 13 15 9 11 2 16 15 1 0 13 3 0 9 11 1 9 0 9 2
20 11 15 1 9 13 13 1 15 2 3 15 1 0 9 1 1 9 1 11 2
24 3 2 9 4 13 9 16 4 9 11 11 11 3 13 15 9 11 1 9 1 9 1 11 2
16 2 3 15 15 4 13 2 7 7 11 2 2 13 4 11 2
25 3 2 9 9 9 9 1 9 9 11 11 4 4 0 11 2 15 4 4 9 9 1 0 9 2
7 11 4 3 13 15 9 2
26 7 12 9 4 13 3 4 9 13 1 9 7 9 0 9 2 7 4 13 16 4 15 13 1 9 2
13 1 0 0 9 2 1 11 4 0 3 12 9 2
19 0 9 9 13 15 1 12 7 12 9 2 16 3 12 9 9 4 9 2
14 11 13 12 0 9 2 1 15 15 13 12 9 11 2
11 9 13 12 0 9 2 16 0 9 12 2
16 16 4 4 0 1 11 2 0 9 13 13 1 12 9 9 2
7 9 3 1 9 9 1 11
19 0 9 11 3 4 13 7 13 9 2 15 4 3 4 1 9 0 9 2
22 3 1 12 9 1 11 13 4 1 9 2 12 9 2 0 9 12 9 0 0 9 2
17 9 13 9 9 7 9 9 2 1 15 4 3 4 0 9 9 2
14 15 9 3 4 4 0 13 9 9 7 13 15 9 2
12 1 15 9 0 4 0 9 0 9 1 11 2
16 9 9 13 4 9 9 0 9 2 2 11 11 7 11 11 2
52 3 4 0 11 11 2 0 9 11 12 2 2 11 11 2 9 1 11 2 7 11 11 2 9 1 11 2 2 9 9 9 0 9 2 2 0 11 2 9 11 2 2 11 11 7 11 11 2 9 11 2 2
19 2 3 15 13 9 0 0 9 1 11 2 2 13 4 9 9 11 11 2
19 2 13 15 16 4 9 2 15 0 9 13 9 9 2 13 0 9 2 2
12 13 4 16 15 9 1 9 9 13 9 9 2
37 2 9 0 1 0 9 13 0 9 2 16 4 9 9 15 13 13 7 13 9 7 9 0 9 2 2 13 4 11 11 2 9 9 0 1 9 2
14 13 4 16 4 9 1 9 9 0 1 9 16 9 2
23 9 0 9 9 4 4 0 1 9 1 0 9 2 16 9 9 15 13 9 13 4 9 2
18 9 9 7 9 0 9 3 4 9 9 2 15 4 3 13 12 9 2
12 15 0 9 13 0 9 1 9 1 0 9 2
19 9 0 9 1 3 4 13 9 2 7 15 13 16 4 15 9 3 0 2
4 11 13 0 9
29 0 9 1 11 0 4 9 15 4 13 9 1 11 2 2 15 4 9 15 4 1 9 11 13 0 9 1 9 2
19 0 9 13 4 0 9 16 4 13 9 12 9 1 11 2 1 9 9 2
24 0 9 13 16 4 13 9 1 15 9 2 7 15 4 0 9 9 7 15 13 1 0 9 2
11 1 9 9 9 2 9 4 13 15 9 2
28 1 0 9 1 9 2 12 9 2 2 9 0 9 13 4 16 4 15 9 0 9 15 4 13 9 1 11 2
23 1 9 9 9 0 9 11 11 2 1 11 4 13 1 9 7 13 9 1 9 1 9 2
10 1 9 4 13 1 0 9 7 9 2
19 9 9 1 11 13 4 0 1 0 7 0 9 7 13 4 0 1 9 2
9 1 12 9 13 4 13 0 9 2
28 11 13 4 11 1 15 9 7 13 9 16 4 15 9 13 0 9 1 9 1 11 1 9 16 13 0 9 2
47 2 1 0 9 12 9 1 3 2 11 4 13 0 9 1 9 0 9 9 2 1 9 1 9 1 9 1 12 9 7 0 9 7 9 2 2 13 4 9 11 1 11 11 2 11 11 2
17 9 9 9 12 4 1 9 15 15 13 13 1 9 1 9 11 2
23 1 12 9 2 3 4 0 0 9 1 9 2 12 9 13 4 9 2 16 4 0 0 2
28 1 12 9 0 0 9 2 3 15 4 13 1 11 2 0 0 9 11 7 11 11 2 11 2 11 7 11 2
16 9 9 2 0 9 13 4 16 4 9 13 12 0 0 9 2
25 1 9 9 11 8 11 2 9 0 9 1 9 11 11 2 11 11 2 13 4 13 9 1 11 2
14 3 2 3 4 9 13 9 1 9 2 13 15 4 2
11 11 13 11 12 9 16 13 0 9 1 11
31 11 13 13 15 0 7 0 9 1 9 1 11 1 12 9 7 15 13 1 0 9 9 1 9 2 13 4 1 9 11 2
21 2 16 14 4 9 7 11 14 13 15 9 2 11 13 4 13 9 1 9 9 2
18 15 4 0 9 7 13 4 0 9 2 2 13 4 0 9 11 11 2
35 11 4 1 9 2 12 9 2 0 16 1 0 9 9 13 9 1 13 15 0 9 1 11 7 15 13 1 0 9 9 1 9 1 11 2
24 2 9 13 2 2 13 4 1 12 9 1 11 0 9 11 11 2 15 9 13 0 9 11 2
21 2 16 14 4 9 7 11 14 13 15 9 2 11 13 4 13 9 1 9 9 2
11 15 4 0 9 7 13 4 0 9 2 2
33 3 9 1 0 9 9 1 9 1 11 1 9 12 9 2 11 4 13 9 1 9 0 9 1 11 1 0 9 9 2 3 11 2
43 3 2 11 1 3 13 13 9 7 9 0 11 9 1 15 9 2 3 9 1 15 0 9 2 11 13 16 11 3 13 15 9 1 12 9 1 9 0 9 9 0 11 2
38 11 4 0 1 0 9 1 12 9 2 3 4 11 13 9 9 1 9 9 1 0 9 0 11 2 0 1 9 11 2 15 15 13 9 11 1 11 2
20 9 9 2 0 9 2 11 2 13 4 3 0 9 1 9 11 1 9 9 2
25 11 4 0 1 0 9 7 9 9 9 1 0 9 2 7 11 4 13 9 7 9 9 1 9 2
11 13 15 16 4 9 13 15 9 12 9 2
26 9 9 11 13 4 9 12 9 3 2 3 15 4 13 1 9 1 9 11 1 11 12 7 12 9 2
19 11 2 14 13 13 9 11 2 1 9 9 11 2 13 4 11 1 9 2
8 2 9 4 4 0 1 15 2
12 0 9 4 1 16 15 9 13 15 9 2 2
27 9 11 1 9 11 11 2 15 3 9 13 1 0 2 9 2 1 9 1 11 2 13 4 9 0 9 2
25 2 4 15 0 3 12 9 1 11 16 12 7 12 9 2 2 13 4 11 1 0 9 1 9 2
30 2 0 9 9 13 4 15 12 9 2 0 15 2 15 4 13 4 0 9 1 9 9 4 14 11 13 15 9 2 2
13 1 9 2 11 4 13 16 14 13 13 15 9 2
27 2 13 1 9 1 15 4 2 2 13 4 1 9 0 9 9 7 9 9 11 11 2 16 13 9 11 2
9 2 9 11 3 4 0 7 0 2
11 9 11 4 15 15 4 13 15 9 2 2
12 11 2 11 7 11 13 9 1 9 9 0 9
31 11 2 11 7 11 13 4 15 1 9 0 0 9 15 4 15 2 3 13 0 12 9 2 1 9 2 13 9 1 11 2
32 1 3 1 12 9 9 1 9 9 11 2 11 2 11 2 11 7 11 13 4 12 9 9 1 9 2 3 9 1 9 9 2
29 9 9 11 7 11 11 11 7 11 11 2 13 4 9 3 1 0 9 9 7 9 11 11 1 9 0 1 11 2
19 2 15 4 3 0 0 9 1 9 15 0 0 9 2 2 13 4 11 2
33 9 0 12 9 9 13 9 9 9 12 9 15 4 15 0 0 9 13 1 0 9 11 1 0 9 1 11 2 1 0 9 11 2
27 9 4 4 0 1 0 9 11 7 1 0 9 0 1 11 2 3 4 11 13 0 9 1 12 9 9 2
15 9 4 3 9 4 0 1 11 2 7 3 1 0 11 2
33 9 2 15 4 2 3 15 13 2 13 0 12 9 2 13 4 11 9 0 0 9 1 11 2 3 15 9 3 13 1 3 9 2
14 3 2 3 9 0 9 9 13 15 1 15 0 9 2
17 13 15 16 4 15 0 9 13 0 2 0 7 0 9 0 9 2
8 9 4 4 9 12 9 3 2
12 0 0 9 1 0 9 9 13 12 9 9 2
34 15 9 3 4 13 4 0 1 12 9 9 1 0 9 7 12 9 9 1 0 9 2 1 9 0 9 1 12 9 9 0 9 3 2
24 0 9 1 9 13 4 12 9 2 7 4 13 3 13 1 9 12 9 1 0 7 0 9 2
35 1 9 0 7 0 9 0 9 2 15 4 12 9 13 0 9 11 2 0 4 16 4 9 11 2 11 4 0 2 0 7 3 0 9 2
20 2 9 4 13 1 15 4 15 1 0 13 1 0 9 2 2 13 4 11 2
43 3 9 0 9 2 0 9 11 11 13 15 4 16 2 0 9 2 15 15 13 9 1 9 9 1 0 9 14 3 1 9 15 4 1 15 0 2 3 7 1 0 9 2
26 7 12 1 12 9 4 13 9 1 9 9 2 2 15 4 13 9 15 4 0 1 9 7 9 9 2
16 0 0 9 11 2 0 0 9 11 2 13 4 9 9 9 2
32 1 0 9 2 1 9 9 2 13 15 0 11 11 2 0 9 11 8 8 8 2 0 9 11 7 11 2 7 0 9 11 2
7 11 13 0 9 1 9 11
26 12 9 1 3 4 9 13 0 9 11 1 0 9 2 0 9 0 1 9 1 9 13 4 1 9 2
23 11 13 1 9 16 4 1 0 9 13 9 0 9 11 11 1 9 9 1 0 0 9 2
30 1 9 2 12 9 2 9 11 11 11 2 9 0 9 7 9 9 13 4 9 0 9 11 11 1 0 9 15 9 2
23 11 15 13 9 0 9 2 9 7 0 9 2 15 4 13 9 1 15 9 7 13 9 2
20 9 11 11 3 4 13 9 0 9 1 9 15 4 0 1 9 3 4 0 2
21 11 4 0 1 12 9 1 9 11 11 2 3 3 9 1 0 9 9 1 15 2
26 0 9 0 9 1 0 9 11 11 7 9 0 9 2 2 0 0 9 2 2 13 15 1 9 9 2
17 0 9 1 9 2 13 15 1 9 2 0 4 1 0 11 9 2
21 1 9 4 0 0 0 9 1 0 0 9 2 7 9 4 0 7 9 9 9 2
29 16 15 15 1 15 15 13 16 4 3 0 1 9 13 1 9 2 9 3 3 13 13 15 4 13 7 13 9 2
16 0 9 0 4 1 9 1 0 9 7 9 1 15 0 9 2
22 1 15 15 11 0 13 9 12 9 12 9 2 13 4 9 16 4 4 0 0 9 2
19 15 9 3 4 13 9 0 9 0 9 11 11 1 11 12 9 12 9 2
18 3 2 11 13 4 15 9 1 9 2 3 16 15 13 16 0 9 2
31 3 15 1 0 9 1 11 11 4 3 13 16 2 3 13 2 1 9 2 3 16 4 1 15 13 2 3 13 9 2 2
16 1 15 4 0 0 9 2 13 4 11 2 3 13 1 9 2
35 0 9 2 1 11 11 2 13 4 0 9 1 9 2 3 9 9 11 7 11 11 2 0 9 7 9 9 7 9 2 16 13 1 9 2
22 3 15 7 11 2 15 15 3 13 1 11 1 0 9 15 9 2 13 1 9 9 2
33 9 0 9 13 4 3 9 15 4 13 11 2 7 9 2 2 3 0 9 0 9 11 11 2 2 13 16 9 4 0 0 9 2
19 2 4 4 0 9 7 9 2 2 13 9 11 11 2 9 9 1 9 2
23 3 2 13 16 4 3 16 4 9 4 0 1 0 2 0 9 0 0 9 3 0 11 2
13 9 3 13 9 9 0 9 1 11 2 1 11 2
13 9 3 13 13 1 9 9 16 15 13 9 9 2
17 1 15 2 9 0 9 11 11 2 9 7 0 13 4 0 9 2
6 9 11 2 11 9 9
19 0 0 9 1 11 7 11 3 4 0 1 12 9 9 0 9 1 9 2
19 0 9 0 9 0 4 16 9 0 9 1 9 9 1 15 9 0 11 2
16 1 12 9 9 2 0 9 1 11 7 11 0 4 12 9 2
19 0 9 0 9 0 4 16 9 0 9 1 9 9 1 15 9 0 11 2
8 3 2 0 4 3 0 9 2
13 3 2 9 0 9 3 13 13 7 9 0 9 2
31 2 0 9 13 0 9 2 2 13 11 11 15 13 9 1 11 1 15 9 1 0 9 2 16 7 1 0 7 0 9 2
11 2 3 2 0 9 13 15 3 0 9 2
9 3 4 13 9 7 13 9 2 2
25 9 9 15 4 13 7 9 9 3 4 13 1 9 0 9 2 15 4 9 15 15 9 13 3 2
14 0 9 13 4 16 4 15 9 13 1 9 9 9 2
9 3 2 0 9 13 12 9 3 2
20 1 9 9 1 0 9 1 11 2 0 7 0 9 13 15 1 0 9 11 2
15 9 13 1 11 1 12 2 12 3 7 12 2 12 3 2
25 13 15 1 9 11 9 2 11 11 2 11 2 11 2 11 7 11 9 2 3 15 9 1 11 2
25 0 0 9 9 11 2 11 0 4 1 9 0 9 2 3 4 9 9 0 9 13 9 1 11 2
27 3 2 13 15 16 4 3 13 2 16 3 3 4 4 0 9 9 9 7 9 2 7 13 4 7 9 2
11 16 9 15 13 4 1 9 9 0 9 2
14 3 1 3 12 9 0 4 9 2 7 9 3 13 2
23 16 13 0 9 2 0 7 0 9 0 9 4 4 0 1 11 2 3 12 9 1 9 2
16 9 7 9 2 11 9 11 13 1 9 1 9 1 0 0 9
15 11 11 1 11 13 4 0 9 1 9 1 9 1 9 2
22 3 1 9 15 9 2 13 0 9 0 9 2 7 1 11 0 0 0 0 9 9 2
33 11 11 1 11 13 9 1 9 9 1 9 1 9 1 9 2 12 9 2 1 12 11 0 0 9 15 4 0 1 11 1 11 2
27 11 11 11 13 4 1 9 2 12 9 2 0 9 1 9 1 9 1 9 1 12 11 0 9 1 11 2
5 13 4 12 9 2
22 0 9 11 4 13 0 9 1 0 9 1 9 1 9 1 0 15 4 0 1 11 2
18 0 0 9 0 9 0 4 1 9 2 12 9 2 1 11 1 11 2
30 9 2 15 15 13 1 9 2 9 12 9 2 2 13 0 9 9 2 7 1 9 4 4 0 0 9 1 0 9 2
18 11 15 1 9 2 12 9 2 13 1 9 9 7 0 9 3 9 2
12 0 9 1 11 13 4 3 12 9 1 9 2
34 0 0 9 9 1 11 0 4 1 9 2 12 9 2 1 11 2 7 1 15 4 13 9 1 11 2 11 2 11 7 0 0 9 2
12 9 9 13 16 13 3 12 15 9 1 9 2
31 9 2 11 2 2 9 2 0 9 11 11 13 4 1 9 2 12 9 2 9 1 0 9 1 12 9 0 9 1 11 2
25 11 11 1 9 2 11 2 13 4 9 1 0 9 1 9 2 15 4 13 1 12 9 1 9 2
40 0 0 0 9 2 0 0 9 1 11 2 13 4 1 9 2 12 9 2 2 7 1 15 4 4 0 3 12 0 0 9 2 12 0 9 7 12 0 9 2
18 9 2 15 15 13 1 9 2 12 9 2 2 0 4 1 0 9 2
24 11 11 13 4 11 2 15 4 1 9 9 0 9 1 9 11 2 1 15 9 2 8 2 2
18 11 4 13 1 9 9 11 12 15 4 0 1 9 2 12 9 2 2
24 0 9 2 9 2 9 2 9 11 11 11 13 4 1 9 1 9 11 15 4 0 1 11 2
23 0 9 13 4 1 9 2 12 9 2 0 9 1 9 9 0 9 9 0 9 11 11 2
21 9 9 15 4 0 9 4 4 0 9 11 2 0 9 7 0 9 1 0 9 2
11 11 13 11 1 9 9 1 0 9 7 9
31 11 0 9 13 13 0 9 1 9 0 9 7 9 1 0 9 7 9 2 13 4 1 9 1 11 0 9 11 1 9 2
7 0 9 0 9 11 11 2
42 3 9 1 9 0 9 0 9 2 11 2 1 9 11 1 9 1 11 2 0 0 9 13 4 1 9 2 12 9 2 11 1 9 9 1 9 9 15 3 13 11 2
41 2 11 13 16 4 1 11 13 1 0 9 1 9 0 9 1 9 0 9 2 7 3 3 13 9 15 13 0 9 2 2 13 4 0 9 11 1 9 11 11 2
55 1 15 0 9 9 11 1 9 2 15 4 0 1 9 2 11 13 4 16 15 9 2 16 15 13 13 11 1 9 12 9 2 13 3 13 1 9 1 9 1 9 9 2 9 2 9 2 0 9 2 9 7 0 9 2
20 0 0 9 2 15 13 4 0 12 9 2 13 4 9 0 0 9 0 9 2
30 3 4 4 0 9 13 14 11 13 1 11 12 9 12 9 2 7 13 13 15 9 1 9 9 1 9 1 0 9 2
12 9 11 13 4 1 9 9 1 9 15 9 2
37 11 13 13 0 2 0 9 1 9 0 9 2 9 9 0 9 7 1 9 1 0 9 7 9 2 13 4 11 1 9 1 9 0 9 11 11 2
33 1 9 1 9 11 11 2 9 11 13 4 11 1 0 9 15 4 13 1 9 2 3 9 0 9 0 9 7 9 0 0 9 2
18 3 2 13 4 16 4 0 9 0 1 9 9 9 2 9 7 9 2
20 11 4 3 13 9 1 9 9 16 13 9 1 0 9 15 13 13 1 9 2
55 1 9 2 0 9 11 11 11 7 9 9 7 0 9 11 11 7 11 11 13 4 15 1 9 11 1 9 11 11 1 9 1 11 2 3 13 15 16 9 13 0 9 1 9 15 9 1 9 9 1 0 9 7 9 2
36 11 2 15 4 13 9 3 3 1 9 9 2 13 4 11 1 0 0 9 1 9 2 3 3 16 4 0 9 4 0 9 1 0 9 9 2
29 3 12 9 0 4 1 11 1 12 9 1 9 0 9 7 0 9 2 7 1 3 15 4 0 1 15 0 9 2
8 9 9 1 4 13 1 0 9
26 16 9 7 0 9 13 13 9 7 13 15 1 9 2 9 13 1 9 16 12 1 9 1 9 9 2
15 14 3 7 3 0 9 13 11 16 4 13 1 0 9 2
20 9 15 13 1 9 12 9 2 7 9 0 9 3 4 0 13 9 1 9 2
18 0 1 9 2 3 1 0 2 15 9 3 13 1 9 7 9 0 2
13 0 4 16 12 9 15 0 9 14 13 1 9 2
25 2 9 0 2 2 7 2 9 9 2 2 3 4 15 1 9 1 0 9 0 1 9 3 9 2
21 9 9 1 15 15 13 9 7 0 0 9 3 15 13 1 9 2 3 0 9 2
42 15 9 2 1 9 1 0 9 2 11 2 2 13 16 3 13 9 9 1 15 4 0 9 2 2 1 0 9 9 9 2 2 13 1 0 9 1 15 15 13 0 2
22 15 9 4 4 0 2 1 15 0 9 7 9 9 2 2 13 4 9 11 11 11 2
14 0 2 1 0 9 1 11 2 0 4 0 9 9 2
26 9 9 11 11 13 4 9 16 13 15 9 0 2 7 3 0 1 0 9 7 9 0 1 0 9 2
30 2 1 0 11 3 4 13 15 2 9 2 0 1 9 0 0 9 2 16 7 0 1 0 9 2 2 13 4 11 2
9 9 9 0 4 1 9 0 9 2
22 9 11 11 13 16 9 9 9 13 13 15 9 2 7 4 3 0 16 13 0 9 2
21 2 15 4 13 1 9 7 9 9 2 3 1 9 1 9 15 15 13 1 9 2
13 13 3 15 0 9 2 2 13 4 11 1 11 2
17 0 2 13 4 2 3 4 0 1 9 9 7 9 9 15 9 2
12 2 13 9 2 3 0 9 2 2 13 4 2
17 1 15 9 2 3 4 3 0 9 16 3 15 15 13 1 9 2
14 16 2 9 0 7 9 1 0 9 3 3 4 0 2
10 2 15 4 0 9 2 2 13 4 2
32 3 16 4 9 13 13 0 0 9 1 9 7 9 2 9 13 0 0 9 16 4 13 1 9 2 3 0 0 9 9 11 2
19 0 0 9 1 9 0 2 11 2 7 15 9 3 13 15 9 1 11 2
19 1 15 2 15 9 13 0 9 9 3 9 3 13 13 15 9 7 9 2
22 3 2 9 9 9 9 2 7 3 7 3 4 13 9 2 13 1 11 9 11 11 2
18 2 11 15 1 11 13 3 3 1 9 1 0 9 7 0 0 9 2
21 15 15 13 9 1 11 3 4 15 15 4 3 13 16 13 2 2 13 4 11 2
13 3 2 13 4 2 15 4 0 9 3 1 9 2
21 11 4 3 13 9 1 0 9 1 9 0 9 2 11 2 7 0 9 1 11 2
33 0 4 9 9 15 4 13 0 9 11 11 2 7 15 13 11 15 4 13 13 9 16 13 16 15 13 1 0 9 9 9 11 2
23 11 13 15 16 4 15 9 9 2 9 9 9 9 9 2 7 9 0 9 11 11 2 2
28 2 2 11 2 13 13 9 9 0 9 2 1 15 2 16 9 0 9 2 2 13 4 0 9 11 11 11 2
32 0 9 0 1 9 13 4 16 4 0 9 9 2 0 2 0 2 0 7 0 2 2 0 1 9 1 0 0 7 0 9 2
15 13 4 16 11 0 3 15 15 14 13 13 16 4 13 2
20 1 15 2 0 9 13 4 9 1 11 1 0 9 1 9 2 9 2 8 2
18 1 9 2 15 9 1 11 13 9 16 4 13 15 0 9 7 9 2
17 1 0 9 9 4 0 9 11 11 7 9 9 0 9 11 11 2
22 11 1 11 3 13 9 1 15 9 2 3 1 0 9 7 3 3 0 9 3 11 2
5 11 13 9 1 9
11 0 9 13 4 9 7 9 9 1 9 2
10 9 1 9 13 4 0 9 1 11 2
20 1 9 16 0 9 13 9 9 2 9 1 0 9 13 15 3 13 1 9 2
30 1 9 16 4 9 1 0 9 2 15 13 16 4 9 1 0 9 2 2 3 9 7 0 0 9 2 2 13 0 2
43 9 9 9 7 0 9 11 11 13 4 1 11 16 14 13 0 9 1 11 1 9 2 9 2 2 9 15 15 13 1 9 0 9 1 12 9 1 9 9 7 9 9 2
15 15 13 13 4 15 2 1 0 9 7 9 1 9 9 2
14 2 1 9 2 9 4 13 0 0 9 1 9 9 2
30 1 9 15 13 2 0 4 9 9 9 2 0 15 4 1 9 9 7 15 15 4 1 9 1 9 2 2 13 11 2
17 12 1 9 4 15 15 4 9 3 3 13 2 7 3 3 13 2
26 1 15 9 2 0 9 3 15 13 2 12 9 9 15 13 1 9 1 0 9 2 2 13 4 11 2
35 15 4 2 9 9 1 9 2 9 0 9 1 9 2 0 9 2 9 15 15 13 1 0 9 7 9 2 9 0 9 7 9 15 9 2
26 11 4 3 0 9 1 11 15 4 13 9 1 9 2 16 4 1 15 0 9 15 9 0 0 9 2
16 2 9 9 9 4 0 9 1 9 7 0 2 1 0 9 2
26 1 3 4 9 1 9 1 0 9 4 0 2 1 9 16 15 0 13 13 9 2 2 13 4 9 2
29 16 15 13 0 9 2 13 4 2 9 4 13 4 0 9 1 12 9 1 12 9 2 1 3 7 1 9 9 2
15 3 4 13 15 4 2 7 15 4 9 2 13 4 11 2
21 2 0 15 3 13 1 9 7 9 2 3 16 4 15 9 9 9 2 7 4 2
11 15 4 0 9 1 9 2 2 13 15 2
21 9 13 16 4 3 13 9 1 9 2 16 13 3 4 15 13 9 1 0 9 2
28 2 13 16 4 9 13 3 1 9 2 16 0 13 1 15 16 4 15 9 7 9 13 1 9 15 15 13 2
33 15 15 4 13 13 9 2 1 9 16 4 1 15 7 13 1 9 7 4 13 1 9 16 13 1 9 2 2 13 0 11 11 2
17 11 11 2 12 2 13 16 4 9 4 3 0 1 9 9 9 2
38 2 9 4 1 9 3 13 9 2 16 15 2 15 4 9 1 9 9 1 11 2 14 13 16 15 9 1 9 14 13 3 13 2 2 13 4 11 2
12 9 7 9 2 0 0 9 13 4 0 0 9
21 0 0 0 9 0 0 9 11 12 2 0 9 2 13 4 0 9 1 9 9 2
10 3 1 9 2 11 13 0 0 9 2
27 0 9 9 0 2 0 9 9 9 0 0 9 9 12 1 11 11 2 13 13 0 0 9 1 9 9 2
27 1 9 9 2 11 4 13 0 9 3 11 9 9 2 15 4 0 0 9 13 15 15 4 13 9 9 2
15 11 4 1 9 2 12 9 2 13 9 1 0 0 9 2
13 11 13 13 9 1 9 1 15 9 1 12 9 2
11 9 13 13 15 9 1 11 1 12 9 2
20 0 9 13 9 3 12 9 0 9 1 3 12 9 9 1 3 1 12 9 2
22 0 9 13 13 12 0 9 1 0 9 16 4 13 9 1 9 9 7 9 1 9 2
15 9 4 3 13 0 9 1 9 0 9 7 13 9 9 2
37 0 9 1 9 11 2 1 9 1 9 9 7 9 9 2 13 4 9 9 0 9 2 9 2 9 9 7 9 1 9 15 15 3 13 16 9 2
10 15 9 0 4 9 9 3 1 9 2
32 0 9 2 3 2 13 13 1 9 9 7 9 2 1 9 9 9 2 15 4 0 9 0 9 2 16 7 1 9 0 9 2
22 3 12 9 7 9 9 4 0 9 2 13 4 1 9 2 12 9 2 0 9 11 2
17 1 9 9 2 11 13 1 2 9 9 2 2 16 7 9 11 2
27 0 9 1 0 7 9 1 0 9 1 11 13 4 1 9 2 12 9 2 1 0 11 9 1 12 9 2
7 9 15 13 1 11 9 2
9 9 9 4 8 9 1 0 11 2
21 0 9 2 0 9 7 0 0 9 2 0 4 1 9 2 12 9 2 1 11 2
11 1 9 4 0 1 0 9 7 9 9 2
19 9 4 13 9 0 9 2 9 11 11 7 9 1 9 7 9 1 11 2
7 11 2 9 2 7 14 9
25 9 1 0 9 14 13 0 9 9 7 3 13 9 9 2 13 1 11 9 9 0 9 11 11 2
11 9 3 0 9 11 13 9 1 9 11 2
33 11 11 2 9 9 0 9 1 9 1 11 2 11 7 11 2 11 2 11 11 7 11 2 13 1 11 1 0 9 1 9 11 2
12 11 2 13 14 13 9 1 11 1 9 11 2
22 11 11 2 1 0 2 9 7 9 9 1 9 11 14 13 16 9 0 9 4 0 2
34 11 4 1 15 13 9 2 1 9 16 15 13 0 9 2 15 4 3 13 11 7 11 9 1 15 0 9 2 16 7 1 9 9 2
12 1 15 2 13 9 1 9 7 9 1 11 2
5 15 4 3 0 2
16 15 13 9 13 2 3 2 15 9 13 4 0 1 0 9 2
12 9 1 0 9 0 4 9 15 15 13 13 2
16 11 2 16 4 15 0 9 7 11 13 13 1 15 0 9 2
33 11 2 11 4 13 9 1 15 15 15 13 1 9 2 12 9 2 7 13 16 4 15 9 15 4 13 9 1 11 13 13 9 2
32 15 15 11 7 11 13 2 7 12 7 0 4 13 13 0 9 1 0 9 9 1 9 7 9 9 9 7 9 1 15 9 2
34 3 2 13 4 13 0 9 15 15 4 0 1 9 1 15 16 4 15 9 0 14 3 1 15 0 2 3 7 1 9 11 7 11 2
28 11 2 0 9 1 11 7 11 1 11 0 4 1 9 2 3 4 15 2 1 15 9 2 13 9 1 9 2
18 11 2 14 13 16 4 13 13 1 15 15 4 4 0 9 9 9 2
23 3 2 14 13 16 4 0 0 9 1 11 7 11 13 0 9 1 15 3 15 15 13 2
13 0 4 16 4 13 0 9 7 9 1 12 0 2
23 3 4 16 4 9 16 15 0 0 9 2 16 4 15 12 9 13 7 13 1 0 9 2
8 14 13 16 4 15 15 13 2
28 3 2 13 13 16 0 9 13 0 9 9 7 13 15 0 9 1 9 9 1 9 11 7 11 7 1 9 2
15 11 2 11 4 13 1 9 1 9 1 0 9 1 9 2
26 3 4 2 1 15 9 2 11 7 11 13 1 15 9 7 3 4 15 0 9 13 13 1 0 9 2
27 11 2 3 3 2 14 4 13 13 1 0 9 2 16 13 16 4 15 1 9 13 13 0 7 0 9 2
27 9 4 13 4 1 9 0 9 2 16 4 1 15 9 9 11 9 1 9 11 2 11 7 0 0 9 2
41 3 2 1 15 9 11 4 13 3 13 1 15 0 9 2 7 15 4 16 15 13 9 1 0 0 9 15 13 9 11 7 11 7 2 1 0 9 2 0 9 2
17 11 2 15 4 9 0 9 13 1 9 9 11 7 11 1 11 2
17 15 11 1 15 9 13 13 16 4 13 9 9 7 13 15 11 2
23 11 2 16 15 4 3 13 2 0 9 9 2 3 1 0 9 2 0 4 1 0 9 2
24 9 1 12 9 13 13 9 7 13 9 16 15 9 13 2 7 4 15 13 9 9 15 9 2
16 11 7 11 4 13 3 13 15 9 7 13 15 9 13 13 2
26 16 4 15 0 9 2 3 4 13 13 16 4 0 2 1 0 2 13 0 7 0 9 1 9 11 2
9 9 2 9 9 4 13 9 9 11
32 9 9 9 11 13 4 1 9 0 9 9 9 1 11 7 13 16 4 15 0 9 4 0 3 9 1 9 9 1 9 9 2
21 9 9 9 11 13 4 1 11 1 9 2 12 9 2 2 1 0 9 9 9 2
22 9 9 2 0 9 1 11 11 11 13 4 16 15 9 9 0 9 11 14 13 13 2
27 2 9 1 0 9 3 14 4 13 4 9 0 9 2 2 13 4 11 1 0 9 0 1 9 1 11 2
16 12 9 11 13 4 1 11 1 9 1 9 1 9 1 11 2
14 9 9 13 4 11 2 12 1 12 0 9 9 9 2
29 11 13 11 1 15 9 9 1 9 11 15 4 13 0 0 9 11 11 2 7 15 15 13 1 2 0 9 2 2
13 11 15 13 9 7 13 1 9 0 9 1 9 2
18 11 11 13 4 1 9 9 3 15 1 2 0 9 2 16 0 9 2
21 0 11 2 2 15 13 12 9 1 3 12 9 9 9 2 2 13 4 0 9 2
22 9 15 9 2 15 4 15 13 1 9 11 2 13 4 9 16 4 15 13 15 9 2
16 0 9 11 11 13 4 9 16 4 9 9 13 9 0 9 2
28 2 3 4 13 3 11 13 4 0 7 3 14 13 4 0 9 2 2 13 4 11 2 7 13 9 1 9 2
16 2 1 15 9 9 4 1 9 1 9 11 2 2 13 4 2
22 9 9 1 9 9 11 13 4 9 0 9 11 2 0 9 11 7 0 9 9 11 2
18 9 4 3 13 11 11 2 3 4 0 9 12 9 13 12 0 9 2
31 11 11 2 0 11 15 4 13 12 9 15 0 9 13 2 2 13 15 16 4 15 13 15 15 4 11 13 3 2 2 2
8 14 13 3 13 1 15 2 2
29 1 9 8 8 8 1 9 0 4 9 9 11 11 16 13 16 4 11 4 1 9 13 9 2 1 9 9 2 2
39 2 15 9 15 4 0 7 9 15 4 13 9 2 9 7 12 9 0 4 3 2 7 15 13 4 7 3 0 13 9 15 0 9 2 2 13 4 11 2
13 9 0 0 9 11 11 3 13 0 9 16 11 2
30 0 9 13 4 1 9 1 11 1 9 16 4 9 0 9 1 11 13 3 1 15 15 9 9 9 13 1 9 11 2
12 3 4 13 9 16 4 11 3 13 15 9 2
22 2 13 15 16 11 13 16 4 11 4 0 1 15 7 15 9 2 2 13 4 11 2
38 2 15 4 7 4 0 1 0 2 0 9 15 15 13 9 0 9 7 4 1 15 13 1 0 9 7 3 4 13 0 11 2 15 4 4 0 2 2
6 11 3 13 0 0 9
14 1 3 1 9 0 9 9 11 2 9 4 3 0 2
14 9 13 16 4 15 0 9 2 16 9 4 3 0 2
20 11 4 13 15 0 0 9 1 9 9 11 1 12 0 9 1 0 12 9 2
40 9 2 0 1 9 9 7 9 2 13 4 9 0 2 15 13 16 4 0 9 13 13 1 9 9 0 9 2 1 15 15 4 13 9 16 15 15 4 13 2
48 1 9 0 12 9 9 2 15 4 0 12 9 1 9 1 9 9 7 9 7 9 0 9 11 8 2 12 9 9 11 13 15 9 2 15 4 1 9 11 11 2 0 9 0 0 11 9 2
39 1 0 9 2 0 9 11 11 11 11 13 4 16 9 13 13 3 9 9 1 0 9 1 0 9 9 2 7 16 4 0 9 4 0 3 12 9 9 2
30 2 9 11 11 13 0 9 15 9 7 9 1 0 9 2 3 0 7 0 11 2 2 13 1 9 15 9 0 11 2
9 1 11 4 13 13 4 15 9 2
21 9 13 3 9 0 1 9 9 9 1 12 0 9 2 1 11 2 11 7 11 2
25 15 9 13 16 0 9 4 13 0 9 9 1 0 12 9 2 7 16 4 13 15 9 7 9 2
27 1 15 2 9 4 13 15 9 1 9 1 0 12 9 7 4 15 4 0 13 0 9 7 9 1 9 2
10 3 4 13 13 12 9 0 9 3 2
23 0 9 4 9 0 0 9 0 1 11 7 15 9 7 9 9 0 1 9 1 12 9 2
41 1 15 2 9 9 11 13 4 3 1 15 4 0 16 4 9 0 9 9 2 3 16 4 9 1 9 11 4 0 1 9 11 11 2 15 4 4 0 0 9 2
20 3 4 13 16 4 9 15 4 0 9 13 13 1 9 9 15 0 9 0 2
23 9 4 3 13 9 16 2 1 0 9 9 9 2 15 14 13 11 11 16 13 15 9 2
15 7 3 2 11 11 4 4 0 0 9 1 0 9 9 2
23 1 0 9 9 9 13 4 3 12 9 2 2 8 8 8 2 2 15 4 4 0 9 2
21 11 4 1 9 13 15 9 2 1 9 16 4 4 1 9 1 0 9 15 9 2
30 1 0 9 1 9 7 9 1 9 0 9 2 9 13 16 4 15 9 0 1 11 2 3 3 1 9 9 1 9 2
21 1 9 11 11 2 0 9 1 9 1 0 9 2 2 15 0 9 4 0 2 2
25 2 3 4 16 4 4 0 9 7 0 9 16 4 9 0 0 4 9 2 2 13 4 1 11 2
17 9 4 13 2 0 2 3 15 13 1 9 2 16 4 3 0 2
31 2 9 12 9 11 13 12 9 9 2 1 15 9 15 4 13 12 9 1 12 9 9 2 15 4 0 9 2 2 13 2
7 11 4 13 9 1 9 12
14 1 0 9 11 0 4 0 9 15 3 0 9 9 2
27 11 4 13 9 1 12 9 9 1 11 1 9 9 0 0 9 12 9 2 9 2 15 13 1 15 9 2
25 9 4 4 0 1 9 9 0 9 9 1 9 12 9 2 1 11 11 7 11 2 1 9 9 2
19 15 4 15 3 13 7 9 0 9 2 16 7 9 9 1 0 9 9 2
31 2 9 9 9 1 9 12 9 2 11 4 13 9 1 15 0 0 9 2 2 13 4 9 9 9 11 11 1 9 9 2
16 9 9 13 2 0 9 1 9 9 0 9 2 2 13 4 2
21 9 9 1 0 4 9 1 0 9 2 16 7 1 0 9 1 9 2 13 9 2
9 2 9 12 0 4 0 0 9 2
42 11 4 13 15 9 9 16 1 0 2 16 7 1 0 9 1 11 2 11 2 11 7 11 2 1 9 1 3 12 9 9 2 2 13 4 9 11 1 9 11 11 2
21 9 7 9 0 9 13 4 9 12 9 2 16 4 0 9 4 0 1 12 9 2
47 2 1 9 9 2 2 2 9 9 0 4 1 9 7 9 12 0 0 9 7 9 12 0 1 11 2 11 2 11 11 7 11 2 2 13 4 1 11 11 11 2 9 0 9 1 9 2
15 13 4 16 4 9 3 13 9 9 9 1 9 0 9 2
17 9 1 9 0 9 13 4 4 0 1 9 12 9 2 13 4 2
23 1 3 0 9 2 0 9 13 13 1 9 1 9 9 9 2 16 3 16 9 15 9 2
20 11 15 13 16 4 9 9 13 9 9 1 9 9 7 0 0 9 1 9 2
18 2 15 9 15 4 9 13 9 9 9 1 9 0 9 1 9 12 2
26 0 9 2 13 4 9 2 0 9 2 1 11 2 2 13 11 11 2 9 9 1 9 1 9 9 2
22 9 9 13 9 9 1 12 9 2 9 9 9 1 12 9 7 0 9 1 12 9 2
8 0 9 13 15 9 3 0 2
26 2 0 9 1 15 9 0 4 9 9 1 11 2 15 4 0 0 12 9 9 2 2 13 4 11 2
15 11 4 13 3 12 9 9 1 11 1 9 0 9 11 2
21 0 0 9 13 4 3 12 9 9 2 16 4 9 13 12 9 1 0 9 11 2
7 0 9 13 1 9 0 9
18 9 3 11 13 15 7 13 9 0 9 0 1 9 7 9 15 9 2
45 0 9 13 0 9 1 11 7 2 2 1 0 9 9 1 0 0 9 7 9 9 2 2 15 9 2 1 9 13 3 0 7 13 15 16 9 13 3 9 7 9 15 13 2 2
44 3 1 15 9 2 11 11 2 15 4 1 9 0 9 11 1 11 2 13 4 16 4 0 9 13 9 15 13 11 2 11 2 11 2 11 7 11 7 13 1 15 0 9 2
41 2 13 4 9 7 9 1 9 1 11 7 4 0 2 0 2 9 1 9 9 2 1 9 9 1 11 2 1 9 1 0 9 9 2 2 13 4 11 1 11 2
14 13 4 16 15 0 9 13 1 9 2 9 7 9 2
31 9 15 4 13 1 15 9 13 4 0 9 11 11 2 9 0 9 1 11 2 15 4 3 13 0 9 1 9 0 9 2
9 9 4 0 0 9 7 0 9 2
43 2 13 4 15 9 3 9 0 7 0 9 0 9 2 15 9 2 9 2 9 2 9 2 9 2 15 4 13 9 0 9 1 9 9 9 1 11 2 2 13 4 11 2
29 11 11 2 9 0 0 9 11 2 13 16 11 13 0 0 9 1 11 2 7 13 11 2 11 2 11 7 0 2
55 9 2 14 13 3 13 9 1 15 4 4 0 13 7 2 13 2 15 9 2 16 15 13 16 4 0 9 9 7 9 7 3 3 0 2 7 15 9 14 13 3 3 4 15 13 1 0 9 2 2 13 4 1 11 2
28 11 11 2 9 9 0 1 0 9 1 11 2 13 4 16 2 3 12 9 11 1 11 7 11 13 0 9 2
24 0 9 9 15 0 9 4 9 1 9 9 9 1 9 7 9 9 2 2 13 4 1 11 2
16 9 4 0 1 11 2 3 4 0 9 13 9 1 12 9 2
10 2 15 9 4 16 15 4 4 3 2
13 15 2 11 2 3 13 13 15 4 4 9 11 2
23 14 13 16 15 13 9 7 14 13 15 13 2 2 13 4 1 11 11 1 11 11 11 2
16 11 11 2 9 0 9 9 1 0 9 2 13 0 0 9 2
26 2 0 4 9 1 0 9 0 1 0 9 2 2 7 4 3 2 1 15 9 3 0 1 0 9 2
28 0 9 0 4 9 1 0 9 11 2 7 15 4 9 1 0 2 0 7 0 9 2 2 13 4 1 11 2
10 1 0 9 1 11 2 11 4 9 2
14 2 16 13 13 15 2 16 9 2 2 13 15 13 2
16 15 15 15 4 13 16 14 13 2 2 13 4 9 11 11 2
34 1 11 4 13 16 4 0 9 9 9 9 11 2 9 1 9 9 1 11 7 11 2 16 7 0 9 9 0 7 15 9 1 11 2
17 11 1 11 13 16 11 3 13 13 9 1 9 0 9 1 11 2
29 2 11 13 13 15 9 2 16 4 13 1 9 11 7 13 13 1 11 7 15 4 15 13 13 2 2 13 4 2
9 11 11 4 9 0 9 1 11 2
27 2 14 13 15 16 9 0 9 2 16 4 3 15 15 15 3 13 13 16 4 2 2 13 4 1 11 2
40 11 11 1 0 9 1 11 13 4 1 11 16 9 13 1 9 1 11 2 16 4 9 1 15 2 15 4 15 7 15 4 15 2 1 15 9 4 11 2 2
10 14 0 9 0 9 13 9 1 0 9
21 1 0 9 2 14 0 9 9 13 15 9 7 15 13 1 0 9 1 0 9 2
36 9 1 11 13 14 0 9 1 9 7 9 9 2 2 16 7 1 9 0 9 1 9 7 1 9 3 2 1 0 0 9 1 15 9 9 2
33 1 9 0 9 0 9 2 12 9 0 9 3 4 1 9 9 15 15 7 13 2 16 3 12 1 12 9 0 9 13 0 9 2
18 9 9 7 9 13 4 0 9 1 9 15 9 2 3 1 0 9 2
19 2 1 12 9 15 4 0 1 12 9 2 12 3 13 7 4 15 13 2
39 15 9 0 4 0 9 7 3 4 9 13 13 9 9 0 9 2 16 15 4 3 0 1 11 2 2 13 4 1 11 11 11 2 9 9 0 9 11 2
34 1 12 9 4 4 12 9 9 9 1 0 11 2 7 12 9 2 15 4 13 0 9 1 9 0 1 9 2 1 12 7 12 9 2
14 9 4 3 13 1 12 9 2 15 4 13 12 9 2
23 15 9 4 12 1 12 9 3 9 2 7 7 12 0 9 15 13 9 4 13 1 9 2
51 2 3 4 9 9 2 7 13 1 9 0 9 9 2 1 9 1 9 1 0 9 12 2 12 9 2 16 7 1 9 9 9 1 0 9 2 2 13 4 1 11 11 11 2 9 11 9 9 0 9 2
24 1 11 2 12 9 9 13 16 3 13 13 9 7 4 0 2 7 12 9 13 13 0 9 2
39 2 15 4 3 3 9 2 16 13 16 15 0 9 13 13 2 13 7 13 15 9 1 0 9 15 9 2 2 13 4 1 11 11 11 1 9 0 9 2
27 0 9 11 11 2 15 4 0 1 0 0 9 1 11 12 9 2 13 4 1 11 16 9 4 4 0 2
28 13 4 15 0 9 2 2 9 11 2 2 1 12 9 2 1 9 1 9 1 9 11 2 16 7 0 9 2
23 2 4 4 9 3 4 13 0 9 2 16 4 13 16 4 13 13 9 2 2 13 4 2
10 3 4 11 13 13 3 9 9 3 2
17 2 13 4 1 0 9 2 3 0 2 7 3 3 15 4 9 2
38 3 3 2 9 1 15 9 13 4 15 1 9 7 16 9 2 13 4 15 3 9 2 3 16 15 13 15 9 7 9 2 2 13 4 11 1 11 2
27 9 1 11 3 13 9 1 9 7 0 9 2 7 14 3 13 9 1 9 9 2 9 2 9 7 9 2
25 9 1 0 9 13 4 16 9 0 9 9 13 9 2 2 15 4 3 3 0 9 1 12 9 2
37 3 2 1 11 4 15 0 9 2 16 7 3 14 13 9 7 9 1 9 9 0 9 1 9 9 2 7 13 0 9 1 9 9 15 13 9 2
31 9 9 1 9 2 11 2 12 4 1 0 9 15 2 3 1 0 9 11 2 3 13 0 9 9 9 7 9 0 9 2
28 2 1 0 9 9 13 0 9 2 7 9 13 3 0 9 0 9 9 2 2 13 4 9 9 11 11 11 2
20 1 9 11 2 9 1 11 3 15 13 9 2 7 3 9 2 9 7 9 2
9 3 12 9 15 13 1 0 9 2
10 9 2 11 13 16 9 13 13 1 9
24 1 9 11 2 0 9 13 4 9 1 9 1 11 7 13 9 0 11 16 13 9 1 15 2
19 3 15 9 2 0 9 11 11 13 1 9 11 11 16 4 13 0 9 2
26 0 9 11 11 2 3 2 13 1 15 0 9 11 11 1 15 9 1 11 1 9 2 12 9 2 2
18 11 4 13 16 4 12 9 0 9 1 0 9 0 11 1 9 11 2
27 0 9 11 11 13 4 1 9 2 12 9 2 1 11 16 4 13 9 9 15 4 13 9 0 9 11 2
18 3 15 13 1 9 11 11 2 9 11 11 7 9 0 9 11 11 2
16 3 1 9 2 11 4 13 9 0 11 16 13 9 1 15 2
29 13 4 16 9 1 9 1 11 13 9 0 7 0 9 2 16 7 9 1 9 1 0 9 2 0 9 7 9 2
24 0 9 11 11 13 4 1 9 2 12 9 2 1 11 11 16 4 13 0 9 1 15 9 2
29 3 1 0 9 2 13 4 16 4 11 13 12 0 9 1 0 9 7 13 0 9 1 0 9 1 9 0 9 2
22 9 9 7 9 9 11 11 7 9 9 1 0 9 11 11 3 4 15 13 9 9 2
40 9 9 9 4 15 13 1 11 12 9 16 15 4 15 4 3 0 2 13 4 1 9 2 12 9 2 8 8 2 3 16 4 9 0 1 9 7 9 9 2
23 9 1 9 3 4 4 13 9 11 11 11 2 9 11 11 11 7 9 11 11 11 11 2
25 1 9 9 11 11 0 4 16 4 0 9 15 4 13 11 15 9 4 0 9 1 9 11 11 2
21 0 9 11 8 11 13 15 1 9 2 12 9 2 1 0 9 0 9 11 11 2
13 9 4 4 0 1 0 9 7 9 1 0 9 2
28 11 15 1 9 13 1 9 11 11 16 4 13 9 9 2 3 9 1 9 2 9 2 9 2 9 7 9 2
21 0 9 11 11 13 4 1 9 2 12 9 2 9 0 0 9 1 11 11 11 2
8 0 9 13 15 11 1 9 2
20 11 4 13 9 11 1 9 12 9 7 13 0 9 1 11 1 9 0 9 2
23 9 11 1 9 1 11 11 11 13 15 1 9 2 12 9 2 1 9 11 11 1 11 2
7 11 4 13 11 12 9 2
6 11 1 9 1 9 11
29 9 11 13 14 13 9 9 15 4 13 1 9 0 9 11 7 13 9 2 7 13 9 1 15 9 1 9 11 2
9 9 9 11 11 7 9 13 9 2
11 9 1 9 0 0 0 9 1 9 11 2
43 11 13 13 13 14 13 9 0 9 11 1 0 9 16 14 4 0 0 0 9 2 7 13 9 2 13 4 1 9 2 12 9 2 0 9 9 2 9 7 9 11 11 2
29 15 9 13 4 3 1 12 9 1 15 4 11 13 12 9 9 1 9 9 15 4 13 4 0 1 9 12 9 2
26 11 4 13 4 15 0 7 0 9 1 9 15 9 2 13 4 11 1 9 1 0 9 9 11 11 2
23 9 2 0 12 9 1 11 2 3 4 13 11 11 2 9 11 2 0 9 0 0 9 2
34 3 9 16 2 0 2 2 11 4 3 13 1 9 16 11 7 13 15 13 2 2 7 4 0 2 2 13 3 9 1 3 0 9 2
24 11 11 2 9 0 0 9 2 9 0 9 2 11 2 2 0 4 9 9 7 9 1 11 2
33 2 2 0 2 11 13 15 1 0 0 9 2 3 15 9 13 0 0 9 2 2 13 4 11 0 9 3 1 0 9 9 11 2
16 2 11 4 13 13 9 15 15 13 0 0 9 1 11 2 2
27 9 11 2 2 9 0 9 1 9 2 2 13 4 16 11 13 3 12 9 15 0 9 1 0 9 9 2
11 14 13 9 1 0 0 9 2 13 4 2
12 3 9 2 13 4 2 15 13 0 0 9 2
24 9 1 9 0 9 3 15 3 13 15 2 3 16 15 9 11 13 1 9 1 0 0 9 2
24 11 15 3 3 13 1 9 13 14 13 9 1 9 9 3 4 1 3 13 1 9 7 13 2
15 7 2 13 4 11 1 9 0 0 11 2 13 0 9 2
11 3 4 2 3 15 13 2 11 15 9 2
34 11 4 1 9 13 9 16 4 15 9 2 16 15 13 9 1 9 9 11 2 3 13 1 9 0 9 15 4 13 13 3 9 9 2
26 16 15 13 9 11 2 13 4 2 9 4 4 0 1 9 2 2 16 15 4 4 2 2 1 11 2
13 2 15 4 9 15 4 13 9 2 2 13 4 2
24 11 4 13 16 4 9 11 13 12 9 9 1 9 11 2 15 4 9 13 13 12 9 9 2
20 9 4 16 11 13 12 1 12 9 9 1 9 1 9 1 3 12 9 9 2
25 3 2 1 9 0 9 1 0 9 13 15 16 4 9 3 1 9 13 13 12 9 9 1 9 2
37 2 13 9 16 0 9 13 15 9 2 7 16 11 13 14 13 15 2 11 4 13 0 9 7 13 0 9 1 15 2 2 13 4 0 9 11 2
12 11 4 3 1 9 0 1 0 9 7 9 2
21 16 15 9 11 13 2 13 4 13 0 9 11 1 0 9 15 4 1 9 11 2
9 11 13 9 9 9 1 11 7 11
35 3 16 15 15 9 13 3 12 9 9 1 9 0 7 0 9 2 9 0 9 11 11 11 13 13 9 11 7 11 1 15 7 0 9 2
36 9 0 9 11 11 11 13 4 1 9 2 12 9 2 1 11 16 4 13 1 0 9 9 11 7 11 15 4 15 13 1 0 7 0 9 2
19 0 9 3 4 4 0 1 12 9 1 11 2 7 4 0 1 9 11 2
27 11 4 1 9 13 3 0 9 1 11 16 7 9 11 2 3 4 13 1 9 7 0 9 0 0 9 2
30 15 9 9 4 9 9 0 9 1 9 9 11 7 11 1 0 9 1 0 7 0 9 2 9 0 9 7 0 9 2
14 1 15 4 13 12 9 1 15 4 0 0 0 9 2
33 12 9 13 4 15 1 0 9 0 1 9 0 7 0 9 2 16 15 7 3 13 1 0 9 2 3 7 15 15 13 13 9 2
17 3 4 9 1 0 9 9 2 12 9 13 3 0 1 15 9 2
29 0 9 13 4 1 9 0 0 9 1 0 9 7 9 1 11 2 16 15 11 13 9 2 9 2 1 0 9 2
29 2 4 4 9 9 1 9 0 7 0 9 7 1 9 9 2 7 4 13 13 9 12 9 2 2 13 4 11 2
16 3 4 13 0 9 1 9 15 9 9 9 15 4 13 11 2
12 2 0 4 12 9 2 9 9 7 0 9 2
13 3 2 13 13 0 9 15 9 2 2 13 4 2
39 0 9 13 1 9 0 9 11 11 11 1 9 9 9 9 2 3 4 15 2 3 15 13 2 13 9 0 11 7 11 16 13 0 9 11 3 15 9 2
27 3 3 0 9 11 2 11 4 1 9 11 1 0 9 11 12 9 15 4 13 0 9 1 9 1 9 2
20 0 9 1 11 1 0 9 13 9 2 16 11 13 15 9 0 9 1 9 2
34 0 9 1 11 11 11 13 4 15 9 16 4 9 2 12 1 0 9 2 2 7 16 11 4 13 9 0 9 3 16 4 15 0 2
25 12 9 13 4 13 9 2 13 4 11 2 3 16 4 9 11 16 15 9 13 13 1 9 9 2
15 7 11 7 11 4 13 13 0 15 13 2 13 4 11 2
9 11 11 13 13 2 0 0 9 2
17 0 0 9 11 11 13 4 9 1 15 0 0 9 2 11 2 2
12 15 4 0 0 9 2 7 13 3 0 9 2
17 0 0 9 11 11 13 4 9 1 15 0 0 9 2 9 2 2
11 0 9 0 4 12 9 1 0 9 11 2
30 15 4 4 0 0 9 11 15 4 1 9 4 0 1 11 2 16 4 11 2 11 2 11 7 11 9 1 15 9 2
10 2 0 4 12 9 2 2 13 9 2
33 2 3 2 16 15 13 0 9 15 4 13 9 1 9 9 2 7 3 16 15 13 1 9 15 4 15 13 9 0 0 9 2 2
26 9 2 15 13 9 9 9 7 11 2 0 4 0 9 1 0 9 15 15 13 1 9 1 0 9 2
22 13 15 16 4 9 4 0 1 9 9 2 7 9 4 13 4 0 1 9 0 9 2
8 9 9 3 4 13 1 9 2
17 12 1 15 2 0 11 11 11 3 4 13 1 9 16 0 9 2
12 9 4 13 12 9 7 13 15 1 12 9 2
22 9 15 3 13 1 11 2 16 4 1 15 7 11 2 11 2 11 9 7 9 11 2
12 9 9 11 11 12 4 1 0 9 1 11 2
33 0 9 11 11 2 0 1 9 1 9 11 11 2 0 4 1 9 2 7 11 11 15 4 13 1 9 9 2 9 2 1 9 2
21 11 15 13 9 2 1 9 2 15 4 12 9 13 0 9 1 0 9 1 11 2
15 1 15 0 9 2 9 2 0 9 4 4 0 0 9 2
9 9 11 11 11 2 13 2 0 9
36 11 11 2 0 0 9 15 4 13 9 2 13 4 0 9 9 0 9 11 15 4 15 3 13 9 0 9 1 9 2 2 0 9 0 9 2
28 0 11 9 11 11 2 15 4 13 1 11 11 2 11 11 7 11 11 2 13 4 0 9 1 9 0 9 2
28 15 9 0 4 1 11 1 9 9 1 0 9 2 15 4 13 13 9 0 9 0 9 1 0 9 0 9 2
36 3 15 15 4 3 13 4 0 9 2 13 15 9 16 15 9 13 15 15 13 9 9 15 9 2 15 4 0 1 15 15 4 1 9 9 2
25 1 9 0 9 2 9 4 13 0 9 13 9 9 2 1 0 9 1 0 9 1 0 9 9 2
16 4 0 13 14 0 9 11 7 0 0 9 11 7 9 9 2
27 9 9 9 15 4 0 0 9 0 4 9 0 9 15 13 0 7 0 9 7 0 9 0 9 11 11 2
37 0 9 13 4 16 4 15 0 2 3 16 4 9 9 0 9 1 9 9 11 11 2 15 3 4 0 13 9 15 13 1 15 0 9 1 9 2
24 3 0 11 3 4 9 13 12 9 1 9 2 3 16 4 13 1 0 9 7 13 4 15 2
11 3 2 13 4 16 15 4 15 0 9 2
17 1 9 12 0 0 9 2 9 0 9 0 4 1 12 9 9 2
19 1 11 2 1 9 0 9 0 4 8 8 8 2 16 7 15 0 9 2
24 11 13 12 9 1 9 2 7 1 9 0 9 2 16 0 9 3 3 4 3 13 15 9 2
16 9 1 9 0 9 1 0 9 9 7 9 1 9 4 9 2
31 3 2 15 4 0 1 11 2 3 16 9 7 9 9 13 0 9 1 9 16 4 13 0 9 16 13 15 9 1 9 2
10 15 4 4 0 0 9 1 0 9 2
16 1 15 2 13 4 13 9 0 0 9 1 11 2 11 11 2
17 3 2 0 4 15 13 3 9 1 0 9 2 9 7 0 9 2
12 9 4 1 9 13 9 1 9 1 0 9 2
9 14 13 9 9 1 9 0 9 2
27 11 13 3 13 7 13 9 7 4 13 13 9 16 4 11 2 1 15 13 9 2 3 13 15 1 11 2
6 11 7 11 13 0 9
21 11 13 9 11 1 9 1 9 1 11 2 16 7 9 0 9 1 15 0 9 2
28 3 9 9 11 1 9 1 11 2 11 4 1 9 2 12 9 2 13 9 9 15 0 9 1 9 1 9 2
12 11 4 1 9 15 9 13 0 9 1 9 2
26 1 9 2 11 4 1 0 9 12 9 13 9 1 9 2 3 16 15 12 9 12 9 3 13 11 2
36 3 2 11 4 13 11 16 15 13 13 1 0 9 0 9 2 3 9 1 0 9 7 9 0 9 2 16 13 13 16 14 13 1 9 9 2
18 9 11 3 4 13 11 1 9 0 9 1 9 9 7 9 1 9 2
51 0 9 11 11 11 11 13 4 1 9 16 4 15 9 13 11 1 9 9 11 2 3 15 1 15 9 3 13 9 0 9 7 3 1 15 15 9 1 9 9 9 7 0 9 2 13 4 0 9 11 2
18 3 4 13 9 0 9 1 11 2 3 1 9 9 2 9 7 9 2
31 2 13 4 9 0 9 2 2 13 4 11 1 0 0 9 1 9 11 11 2 15 4 1 9 13 1 0 0 9 11 2
24 3 1 15 1 11 4 13 7 9 9 11 11 2 9 0 9 11 11 7 9 9 11 11 2
31 9 0 9 2 15 4 3 1 9 9 11 2 13 4 3 9 7 13 1 0 9 1 15 4 0 1 9 15 13 11 2
38 0 9 13 4 2 3 15 13 2 9 1 12 0 9 2 15 2 3 4 15 13 9 0 9 11 11 2 13 12 9 0 0 9 2 11 2 11 2
34 12 1 0 9 9 2 13 4 11 1 9 2 4 4 9 12 9 1 9 2 0 9 2 16 4 15 13 9 11 1 11 12 9 2
30 9 2 3 15 13 2 13 9 0 0 9 1 9 9 12 9 1 0 9 1 0 9 11 2 1 15 9 1 9 2
23 11 7 15 0 9 11 11 11 1 9 4 13 9 1 9 1 9 9 0 9 12 9 2
35 1 0 9 0 9 2 11 4 0 9 2 9 11 2 2 15 15 13 0 9 9 15 4 0 1 11 2 1 15 9 9 0 0 9 2
11 2 3 4 0 0 9 15 15 4 0 2
25 1 15 9 11 13 9 0 9 2 9 2 9 2 9 7 9 2 2 13 4 0 9 3 9 2
24 11 2 0 0 9 2 13 4 9 1 9 1 11 2 8 16 15 1 3 9 13 1 11 2
13 0 9 2 11 7 11 11 13 1 9 13 1 11
35 9 0 0 9 11 11 13 15 1 9 1 9 11 7 11 11 2 3 16 0 9 9 13 1 9 15 0 9 2 1 0 9 1 11 2
36 9 0 0 9 11 11 13 4 0 9 11 7 11 11 1 11 16 15 9 3 13 9 1 0 9 1 0 0 9 1 0 11 2 11 2 2
20 1 15 9 2 9 11 7 11 11 1 9 0 9 13 1 9 15 0 9 2
23 11 4 13 16 9 11 11 7 9 0 7 0 9 13 4 0 1 11 14 4 3 3 2
17 11 4 12 9 0 1 9 3 9 9 1 11 1 11 7 11 2
14 9 9 9 13 1 0 9 0 1 0 11 12 9 2
41 11 4 1 9 2 12 9 2 1 11 13 1 9 11 11 11 11 2 9 11 11 11 2 9 11 7 11 11 11 11 7 9 0 9 11 7 11 11 11 11 2
33 11 4 13 16 3 3 13 16 4 11 13 13 9 9 9 1 11 2 7 3 16 15 15 13 2 15 9 15 13 13 1 11 2
12 1 15 9 2 9 7 9 11 3 4 0 2
30 2 16 0 9 2 11 4 13 9 9 1 9 9 9 2 3 16 4 2 3 0 9 15 9 7 9 1 11 2 2
23 11 4 13 9 1 0 0 9 11 11 7 11 11 7 0 0 9 11 11 7 11 11 2
13 13 15 16 4 11 2 11 7 11 0 0 9 2
23 11 4 13 1 11 3 1 9 9 9 12 9 2 7 0 9 4 0 3 15 3 13 2
21 0 9 13 4 4 0 11 1 0 9 2 7 1 15 15 3 13 13 0 9 2
37 1 9 13 14 16 0 9 13 0 15 4 1 15 9 1 9 7 9 11 2 11 4 13 2 2 3 3 15 13 13 2 16 11 13 4 0 2
17 15 13 13 1 11 7 0 9 13 4 0 1 9 15 9 2 2
19 9 0 9 11 11 13 4 16 15 9 16 15 11 13 1 11 13 3 2
19 9 11 7 11 11 13 4 9 11 1 15 9 16 11 13 0 0 9 2
12 0 0 9 13 4 1 9 1 11 0 9 2
19 11 4 3 13 16 15 9 9 15 9 2 13 13 1 9 9 9 2 2
19 2 0 9 4 9 15 4 3 13 0 9 0 9 2 2 13 4 11 2
8 0 9 11 13 0 9 1 11
34 0 9 11 11 13 4 0 9 1 9 11 1 0 9 1 11 2 3 9 11 16 4 11 13 0 9 1 9 1 9 1 12 9 2
34 3 0 9 1 0 0 9 1 0 11 2 11 2 2 0 9 11 11 13 4 9 0 9 11 1 9 11 9 9 1 9 1 9 2
18 11 2 15 3 3 4 13 9 9 2 13 15 9 11 1 12 9 2
26 2 13 0 7 0 9 1 9 2 2 13 4 11 1 9 2 12 9 2 1 15 0 0 9 11 2
39 0 4 14 0 13 0 0 9 11 11 2 12 1 9 0 9 1 0 9 1 9 11 2 11 4 13 2 3 13 0 9 2 3 7 13 0 9 2 2
19 11 4 0 9 1 9 13 16 0 9 1 9 9 11 1 9 1 9 2
15 0 9 15 11 13 13 13 0 9 7 9 9 0 9 2
35 2 15 4 13 9 1 9 0 9 2 15 13 9 15 9 2 2 13 4 11 3 9 1 9 3 9 0 9 1 9 0 9 1 9 2
11 2 15 4 9 15 0 9 0 9 2 2
20 9 3 13 9 1 11 1 9 0 9 1 11 1 0 0 9 1 0 11 2
36 2 13 4 9 3 3 15 4 13 7 0 9 2 2 3 15 13 2 2 2 13 4 9 9 0 9 2 11 2 11 11 1 9 1 11 2
32 2 14 13 15 13 1 4 15 0 9 2 7 4 3 0 1 9 0 9 2 2 13 4 11 2 16 4 11 13 1 15 2
48 3 11 16 4 2 4 0 9 1 9 0 9 2 1 11 2 11 4 13 16 4 15 9 0 9 12 9 13 1 9 2 16 7 16 4 15 15 1 3 9 13 1 0 9 2 11 11 2
26 11 4 13 0 9 3 3 1 9 9 2 1 9 15 0 0 9 2 11 2 1 0 9 1 9 2
27 11 4 13 9 1 9 1 9 11 1 9 12 2 7 13 15 0 9 0 9 1 0 9 1 9 9 2
23 15 4 15 13 9 1 9 9 0 9 1 9 1 11 7 9 9 1 9 9 1 9 2
21 2 13 15 0 9 9 1 9 12 7 9 12 9 2 2 13 4 11 1 11 2
22 3 15 13 9 9 15 9 2 11 4 13 0 0 9 15 4 13 9 11 1 11 2
22 15 15 13 1 0 9 11 11 2 15 4 9 3 9 9 9 11 2 1 0 9 2
11 11 4 13 9 9 11 1 9 1 11 2
12 11 15 3 13 1 9 1 9 11 11 11 2
20 1 9 1 9 2 9 9 11 2 11 2 13 4 9 1 9 7 9 9 2
12 9 4 13 13 9 9 0 9 1 9 9 2
21 11 15 13 1 9 0 9 1 9 1 0 0 9 15 15 13 1 0 9 9 2
24 2 0 9 4 13 9 9 7 13 0 9 1 9 0 9 2 2 13 4 9 11 11 11 2
11 9 7 9 2 0 9 7 9 13 9 11
21 3 9 11 2 0 9 13 4 9 1 0 9 7 9 15 15 13 9 1 11 2
17 9 11 1 11 13 4 9 1 0 9 7 9 15 15 13 9 2
17 3 0 9 7 9 13 4 9 11 1 9 1 9 9 1 9 2
29 11 11 13 4 9 1 0 9 1 0 9 1 9 1 9 11 2 1 15 9 3 4 0 11 11 7 11 11 2
27 11 11 13 4 9 1 0 9 2 9 4 1 15 9 2 2 16 4 11 11 13 9 1 0 9 9 2
8 9 1 9 13 4 11 11 2
12 9 11 13 4 9 1 9 9 9 9 11 2
28 11 11 11 13 4 12 0 9 1 12 0 9 1 0 9 15 4 1 12 1 12 9 0 1 11 1 11 2
23 11 4 13 9 0 9 1 9 1 9 7 9 2 7 13 1 0 9 1 9 1 9 2
21 0 0 9 2 11 11 11 2 13 4 0 9 1 9 1 9 7 0 1 9 2
20 1 0 9 1 9 0 11 2 11 11 11 13 4 0 9 1 9 1 9 2
22 11 4 13 16 4 11 13 12 9 1 9 0 0 9 11 7 9 11 1 9 11 2
12 15 9 13 4 9 1 9 1 9 15 9 2
16 0 0 9 11 11 13 4 12 9 1 11 1 12 9 9 2
30 11 2 15 4 9 1 11 2 13 15 1 9 1 11 12 9 7 3 13 12 1 0 7 0 9 1 0 0 9 2
12 4 4 9 0 0 9 1 11 7 1 9 2
22 0 0 9 11 11 13 4 9 11 12 1 0 0 9 0 0 9 1 11 1 11 2
15 0 4 4 11 11 11 2 7 0 11 11 1 0 11 2
35 9 0 9 11 11 8 11 2 9 0 2 13 4 7 9 0 9 7 9 1 0 0 9 1 12 11 9 9 2 15 4 0 12 9 2
20 9 0 9 11 11 2 12 2 12 3 1 11 2 13 4 0 9 0 9 2
11 11 2 11 7 11 11 13 9 1 0 9
15 9 12 0 9 3 13 9 0 0 9 1 0 0 9 2
40 1 9 9 9 0 9 12 9 1 11 2 11 2 11 7 11 11 13 4 9 15 15 9 15 12 9 13 9 1 9 7 0 0 9 1 9 15 12 9 2
36 0 9 0 9 11 11 13 4 16 4 15 9 13 7 13 9 9 2 9 9 7 9 1 9 7 9 0 0 9 1 9 9 1 11 9 2
35 2 9 4 1 3 0 9 3 2 16 15 3 13 1 9 9 0 9 1 9 2 15 13 0 2 9 15 4 15 13 7 1 0 9 2
19 0 0 9 15 13 1 0 9 1 0 9 15 9 2 2 13 4 11 2
17 15 0 9 11 11 13 4 9 15 4 15 13 0 9 1 11 2
44 2 15 4 0 9 15 4 13 9 1 9 15 12 9 7 13 9 9 16 4 15 13 0 9 2 9 9 9 7 9 0 9 15 12 9 9 1 11 2 2 13 4 11 2
32 0 9 0 9 11 11 13 4 2 2 15 9 2 1 0 9 2 13 4 9 15 9 1 12 0 9 2 0 9 7 9 2
15 13 0 9 2 9 2 7 7 0 9 0 1 11 2 2
30 15 15 13 1 0 9 11 3 4 13 9 2 3 16 13 9 7 0 9 1 0 9 7 9 1 11 7 11 11 2
16 11 11 2 9 1 11 2 15 9 13 9 1 11 7 11 2
16 1 11 4 13 16 15 9 13 16 4 13 3 9 3 13 2
11 2 3 4 13 13 1 11 11 1 9 2
20 16 13 9 2 3 4 0 16 4 15 3 13 16 4 15 13 7 15 15 2
20 3 2 3 4 1 0 9 3 2 16 15 13 13 7 15 9 15 13 9 2
15 11 11 4 0 9 1 15 7 15 9 2 2 13 11 2
29 11 11 2 9 1 11 9 2 13 4 1 11 16 4 15 0 9 2 7 4 0 1 9 0 9 1 9 9 2
21 2 1 15 4 9 3 16 9 1 9 13 13 1 11 2 7 4 3 0 3 2
25 0 9 13 9 9 2 7 3 15 7 12 9 9 14 4 4 0 13 9 9 2 2 13 11 2
15 13 4 16 9 9 14 13 0 9 1 4 15 1 9 2
58 2 9 13 9 3 1 0 0 9 2 15 13 16 15 1 0 9 4 4 1 9 13 9 2 2 15 15 13 2 0 9 3 1 9 9 7 3 15 2 16 15 0 9 1 11 7 11 11 13 3 2 2 13 4 11 1 11 2
25 13 15 16 4 11 13 0 9 1 11 7 11 11 2 13 11 11 2 9 1 11 9 1 11 2
14 1 11 4 13 16 9 1 0 9 1 11 15 13 2
10 2 3 3 9 13 15 9 1 11 2
26 9 1 0 9 1 11 13 9 1 0 9 2 7 3 4 2 0 2 0 9 1 15 3 4 0 2
19 9 4 16 11 1 11 7 11 11 13 9 1 15 9 2 2 13 11 2
44 11 4 0 9 2 1 9 0 9 1 9 2 9 7 9 2 13 9 9 0 9 1 9 9 2 3 2 0 0 9 2 2 0 0 9 9 9 0 9 1 9 1 11 2
11 0 15 9 3 13 7 1 11 7 11 2
43 11 4 9 13 15 9 16 13 0 9 1 9 1 0 9 9 1 0 9 2 7 9 4 13 16 4 13 7 1 0 9 1 0 9 1 9 0 9 1 9 9 11 2
15 11 13 1 0 9 9 11 1 11 7 0 9 1 0 11
23 11 13 16 11 13 0 9 1 9 11 2 7 13 9 1 0 11 0 9 9 1 9 2
43 0 9 13 4 13 9 1 11 1 0 9 3 12 9 2 16 4 13 0 9 9 1 9 15 9 0 9 2 13 4 1 9 2 12 9 2 0 9 0 9 11 11 2
45 2 13 16 4 3 9 1 0 9 1 0 9 9 2 7 3 1 11 2 2 13 4 0 9 9 1 9 15 4 13 9 1 0 9 2 11 2 2 0 9 1 9 1 11 2
14 2 13 13 1 0 9 15 4 15 9 1 11 2 2
39 1 9 9 2 1 15 4 15 13 1 9 15 4 13 9 1 9 0 9 2 13 4 3 4 0 9 11 7 0 0 9 1 15 9 2 13 4 11 2
32 0 9 3 4 13 13 2 0 9 1 9 11 11 2 1 9 2 3 2 16 9 9 7 11 13 0 9 2 2 13 4 2
46 11 4 13 9 1 9 1 9 12 9 2 7 4 15 9 1 9 13 3 2 1 0 9 1 0 9 9 7 9 11 16 13 15 0 7 0 9 1 9 1 9 9 11 2 11 2
31 1 15 2 15 0 9 9 13 4 16 11 13 4 0 2 0 9 2 1 0 9 2 15 4 9 15 11 13 1 9 2
15 2 14 13 1 9 9 15 15 9 13 2 2 13 11 2
18 2 15 15 13 4 16 15 14 4 0 9 9 7 9 9 1 9 2
15 9 15 15 13 13 13 16 9 1 0 9 13 13 0 2
35 9 0 9 1 11 13 4 15 16 0 9 1 0 9 1 11 2 7 4 15 9 13 13 1 9 9 0 9 1 15 9 2 13 4 2
17 2 14 4 0 9 0 2 14 11 13 0 2 2 13 4 11 2
26 16 15 0 9 9 13 0 9 15 3 0 9 1 11 2 15 9 13 4 15 13 16 11 13 9 2
26 2 13 16 3 15 15 9 4 13 0 9 1 3 9 2 4 4 1 0 11 2 2 13 4 11 2
17 2 15 4 4 9 1 0 11 15 13 0 0 7 9 0 9 2
20 11 15 13 0 9 0 15 9 7 13 9 0 9 15 13 1 15 9 2 2
36 3 2 3 4 13 16 15 11 14 13 13 9 1 11 14 16 13 9 0 9 0 1 9 11 2 7 16 0 11 13 13 13 9 9 11 2
40 11 2 15 9 13 13 0 0 9 11 1 11 12 9 12 9 2 3 13 9 9 9 0 9 2 1 2 9 1 9 2 15 15 3 13 1 0 9 9 2
34 0 0 9 9 1 0 9 12 9 13 15 0 9 0 9 9 0 11 7 9 0 9 2 15 4 0 9 9 15 13 13 15 9 2
34 12 9 3 2 11 4 1 9 9 9 16 15 12 9 1 12 9 2 16 15 0 9 9 15 15 13 9 13 1 0 9 9 9 2
37 11 4 13 16 4 15 2 1 9 9 11 12 9 2 11 13 1 0 0 9 2 9 0 9 1 9 7 0 9 1 9 9 0 11 1 9 2
21 3 13 9 11 2 11 4 13 16 4 11 13 13 9 9 12 9 16 0 9 2
23 3 2 13 4 16 9 9 14 13 7 16 4 3 15 9 13 9 16 14 13 0 9 2
26 11 4 3 13 16 4 2 1 0 0 9 2 11 13 13 0 9 1 9 9 9 1 15 0 9 2
7 11 13 11 11 1 0 9
25 9 9 11 11 7 11 8 1 0 9 2 11 4 13 12 9 1 9 15 13 9 1 0 9 2
57 11 4 0 9 13 9 15 0 9 11 11 1 0 9 2 16 9 4 13 16 4 1 9 9 3 13 7 11 11 2 15 13 11 11 1 9 9 2 11 1 0 9 2 11 11 1 9 7 11 1 0 9 2 1 0 9 2
16 11 4 3 13 12 1 12 9 15 13 0 9 1 0 9 2
32 1 9 9 15 0 9 2 15 4 13 15 0 9 2 0 0 9 2 1 0 9 1 9 0 9 2 4 4 0 1 0 2
15 1 9 9 11 4 13 1 0 9 7 11 9 1 11 2
26 0 9 0 4 9 15 15 13 1 0 9 9 9 9 7 11 2 13 11 11 2 9 11 1 11 2
44 13 15 16 4 0 9 9 1 11 1 12 9 9 15 13 0 9 7 15 4 3 9 15 3 12 1 12 9 11 13 11 2 16 9 0 9 13 16 4 9 9 9 0 2
35 9 1 0 9 9 4 0 9 15 4 9 13 1 0 9 2 16 15 1 9 13 9 9 0 9 1 9 2 16 7 9 9 0 9 2
22 16 9 9 2 9 4 13 3 12 0 9 0 9 2 1 0 9 3 12 9 9 2
29 15 9 13 15 0 9 1 9 9 1 9 7 9 0 9 2 15 4 0 9 15 13 1 9 11 1 9 11 2
26 1 9 9 9 15 4 12 9 13 11 0 4 16 1 11 1 12 9 3 12 13 0 9 11 9 2
18 9 9 11 1 0 9 13 4 3 16 15 9 15 0 9 3 13 2
9 0 0 9 13 0 0 9 0 9
23 12 0 9 1 11 7 11 11 2 11 7 11 7 11 13 4 9 1 9 0 0 9 2
14 15 9 4 0 1 9 1 9 0 9 1 0 9 2
24 12 0 9 1 11 7 11 11 2 11 7 11 2 4 2 7 11 13 13 0 0 0 9 2
17 9 15 0 9 4 9 9 9 1 9 9 1 11 1 0 9 2
48 2 13 15 16 4 15 9 13 0 9 0 9 9 7 9 15 15 13 0 9 9 9 1 9 2 2 13 4 0 9 1 0 0 2 11 2 1 9 0 12 9 1 15 4 0 0 9 2
25 9 4 12 1 9 9 11 2 0 0 9 2 11 2 7 0 9 11 2 9 1 9 1 9 2
19 9 1 9 1 9 9 15 4 15 13 0 9 0 4 9 12 0 9 2
25 16 13 0 9 2 0 15 13 9 16 9 9 2 16 9 0 9 9 2 13 0 9 1 9 2
46 1 9 15 4 11 2 11 7 11 13 1 9 12 9 2 9 4 15 13 13 7 13 15 9 1 9 7 9 9 1 9 1 0 2 3 9 9 0 9 1 9 7 3 9 9 2
37 0 9 0 9 13 9 0 9 9 1 0 9 2 9 9 1 0 9 15 15 13 1 9 2 9 9 9 2 7 0 9 9 7 9 0 9 2
45 2 13 16 4 9 9 2 9 9 7 9 9 1 9 0 9 9 1 0 9 7 9 9 1 9 2 2 13 4 0 9 11 11 11 2 13 15 1 9 15 9 0 1 9 2
38 1 9 9 11 11 11 2 0 9 13 4 16 4 2 9 0 9 2 3 0 9 7 0 9 0 0 9 1 9 0 11 2 0 9 1 0 9 2
28 1 9 9 9 1 9 2 9 11 11 11 13 4 16 0 9 9 13 3 3 13 1 9 9 1 0 9 2
49 2 13 15 1 0 1 0 7 9 2 7 7 1 15 1 15 15 13 9 0 7 0 9 2 16 9 15 4 0 4 3 4 9 0 9 2 16 4 0 1 9 0 9 7 0 9 2 2 2
51 13 15 15 16 4 3 0 13 15 3 13 9 1 9 1 0 9 15 9 2 15 13 1 15 9 9 2 7 3 15 1 15 13 13 0 9 1 3 0 9 15 3 1 15 13 2 2 13 4 11 2
32 1 9 15 0 9 2 1 9 0 9 1 9 1 9 2 12 0 9 13 0 9 1 0 9 7 9 0 9 1 12 9 2
46 9 4 13 9 2 9 7 9 1 0 9 2 16 15 4 0 7 0 9 2 9 1 9 9 2 0 9 2 9 2 0 0 9 7 9 11 2 7 9 1 0 9 1 0 9 2
19 0 0 7 0 9 1 9 0 9 7 9 1 9 13 4 9 7 9 2
15 0 9 13 16 4 9 1 9 1 9 9 1 11 4 0
35 1 9 0 9 0 9 0 0 9 3 4 13 9 1 9 1 9 9 15 4 0 0 9 2 15 13 0 9 1 9 11 7 11 11 2
15 9 15 9 4 4 0 2 13 4 9 0 9 11 11 2
43 9 0 9 2 11 2 1 11 7 11 2 11 2 13 4 1 9 2 12 9 2 16 4 9 9 0 11 1 9 1 0 9 1 9 9 13 13 9 9 1 9 11 2
31 12 0 9 1 11 2 3 0 0 9 2 11 2 2 13 4 12 9 9 1 9 1 0 9 9 9 15 4 13 11 2
15 1 9 4 9 1 9 0 9 9 7 9 9 0 9 2
12 9 9 4 0 9 1 9 11 1 9 11 2
26 9 0 9 13 12 9 13 1 11 16 4 13 9 1 9 12 9 0 1 9 9 11 1 15 9 2
30 0 9 13 4 9 9 9 1 11 1 9 1 9 7 9 2 11 2 2 15 4 0 0 9 1 0 9 1 9 2
48 3 2 0 9 13 4 1 9 16 4 0 9 11 13 13 15 1 9 0 1 9 11 0 9 2 3 16 4 0 9 15 15 0 9 13 9 9 15 13 9 0 2 11 2 7 9 11 2
32 3 15 9 16 2 0 2 2 11 4 1 9 13 16 4 2 16 4 15 9 2 2 9 4 0 1 11 7 0 11 2 2
27 16 4 11 13 15 9 2 15 4 13 16 4 13 13 9 9 1 9 3 1 9 1 11 2 13 11 2
45 9 11 1 9 11 11 13 4 1 9 16 4 1 11 4 3 3 13 16 4 11 13 2 0 9 2 1 9 9 9 16 14 13 0 0 9 1 9 1 9 15 4 13 11 2
34 16 4 11 13 13 9 9 7 0 15 0 9 11 2 15 9 7 9 0 11 13 4 2 9 9 7 9 2 2 13 4 0 9 2
47 2 15 4 13 15 9 2 7 0 11 2 1 9 15 9 2 3 13 9 13 9 1 0 11 7 0 15 15 13 13 1 9 0 9 2 9 9 2 9 7 9 2 2 13 4 11 2
9 0 9 1 11 13 4 0 9 2
32 3 9 1 9 11 16 2 3 0 2 2 0 9 4 13 16 15 15 2 1 0 9 13 9 1 9 1 11 1 11 2 2
9 0 9 1 11 13 4 9 12 9
41 11 2 11 7 11 2 11 2 2 11 11 2 9 0 9 0 9 13 4 1 9 2 12 9 2 16 4 0 9 0 13 9 15 4 0 12 0 9 1 11 2
49 11 4 13 9 0 9 16 4 9 7 0 9 13 9 1 9 0 0 9 0 1 9 1 15 2 9 0 0 9 11 11 11 7 9 9 0 2 11 2 11 11 15 4 1 9 9 0 9 2
11 9 4 0 9 12 9 1 12 9 9 2
9 3 2 11 13 13 1 15 9 2
23 13 4 0 9 16 4 2 0 9 11 15 13 15 1 11 7 0 7 0 9 15 13 2
5 0 0 4 9 2
11 15 1 11 11 14 13 4 15 9 2 2
27 1 9 1 9 2 9 1 11 13 4 9 11 11 7 11 11 1 0 0 9 1 0 9 0 1 11 2
8 9 9 4 4 9 0 9 2
8 0 9 7 9 13 15 1 9
17 9 7 15 9 13 15 1 0 9 2 7 9 4 7 1 9 2
20 9 11 13 1 9 1 11 2 7 9 4 15 9 13 3 0 9 7 9 2
28 2 3 4 1 12 9 13 9 16 4 13 1 0 9 2 7 3 4 13 15 9 1 15 4 15 3 13 2
16 13 4 15 13 2 13 0 9 2 0 9 2 13 0 9 2
23 3 4 1 9 13 13 9 2 7 4 13 3 12 9 2 2 13 4 11 11 1 11 2
11 9 4 13 3 12 9 16 13 0 9 2
12 1 9 4 3 13 13 0 9 1 15 0 2
9 15 4 3 0 9 1 9 11 2
16 1 9 3 13 2 9 3 13 16 4 15 0 3 3 9 2
8 3 2 9 1 15 4 0 2
8 7 9 13 9 11 7 11 2
36 1 0 9 0 9 11 0 4 16 9 0 9 13 3 1 12 9 9 2 9 4 0 12 9 9 2 16 9 1 9 13 3 1 12 9 2
29 2 16 4 13 0 15 9 2 0 4 0 9 11 13 13 3 3 12 9 2 2 13 4 1 11 9 11 11 2
39 0 9 2 15 4 0 1 9 0 9 1 9 2 13 4 16 4 2 16 4 13 15 9 2 11 13 1 0 9 13 12 9 9 2 3 12 15 11 2
36 2 13 16 4 9 9 1 9 15 9 13 9 1 12 11 2 15 4 3 16 15 13 9 2 2 13 4 1 11 11 11 2 9 0 9 2
31 1 11 2 9 4 3 13 12 9 2 9 1 0 9 7 9 1 0 9 2 15 13 16 0 9 14 13 13 12 11 2
25 3 2 14 13 9 7 9 15 4 9 13 16 15 13 15 9 2 7 15 4 9 13 1 9 2
24 2 11 4 13 13 0 9 0 9 16 4 15 9 13 1 3 0 9 2 2 13 4 11 2
27 0 9 1 9 9 11 11 13 4 1 11 16 2 16 9 13 9 2 15 3 3 14 13 1 0 9 2
22 2 16 4 0 9 13 9 9 9 2 15 15 3 13 7 13 9 11 3 1 9 2
16 13 1 9 15 9 13 1 12 9 9 2 2 13 4 11 2
22 1 9 9 2 1 0 9 0 11 2 3 11 7 11 7 11 13 0 9 1 11 2
38 2 11 4 0 9 1 11 7 11 13 13 1 9 1 9 15 4 15 13 1 9 2 7 3 13 9 7 3 9 13 1 9 2 2 13 4 11 2
20 16 9 0 9 13 13 1 9 7 1 15 13 9 2 0 9 13 15 9 2
12 15 9 13 3 1 9 0 9 7 0 9 2
10 7 3 4 7 15 9 4 3 13 2
18 1 9 0 9 2 9 9 3 13 12 9 9 3 16 1 9 9 2
9 0 9 2 11 1 0 9 1 11
22 9 1 11 16 0 9 14 14 13 2 3 1 9 0 9 1 9 1 9 7 9 2
12 3 2 9 15 7 3 13 1 15 0 9 2
27 2 3 14 0 4 2 0 9 12 4 1 0 1 11 2 2 13 4 1 9 0 9 11 11 11 11 2
37 0 0 9 9 3 11 13 4 15 9 1 12 1 0 1 11 2 13 15 1 9 0 9 1 9 1 9 7 9 2 11 2 0 3 15 9 2
45 9 0 9 1 9 2 16 15 4 9 2 9 7 9 2 16 7 0 0 9 1 9 7 9 2 3 4 0 1 0 9 16 1 0 11 2 13 15 1 9 11 1 12 9 2
27 2 3 14 0 4 2 0 9 12 4 1 0 1 11 2 2 13 4 0 9 11 11 11 11 1 9 2
19 0 9 3 13 1 0 0 9 7 9 15 4 13 1 3 0 9 11 2
28 0 9 2 3 1 11 2 13 4 0 9 9 2 16 4 9 9 0 9 1 9 13 9 7 13 9 9 2
36 2 11 15 13 1 9 1 15 4 9 2 0 9 7 9 13 9 1 9 9 7 9 9 2 9 2 9 7 9 2 2 13 15 1 9 2
24 1 11 2 9 9 3 4 0 2 7 3 7 0 2 1 15 15 13 1 4 15 0 9 2
29 2 0 4 0 9 0 9 15 4 13 9 7 3 2 7 15 4 13 11 0 9 2 2 13 4 11 1 11 2
11 0 9 3 13 16 0 9 2 13 11 2
6 9 9 1 9 4 2
9 9 9 7 9 9 3 3 13 2
24 3 2 0 9 2 1 2 9 2 9 7 0 9 2 13 0 9 1 9 2 13 4 11 2
18 2 9 1 9 13 13 9 7 9 1 9 7 9 2 2 13 4 2
42 1 9 15 11 13 16 9 1 0 9 9 9 2 12 9 9 13 4 9 1 12 9 2 1 12 9 1 15 4 9 0 2 15 4 3 1 0 9 1 12 9 2
15 11 4 13 16 4 9 2 0 9 9 12 2 1 11 2
13 9 7 9 2 11 11 13 9 1 9 1 0 9
15 11 11 11 13 4 15 0 9 1 0 9 1 12 9 2
32 3 1 9 9 1 9 7 9 1 15 9 2 0 9 11 11 13 0 9 1 9 2 12 9 1 0 11 13 4 9 11 2
51 2 1 9 2 11 11 1 11 2 0 9 2 2 11 11 1 11 2 0 9 2 7 11 11 1 11 2 0 9 2 13 9 1 9 1 0 9 11 0 0 9 15 4 1 9 0 1 11 1 11 2
28 0 0 9 11 11 13 4 0 9 1 9 1 0 9 11 0 0 9 15 4 12 9 0 1 11 1 11 2
13 4 4 15 0 9 11 1 0 9 1 12 9 2
27 12 9 1 0 11 0 4 1 9 12 9 15 4 13 0 9 1 9 1 9 9 11 2 11 2 11 2
53 9 11 13 4 9 0 9 11 11 2 9 7 0 9 2 2 9 2 9 4 0 7 9 4 1 9 2 2 0 9 11 11 7 9 0 9 11 11 2 1 9 2 2 9 11 2 11 2 11 7 11 2 2
27 0 9 11 11 13 4 12 9 0 9 1 9 1 12 9 9 9 1 0 0 9 1 0 9 1 8 2
14 11 4 13 1 0 9 1 9 1 12 9 0 9 2
21 4 4 15 0 0 7 3 12 9 15 4 11 13 1 0 0 9 1 0 9 2
17 9 9 0 9 11 11 0 4 1 9 2 12 9 2 1 11 2
14 9 2 15 4 13 0 9 2 13 4 1 12 9 2
35 0 9 11 11 13 4 0 9 1 9 1 9 15 4 1 9 2 12 9 2 0 1 11 2 7 15 4 13 12 9 7 0 0 9 2
48 11 4 15 0 9 11 13 2 0 0 9 2 3 16 15 4 15 11 13 1 8 2 11 2 11 1 11 7 11 1 11 2 2 13 4 9 11 11 1 9 1 9 0 9 9 9 9 2
16 1 11 4 1 9 2 12 9 2 0 12 0 0 0 9 2
14 0 9 3 4 13 9 0 0 9 7 0 9 9 2
30 15 9 1 9 13 12 0 0 9 2 11 11 1 11 2 11 11 1 11 2 11 11 1 11 7 11 8 1 11 2
29 0 9 11 2 3 1 11 2 4 4 0 0 9 9 1 12 9 1 9 9 15 4 9 11 13 3 15 9 2
33 1 9 9 0 9 2 11 12 2 2 0 9 11 13 4 1 9 0 9 9 12 0 9 2 7 3 12 9 2 0 15 9 2
4 0 9 13 11
20 1 15 4 3 0 0 9 1 0 9 2 0 9 1 11 13 4 15 9 2
8 9 11 13 1 9 1 9 2
20 1 9 2 12 0 0 9 1 11 3 4 13 15 9 1 0 9 12 9 2
53 1 9 1 9 2 12 9 2 1 9 9 2 0 9 3 1 9 2 15 13 9 11 11 11 2 13 4 9 9 11 2 8 8 8 8 2 2 16 9 1 0 0 9 2 8 8 8 2 2 0 11 9 2
11 3 12 9 7 9 13 4 9 11 9 2
25 3 15 0 2 9 11 11 13 4 9 16 4 2 3 4 0 2 13 0 9 9 1 15 9 2
11 9 0 9 13 0 9 2 13 4 11 2
9 3 4 13 9 9 7 9 9 2
23 11 4 3 13 9 9 0 9 11 11 2 15 4 4 9 11 1 0 9 1 9 11 2
30 1 9 2 3 1 9 3 1 9 2 11 4 13 16 4 3 0 0 9 2 1 0 9 7 0 9 1 15 9 2
21 4 4 3 13 15 9 2 13 4 11 2 15 15 13 1 0 9 1 9 9 2
14 3 2 1 0 9 2 3 13 0 9 2 13 4 2
19 9 9 4 4 0 9 1 15 4 13 1 9 1 3 11 0 9 11 2
27 1 9 0 9 2 9 4 13 12 9 1 9 9 9 0 9 11 11 1 0 0 9 9 1 0 9 2
7 11 15 13 1 0 9 2
15 0 9 11 11 13 4 0 9 9 11 9 0 1 9 2
18 13 4 9 16 13 15 9 7 13 0 9 2 7 0 7 0 9 2
25 1 9 2 0 0 9 11 2 11 13 4 15 0 0 9 15 4 0 9 1 12 1 12 9 2
37 1 9 15 13 16 15 12 1 9 1 0 9 2 2 2 2 13 9 9 9 9 1 9 9 1 15 9 13 0 0 9 2 7 1 9 2 2
40 2 16 4 9 15 9 3 3 0 1 9 9 2 15 15 13 9 1 9 15 0 9 1 0 9 2 3 16 15 13 9 1 9 2 2 13 11 2 11 2
13 11 13 16 4 15 9 9 11 0 1 9 0 9
28 0 9 11 11 11 13 4 1 9 0 9 9 11 16 4 0 9 15 9 1 11 9 0 9 0 0 9 2
21 13 15 16 9 11 11 11 13 15 9 9 11 1 9 2 12 9 2 1 11 2
45 3 15 9 1 9 9 9 11 16 2 0 7 0 2 2 0 9 11 11 11 13 4 1 9 2 12 9 2 16 4 15 0 9 4 9 16 0 9 1 9 13 3 1 9 2
38 3 15 0 9 9 11 2 11 2 1 11 1 11 2 11 4 13 16 15 9 13 9 0 0 9 11 7 11 2 15 4 13 3 3 1 9 9 2
11 15 9 13 9 1 0 9 2 13 4 2
19 2 15 9 9 3 4 0 1 9 0 9 2 13 4 11 15 0 9 2
29 2 15 13 9 1 0 7 0 11 1 15 4 9 7 9 0 9 3 0 7 0 1 9 9 0 1 9 9 2
19 15 3 13 0 0 0 7 0 9 1 9 0 0 0 9 1 11 2 2
21 3 3 3 9 11 2 11 4 1 9 11 1 9 9 1 9 12 2 12 9 2
23 0 11 2 15 13 3 12 9 0 9 9 1 3 12 9 9 2 13 0 9 1 11 2
22 3 11 16 0 9 9 15 9 2 0 9 13 16 4 0 1 15 13 13 0 9 2
19 3 4 0 9 16 4 0 9 4 0 15 9 9 9 0 1 9 11 2
28 2 12 1 0 9 1 15 9 4 4 13 9 7 9 0 9 0 9 1 11 2 2 13 4 11 9 11 2
29 2 0 4 0 0 0 9 2 2 2 2 15 4 9 4 9 9 9 2 7 15 4 3 4 0 9 11 2 2
26 16 4 0 0 9 13 0 9 1 9 9 2 0 9 1 15 4 4 1 0 9 2 13 4 11 2
23 2 4 4 3 0 16 15 11 1 9 7 3 13 9 0 9 0 9 2 2 13 4 2
10 2 11 15 4 4 3 9 0 9 2
15 11 3 13 13 0 9 7 0 9 16 4 13 9 2 2
31 9 11 13 4 1 9 15 9 9 1 11 0 9 0 9 9 15 13 11 2 11 2 11 2 11 2 11 7 0 9 2
27 9 9 3 9 4 13 11 7 11 2 15 4 15 9 2 3 15 13 2 13 1 0 9 3 0 9 2
32 2 15 9 4 13 12 0 1 9 9 2 16 13 13 14 15 0 9 2 2 13 4 1 9 11 2 7 13 0 9 11 2
13 2 4 13 3 7 3 13 1 9 15 4 0 2
23 1 15 9 9 13 13 15 9 7 13 15 9 9 11 3 3 13 0 9 15 9 2 2
9 0 12 9 1 9 1 9 1 11
24 0 9 13 4 1 9 2 12 9 2 16 4 13 12 9 1 9 1 9 9 9 11 11 2
18 3 9 1 9 11 11 2 0 1 9 1 0 9 4 4 0 3 2
29 11 4 13 9 1 12 9 1 9 1 9 1 9 9 11 11 2 3 7 12 9 15 4 3 3 0 1 9 2
24 1 9 0 1 9 2 12 9 2 9 0 9 13 4 11 11 0 0 1 9 1 9 11 2
22 0 9 0 9 2 0 16 0 9 0 0 9 11 11 2 3 3 15 13 1 9 2
10 13 15 16 4 9 0 13 9 9 2
20 0 9 13 4 16 15 11 7 0 0 15 3 3 4 0 2 13 1 9 2
12 15 4 0 9 0 1 9 1 9 1 11 2
21 1 9 12 9 2 9 4 13 0 9 7 13 0 9 0 9 0 1 0 9 2
46 0 4 3 1 12 9 2 3 7 3 9 3 0 9 1 0 9 2 11 2 2 0 9 9 0 9 2 0 1 0 9 0 1 9 1 11 7 11 7 11 2 7 0 0 9 2
37 11 2 15 4 3 0 7 16 9 2 13 15 2 9 2 9 1 9 11 7 13 15 16 4 9 13 3 1 0 9 0 0 9 2 0 9 2
29 11 11 2 9 9 11 2 0 4 3 9 1 9 7 3 4 0 13 4 16 4 15 13 9 15 4 13 11 2
10 9 15 4 0 9 0 4 15 3 2
23 11 2 12 2 4 0 1 0 9 1 9 3 4 13 1 15 9 1 9 9 1 11 2
20 15 0 9 4 13 0 9 1 9 15 4 13 1 9 11 1 9 12 9 2
12 16 9 9 15 4 13 1 0 9 1 11 2
21 15 9 2 16 7 9 0 9 2 15 4 15 13 2 13 4 9 0 0 9 2
27 1 9 9 2 9 4 13 3 9 2 3 9 11 11 7 11 11 2 9 1 9 0 9 11 11 11 2
15 9 13 16 4 9 9 13 9 16 9 4 13 1 9 2
11 11 4 2 3 4 0 2 0 0 9 2
43 13 15 16 4 0 9 0 0 9 11 11 4 1 9 1 9 11 2 7 1 9 0 9 1 9 0 4 16 4 9 1 11 2 0 2 2 14 3 4 15 9 9 2
16 0 9 9 11 13 4 16 4 9 1 11 0 1 12 9 2
29 0 9 0 9 2 11 4 3 9 1 9 11 13 1 11 16 4 15 15 13 1 0 0 9 1 9 1 11 2
13 9 0 9 9 4 13 0 9 0 9 1 11 2
26 1 9 2 11 11 1 9 4 13 9 1 15 15 0 9 13 1 0 0 9 1 9 9 1 11 2
50 15 4 13 9 12 0 9 9 2 11 11 2 9 9 9 11 1 15 4 11 0 2 11 11 2 9 9 9 9 0 9 11 7 11 11 9 9 1 9 11 2 13 15 1 9 9 0 9 11 2
4 9 1 11 11
15 12 1 0 9 0 11 0 15 4 9 1 11 13 9 2
24 11 11 4 4 12 1 0 9 1 0 11 7 12 1 3 3 15 4 13 13 0 0 9 2
18 1 0 4 9 4 0 11 2 7 13 4 0 2 0 7 0 9 2
11 11 4 12 9 1 15 0 9 13 9 2
18 0 4 9 15 9 13 1 9 1 9 16 4 3 3 4 3 0 2
21 1 9 1 0 9 9 2 9 15 4 0 1 9 11 2 3 1 0 9 11 2
20 9 1 11 7 11 13 4 9 11 2 15 4 4 0 9 1 11 7 11 2
33 11 11 2 9 7 9 1 0 9 1 0 9 11 2 13 4 1 11 16 11 2 1 0 12 9 3 4 13 9 2 15 9 2
35 2 4 4 0 9 7 9 2 7 0 7 0 9 2 7 1 15 4 13 9 15 4 13 9 9 0 7 0 9 2 2 13 4 11 2
28 11 15 13 1 0 9 1 9 9 1 0 9 2 7 4 4 9 11 1 0 9 0 11 2 13 4 9 2
31 2 11 4 9 1 9 1 15 4 13 7 9 15 4 13 1 15 9 13 0 9 1 9 0 11 2 2 13 4 11 2
25 11 11 2 9 0 0 9 1 11 2 13 4 1 11 16 4 11 13 2 0 2 9 0 9 2
22 2 13 4 0 16 15 1 9 9 9 11 13 1 2 0 9 2 16 9 0 9 2
30 11 4 9 11 1 9 9 9 13 9 7 13 0 9 1 15 9 11 15 4 13 0 0 9 2 2 13 4 11 2
25 1 12 1 0 9 0 9 2 0 11 13 1 9 7 13 9 0 9 3 2 11 2 11 2 2
10 9 9 1 0 9 13 2 13 2 2
33 3 1 9 1 0 9 2 15 9 7 0 0 9 9 11 11 13 4 16 4 3 13 1 11 2 1 15 4 13 15 0 9 2
19 2 11 4 4 0 11 1 11 7 0 11 1 11 2 2 13 4 11 2
16 11 4 13 1 0 0 9 1 0 11 7 13 0 0 9 2
25 13 4 1 9 7 1 0 0 9 2 3 1 11 2 3 4 13 0 3 9 9 2 11 2 2
6 9 9 1 11 1 9
18 16 4 7 3 1 0 1 9 2 13 9 9 1 11 1 0 9 2
26 1 0 9 9 0 9 1 11 1 9 9 2 11 4 3 0 1 3 0 9 9 7 0 9 9 2
35 3 2 1 3 0 9 9 0 9 2 11 15 13 1 9 0 9 9 2 16 4 1 9 1 15 0 9 1 9 7 3 1 9 9 2
18 3 16 4 12 9 4 12 9 2 9 9 1 9 3 4 1 9 2
16 9 9 11 11 13 16 0 9 1 11 13 9 9 1 9 2
19 13 1 9 0 9 16 1 0 9 15 14 3 9 13 13 3 12 9 2
12 11 3 13 9 9 0 9 2 3 1 9 2
28 9 1 9 7 9 1 0 9 15 4 15 13 13 9 2 15 13 1 9 9 2 13 9 1 9 7 9 2
24 0 9 3 13 13 9 1 15 9 2 15 4 3 12 9 1 15 13 13 9 2 13 11 2
20 9 1 9 9 13 9 9 9 1 0 9 2 7 3 1 9 9 7 9 2
10 1 0 3 12 9 9 13 4 11 2
11 1 9 11 9 15 4 4 1 0 9 2
12 16 4 11 13 9 1 0 2 3 15 13 2
15 9 1 11 0 4 3 9 13 1 9 0 7 0 9 2
14 0 9 13 16 0 9 13 0 9 3 3 0 9 2
9 9 4 3 0 1 0 0 9 2
21 0 9 1 9 1 11 13 16 4 0 9 0 9 15 4 0 13 0 9 9 2
15 3 9 11 13 15 9 2 0 9 1 12 9 1 9 2
10 3 2 15 9 4 3 9 0 9 2
33 1 0 9 2 15 9 13 15 1 9 9 7 13 16 4 9 9 2 15 2 1 15 9 2 13 3 0 9 1 0 3 9 2
26 0 9 9 9 1 11 2 3 1 9 0 7 0 9 9 2 13 4 0 0 9 9 1 12 9 2
18 0 0 9 13 15 1 12 1 12 9 7 12 3 4 13 12 9 2
18 9 9 1 11 2 1 15 9 1 0 9 2 13 1 0 1 9 2
51 1 9 1 9 0 11 2 9 9 1 11 0 4 1 9 2 3 1 11 2 7 13 4 11 7 11 11 2 3 1 9 15 4 13 0 0 0 9 12 9 1 15 0 9 8 8 15 4 0 9 2
14 11 7 9 13 15 1 9 0 0 9 2 0 0 9
10 11 7 15 9 13 9 0 0 9 2
15 9 13 16 4 0 0 9 16 4 15 9 13 13 9 2
7 9 1 9 1 9 11 2
17 9 1 11 7 0 0 9 13 16 0 0 9 13 1 0 9 2
16 0 9 15 15 13 13 4 1 11 2 16 7 1 15 9 2
21 0 0 9 2 15 4 13 9 1 0 9 15 15 13 2 13 4 13 9 9 2
15 9 9 13 4 11 16 4 3 1 9 13 12 9 9 2
29 9 9 2 9 11 13 4 15 9 1 0 12 9 2 1 15 4 2 3 13 9 2 0 9 4 12 9 9 2
24 9 9 7 9 11 11 13 16 4 9 13 1 9 12 9 9 16 9 9 1 9 0 9 2
25 9 9 7 9 11 11 13 4 0 0 9 8 16 0 9 13 9 1 9 16 15 13 1 11 2
14 3 12 9 9 0 0 9 9 4 9 9 0 9 2
33 1 9 8 8 11 1 9 2 12 9 2 2 0 9 13 16 4 2 3 12 9 2 1 3 12 0 9 1 11 2 0 2 2
15 11 11 1 0 9 11 13 4 9 16 9 2 9 2 2
24 1 0 11 2 9 11 11 13 4 11 11 16 4 0 0 9 7 9 15 13 9 13 9 2
26 3 0 9 2 0 9 11 13 16 4 0 9 15 13 1 11 13 9 15 13 13 1 15 0 9 2
20 1 0 9 11 2 11 13 9 9 9 9 7 9 2 12 15 0 0 9 2
34 0 9 11 11 13 9 9 11 1 12 9 1 12 9 2 15 4 2 3 4 13 2 1 9 1 0 0 9 11 11 1 12 9 2
25 11 11 2 0 9 15 13 1 9 8 2 8 8 2 1 15 4 9 15 13 0 9 0 9 2
38 1 15 4 2 0 9 9 0 7 0 9 15 13 2 2 9 2 0 9 1 9 0 2 7 2 9 1 0 0 0 9 1 9 1 0 9 2 2
11 11 13 0 9 1 9 11 1 9 9 9
34 0 9 1 0 9 13 4 1 9 0 0 0 9 9 7 15 9 1 9 9 16 4 13 13 0 9 1 9 0 0 9 11 11 2
22 11 4 13 0 0 9 9 11 11 2 3 2 7 15 9 11 11 1 9 9 9 2
50 0 0 9 9 11 11 7 15 9 11 11 0 4 0 1 9 9 7 0 4 15 0 9 1 9 1 12 2 3 12 9 2 13 4 1 9 2 12 9 2 0 0 9 1 0 11 2 11 2 2
43 9 4 2 0 0 16 4 15 3 7 3 13 1 9 9 3 1 9 15 4 9 4 0 2 2 7 15 4 13 1 9 0 0 9 11 11 2 13 15 1 9 9 2
49 1 9 15 4 1 9 13 0 0 9 11 11 13 15 16 4 1 9 12 9 11 13 11 16 13 1 9 1 15 13 15 0 9 2 1 0 9 0 16 9 12 2 7 13 15 16 14 13 2
32 11 2 15 4 4 0 9 9 9 9 7 0 9 0 9 8 8 2 13 4 9 12 7 13 2 12 0 9 1 15 2 2
12 9 4 3 13 12 9 2 13 15 1 9 2
30 2 0 9 13 4 16 4 9 0 1 15 9 2 16 4 11 2 13 15 9 2 1 11 2 13 15 1 9 11 2
29 11 4 13 0 9 7 13 15 9 16 13 9 1 9 12 2 3 15 16 4 0 15 4 13 1 11 3 0 2
27 9 4 3 13 16 4 0 9 7 9 0 9 1 9 11 11 13 0 9 2 7 9 9 13 4 9 2
31 9 4 13 16 15 11 13 9 12 15 4 13 1 9 7 1 9 13 1 11 7 9 0 9 0 9 11 2 11 2 2
6 9 4 0 9 9 2
27 11 7 0 9 11 11 0 4 0 9 1 0 9 2 16 4 0 9 2 11 11 2 0 0 0 9 2
12 9 1 11 7 0 3 4 1 0 9 11 2
7 13 9 2 0 9 1 11
22 9 1 0 0 11 13 9 2 0 9 1 9 0 9 7 9 1 9 1 0 9 2
12 0 9 13 9 1 0 9 9 9 1 11 2
21 0 9 13 4 12 9 2 7 0 4 1 9 1 9 0 9 7 0 0 9 2
13 9 4 13 12 9 2 3 7 0 9 11 11 2
23 1 9 4 0 9 13 12 0 0 0 9 2 11 11 7 11 2 15 4 0 0 9 2
36 11 4 0 9 13 9 0 9 15 3 13 16 4 4 0 2 1 9 7 0 2 7 3 13 9 1 9 0 7 13 9 0 9 7 9 2
17 4 9 16 15 9 1 11 13 3 13 7 3 13 0 0 9 2
22 0 9 15 13 9 0 11 3 13 16 4 9 3 0 9 7 9 1 9 3 0 2
15 0 9 13 9 0 9 11 8 8 11 1 0 9 9 2
11 0 9 7 0 9 1 11 3 3 13 2
20 0 4 9 15 4 3 4 0 0 9 11 13 15 9 1 0 9 11 11 2
17 9 0 1 8 8 7 12 9 11 13 4 9 0 9 7 9 2
23 13 4 0 9 0 9 2 3 11 11 2 9 8 2 8 8 2 11 2 7 11 11 2
9 0 9 11 11 4 4 0 9 2
27 2 9 4 15 0 9 16 15 13 9 9 2 2 13 4 9 9 11 11 7 11 11 11 1 9 11 2
28 15 9 2 0 4 13 15 11 2 0 4 0 9 11 11 2 11 1 9 9 2 7 15 4 0 9 11 2
23 11 2 15 13 9 11 11 7 11 11 2 13 4 9 0 0 9 2 9 2 1 9 2
9 0 9 3 13 11 2 11 11 2
29 0 4 12 9 0 9 9 11 2 11 2 13 9 1 0 9 2 7 12 4 15 0 9 13 1 9 7 9 2
24 2 13 4 14 3 1 9 0 9 2 3 7 1 9 0 9 2 2 13 4 9 11 11 2
14 0 4 9 1 0 9 11 9 9 13 9 9 9 2
26 9 0 9 9 13 4 0 9 11 11 2 3 0 9 15 4 13 11 9 3 15 1 9 0 9 2
16 0 4 9 13 11 11 2 9 1 11 2 11 9 0 9 2
8 9 13 9 1 0 9 9 2
28 0 9 9 2 15 4 15 9 9 4 2 9 9 2 2 12 4 1 0 1 9 2 7 13 15 9 9 2
9 0 9 0 4 9 1 9 0 2
7 1 12 0 4 9 9 2
17 0 9 11 3 4 13 0 9 9 1 9 1 0 0 0 9 2
26 3 0 9 13 9 13 15 9 2 7 0 9 13 9 13 15 1 9 9 7 13 15 9 0 9 2
15 1 11 15 9 13 1 15 4 9 13 9 1 15 9 2
26 0 4 9 14 0 7 13 0 9 1 9 2 1 9 2 7 15 4 0 2 7 1 9 0 9 2
13 9 8 8 8 11 11 1 11 13 4 15 9 2
8 0 0 9 13 4 15 1 9
21 16 15 13 0 9 2 0 0 9 13 4 2 3 15 13 2 0 9 9 9 2
17 9 11 11 11 11 13 9 16 2 0 9 9 7 0 9 2 2
39 9 0 9 2 11 2 11 11 11 13 4 1 9 2 12 9 2 9 15 0 9 2 3 9 16 4 0 9 1 0 9 13 1 9 11 1 0 9 2
46 2 1 9 9 15 4 13 9 9 2 13 4 13 9 15 13 13 0 9 7 0 9 1 9 1 0 9 1 15 15 11 3 13 2 2 13 4 0 0 9 1 0 9 1 11 2
28 11 2 15 4 13 12 9 11 1 9 12 9 2 13 4 12 9 9 0 9 2 11 2 1 0 0 9 2
28 2 0 4 16 4 15 9 4 0 1 9 11 1 9 7 0 0 0 9 15 13 1 0 2 2 13 4 2
27 12 1 0 9 0 11 12 9 2 4 4 9 0 9 15 13 0 9 2 2 15 13 1 9 1 9 2
13 12 12 0 9 2 3 12 9 2 13 13 11 2
34 1 9 9 0 9 2 15 4 1 12 13 12 9 9 2 9 9 13 9 0 9 2 16 7 9 16 9 9 13 9 7 9 11 2
53 0 9 11 13 4 9 0 0 9 1 11 2 12 2 3 11 2 1 0 0 0 9 2 11 2 2 12 1 0 3 0 7 0 9 2 11 2 7 12 1 0 9 9 7 9 2 11 2 2 9 0 9 2
19 12 0 9 4 4 9 11 1 9 2 16 7 12 4 13 1 9 9 2
18 9 11 1 9 1 9 11 11 13 4 9 9 1 0 7 0 9 2
14 15 0 9 13 9 0 9 7 9 9 0 9 9 2
17 11 4 13 11 11 2 0 9 1 0 9 7 0 9 1 11 2
15 11 4 4 0 1 9 2 16 7 1 9 9 1 9 2
42 3 12 0 9 1 9 13 4 11 11 1 11 2 15 4 0 1 0 9 1 9 7 0 9 2 16 4 0 9 0 9 11 11 4 0 1 0 9 7 0 9 2
12 12 0 9 0 11 13 4 9 1 0 11 2
41 11 11 1 11 0 4 1 0 9 1 0 9 7 9 2 16 4 9 1 9 1 9 2 11 11 1 11 2 4 1 9 9 1 9 2 9 2 9 7 9 2
6 0 9 11 13 1 9
13 3 7 1 0 9 2 11 11 11 4 4 0 2
13 1 0 9 2 9 9 1 9 0 4 1 9 2
13 0 9 11 11 13 4 15 9 1 9 7 9 2
17 3 4 13 0 9 1 11 2 11 4 3 3 4 1 0 9 2
29 3 15 1 9 15 9 2 9 4 3 13 13 15 9 2 3 0 9 12 9 7 3 13 0 9 9 9 3 2
23 0 9 13 4 1 11 1 9 12 9 2 7 3 4 13 9 0 9 1 0 9 11 2
16 0 9 11 11 2 0 0 9 2 13 15 13 9 1 9 2
37 3 2 9 4 15 7 9 15 0 9 4 0 16 4 9 13 13 9 9 11 11 2 0 9 15 4 9 7 0 11 13 11 0 9 1 11 2
21 2 11 4 13 0 9 1 9 9 2 2 13 11 11 2 0 9 9 9 9 2
12 2 9 1 9 1 2 13 11 2 0 4 2
19 7 0 9 4 4 3 0 7 0 16 15 9 4 13 9 1 9 2 2
25 11 11 2 9 1 12 0 9 1 11 2 13 4 3 12 9 3 4 15 13 9 1 15 9 2
13 0 4 12 9 12 9 2 9 3 4 13 11 2
31 1 9 2 0 9 4 13 9 15 9 3 12 9 2 3 4 4 9 9 13 4 15 0 15 9 1 9 1 0 9 2
6 3 4 4 0 15 2
19 3 4 2 9 3 3 0 2 7 3 0 1 15 9 2 2 13 11 2
6 9 4 3 13 3 2
10 9 7 9 13 4 9 1 0 9 2
25 9 0 9 2 15 4 13 0 9 2 0 4 3 7 11 4 13 9 2 15 4 13 0 9 2
23 3 7 3 2 13 0 9 2 7 15 9 0 2 13 15 9 2 2 3 1 9 9 2
27 11 4 2 13 13 9 2 7 4 13 1 0 9 15 4 0 15 13 2 2 13 9 0 9 11 11 2
14 3 2 3 7 1 9 1 9 11 13 0 1 9 2
32 2 0 9 2 0 0 0 9 2 11 11 2 3 2 9 13 2 2 13 15 0 2 13 4 8 8 11 9 9 11 11 2
20 2 15 4 0 9 15 13 2 15 4 9 11 7 0 9 0 0 9 2 2
11 9 0 0 9 13 9 11 16 13 0 9
29 9 0 0 9 11 11 13 4 9 1 11 7 11 1 9 16 4 9 13 1 0 9 16 14 13 0 0 9 2
12 9 0 0 9 11 11 13 4 1 9 11 2
47 11 7 11 2 11 2 13 15 1 9 9 9 2 16 9 9 14 13 13 1 0 9 2 13 4 1 9 2 12 9 2 9 0 0 9 11 11 1 11 2 0 9 15 0 9 11 2
29 2 3 4 0 1 9 15 13 15 9 2 15 9 7 9 15 9 2 2 13 4 11 1 9 3 0 9 11 2
14 0 0 9 1 12 9 0 4 12 7 3 9 9 2
28 3 2 1 0 12 9 13 4 1 9 0 9 15 13 9 12 0 0 9 9 1 9 15 9 1 9 9 2
15 2 3 4 15 13 1 15 9 2 2 2 13 4 11 2
6 2 15 13 13 2 2
25 1 0 9 2 9 15 13 13 1 9 15 4 13 9 9 1 15 9 1 0 9 2 13 4 2
26 0 9 7 9 1 9 9 13 4 1 9 1 9 1 9 7 9 15 4 13 1 11 1 9 12 2
15 2 13 13 15 9 1 11 7 13 0 9 2 2 2 2
11 1 0 9 13 4 1 0 9 1 11 2
15 1 0 9 2 13 4 1 0 9 2 2 13 4 11 2
21 3 4 13 9 11 1 9 1 0 9 16 4 13 0 9 1 9 1 0 9 2
35 0 9 4 4 0 16 9 12 0 9 2 9 0 2 11 2 15 13 0 11 7 9 11 1 15 13 11 7 11 2 0 0 0 9 2
22 9 0 11 13 4 16 4 13 1 9 11 2 16 4 15 0 9 13 1 9 9 2
23 2 13 0 9 13 16 9 15 9 13 13 13 0 0 7 0 9 2 2 13 4 11 2
14 3 4 13 9 11 13 11 1 9 1 15 9 9 2
27 2 9 2 11 2 0 4 16 4 9 15 9 0 9 1 9 4 0 9 0 11 2 2 13 4 11 2
14 2 0 0 9 13 4 15 16 13 1 0 9 2 2
42 3 1 11 2 1 9 15 4 13 1 0 9 11 7 0 0 9 1 11 2 4 4 0 9 11 1 0 9 7 9 11 11 7 0 9 7 0 9 11 11 11 2
31 11 2 0 0 9 15 4 13 11 1 3 4 15 13 9 11 11 12 9 2 13 4 7 1 11 1 9 11 1 9 2
7 0 9 13 4 9 1 9
20 0 9 13 4 9 15 15 13 9 9 9 9 0 1 0 9 1 12 9 2
40 1 9 2 15 4 0 1 0 9 12 9 2 0 9 13 13 9 9 2 3 9 2 9 2 9 2 9 7 9 1 0 9 2 15 4 13 1 12 9 2
16 9 0 0 9 3 4 4 0 1 15 9 9 13 0 9 2
38 2 16 7 0 0 2 7 15 13 1 9 15 4 4 0 0 0 9 1 15 9 2 2 13 4 9 11 11 11 1 9 1 9 0 7 0 9 2
18 16 4 13 9 2 0 9 13 13 9 0 9 1 9 1 9 9 2
21 15 9 13 13 9 2 1 15 4 9 4 0 1 9 9 1 9 9 1 9 2
15 9 1 11 16 9 0 4 0 0 2 0 7 0 9 2
51 0 9 1 9 2 15 4 0 12 9 2 0 4 16 0 9 13 13 0 9 2 15 13 0 9 7 0 9 15 13 2 16 4 12 9 2 1 0 9 0 9 2 0 9 0 9 7 9 0 9 2
28 9 4 12 9 13 9 1 9 2 3 9 0 0 9 16 4 13 13 0 9 7 13 9 15 15 4 0 2
36 3 2 2 16 9 1 12 4 0 9 0 9 2 9 4 13 2 7 9 9 0 0 9 0 4 0 2 2 13 9 11 11 1 9 11 2
27 0 9 7 9 9 9 11 9 1 0 7 0 9 2 11 2 11 11 13 16 4 0 9 9 15 9 2
36 2 1 0 2 9 4 13 15 9 1 0 9 1 0 9 2 15 13 16 14 13 13 16 15 15 0 9 13 1 0 9 2 2 13 4 2
37 11 4 13 16 13 9 15 4 2 0 0 9 1 9 2 14 0 2 3 0 2 14 0 3 0 2 14 0 3 0 7 14 0 3 0 2 2
25 1 11 2 0 11 13 13 0 9 1 0 9 7 15 9 2 15 15 3 13 1 9 0 9 2
42 2 13 16 4 15 9 3 4 0 9 15 13 0 9 2 9 11 13 13 2 0 9 2 1 0 2 0 7 0 9 2 15 15 3 13 16 9 2 2 13 11 2
34 9 9 15 9 3 13 9 9 16 13 9 11 2 0 9 1 0 9 2 11 2 7 0 9 2 15 4 9 13 9 1 15 9 2
47 1 9 1 9 11 1 12 9 2 15 4 13 0 9 2 11 13 16 15 0 9 1 11 13 9 9 0 7 0 0 9 2 1 9 9 16 15 13 0 9 0 9 0 0 0 9 2
28 16 15 9 3 4 13 9 9 9 2 13 11 2 13 4 15 9 9 0 9 1 9 15 15 13 1 11 2
28 9 13 16 4 0 0 9 13 4 9 9 9 0 9 15 4 13 9 2 3 9 9 9 0 9 7 9 2
4 9 9 1 9
16 9 9 1 0 11 1 9 9 2 9 7 9 1 12 9 2
18 11 11 2 0 0 9 7 9 13 4 1 12 9 9 1 0 9 2
29 12 1 9 0 9 2 12 1 0 9 15 15 13 1 9 1 12 9 2 11 4 0 9 4 0 9 1 11 2
12 1 12 1 12 9 4 4 9 1 0 9 2
18 0 9 9 11 11 0 1 11 1 15 9 0 4 12 9 1 11 2
20 11 15 13 7 13 1 11 13 4 9 1 0 9 1 11 7 11 0 9 2
15 1 0 0 9 11 0 4 12 9 12 0 0 9 11 2
13 0 9 13 1 12 9 2 0 9 7 0 9 2
10 1 9 9 3 15 13 12 0 9 2
13 1 11 1 11 0 4 12 9 12 9 0 9 2
32 1 9 15 4 13 9 9 0 4 9 9 1 11 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 7 8 11 2
13 1 11 1 11 7 11 0 4 12 0 0 9 2
15 11 13 1 9 9 9 3 4 0 1 0 9 1 11 2
11 1 0 9 13 4 12 9 1 12 9 2
24 11 1 9 2 0 9 11 1 9 0 11 2 0 4 1 12 1 12 9 1 11 1 11 2
34 1 9 9 15 4 3 13 11 9 9 7 0 9 11 11 13 4 0 0 9 2 9 7 9 1 11 2 11 7 11 7 11 11 2
22 0 0 0 0 0 0 9 11 13 4 12 7 12 9 9 1 9 11 11 1 11 2
11 1 9 4 4 9 0 0 7 0 9 2
8 9 9 3 3 0 9 1 11
22 9 9 11 1 11 11 11 13 4 9 1 0 9 1 9 1 9 9 1 15 9 2
31 9 9 1 11 13 0 9 1 9 11 2 13 4 9 9 15 9 1 15 9 1 9 15 4 0 0 9 11 1 11 2
24 1 0 9 2 9 9 13 1 0 9 1 9 7 0 9 2 15 13 0 9 15 9 13 2
30 2 9 1 15 15 9 9 13 1 9 9 7 9 9 1 9 1 9 9 0 9 13 0 9 2 2 13 4 11 2
15 15 4 3 13 1 9 1 15 15 15 0 9 13 13 2
50 2 0 9 1 9 1 9 0 9 2 3 9 9 9 2 7 9 0 9 2 7 9 16 15 4 9 9 1 9 1 9 2 3 13 9 9 2 11 2 2 15 4 13 1 9 13 15 9 2 2
20 0 9 1 9 9 0 9 3 4 13 1 0 9 9 1 9 9 7 9 2
36 0 9 1 0 9 13 4 1 12 9 1 9 9 7 9 15 9 1 0 13 1 9 0 9 7 9 2 16 7 1 9 9 1 9 2 2
35 11 11 2 15 13 15 9 2 13 16 4 15 9 9 0 9 9 1 9 9 2 9 2 15 1 9 13 3 13 15 9 1 0 9 2
20 0 9 8 8 8 7 9 8 8 2 9 11 11 2 15 13 9 15 9 2
28 9 11 11 13 4 11 2 0 7 0 9 1 9 0 9 9 2 1 2 0 9 0 1 9 15 9 2 2
24 11 13 16 4 9 9 2 9 9 1 9 2 1 9 16 4 13 13 1 9 1 9 2 2
25 9 15 4 11 13 1 9 9 4 0 1 0 9 0 9 7 9 1 15 15 11 3 13 13 2
17 0 9 9 11 11 7 9 11 11 3 4 13 9 1 15 9 2
25 1 9 2 9 0 9 11 8 0 4 0 9 1 0 9 7 4 0 13 12 9 9 0 9 2
21 1 0 9 2 9 1 9 0 0 9 11 8 13 0 9 16 2 0 9 2 2
18 1 9 15 9 0 4 16 4 1 11 13 0 9 2 7 14 9 2
25 11 11 2 0 7 0 9 9 11 2 13 16 15 3 13 0 9 1 9 2 9 7 9 9 2
7 9 11 11 13 9 9 9
31 3 9 1 9 9 1 0 9 9 1 11 1 9 9 11 2 9 9 13 4 16 4 1 0 9 9 13 13 12 9 2
15 2 0 4 0 11 2 2 13 4 0 0 9 11 11 2
11 2 13 4 3 1 12 7 0 9 2 2
38 11 4 13 3 13 9 1 11 12 9 2 13 4 1 9 2 12 9 2 9 11 11 2 3 16 9 9 1 9 9 1 9 11 9 11 4 13 2
31 9 4 0 3 9 1 9 9 1 0 9 9 1 11 1 9 9 1 9 9 11 2 15 4 0 0 9 11 7 11 2
44 3 2 1 0 9 1 9 9 1 9 2 9 12 9 15 4 13 9 2 11 2 11 2 11 2 11 2 11 7 0 9 2 1 9 4 13 13 13 14 9 13 1 9 2
29 2 3 3 13 9 1 9 9 7 15 9 13 16 4 9 15 9 0 9 2 2 13 4 0 9 11 11 11 2
11 2 13 3 13 16 4 13 9 1 9 2
42 3 2 13 16 4 3 0 13 16 9 4 13 1 9 7 13 13 15 9 3 3 16 4 9 9 2 1 9 2 7 4 3 3 16 4 15 0 9 0 9 2 2
20 11 4 13 0 0 9 15 4 1 0 3 9 13 0 9 7 15 0 9 2
29 9 4 13 16 15 0 9 3 13 9 15 4 13 0 9 11 11 11 2 1 15 4 11 13 4 0 0 9 2
19 3 16 13 13 15 9 9 1 9 2 11 4 3 13 9 16 0 9 2
13 11 4 13 16 4 13 15 9 15 4 0 11 2
26 1 11 2 0 9 0 4 12 9 9 1 11 7 11 2 1 15 4 9 9 13 9 1 15 9 2
19 9 15 3 3 11 13 0 9 0 0 9 15 4 13 9 1 0 9 2
19 3 3 9 11 2 11 4 8 8 1 9 11 1 9 9 12 2 12 2
50 9 0 9 11 11 9 13 4 3 15 9 16 4 2 7 15 11 13 13 9 2 0 9 9 2 15 4 9 11 2 11 2 11 2 11 2 11 7 0 9 2 3 1 15 13 9 9 9 2 2
22 0 4 16 4 15 9 9 9 13 1 9 9 2 2 13 4 11 0 9 1 9 2
29 2 13 13 3 7 13 9 1 12 9 2 2 2 1 9 9 11 2 7 4 1 9 9 13 15 15 13 2 2
8 9 9 13 15 13 1 9 2
37 1 9 2 0 0 9 11 11 2 15 4 9 13 0 9 0 9 2 3 4 13 1 9 16 4 11 1 9 13 0 2 1 12 7 0 9 2
15 2 0 4 0 11 2 2 13 4 9 1 9 1 11 2
11 2 13 4 3 1 12 7 0 9 2 2
23 11 15 13 13 1 11 1 11 1 9 2 1 0 0 9 0 11 1 9 1 9 9 2
15 0 9 1 9 13 16 13 13 0 9 1 3 0 9 2
20 2 3 4 4 13 9 1 9 9 11 2 2 13 4 0 9 11 11 11 2
16 2 16 15 9 14 13 2 11 4 13 13 9 15 9 2 2
39 11 11 2 9 0 9 11 7 9 0 0 9 2 13 4 15 9 1 9 2 3 16 4 9 11 13 2 13 15 9 1 9 11 9 9 1 11 2 2
9 9 7 9 2 11 9 9 1 11
13 0 9 1 11 7 0 9 4 4 0 1 11 2
25 3 1 9 1 9 2 0 9 11 4 4 9 9 1 0 9 2 7 1 11 0 9 0 9 2
12 11 4 4 9 0 9 1 11 7 0 9 2
33 11 2 1 11 2 4 4 12 7 12 9 9 0 0 9 1 11 7 0 9 2 13 4 1 9 2 12 9 2 0 9 11 2
17 9 4 13 0 9 2 9 2 9 2 16 7 0 7 0 9 2
13 9 9 4 4 0 1 0 9 2 9 7 9 2
26 0 9 13 4 9 11 1 9 9 1 9 9 11 2 13 4 1 9 2 12 9 2 0 9 9 2
22 1 9 2 9 11 1 9 11 11 13 4 9 9 1 9 9 11 1 9 0 9 2
18 0 9 11 0 4 1 9 9 9 11 1 9 1 12 9 1 9 2
26 0 9 11 4 4 1 12 9 1 9 2 12 9 2 9 0 9 1 0 9 2 13 4 9 11 2
20 9 1 0 9 13 4 9 2 0 9 1 15 9 15 4 3 0 1 11 2
18 1 9 1 15 15 13 4 4 9 9 7 9 11 0 1 0 9 2
12 9 0 9 0 4 1 9 0 9 1 11 2
14 1 9 9 2 1 9 4 12 1 0 9 1 11 2
16 9 13 16 4 9 4 0 1 12 9 7 0 1 12 9 2
5 9 4 3 0 2
13 11 1 11 4 4 12 9 9 0 9 0 9 2
12 0 4 4 0 9 15 13 1 0 0 9 2
20 9 0 9 0 9 1 11 13 4 0 9 1 0 0 9 1 0 0 9 2
15 11 11 13 4 0 9 15 9 9 0 9 9 0 9 2
17 15 4 3 13 11 1 0 9 1 0 9 15 15 13 1 11 2
9 0 9 13 1 9 1 9 1 11
18 9 9 1 9 9 0 9 1 9 1 15 13 0 9 13 4 9 2
12 0 9 0 9 11 13 4 0 9 1 9 2
23 1 15 9 1 12 9 2 9 4 13 9 1 9 9 0 9 1 9 0 9 1 0 2
14 9 0 0 9 15 9 3 4 13 9 1 9 9 2
17 9 0 9 11 11 7 9 11 11 13 4 16 4 9 3 0 2
21 2 16 9 0 9 11 14 13 13 15 9 7 3 13 9 2 2 13 4 11 2
16 9 1 15 9 0 4 0 9 1 15 15 4 9 3 13 2
37 1 0 9 9 0 4 16 9 1 15 13 0 9 4 3 13 13 15 9 1 7 1 0 9 2 0 9 7 1 9 1 0 7 0 0 9 2
18 3 2 1 0 9 0 12 9 2 9 4 13 16 15 4 3 0 2
36 9 4 13 16 4 13 3 9 15 4 0 9 0 9 1 9 1 0 0 9 1 9 7 13 9 16 13 13 14 15 0 9 13 7 14 2
24 1 9 3 4 0 16 4 0 13 9 9 3 1 9 3 9 13 0 9 2 3 0 9 2
11 1 9 2 13 9 16 4 9 3 13 2
27 0 0 0 9 2 0 9 1 9 2 11 2 2 13 4 16 4 13 9 7 4 13 15 9 9 9 2
18 3 2 0 9 11 2 9 0 9 2 13 16 11 7 11 13 9 2
12 2 9 0 9 13 4 0 9 11 7 11 2
22 15 4 15 9 1 9 9 1 11 7 9 9 7 9 0 9 2 2 13 4 9 2
15 1 9 12 9 2 9 14 4 13 13 1 9 9 9 2
12 2 13 0 9 0 9 15 3 3 4 0 2
15 9 4 13 13 7 13 1 9 2 2 13 4 11 11 2
11 0 9 2 0 9 13 4 9 1 0 11
17 11 13 13 12 9 9 1 0 9 2 3 1 11 7 1 11 2
14 3 15 9 2 0 9 13 4 3 12 9 1 11 2
14 9 4 4 0 1 9 0 9 1 11 7 1 11 2
20 0 9 9 7 9 2 11 2 13 13 12 9 9 1 9 9 1 0 11 2
21 1 9 4 13 1 12 7 12 9 2 3 1 9 0 9 1 11 7 1 11 2
33 0 9 13 4 0 9 0 9 1 9 9 1 9 12 9 9 7 12 9 9 9 0 9 2 1 9 0 9 9 9 1 11 2
10 0 9 9 0 4 1 12 9 9 2
49 9 9 1 11 7 11 13 4 13 12 9 9 1 9 15 9 7 3 15 13 1 12 9 9 1 12 9 2 13 4 0 9 11 11 11 1 11 0 9 0 1 9 2 12 9 2 1 11 2
17 9 9 1 0 12 9 12 9 0 4 1 12 9 1 0 9 2
20 0 9 9 1 9 2 11 2 13 9 9 9 1 9 9 1 11 1 11 2
20 11 3 13 9 1 9 9 7 9 1 11 2 15 4 13 12 9 0 9 2
36 11 4 3 13 13 9 1 0 9 2 1 9 3 4 0 2 1 0 9 0 0 9 2 13 4 1 9 2 12 9 2 9 9 11 11 2
28 9 9 1 9 1 11 7 11 2 11 2 13 4 4 12 9 9 1 9 2 13 9 9 1 9 9 11 2
13 0 9 9 0 4 1 12 9 9 7 12 9 2
13 1 9 2 0 0 9 1 9 13 12 9 9 2
7 11 9 0 1 9 7 9
28 0 0 9 11 2 0 1 11 2 13 4 12 9 7 0 9 2 3 11 11 2 11 2 11 11 7 11 2
26 9 2 3 0 1 9 0 0 9 1 0 9 2 3 4 13 16 9 1 9 9 1 0 0 9 2
31 3 2 15 4 9 0 9 2 9 1 9 9 1 11 7 9 0 9 1 0 9 2 0 1 9 0 9 7 0 9 2
47 0 0 9 0 11 2 0 1 12 1 12 9 1 0 0 9 11 2 13 4 3 1 12 9 2 1 9 9 7 1 12 0 9 1 0 9 2 3 7 0 0 9 1 11 7 11 2
36 0 9 4 13 9 9 2 12 9 15 4 13 1 9 3 2 8 8 8 8 8 8 2 2 0 4 3 3 13 2 1 11 11 1 11 2
41 1 0 4 9 1 9 4 7 8 8 2 11 2 11 11 2 11 11 2 11 2 11 2 11 2 7 11 1 11 11 2 11 8 11 7 0 9 11 11 11 2
51 9 1 0 9 2 16 7 1 11 11 2 11 2 11 7 0 9 11 2 13 4 1 0 11 16 4 13 0 9 0 9 2 3 8 9 2 9 2 9 2 9 2 8 8 2 9 2 9 7 9 2
8 9 9 13 15 1 0 9 2
8 15 4 3 4 0 11 9 2
12 0 4 2 0 2 11 9 0 1 9 12 2
11 13 4 12 9 7 13 9 9 1 11 2
19 0 4 0 11 9 0 12 1 11 2 7 13 15 4 3 1 12 9 2
23 1 3 4 11 13 3 0 9 1 8 11 2 11 7 11 11 2 16 7 3 0 11 2
36 1 9 1 9 9 2 4 3 13 9 12 1 0 9 1 11 11 2 15 4 11 9 13 16 2 0 1 11 2 7 1 3 1 9 2 2
13 0 9 15 9 13 1 9 15 4 11 3 13 2
33 4 16 4 4 9 1 9 1 9 7 1 9 2 7 7 9 9 9 9 1 9 11 2 9 4 3 13 0 9 1 0 9 2
24 9 4 13 9 1 0 9 2 7 1 11 11 2 11 7 11 2 16 7 1 0 9 11 2
16 3 2 15 4 9 9 0 1 0 9 0 9 7 0 9 2
35 9 4 13 9 9 1 9 9 1 11 2 1 15 4 13 9 11 11 2 8 8 8 8 8 2 2 3 4 13 9 2 7 0 9 2
31 2 12 9 3 2 13 15 9 7 9 15 9 16 15 11 2 11 2 11 2 11 2 11 2 11 7 0 11 4 13 2
8 3 2 2 2 13 4 9 2
25 16 9 4 13 4 0 1 15 4 0 9 13 1 0 9 1 9 16 1 9 4 0 0 9 2
45 16 16 15 4 4 0 2 0 0 9 2 15 4 1 9 1 9 0 11 2 13 4 9 9 9 9 9 11 11 16 2 11 4 4 0 9 16 15 13 13 9 9 11 2 2
13 8 8 4 4 12 1 9 15 4 13 1 11 2
10 1 9 1 9 9 13 4 9 9 2
26 0 4 9 0 9 1 0 9 9 9 1 15 4 13 2 14 13 13 2 2 9 1 9 1 11 2
33 3 4 4 9 3 1 9 1 11 2 3 1 9 1 11 1 0 9 9 0 1 11 2 11 7 11 2 7 11 7 0 0 2
24 4 4 9 1 12 9 1 9 7 14 13 16 15 15 3 13 4 0 2 2 13 4 11 2
17 9 4 3 13 16 4 0 13 9 9 7 13 9 1 0 9 2
34 1 9 9 1 0 9 2 9 0 11 11 11 2 9 0 0 9 2 13 15 1 11 1 0 9 9 2 3 15 7 3 1 9 2
15 0 9 1 0 11 3 4 13 9 2 16 7 0 9 2
19 13 9 16 4 0 9 1 0 9 13 7 9 1 9 9 1 0 9 2
9 0 9 2 0 9 0 9 13 11
21 9 0 9 0 9 11 11 13 15 1 9 1 9 11 11 11 7 9 11 11 2
18 3 1 0 9 2 0 9 11 11 11 13 1 11 1 9 9 9 2
41 9 0 9 0 9 11 11 13 4 0 9 11 11 1 9 1 9 2 12 9 2 1 11 16 4 15 9 2 13 1 9 9 11 1 9 1 0 9 11 2 2
40 1 15 2 11 4 13 9 9 11 1 9 12 0 9 1 11 16 4 13 9 11 7 13 16 16 4 0 9 13 1 9 11 2 16 15 4 13 1 11 2
21 11 15 3 13 1 9 11 11 11 2 9 9 11 11 7 9 9 11 11 11 2
38 11 13 9 9 0 9 7 9 0 1 0 9 2 13 4 1 9 2 12 9 2 0 9 0 9 11 11 2 1 9 1 0 9 11 11 1 11 2
22 9 9 13 4 0 9 1 9 12 9 2 3 15 9 1 0 9 1 9 12 9 2
17 0 9 11 11 13 4 1 11 1 9 2 12 9 2 7 9 2
20 4 4 0 9 0 0 9 2 3 9 1 9 9 1 9 9 11 2 11 2
25 0 9 11 11 11 13 4 1 9 2 12 9 2 1 0 9 11 1 9 9 11 11 11 11 2
16 11 4 13 1 0 9 9 9 15 15 13 1 9 7 9 2
17 13 15 9 1 12 9 1 12 9 2 3 0 9 11 11 11 2
25 0 9 0 9 11 11 13 4 1 9 2 12 9 2 1 11 3 4 13 1 0 9 11 11 2
22 13 4 15 16 4 0 9 9 1 9 7 9 1 11 7 11 4 1 0 9 0 2
21 11 4 3 13 16 9 9 13 1 0 9 11 1 9 11 1 0 9 1 11 2
28 9 9 9 0 2 11 2 11 11 7 15 0 9 11 11 13 4 1 9 2 12 9 2 9 1 0 9 2
21 9 4 0 9 1 12 9 2 3 9 2 9 0 9 2 0 9 7 0 9 2
14 0 9 11 1 11 2 9 0 9 1 11 7 11 11
18 1 12 1 12 9 2 11 4 16 9 0 9 11 4 9 9 11 2
44 0 9 11 11 4 2 3 1 9 9 9 11 2 13 16 9 1 9 0 9 9 1 11 13 2 0 9 1 15 3 9 13 16 11 7 11 11 13 9 1 0 9 2 2
26 9 11 11 11 13 4 0 9 1 11 7 11 11 2 3 16 4 9 13 0 9 1 0 12 9 2
24 13 4 16 15 11 3 13 1 9 2 9 9 9 2 0 9 2 7 13 9 11 1 9 2
14 9 1 0 9 11 13 12 9 1 0 9 1 11 2
19 11 4 1 11 13 15 12 0 9 0 9 15 12 9 9 7 0 9 2
32 0 9 11 2 0 1 11 1 12 1 12 9 2 4 4 0 0 9 15 15 1 0 12 9 13 1 9 11 7 11 11 2
24 3 12 9 2 3 12 0 9 7 9 0 0 9 7 0 9 2 13 15 1 15 0 9 2
21 9 4 13 0 9 2 0 9 9 0 9 9 9 2 7 9 9 9 9 9 2
10 1 15 2 0 4 7 12 0 9 2
40 0 9 11 11 4 1 9 1 9 11 11 11 13 16 4 9 0 0 9 1 11 9 0 9 9 1 11 2 7 13 9 0 9 16 13 1 15 0 9 2
38 3 4 13 16 9 11 16 13 9 1 11 13 9 0 9 2 15 4 1 0 9 1 9 1 0 9 9 1 9 1 9 7 9 1 11 0 9 2
26 11 4 1 15 9 13 1 0 9 1 11 7 11 11 2 3 16 4 9 3 13 1 0 12 9 2
26 13 4 16 15 11 3 13 1 9 2 0 9 9 2 3 0 9 2 7 4 13 9 11 1 9 2
8 2 9 11 4 3 0 9 2
13 11 7 11 11 0 4 9 1 9 1 1 9 2
37 1 9 15 13 16 13 0 9 1 15 9 7 15 9 9 2 9 0 0 9 7 9 1 9 9 0 15 2 2 13 4 11 3 15 0 9 2
23 11 7 0 0 9 4 1 9 9 13 16 4 1 11 13 0 12 11 2 9 15 9 2
40 11 3 13 12 1 0 9 1 11 7 11 11 2 0 4 3 12 11 2 9 1 12 9 2 7 0 4 7 3 12 9 9 1 9 9 9 3 0 11 2
17 11 7 9 3 4 13 0 9 1 9 0 1 9 9 1 11 2
25 9 4 4 0 12 11 2 9 1 9 9 2 7 3 12 11 2 9 1 9 0 7 0 9 2
13 0 9 15 9 13 7 0 12 12 9 0 9 2
27 1 9 1 15 2 9 0 9 11 11 13 4 12 9 16 0 9 13 16 4 0 9 0 1 0 9 2
13 2 3 4 3 0 7 0 9 1 0 9 2 2
34 1 0 9 0 0 9 7 9 3 9 0 4 9 16 4 1 0 9 13 4 0 9 2 3 1 9 1 0 9 2 9 1 11 2
11 0 9 13 13 1 9 9 1 0 9 2
22 2 4 4 9 1 0 0 0 9 2 3 3 1 0 7 0 9 2 7 0 9 2
35 13 16 4 15 1 15 9 0 9 13 0 9 2 1 9 16 4 1 9 0 16 15 13 9 3 2 2 13 4 0 9 9 11 11 2
32 1 9 2 9 11 11 11 11 2 13 4 16 0 11 13 1 9 0 9 2 15 1 0 13 7 9 11 1 9 1 11 2
10 11 4 13 0 9 16 15 0 9 2
25 9 11 2 0 4 9 1 15 16 9 13 1 11 7 11 11 1 0 9 0 9 2 13 4 2
28 2 11 7 11 11 4 15 9 13 16 15 13 0 9 2 2 13 4 11 9 9 9 2 3 0 3 0 2
17 13 4 16 4 9 0 1 11 7 11 11 9 3 13 9 9 2
33 0 9 9 9 0 1 9 7 9 1 11 2 7 15 4 11 13 12 9 2 13 4 2 3 0 9 9 2 2 13 4 11 2
13 2 9 15 0 9 1 11 13 9 9 0 11 2
48 15 4 9 2 13 1 0 0 9 2 7 1 0 9 7 9 2 3 0 0 9 1 15 13 9 15 4 13 0 9 9 2 15 15 13 13 1 3 0 9 1 15 9 2 2 13 4 2
30 11 4 13 16 4 11 13 1 9 0 0 9 2 9 9 1 0 9 7 9 0 9 9 0 7 0 9 0 11 2
17 15 15 4 3 13 1 11 13 4 3 7 13 16 15 9 14 13
23 9 8 8 11 11 11 1 0 7 0 9 15 9 13 13 9 11 7 11 2 11 2 2
21 0 9 16 4 15 0 9 13 13 1 11 7 11 2 11 2 4 13 0 9 2
28 9 4 13 13 1 0 0 9 7 0 9 2 3 0 0 7 0 9 2 1 15 0 9 1 0 9 9 2
28 15 1 9 1 15 13 0 9 13 0 0 9 7 3 4 3 3 2 16 14 7 3 2 13 3 0 9 2
25 0 9 2 0 16 4 15 13 9 7 13 16 9 1 9 2 13 4 13 0 9 7 0 9 2
16 9 4 0 0 9 11 2 7 4 0 9 15 9 1 9 2
13 15 4 11 7 11 0 0 9 1 0 9 11 2
15 3 2 0 9 3 4 4 9 9 16 9 1 0 9 2
33 3 12 9 1 9 9 2 0 9 1 15 15 13 0 9 7 3 15 13 1 12 0 9 2 13 14 7 4 4 0 9 11 2
8 2 13 15 13 12 1 0 2
5 3 4 13 9 2
18 15 4 15 13 13 7 13 11 2 16 4 9 1 9 13 0 11 2
10 13 4 9 1 11 15 4 0 13 2
24 15 3 4 13 7 9 1 15 9 15 4 13 1 11 2 2 13 0 9 9 11 11 11 2
44 16 0 9 15 4 3 1 9 9 9 13 13 9 11 16 0 9 2 0 9 0 4 9 0 9 2 11 2 2 9 15 13 0 9 0 9 7 13 9 0 0 0 9 2
18 11 4 1 0 9 13 0 9 7 1 9 4 13 3 16 0 9 2
21 3 4 13 9 0 9 15 9 2 15 4 15 13 13 16 4 15 9 13 3 2
9 0 9 13 4 1 9 12 9 2
23 1 9 1 11 11 4 0 9 1 9 9 7 0 9 7 9 9 15 13 9 0 9 2
7 15 9 13 4 9 9 2
32 0 0 9 0 16 9 0 9 13 4 9 0 0 9 1 9 2 0 0 9 2 0 9 2 7 15 4 0 2 0 9 2
15 11 4 3 13 3 0 9 1 9 9 2 3 9 9 2
25 0 9 13 15 13 3 2 1 0 9 3 9 16 4 0 9 13 0 9 1 9 9 0 9 2
17 3 4 13 9 1 9 1 15 9 13 0 9 1 0 0 9 2
15 11 4 13 0 9 9 2 3 9 1 0 9 0 9 2
18 0 9 15 9 4 9 0 0 9 9 11 2 15 4 11 13 0 2
19 1 9 1 9 15 1 0 9 2 15 13 0 9 1 15 4 13 13 2
37 9 3 2 1 15 9 0 9 2 3 4 4 9 1 0 15 15 4 0 1 3 2 7 16 15 4 13 0 9 11 11 2 9 1 9 9 2
17 13 3 9 15 15 13 13 1 9 1 11 2 7 12 4 0 2
27 16 0 2 9 9 9 3 13 0 7 0 7 15 15 13 2 7 15 4 0 16 1 9 4 0 9 2
34 16 0 2 9 0 0 9 13 4 4 3 0 16 4 13 13 0 9 1 0 9 2 7 1 15 9 13 4 4 0 1 0 9 2
29 7 16 0 2 9 0 1 0 9 13 4 0 7 13 4 0 0 0 9 2 16 15 0 9 13 13 0 9 2
9 11 13 1 9 9 1 9 9 11
26 0 0 9 13 4 9 15 15 0 9 11 11 11 13 1 0 9 15 9 0 1 9 0 9 11 2
17 1 9 15 3 13 11 1 9 9 11 7 9 15 9 1 9 2
32 0 0 9 2 11 2 13 4 1 9 2 12 9 2 1 9 9 11 1 9 9 9 11 7 1 0 9 11 1 15 9 2
36 1 9 15 4 13 1 15 0 9 1 11 2 11 4 13 0 9 11 11 11 1 2 9 15 9 1 9 9 0 1 0 9 1 11 2 2
33 9 2 15 4 13 9 0 9 0 11 0 9 2 11 11 2 3 15 13 11 2 1 0 9 1 0 9 1 9 9 11 2 2
35 11 13 12 0 7 0 9 1 12 9 7 3 1 0 9 13 12 9 1 0 9 15 13 12 9 2 15 4 13 0 0 9 1 9 2
37 0 0 9 1 9 9 11 0 4 9 1 9 12 9 2 3 4 0 11 0 9 13 0 9 1 9 0 9 2 16 15 4 9 0 11 13 2
21 1 9 4 3 3 0 9 0 9 1 9 0 11 13 1 11 12 9 0 9 2
8 0 9 0 9 13 3 11 2
33 11 4 0 1 0 0 9 12 9 15 4 13 1 0 9 0 11 15 4 13 11 2 7 15 4 1 9 13 9 9 1 11 2
28 11 4 1 15 9 13 11 16 2 13 1 0 9 15 9 3 0 9 11 7 1 9 1 0 0 9 2 2
30 11 15 3 13 16 1 9 13 7 13 9 15 15 15 0 9 1 11 13 1 0 12 9 9 2 7 13 9 11 2
14 11 4 13 16 9 0 9 4 0 9 9 0 11 2
43 0 0 9 2 3 9 11 11 11 2 1 3 9 3 4 13 16 4 0 9 7 0 9 1 9 13 0 1 9 7 9 0 11 14 16 9 0 11 4 13 1 9 2
7 9 1 9 0 9 1 11
21 9 9 1 9 1 0 9 1 9 0 9 13 4 9 9 1 2 0 9 2 2
17 0 9 11 11 13 4 16 4 9 9 0 9 1 9 9 9 2
26 9 9 15 4 13 0 0 9 2 11 2 2 1 9 1 9 11 11 2 13 4 0 9 0 9 2
23 9 0 9 13 4 12 9 2 3 4 9 9 13 9 0 0 0 9 0 15 1 9 2
20 1 15 9 0 4 0 0 9 1 9 9 9 9 9 7 15 3 0 9 2
18 3 2 0 9 13 15 12 9 2 3 4 11 4 0 13 1 9 2
20 3 3 15 13 1 9 2 13 9 2 11 13 3 12 9 2 0 9 2 2
21 11 4 13 15 9 3 16 3 13 0 9 11 16 4 13 1 0 9 0 9 2
9 2 4 0 16 9 13 0 9 2
18 13 4 16 4 1 0 9 2 0 7 1 9 2 2 13 4 11 2
15 2 12 9 15 4 13 1 0 0 9 13 4 1 12 2
9 13 4 9 3 15 0 9 9 2
7 3 13 0 9 9 2 2
10 0 9 11 11 14 13 15 1 15 2
13 2 2 9 2 2 2 2 4 9 0 9 9 2
17 0 9 13 15 3 1 0 9 3 4 1 9 9 9 7 9 2
13 15 9 1 9 13 9 9 7 9 15 15 13 2
13 13 15 16 4 9 15 13 9 1 9 7 9 2
15 15 4 15 15 4 0 1 0 9 2 2 13 4 11 2
16 9 0 4 4 0 9 2 15 3 13 0 9 1 0 9 2
9 0 4 15 13 9 1 0 9 2
16 2 1 9 9 9 0 4 16 9 2 9 2 13 15 9 2
41 3 0 9 2 9 7 9 3 15 13 1 9 2 4 16 15 13 1 9 15 13 0 9 7 1 15 1 9 0 9 2 2 13 4 9 0 0 9 11 11 2
22 1 15 9 2 0 4 0 9 7 0 0 9 16 4 15 13 9 9 1 0 9 2
12 9 4 16 15 13 0 9 9 2 13 11 2
5 9 13 9 1 11
22 11 13 1 0 9 0 9 16 9 0 9 0 11 2 7 14 13 15 0 9 9 2
28 16 15 0 9 13 1 9 7 9 9 13 2 9 4 3 13 1 9 1 9 1 3 12 0 9 2 9 2
8 0 9 13 0 9 9 11 2
19 1 0 0 9 2 9 0 9 12 4 1 0 9 0 9 9 1 9 2
46 9 13 16 4 14 16 9 14 13 9 2 9 13 12 9 2 3 15 13 1 9 15 9 2 7 3 4 0 16 4 13 1 12 9 2 15 4 1 9 9 9 1 0 9 9 2
22 11 13 9 0 9 1 0 9 1 12 9 9 2 15 4 15 13 12 1 9 9 2
27 13 15 16 15 9 9 1 9 4 13 3 3 4 15 13 1 12 9 2 15 4 4 0 0 0 9 2
14 11 13 13 15 1 9 1 0 9 9 2 0 9 2
10 3 2 0 9 1 11 3 4 0 2
19 3 1 9 12 9 2 1 3 9 9 2 9 4 13 9 1 9 9 2
31 13 15 16 4 0 9 4 3 0 2 16 7 15 0 9 1 12 9 2 1 15 15 7 1 12 9 14 13 0 9 2
20 11 4 0 9 13 0 9 2 7 13 1 13 13 14 15 13 4 15 9 2
25 9 13 16 4 0 9 15 13 9 2 7 9 9 7 9 3 0 2 16 4 15 15 3 13 2
24 9 11 0 4 0 9 9 15 15 13 0 0 9 2 3 0 9 2 0 9 7 0 9 2
17 3 2 0 9 0 1 9 2 3 1 0 9 2 13 0 9 2
14 0 0 9 3 13 9 2 13 9 0 9 1 11 2
24 2 2 9 2 3 13 9 3 9 9 2 9 2 9 9 9 2 7 3 9 9 15 0 2
20 15 9 3 3 13 9 9 0 9 2 2 13 11 11 2 15 13 9 9 2
20 0 9 2 11 11 2 13 1 9 9 2 15 9 13 0 9 9 0 9 2
21 12 9 2 12 9 0 0 9 11 2 1 9 4 12 9 2 0 0 9 11 2
22 1 0 9 2 13 3 12 0 9 2 0 11 2 0 9 11 11 7 0 8 8 2
22 0 9 0 9 1 9 4 0 9 2 1 15 4 0 9 9 2 0 9 1 11 2
23 0 9 11 1 11 2 11 11 2 3 13 16 9 13 13 0 9 1 9 1 0 9 2
17 9 1 0 9 7 0 3 4 0 9 1 15 9 2 13 11 2
26 9 9 11 11 7 9 9 11 11 11 3 4 12 9 13 9 2 7 4 0 0 9 1 15 9 2
17 14 16 9 14 13 15 9 9 2 13 9 2 9 4 13 0 2
6 11 11 0 1 9 9
36 11 2 11 2 9 4 13 13 9 1 9 11 11 11 11 2 16 4 15 13 15 9 2 13 4 1 9 2 12 9 2 9 9 11 11 2
25 9 4 0 2 1 9 7 0 9 1 9 9 2 1 15 4 0 9 9 1 12 1 12 9 2
8 0 9 13 4 13 12 9 2
10 9 3 13 16 15 11 13 1 9 2
14 0 0 9 1 9 4 1 12 9 7 13 1 11 2
21 3 4 4 0 1 9 15 9 1 0 9 9 1 0 9 9 15 9 12 9 2
6 11 13 1 9 1 11
21 16 4 11 3 1 0 9 1 11 2 1 9 4 1 9 0 9 1 15 9 2
31 1 9 2 12 9 2 2 9 1 12 0 9 13 4 1 9 1 9 1 11 2 3 16 15 0 9 3 13 1 9 2
26 2 11 4 1 1 9 13 16 2 3 4 13 0 9 11 2 2 15 13 16 15 3 4 13 11 2
35 2 0 11 2 9 4 11 15 4 13 15 9 7 13 15 0 7 0 9 1 15 2 2 13 4 9 1 9 15 4 13 9 11 11 2
29 3 0 9 2 15 9 13 1 0 0 9 11 2 4 3 13 7 3 15 3 13 16 4 15 13 9 1 11 2
30 1 15 9 2 0 9 1 9 11 4 9 9 1 0 11 12 9 1 15 4 13 2 3 15 13 2 3 12 9 2
28 15 9 13 4 16 4 0 15 9 0 1 0 9 9 1 9 1 9 9 0 9 9 11 12 9 1 11 2
31 1 9 15 13 16 11 2 13 9 15 4 11 3 13 1 9 9 1 9 2 2 16 0 9 4 4 0 1 15 9 2
12 9 13 16 15 9 9 11 13 9 1 11 2
24 9 1 0 9 7 9 13 4 12 9 12 9 9 9 15 13 16 4 12 9 9 1 9 2
9 3 15 12 9 13 1 15 9 2
17 9 9 11 11 2 3 2 13 16 4 3 16 15 11 13 11 2
60 2 3 4 16 15 14 13 9 1 11 16 9 1 9 11 1 11 2 7 4 3 3 16 16 13 13 9 0 9 1 11 2 13 13 0 0 9 2 2 13 4 11 0 9 8 2 3 16 14 13 0 9 1 11 16 4 15 13 11 2
30 3 2 0 0 9 11 11 2 3 9 0 0 0 9 2 13 4 16 4 9 11 11 13 9 11 2 15 0 9 2
13 11 4 3 13 9 11 1 9 11 16 0 9 2
12 0 9 11 4 7 3 1 11 7 13 9 2
14 11 4 13 9 0 9 9 1 9 1 9 12 9 2
20 0 9 11 11 11 11 13 4 1 9 12 9 16 9 13 16 11 13 9 2
17 1 9 12 9 2 11 4 13 0 9 1 9 15 4 13 9 2
6 3 1 9 1 11 11
11 11 13 9 2 7 9 2 9 1 9 2
14 9 9 13 4 11 0 9 2 7 1 9 7 9 2
12 3 2 1 0 4 9 4 7 0 7 0 2
23 3 1 0 1 0 11 2 9 11 11 13 4 1 0 9 1 9 3 4 13 0 9 2
8 15 4 13 3 15 11 13 2
13 2 13 4 16 4 13 0 9 9 2 0 9 2
22 1 0 9 11 4 13 0 9 15 4 4 0 15 1 11 2 2 13 15 11 11 2
23 16 4 0 9 13 9 1 2 0 9 2 0 4 13 16 4 9 1 9 9 1 11 2
6 3 4 0 13 3 2
32 11 4 13 1 9 16 15 9 13 2 7 15 9 13 4 1 9 0 9 1 12 7 12 9 2 15 4 0 16 0 9 2
21 3 2 0 11 13 3 16 3 2 13 11 2 12 2 9 9 7 0 9 9 2
15 15 9 2 11 11 2 4 4 9 11 1 9 15 9 2
27 2 9 9 13 4 0 9 3 2 2 13 15 2 3 0 9 1 9 1 9 2 12 1 0 1 11 2
20 2 4 4 0 9 2 4 4 9 2 4 4 3 3 9 7 1 0 9 2
18 0 4 4 3 2 3 0 2 7 13 15 16 4 15 13 9 2 2
11 0 9 13 4 2 3 2 1 0 9 2
22 11 11 4 4 0 0 9 7 13 4 1 0 0 9 15 4 13 9 1 0 9 2
13 11 4 1 9 13 9 15 4 13 12 9 9 2
14 9 2 0 11 11 2 13 4 9 1 11 16 9 2
19 9 9 2 13 4 15 2 13 4 9 7 13 0 9 7 13 9 9 2
5 15 15 4 13 2
22 11 11 2 0 9 9 9 7 0 9 2 12 9 13 4 9 13 9 1 15 9 2
16 1 9 4 14 11 3 0 2 3 15 13 7 13 0 9 2
16 2 0 9 2 0 7 0 2 3 4 0 13 1 9 2 2
24 1 11 11 2 9 9 9 2 0 11 3 13 16 3 3 3 13 1 9 7 0 9 9 2
25 2 12 9 3 0 9 4 1 9 2 1 9 16 4 9 13 1 12 0 9 2 2 13 4 2
40 2 2 0 2 9 3 3 4 1 9 0 2 16 15 7 3 13 2 16 1 0 9 2 16 15 9 14 13 13 2 16 4 15 3 3 4 13 4 2 2
14 9 1 9 2 13 11 2 13 4 1 9 0 9 2
45 2 16 15 15 9 13 2 3 16 15 9 13 3 0 9 1 9 11 11 2 7 4 0 16 4 15 15 3 13 2 15 11 13 4 13 16 13 4 3 0 2 2 13 11 2
9 9 2 2 0 9 2 9 1 11
15 16 15 9 3 9 3 13 2 9 0 9 13 0 9 2
17 11 15 13 1 2 0 2 1 2 3 0 2 9 1 0 9 2
41 0 9 1 9 9 0 9 7 0 9 1 12 9 13 4 9 9 3 9 2 13 4 0 9 1 9 9 8 8 1 15 0 9 0 1 9 2 12 9 2 2
30 2 15 4 0 0 9 9 0 9 1 3 0 9 2 9 9 1 9 2 15 4 15 9 0 12 9 7 12 9 2
51 9 0 9 13 4 0 9 1 12 1 12 7 13 15 0 9 1 12 9 2 13 15 1 9 7 13 16 4 13 1 9 0 9 1 12 9 1 11 2 0 11 2 1 0 9 7 1 0 0 9 2
47 2 9 4 0 7 13 1 9 1 0 7 0 9 2 9 15 4 3 13 9 2 0 2 9 7 0 4 0 9 0 9 7 0 9 2 2 13 4 11 11 2 9 15 9 1 9 2
21 2 16 9 4 0 2 0 0 9 13 4 0 2 0 1 0 9 7 0 2 2
18 8 8 13 15 0 9 9 0 9 7 0 9 1 9 1 12 9 2
27 16 4 13 9 2 8 8 13 0 9 2 0 9 7 9 9 16 7 9 9 2 9 9 7 9 9 2
39 1 9 9 15 9 1 9 1 12 9 2 1 15 16 12 13 0 2 7 12 0 2 15 9 7 9 0 4 1 9 0 9 0 2 3 0 7 0 2
34 3 0 9 13 15 1 0 9 1 12 1 12 9 2 7 11 2 11 2 11 2 11 11 7 11 13 15 1 15 15 4 13 9 2
19 2 12 9 0 11 13 4 1 9 1 12 9 2 2 13 15 1 9 2
44 2 1 0 9 13 4 1 11 2 15 4 13 1 9 0 1 9 3 0 9 2 1 15 4 0 9 1 15 4 0 16 4 1 9 1 0 9 7 1 9 9 9 2 2
48 16 4 1 9 11 11 2 0 9 0 0 9 2 9 1 9 9 1 9 7 0 9 13 4 16 15 15 9 1 0 9 13 1 12 1 12 2 7 15 15 9 13 1 3 0 1 0 2
24 11 7 11 13 4 9 1 0 9 1 1 12 9 2 1 12 1 12 3 1 12 1 12 2
12 9 11 9 4 0 9 0 0 7 0 9 2
9 3 4 0 0 7 0 0 9 2
23 16 7 1 0 9 2 9 9 15 4 0 16 0 13 12 2 15 4 12 9 0 9 2
24 12 9 0 11 2 11 2 11 2 11 2 11 2 11 11 2 11 7 11 2 13 15 9 2
26 11 2 11 7 11 2 11 7 11 13 15 1 12 3 0 9 2 15 13 12 9 0 9 1 9 2
8 9 0 9 13 15 1 12 2
12 15 3 13 12 9 2 3 12 9 0 9 2
15 3 1 9 15 9 13 1 11 2 15 3 13 15 9 2
7 9 1 9 11 13 0 9
11 4 14 0 9 11 9 9 7 9 9 2
21 9 11 13 4 1 9 0 9 1 9 9 9 1 16 15 4 3 0 12 9 2
26 9 9 15 4 13 13 4 15 9 1 9 2 7 9 4 13 3 1 3 9 16 4 9 4 0 2
12 1 9 2 9 11 13 7 0 7 0 9 2
23 0 4 16 4 11 13 0 9 1 9 9 1 9 2 7 16 4 9 7 3 3 0 2
19 1 0 9 2 11 4 13 16 4 0 0 9 13 3 0 9 1 11 2
15 3 2 15 4 0 9 1 9 1 9 9 1 12 9 2
15 0 9 2 0 0 9 1 0 9 2 0 4 0 9 2
18 1 0 0 9 3 3 3 13 3 1 12 0 1 0 9 16 13 2
9 0 9 7 3 4 1 0 9 2
22 3 4 1 0 9 8 8 2 11 4 3 13 16 13 4 0 3 1 9 9 9 2
29 2 16 13 9 13 16 4 9 0 16 0 9 7 15 1 15 13 9 11 2 2 13 4 9 0 9 11 11 2
20 2 1 9 15 3 13 16 4 11 13 0 9 1 9 7 9 1 11 2 2
18 11 11 2 1 3 0 9 0 9 2 11 2 2 13 3 0 9 2
10 2 9 13 16 1 11 14 13 9 2
17 15 13 16 9 4 13 13 9 1 9 1 9 1 12 9 2 2
34 16 9 13 0 9 2 15 4 3 15 11 4 13 16 4 0 16 9 1 0 9 2 13 11 11 1 9 1 0 11 2 11 2 2
10 2 13 0 9 2 2 13 4 11 2
32 2 12 9 0 4 1 15 9 2 15 4 3 0 0 9 2 7 15 4 9 7 9 2 1 15 4 15 9 3 0 2 2
24 2 3 4 16 13 0 9 2 7 15 14 13 13 16 9 4 0 1 9 2 2 13 4 2
28 9 13 11 2 13 11 11 1 9 1 9 11 2 11 2 2 3 16 4 15 9 11 2 13 12 9 2 2
29 9 1 11 0 4 9 9 2 1 8 8 2 0 9 1 8 8 2 1 15 15 13 1 0 9 0 9 11 2
22 2 9 13 0 9 1 11 2 2 13 4 1 11 11 11 1 0 9 1 0 9 2
21 2 11 4 13 16 4 13 0 9 2 7 15 14 13 13 16 9 1 0 9 2
21 1 15 2 13 4 15 13 1 9 9 7 9 1 9 15 9 15 4 0 2 2
27 2 13 4 0 1 9 9 2 2 13 4 11 2 3 16 4 9 1 0 9 0 9 9 1 0 11 2
11 9 15 2 13 4 2 13 13 1 9 2
17 2 7 0 9 7 9 13 13 1 9 9 2 2 13 4 11 2
8 0 9 2 0 9 11 13 11
23 11 4 0 13 15 9 15 4 13 1 15 0 0 9 2 13 4 9 15 9 0 9 2
13 3 15 9 2 0 9 13 9 1 9 11 11 2
25 0 9 11 11 13 4 15 9 1 11 3 4 13 0 9 1 9 11 7 13 15 1 0 9 2
18 11 4 1 9 2 12 9 2 13 0 9 1 15 9 9 9 9 2
39 2 11 4 4 1 0 9 15 4 13 9 11 2 16 13 16 4 15 9 1 11 2 2 13 4 11 3 16 4 11 0 13 9 1 15 0 0 9 2
20 0 9 13 4 9 1 9 11 11 2 13 4 9 1 9 2 12 9 2 2
10 11 4 13 12 9 15 4 13 9 2
19 9 0 9 11 11 13 4 1 9 2 12 9 2 0 9 11 7 11 2
19 11 4 1 11 13 9 11 9 11 11 2 3 16 9 2 13 9 2 2
22 4 4 2 3 2 15 15 9 4 13 9 1 9 1 11 1 0 9 2 13 4 2
21 1 9 4 13 1 11 1 9 1 9 11 11 2 9 9 9 7 9 9 11 2
23 9 0 9 11 11 13 4 1 9 2 12 9 2 1 11 3 0 9 9 1 15 9 2
14 9 0 9 11 11 13 15 1 11 7 13 9 9 2
12 2 11 13 0 9 1 9 2 2 13 4 2
29 0 9 11 11 13 15 1 9 2 12 9 2 1 0 9 1 11 11 11 1 15 4 13 1 0 7 0 9 2
14 13 4 15 1 9 9 16 4 15 13 9 9 9 2
15 2 9 9 13 9 0 9 1 9 2 2 13 4 11 2
10 9 1 9 0 9 13 0 7 0 9
21 9 0 9 0 1 11 15 13 11 13 1 0 9 0 1 9 1 9 1 11 2
14 1 11 4 0 9 9 1 9 9 1 0 0 9 2
20 3 12 0 9 4 4 0 1 9 0 9 1 9 1 11 2 13 0 9 2
46 0 2 0 9 9 9 15 4 3 13 11 2 2 9 4 0 1 9 1 0 9 1 12 0 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 7 11 2
23 3 4 0 9 12 0 9 1 0 9 0 0 9 2 11 2 7 12 1 9 9 11 2
13 0 9 0 4 12 9 2 3 3 11 7 11 2
14 15 9 0 4 16 4 13 1 12 9 9 1 9 2
16 8 3 0 9 0 4 1 11 2 13 15 1 9 0 9 2
30 0 9 1 0 11 7 0 11 15 4 0 1 9 2 7 15 4 11 13 12 2 1 9 4 2 13 0 9 11 2
16 3 12 9 0 0 0 9 2 0 9 2 13 15 1 9 2
20 11 11 2 9 0 9 11 1 11 2 13 4 16 4 12 9 0 13 9 2
5 13 4 12 9 2
17 11 3 13 16 4 9 9 11 4 0 1 9 9 1 9 12 2
6 9 4 0 1 9 2
20 2 16 15 4 4 9 2 15 15 4 13 9 1 9 2 3 13 1 9 2
15 15 4 9 1 9 15 9 2 2 13 4 11 9 11 2
19 1 9 11 2 0 0 9 13 4 0 9 9 1 9 9 1 0 9 2
14 9 4 13 9 1 0 9 16 3 13 9 1 9 2
31 9 9 11 11 13 16 1 0 9 9 3 3 14 13 0 9 1 9 9 2 7 13 9 0 9 11 2 9 0 9 2
18 11 13 16 4 11 13 0 9 1 9 1 9 2 3 9 7 9 2
7 2 0 4 9 0 9 2
9 15 4 15 9 2 2 13 4 2
18 1 11 7 11 2 12 9 1 0 7 0 9 3 4 3 4 0 2
23 9 9 13 4 11 1 9 0 9 1 9 12 0 9 1 9 9 0 9 1 8 9 2
21 11 4 2 1 15 2 13 0 0 9 1 12 0 0 9 15 4 1 15 9 2
23 9 0 9 3 3 4 9 9 2 7 1 0 9 0 9 1 9 2 9 4 13 0 2
14 11 13 16 15 12 9 9 13 1 0 9 15 9 2
9 1 0 9 9 0 9 1 9 11
23 9 11 12 7 9 9 9 1 9 1 0 0 4 4 15 0 9 0 1 11 15 9 2
20 0 9 9 2 11 2 13 4 15 9 13 0 9 15 15 13 1 9 11 2
31 9 4 0 1 15 13 14 9 9 0 9 1 0 0 2 4 14 0 0 9 11 2 7 13 14 9 12 11 9 9 2
27 11 4 1 9 2 12 9 2 13 9 11 2 11 7 11 2 9 1 15 4 15 13 7 0 0 9 2
6 11 4 13 0 9 2
39 9 9 4 0 9 0 9 2 13 4 0 9 9 9 11 2 11 2 3 15 15 15 9 13 3 1 9 12 9 2 7 14 1 9 1 9 7 9 2
41 9 11 11 11 11 13 4 9 16 15 15 0 9 3 13 1 15 9 1 11 12 9 2 3 16 9 9 4 2 0 1 15 2 2 9 9 0 0 9 2 2
29 9 9 1 9 11 13 4 16 2 9 3 0 9 2 3 1 9 0 9 2 15 4 0 9 9 9 9 2 2
37 11 4 2 1 9 2 13 16 15 7 11 7 0 11 14 13 13 0 9 0 0 9 11 2 7 0 15 4 2 8 8 2 13 9 1 11 2
13 1 9 2 0 0 9 7 11 13 4 0 9 2
46 0 9 11 11 11 13 4 16 4 9 9 11 1 9 1 9 12 11 2 1 15 15 2 3 4 13 2 2 13 2 1 9 2 16 4 9 13 4 0 9 1 0 9 11 2 2
23 1 9 15 2 3 15 14 13 1 0 9 0 9 11 1 0 9 2 2 13 4 11 2
23 1 15 2 13 4 2 9 3 13 4 15 9 16 4 11 9 11 2 1 9 1 11 2
25 3 15 1 9 11 2 9 11 11 11 13 4 16 4 9 11 3 4 2 0 16 9 9 2 2
21 9 12 2 13 4 2 14 13 4 0 3 16 13 2 9 12 9 0 9 2 2
20 3 2 13 4 11 2 15 4 4 12 1 9 1 15 4 11 13 1 9 2
14 0 9 1 11 2 13 4 2 2 3 3 13 2 2
24 3 12 9 2 1 11 7 11 2 13 4 15 0 9 1 9 2 3 15 13 15 9 9 2
52 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 1 9 4 15 15 13 1 11 2 16 4 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 0 11 13 1 9 9 11 2
20 1 9 2 11 4 13 0 9 0 11 15 4 13 15 9 1 0 9 9 2
29 11 4 13 16 4 11 13 0 9 1 0 11 2 7 4 9 11 16 4 15 9 0 11 2 1 0 9 2 2
7 9 1 0 9 9 1 11
20 9 1 0 9 1 11 13 1 9 0 9 9 9 2 13 15 1 0 9 2
20 9 0 9 1 11 7 11 13 4 0 9 9 1 9 7 9 9 1 11 2
11 1 9 4 0 16 4 9 7 3 0 2
30 2 9 9 1 9 7 9 4 4 7 13 12 1 0 9 1 0 9 1 11 2 2 13 4 9 9 11 11 11 2
32 2 1 0 9 7 0 9 9 9 9 1 0 9 2 9 9 15 4 0 13 1 9 7 3 4 3 0 2 2 13 4 2
13 2 9 9 9 13 15 3 2 2 13 4 11 2
35 1 9 2 9 9 9 1 11 13 4 0 9 15 15 13 0 9 1 0 9 9 9 2 3 2 7 4 0 2 9 9 7 15 9 2
17 0 4 9 0 9 15 4 13 3 0 9 2 13 15 1 9 2
21 0 9 13 4 4 3 0 1 0 9 9 1 15 4 0 2 13 15 1 9 2
29 2 3 14 4 15 0 2 15 9 9 13 4 15 13 1 0 9 1 9 9 1 9 2 2 13 15 1 9 2
44 2 1 0 9 1 9 9 2 1 9 4 14 15 9 7 9 9 2 11 15 14 13 13 4 15 0 9 1 0 9 0 9 7 0 0 0 9 2 2 13 4 11 9 2
13 0 9 13 4 11 11 2 9 0 9 1 11 2
21 2 13 15 16 4 15 9 13 0 9 1 9 9 7 9 9 2 2 13 4 2
36 9 0 9 13 4 16 0 9 1 0 9 13 1 9 15 4 0 13 1 9 0 9 7 13 1 15 9 2 13 4 9 0 9 7 11 2
17 15 9 0 4 7 9 7 9 0 9 4 1 9 13 0 9 2
9 11 7 11 0 1 9 9 0 9
26 9 0 9 7 9 1 9 9 0 4 1 9 11 7 11 1 9 0 9 2 13 4 0 0 9 2
31 11 7 11 2 11 2 13 13 0 9 2 3 7 9 9 2 16 13 13 9 9 1 11 7 11 2 13 4 0 9 2
23 13 4 16 4 9 9 1 0 9 13 13 0 9 9 7 13 1 9 2 9 7 9 2
68 2 0 3 9 2 3 7 9 2 4 4 1 0 9 1 9 11 2 2 13 15 1 9 9 0 9 0 1 9 2 12 0 2 2 7 13 16 0 0 9 1 11 11 11 2 3 13 16 9 1 11 2 7 3 1 11 2 13 0 9 11 1 0 9 7 9 2 2
34 2 9 11 7 9 3 4 0 1 11 15 9 13 13 13 14 13 9 13 0 9 1 11 7 0 0 9 2 2 13 15 1 9 2
36 1 11 4 1 9 9 9 9 15 1 9 13 9 9 11 1 9 9 1 9 9 1 9 7 9 1 9 2 15 4 0 9 1 0 9 2
26 1 9 4 0 9 9 9 9 11 1 9 0 9 11 1 15 4 15 13 1 9 9 1 9 9 2
28 0 9 11 1 0 9 7 9 11 11 13 4 16 4 9 0 9 1 0 9 1 9 11 16 15 13 11 2
28 2 11 4 3 13 11 15 9 2 2 13 4 11 1 9 0 0 9 0 9 2 7 13 0 9 8 8 2
11 2 16 13 9 2 9 11 4 4 0 2
25 16 13 9 2 13 4 15 1 9 9 11 1 9 0 9 2 9 7 9 2 2 13 4 11 2
33 3 0 9 1 0 9 9 0 9 1 11 1 9 9 2 11 4 13 2 16 4 1 15 9 9 11 4 3 7 3 0 2 2
22 9 1 9 13 9 0 9 12 9 1 11 1 0 9 2 9 0 0 7 0 9 2
23 0 9 13 9 9 9 1 9 9 7 0 9 1 15 9 4 4 12 9 7 12 9 2
14 9 11 4 4 0 0 9 9 0 9 7 9 9 2
36 1 0 9 1 9 9 15 4 13 1 12 1 12 9 2 9 12 9 1 9 13 4 0 9 7 13 0 9 1 12 9 2 9 7 9 2
41 3 15 9 7 11 7 9 11 2 9 9 11 11 13 4 16 4 9 9 9 0 9 1 9 11 9 11 9 1 9 15 9 2 15 13 0 9 1 9 9 2
19 1 9 9 1 9 9 1 11 2 1 9 1 11 13 4 13 12 9 2
20 0 0 9 0 9 13 15 9 2 3 16 15 15 14 13 9 12 0 9 2
20 1 9 2 1 9 4 0 9 9 11 1 11 2 1 9 1 9 9 9 2
50 3 4 0 7 9 9 1 9 9 2 15 4 1 0 9 2 3 4 13 11 2 2 13 4 14 0 9 1 11 0 13 0 9 7 0 9 7 13 9 3 0 1 9 9 1 9 0 9 2 2
9 9 15 13 9 2 9 13 0 9
23 0 9 9 2 0 9 7 9 9 1 9 0 9 1 0 0 9 13 1 9 0 9 2
10 0 9 3 4 12 1 0 0 9 2
17 0 1 9 11 7 11 2 0 9 12 4 1 0 0 9 9 2
13 0 4 1 3 15 2 1 15 9 3 13 9 2
18 3 12 0 9 9 13 1 9 0 0 9 1 0 0 9 7 9 2
8 3 2 1 0 9 13 9 2
18 1 15 2 0 4 9 2 0 7 3 0 9 15 13 1 0 9 2
10 9 15 9 13 9 7 9 3 0 2
19 9 13 16 4 9 7 9 2 3 0 1 9 1 9 7 15 9 2 2
15 3 16 0 0 9 13 0 9 2 13 1 0 0 9 2
32 9 9 1 0 9 7 0 9 9 1 9 13 4 1 0 9 0 9 9 7 9 7 9 0 9 1 9 9 2 13 9 2
27 9 1 12 0 9 2 7 1 9 1 0 9 2 1 9 13 3 1 9 2 7 3 7 0 9 9 2
12 0 4 9 0 9 2 16 4 0 3 0 2
12 9 13 16 4 0 9 9 13 14 0 9 2
34 2 1 16 9 13 12 9 1 9 2 9 4 15 13 3 1 9 2 2 13 4 9 9 1 11 11 11 2 0 9 1 9 11 2
10 2 3 4 13 0 9 7 13 0 2
7 7 15 4 13 9 2 2
17 1 9 9 2 0 9 11 13 0 9 15 13 0 9 0 9 2
29 2 13 14 15 4 15 13 15 9 15 13 9 1 9 0 9 2 2 2 13 4 9 9 11 11 2 0 9 2
35 1 12 0 9 1 3 1 12 9 2 11 7 3 12 3 13 9 1 9 0 9 2 13 0 9 9 1 9 0 16 9 1 9 11 2
23 2 9 1 9 0 7 9 0 9 1 9 3 15 13 1 12 9 9 2 2 13 15 2
28 2 0 9 1 3 12 9 13 4 0 16 4 15 13 9 9 7 9 4 0 2 16 9 3 4 13 2 2
6 9 9 0 4 9 2
16 9 1 9 0 9 1 0 12 9 14 13 9 2 13 9 2
40 1 9 1 9 1 9 11 2 11 4 12 13 3 4 1 9 15 9 0 9 13 1 9 1 0 9 2 13 4 9 9 9 11 11 1 9 0 0 9 2
16 3 2 0 12 9 3 4 13 15 9 0 1 9 15 9 2
22 1 15 2 9 4 9 0 1 9 0 9 2 15 4 9 4 15 9 0 1 11 2
32 3 16 0 9 13 0 0 9 1 14 0 9 15 9 2 11 13 1 15 16 4 11 4 1 9 13 9 1 0 12 9 2
18 0 9 0 9 0 0 9 13 0 9 0 9 2 3 9 7 9 2
13 9 15 9 13 9 9 2 15 13 9 0 9 2
9 0 9 9 13 4 0 9 9 2
23 13 15 16 4 9 2 3 15 15 9 13 2 3 13 9 0 9 7 9 9 15 9 2
33 0 9 0 9 9 2 9 7 0 9 2 9 3 0 0 9 2 9 0 9 7 9 0 9 1 9 0 4 16 0 0 9 2
31 1 9 11 1 12 13 15 16 12 0 9 13 3 12 0 9 0 7 0 9 15 13 1 0 9 16 9 0 0 9 2
23 2 9 15 9 2 16 7 3 0 1 0 12 2 1 9 13 9 11 2 2 13 15 2
34 9 4 0 12 9 1 15 4 12 1 11 0 9 1 9 0 9 1 9 2 15 12 0 9 13 15 9 9 9 7 0 9 9 2
43 9 9 1 11 2 3 12 3 0 9 1 9 0 9 9 2 9 9 7 1 0 9 1 9 9 2 1 9 9 2 13 9 1 0 9 2 15 15 9 13 1 11 2
11 9 15 13 1 9 9 1 9 0 9 2
26 3 2 7 3 4 3 0 1 9 1 0 0 7 0 9 2 13 9 2 3 11 16 0 9 9 2
30 2 9 1 9 9 9 3 4 0 9 0 9 7 9 0 9 2 7 14 0 9 9 2 2 12 4 1 9 11 2
18 2 13 4 3 9 16 15 9 9 9 1 9 13 1 0 9 2 2
32 9 4 13 7 3 0 9 1 0 0 9 2 1 15 15 13 16 4 0 3 1 15 9 2 7 4 13 9 9 0 9 2
20 13 4 7 16 13 0 9 1 9 1 9 7 0 9 1 9 9 7 9 2
17 2 3 12 0 9 13 4 13 0 9 1 0 9 2 2 13 2
8 0 9 2 0 9 9 1 11
16 9 0 9 1 11 0 4 1 12 9 1 0 9 12 9 2
14 3 1 0 9 15 9 2 0 9 13 0 9 11 2
10 9 0 9 1 11 0 4 12 9 2
31 9 0 9 1 11 0 1 12 9 1 0 9 12 9 2 13 9 15 4 1 9 2 12 9 2 13 9 0 9 9 2
17 11 13 0 1 0 9 2 3 11 2 15 4 3 9 4 0 2
20 11 4 3 13 1 0 9 2 16 4 1 0 9 12 9 0 9 13 11 2
25 11 4 1 9 13 3 12 9 9 9 0 9 7 0 0 9 2 13 4 12 9 9 11 11 2
13 15 9 4 4 0 1 3 12 0 9 1 9 2
23 11 15 13 16 4 4 0 1 9 3 0 9 7 1 15 4 0 16 9 1 0 9 2
36 9 0 9 1 11 2 11 11 2 13 4 16 4 9 13 0 9 15 9 1 9 15 1 9 13 9 0 9 1 9 7 9 0 9 11 2
12 0 9 9 3 3 4 0 2 13 4 11 2
14 15 9 0 9 4 4 0 1 9 9 1 9 9 2
25 0 9 1 9 7 9 11 13 4 0 9 1 9 12 9 9 2 13 15 1 0 9 0 9 2
45 8 8 8 2 8 2 8 8 2 8 8 2 8 2 0 9 11 7 8 8 0 4 0 9 15 4 13 9 2 15 4 9 9 12 9 1 9 12 9 9 1 1 9 9 2
22 0 0 9 11 13 15 1 9 7 9 1 12 9 1 0 9 2 3 12 9 9 2
17 9 0 0 9 15 13 9 9 1 11 16 9 9 11 1 9 2
39 1 0 12 9 15 9 2 9 4 13 12 9 9 2 3 9 1 12 9 1 0 9 2 16 4 9 0 1 12 9 1 0 9 2 1 12 9 9 2
23 0 0 9 11 13 4 12 9 9 1 0 9 1 0 12 9 2 13 4 12 9 9 2
30 0 0 9 11 13 15 1 9 9 9 9 11 9 2 9 0 9 9 11 11 9 2 16 7 9 9 9 1 11 2
7 0 9 2 0 9 13 11
11 9 11 8 11 13 4 1 9 1 11 2
20 3 1 0 9 2 0 9 11 11 13 15 1 0 9 0 9 11 11 2 2
28 0 9 11 11 2 8 2 7 9 0 11 11 13 9 0 9 1 9 11 1 11 1 9 2 12 9 2 2
23 0 9 11 11 4 4 1 9 2 12 9 2 9 0 9 1 9 0 9 11 8 11 2
25 11 4 4 0 9 15 9 9 15 4 13 12 9 1 15 4 3 4 11 11 2 11 7 11 2
26 1 0 9 2 11 4 13 16 4 7 11 7 0 11 13 0 9 2 7 4 15 9 13 13 9 2
34 0 9 0 9 11 11 7 15 0 9 11 11 15 4 13 1 9 11 13 4 1 9 2 12 9 2 9 1 9 1 9 9 9 2
17 3 4 13 1 9 16 0 9 13 9 0 9 1 9 1 11 2
25 9 0 9 11 7 11 2 11 2 11 11 13 1 0 9 0 11 1 9 0 9 7 0 9 2
15 11 15 1 9 2 12 9 2 13 1 0 9 11 11 2
10 0 9 15 9 4 9 7 0 9 2
49 3 1 0 9 1 11 1 15 0 9 11 11 0 1 9 2 12 9 2 2 0 9 11 11 13 4 9 16 4 15 9 4 1 9 13 9 1 11 2 7 4 13 16 4 1 9 0 9 2
13 11 4 3 13 9 9 7 9 11 1 15 9 2
31 0 9 0 9 11 11 13 4 11 7 11 2 11 2 1 9 2 12 9 2 16 14 13 1 15 9 1 9 1 11 2
23 1 9 11 13 1 0 9 11 11 11 2 15 0 9 11 11 7 9 0 9 11 11 2
41 0 9 11 11 13 4 1 9 2 12 9 2 9 9 0 9 11 11 11 16 4 9 1 0 9 1 11 1 11 7 9 11 1 0 11 4 0 1 0 9 2
24 11 2 15 4 13 1 11 1 9 9 0 9 2 13 4 0 9 1 0 9 0 1 11 2
39 1 9 1 0 9 11 11 1 9 2 12 9 2 1 11 2 0 9 0 9 11 11 13 4 16 3 3 13 0 9 1 9 9 1 9 11 1 9 2
24 2 13 13 0 0 9 7 13 11 7 11 1 9 9 7 9 1 9 2 2 13 4 11 2
18 9 9 11 11 7 11 13 4 1 9 2 12 9 2 9 1 9 2
28 1 9 4 0 9 0 7 0 9 16 4 15 13 9 7 9 1 9 2 1 9 9 9 0 9 11 11 2
8 9 15 13 1 9 9 1 11
16 0 4 15 9 1 3 1 12 0 13 1 9 13 0 9 2
16 12 3 0 9 13 15 16 4 15 13 1 9 1 0 9 2
30 9 13 1 0 9 2 9 0 0 9 3 1 9 2 7 1 9 9 1 3 0 0 9 7 15 0 9 0 9 2
14 0 9 9 13 13 0 9 1 9 16 4 13 9 2
25 11 2 9 11 11 2 4 4 12 0 0 9 0 1 9 2 7 4 13 12 9 1 0 9 2
32 1 0 4 0 9 3 3 3 9 2 7 9 13 3 9 2 0 0 9 11 7 9 9 1 9 9 0 9 2 11 2 2
18 11 4 1 9 13 9 11 11 7 11 11 2 7 13 0 9 9 2
19 2 9 7 9 1 9 11 1 0 4 9 2 2 13 4 11 1 11 2
16 2 0 4 15 0 9 2 0 9 7 9 1 9 9 2 2
18 3 4 0 9 9 0 9 2 9 0 1 9 2 1 9 1 9 2
23 11 13 0 9 2 0 9 2 0 9 1 0 7 0 9 2 3 0 9 1 0 9 2
9 9 13 7 0 9 1 0 9 2
7 2 11 15 13 1 9 2
41 1 9 9 2 11 4 15 9 13 1 0 9 2 9 1 9 7 0 9 2 7 15 4 9 15 0 9 4 4 1 9 13 1 9 2 2 13 11 1 11 2
26 9 11 2 15 4 13 11 11 2 13 0 9 7 0 4 1 0 9 0 9 1 11 7 0 9 2
45 2 13 16 11 4 0 0 9 2 7 15 13 9 7 0 9 2 9 14 13 4 7 13 0 9 2 15 13 9 15 4 0 1 15 9 2 7 14 1 11 2 2 13 11 2
21 15 4 3 0 0 9 1 11 15 15 9 13 9 9 2 15 3 13 7 9 2
23 2 13 9 15 15 13 15 9 2 7 14 9 15 15 13 9 2 2 13 11 1 11 2
22 9 14 13 13 9 16 13 1 15 9 16 4 1 9 13 0 9 1 9 9 9 2
56 2 14 13 9 7 9 1 9 1 9 2 7 3 4 16 15 4 13 1 9 7 9 9 1 0 9 2 7 13 16 4 9 14 0 15 0 9 2 7 3 3 7 0 9 4 15 9 2 3 16 15 9 13 13 2 2
25 11 7 11 13 15 16 9 15 9 13 1 9 7 0 9 2 16 15 4 0 9 11 11 11 2
24 2 9 1 9 13 2 0 2 9 16 4 0 16 0 9 3 13 1 9 2 2 13 11 2
30 2 9 4 0 16 13 16 15 9 3 13 2 16 4 9 11 1 0 9 2 3 16 7 9 9 2 2 13 11 2
32 11 13 16 4 9 1 9 0 1 0 9 2 7 9 9 13 4 0 1 9 7 0 9 2 7 14 1 0 9 7 9 2
28 11 13 16 4 15 9 3 0 9 0 9 9 9 1 9 9 0 9 2 9 2 0 9 11 7 0 9 2
24 0 9 0 9 2 15 4 13 15 0 9 2 3 4 13 9 16 15 1 9 2 13 11 2
12 2 0 9 3 4 9 1 9 16 1 9 2
7 1 9 4 0 9 0 2
4 3 4 0 2
20 9 11 3 15 3 13 1 0 9 2 7 0 9 3 4 9 1 9 2 2
20 11 13 0 0 9 2 1 15 13 16 4 13 9 2 7 15 13 9 9 2
46 2 0 9 13 1 9 1 15 9 4 0 1 9 1 0 2 1 9 15 13 0 9 1 9 1 9 0 9 2 16 9 4 0 1 9 2 7 1 9 13 9 2 2 13 15 2
16 11 13 16 4 13 1 15 16 15 13 0 0 9 7 9 2
7 9 1 11 14 13 9 2
12 1 15 2 9 13 16 4 3 0 0 9 2
15 11 13 16 4 1 11 3 16 13 13 1 15 1 11 2
30 11 13 16 4 9 2 15 4 13 1 9 7 9 0 9 2 4 1 0 9 0 1 9 11 1 0 9 1 11 2
20 2 9 15 9 0 4 9 11 2 7 14 9 11 1 11 2 2 13 11 2
25 2 1 15 2 11 4 0 16 1 15 9 13 0 9 1 11 2 1 9 0 2 1 11 2 2
35 15 13 9 9 2 7 1 0 9 13 0 11 9 2 15 4 15 9 13 1 9 1 9 9 9 11 3 7 15 9 1 0 9 2 2
29 0 4 9 1 0 9 13 9 3 4 3 13 15 9 7 4 14 13 0 9 16 4 15 0 9 1 0 9 2
29 0 9 9 2 15 4 13 9 11 11 2 13 16 11 13 9 12 2 12 9 2 16 11 13 15 12 2 12 2
10 9 7 9 2 0 9 0 1 9 11
11 9 11 13 4 9 1 9 11 1 11 2
22 3 1 9 1 9 2 11 9 12 0 0 9 2 7 11 7 11 13 9 1 9 2
12 11 11 2 1 9 2 3 4 9 9 11 2
22 9 11 1 11 3 4 1 9 2 12 9 2 13 0 9 11 11 2 13 4 9 2
9 0 12 9 9 4 13 9 9 2
32 0 9 2 9 1 8 11 7 9 0 0 9 2 13 4 16 4 3 13 9 7 3 15 13 1 9 12 9 16 0 9 2
10 9 9 13 1 9 9 16 0 9 2
17 1 11 4 15 1 12 9 1 9 15 9 13 12 0 0 9 2
40 1 9 4 13 3 0 9 1 11 11 2 9 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 9 11 11 2 11 11 7 0 0 9 8 11 2
9 9 13 0 9 1 9 7 9 2
48 11 7 11 13 4 9 1 9 1 9 2 9 2 0 9 2 0 9 2 0 9 0 9 7 9 0 7 0 9 1 9 15 15 13 1 12 9 2 13 4 1 9 2 12 9 2 11 2
6 9 4 0 1 11 2
20 9 0 0 7 0 9 2 11 2 13 15 1 9 2 12 9 2 1 11 2
23 1 9 2 15 13 12 9 2 3 4 13 9 1 11 2 11 2 11 2 11 7 11 2
25 0 0 0 9 13 4 0 9 11 12 15 4 1 12 9 1 9 2 12 9 2 0 1 11 2
9 1 0 9 2 9 4 13 11 2
14 0 9 11 11 2 12 2 0 4 0 9 1 9 2
23 11 11 0 4 1 9 2 12 9 2 1 9 0 9 11 1 9 9 1 0 0 9 2
10 4 4 0 9 15 4 13 0 9 2
21 0 9 2 11 11 11 2 13 4 9 1 9 11 1 11 12 2 12 0 9 2
9 11 13 9 15 0 9 1 9 11
19 11 4 13 9 0 9 1 15 0 9 1 9 11 2 1 9 11 11 2
13 11 11 13 4 1 9 1 9 2 12 9 2 2
34 11 4 1 9 2 12 9 2 13 9 0 9 11 11 1 15 0 9 1 9 11 2 1 15 4 0 9 11 11 13 16 15 13 2
29 2 0 4 1 9 9 1 9 7 0 9 7 0 4 16 13 3 13 9 9 11 2 2 13 4 11 1 9 2
14 9 4 13 1 9 0 9 1 0 9 7 9 11 2
24 15 4 1 9 13 9 9 11 11 3 1 15 16 13 15 9 2 1 0 9 2 15 13 2
39 0 9 0 9 2 11 2 2 11 4 0 1 9 0 9 1 0 9 9 1 0 9 11 2 11 2 2 9 0 9 2 1 0 9 1 9 12 9 2
41 0 9 2 0 4 9 11 1 9 1 0 9 2 11 2 1 0 9 9 11 11 11 7 1 9 4 0 1 0 9 11 1 0 9 2 0 9 7 9 9 2
17 11 4 3 0 1 9 0 0 9 2 11 2 15 4 11 9 2
32 1 0 9 1 15 9 12 9 2 11 4 0 1 9 0 7 0 9 11 1 9 1 9 16 4 13 15 9 1 0 9 2
21 15 9 1 0 9 0 1 9 3 4 13 9 1 15 9 1 9 1 0 9 2
42 0 9 11 2 1 15 4 0 13 9 11 1 8 8 8 2 2 0 0 9 15 4 13 1 9 1 9 2 13 4 1 9 16 4 4 15 0 9 1 15 9 2
19 1 15 2 13 15 9 1 15 9 2 15 4 13 9 11 1 0 9 2
14 0 9 9 1 9 4 13 13 0 9 1 15 9 2
26 1 9 11 2 9 11 13 9 13 9 1 9 1 15 0 9 7 13 0 9 2 7 14 9 3 2
25 9 0 9 1 0 0 9 12 9 3 4 13 0 7 0 9 11 11 7 11 11 1 9 9 2
27 1 9 11 1 9 2 9 11 11 11 13 4 16 4 9 1 0 11 4 0 1 12 9 1 12 9 2
25 9 1 9 11 0 4 1 12 9 2 15 15 13 12 9 3 16 0 9 1 9 1 9 11 2
29 0 9 7 9 2 15 15 13 0 9 12 9 2 3 4 1 9 13 1 9 0 9 2 7 3 1 0 9 2
32 16 9 1 0 9 1 9 12 2 12 2 13 4 9 1 0 9 9 1 0 9 7 13 9 1 12 9 9 1 0 9 2
25 11 4 3 4 9 1 11 1 12 9 2 3 4 13 9 1 9 7 9 1 9 0 9 9 2
15 0 4 1 9 7 0 9 9 0 9 1 9 12 9 2
25 1 9 0 9 11 1 9 3 2 11 4 13 15 0 9 1 9 9 11 1 9 9 0 9 2
26 1 9 4 13 16 4 15 13 0 9 9 11 11 2 15 4 15 0 9 13 15 9 9 11 11 2
29 11 4 3 13 16 13 0 9 9 9 7 13 15 0 9 11 11 2 9 1 0 0 9 8 2 1 15 9 2
6 15 9 13 13 9 2
7 9 11 13 0 9 1 11
14 9 0 16 13 0 9 13 4 15 1 11 7 11 2
22 0 9 0 9 11 11 2 3 2 1 9 9 11 11 11 2 13 4 11 1 9 2
31 0 9 0 0 9 2 3 0 9 1 9 9 1 9 16 13 0 9 2 13 4 0 9 1 11 7 11 2 11 2 2
16 9 9 0 4 1 0 9 11 16 13 9 1 11 7 3 2
24 12 9 4 0 2 9 11 1 11 2 1 3 7 1 3 2 13 0 9 1 15 0 9 2
18 15 13 0 9 2 16 0 13 16 4 15 13 13 0 7 0 9 2
15 11 7 11 4 3 12 9 13 0 9 2 9 0 11 2
25 1 9 0 9 2 3 4 13 9 1 11 1 0 9 2 0 9 0 9 11 11 13 4 11 2
27 15 4 3 13 9 0 9 2 7 13 15 7 1 0 0 9 7 9 2 3 0 9 1 11 11 11 2
20 11 4 1 15 9 3 13 11 16 0 9 1 9 1 9 1 11 7 11 2
21 3 4 13 0 9 1 9 1 9 15 15 13 1 11 7 1 9 0 9 9 2
10 15 9 3 4 0 2 3 1 9 2
13 15 4 0 16 9 0 9 9 11 16 0 9 2
57 9 9 9 0 0 9 1 9 2 11 11 1 9 0 9 2 11 2 2 11 11 1 9 1 11 7 11 2 11 2 7 11 11 1 0 9 2 11 2 2 13 4 9 1 0 9 1 11 9 9 0 11 0 9 1 11 2
7 3 2 9 3 4 0 2
16 3 4 11 13 9 3 16 4 9 9 0 2 7 14 0 2
9 0 9 0 13 4 16 4 13 2
22 3 15 13 16 4 9 1 9 0 7 0 7 0 9 11 1 0 0 9 7 9 2
25 1 15 4 4 0 9 9 9 11 2 11 2 11 7 11 2 16 7 9 11 11 2 0 11 2
29 9 4 4 0 7 0 2 7 9 9 9 11 1 9 0 11 11 13 4 0 9 1 11 9 9 0 0 9 2
29 3 2 9 9 0 9 2 11 2 2 0 9 2 13 4 9 1 15 15 13 0 9 1 11 7 11 1 9 2
41 2 0 4 9 15 4 0 9 13 16 4 13 11 1 9 0 9 2 7 3 13 16 4 15 9 2 3 15 15 13 0 9 2 0 2 2 13 15 1 9 2
21 1 9 11 1 9 2 11 4 13 0 0 0 9 7 9 1 9 1 0 9 2
33 11 4 0 9 4 0 0 0 9 1 11 2 1 12 9 9 2 1 11 2 11 7 11 2 13 4 9 11 1 9 0 9 2
5 0 9 11 13 9
21 0 9 9 2 9 9 2 13 15 1 15 9 1 9 9 9 1 0 11 11 2
8 11 13 13 12 9 9 3 2
30 11 2 3 0 9 1 9 2 4 4 0 15 9 1 9 11 1 0 11 11 1 9 9 1 9 2 12 9 2 2
44 0 9 9 0 12 9 13 15 1 0 9 0 9 12 9 3 4 15 9 9 1 0 9 0 1 9 0 0 9 2 15 15 4 13 16 13 1 9 7 13 1 0 9 2
21 13 15 16 4 15 1 9 9 9 3 13 16 4 11 13 4 0 1 15 9 2
11 9 3 9 13 4 1 0 9 1 9 2
20 2 9 1 9 4 4 0 16 13 1 15 9 2 2 13 4 8 8 8 2
33 2 9 0 9 1 0 9 2 15 4 13 1 9 2 13 4 16 9 13 16 13 9 15 13 0 9 2 2 13 4 8 8 2
17 9 1 11 11 13 4 3 16 4 13 11 3 16 15 14 13 2
28 2 16 15 9 13 7 14 4 13 3 3 2 15 4 15 0 3 13 2 2 13 4 12 1 9 0 9 2
9 2 15 13 9 3 16 0 9 2
51 1 9 16 4 11 13 13 0 0 9 16 13 1 11 2 15 13 0 9 1 11 11 7 13 15 3 12 9 1 9 11 2 0 4 16 15 13 1 9 3 16 15 4 13 9 1 9 3 4 13 2
32 2 11 13 13 3 9 2 7 15 4 3 0 9 9 2 3 14 4 13 9 3 13 2 2 13 4 11 11 2 9 9 2
14 11 4 0 1 15 16 13 7 1 12 9 9 3 2
8 9 1 11 2 9 4 9 2
13 15 4 0 1 9 0 9 7 3 13 15 9 2
19 9 13 13 3 1 0 9 1 0 9 2 16 13 7 0 9 7 9 2
15 3 9 0 9 13 4 15 16 4 11 2 0 9 2 2
13 3 2 11 11 13 4 9 7 9 1 0 9 2
21 2 15 4 0 2 0 9 15 4 13 15 7 15 15 13 2 2 13 4 11 2
25 2 11 14 13 9 1 4 15 2 2 13 4 11 2 2 3 16 15 14 13 7 13 15 2 2
19 7 16 4 15 0 9 4 0 2 11 4 13 1 0 9 7 0 9 2
16 2 14 13 3 13 16 4 15 13 16 13 3 13 7 13 2
21 16 15 13 16 4 15 0 2 3 13 3 12 9 1 15 2 2 13 4 11 2
22 15 7 15 9 2 15 4 9 9 1 9 2 13 4 9 0 9 1 15 0 9 2
10 11 4 13 1 9 1 15 0 9 2
19 1 3 9 0 0 9 13 4 0 9 9 1 11 16 4 4 15 9 2
11 9 9 13 4 3 4 11 13 15 9 2
10 11 13 16 4 9 4 0 1 9 2
16 2 11 15 4 13 1 0 9 2 7 4 15 4 0 2 2
10 8 8 8 13 4 11 16 4 0 2
20 2 9 13 4 0 2 7 3 1 15 15 13 9 16 9 9 3 13 9 2
18 9 4 16 13 14 4 3 0 9 9 2 3 14 13 13 3 2 2
5 0 9 1 0 9
22 3 1 9 9 9 2 9 9 7 9 0 9 2 0 9 1 11 11 3 15 13 2
6 9 1 11 13 0 2
27 1 0 9 9 2 11 9 13 4 1 12 9 1 12 9 2 7 4 1 9 11 15 9 13 12 9 2
21 1 9 16 4 9 13 9 1 0 9 1 12 9 2 11 15 13 1 0 9 2
10 9 7 9 3 13 3 12 9 3 2
8 9 7 9 13 3 12 9 2
28 1 9 2 9 9 13 4 2 9 1 0 9 1 11 13 3 12 9 3 2 15 0 13 9 9 1 9 2
10 1 0 2 15 0 9 4 13 9 2
21 0 9 13 16 4 12 1 0 9 15 15 9 4 13 15 0 7 3 0 9 2
16 3 2 0 0 9 2 9 0 0 9 2 7 3 13 9 2
34 2 0 2 0 7 0 9 1 9 9 0 9 2 9 9 2 9 2 9 2 0 7 0 9 7 0 9 13 4 4 0 0 9 2
33 0 9 1 0 9 13 2 13 2 0 9 2 1 0 9 1 0 9 1 0 9 2 2 13 9 9 1 9 7 9 11 11 2
12 9 4 13 9 0 9 16 4 13 0 9 2
6 0 9 3 15 13 2
27 1 12 1 12 9 13 4 0 9 9 1 11 7 0 11 1 9 1 0 9 2 7 15 3 4 9 2
16 0 4 9 3 0 9 13 4 0 1 9 9 1 9 9 2
40 2 9 1 9 13 2 2 2 9 2 15 4 13 4 0 1 9 9 1 0 9 2 15 4 15 13 0 3 9 2 2 13 4 11 2 3 9 0 9 2
17 11 13 16 0 9 13 0 9 2 7 11 11 4 3 0 9 2
19 12 1 9 4 2 3 2 15 15 4 9 1 9 0 9 3 13 9 2
31 2 3 13 3 12 9 15 4 0 9 13 0 9 2 15 4 0 9 2 2 13 4 0 9 0 9 11 11 1 11 2
15 0 0 9 13 4 16 4 1 9 3 9 4 12 9 2
16 1 9 16 9 4 13 9 2 9 13 16 4 13 13 9 2
7 0 9 9 13 12 9 2
25 3 2 0 9 3 4 3 0 2 3 15 15 15 15 4 13 1 9 1 9 14 13 4 0 2
36 2 0 9 9 2 3 1 0 9 2 4 4 3 12 9 9 1 9 12 9 2 7 1 9 12 13 4 12 9 9 2 2 13 4 11 2
36 3 16 4 11 11 0 9 13 0 9 1 12 9 9 2 9 9 11 11 11 13 16 15 0 9 9 13 3 1 9 16 1 3 0 9 2
7 2 0 9 13 0 9 2
32 11 13 3 13 9 9 1 9 7 3 13 13 14 15 9 4 0 9 2 9 9 7 0 9 2 2 13 4 11 1 11 2
7 0 9 11 13 9 1 9
38 0 9 11 11 11 13 4 1 9 16 4 13 14 13 9 2 7 4 15 1 15 13 1 9 9 1 9 15 4 0 9 7 1 9 15 13 11 2
51 0 9 11 11 11 13 4 1 9 2 12 9 2 16 4 13 1 15 9 1 9 9 2 7 4 1 15 13 1 9 15 9 7 13 15 1 9 9 1 9 0 9 2 16 7 1 9 15 13 11 2
17 2 0 9 14 13 13 15 9 1 0 9 2 2 13 4 11 2
13 2 16 4 3 13 9 15 4 4 9 9 2 2
34 9 4 9 1 9 0 9 13 12 9 2 9 1 15 4 0 9 3 13 0 9 9 15 4 3 0 1 9 11 1 11 12 9 2
21 2 16 4 13 9 4 13 1 9 9 0 9 2 2 13 4 11 9 1 9 2
8 2 13 4 9 0 9 9 2
30 13 4 1 12 9 9 1 2 2 2 9 1 9 9 1 9 2 9 1 11 7 9 9 1 15 4 13 9 2 2
21 1 0 9 2 0 9 9 1 15 4 15 13 1 9 13 4 4 0 1 9 2
16 13 15 16 4 11 1 9 13 9 2 1 9 11 0 9 2
25 15 4 15 13 9 1 0 9 15 9 2 15 4 15 1 15 15 9 11 11 13 3 1 9 2
28 9 2 16 15 13 2 13 16 4 0 9 13 1 9 0 9 0 9 2 15 4 15 13 0 9 0 9 2
44 3 2 9 0 9 9 8 1 9 13 4 9 1 9 0 9 1 9 0 9 15 15 4 0 1 9 9 0 9 2 7 0 9 13 3 4 9 11 3 13 9 0 9 2
30 9 1 11 13 4 9 16 4 0 9 13 13 9 9 1 11 0 1 9 1 11 2 15 15 13 1 9 12 9 2
26 0 9 1 9 1 9 15 4 11 13 1 9 13 11 9 9 1 9 9 16 9 14 13 15 9 2
30 1 9 1 11 1 9 1 11 2 9 11 1 9 11 11 13 4 16 4 11 13 13 16 14 13 1 9 0 9 2
37 2 3 4 0 7 0 9 11 13 15 1 9 2 1 11 2 2 3 16 4 1 9 9 0 9 1 9 7 9 1 9 2 2 13 4 11 2
11 11 4 1 9 1 9 9 13 0 9 2
18 2 15 9 2 15 9 13 4 0 9 1 9 9 2 2 13 4 2
49 2 0 1 11 4 15 13 4 14 9 1 0 9 2 1 0 0 9 15 4 13 2 3 13 1 0 9 2 13 9 9 9 0 1 9 9 0 1 9 11 2 2 13 11 0 0 9 11 2
19 7 0 7 0 9 13 4 2 16 15 13 2 0 9 16 14 13 9 2
37 2 13 9 13 15 1 0 9 1 9 1 11 7 13 9 0 9 2 2 13 4 9 0 0 9 2 0 9 0 9 11 11 2 7 13 11 2
28 1 9 2 11 4 1 9 13 9 1 9 1 9 2 9 1 15 4 0 9 13 15 0 9 1 9 9 2
20 1 9 9 15 4 9 13 0 2 9 4 0 9 13 9 9 1 0 9 2
9 9 0 1 9 1 0 9 1 11
29 15 3 3 4 13 9 1 12 0 9 1 0 9 1 11 2 7 15 15 13 1 0 9 15 13 1 9 11 2
14 0 9 7 0 9 11 13 4 16 4 9 9 0 2
23 0 9 13 4 9 1 9 0 9 1 11 1 15 4 1 9 2 12 9 2 13 9 2
12 12 0 9 1 0 9 1 11 13 4 9 2
22 0 9 1 0 9 1 9 11 2 1 9 11 2 0 4 12 9 1 0 0 9 2
15 12 9 4 13 16 4 0 13 9 0 12 9 1 9 2
26 12 9 3 2 3 12 2 12 3 2 0 9 13 4 9 1 0 9 1 11 11 1 9 9 11 2
8 1 9 4 3 0 0 9 2
9 7 1 12 1 9 4 4 9 2
26 0 9 7 11 2 0 9 11 1 11 2 13 4 9 16 0 2 3 16 15 14 13 13 0 9 2
38 2 9 1 0 9 1 9 11 13 9 12 0 9 2 15 4 3 9 15 1 0 0 9 15 13 1 9 7 1 11 2 2 13 4 9 11 11 2
38 12 0 9 2 9 9 15 15 13 9 0 9 1 0 9 2 7 0 9 9 1 9 11 3 15 9 2 3 4 13 0 9 9 2 13 4 11 2
16 0 13 16 9 3 13 1 9 9 9 11 1 11 7 11 2
46 1 9 1 11 11 13 4 3 9 1 9 0 9 0 9 1 15 15 13 1 9 1 9 11 2 1 15 9 3 3 9 14 13 13 9 1 9 3 0 0 9 15 13 11 11 2
29 9 4 13 3 9 1 9 11 2 7 9 13 13 9 1 15 9 1 9 9 9 9 7 9 9 1 0 9 2
29 9 0 9 13 4 9 16 3 13 9 7 9 1 11 2 7 9 13 16 4 9 9 1 11 7 15 0 9 2
11 3 2 9 1 9 9 3 13 4 0 2
23 1 9 2 0 0 9 1 11 2 1 0 9 11 11 11 2 13 4 9 3 0 9 2
24 11 11 2 9 0 9 1 9 2 13 4 11 1 0 9 2 3 16 4 3 13 0 9 2
8 9 11 16 13 0 9 13 9
17 1 0 9 15 9 2 0 9 13 0 9 9 9 9 1 9 2
42 9 0 1 9 13 15 1 9 2 1 9 0 11 2 7 3 13 0 0 1 9 9 9 1 9 2 15 15 9 13 1 9 15 4 4 0 1 0 0 9 11 2
19 15 4 9 11 13 12 9 9 1 9 9 1 9 7 9 1 15 9 2
15 9 9 13 16 4 15 13 9 9 7 13 9 1 11 2
10 3 2 1 9 4 15 9 1 9 2
20 9 1 15 4 15 13 9 13 2 9 2 11 7 3 4 0 9 15 9 2
24 2 1 0 9 2 15 4 9 13 0 2 2 13 4 1 11 11 11 2 9 1 9 0 2
31 2 9 4 1 15 15 15 2 9 2 13 12 9 2 0 9 11 2 13 9 3 0 9 2 9 9 2 2 13 4 2
21 7 0 0 11 0 9 2 11 2 3 15 3 13 9 9 7 9 9 1 9 2
31 11 13 16 15 9 9 1 9 13 1 9 0 0 9 2 7 14 1 9 7 1 9 9 2 16 15 15 13 13 9 2
58 2 1 9 1 9 7 9 0 0 9 2 9 9 1 9 13 0 0 9 2 15 13 16 4 9 1 9 9 9 1 9 3 0 9 1 9 9 7 9 2 2 13 4 1 11 11 11 2 9 11 7 9 0 9 1 9 9 2
20 2 0 15 0 9 7 9 13 7 1 0 7 1 0 9 2 2 13 4 2
15 2 15 15 9 13 1 0 9 0 9 2 2 2 2 2
22 13 4 0 16 2 1 9 9 15 0 9 2 4 13 1 9 9 2 2 2 2 2
17 3 3 13 16 15 9 9 1 9 13 1 9 9 7 9 2 2
45 2 15 4 15 9 13 13 3 1 15 13 9 0 9 2 9 9 9 2 7 0 9 15 4 15 9 13 2 1 15 9 13 15 9 7 1 15 15 13 9 2 2 13 4 2
25 2 13 9 0 0 9 1 15 9 2 0 9 1 11 2 9 15 13 4 7 9 1 9 9 2
30 3 1 15 9 13 13 9 9 1 9 7 2 4 14 0 1 9 2 3 3 13 13 1 9 2 2 13 4 11 2
43 1 9 16 13 15 9 1 11 2 11 4 1 9 9 1 11 13 16 9 2 1 9 13 9 1 0 9 7 9 15 9 1 9 7 9 9 1 9 9 15 9 2 2
34 15 4 9 1 9 12 9 13 9 1 9 0 9 9 1 11 2 7 13 16 4 1 0 9 1 15 9 13 1 0 9 15 9 2
29 11 4 1 12 7 12 9 13 9 1 9 7 9 9 9 1 9 1 12 9 9 9 1 11 2 11 7 11 2
17 13 15 16 15 1 11 13 15 1 0 9 9 1 9 1 11 2
20 0 9 9 1 9 1 9 2 14 3 11 2 13 15 1 12 9 0 9 2
25 3 1 11 2 3 3 0 9 13 0 9 1 11 2 11 2 11 2 11 2 11 7 0 11 2
26 3 2 11 2 1 15 15 13 16 13 0 9 9 1 9 2 13 4 9 3 16 9 9 1 9 2
7 14 0 9 1 9 1 11
17 0 9 0 4 1 9 16 13 0 9 9 1 9 0 0 9 2
35 16 15 9 1 12 9 13 1 0 0 7 0 9 2 0 4 9 2 3 0 0 9 1 11 2 1 12 9 9 11 13 0 9 9 2
18 15 15 13 1 9 13 15 0 9 9 1 9 0 0 9 11 11 2
19 2 14 13 13 9 15 13 9 9 2 2 13 4 9 0 9 11 11 2
24 9 4 13 0 9 2 7 9 9 13 4 9 1 15 15 1 9 13 16 13 4 15 9 2
11 2 9 4 9 11 11 2 2 2 2 2
22 0 4 11 13 1 15 9 2 3 7 15 2 2 13 4 11 11 2 0 0 9 2
35 9 4 1 0 12 9 13 9 9 2 3 15 13 3 0 9 7 9 9 2 7 0 0 9 9 8 8 13 9 7 1 9 1 9 2
34 3 4 0 9 13 15 0 9 9 9 2 14 1 15 15 13 0 9 2 3 3 15 13 16 4 9 3 3 3 13 1 0 9 2
14 12 15 1 9 13 7 4 13 9 9 1 15 9 2
17 2 14 13 13 16 4 9 3 0 0 7 0 9 13 4 0 2
16 15 4 12 1 0 9 1 11 2 2 13 4 9 11 11 2
16 9 15 13 9 0 4 9 15 14 13 16 4 4 0 9 2
35 11 11 2 9 9 11 2 1 11 13 16 4 9 4 0 0 9 1 15 4 9 2 3 0 2 13 15 9 1 9 2 9 7 9 2
14 2 1 0 9 9 9 13 9 3 0 0 9 2 2
22 2 15 4 9 9 7 9 0 9 7 0 9 2 2 13 4 9 11 11 1 11 2
27 2 4 9 1 15 16 13 12 0 9 15 13 16 9 14 4 13 13 2 16 0 13 16 15 13 13 2
25 3 4 9 1 9 15 13 2 13 14 15 9 2 2 13 4 1 11 11 11 2 0 9 11 2
7 9 13 9 9 9 1 11
18 0 13 9 3 4 9 9 1 9 1 9 9 0 9 7 0 9 2
25 0 9 13 9 3 15 15 9 1 0 9 1 9 9 12 9 13 1 9 1 9 7 9 9 2
25 9 2 15 4 3 0 2 13 4 1 9 0 9 2 3 0 0 9 9 0 9 0 0 9 2
18 9 4 15 13 15 2 16 4 15 2 16 13 2 13 1 0 9 2
38 9 4 13 1 11 2 16 9 11 11 2 9 0 9 7 9 0 9 11 2 15 4 2 1 15 9 2 3 13 9 1 9 0 9 1 9 9 2
30 3 2 0 9 13 4 15 1 9 16 4 15 15 13 0 9 3 1 9 15 15 15 15 13 9 1 9 13 9 2
32 9 0 9 3 4 15 13 0 7 13 9 0 9 2 9 9 2 9 1 0 9 2 9 1 9 2 7 13 0 9 9 2
34 2 11 14 13 13 2 2 13 4 12 1 9 2 15 15 13 3 16 11 7 13 16 4 9 16 4 9 13 13 0 9 4 9 2
20 2 15 4 4 3 0 2 16 4 2 9 2 2 9 2 13 7 13 9 2
30 1 15 2 0 9 9 13 4 16 15 9 9 14 13 15 9 9 7 9 9 1 15 4 0 2 2 13 4 11 2
9 11 11 13 4 13 9 9 9 2
38 2 15 4 13 2 11 2 2 9 7 9 2 9 2 9 2 9 2 2 0 9 9 9 2 11 11 2 0 15 13 1 9 2 9 1 9 2 2
16 2 3 4 13 2 3 2 4 7 3 13 2 2 13 4 2
20 0 9 2 11 2 13 15 7 13 16 4 0 7 3 0 9 13 0 9 2
19 2 9 2 9 2 2 2 0 7 14 2 15 9 0 4 1 0 9 2
29 15 4 13 9 1 9 7 13 9 1 9 2 7 0 9 13 1 9 16 4 0 9 13 13 1 0 9 2 2
18 15 0 9 15 9 4 4 0 1 9 1 9 0 9 2 13 11 2
36 0 9 2 11 2 13 4 15 1 9 15 4 13 9 9 2 3 3 16 15 4 3 15 9 15 4 7 3 1 9 16 4 13 0 9 2
8 2 9 15 4 13 1 15 2
27 9 15 4 15 1 9 2 7 7 1 0 9 2 0 1 15 15 15 3 13 1 11 7 1 0 9 2
12 1 15 9 4 15 13 13 2 2 13 4 2
13 1 9 9 7 9 2 11 13 9 1 0 9 2
8 2 3 4 15 9 13 9 2
18 13 4 9 9 2 13 4 15 16 4 3 3 7 16 15 13 13 2
8 0 9 0 4 1 9 9 2
13 15 4 9 3 1 3 0 9 2 2 13 4 2
6 11 11 15 13 1 11
22 1 9 0 1 9 2 0 9 7 9 11 11 13 15 9 7 13 15 9 0 9 2
27 11 11 2 0 9 2 9 7 12 1 0 9 0 9 2 13 15 1 11 12 9 1 12 9 1 9 2
22 9 11 2 9 11 7 9 9 7 9 11 2 13 9 1 9 11 1 15 0 9 2
26 11 2 9 7 0 0 9 0 0 9 2 13 4 1 11 1 9 12 9 2 1 0 9 12 9 2
22 1 11 4 0 1 15 0 9 7 9 2 7 13 9 1 11 2 3 1 3 13 2
21 9 0 9 2 3 9 11 11 11 2 13 4 11 1 9 7 13 15 0 9 2
44 0 1 15 0 9 0 9 7 16 9 0 9 11 2 11 13 13 9 1 0 9 2 14 16 0 9 2 3 16 0 9 15 15 13 1 0 7 0 9 9 11 1 11 2
24 3 2 11 7 3 13 0 9 11 2 15 15 13 1 9 2 7 3 4 0 1 0 9 2
28 3 1 11 2 9 9 11 11 11 13 16 4 11 4 0 9 1 0 9 2 16 13 4 3 9 9 11 2
27 1 11 2 2 11 4 2 16 9 15 13 9 2 13 1 0 0 9 1 11 15 15 13 1 9 2 2
43 11 11 1 0 9 0 9 0 9 13 16 2 0 9 1 11 2 7 0 1 11 2 2 3 16 4 0 2 0 7 0 9 11 2 16 3 0 2 13 9 15 9 2
24 11 4 13 0 9 1 11 2 3 9 15 9 16 2 9 9 0 1 0 9 0 9 2 2
26 2 13 13 15 15 13 9 15 9 2 7 15 15 13 13 15 0 9 13 4 13 2 2 13 4 2
27 11 4 13 0 0 9 1 9 2 0 9 2 0 9 2 15 4 3 13 1 15 9 3 3 12 9 2
20 13 15 3 4 13 2 0 9 2 1 9 16 13 9 1 9 0 9 11 2
32 0 0 9 1 0 0 0 9 9 11 8 11 13 9 3 4 3 11 13 1 9 2 0 9 2 1 15 9 1 12 9 2
36 1 9 3 15 3 13 1 2 0 9 2 7 2 9 1 9 0 9 2 2 9 11 11 1 9 11 13 16 4 9 9 1 11 0 9 2
30 2 13 15 1 9 9 7 9 2 7 9 1 11 13 15 13 1 15 9 1 15 4 13 2 2 13 4 1 11 2
23 9 11 11 2 9 0 9 1 9 2 13 15 16 4 1 0 9 13 1 3 0 9 2
33 2 3 4 9 1 0 9 4 0 13 1 9 2 7 9 9 9 13 15 1 9 9 0 9 1 11 2 2 13 11 1 11 2
28 3 2 1 9 1 0 9 1 0 9 2 13 9 3 4 0 9 11 7 13 14 4 1 9 13 15 9 2
32 0 9 0 9 2 11 2 15 13 11 2 13 15 4 16 15 15 13 2 16 1 11 7 0 0 0 9 7 3 13 9 2
31 11 11 11 1 9 1 0 9 13 16 3 13 13 0 9 1 0 9 2 7 13 3 0 16 4 11 13 9 1 11 2
33 2 16 15 14 13 2 15 4 0 9 3 0 7 9 4 15 15 1 0 9 13 1 9 0 0 9 2 2 13 4 1 11 2
6 0 9 2 9 13 11
11 9 9 13 15 1 11 13 9 11 12 2
27 3 1 0 9 2 0 9 11 13 15 1 9 11 2 7 0 9 0 9 11 13 9 11 0 1 11 2
8 11 4 4 9 9 11 12 2
19 9 11 12 13 4 1 0 9 11 15 4 13 1 9 2 12 9 2 2
23 13 4 9 16 15 9 13 13 2 3 16 4 1 15 9 4 9 2 0 9 2 9 2
26 9 11 11 13 15 1 11 1 9 7 13 0 9 16 13 9 1 11 16 13 15 9 0 9 9 2
32 0 9 11 11 13 15 1 9 2 12 9 2 1 9 0 9 11 7 11 2 11 2 16 4 13 1 0 9 7 0 9 2
9 11 4 13 9 11 0 9 11 2
32 13 4 16 4 3 9 4 0 9 11 9 7 9 9 11 2 3 15 16 9 1 9 1 0 9 7 9 9 15 1 15 2
45 11 4 1 9 11 7 9 9 13 4 4 0 1 9 15 9 7 9 12 9 2 13 4 1 9 2 12 9 2 0 9 0 9 11 11 11 2 15 9 4 0 0 9 11 2
31 11 4 13 0 0 0 9 1 0 9 7 13 0 9 9 1 9 15 9 2 13 4 0 9 11 11 1 9 1 11 2
23 11 4 13 1 11 1 11 7 11 2 3 4 13 1 9 11 2 0 11 1 0 9 2
21 0 9 11 11 13 15 1 9 2 12 9 2 1 11 1 15 0 9 11 11 2
10 13 4 1 0 9 1 9 0 9 2
20 1 9 0 9 2 11 15 3 13 1 9 11 11 7 0 0 7 0 9 2
27 0 9 9 11 11 7 15 0 9 11 11 13 4 1 9 2 12 9 2 1 11 0 9 1 0 9 2
10 11 15 1 9 13 1 9 11 11 2
6 9 13 0 9 1 11
22 13 15 16 1 9 1 0 9 1 11 1 15 4 13 1 9 3 3 13 0 9 2
16 9 9 1 9 9 13 9 1 9 1 9 0 9 1 11 2
17 1 0 9 1 9 1 9 0 4 0 9 2 7 0 4 4 2
22 0 9 13 4 9 0 9 1 11 3 9 1 9 0 9 1 9 2 12 9 2 2
26 9 2 0 16 0 9 1 9 0 9 1 0 3 12 9 2 13 15 0 9 15 15 13 0 9 2
36 2 0 9 0 4 1 12 2 12 3 2 12 11 2 1 0 9 2 3 0 9 1 0 9 7 9 2 2 13 15 1 9 9 0 9 2
34 0 9 2 3 15 13 2 13 1 9 0 9 2 3 9 9 0 9 9 11 11 1 9 0 9 7 9 1 9 9 3 12 9 2
35 15 9 13 4 0 0 9 1 11 1 3 4 0 0 9 12 9 2 15 4 13 0 9 9 1 12 9 2 3 16 4 0 7 0 2
22 1 9 12 9 3 4 9 0 9 2 0 0 9 16 9 0 9 0 9 11 11 2
36 3 16 15 4 0 1 2 3 0 9 2 1 9 3 2 0 9 1 11 11 11 13 4 16 14 13 13 2 9 1 15 0 9 9 2 2
30 9 0 9 2 15 15 13 1 0 12 9 1 9 11 7 0 4 0 9 2 12 4 1 0 9 1 0 9 11 2
29 1 0 9 0 4 16 4 9 13 9 1 9 0 9 7 13 1 9 1 0 9 2 3 15 3 13 9 9 2
18 9 4 13 16 4 0 12 7 12 9 2 7 4 0 9 1 9 2
10 1 9 4 3 0 9 1 0 9 2
21 3 1 9 2 12 0 9 13 4 9 1 9 9 2 3 9 0 9 7 9 2
19 0 9 11 13 4 16 4 9 13 0 9 7 0 9 1 9 1 9 2
11 11 4 13 9 1 9 3 7 13 9 2
29 2 9 16 15 4 15 3 4 13 2 11 2 1 0 2 0 9 7 1 9 9 2 2 13 4 9 0 9 2
26 2 11 9 0 4 13 0 9 2 15 4 13 7 1 9 2 16 15 14 4 13 9 15 9 2 2
27 1 9 12 9 9 15 13 1 9 0 0 9 15 4 13 0 9 1 12 0 9 7 3 0 9 2 2
7 11 15 13 0 9 1 9
22 0 9 1 11 13 4 1 0 9 11 1 15 4 0 0 9 9 1 9 0 9 2
10 9 9 11 13 4 1 0 9 9 2
22 1 11 4 12 9 0 0 9 2 9 0 9 2 9 7 9 15 13 0 9 11 2
9 9 4 0 12 9 9 9 9 2
8 9 9 4 4 9 0 11 2
21 9 0 9 7 0 9 13 4 9 15 15 0 9 13 1 9 1 9 9 9 2
23 9 9 4 15 13 1 9 0 9 15 4 13 1 9 2 3 0 2 0 7 0 9 2
19 2 0 9 2 13 15 15 9 7 0 9 2 13 4 0 7 13 13 2
15 15 0 9 4 0 2 0 2 0 7 0 9 0 9 2
8 9 15 9 4 9 9 9 2
31 9 9 4 9 9 15 14 13 9 2 7 0 9 15 0 13 13 2 2 13 4 9 9 11 11 11 1 9 9 9 2
22 9 9 0 4 1 9 9 0 11 2 1 0 9 16 4 1 9 0 9 0 9 2
12 11 4 13 16 9 4 13 4 15 0 9 2
9 9 1 9 9 4 13 9 9 2
14 0 9 4 0 1 0 7 0 9 1 9 7 9 2
22 1 0 9 13 15 12 0 9 2 15 13 12 9 1 9 2 11 2 11 7 11 2
7 9 3 13 9 9 11 2
7 9 1 0 9 4 0 2
22 9 0 9 11 2 11 2 13 4 1 9 2 3 16 15 15 9 11 13 9 9 2
16 11 4 13 16 4 9 4 0 16 4 0 7 13 9 9 2
17 11 2 4 3 0 9 2 2 13 11 11 2 9 9 0 11 2
17 15 13 2 9 7 9 0 9 0 9 11 2 2 13 4 11 2
30 9 4 1 9 3 13 9 15 15 9 15 4 4 0 13 9 1 9 1 12 7 12 9 13 1 9 1 15 9 2
12 9 4 3 13 0 9 0 9 9 7 9 2
9 11 11 13 9 9 1 9 1 11
25 11 2 11 2 9 11 13 4 1 9 2 12 9 2 3 13 11 11 9 9 1 9 1 11 2
34 0 9 2 11 2 13 4 9 9 16 15 15 13 2 7 4 3 13 15 0 9 15 4 0 13 9 1 9 1 0 9 1 11 2
20 1 15 9 4 9 9 2 9 9 7 0 9 7 9 1 0 9 7 9 2
17 15 9 1 9 13 4 9 16 4 15 9 11 11 13 3 13 2
12 0 9 2 0 11 13 4 12 0 9 1 11
10 11 13 12 0 9 1 0 0 9 2
26 3 1 0 9 2 0 9 1 11 7 0 0 9 1 11 13 4 9 2 7 11 9 0 9 9 2
27 0 0 9 11 13 13 12 0 0 9 1 11 1 12 9 2 13 4 1 9 2 12 9 2 0 9 2
36 9 4 1 3 1 15 9 13 3 12 9 9 1 11 2 7 1 12 9 13 13 9 0 9 9 2 1 9 1 3 12 9 1 15 9 2
31 11 4 9 0 9 9 1 15 4 0 9 9 1 9 9 7 9 9 1 9 2 9 1 9 9 7 0 9 1 9 2
11 9 13 1 9 2 12 9 2 1 9 2
16 11 4 0 9 9 15 9 2 1 9 9 11 7 11 11 2
39 0 9 1 11 7 0 0 9 1 11 13 4 1 9 2 12 9 2 9 1 9 2 1 9 9 9 1 0 9 9 7 9 7 9 9 1 9 9 2
26 0 0 0 0 9 11 13 4 3 0 1 9 2 12 9 2 2 15 4 0 9 9 1 0 9 2
18 0 0 9 13 9 9 12 0 9 7 13 4 13 12 9 9 3 2
21 9 9 13 3 12 9 9 7 13 9 2 11 9 7 3 0 9 1 0 9 2
17 0 9 11 11 13 4 9 1 9 0 9 1 11 2 1 11 2
17 0 0 9 1 9 11 11 13 4 9 1 0 0 9 12 9 2
6 9 4 13 12 9 2
16 0 0 9 16 15 4 11 7 11 15 4 1 9 11 11 2
24 0 9 13 4 9 1 12 9 1 9 1 9 1 9 12 2 1 9 1 0 9 0 9 2
17 0 9 9 13 4 9 1 12 9 9 1 0 12 9 15 9 2
7 11 15 13 1 0 0 9
23 0 9 7 0 9 13 16 4 0 9 2 9 1 9 11 7 0 9 2 13 13 9 2
21 9 15 4 13 1 9 1 0 9 11 0 4 9 0 9 2 1 3 0 9 2
26 0 9 9 11 11 13 16 4 15 15 15 13 1 9 13 13 14 3 0 0 9 2 3 7 9 2
33 2 13 15 16 4 2 3 4 1 9 9 1 9 11 2 15 13 4 9 1 9 3 9 2 2 13 4 11 9 11 9 9 2
25 0 13 14 9 11 13 11 2 11 4 13 16 4 9 11 16 15 1 11 13 0 7 0 9 2
18 9 0 9 11 11 13 15 16 9 1 0 3 9 13 0 0 9 2
24 1 9 1 15 2 1 11 4 13 16 4 9 11 1 0 9 15 15 13 13 1 0 9 2
11 2 9 0 7 0 0 9 13 4 0 2
11 11 4 0 9 7 3 1 15 13 13 2
22 13 15 16 4 0 9 7 9 11 1 11 1 0 9 13 1 15 2 2 13 4 2
8 13 0 9 16 3 0 9 2
37 2 0 9 14 13 13 16 9 1 0 0 9 7 1 15 9 2 2 13 4 11 2 3 16 0 9 14 13 9 7 3 13 0 9 1 11 2
23 11 11 2 9 1 0 9 1 0 9 2 14 13 16 9 11 13 1 0 9 1 11 2
21 2 0 9 3 14 13 15 7 14 13 16 4 9 7 9 13 1 9 1 11 2
27 9 4 13 1 0 9 1 9 11 12 9 7 14 13 16 4 15 13 3 2 2 13 4 11 1 11 2
27 13 16 2 1 0 9 1 9 11 2 13 7 0 2 3 0 9 2 0 9 2 3 9 9 7 9 2
18 2 14 13 0 9 1 0 7 0 9 2 0 9 13 15 1 11 2
16 15 13 0 9 16 15 3 13 7 13 2 1 9 1 9 2
24 3 4 1 11 0 9 9 9 2 7 1 0 4 4 7 11 7 11 2 2 13 4 11 2
17 3 12 0 0 9 1 11 2 13 4 1 11 2 4 0 9 2
13 2 9 9 15 13 12 9 3 4 0 0 9 2
26 3 4 13 9 9 7 0 9 13 16 4 0 13 1 0 9 2 7 3 7 9 2 2 13 4 2
11 0 9 11 13 1 0 9 1 9 1 9
41 0 9 13 4 13 9 1 11 16 15 13 1 9 9 9 16 15 13 15 9 1 0 9 2 13 4 1 9 9 11 11 2 1 0 9 1 9 0 9 11 2
5 0 9 11 11 2
45 0 9 11 11 13 4 1 9 2 12 9 2 0 9 1 0 9 11 1 0 9 1 11 1 9 16 15 1 15 13 9 4 15 0 1 9 7 9 1 9 9 1 0 9 2
35 2 15 9 15 14 13 9 11 0 4 2 2 13 4 11 2 3 3 16 4 15 9 1 9 9 1 0 9 13 13 11 1 9 9 2
22 2 1 4 15 9 1 15 15 13 15 9 13 4 15 9 7 15 9 1 15 9 2
46 16 13 3 13 9 15 13 3 4 15 0 15 13 2 2 13 4 11 1 9 1 9 11 11 2 9 9 0 9 11 1 11 2 1 15 4 0 1 0 9 7 9 9 9 11 2
57 0 9 4 4 0 1 9 0 9 9 15 13 11 2 11 2 11 2 11 2 11 7 0 9 2 7 15 4 13 9 9 2 0 9 1 11 11 11 2 0 9 11 11 7 11 11 11 15 13 11 2 1 9 1 15 9 2
33 11 4 4 3 0 1 9 1 9 11 0 1 9 15 4 13 11 2 7 15 4 13 3 1 9 9 7 3 4 13 15 9 2
10 11 4 0 9 13 9 9 16 9 2
25 2 9 9 13 4 0 9 2 2 2 16 13 9 11 2 2 13 4 11 1 9 9 0 11 2
22 2 3 4 13 15 9 2 13 16 4 15 3 0 9 7 13 4 13 15 15 2 2
35 0 9 9 13 13 1 9 2 3 4 9 9 9 13 1 11 2 3 4 15 13 1 0 9 2 7 3 1 9 13 0 9 1 11 2
23 1 9 2 9 15 1 9 1 11 13 1 9 12 9 9 9 1 15 4 13 9 9 2
15 2 15 4 0 9 2 2 13 4 9 0 9 0 9 2
15 2 9 4 9 9 15 0 9 7 9 1 9 9 2 2
33 9 9 9 11 0 4 0 9 1 9 9 2 1 15 4 0 9 13 9 9 9 9 11 1 11 1 9 11 16 4 13 9 2
29 0 11 15 13 12 9 1 3 12 9 9 9 13 4 9 2 16 14 4 3 13 0 9 1 11 15 4 13 2
14 3 2 9 7 9 1 9 13 4 9 1 0 9 2
20 0 0 9 0 11 13 4 1 9 1 0 0 9 1 9 7 0 0 9 2
26 2 13 4 0 16 15 1 9 13 9 2 2 13 4 9 9 11 11 11 0 9 11 2 13 11 2
11 2 9 11 13 9 13 9 1 15 9 2
10 13 9 16 4 13 0 1 9 11 2
37 14 3 3 4 1 9 9 2 12 2 12 2 2 9 7 9 2 16 0 15 4 13 1 0 12 9 2 2 2 3 16 4 13 9 9 2 2
7 0 9 11 14 13 0 9
18 0 9 13 4 13 0 9 2 15 4 13 15 9 0 1 0 9 2
7 3 2 9 3 13 9 2
10 9 0 9 11 11 11 13 13 9 2
15 3 9 13 15 0 9 1 9 0 9 1 9 1 9 2
18 12 9 13 13 0 9 15 4 13 11 13 1 9 7 13 0 9 2
12 0 2 0 9 9 2 13 9 0 9 9 2
21 1 9 2 0 9 13 4 9 9 2 16 4 15 15 13 13 9 0 1 9 2
14 9 15 15 13 1 9 9 3 4 1 0 13 9 2
18 9 9 0 9 3 4 13 2 3 9 1 12 9 1 9 12 9 2
12 16 4 9 7 9 13 2 9 4 4 0 2
19 9 4 13 16 4 0 9 13 13 9 7 15 13 9 3 0 0 9 2
17 0 1 3 0 9 2 15 9 13 9 9 16 15 9 14 13 2
14 9 9 2 9 15 13 1 0 9 1 3 12 9 2
9 3 2 9 7 15 9 4 0 2
10 13 4 16 0 9 3 13 9 9 2
15 11 11 2 9 0 9 2 14 13 9 1 9 0 9 2
31 15 15 4 3 13 4 9 2 13 11 2 4 9 0 9 1 0 7 0 9 2 15 4 13 0 9 7 0 0 9 2
20 9 0 9 11 7 9 11 11 2 15 4 9 13 0 0 9 2 4 0 2
8 0 9 0 9 0 4 9 2
30 9 13 16 9 2 16 13 13 9 2 13 13 9 2 13 9 9 7 0 9 2 7 14 13 15 9 1 0 9 2
11 13 15 16 0 9 13 1 9 0 9 2
20 1 9 2 0 9 13 15 1 9 15 4 9 13 3 0 2 7 9 13 2
24 1 0 12 9 15 9 2 9 4 13 1 12 9 2 16 4 9 3 13 9 1 12 9 2
19 1 9 15 4 15 3 13 4 9 2 9 2 0 9 2 9 7 9 2
17 1 9 4 13 9 2 0 9 2 9 2 9 2 9 7 9 2
15 0 9 14 13 9 16 0 9 15 15 13 0 0 9 2
17 13 16 4 9 3 0 1 0 9 2 9 9 7 9 1 9 2
20 0 0 9 7 3 4 0 2 1 9 1 12 9 1 0 3 9 15 9 2
16 0 9 2 1 9 1 9 9 1 0 9 13 4 15 9 2
29 3 0 2 13 0 9 2 9 0 9 4 0 2 16 4 3 9 13 9 9 0 9 7 3 13 1 0 9 2
16 11 15 3 3 13 3 4 1 9 13 0 9 1 15 9 2
9 3 4 15 15 13 9 15 9 2
5 11 13 9 11 9
14 9 13 0 9 1 0 15 4 0 13 0 0 9 2
12 3 2 9 15 13 1 9 9 7 0 9 2
15 13 9 9 9 1 11 2 7 0 9 7 3 13 9 2
27 11 15 4 0 13 15 0 9 13 13 0 9 1 9 0 0 9 1 9 2 11 2 9 0 9 2 2
14 0 9 9 3 4 13 12 9 0 0 9 7 9 2
11 9 15 13 12 9 3 7 13 9 9 2
15 9 15 13 9 9 1 11 2 11 2 11 7 1 9 2
27 2 9 15 11 9 9 4 9 9 11 2 0 9 2 8 9 7 9 2 2 13 4 9 9 11 11 2
33 2 0 4 7 13 0 9 1 9 2 7 4 15 3 0 2 16 13 9 9 3 1 9 9 2 2 13 11 2 9 1 11 2
19 3 12 9 15 9 13 1 0 9 2 16 0 13 1 0 9 3 11 2
11 12 9 13 15 9 2 3 7 11 9 2
13 9 15 13 1 9 11 9 7 0 9 1 9 2
11 1 9 2 9 3 13 9 0 9 9 2
9 11 4 13 3 4 13 9 9 2
16 15 9 15 15 13 1 9 1 9 9 13 15 1 9 9 2
33 1 15 2 9 15 13 1 9 16 13 11 9 1 0 9 2 3 2 9 1 0 9 9 4 9 8 2 8 2 2 13 2 2
21 3 0 9 15 4 13 11 2 7 13 8 9 2 13 4 9 9 9 1 11 2
14 1 9 1 0 9 2 9 9 0 4 1 12 9 2
33 3 2 0 9 0 9 7 0 9 9 9 13 0 9 2 7 3 12 9 9 13 4 0 9 16 9 15 15 13 1 9 9 2
9 0 9 1 11 2 13 9 1 9
28 0 9 1 11 7 11 13 4 3 9 13 16 9 16 15 4 0 9 1 9 0 0 9 4 0 0 9 2
43 12 9 1 0 9 1 9 0 0 9 1 11 2 0 9 0 9 11 2 11 2 13 3 13 15 9 7 13 9 16 4 0 9 3 13 9 7 9 15 13 1 9 2
31 2 9 2 9 7 9 14 13 13 0 9 7 9 2 7 16 15 15 9 3 13 2 3 15 13 0 7 0 9 9 2
16 9 1 9 9 9 4 1 9 2 2 13 15 1 9 11 2
33 3 16 15 11 3 13 9 0 9 9 2 9 7 9 2 0 15 13 16 15 15 9 13 13 1 9 1 15 0 9 13 9 2
22 16 4 11 13 0 9 9 3 1 9 12 9 2 0 9 9 7 3 4 0 9 2
26 2 9 15 14 13 1 0 9 9 4 15 9 7 14 13 0 9 9 0 9 2 13 9 0 9 2
37 16 4 15 3 2 4 3 13 0 0 9 2 7 15 4 0 1 11 2 15 7 1 9 13 3 0 9 2 2 13 1 11 9 11 11 11 2
37 2 9 4 7 13 15 15 2 7 9 0 9 14 13 3 4 0 1 9 2 16 4 15 9 1 9 2 2 13 4 1 11 9 11 11 11 2
25 9 13 16 4 4 15 0 9 9 0 9 9 13 1 9 16 9 2 9 4 1 9 7 9 2
36 9 9 11 9 11 11 16 13 9 0 9 7 0 9 1 11 7 1 9 2 15 15 13 9 7 9 1 9 9 2 3 4 15 0 9 2
19 0 9 0 4 1 9 1 9 0 9 2 9 1 0 0 9 11 11 2
27 2 9 16 15 9 7 9 13 1 9 7 0 9 13 15 9 0 7 0 2 16 13 13 15 0 9 2
29 13 16 1 11 1 9 7 1 9 13 0 2 0 7 0 9 7 9 15 7 15 9 2 2 13 15 1 9 2
35 2 15 13 9 7 9 1 15 15 3 13 2 0 3 1 9 9 2 3 9 7 15 9 1 9 0 9 9 2 2 13 15 1 9 2
13 9 0 9 2 9 11 11 2 13 4 0 9 2
21 2 9 15 13 3 0 9 7 13 15 0 0 9 13 9 2 2 13 4 11 2
26 11 11 2 0 9 0 9 11 0 11 2 3 4 13 9 1 9 7 13 9 16 15 13 0 9 2
33 2 15 9 13 16 1 9 13 9 15 0 9 2 7 13 4 13 1 15 14 16 4 15 15 13 9 16 9 3 15 13 9 2
26 13 15 1 15 9 7 9 2 11 2 15 3 4 13 9 3 15 13 1 9 2 2 13 4 11 2
9 9 1 9 9 1 11 13 15 9
19 9 11 11 13 16 9 13 15 9 9 1 0 9 11 7 13 0 9 2
32 9 11 11 2 0 9 12 9 3 1 11 2 1 9 1 11 7 11 2 13 4 0 9 9 3 16 9 9 13 15 9 2
26 9 4 13 1 15 4 9 13 16 4 11 11 2 0 11 2 3 1 9 9 13 9 1 0 11 2
45 3 2 13 12 9 9 1 11 2 11 2 11 7 0 0 7 0 9 15 13 1 9 1 9 1 11 11 2 7 0 0 9 13 16 4 3 1 15 9 15 3 13 1 9 2
31 2 13 15 3 2 1 9 4 7 3 7 3 7 14 13 15 4 15 9 2 2 13 4 1 11 9 15 9 11 11 2
20 9 1 9 13 3 9 7 1 15 4 4 0 9 9 1 9 1 0 11 2
29 1 0 12 9 2 3 2 13 14 0 9 9 1 11 7 11 15 13 1 9 7 9 7 13 13 1 0 9 2
38 2 13 4 9 0 9 16 15 13 1 9 1 0 9 9 2 7 15 4 13 4 15 16 4 15 13 2 2 13 4 1 11 9 9 11 11 11 2
14 11 11 4 0 9 1 3 0 9 7 13 12 9 2
12 1 9 9 1 9 1 9 13 4 12 9 2
22 2 11 4 0 1 3 9 2 2 13 4 1 11 11 11 2 9 0 9 1 9 2
29 11 4 13 16 4 3 0 0 9 1 9 1 11 2 16 15 9 9 9 1 11 13 12 9 1 0 12 9 2
31 2 13 16 15 9 15 13 9 13 1 0 9 11 7 2 1 2 9 0 9 2 2 13 4 1 11 9 11 11 11 2
17 0 9 14 13 15 9 16 13 1 9 2 16 13 1 15 9 2
16 1 3 12 9 1 0 9 1 15 9 2 3 12 13 9 2
25 9 9 1 9 13 4 16 9 1 11 11 4 4 0 2 7 16 9 13 1 9 1 9 0 2
30 2 13 4 1 9 9 16 13 15 0 9 15 4 13 1 9 1 9 2 2 13 4 1 11 9 1 9 11 11 2
26 11 13 16 15 1 9 1 11 11 13 13 0 9 2 1 15 4 9 9 13 13 9 16 13 13 2
19 9 1 9 9 9 13 4 16 4 13 9 1 9 9 7 9 9 9 2
19 9 4 13 9 16 4 13 0 9 15 4 13 9 9 1 9 15 9 2
21 9 13 16 9 9 11 11 13 15 1 9 9 2 7 12 9 13 9 7 9 2
42 2 1 9 1 9 9 15 9 4 13 3 0 9 2 14 13 4 14 0 16 4 15 13 13 2 2 13 4 1 11 0 9 9 1 9 7 9 9 9 11 11 2
26 11 4 13 16 4 9 13 7 13 9 9 2 7 15 3 3 13 1 9 2 3 3 13 13 9 2
32 11 4 3 13 16 0 9 3 4 4 0 1 9 9 9 2 7 16 9 7 3 4 13 4 15 9 1 9 9 0 9 2
20 11 15 13 1 0 12 9 1 9 1 9 9 1 9 2 1 11 7 11 2
13 11 13 1 9 1 9 11 2 7 3 9 1 9
20 1 9 1 9 11 2 1 9 11 2 12 9 4 13 2 7 12 4 0 2
32 12 11 13 4 2 7 3 9 4 0 1 15 4 15 9 11 7 11 13 1 9 11 1 9 11 1 9 2 12 9 2 2
17 9 9 1 9 4 9 13 15 9 2 7 4 4 9 1 9 2
21 0 9 0 9 11 11 13 4 16 4 9 4 0 2 7 16 15 9 13 9 2
16 2 2 13 2 0 9 1 11 2 2 13 4 11 1 11 2
14 2 15 15 4 0 4 16 15 9 13 7 13 2 2
21 11 4 0 9 1 15 4 9 0 1 3 4 11 13 13 15 9 1 9 11 2
13 9 11 11 11 13 4 9 7 13 15 9 11 2
33 2 3 2 16 13 0 9 7 16 13 9 9 1 9 11 2 14 15 15 13 11 1 11 7 1 11 2 2 13 4 1 11 2
24 9 11 11 11 13 4 1 11 16 4 1 9 13 16 4 9 9 13 13 9 1 15 9 2
16 2 3 4 13 1 9 2 12 9 4 0 2 12 4 13 2
13 11 3 4 4 0 2 2 13 4 11 1 11 2
8 13 4 16 4 9 3 0 2
8 2 13 15 16 4 13 3 2
17 9 4 13 13 9 1 16 13 9 2 2 13 4 11 1 11 2
17 0 9 1 11 11 11 13 4 1 11 16 13 9 1 0 9 2
19 11 4 9 13 2 0 9 2 2 15 4 2 13 4 0 14 3 2 2
24 9 15 13 1 9 0 9 1 9 0 9 11 2 3 4 11 9 2 7 0 9 13 9 2
35 3 1 9 2 9 0 11 1 11 13 4 9 16 4 13 12 9 15 4 13 13 1 0 9 3 1 11 12 1 9 0 0 9 11 2
16 11 4 13 16 4 9 9 4 2 0 2 0 7 0 2 2
38 0 9 11 13 4 9 9 11 1 9 2 11 11 2 15 4 13 16 4 11 1 9 13 2 0 2 9 2 16 13 2 9 0 9 1 0 9 2
32 11 4 13 16 4 11 13 9 2 1 9 2 2 7 16 2 9 14 13 9 11 7 0 0 9 2 3 3 9 11 2 2
17 11 11 2 9 0 9 2 13 4 1 11 16 13 9 0 9 2
10 0 9 4 0 1 9 11 1 9 2
6 2 4 4 0 9 2
21 15 4 9 2 11 2 15 15 13 0 7 0 9 2 2 13 4 11 1 11 2
21 9 1 9 11 13 4 9 0 9 11 11 11 2 15 4 13 1 0 9 11 2
13 2 0 2 0 9 13 9 9 7 9 1 9 2
17 0 4 2 2 2 1 9 0 9 3 11 2 2 13 4 11 2
24 13 4 11 7 11 16 13 1 9 7 9 2 7 13 13 9 1 9 2 15 3 4 0 2
13 9 7 9 2 0 0 9 4 4 1 9 0 9
16 0 0 9 11 11 4 4 1 9 0 9 1 0 9 9 2
38 3 1 9 1 9 7 9 2 9 9 0 11 11 13 9 0 9 9 7 9 2 7 0 9 13 16 4 0 9 0 9 13 4 9 9 1 9 2
29 0 0 9 11 11 13 4 9 0 9 7 0 9 9 1 12 7 12 9 2 13 4 12 9 0 9 0 9 2
17 0 9 13 4 0 9 1 9 9 15 4 12 9 0 1 11 2
19 9 9 0 11 11 13 4 12 9 9 1 9 1 0 9 9 7 9 2
14 9 4 0 1 11 2 1 11 2 1 0 9 9 2
31 1 9 0 9 1 9 11 11 0 4 16 0 9 15 13 0 9 13 4 9 9 1 9 2 13 4 12 9 9 11 2
19 1 9 2 0 9 15 13 0 9 3 4 0 7 13 4 9 0 9 2
28 0 9 1 9 1 9 9 1 0 9 11 1 11 13 4 12 9 0 9 3 0 9 8 1 9 0 9 2
21 1 9 2 9 4 13 9 3 9 1 0 9 1 0 9 16 4 13 0 9 2
25 9 0 9 13 4 9 0 9 15 3 1 3 4 4 0 1 11 2 13 4 12 9 0 8 2
20 0 9 2 9 4 13 3 12 9 15 0 9 9 15 4 4 0 1 9 2
37 3 12 9 9 1 11 13 9 9 2 1 9 1 12 9 9 2 13 9 15 4 13 0 9 1 9 7 9 1 9 9 0 9 9 12 9 2
25 9 13 16 4 9 0 9 15 13 9 2 12 9 2 3 0 1 9 11 2 15 13 12 9 2
7 0 0 0 9 0 9 11
16 0 0 9 0 9 11 7 11 13 9 12 0 0 9 11 2
11 9 4 13 0 7 0 0 9 7 9 2
40 1 9 0 9 2 0 9 2 0 9 7 9 1 11 2 9 9 11 7 11 2 11 2 13 4 1 9 2 12 9 2 1 11 0 0 9 0 9 11 2
25 0 9 0 9 11 9 4 9 9 15 13 12 9 2 9 7 0 9 1 12 0 0 9 11 2
14 9 4 13 7 13 9 0 0 7 0 9 7 9 2
23 1 9 0 9 9 11 11 11 2 13 15 16 4 0 9 4 0 12 9 1 0 9 2
13 13 15 16 4 9 9 7 9 13 3 12 9 2
28 1 9 0 9 11 13 15 9 9 0 2 11 2 7 9 9 2 11 2 1 15 12 9 2 0 7 0 2
29 1 0 9 9 2 15 15 13 15 9 2 0 9 0 4 12 0 0 9 1 0 9 9 11 7 0 9 11 2
23 0 9 13 12 9 2 12 9 7 12 9 2 15 4 0 1 15 9 1 11 7 11 2
28 1 9 9 1 0 0 9 1 11 2 9 4 13 0 0 9 15 0 9 2 7 1 9 11 1 0 9 2
39 0 9 1 0 9 13 4 16 4 0 9 11 11 11 2 9 0 9 15 4 13 9 2 13 1 0 9 9 11 2 11 11 2 0 9 1 9 9 2
22 16 15 4 11 13 16 13 9 2 11 4 13 9 9 11 11 11 2 9 0 9 2
19 15 4 0 9 1 9 1 11 16 4 9 11 3 13 0 9 0 9 2
29 2 15 1 3 4 13 0 0 9 1 9 15 4 13 0 9 1 9 7 9 1 15 9 2 2 13 4 11 2
17 2 3 4 13 15 9 7 1 9 1 0 9 1 9 13 9 2
6 9 4 9 0 9 2
19 3 2 12 9 12 4 15 0 9 1 9 9 2 9 9 7 9 2 2
29 9 1 11 13 4 0 12 9 9 1 12 9 2 13 4 1 9 9 2 3 9 1 9 9 7 1 0 9 2
40 15 9 0 4 9 1 9 1 11 2 7 9 1 9 0 9 13 4 13 0 9 9 1 12 9 2 13 4 9 1 15 9 0 1 9 2 12 9 2 2
28 1 12 9 2 9 4 13 0 12 9 9 2 13 4 0 9 0 9 1 9 11 11 2 13 15 1 9 2
37 2 13 16 4 1 0 9 0 9 13 3 12 9 9 2 7 15 3 13 1 15 9 16 13 0 9 1 9 9 1 0 9 2 2 13 4 2
27 0 9 2 1 0 9 2 9 4 9 1 9 0 9 2 16 4 15 13 9 0 0 9 7 15 9 2
30 1 0 9 9 13 4 2 1 0 9 2 4 0 0 9 2 13 4 11 2 15 4 3 9 0 9 1 0 9 2
41 0 9 15 4 13 13 9 9 0 4 9 1 9 2 15 15 3 13 9 0 9 15 15 13 13 1 9 7 3 13 0 9 0 1 15 9 2 13 4 11 2
43 2 1 9 0 9 13 4 0 16 4 1 9 9 1 0 0 9 13 1 12 1 12 9 2 16 4 3 15 4 0 1 9 1 12 1 12 9 2 2 13 4 9 2
19 1 0 9 2 9 4 13 9 9 7 13 15 3 1 9 1 9 9 2
23 2 0 9 2 3 1 9 4 4 1 9 13 9 2 15 4 13 1 0 9 9 2 2
43 11 2 15 4 9 1 9 0 9 0 1 9 0 9 3 15 9 2 13 16 4 9 0 9 1 9 9 2 7 9 15 9 9 2 13 9 0 9 1 0 12 9 2
23 1 9 9 9 1 9 11 11 2 9 11 1 9 12 9 15 9 13 4 12 9 9 2
9 0 9 13 4 3 12 9 9 2
29 1 0 9 0 9 15 9 2 12 4 0 3 9 2 12 1 9 2 7 12 9 0 9 0 4 1 9 9 2
29 2 1 12 9 13 9 12 9 1 9 2 9 12 9 7 9 12 9 9 1 9 0 9 2 2 13 4 11 2
25 1 0 9 0 1 9 1 9 13 15 9 9 1 9 11 2 0 9 7 3 0 7 0 9 2
8 15 1 0 9 13 9 1 11
19 12 15 0 9 15 9 13 11 7 13 0 9 9 1 11 16 0 9 2
16 9 7 0 0 9 9 11 11 13 1 9 15 9 1 9 2
15 9 1 11 7 11 12 4 0 9 9 0 0 9 1 12
26 9 1 15 12 0 9 13 9 9 0 9 7 0 9 2 7 9 15 13 0 7 0 9 9 9 2
16 3 4 13 16 15 9 11 13 9 1 0 7 0 9 9 2
19 9 13 9 0 9 15 13 16 4 9 13 0 9 0 9 7 0 9 2
22 0 9 15 3 13 13 0 0 9 2 15 4 0 1 9 0 9 7 9 9 9 2
19 1 0 9 2 0 9 13 0 9 9 7 13 1 9 0 7 0 9 2
17 3 2 3 4 13 15 1 15 9 9 1 11 13 1 0 9 2
11 9 3 4 15 15 4 4 1 0 9 2
11 0 0 9 2 0 9 2 3 14 13 2
18 9 4 15 16 4 9 0 0 9 13 0 2 16 7 9 0 9 2
9 3 4 3 13 1 9 9 9 2
19 1 9 15 3 13 1 0 9 9 2 13 15 16 4 0 9 0 9 2
14 9 13 0 9 9 2 1 15 1 11 13 0 9 2
29 9 14 13 13 9 1 9 0 0 2 0 7 0 9 0 9 2 16 15 15 9 13 2 13 15 7 9 9 2
18 1 0 9 2 9 1 11 3 4 12 1 9 15 13 13 0 9 2
19 1 9 4 9 9 15 4 9 9 2 16 13 4 0 9 1 0 9 2
32 1 0 9 2 0 9 1 11 2 0 9 2 13 13 15 0 0 2 0 7 0 9 16 14 4 13 1 9 9 15 9 2
29 15 13 1 9 1 9 0 9 9 2 16 4 15 13 1 0 9 2 7 11 3 3 13 0 8 8 8 9 2
31 3 4 16 12 1 9 13 1 9 2 0 9 2 15 4 13 1 9 0 9 2 7 1 14 0 9 13 1 0 9 2
16 3 2 15 4 9 3 0 1 9 0 0 9 7 0 9 2
20 1 15 9 2 15 9 13 9 1 9 0 9 2 15 4 3 0 1 11 2
28 9 15 4 9 9 11 2 11 2 15 4 13 9 9 0 9 1 15 4 11 13 11 9 1 9 0 9 2
29 11 2 11 7 11 13 13 1 9 1 11 1 9 1 9 1 11 2 1 15 0 13 0 9 0 9 7 9 2
15 9 1 9 11 13 9 9 1 15 9 7 13 0 9 2
8 0 9 12 13 15 9 9 2
24 1 0 11 9 1 11 13 0 9 9 2 7 13 1 9 0 0 9 7 9 1 0 9 2
17 3 2 11 7 1 15 9 13 14 0 9 0 9 7 0 9 2
10 9 4 7 0 9 0 9 15 9 2
13 9 1 11 3 13 0 9 1 0 9 0 11 2
15 3 2 1 14 0 0 9 2 9 9 14 13 0 9 2
20 3 2 7 9 1 11 2 7 1 11 2 14 13 13 0 7 0 0 9 2
18 9 4 16 0 0 9 7 9 9 9 1 0 9 13 1 0 9 2
10 0 9 1 9 13 13 1 15 0 2
5 9 9 11 7 11
25 9 11 1 9 11 3 4 15 13 1 0 3 9 16 4 1 11 0 9 1 9 1 0 9 2
42 11 9 11 11 7 15 0 9 11 11 13 4 9 1 9 2 12 9 2 1 15 16 13 3 1 0 0 9 1 12 9 2 15 4 0 9 9 11 1 9 11 2
30 1 3 9 9 3 4 9 0 2 11 7 11 13 4 0 9 1 0 9 1 9 0 9 7 13 15 3 13 9 2
33 2 0 9 13 4 0 9 1 0 9 7 9 11 16 11 13 9 9 11 1 9 11 2 2 13 4 9 9 1 9 1 9 2
14 11 4 3 13 0 9 11 2 0 0 0 9 11 2
51 2 7 12 9 7 0 9 1 12 9 12 9 2 3 4 12 9 13 9 1 0 11 2 13 4 15 0 9 1 9 0 9 2 16 1 0 9 3 7 1 9 1 9 11 2 2 13 15 1 9 2
21 2 15 4 9 1 15 0 13 2 2 13 4 11 2 3 16 4 3 0 9 2
17 2 15 13 9 7 9 9 1 0 9 12 9 7 15 9 2 2
28 11 15 13 16 4 9 9 11 13 0 9 7 4 11 13 9 1 9 7 13 9 1 9 9 7 9 9 2
18 11 4 13 16 4 12 9 0 13 9 9 0 9 7 1 9 11 2
20 15 9 13 4 0 9 9 11 2 9 11 1 9 11 11 7 0 0 9 2
24 11 4 13 16 4 0 13 1 0 9 9 2 15 13 9 1 0 9 9 1 9 12 9 2
35 2 9 11 7 11 13 4 0 9 9 0 9 2 2 13 4 0 9 11 11 2 3 16 15 9 2 13 9 9 0 9 7 9 9 2
15 15 4 13 0 9 7 13 16 9 1 0 0 11 2 2
10 11 2 9 4 15 13 9 1 0 9
27 9 11 1 11 13 16 4 15 9 0 1 0 9 13 9 1 9 9 9 7 16 15 14 13 9 11 2
31 0 9 11 13 4 1 9 2 12 9 2 9 1 0 9 0 9 2 15 4 0 9 9 1 9 1 0 9 7 9 2
13 9 4 13 0 11 15 13 16 4 0 9 11 2
14 3 2 11 13 16 1 9 14 13 4 15 0 9 2
18 2 9 1 0 9 1 11 0 4 9 2 2 13 15 1 9 9 2
11 2 9 15 4 9 1 0 9 7 9 2
11 15 4 4 0 1 0 9 1 11 2 2
27 16 4 15 9 13 2 13 15 13 7 13 9 3 9 7 13 15 13 9 1 9 15 2 13 4 11 2
19 2 0 9 4 4 1 0 9 0 1 9 9 2 2 13 15 1 9 2
24 9 13 0 9 12 9 9 11 7 13 15 0 9 1 9 9 9 9 1 11 2 13 9 2
24 9 0 11 7 3 4 0 1 15 16 13 16 15 13 1 9 11 1 9 15 0 0 9 2
8 9 1 11 4 13 15 9 2
20 9 11 11 7 9 11 11 13 4 1 9 0 9 3 16 11 4 9 9 2
18 9 4 13 4 15 9 1 9 2 9 7 0 9 11 2 13 4 2
7 9 9 4 4 3 0 2
18 9 0 9 13 4 1 9 9 1 9 3 16 4 13 9 12 9 2
9 2 3 4 13 14 9 9 11 2
16 15 4 14 11 2 7 14 11 2 2 13 4 1 0 9 2
36 0 9 11 11 13 4 1 9 9 2 9 7 9 11 16 15 13 1 9 9 9 2 1 16 15 13 1 9 16 15 4 9 1 0 9 2
9 9 4 3 3 0 2 13 4 2
11 2 11 4 0 9 2 2 13 4 11 2
16 2 14 14 13 3 13 15 16 4 11 9 7 13 3 2 2
8 11 13 0 9 8 9 1 11
23 11 2 11 2 9 11 13 4 1 9 2 12 9 2 0 7 0 9 8 9 1 11 2
20 1 9 11 11 2 9 9 1 9 2 9 4 13 16 4 11 13 15 9 2
25 11 4 1 3 1 11 13 12 9 9 1 9 9 0 9 1 9 1 12 9 9 0 12 9 2
10 11 7 11 13 1 9 9 1 0 9
14 9 12 9 0 4 1 3 4 11 0 9 13 11 2
34 16 4 9 11 7 11 1 0 9 2 9 9 12 9 13 4 1 9 1 11 1 9 2 12 9 2 2 9 13 9 7 0 9 2
25 0 9 9 11 11 13 15 1 3 0 9 2 3 9 11 11 2 9 11 11 7 9 11 11 2
20 11 7 11 13 4 0 9 1 0 9 7 13 16 4 0 9 9 12 9 2
26 2 13 1 9 0 9 2 0 9 7 9 2 16 7 0 9 7 9 0 9 2 2 13 4 11 2
16 2 0 9 1 9 13 0 9 2 9 1 9 0 9 2 2
20 1 9 11 2 13 3 3 15 1 13 2 3 9 0 9 7 9 0 9 2
36 13 4 16 13 3 9 1 9 1 0 0 9 7 9 9 2 15 4 1 0 9 2 7 13 16 4 0 9 1 11 4 0 1 0 9 2
14 9 12 9 0 4 1 3 4 11 0 9 13 11 2
8 11 4 1 15 13 0 9 2
18 3 2 1 0 9 9 2 9 11 11 11 4 0 1 0 9 11 2
28 11 4 3 13 9 1 0 9 2 7 15 4 13 2 16 4 1 9 0 9 1 0 9 0 1 0 9 2
23 0 0 9 13 4 0 9 11 11 2 15 4 13 16 11 7 11 13 3 13 0 9 2
18 1 9 1 9 2 11 4 13 16 15 11 13 1 0 9 0 9 2
16 2 13 4 13 16 15 11 7 11 14 13 1 9 0 9 2
32 3 2 13 15 16 15 9 13 4 3 1 9 9 7 1 0 4 9 16 15 15 9 3 13 2 16 15 15 13 11 2 2
7 9 9 11 0 1 9 9
32 11 2 11 2 9 4 1 9 2 12 9 2 13 11 11 2 0 9 0 0 0 9 11 2 1 9 9 16 4 13 9 2
9 0 4 15 9 7 9 1 11 2
20 0 9 13 4 16 4 15 9 0 1 9 3 4 4 9 11 2 9 11 2
5 9 3 2 13 2
15 0 0 9 13 1 9 1 15 4 0 12 9 1 11 2
21 9 9 0 0 9 11 11 11 9 4 13 0 1 9 11 11 1 0 9 11 2
16 3 2 1 0 9 15 15 13 2 16 4 9 13 9 11 2
12 9 13 13 9 7 13 15 1 9 1 9 2
7 15 4 4 0 9 9 2
24 0 12 9 1 11 1 11 16 4 4 9 0 9 2 12 9 0 9 13 4 11 12 9 2
10 9 4 15 13 12 9 1 9 11 2
16 0 4 1 9 12 9 7 0 12 2 1 3 15 4 13 2
19 11 4 13 9 1 15 9 12 9 2 3 3 12 9 9 1 0 9 2
45 9 4 3 13 16 9 1 9 0 9 7 0 9 2 3 0 9 11 11 2 0 9 11 11 2 0 0 9 11 11 2 0 0 9 11 11 7 0 9 11 11 7 11 11 2
8 11 4 13 9 1 12 9 2
15 2 9 4 0 1 9 15 15 4 15 13 1 0 9 2
16 9 4 15 13 1 9 9 2 2 13 4 9 11 11 11 2
13 13 15 16 4 9 9 13 3 1 12 9 9 2
7 3 2 9 4 13 3 2
30 9 4 0 7 0 1 9 3 16 9 2 0 9 11 11 11 2 4 13 0 9 9 11 2 3 4 13 13 9 2
21 9 11 13 4 9 12 9 16 4 13 9 9 2 7 9 4 3 3 1 9 2
13 9 4 13 13 0 1 0 9 7 13 0 9 2
18 9 4 15 13 13 1 9 2 13 9 7 13 1 9 15 0 9 2
5 13 14 11 0 2
21 9 11 11 11 13 16 11 13 13 0 9 1 9 11 2 7 9 13 1 15 2
12 0 9 1 11 13 9 1 3 0 0 9 2
15 1 3 9 9 4 13 13 9 1 11 1 9 12 9 2
32 9 11 11 11 3 15 13 9 11 15 4 15 13 9 7 13 0 2 16 7 13 9 1 0 9 7 13 0 9 1 9 2
20 2 16 15 13 9 11 15 4 1 9 1 9 11 2 13 4 15 2 2 2
10 15 13 16 15 9 9 4 0 9 2
11 15 4 0 2 2 13 4 11 9 11 2
30 16 9 13 16 4 0 9 13 13 0 9 2 11 13 1 15 9 2 3 16 4 11 1 9 13 15 9 0 9 2
41 3 9 0 0 9 2 9 11 2 9 1 9 1 11 2 13 4 9 1 12 1 12 9 2 1 0 9 9 1 12 9 2 3 15 1 3 12 9 0 9 2
26 1 15 9 2 11 2 15 13 3 1 12 9 9 2 12 9 4 4 0 1 12 0 9 1 9 2
10 3 2 9 0 0 9 13 4 11 2
28 9 4 0 1 0 12 9 1 9 2 16 4 9 1 9 4 3 12 9 0 1 9 1 0 9 0 9 2
20 9 13 16 4 0 9 13 13 1 9 2 3 9 1 12 9 1 12 9 2
14 15 9 13 16 4 11 1 11 9 1 9 0 9 2
24 16 11 7 11 13 13 9 2 13 15 16 4 11 13 1 0 9 1 12 7 12 9 9 2
21 3 2 9 4 13 7 9 15 9 2 15 4 13 4 0 1 0 9 7 9 2
12 9 1 2 0 9 2 11 13 4 0 9 2
22 0 9 0 9 7 9 2 11 2 2 16 7 0 9 2 13 1 0 9 1 11 2
12 9 2 1 0 9 2 13 1 9 15 9 2
34 2 15 4 0 9 1 11 2 7 15 4 0 9 7 14 13 15 13 3 2 2 13 4 11 11 2 0 11 9 9 2 11 2 2
34 1 9 11 2 11 4 0 9 13 9 0 9 2 1 9 9 12 0 0 9 2 9 9 1 0 9 9 7 9 0 0 9 9 2
14 4 3 13 14 15 9 0 1 15 13 0 0 9 2
29 9 9 0 9 11 11 11 13 4 0 9 2 7 4 13 16 13 9 1 9 2 16 14 4 0 9 1 11 2
15 2 1 0 9 0 9 2 13 15 0 9 1 0 9 2
23 3 15 13 0 9 1 11 2 15 4 15 0 9 13 1 0 9 2 2 13 4 11 2
24 2 1 12 9 0 9 1 9 7 11 2 3 4 0 15 9 3 13 15 4 3 3 2 2
5 11 7 11 13 11
35 0 9 1 0 9 2 11 2 1 11 7 11 2 15 13 1 9 1 9 2 13 4 2 16 15 13 2 3 12 9 9 1 0 9 2
11 9 15 1 9 13 1 9 0 9 9 2
27 1 12 9 12 9 11 7 11 2 11 2 4 13 9 1 0 9 2 11 2 1 0 9 1 12 9 2
17 16 9 15 11 14 4 4 0 9 1 11 15 13 15 9 9 2
20 13 15 16 4 9 9 13 0 9 0 12 9 9 2 16 7 13 0 9 2
23 1 9 9 13 1 0 0 9 1 15 4 0 9 7 0 9 13 9 1 0 0 9 2
26 15 4 13 16 4 0 0 0 9 2 16 15 4 9 2 9 2 9 7 9 2 13 4 0 9 2
25 9 9 9 0 2 11 2 13 4 9 1 9 12 9 11 2 1 9 1 9 1 0 0 9 2
17 11 7 9 0 9 0 4 3 16 4 0 0 9 13 9 11 2
22 11 15 13 1 9 9 2 1 15 0 0 9 13 16 4 13 9 9 1 12 9 2
30 0 9 15 9 3 4 13 0 7 15 1 0 9 2 7 0 9 11 11 13 9 1 9 9 16 4 13 15 9 2
36 2 11 4 13 9 1 0 3 9 16 7 1 0 9 9 7 1 15 4 1 9 4 3 13 15 9 16 4 13 0 2 2 13 4 11 2
30 9 1 12 9 11 13 4 16 4 1 9 9 9 11 4 0 3 12 9 9 2 7 9 9 13 16 15 4 3 2
34 2 16 3 13 13 9 16 13 11 4 4 3 16 9 7 9 13 15 0 9 7 0 9 2 2 13 4 9 9 9 11 11 11 2
32 9 9 11 13 4 16 15 9 7 9 13 0 9 2 1 9 9 16 4 4 1 9 13 1 9 1 0 9 3 0 9 2
23 3 2 0 9 13 4 0 9 1 15 9 2 3 16 15 14 4 13 13 1 9 11 2
