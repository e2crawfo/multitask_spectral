557 11
59 9 1 12 9 12 13 1 11 11 1 9 11 12 7 12 9 0 13 1 0 15 13 1 13 9 1 9 11 2 11 0 9 13 11 3 13 0 1 9 9 9 2 13 1 9 0 1 11 11 7 13 1 9 12 11 1 9 0 2
11 11 13 9 15 13 1 11 11 2 11 2
13 0 9 9 11 11 11 15 3 13 1 9 10 2
11 9 7 9 3 3 3 13 1 9 10 2
20 1 12 9 1 9 11 11 12 13 2 15 3 13 13 9 1 9 9 11 2
13 11 11 13 9 1 10 9 9 7 9 9 9 2
17 15 3 13 3 10 9 10 3 9 7 10 9 10 3 3 9 2
29 11 3 13 1 13 9 2 7 10 9 9 1 9 2 9 2 9 2 9 2 9 2 7 9 3 3 13 0 2
11 16 15 13 3 13 7 13 9 1 11 2
21 3 0 2 11 13 9 1 11 2 15 3 13 9 2 11 13 9 0 11 2 2
37 1 11 2 11 11 9 3 13 9 15 14 3 13 2 16 9 9 9 15 3 13 1 0 7 1 9 9 13 0 16 11 11 14 3 13 9 2
24 1 0 9 12 2 13 11 11 12 2 12 1 9 9 9 0 15 13 1 11 2 11 11 2
14 11 13 10 9 2 9 2 7 3 9 9 0 11 2
9 11 13 3 11 11 13 13 9 2
68 3 11 11 11 13 9 11 11 3 11 9 11 13 11 11 15 13 1 1 11 11 9 10 14 13 0 16 9 11 11 12 2 3 1 9 9 3 1 3 13 10 9 9 7 9 9 1 11 1 9 16 11 3 13 10 9 11 1 13 13 3 13 10 9 0 11 11 2
25 3 13 13 1 9 11 2 9 2 2 11 2 9 2 2 11 2 9 2 2 11 2 9 2 2
11 7 10 2 10 9 13 10 9 9 9 2
40 11 11 11 2 11 2 13 9 9 9 0 15 13 10 9 5 9 9 2 9 9 9 9 9 5 9 5 9 2 9 0 2 7 9 2 9 1 10 11 2
8 15 3 9 15 0 10 11 2
19 9 10 3 3 13 1 11 11 2 7 10 9 0 1 11 11 7 11 2
9 9 0 1 9 10 13 11 11 2
18 13 1 12 9 9 0 15 13 1 9 9 7 9 9 1 9 11 2
14 16 15 13 15 15 13 2 16 10 9 0 2 0 2
36 11 10 13 1 11 15 3 13 9 0 2 11 11 1 9 13 1 9 9 15 13 12 5 2 11 11 9 13 9 9 15 13 13 12 5 2
6 11 10 13 9 12 2
46 1 11 11 11 11 11 11 11 11 9 11 3 11 11 11 9 2 13 2 2 16 9 11 11 12 9 9 9 9 3 13 1 10 9 9 2 10 9 0 15 13 7 13 9 2 2
67 9 2 9 9 15 3 0 1 9 9 7 11 11 1 11 11 13 1 9 2 9 0 0 1 11 11 2 1 9 9 11 2 2 9 11 2 9 9 11 11 2 2 11 2 11 7 11 2 16 13 1 9 11 16 1 9 11 2 3 13 9 2 5 1 11 2 2
17 1 12 15 13 1 15 3 13 2 1 9 9 1 13 2 2 2
11 11 11 3 13 11 11 15 13 11 11 2
30 15 13 9 1 11 11 2 7 13 1 9 0 1 9 12 2 12 2 7 9 9 1 9 13 9 1 9 9 0 2
14 15 13 9 1 9 2 15 13 1 9 0 13 11 2
35 9 1 9 2 11 11 2 7 9 1 9 11 2 9 10 3 13 1 9 12 2 7 1 12 2 9 10 13 1 9 9 1 9 9 2
15 9 1 9 11 9 11 12 3 13 1 9 9 9 10 2
11 11 11 11 11 11 13 9 1 12 12 2
18 11 11 13 10 10 9 1 11 11 2 11 11 2 11 11 2 11 2
15 2 16 1 3 9 15 13 1 9 2 9 9 9 10 2
10 1 0 3 3 13 7 9 2 9 2
15 16 9 10 13 1 9 11 16 11 13 7 13 1 9 2
63 9 10 13 9 12 2 12 1 9 11 2 9 10 13 1 12 9 15 13 11 11 11 2 11 11 11 11 2 11 11 9 11 2 7 11 11 11 11 2 2 15 13 12 9 9 2 1 11 11 11 2 11 11 2 7 11 11 11 13 12 9 0 2
29 11 13 1 11 11 1 11 11 2 11 11 11 2 11 2 11 2 1 12 1 10 9 2 3 9 13 9 9 2
32 1 13 2 9 13 1 9 13 9 9 0 2 9 9 9 2 7 9 15 13 13 9 2 9 0 2 7 9 9 1 9 2
19 16 13 9 11 2 16 9 9 1 11 11 11 11 2 11 2 3 0 2
14 11 13 1 11 11 1 12 7 13 9 1 9 9 2
19 11 11 2 2 11 11 2 2 13 9 15 13 1 11 1 11 2 11 2
19 11 13 10 9 9 1 9 11 11 2 9 11 2 11 11 11 2 11 2
7 16 3 15 13 9 3 2
21 15 13 9 7 9 2 9 1 13 7 13 9 11 1 10 9 9 9 7 9 2
24 11 13 10 9 13 12 9 15 13 1 9 11 2 11 11 2 9 11 2 1 1 9 11 2
21 16 14 9 15 3 13 11 13 2 7 13 2 9 9 2 15 3 15 3 13 2
21 12 2 9 13 11 1 11 2 10 9 0 13 16 9 10 2 13 1 9 2 2
20 16 16 9 2 9 13 13 9 9 2 11 13 3 1 11 9 12 2 12 2
23 9 9 7 9 11 1 9 12 1 11 7 1 9 0 3 3 15 13 16 9 9 9 2
19 9 13 2 9 2 1 9 7 9 2 9 15 13 1 9 13 9 9 2
8 0 9 11 2 11 7 11 2
10 1 9 10 2 11 13 13 11 11 2
25 15 13 0 3 13 2 0 15 10 9 15 3 15 13 1 15 15 3 13 9 9 10 9 0 2
13 9 10 3 13 1 10 10 9 1 9 1 11 2
32 11 3 3 13 1 9 9 9 11 2 16 15 13 10 9 1 13 1 3 0 7 3 0 1 9 9 9 7 9 9 9 2
29 12 9 0 13 12 2 12 2 12 2 12 2 12 2 12 2 7 12 2 12 13 1 9 12 9 1 9 12 2
16 11 13 9 9 1 10 9 11 16 9 13 1 13 9 9 2
13 9 10 13 9 2 9 15 13 1 9 9 11 2
12 11 11 13 9 1 10 9 0 15 13 9 2
24 15 13 9 1 11 11 1 9 13 9 1 11 2 5 11 11 13 10 9 9 0 1 11 2
20 11 13 9 0 13 1 9 2 9 2 9 9 2 9 7 9 2 9 0 2
12 9 10 13 2 13 2 7 13 1 11 11 2
10 3 9 13 9 11 10 2 16 13 2
26 11 11 7 9 9 2 9 13 9 9 15 13 1 12 9 9 9 1 10 10 9 9 9 2 9 2
11 11 11 13 1 9 1 2 12 7 12 2
19 9 9 12 9 13 1 10 9 11 13 11 11 1 0 9 10 2 12 2
25 0 2 0 10 2 9 3 13 9 2 9 2 11 11 2 7 10 9 15 13 11 11 1 9 2
27 1 9 15 13 1 11 11 11 2 9 15 3 0 13 1 9 2 10 9 7 15 0 1 9 9 0 2
18 15 13 15 11 2 11 15 0 15 13 9 9 12 9 12 2 12 2
12 11 13 10 9 1 11 11 2 11 2 11 2
20 14 9 3 3 3 13 9 1 9 10 9 0 3 13 1 9 9 0 11 2
13 1 11 11 2 11 3 13 9 0 1 9 10 2
14 1 9 13 9 11 11 9 2 9 15 0 7 0 2
10 11 13 9 9 2 9 0 7 13 2
19 11 3 13 9 2 15 3 13 11 13 7 13 1 11 2 11 11 11 2
12 11 10 13 12 9 7 12 9 15 3 0 2
23 11 11 11 2 11 11 13 11 1 12 1 13 9 11 11 1 11 11 11 1 11 11 2
13 15 13 9 9 1 9 9 11 11 11 11 11 2
25 3 10 9 10 13 2 1 10 9 11 2 15 13 1 9 1 9 9 13 9 9 1 9 12 2
9 9 9 9 15 3 13 9 10 2
14 16 11 11 13 9 9 12 2 11 11 13 15 0 2
18 11 2 9 2 9 7 9 0 13 1 11 1 13 9 1 9 11 2
52 16 1 2 11 11 11 11 11 12 9 10 13 1 11 12 11 2 1 9 11 11 11 11 12 15 13 9 9 11 2 12 11 12 2 11 3 13 1 11 11 11 11 12 7 11 13 11 11 11 11 12 2
49 11 12 9 3 13 1 9 11 11 15 13 9 3 0 1 11 12 7 11 12 2 11 13 9 9 9 15 13 1 11 13 9 9 13 9 1 9 12 15 13 0 2 7 1 9 15 14 0 2
22 9 9 9 13 12 9 2 7 13 12 9 0 2 15 9 3 13 1 9 9 9 2
12 3 11 11 7 11 11 13 13 9 15 13 2
15 3 11 13 9 1 9 2 16 15 3 0 13 3 0 2
23 1 9 10 2 15 13 9 9 15 13 13 11 13 9 0 7 13 9 10 13 9 11 2
26 1 9 10 12 9 9 10 13 3 0 1 9 12 7 12 1 9 9 2 1 9 1 9 0 0 2
52 1 1 9 9 12 2 12 2 11 11 13 16 11 11 13 1 1 9 1 1 9 13 1 11 2 16 13 9 15 3 0 1 9 11 7 3 9 9 0 13 1 1 9 11 7 13 1 1 9 11 11 2
19 11 11 13 9 1 12 9 2 11 1 9 12 2 13 9 1 12 9 2
25 16 11 3 13 0 2 11 0 13 11 11 2 11 11 2 2 9 9 11 15 13 13 9 11 2
9 11 11 13 1 11 1 9 12 2
20 1 9 9 2 9 13 9 0 12 2 12 9 1 9 0 7 0 15 0 2
31 3 14 13 2 9 12 2 1 12 9 2 3 12 9 1 1 3 13 2 1 0 12 9 13 9 7 12 9 13 9 2
24 11 11 11 13 1 1 9 11 11 7 9 3 13 1 9 11 2 11 2 15 13 9 11 2
18 11 13 9 1 9 0 0 0 15 13 9 11 1 9 11 11 11 2
14 11 11 13 10 9 1 11 11 2 11 11 2 11 2
70 9 10 3 13 1 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 11 11 2 7 9 9 11 13 1 9 9 1 9 9 11 1 1 11 11 9 9 2
34 11 2 11 11 11 2 15 13 13 11 11 7 11 11 11 2 9 3 13 10 9 10 7 3 13 1 9 2 15 0 3 13 9 2
14 9 9 15 11 2 12 9 7 12 9 2 14 0 2
24 13 10 9 1 13 9 2 9 15 13 2 10 2 10 3 13 16 14 3 13 12 7 0 2
7 9 10 3 9 1 9 2
19 11 11 13 10 10 9 1 9 11 11 2 11 11 2 11 11 2 11 2
26 7 3 2 1 9 2 9 10 9 9 9 3 13 1 9 9 2 9 1 9 9 11 7 9 9 2
28 15 13 9 9 9 11 11 11 2 13 0 16 14 0 1 9 9 11 9 2 11 11 2 15 13 1 9 2
25 11 11 9 2 13 9 9 11 11 2 13 9 9 9 0 1 11 15 13 1 11 11 11 11 2
14 3 13 9 2 12 9 10 13 2 1 13 9 15 2
26 11 9 3 13 3 9 13 9 2 9 2 7 9 15 1 9 9 1 9 0 15 13 9 1 0 2
51 9 9 13 1 9 11 13 9 9 2 15 13 11 11 1 11 2 11 11 13 9 11 9 11 5 9 2 11 7 9 10 3 13 1 9 2 3 13 1 9 9 9 2 9 2 9 7 9 2 9 2
5 3 9 15 13 2
17 9 0 2 11 13 7 13 11 3 13 1 9 1 11 7 11 2
16 9 3 13 1 12 9 1 11 2 12 1 11 7 12 11 2
8 11 13 11 16 9 14 13 2
23 11 11 13 9 0 1 9 15 3 13 9 2 9 1 9 9 1 9 7 0 2 9 2
12 9 9 3 3 13 1 11 11 1 13 9 2
20 11 13 10 9 1 9 2 9 7 1 3 0 9 13 1 9 2 9 13 2
17 16 3 13 11 11 2 9 3 13 9 9 11 11 1 9 12 2
11 15 13 1 11 11 2 11 2 15 0 2
10 3 13 1 9 0 1 9 11 12 2
33 1 10 9 1 11 11 1 9 12 11 12 2 11 13 1 2 2 3 15 13 2 9 10 15 13 1 9 2 9 9 9 2 2
24 9 10 3 13 1 13 9 15 13 1 9 0 7 13 1 13 3 9 15 13 1 9 15 2
8 12 9 9 13 1 11 12 2
29 2 11 2 3 9 2 9 13 9 9 7 9 0 1 9 2 9 2 7 9 1 9 15 13 1 9 15 0 2
18 1 9 1 9 0 2 15 13 13 9 9 2 9 1 13 9 9 2
105 1 9 9 2 11 11 11 11 13 9 9 1 10 9 2 9 9 2 12 9 9 9 2 1 9 7 1 9 2 2 9 2 9 9 2 9 15 13 1 9 0 1 11 5 11 1 11 11 2 9 2 9 9 2 9 2 9 7 9 1 10 9 2 9 2 9 1 11 11 11 11 11 2 3 2 11 2 11 2 11 2 2 11 2 11 11 2 11 2 11 2 11 2 7 11 2 7 9 9 9 2 9 2 9 2
26 3 9 13 1 11 1 9 12 2 16 9 2 15 13 11 11 2 9 9 11 7 11 11 11 2 2
4 3 9 0 2
27 13 7 9 15 13 9 9 2 9 11 2 16 13 1 9 15 0 2 3 13 1 9 9 2 9 0 2
23 9 9 9 9 13 0 9 9 9 1 9 9 9 2 9 2 9 2 9 2 7 9 2
5 15 13 1 9 2
14 9 10 13 1 9 9 11 11 11 2 0 11 11 2
13 11 11 7 11 3 13 9 1 9 0 9 10 2
13 16 13 9 2 11 13 9 9 7 3 13 0 2
32 16 1 13 1 10 9 2 3 13 9 1 13 9 15 13 11 11 2 11 11 2 1 12 9 12 9 2 12 11 12 2 2
19 11 3 13 9 9 15 13 11 11 7 11 11 2 9 15 13 9 11 2
11 3 13 9 15 13 9 1 11 1 11 2
19 12 9 0 13 1 0 2 16 9 12 2 12 13 1 9 11 2 11 2
5 15 13 1 9 2
11 16 13 12 2 11 11 11 13 11 11 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
33 11 9 13 1 9 2 12 9 1 9 9 15 13 9 1 13 13 2 7 9 13 1 9 11 2 7 3 13 1 10 9 2 2
33 9 0 11 2 11 11 11 2 2 11 11 11 2 2 2 15 13 1 9 12 2 13 10 10 9 1 9 9 0 1 9 0 2
57 9 1 9 13 1 9 9 9 2 9 9 13 1 10 9 2 11 2 13 9 9 9 9 0 3 13 9 11 15 13 1 9 2 1 2 11 9 2 13 9 11 9 1 0 7 1 9 9 9 15 13 1 13 9 0 0 2
23 16 9 9 13 14 13 13 9 2 16 11 13 13 9 10 9 2 13 9 1 13 9 2
12 16 2 11 13 9 11 11 0 3 1 9 2
11 9 9 13 9 1 9 9 1 9 0 2
15 11 11 13 9 1 11 11 2 11 2 11 11 2 11 2
26 1 1 11 11 2 13 11 11 15 13 9 11 11 7 3 13 11 11 13 12 9 2 9 7 9 2
3 13 15 2
11 15 3 13 1 9 0 1 9 9 11 2
21 13 1 11 11 11 11 11 1 9 12 2 9 10 3 0 1 3 1 12 9 2
5 3 9 1 11 2
20 9 9 11 1 11 7 11 1 9 12 13 9 15 13 1 9 15 11 12 2
34 11 13 1 1 12 9 15 13 1 11 11 11 2 11 12 7 3 3 13 11 11 15 13 1 10 9 15 13 1 9 11 11 11 2
19 3 1 12 9 13 1 12 9 9 15 13 0 1 9 7 0 1 9 2
22 9 9 11 13 11 11 11 11 15 13 11 2 11 2 2 11 2 11 2 7 11 2
26 9 10 13 1 9 9 15 3 0 13 9 9 1 13 9 2 9 0 1 10 10 9 0 2 11 2
13 3 9 1 9 3 13 1 1 10 9 1 11 2
11 11 3 13 10 9 9 1 9 9 9 2
14 1 9 12 2 9 13 9 9 15 0 0 1 9 2
12 11 13 7 11 13 9 0 2 14 3 13 2
14 16 9 10 0 2 7 0 2 3 9 9 1 9 2
24 11 11 11 11 13 9 9 9 11 2 11 1 9 11 11 2 13 12 5 1 1 9 11 2
11 11 11 3 13 13 9 1 11 11 11 2
12 10 9 1 11 13 2 9 0 2 9 10 2
18 11 11 2 13 9 0 0 1 9 2 9 2 15 13 1 9 12 2
24 1 11 3 13 12 9 9 9 15 13 2 16 9 9 2 9 15 14 13 7 9 9 9 2
23 1 11 2 15 13 16 11 11 13 13 1 11 11 11 2 16 11 11 7 11 13 9 2
16 11 11 13 9 11 11 15 12 2 12 1 10 9 11 11 2
20 1 9 9 2 11 11 13 1 11 2 11 3 13 10 9 1 9 9 12 2
16 11 11 2 2 13 10 9 9 9 9 15 13 1 9 9 2
16 13 1 11 13 2 2 15 13 11 13 10 9 9 2 14 2
21 11 2 11 2 11 11 11 11 2 2 13 1 12 11 12 1 0 1 11 11 2
10 15 13 11 11 13 11 11 11 11 2
19 15 13 9 0 1 9 1 9 12 11 2 1 9 12 2 12 1 11 2
23 1 9 12 2 11 11 11 13 9 11 3 2 3 13 15 15 13 13 1 9 0 2 2
24 11 11 3 13 1 11 11 2 13 10 9 13 11 2 7 3 13 1 12 9 1 11 11 2
41 1 9 2 9 11 2 7 9 2 9 0 2 12 9 13 11 1 3 2 3 1 9 1 9 1 13 9 11 1 9 9 11 2 9 11 2 7 10 9 0 2
21 11 11 13 9 15 3 13 1 9 0 15 13 1 9 11 15 0 1 9 9 2
18 9 9 10 13 11 2 15 13 11 7 9 13 9 0 1 9 10 2
24 11 11 13 10 10 9 15 13 1 11 11 11 2 9 11 11 11 2 11 11 11 2 11 2
9 11 11 13 9 11 1 12 9 2
34 15 3 13 9 9 11 11 1 9 13 11 2 9 7 11 2 11 11 2 11 11 2 11 5 11 1 11 11 7 11 11 11 11 2
14 11 13 9 10 7 1 0 13 9 9 9 1 9 2
12 9 9 9 11 13 3 13 1 0 9 11 2
16 1 10 2 9 15 3 15 13 1 9 15 13 9 9 0 2
40 3 7 2 1 9 15 0 2 9 1 9 2 11 11 7 9 9 2 9 11 2 13 13 9 11 7 13 15 2 13 1 11 13 15 7 13 11 1 11 2
15 3 9 15 3 15 13 1 9 7 9 10 3 15 13 2
14 1 11 2 11 13 1 11 11 2 15 14 3 13 2
15 15 13 10 10 9 15 3 13 13 10 9 15 13 11 2
8 3 9 9 0 10 13 15 2
20 11 13 11 11 1 9 0 1 11 1 9 9 11 7 9 13 15 13 11 2
15 11 13 10 9 1 11 11 11 11 2 11 11 2 11 2
12 1 13 1 9 11 2 15 13 1 11 11 2
16 16 11 11 13 9 15 3 0 1 9 2 11 3 13 9 2
25 11 10 13 1 9 1 9 9 9 11 11 11 7 11 11 16 13 13 11 11 11 1 11 12 2
10 10 9 15 3 13 3 13 1 9 2
32 16 16 1 9 10 13 12 12 9 15 13 1 12 12 9 15 13 2 16 9 10 13 9 2 15 9 13 9 0 0 3 2
16 1 10 9 13 2 11 13 9 1 9 15 0 1 9 15 2
31 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 13 10 9 9 0 1 9 10 2
15 1 13 1 9 2 10 11 3 13 7 13 9 9 3 2
25 9 10 13 1 9 13 12 7 3 13 9 9 2 9 9 2 7 13 1 9 0 9 2 9 2
11 3 1 9 11 1 3 13 9 0 10 2
50 3 2 11 11 10 3 0 13 1 9 11 11 1 11 11 2 1 10 13 3 9 11 11 11 11 15 3 3 13 9 11 11 2 11 11 11 1 0 15 13 13 1 9 11 2 0 11 9 2 2
9 11 3 13 9 1 9 9 9 2
39 2 12 2 9 11 13 9 9 1 9 13 2 13 9 9 1 9 2 1 9 2 9 2 9 2 9 2 9 0 2 9 7 9 2 12 2 9 9 2
33 11 11 13 9 9 1 9 15 13 1 11 7 9 2 9 0 13 9 2 0 1 9 2 9 9 9 2 9 2 9 7 9 2
16 11 2 11 11 2 11 13 9 1 11 11 11 11 2 11 2
31 1 11 12 2 11 2 11 2 7 11 3 13 9 11 11 1 13 11 1 13 11 16 13 9 1 11 7 11 1 11 2
10 11 11 0 1 9 9 1 9 11 2
24 11 9 1 13 2 9 9 13 1 9 2 9 0 2 16 14 13 9 7 9 9 15 13 2
22 1 9 3 1 9 9 15 15 13 2 11 13 16 15 13 1 10 9 15 3 0 2
49 9 9 10 15 13 1 10 9 1 10 9 1 13 10 9 9 0 1 9 2 9 1 9 1 13 9 2 9 9 2 9 2 9 2 9 9 2 9 0 2 0 2 9 2 9 9 7 9 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
6 7 7 2 11 13 2
22 11 11 2 2 13 10 9 9 9 13 11 15 13 1 9 11 3 13 1 9 9 2
87 15 0 13 1 9 12 11 11 11 1 9 11 11 11 2 11 2 11 11 2 7 11 11 11 11 7 3 13 9 9 15 1 13 9 11 2 11 11 1 9 0 11 7 3 13 12 9 13 11 11 11 11 7 11 11 11 12 15 3 13 7 13 1 10 9 0 1 11 2 11 11 2 11 11 2 11 11 2 11 2 11 11 11 2 7 11 2
2 0 2
18 2 11 11 2 1 9 1 9 9 16 13 1 9 2 9 9 11 2
13 15 3 13 2 15 13 0 1 1 9 2 11 2
21 1 10 9 13 13 9 9 12 1 9 12 2 12 2 12 2 12 2 7 12 2
16 9 9 9 0 3 13 9 9 9 9 10 15 9 12 9 2
25 1 11 2 11 13 9 13 10 9 0 1 11 2 11 11 2 7 10 9 15 0 7 9 9 2
12 11 11 13 0 1 9 7 9 15 9 0 2
7 11 9 13 1 9 9 2
12 1 12 9 9 10 2 12 9 11 3 13 2
18 11 11 15 0 1 0 13 0 9 9 2 9 12 5 10 9 9 2
17 11 13 9 9 2 11 11 2 2 1 10 9 0 15 13 0 2
27 9 9 9 13 13 1 12 2 10 7 12 2 10 16 10 9 9 7 9 7 9 9 13 1 9 0 2
23 11 11 3 2 11 11 13 9 15 1 9 2 7 15 3 3 3 13 1 11 1 9 2
21 9 10 3 13 1 13 1 9 9 2 7 1 9 1 0 2 1 13 9 9 2
18 11 13 10 10 9 1 9 11 11 2 11 11 11 2 11 2 11 2
9 11 9 13 9 9 1 9 11 2
9 16 9 15 3 13 9 9 15 2
10 7 2 14 13 9 15 13 9 10 2
11 1 12 11 12 2 9 13 1 12 12 2
3 3 9 2
18 11 3 13 16 13 1 9 2 9 2 7 11 11 1 9 9 9 2
12 9 0 9 13 10 2 9 2 1 0 9 2
11 1 15 11 0 11 11 13 1 9 10 2
10 3 10 15 13 9 2 9 15 15 2
14 1 9 11 2 3 3 13 15 13 11 3 13 9 2
26 11 11 2 15 3 13 1 13 13 9 2 15 16 3 3 15 13 13 9 7 14 13 1 11 11 2
56 1 11 2 15 13 1 10 9 9 1 11 2 11 11 2 15 3 13 1 9 1 9 9 11 2 11 3 13 13 9 1 9 1 9 9 11 2 1 10 2 11 3 13 9 0 9 2 9 11 11 2 15 13 1 9 2
14 16 9 15 13 10 9 3 13 9 9 11 7 13 2
9 1 11 13 9 2 11 3 13 2
16 11 11 7 13 2 11 11 11 11 2 7 2 11 11 2 2
16 9 10 13 1 9 12 9 9 1 9 2 9 10 13 12 2
25 1 9 12 2 11 2 11 2 7 11 2 2 15 13 13 1 11 7 13 9 1 9 7 9 2
14 11 11 3 3 0 1 13 1 10 10 9 9 11 2
12 9 9 3 13 0 9 1 9 2 9 2 2
35 9 9 13 11 11 11 11 11 11 11 11 2 11 2 16 9 9 13 2 11 11 2 2 15 13 1 11 7 13 9 1 9 12 9 2
11 11 11 13 10 10 9 15 13 9 10 2
21 1 10 9 0 2 11 11 3 13 9 0 13 9 2 9 9 13 9 7 9 2
16 10 9 14 13 9 11 11 2 16 15 13 13 1 9 0 2
31 1 9 12 2 11 11 13 16 9 0 9 11 11 13 12 5 7 12 12 1 9 9 0 15 13 1 9 15 13 9 2
22 16 11 13 9 9 15 3 3 13 2 16 13 11 7 11 2 15 3 3 13 9 2
22 3 2 1 9 0 1 9 0 9 13 2 3 3 16 10 9 3 13 9 9 9 2
10 1 1 9 9 13 1 9 1 11 2
19 1 11 0 2 11 11 13 11 11 11 1 10 10 9 9 9 1 11 2
24 9 9 10 13 1 13 9 9 11 1 11 1 13 9 9 15 13 1 9 9 9 9 11 2
12 11 3 13 1 9 0 7 1 9 11 12 2
12 11 3 13 9 1 11 7 13 9 9 10 2
14 1 9 2 9 15 13 0 10 2 13 9 1 9 2
18 11 13 10 9 9 1 9 11 2 11 11 2 11 11 11 2 11 2
6 9 9 10 3 13 2
13 1 10 1 9 9 9 2 9 2 11 11 2 2
18 11 10 13 13 11 2 11 11 12 11 12 15 13 9 1 11 11 2
21 9 9 2 15 13 1 12 9 2 3 13 16 15 13 1 10 9 15 13 11 2
17 11 9 1 9 10 13 9 1 9 0 2 10 10 13 11 11 2
22 11 12 3 13 16 11 11 13 9 1 9 9 9 13 9 9 3 9 2 9 2 2
21 13 2 13 15 13 13 11 11 11 2 13 12 9 9 15 2 9 2 7 13 2
36 10 11 1 11 13 1 11 11 13 12 9 9 15 13 11 1 2 9 9 7 9 2 9 9 0 2 7 9 11 11 7 11 15 0 2 2
22 11 13 10 10 9 2 9 9 2 11 2 1 9 9 12 2 11 11 11 11 2 2
11 15 13 3 1 9 11 2 11 7 11 2
17 11 13 16 11 3 13 1 0 1 10 10 9 9 16 9 13 2
22 9 12 2 11 11 1 12 9 13 1 9 7 1 9 12 11 11 13 13 9 11 2
21 1 9 12 11 12 11 13 1 9 11 7 1 9 12 11 12 11 13 1 9 2
19 9 9 13 1 9 1 9 9 13 1 9 9 9 1 13 7 13 3 2
12 11 0 11 11 11 7 15 0 13 11 11 2
9 3 10 9 10 13 1 11 11 2
21 3 13 13 11 13 9 9 11 11 7 11 11 2 12 9 12 9 12 11 12 2
12 9 0 9 9 11 11 1 11 13 9 11 2
32 2 12 2 9 9 1 9 11 11 1 11 11 1 13 12 11 11 1 11 2 14 1 11 12 5 11 1 9 11 11 11 2
12 11 13 10 9 2 16 11 13 1 9 11 2
24 3 11 13 1 11 11 11 7 11 11 11 11 11 11 11 11 11 2 11 2 1 11 11 2
32 16 10 9 3 13 2 2 10 9 9 2 2 7 9 9 1 9 9 3 3 13 1 9 2 9 0 2 11 11 2 2 2
9 13 2 11 11 11 13 1 9 2
14 11 2 11 13 2 7 11 13 1 13 10 9 9 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
10 11 9 10 13 9 9 11 7 11 2
23 16 10 9 9 13 2 11 3 13 9 16 9 15 13 9 10 13 2 11 2 9 11 2
24 13 0 2 15 13 1 11 2 7 1 12 2 11 13 1 11 2 16 15 3 13 9 9 2
29 11 11 13 1 12 9 11 2 12 9 11 7 12 9 0 2 15 3 13 1 9 2 9 9 15 13 11 11 2
15 11 11 11 11 13 10 9 11 15 13 1 11 11 11 2
20 11 9 10 13 3 9 15 13 2 13 7 9 9 9 15 14 3 13 0 2
19 16 11 11 11 13 9 9 2 3 9 11 13 11 11 11 1 11 11 2
16 11 9 10 13 9 1 11 11 2 15 3 13 11 7 11 2
11 11 10 13 1 9 12 1 9 11 11 2
59 11 11 11 11 11 7 11 11 11 11 11 1 11 11 11 2 13 9 1 11 11 2 11 11 11 11 2 3 11 11 2 11 11 11 11 13 1 11 11 7 11 11 11 2 11 10 13 1 11 11 11 2 16 11 11 13 1 13 2
42 11 2 0 1 11 11 11 11 11 2 13 9 9 13 1 10 9 9 9 9 12 15 13 2 13 7 13 1 11 2 11 2 0 1 11 11 11 11 11 11 2 2
25 16 14 13 3 13 0 9 15 3 0 13 0 9 11 16 15 14 3 13 9 9 1 9 10 2
8 3 9 15 13 9 15 13 2
22 3 15 13 9 11 7 11 11 11 2 16 1 9 15 13 1 11 11 16 13 13 2
90 9 1 9 9 11 11 1 13 9 9 7 13 9 9 0 1 0 7 0 13 9 0 7 13 9 9 9 11 1 9 9 2 9 9 2 9 7 9 1 13 9 7 9 9 9 11 11 11 2 9 13 1 12 9 15 13 1 11 11 11 2 9 15 3 13 1 1 9 10 13 2 9 15 13 1 1 9 10 13 2 9 15 3 13 1 1 9 10 13 2
32 11 11 11 13 1 12 9 1 11 11 11 11 2 11 11 11 13 1 12 9 1 12 9 2 16 11 11 2 11 7 11 2
17 9 0 9 9 13 1 9 15 13 1 9 9 15 13 3 0 2
21 9 11 11 11 3 13 1 11 1 9 9 9 15 13 1 11 2 11 11 2 2
17 11 11 13 12 9 1 9 12 9 7 12 9 1 9 12 11 2
7 9 9 1 9 0 9 2
9 11 3 13 1 9 11 2 11 2
11 11 13 9 7 13 1 11 11 2 11 2
43 11 11 11 11 2 2 13 11 2 13 9 9 9 1 11 2 7 13 9 1 2 11 13 9 11 1 9 12 7 13 9 1 9 9 1 11 7 10 9 15 3 0 2
14 12 9 15 13 1 9 0 3 13 9 1 9 0 2
12 9 9 1 9 9 9 10 13 1 9 11 2
26 3 2 3 1 10 15 13 1 11 11 2 11 11 11 2 11 11 11 2 11 11 11 11 3 11 2
16 16 15 13 10 10 1 13 9 2 9 9 15 14 3 13 2
17 15 13 1 11 2 13 1 11 2 16 15 13 9 1 11 11 2
22 11 15 13 7 10 13 2 15 15 3 13 11 11 2 7 1 9 9 15 3 13 2
9 11 15 0 7 13 3 1 11 2
22 15 13 1 9 11 7 11 2 11 1 9 12 2 13 9 11 2 11 1 9 9 2
19 1 9 12 11 12 2 11 13 9 13 11 12 13 11 11 11 11 11 2
48 3 13 9 9 9 12 9 2 9 2 9 13 13 9 0 9 3 11 2 7 11 11 2 11 2 11 2 2 9 11 11 2 11 1 9 11 15 13 1 12 2 12 2 9 1 12 9 2
23 11 3 13 1 9 2 9 9 11 7 9 15 0 9 13 9 13 11 11 1 9 12 2
17 13 13 9 9 1 9 9 10 2 16 11 13 3 13 7 13 2
8 15 13 1 11 11 11 11 2
11 3 15 13 15 12 13 12 3 13 12 2
10 1 9 2 15 13 9 0 11 11 2
9 15 3 13 3 9 15 3 13 2
28 1 11 12 2 10 9 1 9 9 1 11 2 1 12 5 1 9 11 2 13 7 9 13 13 1 9 12 2
8 11 13 9 9 1 9 11 2
25 11 2 1 11 2 7 11 1 11 2 13 10 9 1 9 11 2 15 3 2 3 13 10 9 2
48 15 3 13 9 2 9 13 1 9 3 2 11 2 1 11 2 7 9 1 9 16 9 2 9 15 13 9 0 15 0 2 9 2 2 3 13 9 7 9 2 9 16 9 2 9 10 13 2
17 9 15 13 3 2 3 13 0 16 9 3 13 0 1 9 9 2
17 11 11 11 11 12 13 10 9 9 9 11 15 13 1 9 12 2
19 3 11 13 9 10 1 9 1 2 12 7 13 1 1 11 11 1 12 2
16 13 11 2 11 1 10 9 9 13 9 2 9 9 0 0 2
9 12 12 9 3 9 0 13 13 2
40 11 13 9 1 12 12 9 7 11 11 11 1 9 2 7 13 16 9 11 1 9 2 9 11 3 13 1 0 15 13 7 2 3 1 9 7 13 9 2 2
10 1 11 3 13 1 9 7 13 9 2
10 9 9 10 1 0 13 11 13 9 2
43 9 10 3 9 9 1 9 15 3 13 9 11 2 9 9 0 13 9 2 12 10 13 9 15 3 0 2 16 3 13 3 1 12 9 9 2 12 1 9 15 3 0 2
19 9 10 3 0 2 3 13 1 9 1 9 9 7 9 9 2 11 11 2
23 11 13 9 10 10 9 15 13 1 11 11 11 11 2 11 11 2 11 11 11 2 11 2
13 15 13 11 11 1 9 9 1 9 12 11 12 2
19 11 11 11 13 9 1 9 11 1 9 11 15 13 1 13 9 9 0 2
10 9 10 13 9 10 9 0 1 11 2
6 11 13 9 11 11 2
19 9 11 11 11 12 10 13 9 1 11 11 11 12 15 3 13 9 0 2
13 9 10 13 9 1 12 9 13 1 9 11 0 2
17 11 3 3 13 9 0 9 11 11 1 11 3 13 1 11 11 2
17 9 15 3 0 7 0 9 9 15 3 0 13 1 9 9 9 2
13 11 12 5 11 11 13 9 0 11 12 5 11 2
32 1 9 12 2 9 10 13 9 9 1 12 9 7 13 9 9 12 12 2 2 9 10 13 9 9 9 12 9 5 12 2 2
17 11 13 9 10 7 13 1 13 9 10 2 7 7 9 14 13 2
17 11 13 9 15 13 1 9 11 2 11 11 2 11 11 2 11 2
9 15 3 13 3 13 9 1 9 2
13 11 11 2 2 13 10 9 9 9 9 1 11 2
15 10 13 9 1 9 12 11 2 11 2 11 11 11 11 2
13 3 0 11 13 9 9 2 1 15 3 10 9 2
9 9 10 13 1 12 1 11 11 2
20 11 2 11 11 2 12 2 12 2 2 13 9 9 9 1 13 13 1 9 2
63 1 12 2 11 13 1 1 9 12 1 11 11 12 2 13 9 1 11 2 12 2 1 9 15 13 9 1 10 9 11 2 1 1 11 2 15 3 13 1 1 11 11 2 10 13 9 11 1 13 9 9 7 13 9 0 15 13 13 9 2 11 2 2
9 7 15 15 3 13 9 1 11 2
22 1 13 1 9 9 1 9 2 15 3 13 1 9 13 9 9 1 10 9 7 9 2
11 16 2 9 3 15 13 1 9 9 0 2
9 11 7 9 9 13 1 9 9 2
46 11 15 13 1 9 9 13 11 11 11 11 2 9 10 13 1 9 12 7 3 13 10 0 9 15 0 1 1 11 12 11 7 11 11 2 1 9 9 10 13 9 0 1 9 12 2
28 16 9 1 9 13 9 15 3 0 2 16 9 13 14 13 1 11 2 11 2 15 3 13 9 10 2 13 2
34 15 13 1 12 3 1 9 11 11 11 2 7 16 1 9 0 1 9 0 2 11 2 15 13 9 1 13 1 10 9 15 14 0 2
21 2 16 11 13 7 13 1 9 2 2 9 9 15 1 9 15 0 3 13 10 2
14 11 13 0 1 9 2 13 9 9 13 11 1 11 2
19 1 9 12 2 9 9 11 13 1 3 13 0 13 9 1 12 11 12 2
22 9 10 13 1 12 2 12 13 9 1 9 12 2 12 2 5 12 7 9 14 13 2
25 3 10 9 0 1 11 13 7 13 1 11 2 11 0 11 13 1 11 11 11 11 11 1 11 2
8 1 9 12 15 13 9 9 2
18 15 13 12 9 11 2 13 9 1 0 2 7 3 13 1 11 11 2
14 11 13 9 11 1 11 11 11 11 1 12 2 12 2
18 11 11 11 13 10 9 9 1 11 11 15 13 9 0 9 9 9 2
33 11 9 0 15 13 9 10 2 13 11 2 11 2 11 11 2 11 2 11 2 11 2 11 5 11 2 11 2 11 2 7 9 2
15 11 3 13 1 0 1 9 9 9 15 13 1 9 0 2
12 3 13 11 11 11 11 3 0 1 9 11 2
19 7 9 9 3 11 2 11 2 11 7 11 9 9 10 13 1 11 11 2
23 15 13 0 16 13 1 9 0 1 11 11 11 11 11 11 2 15 13 1 11 2 11 2
15 11 11 11 11 2 11 11 11 11 11 11 11 2 11 2
25 1 9 12 2 16 13 9 9 2 9 1 9 13 9 9 1 9 9 0 7 13 9 13 9 2
22 11 11 2 13 9 9 9 15 13 1 11 11 7 11 11 11 1 9 9 9 3 2
29 11 9 10 13 1 0 9 11 11 2 11 2 13 1 11 2 11 7 13 9 9 0 7 0 1 9 11 11 2
7 11 3 0 1 9 11 2
11 1 9 12 9 10 13 9 1 12 9 2
18 11 9 13 9 1 13 9 9 9 15 13 1 9 11 2 11 11 2
18 16 15 13 7 13 11 13 1 1 9 2 16 9 9 0 3 13 2
63 11 9 15 13 1 13 9 12 11 12 0 13 1 9 2 9 13 2 16 2 11 11 11 11 2 11 5 11 11 2 11 11 11 2 11 11 7 11 7 11 11 12 5 11 11 11 12 2 15 13 1 13 9 9 5 9 2 9 9 7 9 0 2
22 15 12 9 13 1 9 11 1 9 9 12 13 11 15 3 3 13 11 1 10 9 2
30 1 9 0 1 12 9 2 11 13 9 1 9 2 9 0 2 3 1 11 11 2 13 9 11 2 11 2 7 11 2
23 9 10 13 1 9 10 11 16 11 13 11 2 13 10 10 11 2 1 9 9 1 11 2
22 11 11 13 10 10 9 15 13 1 9 11 2 9 11 11 2 9 11 11 2 11 2
17 11 11 11 7 11 11 2 11 7 11 2 13 9 9 11 11 2
24 9 15 13 1 0 12 9 13 0 2 9 9 2 9 0 7 9 0 2 9 7 9 11 2
21 11 11 15 0 1 9 0 13 9 9 7 9 15 13 1 9 0 3 0 13 2
12 16 9 3 13 7 3 13 9 9 1 9 2
57 11 11 11 13 3 0 1 9 9 7 9 2 9 11 7 11 13 3 0 1 9 9 7 9 0 0 1 9 9 2 9 0 9 13 9 15 0 3 13 1 12 9 2 9 2 9 7 9 2 9 0 1 9 13 9 10 2
26 1 9 9 13 2 11 13 9 9 1 9 9 7 15 9 10 13 3 3 0 7 0 9 13 11 2
22 1 9 11 2 11 13 16 9 2 9 11 2 7 2 9 11 2 13 1 9 0 2
82 1 10 9 2 11 2 11 11 2 7 11 11 2 11 13 1 9 2 9 0 15 9 3 13 1 9 11 2 1 1 10 9 9 2 9 0 2 13 9 2 9 15 13 1 9 11 1 0 3 13 1 9 1 11 1 10 9 15 13 9 2 15 13 1 2 11 11 2 15 13 1 11 12 2 12 2 11 12 7 11 12 2
13 3 9 2 9 13 9 9 1 9 9 2 9 2
17 11 11 3 13 9 1 11 11 15 13 1 10 9 9 7 9 2
14 9 9 9 9 13 1 9 9 9 2 9 7 9 2
163 2 11 11 2 2 2 1 9 1 15 2 7 1 15 1 9 2 2 9 9 9 13 11 2 11 11 11 15 13 2 13 12 9 0 1 9 2 13 12 9 9 11 2 3 2 3 9 9 14 9 2 2 2 1 10 9 0 7 9 2 3 13 9 9 1 11 11 15 3 2 3 9 10 3 13 9 9 9 1 9 7 9 9 3 2 3 1 3 13 2 7 13 9 0 1 9 3 15 13 2 2 2 9 2 9 1 9 9 2 0 9 7 0 2 0 11 11 2 11 2 12 11 2 11 2 11 2 11 2 11 2 11 11 2 2 12 2 12 2 12 11 2 2 12 2 12 11 11 11 11 13 3 12 9 2 13 9 11 2 15 3 0 2
7 9 1 0 13 9 9 2
27 11 9 0 2 7 9 0 2 13 9 9 11 11 15 3 13 9 12 9 2 7 9 9 1 12 9 2
12 11 2 11 11 13 11 11 9 12 2 12 2
8 9 13 13 12 9 9 0 2
17 9 10 13 9 16 11 13 9 10 16 9 13 9 1 10 9 2
23 11 2 9 2 9 2 13 1 11 11 2 11 2 1 12 9 2 11 13 12 9 2 2
17 11 13 9 9 11 1 9 9 7 9 11 2 15 13 1 11 2
6 15 15 3 13 11 2
13 11 13 11 1 9 11 2 7 11 1 9 11 2
8 9 3 12 9 0 9 10 2
10 3 15 13 9 0 1 9 13 11 2
23 9 9 11 11 13 1 12 9 15 3 13 1 1 12 9 9 9 11 2 1 1 3 2
15 11 13 1 11 7 1 0 13 1 9 2 9 0 11 2
11 11 11 3 13 9 9 1 11 11 12 2
44 11 7 9 11 2 2 13 9 2 9 15 13 9 1 9 13 9 1 9 9 1 9 7 9 9 0 2 7 3 13 9 7 9 1 13 9 15 3 0 7 13 13 9 2
11 3 11 3 13 1 9 9 7 9 9 2
10 11 11 13 12 9 9 1 9 10 2
28 11 11 3 3 13 11 11 2 11 11 2 9 11 7 10 9 2 9 0 13 11 11 11 11 7 11 11 2
15 11 11 13 10 9 15 13 1 11 2 11 2 11 11 2
75 1 9 12 11 12 2 12 9 11 0 13 7 3 1 12 9 0 13 1 11 11 11 1 9 11 11 11 11 12 2 16 10 9 15 13 1 9 1 9 11 11 11 16 15 3 3 13 9 12 9 11 11 11 11 1 11 11 11 2 7 15 3 13 1 9 9 1 9 11 2 11 11 2 11 2
24 11 13 10 10 11 15 13 1 11 11 11 2 11 11 2 11 11 11 2 11 11 2 11 2
13 11 3 13 1 9 15 13 3 11 14 3 13 2
8 3 15 3 13 15 1 13 2
10 10 9 11 13 1 9 0 2 11 2
24 15 15 3 13 15 11 2 10 9 15 13 3 13 13 1 9 0 1 9 9 9 2 11 2
14 10 9 3 2 9 10 3 13 7 3 13 9 15 2
22 11 7 11 13 1 13 0 1 11 9 12 2 16 15 13 1 11 13 11 7 11 2
13 9 10 13 1 9 9 15 13 1 3 7 0 2
16 3 3 9 15 13 1 9 12 13 12 9 13 1 9 12 2
11 15 14 13 9 7 13 9 0 15 0 2
15 3 11 8 3 13 10 10 7 3 3 13 9 15 0 2
22 3 11 11 3 13 9 1 11 2 3 13 10 9 0 1 9 7 13 9 11 13 2
16 9 13 13 7 13 9 7 15 13 1 9 9 3 9 13 2
8 9 11 13 1 0 7 0 2
9 3 11 3 13 1 10 9 9 2
12 15 13 11 11 11 7 13 13 9 11 11 2
4 11 9 10 2
3 3 13 2
8 11 11 13 9 1 12 12 2
20 9 11 15 13 1 12 9 9 13 1 11 11 11 11 11 11 2 11 2 2
22 12 11 11 11 13 10 9 9 0 9 12 15 13 13 9 12 1 11 2 11 11 2
31 1 9 15 0 9 15 13 13 1 9 2 9 7 9 0 1 9 10 2 10 2 0 1 9 11 1 9 11 0 2 2
26 11 13 9 15 13 1 13 9 15 13 2 13 2 13 7 13 0 1 9 9 15 13 3 15 13 2
30 7 9 9 1 9 11 11 7 10 9 9 1 11 5 11 7 10 11 1 10 11 3 13 11 14 3 13 9 10 2
27 11 11 2 11 2 11 11 13 10 10 11 11 11 11 15 13 1 11 11 11 2 11 11 11 2 11 2
31 11 11 11 13 9 9 11 15 13 1 12 9 12 15 13 1 11 11 7 13 1 11 11 2 11 11 2 7 11 11 2
11 11 13 1 11 2 9 10 13 1 12 2
18 11 2 15 3 13 3 0 9 2 7 9 9 2 11 2 11 11 2
12 11 1 9 9 2 7 11 1 9 9 9 2
26 13 9 11 11 11 2 11 2 1 11 11 11 11 11 1 9 9 9 9 2 11 2 9 9 12 2
15 11 3 13 1 13 1 11 7 11 13 1 9 9 11 2
96 11 9 15 3 13 16 11 14 9 15 3 13 1 9 2 13 9 12 2 11 11 7 9 12 2 11 11 2 11 11 1 13 9 11 2 1 9 0 12 2 11 13 15 1 11 11 2 11 11 11 2 2 15 13 9 0 1 11 0 2 15 3 13 10 9 9 11 2 11 13 16 15 3 0 7 3 0 1 9 2 9 9 1 11 2 15 13 11 2 9 9 9 2 1 9 2
36 9 9 9 15 13 1 9 3 13 13 9 1 9 12 7 9 9 13 1 12 9 2 12 9 2 13 12 9 2 12 9 2 1 9 12 2
5 3 13 1 9 2
20 1 9 15 13 11 11 15 0 2 0 2 15 0 13 1 11 11 11 11 2
44 11 11 11 11 13 12 5 1 9 11 11 1 11 11 2 11 9 10 14 3 0 1 9 0 1 11 2 16 9 9 10 13 9 11 2 11 2 11 11 11 2 7 11 2
31 9 0 9 13 9 15 13 1 0 1 9 1 9 0 7 0 1 10 9 2 7 1 9 0 0 7 9 9 0 0 2
11 1 9 10 2 11 13 9 1 12 9 2
12 15 14 13 9 13 9 3 13 1 9 9 2
18 11 11 11 13 9 1 9 11 11 2 11 11 11 2 11 2 11 2
29 9 9 9 3 13 1 9 11 1 13 7 13 9 1 10 9 7 9 15 13 2 3 3 13 1 10 9 9 2
25 11 11 11 2 11 3 13 9 2 9 11 7 11 2 1 9 9 11 11 2 2 16 13 9 2
9 1 9 12 2 9 13 12 9 2
12 16 13 11 11 2 1 9 13 7 3 9 2
24 1 9 11 3 13 1 10 9 1 11 11 2 11 11 2 11 11 2 11 11 7 3 9 2
18 15 3 13 1 9 15 13 9 2 7 16 9 13 7 15 3 13 2
29 1 1 15 15 13 1 2 11 3 13 9 1 11 11 11 11 2 11 2 10 9 9 15 3 13 13 9 9 2
43 9 1 9 9 11 2 1 9 12 2 9 10 13 9 9 3 12 9 7 13 9 9 12 2 12 12 2 2 9 10 13 9 9 9 1 12 2 12 9 5 12 2 2
26 1 13 1 11 2 11 13 9 9 11 9 7 9 9 11 11 15 0 1 9 2 11 11 11 2 2
14 10 0 1 9 2 9 10 13 1 9 12 2 12 2
15 1 9 11 2 13 9 7 10 9 13 10 9 7 9 2
11 1 9 9 2 11 11 13 9 1 11 2
15 11 12 1 11 9 10 13 0 9 9 12 9 9 9 2
18 16 13 1 11 2 11 3 13 7 13 12 10 9 2 11 7 11 2
25 11 11 11 11 13 0 1 9 11 11 15 13 1 1 9 2 16 15 14 13 1 13 9 10 2
18 11 13 10 9 15 3 13 1 9 11 11 1 9 9 7 9 9 2
15 1 12 2 15 13 9 11 11 11 2 11 2 1 9 2
26 11 2 9 2 13 9 12 2 7 9 2 11 11 2 11 11 2 7 14 3 13 1 9 11 0 2
26 16 14 2 9 1 13 3 3 13 9 13 15 1 10 9 0 7 9 9 0 15 3 13 9 10 2
42 11 11 11 13 9 9 9 11 11 9 9 11 11 2 9 13 0 0 10 13 1 12 11 12 7 13 1 0 11 11 2 11 11 2 11 11 2 7 3 3 0 2
40 11 2 11 2 11 11 2 2 13 9 11 15 13 7 3 9 9 9 9 13 11 2 11 2 11 2 11 11 13 9 1 9 2 9 2 11 1 11 11 2
3 11 13 2
30 16 2 9 15 13 1 9 10 13 1 11 11 16 14 13 13 1 9 15 13 9 2 9 2 9 2 7 9 9 2
12 9 9 9 13 1 9 9 7 9 9 9 2
35 9 1 9 15 14 0 13 9 9 15 3 0 2 9 9 1 9 9 2 9 3 0 7 0 7 9 0 2 7 13 9 9 15 0 2
22 1 1 9 13 10 9 2 9 1 9 2 9 9 2 11 11 7 11 11 3 0 2
24 1 9 11 9 10 2 11 3 3 13 13 1 11 2 16 9 3 13 15 0 1 9 9 2
32 13 13 9 9 1 9 11 1 12 9 9 2 1 12 9 12 1 12 11 12 9 12 9 11 11 13 9 9 9 2 9 2
28 11 7 11 13 16 11 11 13 9 16 9 13 9 9 2 7 10 9 0 3 13 9 15 0 1 13 9 2
9 15 3 13 11 11 15 13 9 2
11 11 9 15 14 13 9 10 13 13 9 2
19 11 11 1 9 9 10 13 1 12 9 7 13 1 9 9 7 9 0 2
20 16 1 9 10 9 3 13 9 2 16 9 9 3 13 1 9 9 1 9 2
18 11 11 13 10 10 9 9 15 13 1 11 7 13 1 9 9 9 2
15 1 9 11 12 3 2 15 13 13 12 5 9 11 11 2
13 3 9 10 13 0 1 9 9 1 9 7 11 2
82 16 9 13 9 9 9 16 9 10 3 13 9 15 0 1 9 15 1 13 13 11 11 2 12 11 12 9 12 2 14 13 9 9 1 9 9 0 9 2 9 9 2 9 9 2 9 2 11 9 7 9 9 9 2 9 9 7 9 9 2 7 9 9 9 7 9 9 2 9 9 0 2 7 9 2 9 15 13 10 9 2 2
9 11 13 1 9 9 11 1 11 2
21 11 11 2 11 11 7 11 11 1 11 11 2 7 11 11 1 5 11 2 11 2
21 11 15 0 7 9 15 9 7 9 9 12 9 13 9 15 3 13 1 9 9 2
14 11 13 9 1 11 10 2 11 2 11 11 2 11 2
4 3 9 0 2
12 16 16 9 9 11 11 11 13 9 9 10 2
27 1 10 3 9 9 1 9 9 1 11 7 11 7 9 9 3 13 9 1 9 9 7 13 9 9 9 2
33 12 9 2 11 2 11 2 11 2 11 7 11 2 13 9 1 11 11 11 2 9 15 3 0 2 1 1 9 13 9 9 9 2
16 1 9 12 2 1 9 9 2 3 9 10 13 1 9 11 2
47 1 1 9 11 2 11 11 11 7 11 11 11 2 11 11 2 13 9 9 11 11 2 15 13 13 1 2 9 10 13 1 9 16 1 9 0 9 9 1 11 1 9 11 11 13 13 2
10 3 0 10 10 13 1 9 11 11 2
9 15 3 0 2 16 3 3 13 2
25 1 9 9 9 12 2 16 9 14 13 9 2 9 0 3 13 1 9 9 9 11 15 3 13 2
30 3 11 13 11 13 1 9 9 11 11 2 7 15 13 9 1 13 1 9 9 7 15 13 16 15 13 9 9 9 2
17 9 0 14 13 2 16 11 11 11 11 13 2 16 13 1 9 2
24 11 2 11 2 3 13 1 11 7 11 2 13 9 7 9 0 12 1 9 11 2 11 11 2
14 1 13 9 15 13 2 10 9 3 13 9 13 9 2
49 11 11 11 11 7 13 13 11 11 13 10 9 13 9 13 9 15 13 9 9 1 9 1 9 15 3 0 2 0 1 13 2 7 3 0 1 13 1 9 15 13 1 1 9 9 14 3 13 2
18 9 9 9 13 1 13 9 15 13 1 9 9 9 1 9 9 9 2
14 3 2 9 9 11 13 7 13 9 9 1 9 10 2
16 15 15 3 13 1 9 15 15 3 13 1 9 9 1 15 2
20 9 11 11 13 13 9 16 1 9 10 9 9 9 1 11 3 13 15 13 2
29 11 11 13 2 11 11 11 2 11 2 7 3 2 11 2 13 1 13 12 9 13 1 9 9 15 1 11 11 2
14 9 2 9 0 3 13 1 9 2 9 9 11 11 2
20 9 10 13 12 11 12 2 12 9 16 11 2 11 11 13 1 12 11 12 2
17 12 9 13 1 0 2 7 3 9 3 13 12 12 2 14 13 2
39 16 3 1 9 2 9 9 15 13 1 9 0 3 3 13 9 9 1 9 9 0 1 2 11 2 11 2 11 2 11 11 11 2 11 2 11 7 11 2
15 10 3 9 1 9 15 13 1 9 1 9 13 9 9 2
12 15 13 1 9 16 15 13 9 0 1 9 2
65 13 1 9 1 9 9 1 11 2 11 11 11 2 11 12 1 9 12 1 12 9 2 11 2 11 2 11 2 11 11 11 2 11 2 7 11 2 1 9 1 13 9 2 9 9 9 9 9 15 13 9 15 13 7 13 13 1 13 9 1 9 1 9 9 2
16 9 9 11 14 0 2 16 13 9 1 11 3 0 7 14 2
24 1 10 9 9 15 0 2 11 3 2 3 13 9 0 1 13 9 2 11 2 9 9 13 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
48 3 9 9 7 9 9 15 13 2 16 13 12 9 11 11 2 3 2 1 11 2 13 12 9 9 11 11 2 3 2 1 9 0 1 11 2 10 9 9 0 1 11 2 13 9 13 1 2
14 11 13 13 9 9 9 1 11 11 1 11 11 12 2
47 3 1 12 11 12 11 2 13 9 2 1 9 9 7 13 1 11 11 11 2 12 5 11 5 12 1 11 11 11 11 1 11 11 2 9 11 13 1 12 9 1 0 1 12 11 12 2
10 11 11 11 2 11 11 11 11 2 11
38 9 0 0 13 9 10 13 1 9 9 7 9 9 9 9 11 2 1 9 10 9 10 13 13 9 9 9 9 10 9 11 13 10 9 7 9 9 2
31 1 9 2 13 9 1 10 9 10 2 1 1 9 9 2 9 3 13 1 3 0 2 3 1 9 2 9 0 7 0 2
19 11 11 1 9 16 13 1 9 2 9 9 3 13 9 0 1 9 11 2
11 10 9 13 1 9 2 10 3 1 11 2
21 15 13 1 11 2 11 11 11 12 2 7 15 3 13 9 1 9 9 1 9 2
18 11 10 2 15 13 1 9 9 11 11 2 13 9 9 1 9 9 2
5 3 13 9 9 2
39 11 3 13 1 9 9 12 1 9 0 1 9 12 2 1 11 12 11 11 9 11 2 11 2 13 13 9 9 15 1 9 0 1 9 0 1 12 9 2
12 9 9 15 0 3 13 9 15 0 7 0 2
19 7 11 13 2 2 11 11 2 15 13 10 9 7 9 7 3 9 9 2
