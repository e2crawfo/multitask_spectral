349 17
14 12 9 2 1 12 9 2 12 8 7 3 13 9 2
16 10 0 9 1 9 8 1 10 0 9 13 3 3 0 3 2
24 2 6 2 3 4 15 15 3 3 0 3 2 2 13 15 3 1 10 9 1 11 1 8 2
10 1 10 9 1 11 13 11 0 3 2
6 15 13 1 12 9 2
23 1 15 12 11 1 11 2 13 11 11 0 1 12 7 13 10 13 9 3 3 1 12 2
21 2 10 9 1 11 4 10 0 9 2 2 13 11 2 15 9 15 9 8 13 2
10 2 15 4 3 3 4 16 15 13 2
18 15 13 1 10 0 9 1 8 0 3 10 9 4 1 10 15 9 2
12 10 9 13 1 13 2 13 7 3 3 13 2
24 3 13 3 15 4 16 15 9 7 15 9 1 15 13 8 1 11 1 11 0 1 13 2 2
9 3 13 15 1 4 1 15 9 2
60 7 10 0 9 1 11 13 3 8 9 3 1 10 0 9 1 11 1 15 9 2 10 3 13 9 1 11 2 10 9 1 10 0 9 13 9 2 10 13 9 7 15 13 1 10 9 0 9 1 10 9 11 11 2 11 2 8 7 11 2
17 9 4 16 11 1 10 13 7 0 9 3 15 13 9 13 4 2
19 2 3 13 15 1 9 10 0 9 1 10 9 2 2 13 15 0 0 2
14 2 3 4 11 0 3 15 0 16 15 15 13 2 2
13 3 13 1 10 9 2 9 4 2 1 15 9 2
24 10 0 9 2 1 9 8 0 1 0 9 7 9 11 3 1 10 9 2 13 3 3 8 2
15 6 2 2 3 13 15 3 3 1 10 9 1 12 9 2
23 15 13 15 3 0 1 10 9 2 7 15 13 3 1 10 9 16 8 1 15 9 13 2
27 1 9 13 10 0 9 3 0 3 2 7 1 3 13 9 2 16 3 11 2 13 15 3 3 3 3 2
17 3 13 3 1 8 0 9 1 10 9 7 4 15 13 4 2 2
15 3 13 4 10 9 1 10 9 1 10 0 9 1 11 2
40 1 10 0 9 1 9 11 7 0 9 1 0 9 11 13 3 0 15 9 2 9 7 9 1 10 0 9 1 11 2 1 3 10 0 9 1 10 0 9 2
17 1 10 9 1 11 13 10 9 1 11 3 12 9 1 12 9 2
13 1 10 9 1 11 4 10 9 3 3 15 0 2
24 11 13 11 0 12 9 2 3 13 12 9 2 1 8 7 11 2 1 10 9 1 12 9 2
17 2 3 3 4 10 0 9 10 0 1 15 9 2 2 13 11 2
16 11 13 10 0 9 1 10 9 1 15 0 8 1 12 4 2
6 11 13 10 0 9 2
10 3 1 12 9 13 11 10 9 3 2
9 1 10 0 9 13 11 10 9 2
14 10 0 9 13 10 3 0 2 7 3 0 9 3 2
6 11 13 3 0 3 2
8 9 4 1 10 0 9 0 2
7 3 15 9 4 8 4 2
11 11 13 3 7 13 10 9 1 11 0 2
9 13 9 4 10 11 1 15 8 2
10 10 9 1 11 13 15 0 9 4 2
19 10 9 1 10 11 13 1 10 9 1 11 15 15 1 11 4 2 12 2
11 10 9 13 3 3 0 1 10 9 4 2
9 12 9 4 3 1 10 11 4 2
11 1 8 4 11 10 0 9 1 4 4 2
17 10 0 9 4 10 0 9 1 10 9 1 11 2 8 15 8 2
8 11 13 12 9 1 11 3 2
7 11 13 10 9 1 12 2
8 11 13 1 10 9 1 11 2
11 10 9 13 15 9 1 10 9 1 11 2
11 10 9 1 8 13 1 9 12 9 4 2
9 10 9 13 16 1 0 9 4 2
11 1 10 9 1 8 7 8 13 15 8 2
23 16 10 9 1 11 1 9 4 4 2 13 9 1 10 9 15 9 1 10 9 1 4 2
28 11 7 11 13 15 3 16 0 9 1 10 9 4 1 10 9 1 10 11 9 2 13 9 1 11 7 11 2
18 11 13 1 12 1 11 2 11 13 15 1 9 1 8 2 12 2 2
16 10 9 11 7 11 7 9 11 13 3 3 10 9 1 9 2
18 12 13 10 0 9 1 10 0 9 1 10 9 1 8 1 12 4 2
7 10 11 4 11 1 11 2
8 10 0 9 13 8 1 8 2
14 10 0 9 13 1 9 1 8 2 12 2 7 8 2
8 8 13 10 9 1 11 13 2
8 8 13 15 9 1 11 4 2
28 15 13 10 0 9 3 3 16 11 2 16 0 9 13 2 15 1 15 9 1 9 8 1 10 9 13 4 2
7 2 15 4 15 9 9 2
9 15 13 15 3 3 15 4 4 2
15 15 13 10 9 10 0 9 1 4 1 15 7 15 9 2
14 10 9 1 11 4 3 0 2 7 3 10 0 2 2
11 11 13 1 10 9 1 12 4 1 11 2
15 10 9 13 1 10 0 9 1 10 9 2 13 1 11 2
12 15 4 10 0 9 1 10 0 0 9 8 2
19 1 10 9 13 11 2 13 9 1 10 0 11 2 3 0 1 10 9 2
17 10 9 13 3 0 2 7 3 13 11 2 0 2 1 9 0 2
15 3 10 0 12 9 1 10 0 9 13 15 1 10 9 2
13 11 13 9 8 16 8 16 0 9 0 1 4 2
14 10 0 9 1 11 13 1 10 9 10 0 9 9 2
20 0 9 1 10 0 9 13 3 16 11 10 0 9 4 16 8 3 1 13 2
13 10 9 4 16 12 9 3 1 15 9 1 4 2
15 8 13 10 9 0 9 4 3 1 4 1 10 0 9 2
19 15 13 16 10 9 15 15 4 4 7 3 13 9 3 3 4 4 4 2
9 8 13 15 1 11 3 1 8 2
11 11 13 15 1 10 9 3 1 10 9 2
16 16 0 9 11 1 11 16 0 9 11 13 3 9 1 4 2
18 11 4 12 9 9 1 11 2 3 15 1 8 1 10 0 9 13 2
15 3 4 15 9 3 3 8 4 1 0 9 2 3 0 2
10 8 4 3 1 8 10 0 9 4 2
20 9 2 9 2 9 7 9 13 13 11 3 1 10 9 1 10 11 1 11 2
12 3 12 0 9 7 9 4 1 10 9 4 2
19 10 12 9 13 15 10 15 9 1 10 9 2 8 2 0 7 0 2 2
13 8 1 11 13 10 9 1 11 2 9 13 9 2
15 8 1 15 8 2 9 1 0 9 2 13 10 9 3 2
9 10 9 4 4 1 10 0 9 2
32 9 7 9 13 1 11 4 1 10 9 1 10 9 1 10 9 1 10 9 1 10 12 0 9 7 11 2 9 2 1 11 2
21 3 1 0 9 2 7 1 9 7 13 13 10 0 15 9 1 10 9 4 4 2
25 2 1 1 13 13 15 10 0 0 9 4 2 2 13 10 0 9 8 1 8 2 9 1 0 2
25 2 15 4 3 10 9 16 10 9 1 10 11 3 1 4 1 9 1 15 15 15 9 13 2 2
23 10 2 9 2 1 10 0 13 3 8 1 10 9 1 9 1 10 9 1 10 0 9 2
39 3 13 10 9 2 9 7 9 2 15 0 9 1 0 9 2 9 1 10 9 7 10 9 1 9 2 8 4 2 13 10 9 8 2 15 1 10 9 2
22 10 0 13 4 1 10 0 9 1 10 9 1 10 0 9 1 10 0 1 13 4 2
36 10 9 1 10 9 13 10 9 1 10 0 9 7 4 3 1 9 8 16 15 8 10 0 10 9 1 10 2 9 1 10 9 2 1 4 2
39 2 15 13 16 9 1 0 9 2 15 4 4 16 15 9 7 10 9 1 15 9 1 4 2 3 1 9 7 9 4 4 2 2 13 8 1 15 8 2
25 10 9 13 15 1 9 8 4 1 10 9 1 10 0 9 8 2 15 0 9 1 11 4 4 2
26 15 9 13 0 1 13 1 9 1 15 9 1 10 13 9 8 10 9 3 15 16 9 1 11 13 2
16 9 8 1 11 13 1 8 10 9 1 10 0 8 10 11 2
12 15 13 1 15 3 10 0 9 1 10 9 2
28 15 13 3 1 4 16 15 15 9 8 4 4 1 15 13 1 10 9 1 10 13 9 9 1 10 13 9 2
23 8 2 9 1 10 0 9 1 11 2 1 10 9 1 11 2 13 11 10 9 9 4 2
13 11 13 15 13 12 9 7 12 9 0 1 4 2
11 10 0 9 13 1 12 9 7 12 9 2
12 10 0 9 13 3 1 10 9 1 15 8 2
12 1 10 9 13 10 9 9 4 1 15 9 2
13 11 11 13 10 9 1 9 2 1 10 9 11 2
14 15 13 10 9 11 1 10 9 1 11 1 10 9 2
17 10 9 13 15 3 4 2 15 9 4 7 0 16 12 9 4 2
15 3 4 15 4 16 3 1 10 12 9 10 9 1 4 2
16 15 12 13 13 1 10 9 1 10 9 16 11 10 9 4 2
18 9 8 13 1 15 9 2 8 2 15 8 1 15 13 13 9 4 2
8 13 9 8 13 10 8 9 2
16 10 9 1 10 12 9 9 1 11 13 10 9 1 15 8 2
27 8 1 15 8 1 11 2 15 13 1 9 1 8 2 4 1 10 9 10 0 9 15 1 10 9 13 2
5 15 13 12 9 2
18 8 1 10 9 1 15 8 13 16 10 3 13 9 1 10 9 12 2
21 15 13 16 12 9 3 12 9 9 7 10 9 0 0 9 1 11 7 15 8 2
21 16 1 10 9 10 9 13 2 13 10 9 15 3 1 1 11 2 11 7 11 2
20 10 9 1 11 13 3 1 15 9 1 11 1 11 9 1 12 7 12 9 2
8 9 13 3 0 1 9 3 2
24 10 9 1 15 15 9 4 10 9 1 10 0 9 1 10 9 1 10 9 1 9 7 9 2
14 15 9 13 15 9 15 12 9 7 12 9 7 0 2
38 10 0 9 13 10 9 9 1 11 2 11 7 11 16 1 13 16 10 9 9 15 1 10 12 9 1 0 9 1 15 9 13 2 0 0 4 4 2
24 3 13 10 9 1 11 1 10 0 9 12 13 2 7 13 1 11 7 11 3 12 9 0 2
24 15 1 15 13 10 0 9 4 1 15 7 15 9 1 9 7 9 9 1 10 9 4 13 2
25 15 9 4 3 4 2 10 9 1 11 13 10 9 1 10 9 1 9 15 15 9 13 1 9 2
7 1 10 9 13 15 3 2
40 10 9 1 9 8 2 11 2 8 2 13 16 10 0 9 2 0 15 0 4 15 0 9 1 4 2 2 3 1 15 9 10 9 3 12 9 13 4 4 2
19 10 9 13 15 9 2 1 10 9 7 0 9 2 1 10 0 0 9 2
34 1 10 0 9 2 11 2 13 3 3 8 1 10 9 1 11 12 9 1 9 4 9 2 12 1 9 2 15 12 9 3 13 4 2
18 15 1 15 13 3 3 1 10 0 9 2 7 4 3 1 9 4 2
8 10 9 13 13 3 0 4 2
19 7 16 10 9 15 9 3 13 2 13 15 1 12 9 3 10 0 9 2
11 10 9 13 10 9 1 10 0 9 4 2
12 10 9 15 3 3 1 9 13 4 1 4 2
21 10 9 1 15 9 4 3 4 1 10 0 0 9 1 8 2 11 2 1 11 2
14 10 9 1 10 0 9 1 10 0 9 4 13 0 2
16 15 0 9 13 2 1 9 1 15 10 2 15 13 9 4 2
18 7 8 12 0 0 13 1 15 9 1 11 1 15 9 1 4 4 2
15 9 13 3 10 9 8 4 16 9 15 15 13 0 13 2
10 10 0 9 13 15 13 1 9 4 2
21 11 2 12 2 7 11 2 12 2 1 11 13 3 15 9 3 1 10 0 9 2
29 10 0 9 4 4 1 10 9 1 15 8 2 10 9 1 9 7 9 1 10 9 2 8 9 1 15 0 8 2
27 2 15 13 10 0 9 1 11 3 3 10 9 4 2 1 15 9 1 9 10 0 9 2 2 13 11 2
21 2 12 9 3 13 15 1 11 1 8 3 1 4 2 16 10 9 8 1 13 2
15 3 13 15 0 1 10 9 2 16 0 9 1 13 2 2
30 8 2 10 9 1 15 13 1 10 9 1 12 1 8 2 4 0 10 9 3 4 4 1 10 9 1 9 7 9 2
20 1 11 2 1 2 8 2 9 2 4 1 15 9 11 3 3 15 1 4 2
11 7 15 3 1 0 9 1 10 9 15 2
48 16 10 0 9 3 3 10 9 13 7 10 0 9 1 10 11 0 13 1 10 15 3 3 0 9 1 12 9 2 4 10 9 1 15 8 3 0 1 10 9 15 15 1 10 9 4 13 2
40 3 4 11 2 12 2 1 11 2 15 8 15 8 1 8 13 3 1 4 2 3 0 16 10 9 3 10 0 2 13 9 4 16 15 0 3 10 9 4 2
12 2 10 10 9 13 15 3 4 1 15 9 2
9 15 4 15 0 9 1 10 9 2
9 15 13 15 3 0 13 1 15 2
8 15 13 3 3 15 3 3 2
10 10 0 9 1 10 9 4 3 3 2
20 1 15 1 15 9 3 1 13 2 13 15 10 9 0 3 1 10 9 2 2
8 7 9 4 3 8 1 11 2
34 10 9 1 10 9 13 3 3 15 16 2 9 2 2 7 13 0 2 9 2 7 10 13 9 1 10 0 9 13 15 9 0 4 2
19 16 11 10 0 9 4 4 2 4 1 11 3 3 2 3 13 2 4 2
12 2 15 13 0 16 11 3 15 1 9 4 2
23 9 1 11 13 3 0 3 2 0 16 15 3 3 4 16 15 13 1 15 15 9 2 2
8 3 13 9 11 15 0 4 2
36 1 8 2 8 1 11 9 2 8 2 2 13 15 1 15 9 10 0 9 7 9 7 13 15 3 1 3 15 3 3 1 4 1 15 9 2
13 2 10 0 9 13 0 0 1 4 1 10 9 2
7 3 3 3 2 7 0 2
14 15 13 10 9 4 1 9 16 15 7 15 13 2 2
14 10 9 2 15 12 2 13 10 9 1 10 0 9 2
8 3 13 11 1 3 10 9 2
13 2 0 16 15 0 13 2 13 15 0 4 2 2
15 11 10 9 3 13 8 10 9 10 9 1 15 0 3 2
28 1 9 3 5 10 9 1 15 13 9 13 3 9 1 15 5 13 15 1 9 9 4 2 13 1 10 9 2
36 12 9 3 4 10 13 9 1 10 11 15 2 16 13 16 10 9 0 9 13 4 1 11 2 13 12 9 1 10 0 9 4 16 15 9 2
15 10 9 4 15 0 2 15 9 15 13 4 7 15 4 2
12 7 16 10 10 9 13 10 9 3 3 3 2
28 15 3 13 2 4 10 9 2 0 2 9 2 2 10 9 16 10 0 9 9 13 1 10 9 1 10 9 2
41 15 4 1 15 15 10 13 9 13 16 10 9 1 13 1 9 2 9 2 0 9 1 10 9 7 3 3 15 8 2 1 10 0 9 1 15 15 10 9 13 2
10 3 13 15 4 16 10 13 9 4 2
35 10 9 1 0 9 8 1 10 0 9 11 1 11 4 9 2 13 15 8 10 9 4 7 10 9 3 0 4 1 4 1 15 13 9 2
10 10 9 3 4 0 2 1 10 9 2
14 1 12 13 10 0 9 16 10 9 15 0 9 4 2
28 7 1 10 9 16 10 9 12 9 8 4 4 16 1 13 9 1 4 2 13 10 9 1 12 3 0 3 2
15 10 9 3 13 10 0 9 1 9 15 1 10 9 4 2
11 3 15 9 13 16 9 1 9 4 4 2
12 10 9 1 0 9 13 10 15 9 4 4 2
19 15 13 8 4 3 10 9 4 2 7 13 15 3 3 4 16 15 4 2
8 15 13 1 11 7 10 11 2
21 3 10 9 1 10 0 0 9 13 1 10 9 1 15 15 9 10 9 0 4 2
15 8 2 15 9 11 7 15 9 8 13 8 10 9 4 2
12 7 10 9 3 4 3 0 0 2 13 15 2
7 2 15 13 15 3 4 2
12 15 4 0 2 10 0 9 2 2 13 11 2
13 15 1 9 3 13 4 10 0 9 2 13 15 2
16 15 13 0 4 1 15 9 2 0 10 9 1 11 4 4 2
53 3 13 8 1 15 9 1 0 0 9 3 9 1 4 1 1 10 11 1 11 15 2 8 2 13 2 10 0 9 1 9 1 10 0 9 8 10 9 1 10 9 2 8 2 7 2 15 13 1 10 9 2 2
36 3 10 0 9 1 11 13 3 2 2 15 13 4 15 3 1 15 9 4 4 2 7 1 9 13 15 15 3 3 4 2 2 13 10 9 2
44 10 9 4 3 1 11 7 8 4 2 7 10 9 1 11 4 15 9 10 0 2 16 9 8 2 9 2 3 0 13 15 9 10 9 8 4 4 1 15 13 1 15 8 2
8 15 4 10 0 0 9 8 2
20 2 10 9 15 3 2 9 7 9 3 13 2 2 3 13 8 10 9 3 2
25 8 2 3 1 10 9 12 10 13 9 1 0 7 9 2 13 16 10 9 1 10 0 0 9 2
13 10 0 9 13 12 9 0 7 12 9 0 4 2
23 2 15 13 9 16 15 0 9 2 2 13 8 2 15 0 9 3 1 15 0 4 4 2
12 10 9 13 0 1 4 4 1 10 0 11 2
18 1 8 4 10 9 10 9 4 1 10 1 15 9 2 13 15 3 2
16 2 3 13 3 3 9 3 15 3 4 4 16 15 3 4 2
13 3 13 9 15 0 8 7 13 15 1 10 0 2
24 15 13 3 10 9 15 4 4 1 12 2 16 15 9 9 1 15 15 0 9 10 9 13 2
7 3 13 9 15 15 13 2
22 15 4 3 0 3 16 15 15 9 4 4 2 16 10 9 3 1 15 9 4 2 2
10 1 8 4 1 15 9 15 1 4 2
20 9 11 1 11 13 3 16 15 15 0 4 16 10 9 1 11 4 1 4 2
19 15 13 2 3 3 1 4 16 3 3 15 4 4 4 1 10 0 9 2
25 2 3 13 15 15 9 1 11 7 10 11 3 2 8 16 3 4 4 1 9 1 10 9 2 2
26 9 13 3 9 2 2 15 13 4 4 16 10 9 1 11 9 0 4 1 15 13 1 10 9 2 2
23 1 15 0 9 4 0 11 2 1 10 11 13 1 10 9 1 10 9 2 15 8 3 2
14 2 9 13 10 0 9 4 4 16 15 3 4 4 2
21 3 13 15 1 11 15 13 15 10 9 4 4 2 3 11 1 15 9 4 4 2
9 16 9 8 15 13 4 1 11 2
21 15 13 0 2 16 15 15 3 13 4 2 4 3 3 7 9 1 15 4 2 2
19 10 15 13 9 11 13 10 9 1 15 15 12 9 1 10 0 0 9 2
6 15 13 8 1 11 2
10 10 9 13 15 1 9 1 10 9 2
11 10 9 1 11 13 15 1 10 0 9 2
11 3 0 4 0 16 9 8 0 3 13 2
18 10 9 13 16 11 3 4 2 7 13 0 3 4 1 10 9 3 2
12 1 9 4 4 16 15 1 10 9 4 4 2
17 3 13 9 4 1 10 9 15 10 0 9 1 10 9 13 4 2
18 0 9 13 3 3 3 9 1 10 9 7 13 10 9 1 9 9 2
7 15 13 1 10 0 9 2
15 10 12 9 13 4 4 1 15 2 11 2 8 0 9 2
18 0 0 9 4 3 10 0 9 1 10 11 2 7 3 10 3 0 2
26 11 7 8 4 10 3 0 9 1 11 2 7 15 13 1 10 5 3 13 5 9 1 10 9 4 2
12 1 11 13 1 12 10 0 13 9 15 9 2
21 3 4 11 3 0 9 7 13 1 13 3 16 10 13 9 8 15 13 13 4 2
9 9 12 13 15 12 9 4 4 2
17 0 11 2 16 12 0 9 13 4 4 2 13 10 0 9 4 2
23 12 9 0 4 10 0 9 2 15 15 13 9 1 10 0 9 2 3 0 3 1 4 2
17 9 13 16 3 15 15 1 4 4 16 1 10 2 0 2 11 2
12 3 13 3 15 9 4 1 10 13 0 9 2
28 9 7 9 13 16 3 10 9 3 4 4 7 16 15 3 13 9 3 1 9 4 4 2 15 10 9 13 2
25 1 10 9 1 10 9 11 13 10 9 1 10 0 9 1 9 9 15 16 1 10 9 0 9 2
20 15 16 10 9 3 3 13 16 10 11 0 9 10 9 1 12 9 4 4 2
22 15 9 4 0 0 16 1 15 9 10 9 1 10 9 1 12 12 9 3 1 13 2
14 3 15 0 3 13 4 10 0 9 11 1 9 4 2
7 9 8 13 15 9 0 2
24 1 10 9 11 4 3 4 1 10 0 9 3 10 9 2 0 2 0 7 0 2 13 4 2
14 9 8 13 16 10 13 9 13 7 13 9 3 4 2
8 15 13 11 1 10 9 8 2
24 15 13 16 3 9 4 4 1 10 9 1 10 9 8 2 3 15 13 2 8 2 9 4 2
14 2 15 9 13 1 15 10 9 16 15 3 13 4 2
24 15 13 10 0 9 4 1 15 9 7 15 9 4 1 10 0 0 9 4 2 2 13 11 2
16 10 11 13 3 1 10 0 9 1 9 2 1 10 9 8 2
10 15 13 3 4 16 9 0 4 4 2
19 10 9 4 0 4 1 10 9 15 2 3 0 0 0 9 2 13 4 2
17 10 9 3 1 13 9 13 1 3 3 8 3 2 13 11 3 2
14 2 3 13 15 3 1 10 0 9 13 1 15 3 2
8 0 2 16 15 3 0 13 2
15 15 13 15 1 3 3 3 15 4 7 15 13 0 2 2
13 3 13 9 4 15 0 9 1 12 9 13 4 2
15 8 1 11 13 15 1 15 13 16 10 9 10 9 4 2
7 2 15 13 15 3 4 2
12 15 13 1 9 1 10 9 4 15 0 9 2
17 15 4 0 16 11 15 3 3 4 2 2 13 15 1 10 9 2
14 10 9 13 16 10 9 1 10 9 3 3 4 4 2
11 9 1 9 1 9 7 9 4 0 0 2
15 2 1 15 9 13 3 3 3 15 4 2 2 3 8 2
13 9 11 1 9 4 1 10 9 1 15 9 4 2
24 0 9 13 15 1 10 9 1 15 8 16 10 9 3 2 3 0 9 2 10 9 4 4 2
21 15 4 3 4 16 10 11 1 10 0 9 3 0 4 4 4 8 10 0 9 2
25 3 13 10 9 1 10 9 3 0 1 10 9 15 1 10 9 1 10 11 7 10 9 4 4 2
15 1 15 9 13 16 12 9 1 10 9 1 9 13 4 2
23 16 15 15 16 12 9 1 3 13 13 10 11 1 10 9 1 10 9 1 10 9 4 2
8 7 10 9 13 3 3 4 2
13 1 10 0 9 13 12 9 1 10 9 1 9 2
12 11 13 16 15 1 10 0 9 3 0 4 2
33 1 10 9 1 8 1 10 9 1 15 9 13 3 10 0 9 1 10 11 3 13 4 4 1 10 13 9 1 9 11 7 11 2
13 10 9 9 13 0 9 3 1 10 9 0 9 2
37 3 13 10 0 9 8 2 15 1 10 9 13 9 2 3 3 16 15 1 10 9 4 4 2 15 1 10 0 9 1 10 0 7 8 4 4 2
32 8 2 1 3 1 10 0 9 15 3 0 13 1 10 9 2 13 1 4 16 15 13 3 1 10 9 1 10 11 4 4 2
24 2 15 13 15 1 15 3 2 15 13 3 3 3 4 2 2 13 15 2 13 1 10 9 2
25 1 10 0 9 2 1 10 9 3 9 11 10 9 0 9 13 4 2 4 3 0 15 9 4 2
18 10 9 13 3 3 3 1 4 4 1 10 13 9 15 3 4 4 2
31 10 9 13 15 3 1 4 1 10 9 1 12 9 2 3 3 16 15 1 10 0 9 13 2 3 13 11 11 15 13 2
14 2 15 9 3 1 10 9 2 2 13 15 9 0 2
16 11 1 15 0 9 13 10 15 9 11 1 4 1 10 9 2
17 10 9 4 3 2 16 15 3 13 2 4 4 1 4 13 4 2
17 10 11 13 3 1 10 9 1 10 9 4 16 15 3 3 4 2
31 15 13 15 1 10 9 4 2 7 9 4 15 3 4 16 10 9 9 10 11 0 0 13 4 4 2 7 15 13 3 2
26 0 16 10 9 10 9 1 15 8 13 4 2 13 10 9 0 1 10 9 7 11 9 4 7 9 2
17 9 11 13 10 9 1 10 9 16 10 13 9 15 3 4 4 2
33 16 9 11 15 9 4 2 4 10 9 2 3 1 10 9 2 2 3 11 1 10 9 1 9 1 9 1 11 7 11 7 11 2
36 15 9 4 15 0 3 3 2 11 7 11 13 15 0 16 15 9 4 2 3 16 15 1 15 9 0 4 16 10 9 1 10 9 9 4 2
13 11 9 0 1 9 2 9 11 4 3 3 9 2
19 9 13 3 0 1 10 9 15 11 13 2 9 10 11 2 9 1 11 2
18 15 4 2 0 9 9 11 10 11 2 9 8 2 9 8 2 4 2
18 10 9 1 11 13 3 10 9 11 2 7 15 4 15 9 1 11 2
13 15 9 4 0 1 10 2 0 9 7 9 2 2
12 15 13 3 3 15 4 7 15 4 3 11 2
31 16 10 9 3 13 3 15 9 3 1 4 16 11 1 10 0 9 12 9 1 11 4 4 2 13 1 15 9 9 4 2
17 9 7 11 13 15 3 16 10 9 11 0 0 1 9 4 4 2
9 4 15 10 0 9 1 10 9 2
11 15 4 2 13 10 9 2 8 15 4 2
31 1 10 11 4 3 15 9 0 4 2 10 0 9 13 4 7 4 4 10 9 1 15 1 1 11 1 9 1 4 4 2
16 1 11 4 15 1 9 9 16 10 9 3 15 0 4 4 2
11 3 15 4 1 11 4 2 10 9 4 2
22 11 13 15 4 1 9 2 3 10 11 2 15 3 3 9 13 3 5 0 5 9 2
11 8 10 9 1 9 13 3 1 15 3 2
11 11 4 9 1 4 1 10 9 1 9 2
15 1 10 0 9 13 15 9 9 1 9 1 15 15 9 2
32 3 13 3 1 11 12 0 7 0 9 3 9 1 10 10 9 9 13 1 10 9 2 9 2 9 2 9 2 11 7 11 2
9 9 4 1 15 9 10 0 9 2
23 0 13 9 13 15 3 3 2 3 10 11 2 7 15 13 15 0 16 15 15 8 13 2
9 15 4 3 0 2 7 3 0 2
24 10 9 4 3 0 2 3 3 10 16 12 7 12 9 2 2 10 9 1 9 4 3 0 2
25 10 11 13 3 3 1 13 16 15 3 15 15 4 2 7 13 3 9 3 16 10 9 1 4 2
8 15 13 1 15 13 1 9 2
28 15 13 13 2 7 16 10 9 4 4 13 15 16 10 9 15 13 1 9 1 15 15 9 15 0 4 4 2
22 15 13 10 0 9 8 3 0 3 16 15 9 10 13 12 9 9 4 1 15 8 2
30 15 13 15 3 2 7 4 4 16 15 11 4 4 16 1 15 9 0 9 3 1 13 7 1 12 13 9 1 13 2
17 11 4 1 10 0 9 11 10 0 9 4 7 10 0 9 13 2
16 10 0 9 16 10 9 1 10 0 9 1 10 9 1 13 2
23 10 9 11 13 1 10 0 9 1 15 9 3 12 9 4 16 10 9 1 11 1 13 2
25 1 9 11 13 15 3 1 15 9 1 0 9 8 7 9 1 9 8 10 9 1 10 9 4 2
16 3 13 0 9 1 11 2 11 7 11 13 4 1 10 9 2
13 11 13 8 12 9 1 11 2 1 15 9 13 2
11 15 13 3 3 16 9 4 1 15 9 2
11 0 4 13 1 10 13 9 1 10 11 2
11 3 13 9 4 8 10 9 0 9 4 2
10 3 13 11 15 1 15 2 8 2 2
31 10 9 15 0 11 1 10 0 9 1 11 13 4 4 2 7 0 3 15 4 16 10 9 7 13 1 10 9 1 11 2
18 16 10 9 10 9 1 13 2 13 11 15 0 9 1 10 9 4 2
20 1 15 8 2 9 1 15 8 2 10 0 9 8 7 10 0 0 9 8 2
15 15 0 4 10 13 9 10 9 3 11 1 15 9 4 2
35 15 13 1 12 3 3 1 13 1 10 9 5 10 0 0 9 3 5 3 10 9 1 0 2 15 0 2 9 4 3 10 9 15 9 2
36 1 10 9 1 10 9 8 13 9 11 16 10 9 1 10 9 1 15 8 0 4 4 16 3 3 10 9 4 4 9 16 11 3 1 13 2
21 15 8 4 1 15 15 4 16 15 0 2 7 3 15 16 10 9 7 0 9 2
18 15 13 2 13 11 2 16 10 9 1 9 1 15 8 10 9 13 2
38 10 9 1 10 9 4 3 4 1 10 13 9 1 0 9 7 9 2 15 3 10 13 9 0 13 16 1 10 11 1 10 9 7 10 9 1 13 2
11 7 3 3 15 4 4 2 13 4 4 2
18 11 13 2 8 10 0 9 0 9 2 0 9 7 9 1 10 9 2
13 11 7 15 9 13 10 9 3 4 4 1 9 2
13 1 15 4 10 9 10 0 9 1 10 0 9 2
9 10 9 13 1 15 9 1 11 2
12 2 8 2 2 13 10 0 9 1 10 9 2
5 10 9 13 3 2
