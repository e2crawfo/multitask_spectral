786 17
8 9 1 9 0 1 9 13 9
51 9 12 2 12 2 8 8 2 2 13 9 9 9 9 0 0 1 9 0 1 9 13 12 9 1 9 9 2 9 9 9 2 1 9 9 1 9 9 9 0 0 15 13 1 15 1 15 13 9 9 2
51 7 13 9 9 0 13 7 9 9 2 9 1 9 2 13 12 9 1 15 12 9 2 9 7 9 15 8 8 13 1 9 8 8 7 9 0 14 13 0 1 9 15 13 9 8 1 9 7 9 0 2
29 7 13 8 1 7 9 15 13 0 9 9 1 9 9 9 0 8 8 13 1 9 2 9 0 2 1 9 0 2
13 7 13 2 14 13 1 9 15 1 9 9 2 2
37 7 13 8 0 1 9 12 9 2 13 9 1 9 7 9 9 0 7 13 7 13 8 0 1 15 15 13 1 7 15 9 0 1 9 9 2 2
38 7 13 9 2 9 1 9 2 15 13 15 9 1 12 9 1 9 1 9 1 9 15 9 0 1 10 9 1 9 15 9 1 12 9 2 9 12 2
14 7 13 9 0 1 9 0 1 9 0 1 9 0 2
3 1 9 9
53 8 12 2 12 2 8 8 2 2 1 15 13 9 9 0 1 9 9 2 8 2 8 8 2 8 2 13 9 9 9 8 1 9 15 9 0 1 9 15 15 13 9 9 0 1 9 0 1 9 10 9 0 2
48 1 9 12 8 8 8 2 9 2 8 8 8 2 8 2 13 9 1 9 8 0 1 9 9 0 1 10 9 0 0 1 9 9 7 8 1 9 9 7 1 0 9 9 0 0 1 15 2
4 9 1 9 0
32 8 12 2 12 2 8 8 8 2 2 12 13 8 8 0 9 15 1 9 9 9 8 8 8 8 8 8 2 12 9 2 2
33 7 13 9 8 0 8 0 7 8 8 8 8 8 0 13 1 9 15 1 9 8 15 13 8 9 9 15 1 1 12 12 9 2
37 12 13 8 8 9 9 9 8 7 9 8 8 0 15 13 1 9 0 9 13 1 9 15 1 8 0 1 9 12 9 1 1 7 13 9 9 2
40 7 13 8 2 12 9 2 9 9 9 9 15 1 9 9 0 0 2 7 15 13 12 9 3 1 9 12 15 13 15 8 1 9 7 15 13 1 9 0 2
17 12 13 0 8 8 9 8 0 9 1 9 9 1 9 8 0 2
16 7 13 9 9 8 2 12 9 2 1 12 2 12 12 9 2
24 7 13 8 12 9 0 1 9 9 15 7 13 1 9 8 8 8 0 1 9 15 1 8 2
12 12 9 7 9 9 1 9 0 1 9 9 9
46 8 12 2 12 2 8 8 2 2 13 1 9 0 0 7 9 0 1 9 12 9 1 9 8 13 9 9 9 9 8 1 9 9 7 13 1 12 9 1 0 7 13 1 9 9 2
29 7 13 9 1 9 12 1 9 0 2 12 8 2 1 10 9 15 13 1 9 12 8 9 8 7 13 12 9 2
32 7 14 13 10 9 10 9 1 9 8 7 9 0 7 13 1 9 0 9 0 0 13 1 0 1 9 2 9 1 9 9 2
13 9 9 9 0 1 9 13 9 1 9 9 2 9
40 9 12 2 12 2 8 8 8 2 2 13 9 9 9 0 1 9 8 8 9 1 9 9 2 9 1 9 9 1 0 9 0 7 13 9 1 9 9 0 2
43 7 13 9 1 9 9 9 0 1 9 0 1 9 8 8 1 9 8 8 7 2 9 9 14 13 1 7 15 13 7 15 1 0 7 13 1 12 7 9 9 0 2 2
33 7 13 8 13 1 9 2 9 12 9 1 9 9 7 13 9 1 9 9 9 9 1 9 0 1 9 9 2 9 1 9 2 2
39 7 13 9 15 13 1 9 0 1 9 9 12 9 9 15 1 9 9 0 1 9 10 9 15 13 9 12 9 7 15 13 1 9 2 9 9 15 0 2
9 9 9 0 1 9 0 1 9 9
46 8 2 9 8 2 12 2 12 2 8 8 2 2 8 12 9 0 9 9 9 9 0 1 12 9 1 9 8 1 9 9 1 9 9 7 9 1 9 7 13 9 9 15 13 9 2
44 7 13 9 1 9 9 0 0 1 9 8 8 2 7 9 9 12 0 1 9 9 9 9 0 7 13 9 9 15 1 12 1 12 9 2 13 9 15 1 12 7 12 9 2
32 7 13 9 15 13 1 9 9 9 1 9 8 2 9 9 8 2 2 8 9 0 9 15 13 1 0 0 7 9 0 2 2
38 7 13 7 15 2 13 9 9 9 1 9 9 9 8 7 9 9 15 7 9 9 9 1 15 7 9 1 1 9 0 7 9 1 1 9 0 2 2
49 7 13 2 7 9 1 9 0 14 13 1 9 0 7 9 1 9 7 9 1 1 9 0 7 1 9 7 9 1 9 9 9 7 9 9 12 9 14 13 1 9 0 9 7 1 0 9 2 2
35 7 13 10 9 1 9 9 0 1 9 0 9 14 13 1 9 9 0 0 1 8 8 7 9 9 9 9 0 0 1 12 9 2 9 2
7 9 0 1 8 7 9 8
50 8 12 2 12 2 8 8 2 2 13 9 2 8 2 9 9 9 1 9 0 7 9 0 8 8 13 3 1 9 0 9 8 8 2 12 9 2 9 1 9 2 7 13 15 1 9 15 0 0 2
33 7 13 9 7 8 15 13 9 8 1 9 9 9 0 13 0 9 13 9 0 1 9 2 9 0 2 1 9 0 0 8 8 2
26 7 13 8 9 3 9 0 1 9 8 1 9 9 8 1 9 9 8 7 9 15 7 9 9 15 2
30 7 13 8 8 13 15 9 9 9 8 8 8 9 1 9 1 9 9 8 0 7 0 1 9 8 1 9 9 15 2
35 7 1 0 7 13 8 1 9 15 9 9 1 9 1 9 9 15 1 8 2 12 8 9 9 2 7 14 13 0 7 13 1 9 0 2
36 7 13 8 1 12 9 2 9 0 1 8 1 9 1 9 13 1 9 12 9 1 9 0 1 9 1 9 9 0 1 8 0 1 9 8 2
45 7 13 8 13 1 9 1 12 9 0 2 9 0 1 9 8 1 9 9 15 13 13 15 1 9 15 15 13 9 1 12 9 0 1 9 15 9 1 9 9 0 1 9 0 2
6 9 0 1 9 9 0
36 8 12 2 12 2 8 8 2 2 13 9 0 9 9 7 9 8 8 14 13 9 0 1 9 1 9 9 13 15 3 1 8 0 7 8 2
21 7 13 9 7 9 1 0 7 9 15 14 13 9 2 14 13 8 9 9 9 2
55 7 14 13 1 9 9 14 7 15 13 7 13 9 0 9 1 9 9 12 2 9 0 0 12 7 8 2 0 9 15 1 12 1 12 9 2 9 1 8 2 9 2 7 14 13 1 9 0 1 9 0 1 9 15 2
21 7 14 13 8 3 9 15 9 1 9 9 8 0 2 0 1 12 12 9 2 2
25 7 1 0 7 13 9 0 1 9 15 1 9 9 0 1 9 15 1 9 1 8 0 7 8 2
11 9 9 7 9 0 1 9 1 9 1 8
39 8 12 2 12 2 8 8 2 2 13 9 1 9 0 0 1 9 0 7 9 13 7 13 9 0 1 9 0 3 9 1 9 13 1 9 0 1 8 2
31 7 13 9 7 8 8 2 12 9 2 13 15 9 0 9 9 9 1 9 15 1 9 8 1 9 8 2 9 9 2 2
41 7 13 8 8 2 12 9 2 9 9 9 1 8 9 8 2 9 9 2 0 1 9 15 15 13 12 5 1 9 15 1 9 13 9 1 9 8 2 9 2 2
27 7 13 9 0 2 8 8 2 12 9 2 13 3 9 9 1 8 8 3 1 9 15 9 1 9 0 2
17 7 13 12 9 14 13 0 3 9 1 9 0 7 9 0 9 2
26 7 13 8 8 2 9 9 0 2 7 9 13 1 9 15 7 7 1 9 0 7 13 9 0 2 2
26 7 13 12 9 1 9 9 7 12 9 7 12 9 1 9 0 8 1 3 9 1 9 9 1 9 2
14 9 5 8 5 0 1 9 13 9 9 15 1 9 0
41 8 12 2 12 2 8 8 2 2 13 8 8 9 9 9 5 8 5 1 9 9 3 9 7 9 13 9 1 9 7 8 7 13 1 9 9 15 1 9 0 2
56 7 13 9 9 8 1 8 9 15 7 9 14 13 1 9 0 9 1 9 1 9 9 15 1 9 8 2 12 2 7 13 2 8 13 9 0 1 8 8 2 2 7 15 13 2 7 9 14 13 0 9 1 9 0 2 2
32 7 13 8 1 7 9 0 1 8 0 7 0 15 13 9 15 0 1 9 0 0 2 13 7 13 1 9 7 13 9 9 2
44 7 13 9 5 8 5 3 9 1 8 1 9 9 15 0 1 9 8 2 12 8 2 8 2 8 0 1 0 9 0 7 0 1 9 0 1 0 7 1 9 9 0 0 2
54 7 13 8 7 9 1 9 1 9 9 0 0 0 2 7 9 0 13 9 15 8 2 12 1 9 0 9 7 7 8 13 1 9 9 15 9 2 8 2 2 7 0 9 13 0 1 9 1 0 1 9 8 0 2
37 7 13 9 1 9 15 9 9 9 0 2 8 8 2 7 14 13 9 8 2 12 0 15 13 1 9 9 10 2 7 14 13 9 9 12 9 2
8 9 9 2 9 0 2 2 2
81 9 2 7 13 9 9 9 9 0 1 9 9 1 8 8 15 13 1 9 9 9 9 15 1 9 7 9 7 15 13 7 15 14 13 1 9 9 9 9 15 14 13 9 1 9 7 15 9 9 0 1 9 15 13 1 15 7 13 9 0 1 9 1 9 0 1 9 9 15 1 9 9 7 1 15 8 8 8 8 8 2
58 7 13 3 9 9 0 8 8 15 13 1 9 12 12 9 0 2 12 12 9 2 1 9 0 7 1 9 1 9 9 9 0 0 9 15 13 15 9 9 1 9 15 1 9 9 9 15 0 7 9 0 1 9 9 15 1 9 2
74 7 13 8 9 1 9 9 0 1 12 12 9 7 1 9 15 9 1 15 1 9 1 9 9 1 9 8 8 15 13 8 1 12 9 0 1 9 1 9 15 7 13 0 1 9 9 1 9 9 12 9 9 9 1 15 2 7 13 8 7 15 14 13 7 14 13 8 9 15 15 13 9 15 2
62 7 13 8 13 1 9 9 7 9 0 1 9 1 9 9 1 9 15 1 9 15 7 8 9 15 8 8 8 1 7 9 0 7 9 9 2 7 13 0 1 8 1 9 9 15 9 1 9 9 0 2 8 2 9 1 9 15 13 1 15 9 2
74 7 13 9 8 8 1 9 15 8 8 1 9 7 9 9 1 9 8 8 8 1 9 9 9 9 0 7 13 9 9 2 7 1 9 9 0 1 9 8 9 15 12 9 2 7 7 15 14 13 9 7 13 8 1 9 9 0 1 15 9 1 9 7 13 1 15 9 15 9 15 13 15 8 2
17 7 13 8 13 1 9 0 0 1 8 1 9 9 15 1 9 2
31 7 14 13 13 9 9 8 1 15 9 7 13 9 1 9 15 7 13 9 1 9 9 1 15 0 7 0 0 1 9 2
76 7 0 7 9 8 13 9 8 1 9 1 9 15 9 9 9 1 9 9 9 1 8 11 9 0 8 13 1 9 15 7 13 15 1 0 7 13 9 1 9 15 9 0 7 9 0 7 13 12 9 1 9 9 9 2 7 13 1 9 14 12 1 9 9 9 7 9 9 8 1 9 0 1 9 15 2
52 7 1 9 0 3 2 13 8 9 9 13 1 9 9 9 9 9 9 15 1 9 9 15 13 1 9 1 9 1 0 9 8 8 0 1 9 0 1 9 9 8 2 7 9 9 0 9 1 9 9 3 2
31 7 13 9 9 8 0 1 9 1 9 0 15 13 1 9 1 9 15 7 13 9 15 9 15 1 9 15 9 9 15 2
7 8 8 13 9 1 8 8
60 8 8 12 2 12 2 8 8 2 2 1 9 9 0 1 9 15 15 13 9 0 0 1 8 8 2 13 8 8 9 9 9 1 9 9 15 0 7 13 1 9 9 15 13 1 15 9 15 7 2 9 15 2 0 1 9 0 8 8 2
45 7 13 8 8 1 9 12 9 0 15 13 1 15 9 0 2 1 12 9 1 8 8 8 8 8 8 7 9 0 2 7 9 8 3 1 9 8 8 0 9 1 9 0 2 2
48 7 13 8 15 13 1 15 0 9 1 15 1 9 1 9 0 1 9 2 14 15 3 1 9 9 7 13 1 15 9 2 2 7 13 8 1 9 0 9 0 1 12 9 0 2 9 0 2
18 7 1 9 13 9 15 8 1 9 7 13 15 1 9 15 1 15 2
33 7 13 9 8 2 9 1 9 15 7 1 9 15 1 9 0 7 0 2 9 1 9 8 8 1 10 9 15 13 8 9 2 2
35 7 1 9 15 13 9 1 9 7 9 13 1 9 8 8 9 1 8 8 7 13 9 2 7 13 12 1 12 12 9 0 1 9 9 2
33 8 1 8 8 7 15 9 0 1 9 9 0 1 9 0 0 2 13 9 9 0 1 8 7 9 15 9 9 0 1 9 9 2
100 7 13 9 8 15 9 15 13 13 15 9 8 2 8 0 8 8 9 10 9 1 9 9 8 8 8 9 1 9 0 7 12 2 8 8 8 3 2 7 14 8 9 1 9 2 2 2 2 2 2 7 13 7 2 8 8 7 8 8 14 13 9 1 9 9 7 9 1 9 7 9 7 1 9 9 0 8 8 9 15 2 0 1 8 8 0 1 9 1 9 0 15 14 13 9 0 1 15 9 2
47 7 13 8 9 0 1 8 8 9 2 0 2 2 7 13 7 2 8 8 13 0 1 0 9 0 8 8 1 8 8 0 2 9 7 15 7 9 0 13 7 13 1 9 9 0 2 2
30 7 13 9 0 1 7 15 2 1 8 9 2 2 2 2 2 13 0 0 2 8 8 8 9 7 15 9 0 2 2
26 7 1 9 9 0 2 8 12 2 8 13 0 1 9 9 13 1 15 2 9 0 1 9 8 2 2
28 7 14 13 8 2 12 9 2 1 8 8 9 7 13 1 8 1 9 9 15 0 7 13 9 9 1 9 2
13 7 13 1 15 1 9 15 2 13 9 0 2 2
30 7 13 8 8 8 9 9 1 7 13 9 1 9 1 9 0 1 8 1 8 2 9 2 1 9 9 7 9 0 2
40 7 13 9 0 9 15 9 1 7 13 9 1 9 15 0 8 8 9 1 9 0 15 14 13 1 15 1 9 0 8 8 1 0 1 9 0 2 9 0 2
28 7 13 9 8 9 8 9 8 1 9 15 2 8 8 13 9 1 9 9 7 13 1 9 9 8 8 2 2
38 7 13 12 9 7 12 12 9 7 12 1 9 9 9 1 8 8 1 9 1 9 0 15 13 9 0 1 9 0 1 9 0 1 9 0 2 9 2
14 7 13 1 0 7 13 9 15 0 1 9 1 8 2
10 9 9 9 1 9 12 8 1 9 9
39 8 12 2 12 2 8 8 2 2 8 2 9 2 13 9 9 0 8 8 7 9 0 13 9 9 9 12 9 0 1 9 0 0 8 1 9 9 8 2
28 7 13 9 9 9 9 13 1 9 1 9 9 9 2 7 13 9 9 9 9 9 1 9 9 1 9 9 2
35 7 13 9 9 9 0 9 8 8 13 9 7 9 9 2 14 13 0 1 9 2 7 9 0 7 9 13 0 1 9 1 9 9 2 2
55 9 2 9 2 13 9 9 0 1 9 8 8 9 9 9 8 8 1 9 1 9 2 7 15 1 9 0 1 9 13 1 9 0 2 7 13 8 0 1 9 9 9 2 14 14 13 3 1 9 0 1 9 0 2 2
31 7 13 8 1 7 2 9 0 1 9 1 0 0 1 15 1 9 7 9 7 15 14 13 9 0 7 9 0 0 2 2
49 9 2 9 2 13 9 9 0 8 8 9 7 9 7 9 2 0 2 1 9 1 9 9 2 7 13 8 1 9 1 9 0 0 2 14 15 0 1 9 7 0 7 13 1 0 9 13 2 2
40 7 13 9 15 13 13 1 9 9 1 8 15 13 15 0 2 7 9 13 1 9 9 9 7 9 3 2 1 15 13 7 15 15 9 0 1 9 9 2 2
28 9 2 9 2 9 2 13 8 9 7 9 0 9 8 8 9 8 8 1 9 9 9 9 0 1 9 0 2
38 7 13 8 1 9 1 9 8 8 2 8 8 8 1 10 9 1 12 9 8 8 8 8 9 0 1 9 9 1 9 0 1 9 1 9 9 2 2
43 9 2 9 2 9 2 13 9 15 13 9 0 0 9 1 9 2 7 14 13 9 1 9 9 0 8 8 9 9 1 9 7 15 13 7 13 1 15 1 9 7 0 2
25 7 13 9 15 13 15 9 9 0 8 8 9 1 0 9 7 9 1 9 1 9 9 8 8 2
48 9 2 9 2 13 9 9 0 8 8 9 7 13 9 7 9 1 9 9 13 1 15 9 0 1 9 1 15 2 7 13 9 0 0 7 8 13 7 13 10 9 2 1 9 9 0 2 2
23 7 13 7 9 14 13 1 9 9 0 7 13 1 9 0 0 1 9 9 0 1 9 2
26 7 14 13 12 9 0 1 15 9 7 9 13 13 1 9 1 9 0 9 1 9 1 9 1 9 2
18 8 2 9 2 13 9 9 9 9 8 11 8 8 8 9 1 9 2
60 7 13 9 0 0 8 8 7 9 0 8 8 13 1 9 0 15 7 13 1 15 9 8 1 9 9 13 15 9 9 0 7 0 7 1 1 15 1 9 0 9 9 8 8 8 8 8 8 7 9 9 8 8 8 7 9 9 8 8 2
56 9 2 9 2 0 2 13 9 9 9 1 9 8 8 9 9 7 9 0 1 9 9 1 9 1 9 9 2 7 13 8 1 9 0 1 9 2 1 0 9 1 9 9 9 1 9 9 0 7 9 0 13 1 9 2 2
28 2 13 9 1 9 1 9 0 1 9 0 0 15 13 9 0 1 9 9 7 13 1 9 9 7 12 9 2
40 9 2 9 2 13 9 0 0 9 1 9 1 9 0 8 8 1 9 9 0 9 15 13 15 1 9 7 9 0 8 8 1 9 1 9 9 0 1 9 2
37 9 2 9 2 13 9 9 7 12 9 13 9 1 9 1 9 9 0 0 1 9 8 2 12 9 9 9 2 7 8 2 12 9 1 9 2 2
26 9 2 9 2 13 9 9 9 8 8 8 2 9 9 9 8 8 9 1 9 0 1 9 9 0 2
29 7 13 8 1 9 9 9 2 0 8 2 0 7 9 9 0 15 13 1 15 7 13 9 9 9 1 9 12 2
34 7 9 8 13 0 7 9 9 13 13 7 13 8 8 8 9 9 9 1 10 9 7 15 8 13 9 9 9 1 9 0 1 9 2
14 7 14 13 8 8 9 1 9 9 7 9 1 9 2
31 8 2 9 2 9 2 13 12 9 9 15 1 9 9 9 1 9 9 8 9 7 13 13 9 1 15 1 9 9 0 2
51 8 2 9 2 13 9 9 9 9 7 9 0 8 1 9 15 1 9 7 9 1 9 12 9 1 9 8 0 13 9 1 1 9 12 2 12 8 8 1 9 8 9 9 8 8 13 9 15 1 15 2
11 7 14 13 9 1 9 7 9 1 9 2
36 8 2 8 2 9 2 0 2 13 9 8 8 8 8 9 7 15 13 9 9 0 0 8 8 3 2 1 7 13 9 0 8 8 9 9 2
36 2 13 9 9 0 7 9 0 8 8 13 8 9 1 9 9 9 1 8 1 9 9 2 7 14 13 8 1 9 9 15 0 8 8 8 2
45 8 2 8 2 9 2 1 0 1 12 9 1 9 1 9 9 1 9 8 0 2 14 13 9 9 8 15 13 9 15 9 3 14 1 9 0 9 14 13 1 9 9 9 0 2
37 8 2 9 8 2 0 2 8 2 0 2 13 9 8 0 8 8 8 9 1 9 9 1 9 9 1 0 1 9 1 9 1 9 0 1 15 2
32 7 13 8 1 9 13 15 1 9 9 0 7 12 1 9 1 9 0 1 9 9 1 12 9 1 9 0 1 9 9 0 2
47 2 7 14 13 9 9 8 9 9 0 1 9 9 9 0 7 13 9 0 1 9 0 0 1 9 8 9 7 13 0 9 0 0 13 1 8 0 1 9 0 15 13 1 12 1 12 2
41 9 2 9 2 9 2 13 9 1 9 9 7 9 9 9 7 9 13 1 9 0 1 9 9 9 2 15 13 12 9 7 12 9 7 15 9 9 1 9 0 2
58 9 2 0 2 9 2 9 2 1 9 9 0 1 9 15 15 13 9 0 0 1 8 8 2 13 8 8 9 9 9 1 9 9 15 0 7 13 1 9 9 15 13 1 15 9 15 7 2 9 15 2 0 1 9 0 8 8 2
44 7 13 8 1 12 9 0 2 1 12 9 1 8 8 13 8 8 2 8 7 9 0 2 7 9 15 3 7 13 9 0 1 9 0 2 8 8 2 9 0 1 9 0 2
33 8 2 8 2 13 9 0 0 2 8 8 2 9 7 15 14 13 9 9 9 8 9 2 7 15 9 1 9 1 9 9 0 2
8 9 8 2 9 8 13 1 9
65 8 2 8 2 12 2 12 2 8 8 8 2 2 13 9 9 9 0 0 1 9 9 0 2 12 2 12 8 2 0 8 8 1 9 1 9 0 1 0 1 9 2 1 9 7 13 1 9 0 1 9 8 0 0 1 9 9 9 9 0 12 2 12 8 2
36 7 13 8 15 13 1 9 0 1 9 0 1 12 9 2 9 9 12 1 9 9 0 2 2 13 9 15 0 7 9 13 1 9 15 2 2
51 7 13 9 0 13 8 1 9 9 1 9 2 9 9 0 1 9 9 15 9 1 9 0 1 7 13 9 1 9 1 9 0 3 2 7 1 0 9 1 15 1 9 1 9 9 0 1 8 9 0 2
30 7 13 8 7 13 9 9 9 2 2 13 0 1 9 7 13 1 9 9 2 7 14 13 13 9 1 9 15 2 2
26 7 13 2 13 0 1 9 15 1 8 7 1 7 9 0 14 13 1 9 15 7 9 15 0 2 2
42 7 7 10 9 14 13 7 8 13 9 1 9 0 7 13 1 10 9 2 2 14 13 1 9 15 1 8 1 9 9 9 1 9 1 9 9 15 13 9 15 2 2
39 7 13 8 1 7 9 15 13 15 9 13 0 1 9 1 9 12 0 1 8 2 7 1 7 1 15 9 9 1 9 1 9 15 13 15 1 9 0 2
14 7 14 13 8 9 8 0 1 9 0 9 9 0 2
38 7 13 9 0 9 0 1 9 7 13 9 1 9 12 2 12 8 1 9 7 12 2 12 8 2 1 1 13 12 9 1 9 9 12 2 12 8 2
41 7 13 0 0 0 0 8 9 9 12 2 2 13 9 1 9 0 8 8 2 1 0 9 7 7 9 9 9 12 0 13 1 7 15 13 9 15 0 0 2 2
10 8 13 9 9 0 1 9 9 9 0
43 8 12 2 12 2 8 8 2 2 13 8 1 9 9 0 15 13 9 15 1 15 1 9 1 9 9 9 0 8 0 1 9 9 8 2 7 13 9 9 9 1 8 2
38 7 13 9 1 9 8 9 8 8 7 9 13 1 2 9 9 2 13 1 15 8 1 9 0 2 7 7 15 13 7 9 10 9 2 9 0 2 2
45 7 13 9 1 8 13 9 1 9 15 7 8 14 13 1 9 0 1 9 2 7 7 15 13 9 9 9 1 9 1 9 15 13 7 13 15 1 15 1 9 13 1 15 15 2
33 7 13 9 9 0 8 8 9 1 9 15 0 8 8 0 1 15 9 9 0 7 15 14 13 9 1 9 2 7 13 9 8 2
60 7 13 2 8 7 15 2 9 2 13 8 8 0 1 9 15 2 8 2 2 2 2 2 1 15 7 1 9 15 9 9 9 8 1 9 1 9 15 2 8 8 8 0 1 9 1 9 10 8 7 15 13 8 8 9 1 15 9 2 2
18 7 13 0 15 7 13 9 9 0 13 9 15 1 8 1 9 9 2
27 7 1 9 0 9 0 13 9 9 1 9 0 0 1 9 12 9 9 0 2 1 10 13 9 1 9 2
2 1 9
8 14 13 9 0 9 1 9 2
32 13 9 1 12 1 9 15 1 9 9 1 9 15 1 9 0 7 9 1 9 9 0 1 9 8 0 0 1 9 9 8 2
48 7 14 13 1 15 0 9 9 15 7 13 9 15 1 9 7 1 9 8 8 13 9 1 9 9 1 9 9 7 13 1 9 9 13 1 9 9 7 13 9 15 9 9 0 1 9 0 2
53 7 1 9 0 13 9 9 9 0 8 1 9 9 7 13 9 7 9 9 1 9 9 9 0 1 9 15 7 9 15 1 9 9 0 1 9 0 1 9 1 9 15 7 9 9 1 9 0 0 1 9 9 2
33 7 9 1 15 13 9 9 1 9 13 9 1 15 9 9 9 0 1 9 7 13 1 9 9 9 9 9 7 9 9 7 9 2
57 7 1 15 13 1 9 7 14 9 13 1 15 13 1 9 0 1 9 9 1 9 9 9 15 7 13 9 1 15 1 9 9 0 3 15 13 7 13 1 9 0 7 15 15 13 1 9 9 15 13 9 9 15 1 9 9 2
56 7 13 7 9 13 0 1 9 9 7 13 9 15 7 13 9 9 1 9 15 7 13 1 9 0 0 1 9 2 1 7 13 1 9 2 7 13 9 15 0 1 9 9 7 13 9 15 0 1 9 15 7 13 1 9 2
3 8 2 8
2 1 9
7 8 1 9 7 13 12 9
30 13 9 9 0 1 9 0 1 9 1 9 1 9 9 9 13 1 15 12 9 0 14 13 1 9 9 1 9 9 2
35 9 9 1 9 13 9 13 1 15 0 0 13 1 15 9 15 1 9 9 1 9 9 13 15 9 0 0 13 15 1 9 12 1 9 2
59 7 1 9 9 1 15 13 7 15 13 1 9 0 7 13 1 15 7 1 9 0 13 1 15 7 13 1 9 15 9 0 7 13 15 1 7 15 0 1 9 15 2 8 2 1 9 8 8 8 7 13 1 15 9 15 1 9 10 2
31 7 3 13 9 12 1 9 9 9 13 1 15 9 8 0 1 9 7 15 15 13 9 0 7 13 1 0 1 15 9 2
41 7 13 1 0 1 15 1 9 15 1 9 0 13 1 12 9 1 9 15 1 9 9 0 9 14 13 14 1 9 9 0 1 9 15 0 1 9 8 0 0 2
40 9 7 9 13 1 15 10 9 7 13 9 8 8 7 13 0 9 15 1 9 7 13 7 15 13 1 9 9 7 13 9 1 9 9 7 13 9 1 9 2
36 7 13 9 1 9 7 9 1 9 1 0 1 15 12 7 1 9 9 15 8 7 9 0 13 1 9 9 0 1 9 9 1 9 9 0 2
3 8 2 8
3 9 0 2
9 12 9 0 14 13 9 0 9 9
48 8 2 8 8 2 2 13 9 2 8 2 0 3 7 1 12 9 0 14 13 9 15 1 9 8 1 9 9 0 15 13 1 9 1 9 9 1 9 0 13 15 9 9 9 0 1 9 2
38 7 13 9 7 10 9 13 1 9 12 9 1 9 2 8 8 2 0 0 0 1 9 1 9 9 1 9 9 7 9 0 1 9 8 8 7 0 2
31 7 14 13 9 10 9 1 9 1 9 2 8 12 2 7 13 9 9 0 15 13 15 9 9 9 0 10 1 12 9 2
35 7 13 9 7 9 1 0 9 1 9 13 1 9 15 1 10 9 1 9 9 9 0 1 9 9 15 13 1 15 9 0 1 9 0 2
36 7 13 7 10 9 13 7 13 9 2 8 8 2 1 2 9 0 2 1 9 9 1 9 9 0 1 1 9 1 9 9 9 1 10 9 2
45 7 13 9 1 9 9 9 0 13 0 3 1 9 8 8 7 8 13 9 1 9 0 1 9 9 15 1 9 0 1 9 0 1 9 7 8 13 9 9 15 1 9 7 9 2
33 7 9 1 9 0 1 9 13 9 0 1 9 1 9 1 9 9 15 1 9 9 9 0 8 8 1 9 9 0 1 8 8 2
33 7 13 9 2 8 2 3 1 9 1 9 0 0 14 13 15 9 15 2 3 9 1 9 8 8 1 9 2 0 2 0 2 2
39 7 13 9 9 0 0 3 7 9 9 8 8 1 0 7 13 13 1 9 3 1 9 13 1 15 7 8 13 1 8 9 9 15 1 9 0 1 9 2
2 8 0
2 9 9
22 9 0 13 10 9 1 0 9 0 15 13 1 9 9 0 1 9 3 1 9 9 2
16 9 9 15 9 9 1 9 9 9 9 9 0 1 9 15 2
49 9 9 0 7 9 0 1 9 0 7 9 9 15 10 9 9 9 7 9 15 0 0 1 9 0 1 0 7 0 7 0 7 0 0 1 9 9 0 2 14 8 1 9 7 8 1 9 9 2
98 9 9 13 1 9 0 9 0 1 9 7 9 7 9 8 8 15 1 9 10 13 9 9 0 1 9 1 8 9 1 8 0 9 7 9 7 9 0 13 1 9 9 7 9 9 0 1 0 9 0 1 9 0 7 15 7 14 9 1 9 1 7 13 9 0 9 15 0 7 7 1 9 9 0 8 8 1 0 9 7 14 8 9 1 9 8 9 15 0 1 9 7 9 7 9 7 9 2
77 1 9 9 8 8 8 1 9 9 0 7 9 9 7 0 9 7 7 9 9 9 9 0 15 9 0 0 1 10 9 15 13 1 15 9 7 13 9 9 0 0 2 7 9 14 13 1 9 7 9 7 9 0 7 9 1 9 0 7 1 9 9 7 9 7 14 8 8 1 9 8 9 9 7 9 2 2
35 8 9 7 15 14 8 1 10 9 1 9 10 9 1 9 1 0 15 13 9 15 1 9 1 9 9 0 0 1 9 9 7 9 9 2
11 8 9 15 9 1 8 8 1 9 15 2
13 8 9 15 9 8 8 8 1 9 15 1 9 2
17 8 9 15 7 9 9 8 8 7 1 15 15 1 9 9 9 2
17 9 2 9 9 9 0 14 13 1 9 1 0 1 9 1 9 8
5 8 8 2 8 8
88 13 9 9 0 13 9 1 15 1 9 8 0 7 15 14 13 1 9 15 13 15 9 0 1 3 1 0 1 9 2 9 1 9 9 1 9 1 9 1 15 13 15 9 2 7 7 13 9 9 1 9 9 2 13 9 0 7 9 0 2 7 15 9 0 15 13 1 15 9 1 9 9 1 9 9 2 14 13 1 1 10 9 9 1 9 9 9 2
68 13 9 1 9 15 13 15 9 9 1 9 0 1 3 1 9 9 8 0 15 13 1 15 12 9 2 1 15 12 9 7 12 9 12 1 15 0 2 7 15 13 9 12 0 7 9 1 9 13 1 9 0 7 12 9 1 12 0 9 1 9 15 13 1 15 12 9 2
57 7 13 9 9 8 1 9 9 8 9 12 1 9 9 9 2 1 9 1 9 9 15 1 9 9 9 0 2 2 7 2 9 1 9 9 2 0 7 9 15 13 15 9 9 1 9 9 2 13 9 9 0 1 9 0 2 2
87 7 13 2 2 8 9 9 7 14 8 15 15 9 0 8 8 8 8 9 1 9 1 9 9 7 13 8 9 15 7 13 9 9 1 9 15 2 2 7 13 8 7 13 9 13 9 0 1 9 2 7 13 2 2 13 0 7 13 9 9 1 9 1 10 15 0 7 15 15 0 7 9 13 9 9 9 9 7 9 8 8 9 8 8 9 2 2
36 7 13 9 9 1 9 9 9 9 0 1 3 2 1 9 1 9 9 2 13 1 15 9 9 9 2 0 7 15 2 9 1 9 0 2 2
98 7 13 9 9 9 8 8 1 2 9 2 7 15 2 13 13 1 7 13 9 9 0 1 9 9 15 13 15 9 0 1 9 9 12 9 1 9 7 9 12 0 7 9 7 9 9 1 9 0 2 2 7 13 2 7 9 7 9 0 13 1 9 9 0 1 9 15 13 15 9 2 7 15 13 9 12 0 7 9 12 3 1 9 14 13 1 9 9 2 15 13 15 9 8 9 9 0 2
82 7 13 9 0 1 7 15 2 14 9 1 9 1 9 1 9 9 0 2 7 15 14 13 9 1 9 0 7 7 3 9 13 9 1 15 9 1 9 9 2 2 0 1 2 7 9 13 9 0 0 1 0 1 15 7 15 13 9 0 1 9 15 9 2 1 9 15 1 9 7 9 1 9 9 7 9 15 7 9 15 2 2
65 7 13 9 9 0 2 7 15 9 1 12 9 0 13 9 1 15 1 9 2 1 7 2 9 14 13 1 9 9 9 9 0 1 9 9 7 9 1 9 9 1 10 9 1 9 0 2 2 0 1 7 15 2 14 13 9 1 9 9 14 1 9 0 2 2
60 7 13 8 1 7 15 2 13 9 1 9 9 1 9 7 7 15 9 9 9 2 2 0 1 7 15 2 13 1 9 9 0 13 1 9 1 9 9 1 9 9 2 7 15 15 8 8 1 15 1 9 0 1 8 9 0 1 9 2 2
94 7 1 9 13 9 1 9 0 1 9 1 9 15 1 9 15 13 7 15 2 14 13 1 9 9 8 2 2 7 13 1 9 9 1 2 9 15 13 1 15 8 9 2 7 13 15 1 7 2 9 13 0 1 9 9 2 2 7 13 9 15 13 9 9 15 2 2 14 9 1 9 9 7 9 15 9 9 0 2 2 0 1 7 9 15 13 1 9 2 14 13 0 2 2
81 7 13 9 0 7 9 15 13 1 9 9 1 9 9 0 1 9 1 0 9 0 0 2 7 13 1 12 0 1 15 3 9 1 15 1 9 9 2 7 1 9 9 9 13 9 15 1 9 0 0 7 9 0 14 13 1 9 12 3 2 1 9 15 1 9 0 7 13 1 9 9 12 9 1 9 1 9 9 9 0 2
85 7 13 9 1 7 9 0 15 9 0 15 13 1 15 9 1 9 9 1 9 9 2 7 13 9 7 9 15 13 15 9 1 9 9 2 2 9 13 9 1 9 0 9 15 1 9 9 1 9 2 2 7 13 1 2 7 9 15 13 1 15 9 14 13 1 9 9 7 14 13 9 9 0 7 9 15 13 1 9 9 1 10 9 2 2
13 2 0 1 9 9 2 13 2 9 9 2 1 9
76 9 2 2 9 2 2 13 2 9 0 1 9 9 2 1 9 9 9 13 9 15 1 9 15 0 1 9 15 7 13 9 9 9 9 9 9 2 7 13 9 1 9 9 1 9 9 0 1 9 1 9 0 0 13 9 12 9 13 1 9 9 1 9 9 0 1 9 12 9 1 1 12 1 12 0 2
94 7 13 9 0 9 9 0 1 9 13 1 9 9 0 1 9 9 1 9 9 9 1 9 0 2 7 1 1 9 15 13 15 9 1 0 15 9 9 1 9 15 1 9 1 9 9 7 1 9 9 1 9 2 7 13 9 9 1 9 0 1 9 1 9 15 1 15 7 9 1 15 2 7 13 7 13 9 9 1 9 12 9 2 7 12 9 7 12 12 9 7 9 15 2
10 12 12 9 1 9 9 9 0 2 0
63 9 2 2 9 2 2 13 9 2 9 8 2 8 1 9 7 9 2 11 8 7 9 0 1 9 9 0 1 9 0 1 9 7 9 14 13 0 2 7 14 13 9 15 13 1 9 8 12 12 9 1 9 0 13 1 12 9 0 9 15 12 12 2
61 7 13 7 9 0 13 9 0 1 9 14 13 9 9 0 1 9 1 9 0 1 9 9 0 2 7 13 7 9 13 9 12 1 12 12 9 1 9 0 0 9 1 15 9 15 12 12 9 2 0 1 7 9 13 9 9 15 12 12 9 2
3 8 0 9
2 8 8
43 1 8 13 9 9 0 0 7 8 8 1 9 8 2 7 13 7 9 1 9 1 15 1 15 8 0 1 9 2 7 13 7 15 13 9 2 8 2 1 9 8 8 2
158 7 1 9 15 13 12 9 13 8 8 1 8 0 9 13 1 9 10 9 13 15 9 8 8 1 8 1 9 8 1 12 9 1 9 9 8 1 9 0 8 8 7 1 0 9 0 1 9 2 7 1 15 8 2 7 7 8 13 15 13 9 1 9 15 2 7 14 13 8 1 9 1 9 0 1 9 0 15 13 0 1 8 8 8 2 7 13 9 15 1 9 2 1 9 0 1 9 8 8 2 7 13 1 15 9 1 9 7 9 1 8 7 9 15 2 7 15 13 2 8 8 2 1 9 9 0 1 9 9 0 7 13 1 8 7 13 1 15 1 9 2 9 0 8 8 2 7 13 15 1 9 9 0 1 9 7 9 2
91 7 14 13 10 9 9 8 8 13 15 12 12 9 7 1 15 9 0 0 1 9 15 13 9 8 8 1 8 8 8 1 9 15 14 13 9 15 2 7 1 15 2 7 14 9 1 15 13 1 9 9 0 1 9 13 7 8 13 9 12 2 12 12 9 0 15 9 9 0 1 9 2 1 9 7 9 9 0 1 8 13 1 1 9 0 14 8 12 12 9 2
121 7 13 8 1 9 8 1 9 9 1 9 0 7 0 2 15 13 9 9 0 1 9 9 13 9 9 0 1 7 9 9 1 8 1 9 7 9 0 15 9 0 7 1 0 7 14 9 1 15 13 1 9 9 0 2 7 14 13 8 1 9 0 1 9 9 0 1 9 9 7 1 9 0 7 0 1 8 2 7 15 14 13 1 9 0 1 9 1 8 1 9 0 2 7 14 9 0 13 7 15 13 1 8 7 13 2 9 2 1 9 1 9 9 15 1 9 0 0 1 9 2
172 7 14 13 8 1 10 9 2 7 14 9 9 9 9 9 15 12 12 9 13 7 13 9 1 9 9 1 9 0 7 9 0 1 9 9 2 7 13 9 1 9 9 8 15 13 1 0 9 9 1 9 2 7 14 13 9 9 0 7 13 1 9 1 7 8 2 0 2 1 9 9 1 9 1 9 7 15 13 15 13 1 9 1 9 12 9 0 1 9 9 0 7 13 15 1 9 0 1 9 7 15 2 1 9 1 12 9 2 7 7 13 15 1 9 9 15 1 9 0 1 15 8 13 9 1 9 2 7 1 15 7 14 8 14 13 9 15 1 9 8 7 9 9 15 2 7 3 9 1 7 9 1 9 13 7 0 13 13 1 9 9 9 1 9 1 9 0 9 1 9 9 2
117 7 14 13 9 9 0 9 1 9 9 8 8 8 0 1 9 9 0 0 1 9 9 9 9 7 0 8 8 9 1 9 0 2 8 8 8 9 1 9 13 8 9 9 15 8 9 0 13 1 15 2 9 2 9 7 13 7 15 13 1 9 0 1 9 0 1 15 9 9 2 9 9 2 2 14 7 9 1 9 9 0 13 1 9 9 1 10 9 1 9 7 8 14 13 9 9 9 9 8 0 1 9 0 1 15 1 9 1 9 9 1 15 0 1 9 0 2
111 7 1 9 10 2 9 2 7 14 9 8 14 13 9 1 9 0 2 0 15 13 7 15 13 1 15 13 9 2 8 8 14 13 7 8 14 13 1 9 13 15 1 12 12 9 2 7 14 9 7 8 0 14 13 0 1 9 1 8 7 14 13 8 9 1 9 2 8 2 9 2 9 7 8 8 1 9 9 0 2 7 13 1 9 15 9 9 7 9 0 7 0 1 8 8 14 13 2 1 9 15 9 0 8 7 9 0 1 9 9 2
10 9 0 2 0 1 9 9 9 1 0
2 8 8
23 13 9 7 9 1 9 0 1 9 9 9 1 0 1 9 1 9 2 12 2 12 2 2
38 7 13 9 9 0 0 1 9 0 1 9 0 9 1 15 9 1 9 9 0 7 0 1 9 1 0 2 7 15 1 9 13 1 9 8 1 9 2
33 7 14 13 9 0 9 1 9 9 0 8 1 9 0 8 8 8 8 8 2 7 13 1 8 1 9 0 9 1 12 9 0 2
46 7 13 9 9 0 9 15 9 1 9 8 8 1 9 0 2 7 14 13 9 1 1 8 9 9 7 0 2 1 1 8 8 13 9 0 2 7 13 12 1 12 1 0 8 8 2
41 7 14 13 10 9 9 0 9 1 8 1 9 0 2 0 7 8 8 2 9 1 9 15 0 7 0 2 7 13 9 8 0 1 9 1 9 13 1 9 0 2
5 8 8 7 9 0
74 13 12 9 0 8 8 1 9 8 1 8 1 0 1 9 0 2 9 2 12 1 9 0 0 2 7 13 9 1 9 12 9 0 7 12 0 7 9 12 9 7 12 0 2 7 13 1 9 7 9 12 9 0 0 7 9 9 1 12 9 0 2 7 9 12 9 0 7 9 9 1 12 9 2
19 7 13 9 0 0 1 9 9 0 9 1 9 7 9 15 9 0 0 2
35 7 13 9 0 9 0 1 8 1 0 1 9 2 9 2 8 1 0 1 9 9 15 9 12 15 13 12 12 1 9 7 9 7 0 2
10 9 7 8 13 8 8 9 9 9 8
2 9 8
117 13 9 0 8 9 8 7 9 0 8 9 8 8 8 8 8 9 9 8 1 1 8 9 9 0 15 8 9 8 2 7 13 8 9 8 1 9 9 0 9 9 1 8 7 9 9 8 13 2 9 8 8 13 1 9 15 8 8 0 8 8 0 13 9 8 8 7 13 8 8 1 9 7 9 2 2 7 13 7 9 13 1 9 1 9 0 2 7 13 1 7 8 8 1 9 7 8 2 13 9 0 0 1 8 9 9 8 8 0 8 13 9 9 9 0 2 2
29 7 13 9 0 1 9 9 0 9 1 9 1 9 9 8 8 8 1 9 9 0 1 9 9 0 7 9 0 2
59 7 1 9 15 13 9 0 7 8 8 8 8 1 9 9 2 13 8 8 7 8 9 1 9 8 8 1 9 0 0 1 9 9 9 1 9 13 15 9 0 7 14 13 1 9 9 1 0 15 7 13 1 9 9 15 13 15 2 2
35 7 13 9 0 7 8 9 1 9 9 9 8 8 13 1 2 9 7 9 9 9 0 8 8 9 7 9 8 0 0 1 9 9 2 2
88 8 8 8 13 7 9 14 13 1 9 8 0 2 13 9 0 1 9 0 8 8 2 1 9 15 0 1 9 0 1 9 0 2 9 0 8 8 8 1 2 8 1 9 0 7 9 0 1 8 9 0 8 8 1 9 9 9 2 9 7 9 1 9 0 9 14 13 1 9 15 2 2 8 7 9 9 0 13 1 9 1 2 9 13 15 8 2 2
19 1 9 1 9 9 9 0 2 9 2 9 9 9 1 0 1 9 12 9
2 8 8
44 13 9 9 1 9 1 9 13 15 1 0 1 9 9 1 9 1 0 2 1 9 13 9 9 9 0 1 10 9 1 1 15 9 9 9 1 0 1 9 13 1 12 9 2
25 13 9 0 9 0 1 9 1 9 0 0 7 9 0 1 9 9 0 15 13 9 1 9 0 2
75 7 13 9 0 1 9 1 2 9 2 7 13 1 9 9 0 9 7 9 9 9 7 9 9 7 9 15 13 1 9 0 2 7 13 7 9 14 13 0 1 9 7 0 1 9 9 0 13 1 9 15 9 9 10 13 0 1 9 0 1 9 1 9 9 9 1 9 0 1 9 0 1 9 15 2
128 7 13 9 7 9 13 1 9 15 1 9 9 9 9 9 7 9 9 9 9 1 0 1 15 1 9 13 1 12 9 1 0 2 7 13 9 0 9 15 1 9 9 3 1 9 9 15 13 9 1 9 9 9 7 9 9 2 12 12 1 9 1 12 12 1 9 2 2 7 13 9 1 9 9 9 9 1 8 1 9 9 9 8 8 1 9 1 9 7 9 9 15 2 0 1 7 8 9 0 14 13 1 9 1 9 9 15 7 13 9 15 1 0 0 1 1 9 7 1 9 15 8 8 8 8 8 8 2
48 7 13 9 1 9 9 9 9 15 13 1 15 9 9 1 9 12 12 9 2 12 12 9 2 13 1 15 9 7 13 1 9 2 0 7 2 9 0 1 9 9 0 15 13 15 9 2 2
84 7 13 2 9 2 7 9 9 9 13 3 9 0 1 9 0 13 1 15 1 9 9 1 9 1 9 10 9 2 7 13 1 9 9 2 9 9 14 13 1 9 9 15 9 0 15 13 1 9 0 0 1 9 0 2 7 1 9 10 9 9 9 1 9 7 9 9 0 7 9 1 9 0 1 9 0 0 7 9 15 1 9 2 2
40 13 7 0 1 12 9 9 0 0 1 9 1 9 13 12 12 9 13 9 15 2 7 13 10 9 9 0 9 9 12 1 9 9 0 1 9 12 12 9 2
30 7 13 7 9 9 8 8 7 9 9 8 8 8 13 9 0 1 9 9 1 9 9 7 9 7 9 9 1 9 2
19 13 9 1 9 0 1 8 1 9 12 12 8 2 9 13 9 1 9 9
23 9 2 2 9 2 2 13 9 9 0 1 9 8 8 7 13 9 0 7 9 1 9 2
35 7 13 1 9 1 9 15 9 9 0 1 8 9 0 1 3 1 9 7 15 13 9 1 9 10 9 1 9 9 15 13 1 9 0 2
67 7 13 9 9 0 0 7 0 2 13 9 0 1 12 12 9 2 12 12 9 2 2 7 13 7 13 10 9 1 9 9 0 0 1 1 12 12 9 3 7 1 9 9 9 14 13 1 12 12 9 2 15 13 9 0 9 7 7 3 9 9 13 15 9 1 9 2
154 7 13 9 7 8 9 9 0 7 0 1 9 12 7 15 13 1 9 15 9 0 1 9 9 12 12 8 0 2 12 12 9 2 1 15 12 12 1 9 9 14 13 7 9 1 9 9 0 2 7 13 9 13 15 9 9 0 1 9 1 7 9 14 13 1 9 1 9 9 7 9 7 9 9 7 9 0 7 9 7 9 7 9 1 9 1 9 9 2 8 1 9 0 7 9 0 0 2 7 13 9 3 1 9 0 1 9 9 1 9 0 1 9 1 8 1 9 9 9 9 0 1 9 9 12 7 15 13 1 0 15 9 12 1 12 1 9 0 1 9 0 1 9 1 8 1 12 9 0 2 9 2 12 2
43 7 13 9 0 9 9 1 9 9 12 12 8 2 1 7 13 9 9 1 9 0 1 9 12 1 12 1 9 0 9 1 9 1 9 9 7 9 9 9 7 9 9 2
22 7 13 9 0 3 9 9 10 9 1 7 14 13 12 12 8 13 1 9 9 15 2
25 7 13 8 1 9 9 0 15 13 9 1 9 1 9 9 9 1 9 9 1 9 0 7 0 2
65 7 13 8 7 9 9 9 0 15 13 1 15 9 1 8 1 9 12 7 1 9 13 12 12 8 2 0 1 7 3 9 0 7 0 13 1 15 9 9 12 7 9 15 12 12 8 2 7 13 8 9 0 1 9 9 9 12 2 12 9 15 12 12 8 2
33 7 13 7 9 0 8 1 12 9 2 9 2 9 12 13 1 12 12 9 0 1 1 12 9 9 9 9 15 1 12 12 9 2
26 13 1 9 9 0 1 9 9 0 2 9 0 13 12 12 9 1 9 9 9 7 9 7 9 7 9
2 8 8
49 13 9 0 12 12 9 2 12 12 9 2 1 9 9 9 7 9 7 12 12 2 12 12 9 2 1 9 9 9 7 9 1 9 15 14 13 1 9 12 9 0 0 1 9 9 1 9 15 2
37 13 9 9 9 0 8 8 7 9 14 13 9 9 9 0 15 13 0 1 9 9 1 9 15 7 14 13 9 9 1 9 0 9 1 9 9 2
55 7 13 9 7 9 14 13 1 9 9 1 9 9 10 9 7 9 15 12 9 13 9 0 1 9 0 1 9 0 1 15 1 12 12 9 2 12 12 9 2 1 9 12 12 9 2 12 12 9 2 9 9 10 9 2
121 7 13 7 10 9 0 1 9 2 7 7 9 15 13 1 9 7 9 0 1 9 0 7 1 7 7 14 15 14 13 15 9 9 9 0 1 15 7 4 9 9 1 9 9 15 2 7 14 13 1 9 0 1 9 0 1 9 9 1 10 13 1 9 9 15 13 15 9 0 1 9 0 2 7 14 13 9 15 1 9 7 13 1 9 9 1 7 9 15 0 1 9 1 9 2 7 13 2 2 14 10 9 13 9 15 1 9 9 9 0 15 13 1 9 7 15 1 9 9 2 2
39 7 13 8 9 0 9 0 0 1 9 9 0 1 9 9 0 2 0 7 9 9 1 9 13 1 9 9 0 1 10 9 15 13 9 15 1 9 0 2
41 7 13 7 15 14 13 9 1 9 0 1 9 9 9 9 9 1 9 9 9 9 0 7 14 13 9 9 0 1 0 1 9 9 7 9 9 0 1 9 9 2
33 7 1 9 9 9 13 8 7 3 9 1 9 0 1 9 9 9 9 0 1 9 1 9 9 15 13 15 9 0 7 9 0 2
2 9 0
37 7 13 9 9 9 1 12 9 1 9 12 0 1 9 1 15 13 7 9 9 1 10 9 0 9 1 9 0 15 13 15 9 9 2 9 2 2
88 7 13 9 1 9 1 9 0 1 9 12 9 15 2 8 8 1 9 7 9 9 2 0 1 0 1 9 8 14 13 9 15 1 9 0 2 7 9 2 9 1 9 2 15 13 9 9 12 1 12 1 9 9 15 7 14 13 9 15 1 9 0 2 7 9 2 9 1 9 7 9 2 0 1 0 1 9 15 14 13 9 15 1 9 9 1 15 2
68 7 13 1 7 9 1 9 9 9 9 10 9 1 9 1 9 0 13 1 12 12 9 2 12 12 9 2 2 7 13 9 1 9 9 2 9 8 2 7 9 2 8 8 2 15 14 13 9 1 9 9 0 1 9 9 1 9 9 9 0 15 13 9 9 9 15 0 2
65 7 13 8 2 2 7 9 13 9 1 9 9 1 9 9 7 9 7 9 9 7 9 15 13 1 9 9 9 9 0 1 9 1 15 0 2 9 1 9 9 9 0 7 0 7 9 1 9 1 9 9 0 1 9 13 9 9 1 9 0 1 15 0 2 2
56 7 13 2 2 14 9 0 1 9 9 9 7 9 13 12 12 9 2 12 12 9 2 9 1 9 9 0 1 15 1 9 12 12 9 2 12 12 9 2 1 15 13 7 9 9 0 9 7 13 9 15 12 12 9 2 2
39 7 13 8 1 7 15 13 9 0 1 8 9 9 1 9 12 9 1 9 9 0 1 9 12 12 9 2 8 8 1 9 9 12 12 9 13 1 9 2
40 7 1 9 9 7 9 2 13 2 2 13 0 9 9 9 0 9 1 9 9 7 9 1 9 0 9 15 12 12 9 1 9 9 9 9 0 1 9 2 2
27 7 13 2 2 14 9 9 9 1 9 13 9 9 1 9 12 1 12 1 9 9 15 13 9 15 2 2
45 13 1 7 9 13 9 0 1 9 0 1 9 0 12 2 12 13 9 9 9 7 9 9 0 7 9 9 0 1 1 9 9 9 7 9 9 9 0 7 9 9 1 9 0 2
47 7 13 9 9 9 1 9 9 7 9 9 15 13 9 9 2 7 13 9 1 9 13 9 12 9 7 9 1 9 1 9 0 13 12 12 9 1 9 12 9 13 15 9 1 9 15 2
8 2 9 1 9 2 8 8 8
66 1 9 1 9 9 0 13 3 9 9 1 8 9 0 9 8 9 2 9 1 8 2 8 9 10 1 12 9 12 2 1 9 9 8 1 8 2 13 15 9 9 9 7 9 8 8 8 8 0 9 9 8 7 9 0 9 8 7 9 9 8 8 9 9 8 2
113 13 9 9 9 9 0 1 9 9 0 9 8 8 1 9 7 13 1 9 8 8 2 2 8 8 13 9 9 0 1 9 8 8 1 0 9 15 7 15 9 1 12 9 13 1 9 7 9 0 7 0 13 15 9 1 8 2 7 9 15 15 15 13 1 8 8 0 8 8 9 1 9 8 8 8 8 8 8 1 8 9 8 8 8 8 8 8 8 8 9 2 7 13 7 13 1 9 7 9 9 9 9 8 8 8 8 8 1 9 8 8 2 2
62 13 1 15 9 9 9 9 8 9 7 13 7 9 8 13 1 9 15 1 2 9 0 8 1 9 13 1 15 9 0 9 2 7 15 13 9 9 7 1 9 1 9 7 9 9 1 9 15 0 7 1 9 0 15 13 15 9 0 7 0 2 2
22 7 13 7 9 9 0 13 1 9 0 14 14 0 15 9 9 7 9 9 7 9 2
62 13 1 15 9 8 9 9 7 13 7 9 15 13 8 9 1 9 7 9 2 0 2 8 8 8 8 8 8 0 1 9 1 9 2 2 7 13 8 9 1 8 12 2 9 7 8 2 8 0 8 8 2 9 7 9 8 2 9 7 9 0 2
62 7 13 9 1 9 2 1 15 13 9 1 9 0 9 0 0 1 9 0 1 15 2 9 9 2 2 14 14 13 13 9 1 9 0 0 1 9 9 0 2 14 9 0 0 1 9 7 13 1 15 7 13 1 9 15 7 14 13 9 9 0 2
32 7 13 8 8 8 1 2 9 9 9 1 9 8 8 2 7 9 7 9 9 9 13 1 9 0 1 9 0 7 9 0 2
59 7 13 9 1 2 9 1 9 1 9 9 15 13 9 0 8 8 8 8 9 13 0 8 8 8 13 0 2 7 0 10 13 10 9 1 9 13 1 8 8 1 9 9 0 9 7 1 9 1 9 8 9 1 9 0 9 0 2 2
33 7 13 1 9 8 8 9 8 7 2 13 3 15 15 8 1 9 1 9 1 9 15 13 9 8 8 9 8 8 8 8 2 2
11 7 13 9 9 15 1 8 9 1 9 2
15 8 13 9 8 1 9 0 2 13 9 0 8 8 9 8
72 9 0 1 9 8 9 8 13 3 9 9 1 9 0 1 9 15 13 9 0 13 9 9 0 1 9 9 8 8 8 8 9 8 8 8 8 7 8 8 8 8 8 7 8 8 8 8 0 2 7 13 9 9 9 8 9 15 8 8 8 8 0 1 9 0 1 9 9 8 9 8 2
63 13 9 9 0 2 9 7 9 9 7 9 7 9 7 9 9 8 8 0 1 9 2 7 13 9 0 1 9 9 0 7 9 9 8 8 9 8 8 1 9 1 9 0 7 9 9 2 7 13 3 1 9 0 2 0 9 7 9 14 13 1 15 2
32 7 13 8 7 2 9 13 1 9 9 1 9 0 1 9 9 0 2 7 13 8 8 8 9 1 15 13 9 1 8 2 2
58 7 1 9 13 9 2 9 9 8 1 9 0 1 9 8 8 2 7 13 7 13 9 9 2 2 13 9 0 1 7 2 9 9 8 13 9 0 1 9 8 0 1 9 8 8 9 1 9 0 13 9 0 8 8 9 9 2 2
9 9 2 9 8 8 13 1 15 2
42 2 1 8 8 8 0 13 9 13 1 9 8 8 9 9 7 9 2 7 15 9 8 8 9 9 8 9 8 2 7 15 13 7 14 13 9 9 8 8 7 9 2
31 1 10 9 7 1 9 15 8 8 2 8 1 0 8 8 2 7 8 1 8 9 9 15 8 1 9 9 8 8 2 2
149 7 13 8 9 13 1 15 2 2 7 8 9 13 9 9 10 9 1 9 15 1 9 7 9 7 9 9 8 8 7 9 8 8 3 7 8 0 8 8 8 7 9 9 0 15 9 9 8 8 7 9 8 8 7 1 8 8 7 9 1 8 8 8 0 8 8 2 15 9 15 1 9 15 9 7 1 15 0 1 9 0 13 7 13 8 1 9 8 0 7 13 1 9 9 8 8 2 8 9 8 9 9 8 8 8 8 7 9 9 0 1 9 7 9 1 9 15 7 9 9 15 0 8 8 8 1 9 1 1 9 15 8 7 8 8 1 9 8 8 8 8 1 0 15 8 8 8 2 2
60 13 15 8 13 2 2 13 9 8 9 8 9 8 8 9 0 0 8 8 0 0 8 8 9 9 0 1 9 0 8 8 2 7 8 1 9 13 9 7 9 13 7 13 9 8 8 0 7 0 1 9 8 0 2 8 8 10 9 15 2
56 2 9 9 0 1 8 8 8 8 1 9 8 2 7 9 15 0 8 8 9 2 7 9 9 8 8 1 9 0 0 8 15 9 9 8 8 9 1 9 9 0 0 15 13 1 9 9 9 7 9 9 8 8 8 0 2
19 2 9 1 9 9 13 2 7 14 9 13 15 2 8 8 9 9 0 2
36 2 8 9 1 9 9 0 1 9 2 8 8 0 15 8 9 0 2 7 9 15 1 8 9 1 15 8 9 0 1 1 9 9 1 15 2
21 9 9 1 9 0 8 8 2 7 10 9 13 7 13 9 1 9 1 9 2 2
20 1 9 15 13 8 7 9 15 2 1 9 0 1 9 15 7 9 15 2 2
25 7 13 1 9 9 15 13 1 9 0 8 8 2 7 13 9 9 1 7 15 9 9 9 15 2
63 7 13 8 9 9 2 7 13 2 2 9 13 1 8 13 0 1 9 1 9 9 7 7 15 0 9 1 9 0 2 2 7 14 13 9 1 9 14 13 0 9 2 8 8 13 13 15 9 0 2 7 13 1 15 9 9 9 1 9 7 9 2 2
33 7 13 1 7 9 2 14 13 1 9 9 1 9 2 2 0 7 15 0 2 15 13 0 1 8 8 9 0 8 8 0 2 2
77 7 13 8 7 2 8 8 7 0 8 8 1 15 9 9 9 15 9 1 9 15 2 2 2 2 2 8 8 13 15 9 13 9 1 9 8 8 0 8 8 0 2 8 8 9 7 15 1 8 9 9 1 9 0 7 7 15 1 15 13 9 15 1 7 13 9 1 9 8 8 2 13 1 9 9 2 2
10 7 13 8 8 1 9 9 1 9 2
35 7 13 8 7 2 9 13 9 8 8 9 0 1 9 2 7 9 1 9 8 8 2 2 7 13 9 9 1 15 13 1 9 8 8 2
36 7 13 0 7 15 2 13 1 9 0 7 13 9 7 7 8 9 9 0 13 1 9 9 8 1 9 0 7 1 8 9 1 9 0 2 2
12 8 2 9 9 0 7 9 0 1 9 13 9
51 13 9 9 9 0 8 8 1 0 1 2 9 2 7 8 9 0 1 9 0 1 9 9 15 8 8 8 0 8 8 8 7 9 9 15 1 9 2 7 7 15 14 13 1 9 9 0 0 1 9 2
48 7 13 7 9 0 1 9 0 0 7 0 2 7 13 7 13 9 9 0 0 1 9 13 1 9 15 2 7 9 0 1 9 1 9 7 7 13 9 0 9 9 0 1 10 0 7 13 2
31 7 13 8 9 0 0 9 1 9 9 7 7 9 0 1 9 9 0 1 15 7 7 9 9 0 1 9 13 13 9 2
43 8 14 13 0 1 9 13 9 9 0 8 8 7 9 9 15 14 13 9 15 1 8 8 2 9 0 1 9 9 0 0 2 0 1 7 15 14 13 0 0 1 9 2
32 7 13 8 1 9 1 9 0 1 8 9 1 0 2 1 9 9 1 9 15 13 15 9 8 8 1 15 1 9 0 2 2
103 7 13 2 1 9 8 8 8 9 13 1 9 0 2 9 8 8 1 15 9 0 14 8 9 15 7 8 9 9 0 2 9 13 9 8 8 1 9 7 1 15 2 7 14 15 0 1 9 7 1 15 9 1 9 12 9 1 9 9 9 7 10 9 0 8 8 8 7 8 8 2 2 7 13 2 14 13 8 8 1 9 8 8 2 7 1 9 8 8 7 15 13 9 9 1 9 0 13 9 8 8 2 2
44 7 13 8 7 15 2 13 9 9 1 9 9 9 2 0 1 8 8 2 1 10 13 9 9 1 1 9 2 7 1 0 7 8 9 0 1 9 9 9 0 9 9 2 2
51 7 13 7 15 13 9 1 9 9 9 0 1 0 9 13 2 1 9 9 0 0 13 1 9 9 2 7 9 9 9 2 7 13 9 1 9 9 14 13 0 1 9 1 9 9 9 0 1 9 9 2
6 9 9 0 1 9 9
66 13 9 0 13 1 15 2 9 9 2 1 9 9 0 0 9 1 9 9 9 7 14 13 10 9 1 1 9 0 1 9 9 9 0 7 14 13 9 0 9 0 15 13 14 13 9 1 15 9 1 9 9 1 9 15 13 1 9 9 9 9 12 1 9 9 2
41 7 13 9 9 9 15 1 9 9 1 9 0 7 8 7 9 1 9 9 0 7 0 1 9 0 1 9 0 7 9 15 13 15 9 9 9 1 9 0 0 2
44 13 8 8 9 9 9 0 1 9 8 8 9 9 13 1 15 9 0 1 9 9 0 1 9 9 0 1 9 9 15 13 15 9 9 9 1 7 9 9 0 13 1 9 2
82 7 13 8 1 9 15 7 15 13 9 9 1 9 9 8 8 8 9 0 9 0 1 9 9 15 13 1 9 0 9 1 9 0 1 9 9 0 9 15 13 1 9 0 7 0 7 9 9 15 13 1 9 9 15 13 15 9 9 9 2 7 7 8 14 13 1 15 13 9 9 1 9 1 9 9 0 15 13 15 9 0 2
49 13 8 7 15 13 9 9 0 1 8 1 9 9 0 7 13 15 1 7 13 1 9 15 1 9 9 9 1 9 0 1 9 1 9 0 1 9 0 1 9 9 15 13 7 13 1 9 0 2
58 7 13 9 9 7 9 9 9 1 9 0 13 1 7 9 9 0 13 1 9 9 9 0 15 13 9 9 15 1 9 1 15 1 9 9 15 13 1 9 9 9 9 9 0 15 13 9 15 1 9 15 1 9 15 1 9 0 2
49 7 13 9 9 1 9 15 1 9 9 7 9 13 1 9 9 9 8 7 9 9 0 9 1 9 0 8 1 9 9 15 13 9 9 0 7 9 9 8 8 1 9 1 9 9 10 9 2 2
12 7 13 9 9 9 0 9 1 9 0 0 2
42 7 13 7 9 9 9 1 9 0 13 7 15 1 9 9 9 0 1 9 1 7 13 9 9 8 1 9 9 0 1 9 9 7 9 7 9 7 9 7 9 0 2
31 7 13 9 1 9 9 9 1 9 1 8 7 8 1 9 9 0 1 9 0 9 1 9 9 1 10 9 1 9 0 2
40 7 13 2 9 9 2 7 9 13 9 0 1 9 0 1 9 9 1 9 9 9 0 1 9 7 9 0 14 13 1 15 14 0 7 9 1 0 14 13 2
22 7 14 13 9 9 0 9 1 9 9 9 9 0 9 15 1 8 9 9 0 2 2
16 7 15 1 9 9 1 9 1 0 7 9 0 1 9 0 2
14 9 0 0 0 2 9 9 0 7 9 15 9 1 9
79 13 9 8 8 9 9 0 0 0 1 9 1 2 9 2 9 1 9 9 0 8 8 9 1 9 0 1 9 1 15 1 14 9 0 1 7 3 9 0 0 9 14 13 9 15 1 9 9 1 9 0 7 7 15 14 13 1 9 9 1 9 2 7 7 9 0 13 1 9 7 9 15 13 15 1 9 9 0 2
44 7 13 2 14 14 13 9 9 9 9 9 0 1 9 0 0 15 9 15 13 15 9 9 9 0 1 9 0 7 13 9 9 7 9 3 13 1 15 13 1 15 1 9 2
105 7 13 7 9 13 1 9 15 13 9 9 1 9 0 1 9 0 7 13 1 9 15 1 9 9 7 13 1 9 9 0 1 7 1 9 9 0 7 13 9 15 1 9 9 0 1 9 1 9 0 1 9 15 1 9 0 7 9 9 1 0 1 9 1 15 1 9 0 13 15 9 0 1 9 9 10 13 1 15 1 9 2 7 9 9 1 9 1 9 1 9 9 9 1 15 1 9 9 9 1 9 9 15 8 2
101 7 13 8 7 9 1 10 9 13 1 9 7 1 9 9 8 1 9 9 9 9 1 9 0 13 9 9 7 9 9 7 9 9 1 9 9 0 1 9 9 9 9 1 9 0 7 9 9 8 0 0 1 9 14 13 3 9 0 1 9 0 1 9 1 9 15 13 15 0 1 9 1 9 9 15 7 14 13 8 1 9 9 9 14 13 9 1 9 15 1 9 0 1 9 9 7 9 9 9 0 2
77 7 1 9 9 9 1 9 9 9 1 9 13 9 9 0 0 2 10 9 14 13 9 15 1 9 0 1 9 0 7 7 9 0 13 1 9 13 1 9 9 9 9 7 1 15 7 7 9 9 13 1 9 9 0 9 7 9 14 13 1 9 7 7 1 9 9 15 13 1 9 0 1 9 1 9 15 2
81 7 1 9 0 0 1 9 9 0 7 15 13 1 0 13 15 1 9 9 0 13 7 3 9 1 9 0 7 9 1 9 1 9 10 9 1 9 9 9 0 9 9 7 14 13 1 9 9 9 9 1 9 9 0 2 15 13 1 15 9 2 1 9 0 7 9 1 9 9 9 0 7 9 9 7 9 9 0 7 0 2
97 7 1 9 1 9 9 1 9 9 9 7 9 9 0 1 9 0 7 15 13 15 9 0 1 9 13 8 7 9 13 1 9 9 10 9 7 15 13 9 9 9 0 1 15 12 12 9 1 9 15 1 9 0 7 13 7 3 9 1 9 0 1 9 0 1 9 9 1 9 9 0 1 9 1 15 1 9 7 9 1 9 7 15 13 9 1 10 9 7 14 9 1 10 9 1 9 2
49 7 13 8 8 8 9 9 9 2 8 2 1 9 9 0 0 1 9 9 0 1 9 9 0 0 0 7 9 13 15 13 9 9 9 9 15 13 9 15 7 14 3 9 0 14 13 1 15 2
35 7 13 2 8 8 1 9 9 1 9 1 9 9 0 1 9 7 7 13 9 0 1 9 0 8 8 8 8 3 1 9 9 1 9 2
7 9 9 9 9 1 9 9
36 13 9 8 8 8 9 9 0 9 9 9 9 1 9 9 9 0 0 1 7 15 14 13 9 10 9 1 9 9 0 15 13 1 9 0 2
40 7 13 8 7 3 9 9 1 9 9 9 1 9 2 7 7 9 0 13 9 9 0 0 1 15 9 9 1 9 1 9 0 1 9 9 1 9 0 2 2
23 7 14 13 9 1 9 1 9 15 1 9 9 9 1 9 15 13 1 9 1 10 9 2
89 7 13 9 8 8 14 13 9 1 9 15 0 8 8 9 12 2 12 0 1 9 9 9 9 7 9 9 1 9 9 9 0 1 9 9 1 9 9 8 8 7 0 8 8 1 9 9 8 8 1 8 7 13 8 1 7 9 0 7 0 13 1 9 9 9 0 0 1 9 1 9 9 9 9 0 7 9 1 9 1 10 9 1 9 9 0 1 0 2
4 9 1 9 9
25 1 9 8 2 8 8 2 9 9 2 1 9 9 0 1 9 9 9 2 13 9 0 1 9 2
33 13 9 0 9 0 9 1 9 9 15 13 1 9 1 9 0 1 9 9 7 9 9 9 7 9 9 9 7 9 9 9 0 2
62 13 8 2 8 9 9 9 7 13 1 9 1 9 9 9 0 2 7 13 9 15 1 9 9 9 1 9 15 1 9 1 9 0 1 9 0 2 7 13 2 1 0 9 2 1 9 9 1 9 9 1 1 9 9 0 2 1 1 9 7 9 2
51 7 13 1 9 13 15 9 9 9 9 7 9 9 0 9 12 2 12 0 7 9 9 0 2 15 13 15 9 2 13 1 9 9 2 1 9 7 9 9 0 1 15 2 7 7 1 9 0 2 2 2
87 2 7 1 9 1 9 9 1 9 0 1 9 9 1 9 1 9 15 1 9 9 7 15 13 1 1 12 12 9 2 13 7 3 9 13 9 15 0 1 9 9 9 9 9 1 9 0 1 9 9 0 2 1 9 15 1 9 15 1 9 2 2 2 7 13 9 9 1 9 9 15 1 10 9 2 2 7 15 1 15 13 9 9 9 2 2 2
3 7 13 2
49 2 8 8 14 8 9 1 8 8 0 2 9 9 9 0 0 2 7 3 9 9 9 0 8 8 2 2 1 9 1 15 1 9 0 1 9 0 0 1 9 9 9 0 7 9 9 9 2 2
83 1 9 0 13 8 2 8 8 2 9 0 1 9 9 15 1 9 0 9 1 9 9 1 9 15 1 9 1 9 0 1 9 2 7 9 9 15 13 15 9 0 2 9 8 8 9 9 1 0 9 7 1 9 15 9 9 7 9 7 9 7 9 1 9 2 7 3 8 9 9 9 9 0 7 9 9 1 9 9 9 1 15 2
7 9 9 1 9 9 0 0
35 13 9 9 1 9 9 0 1 9 0 9 12 2 12 0 1 9 9 9 1 9 0 1 15 1 9 2 9 9 9 9 1 15 2 2
40 7 13 9 9 9 9 9 7 9 9 1 9 8 8 8 8 2 2 10 9 13 9 9 2 7 15 13 9 9 7 13 1 9 0 1 9 9 0 2 2
64 7 1 7 9 9 9 0 7 9 1 9 0 8 8 1 9 9 1 9 0 8 8 8 2 7 13 9 1 9 0 1 9 2 8 7 9 9 7 9 0 0 13 7 9 0 1 9 2 13 1 9 9 9 9 0 1 9 1 9 1 9 0 2 2
31 7 1 0 7 13 9 9 0 9 12 2 12 0 2 1 7 13 9 0 1 9 0 1 7 13 9 9 12 9 0 2
18 8 1 9 9 9 0 2 9 14 13 9 1 9 7 13 1 9 15
55 13 9 8 8 9 9 9 9 12 2 12 0 9 0 1 9 0 2 7 13 7 9 9 1 9 0 9 0 7 13 1 9 3 2 7 7 15 9 1 9 0 7 9 1 15 2 7 13 1 9 9 1 9 15 2
33 7 13 9 9 9 1 7 9 0 13 9 9 0 1 12 12 9 1 0 9 9 2 7 13 1 9 9 0 1 9 0 0 2
37 7 1 9 15 2 13 9 8 8 8 9 9 7 9 13 1 9 9 0 1 9 9 0 2 7 7 15 13 0 12 12 9 9 1 10 9 2
23 7 13 9 9 9 8 8 8 7 9 14 13 0 1 9 0 2 7 9 1 9 0 2
6 9 13 9 1 9 9
38 13 8 8 9 9 0 1 9 9 7 9 9 9 0 2 8 2 7 9 13 1 9 0 1 9 1 9 9 2 7 1 9 1 9 0 1 15 2
59 7 13 2 1 9 0 1 2 9 2 7 15 7 14 9 9 14 13 9 2 7 13 1 15 13 15 1 9 9 0 1 9 13 13 9 15 9 12 2 1 9 9 9 0 8 8 2 1 9 9 15 13 9 9 8 8 1 8 2
48 7 13 7 10 9 1 9 1 9 1 9 2 13 7 13 7 14 9 9 7 9 15 1 15 2 7 9 15 1 9 15 13 1 10 9 7 15 14 13 0 9 1 0 9 0 1 9 2
43 7 13 7 9 13 9 0 1 9 0 2 7 14 13 9 0 1 9 7 9 9 15 1 9 2 15 13 0 7 13 9 1 15 1 9 15 1 9 1 9 9 15 2
16 9 9 1 2 8 2 1 9 9 1 9 9 9 1 9 9
35 13 9 9 1 9 1 9 9 1 2 8 2 3 1 9 9 9 9 0 1 9 9 0 15 13 0 9 15 1 12 9 1 9 0 2
49 7 13 9 9 9 0 1 7 13 8 1 9 0 1 9 9 9 0 1 9 12 1 12 9 1 0 9 2 9 2 1 9 9 9 1 9 0 7 15 9 15 13 1 15 9 1 9 0 2
49 7 13 9 2 8 2 1 8 9 9 2 9 2 1 9 9 9 14 7 9 0 1 2 8 2 13 1 8 3 1 7 2 9 14 13 9 9 9 1 9 0 1 9 1 9 2 9 2 2
18 7 13 0 2 2 9 0 7 7 4 3 9 0 1 15 1 2 2
40 1 9 15 13 8 11 8 8 9 9 9 3 2 7 9 8 14 13 1 9 15 0 9 12 9 0 9 9 9 9 9 0 9 1 9 0 7 9 0 2
19 7 13 8 2 2 14 15 14 13 1 9 0 9 0 1 9 0 2 2
35 7 13 9 9 1 9 9 7 10 9 14 13 1 9 1 9 0 1 9 15 1 9 0 2 15 13 15 2 8 2 1 8 9 0 2
35 7 13 8 1 15 7 13 14 13 9 1 9 9 9 9 1 9 12 9 0 1 9 0 9 1 9 7 13 2 14 14 13 9 2 2
20 7 13 7 9 9 1 9 0 1 9 9 14 13 9 0 13 1 9 8 2
27 14 7 9 9 7 9 0 8 8 8 3 13 7 15 14 13 0 9 1 2 8 2 1 9 9 9 2
9 7 13 8 2 14 13 9 9 2
15 14 13 9 1 10 9 1 0 9 7 14 13 15 2 2
34 7 13 0 1 9 0 0 9 9 1 12 9 1 9 9 9 1 9 7 9 9 9 1 9 0 7 9 1 9 9 13 9 9 2
46 7 1 10 9 13 9 9 0 8 8 3 1 9 9 2 8 2 9 9 15 1 12 9 0 1 0 1 9 1 9 15 2 9 8 8 8 2 8 8 9 0 1 9 9 2 2
36 7 13 9 9 0 8 8 1 9 15 1 9 9 9 7 7 15 13 7 15 4 3 0 15 13 1 2 8 2 9 15 1 9 9 9 2
10 7 13 8 2 1 9 8 0 2 2
16 7 9 0 13 9 15 1 9 9 15 13 15 9 0 2 2
23 2 8 2 0 2 0 2 0 13 1 9 1 9 9 9 1 0 8 8 13 12 12 9
48 13 9 0 1 0 3 7 15 13 9 8 0 1 12 9 0 15 2 8 2 8 7 2 8 2 9 0 7 2 8 2 8 2 1 9 9 9 9 1 0 13 9 15 8 12 12 9 2
29 7 13 9 1 9 0 1 9 8 8 2 7 15 8 13 0 9 2 7 13 1 9 1 9 9 1 9 9 2
38 7 13 7 9 13 1 9 0 9 9 1 0 7 13 9 9 1 9 9 13 9 0 1 0 12 12 9 0 1 9 0 7 0 12 12 9 0 2
10 7 13 1 7 9 9 15 12 9 2
50 7 13 9 1 9 0 1 9 2 9 2 12 2 7 9 0 0 2 1 15 2 8 2 8 7 2 8 8 2 9 8 2 8 13 8 8 2 13 1 9 1 9 9 9 1 9 0 1 0 2
23 7 13 0 12 12 9 0 1 9 0 2 7 13 9 15 1 15 1 12 12 9 0 2
30 7 13 9 8 0 0 0 1 9 13 9 0 0 1 9 9 0 1 15 13 9 1 9 9 7 9 0 1 0 2
19 7 13 9 0 8 8 1 9 2 9 0 2 12 2 9 1 10 9 2
53 1 9 15 13 9 9 7 9 0 0 9 8 8 1 9 15 9 0 0 0 1 9 7 9 2 7 10 9 13 9 9 1 9 0 7 9 0 7 9 13 9 1 9 1 9 15 1 9 9 7 9 2 2
82 7 13 9 8 15 13 3 9 0 0 1 9 9 1 9 9 0 8 8 8 15 13 9 1 7 10 9 13 9 0 7 0 1 9 9 7 9 0 2 9 15 13 9 1 9 7 9 9 0 7 1 9 15 1 9 0 2 7 13 1 7 10 9 0 1 9 7 9 0 15 13 9 9 7 9 0 1 9 0 1 0 2
69 7 13 1 10 9 0 1 8 9 1 1 12 9 0 7 0 9 9 8 1 10 13 9 9 7 9 2 1 15 13 9 1 9 1 0 9 7 9 8 1 10 9 7 9 9 7 9 9 0 7 9 8 0 1 10 13 1 9 9 9 9 9 7 9 1 0 7 9 2
78 7 14 13 1 9 10 9 12 9 7 9 0 7 0 13 1 9 9 0 7 9 0 1 9 15 9 1 9 7 9 0 7 9 7 9 7 9 9 0 7 9 9 9 0 7 9 9 0 7 9 9 2 7 13 1 10 9 7 9 7 9 9 0 7 0 1 9 1 0 9 9 0 1 9 9 7 9 2
37 7 13 9 9 0 0 13 9 7 9 7 8 2 1 9 0 1 9 9 0 1 9 9 7 9 2 7 13 9 9 0 1 9 0 1 0 2
7 9 9 8 1 9 9 0
41 13 9 9 0 8 8 2 12 9 2 1 9 0 1 9 13 13 15 1 9 0 1 9 9 7 9 2 7 1 9 9 7 0 9 9 2 9 1 9 0 2
38 7 13 9 0 14 13 9 15 1 9 8 9 15 2 7 13 9 9 8 8 7 9 2 13 1 9 0 2 1 9 15 1 9 1 9 9 2 2
83 7 13 8 0 2 7 13 1 15 8 9 2 7 13 9 0 2 1 7 15 13 9 1 9 15 12 9 2 7 1 9 15 13 7 13 2 7 13 9 9 15 0 15 13 1 9 1 15 1 9 15 1 9 1 9 1 9 0 1 9 0 1 9 2 15 14 13 1 9 15 1 9 9 15 8 8 2 9 9 9 8 8 2
16 7 13 8 1 9 1 12 9 7 13 9 15 1 9 15 2
59 7 13 9 0 7 9 14 13 1 9 1 9 9 9 1 9 9 0 8 1 15 2 2 9 1 9 15 0 1 9 1 9 15 9 0 1 9 0 0 0 1 9 0 1 9 9 15 13 12 8 7 9 1 9 0 1 9 2 2
61 7 1 9 1 7 15 14 13 1 9 0 15 13 9 15 9 1 9 0 2 7 14 9 9 0 13 7 9 2 14 13 1 9 0 1 9 15 0 0 2 7 7 9 0 13 1 9 15 0 2 1 9 0 9 0 1 9 1 15 2 2
24 7 13 7 9 2 14 13 1 9 9 0 0 1 9 0 9 0 7 0 15 13 1 9 2
8 9 9 0 13 9 15 1 9
15 13 9 2 8 2 0 1 0 9 9 0 1 9 0 2
18 13 9 9 0 15 13 9 9 15 0 7 9 9 9 9 1 15 2
19 7 13 1 7 9 9 0 15 1 9 15 1 9 7 9 15 1 9 2
24 13 9 9 14 12 9 9 9 9 7 9 1 9 9 7 9 1 9 3 7 13 1 9 2
10 9 9 2 9 13 1 9 1 9 15
58 13 9 9 9 2 9 9 9 0 8 8 15 13 1 15 7 9 13 9 0 1 9 7 13 1 9 1 9 9 0 2 7 13 2 14 15 9 0 13 1 9 2 7 9 13 1 9 1 10 13 15 7 15 9 9 7 9 2
49 7 13 9 9 8 1 7 9 1 9 13 9 0 7 13 1 9 1 9 1 9 1 2 9 2 7 13 2 2 14 9 9 14 13 9 0 14 1 8 15 13 9 0 0 1 9 0 2 2
60 7 13 9 7 9 10 13 0 1 9 0 7 9 2 9 15 9 1 9 9 1 9 9 9 9 1 2 9 9 2 7 9 1 9 9 1 9 9 0 1 9 1 9 9 1 9 9 7 9 9 0 1 9 9 7 9 9 7 9 2
14 9 9 0 8 2 1 9 9 14 13 1 9 9 9
12 13 9 0 9 12 2 12 9 15 1 0 2
27 7 13 9 0 1 9 9 9 9 8 8 1 9 3 1 9 9 9 8 8 1 0 1 9 1 8 2
16 7 13 9 9 0 8 8 8 1 10 9 1 9 1 9 2
45 7 13 2 8 0 7 0 1 10 9 2 7 13 8 2 15 13 7 13 7 7 13 2 2 7 15 13 7 13 7 7 13 2 8 1 9 9 14 13 1 9 9 9 2 2
24 7 13 8 9 8 9 1 9 0 13 15 8 0 7 13 15 9 1 9 1 9 0 0 2
15 7 13 7 2 8 13 0 7 14 0 1 10 9 2 2
30 7 13 2 8 8 7 13 9 1 9 0 0 7 9 0 2 0 2 7 9 0 9 0 1 9 7 14 9 2 2
28 1 9 15 13 9 9 0 9 8 8 2 14 9 1 0 13 0 7 15 13 0 7 13 9 1 9 2 2
33 7 13 9 8 2 14 9 1 9 0 13 1 9 7 13 0 2 7 9 0 14 13 0 9 1 9 0 7 13 9 15 2 2
61 7 13 8 14 13 9 15 8 1 7 15 13 15 9 9 0 1 1 9 12 1 9 9 9 1 9 9 2 7 9 9 9 8 9 0 1 9 2 13 13 1 9 9 1 9 0 8 8 7 13 9 15 1 10 13 15 1 2 9 2 2
24 7 13 8 2 8 7 8 7 9 8 14 8 8 9 8 8 8 8 8 1 15 9 0 2
11 2 8 2 0 13 9 9 15 12 12 9
43 13 9 2 8 2 0 1 9 7 9 9 9 0 1 9 15 13 15 1 9 12 12 9 2 12 12 9 2 7 15 1 9 12 5 1 0 1 9 1 9 9 9 2
20 7 14 13 8 1 9 9 9 1 9 0 8 8 0 9 7 9 9 0 2
67 7 13 9 1 9 13 15 1 9 7 9 9 1 9 14 13 9 1 9 9 7 13 9 9 9 1 0 9 0 7 0 1 9 2 1 15 9 8 0 2 9 7 9 0 0 7 9 0 0 7 9 9 2 9 9 0 0 2 7 9 0 0 7 9 8 8 2
81 7 13 9 8 1 9 7 9 15 13 9 15 0 12 8 9 2 1 12 8 9 2 14 13 1 9 2 0 1 9 12 12 9 2 12 12 9 2 1 9 0 0 12 5 13 9 12 9 2 7 9 0 1 9 12 12 9 2 12 12 9 2 1 9 0 2 12 5 0 1 9 9 7 9 0 1 9 0 0 2 2
8 9 7 9 9 0 13 9 9
35 13 9 0 2 0 9 0 1 9 0 1 8 9 9 1 9 9 0 0 1 12 9 7 13 9 9 9 1 9 9 0 1 9 0 2
26 7 13 9 9 9 8 2 8 8 8 1 9 9 0 7 14 13 15 9 1 9 9 0 1 9 2
110 13 8 8 2 8 8 9 9 9 0 7 0 1 9 9 0 0 1 7 9 0 1 9 13 9 0 1 9 12 0 7 13 12 8 9 9 12 1 9 9 9 15 12 2 12 5 9 1 9 12 1 9 9 9 0 1 9 1 9 9 9 9 0 7 9 0 1 9 0 7 13 9 9 1 9 9 1 12 8 9 9 12 1 12 8 9 9 7 13 0 9 0 1 9 0 1 9 7 9 7 9 9 15 7 9 8 7 9 15 2
64 7 1 9 8 8 8 1 9 0 7 14 13 12 8 9 9 12 1 9 9 15 12 5 1 9 12 1 9 9 8 8 1 9 7 9 15 7 9 9 8 7 9 15 7 9 0 1 1 13 9 0 1 9 1 9 7 9 0 7 9 7 9 15 2
66 7 13 8 2 8 8 9 0 1 9 0 1 9 0 1 9 0 7 9 13 9 9 0 12 1 9 9 7 3 9 15 13 9 9 15 1 8 1 9 1 9 15 1 8 1 0 9 7 0 9 1 9 9 0 1 8 0 15 9 1 9 9 1 9 9 2
15 9 0 13 7 9 0 2 9 0 2 1 2 9 9 2
60 13 9 13 9 2 9 9 0 7 9 2 1 9 8 0 0 2 13 2 9 2 9 1 15 9 12 2 12 0 1 9 0 2 7 2 9 0 0 2 15 13 8 0 9 15 13 1 9 9 1 9 9 15 2 13 9 1 9 2 2
81 7 13 9 1 9 13 15 9 1 12 9 0 1 9 2 9 0 7 0 1 9 0 2 2 13 1 7 9 13 3 2 1 9 9 8 7 9 9 0 7 9 0 7 9 9 0 7 0 8 7 9 0 2 7 2 9 0 8 2 7 15 13 1 9 7 9 9 7 9 0 9 1 9 9 0 8 1 9 9 0 2
56 7 13 9 15 13 1 9 12 9 0 7 2 9 9 7 9 9 2 0 1 15 8 1 8 2 9 1 9 15 0 7 9 15 0 14 13 1 9 9 0 9 15 15 13 15 7 13 15 9 0 7 9 15 0 2 2
54 7 13 1 9 2 9 0 7 0 1 9 0 2 7 10 9 15 2 13 15 7 13 15 9 9 0 0 13 9 15 0 1 9 9 0 1 9 9 9 7 9 9 7 9 1 15 0 7 9 1 9 9 2 2
62 7 13 2 9 2 7 2 15 13 7 14 13 1 9 9 2 9 1 9 9 0 1 0 0 2 7 9 0 7 9 7 9 0 2 14 13 7 13 1 7 15 9 7 9 7 9 9 2 7 1 15 13 9 0 1 9 1 9 15 0 2 2
21 7 15 9 0 1 7 9 0 15 13 1 9 13 7 13 1 2 9 0 2 2
13 9 13 1 9 9 7 8 9 1 9 1 9 9
22 13 9 0 1 9 0 9 9 9 1 9 9 9 0 2 9 9 9 1 9 9 2
75 7 13 8 1 9 2 1 9 15 9 9 12 2 12 0 1 9 7 1 15 1 8 2 2 7 9 9 9 1 9 1 9 7 13 1 9 0 1 15 7 9 9 2 8 8 8 9 9 15 8 8 1 9 2 2 0 1 2 7 9 8 7 9 13 1 9 7 7 9 13 1 9 9 0 2
15 7 3 9 0 1 9 1 9 9 0 7 8 0 2 2
47 7 13 8 7 15 14 13 1 9 1 9 9 9 0 7 1 8 14 13 1 9 0 1 9 9 15 13 15 8 8 9 0 1 9 0 1 9 1 9 0 1 9 7 9 1 9 2
11 9 9 1 9 9 2 8 8 2 1 9
52 13 8 8 9 9 0 1 9 1 9 9 9 15 13 15 9 0 1 9 0 7 0 1 9 9 9 2 8 8 2 2 8 8 1 7 13 9 9 0 13 0 1 9 15 13 15 9 0 1 9 9 2
22 7 13 9 0 9 7 9 9 15 13 15 9 13 1 12 12 9 1 9 1 9 2
18 7 13 8 8 9 1 9 9 1 9 1 9 0 1 9 0 8 2
12 9 2 8 8 2 1 0 9 0 2 12 9
39 13 8 2 8 8 9 9 9 0 1 9 8 8 7 9 0 1 9 14 13 9 9 0 9 12 9 0 1 9 9 9 7 9 1 9 15 1 9 2
17 13 8 7 9 13 1 10 9 1 7 13 9 9 12 12 9 2
32 13 8 1 9 0 1 2 9 9 2 7 9 13 2 8 2 1 10 9 7 9 9 13 9 9 9 9 0 12 8 9 2
62 7 1 15 7 13 8 0 14 13 1 9 8 8 7 13 1 9 0 13 8 7 9 0 13 1 9 12 1 12 12 9 8 8 1 9 9 0 2 7 13 10 9 1 9 0 2 9 7 9 0 1 9 13 9 7 14 13 9 13 0 9 2
29 1 9 1 9 9 9 0 1 9 1 9 7 9 9 1 1 12 12 9 7 14 13 8 8 10 0 1 9 2
38 13 8 7 15 14 13 3 9 9 0 0 9 12 9 8 8 9 9 9 1 9 0 12 7 9 9 9 9 7 9 9 1 9 9 1 9 9 2
8 9 0 1 9 9 1 9 11
38 13 1 9 0 1 9 0 9 9 9 15 13 15 9 2 8 2 0 1 9 9 1 9 0 2 8 12 2 9 11 1 9 13 1 12 12 9 2
41 7 13 8 8 8 9 9 9 9 2 8 2 7 9 14 13 1 9 12 12 9 0 7 13 9 1 9 9 9 1 9 9 9 7 9 0 8 8 8 0 2
20 7 13 7 9 14 13 1 9 15 1 9 9 1 9 8 8 0 1 9 2
24 7 13 7 9 14 13 1 9 1 12 12 9 0 1 9 0 7 1 12 12 9 1 8 2
26 7 13 7 9 14 13 1 9 1 12 5 1 9 15 1 9 0 0 1 1 7 13 1 10 9 2
11 9 9 9 0 13 9 9 1 9 15 0
21 13 9 12 2 12 0 1 9 9 1 9 1 9 1 9 9 9 0 7 0 2
31 7 13 9 1 9 0 8 8 8 9 9 9 9 2 7 13 15 1 9 0 8 8 9 9 0 1 9 9 9 0 2
34 7 13 8 8 8 7 9 13 1 9 9 0 1 9 7 8 1 9 9 9 7 13 1 9 9 0 7 9 7 9 9 1 9 2
30 7 13 7 9 15 13 9 15 1 9 0 13 1 9 9 7 9 1 9 7 15 1 9 9 9 1 9 9 0 2
28 7 13 7 9 15 13 9 15 1 9 0 13 1 9 15 13 7 13 15 9 1 9 9 9 0 7 0 2
37 7 13 1 9 10 9 15 13 1 9 9 1 9 1 9 0 2 0 1 7 9 0 7 0 13 9 9 0 0 1 9 0 1 9 9 9 2
21 7 13 1 10 9 9 9 1 9 10 9 0 10 13 1 15 1 9 7 9 2
13 0 0 13 9 9 1 9 9 9 9 0 1 9
37 13 12 9 1 9 0 1 9 0 9 9 0 1 9 0 1 9 0 13 1 15 1 9 9 9 0 1 9 0 1 9 9 9 0 1 15 2
26 7 13 0 7 15 13 9 9 0 1 10 9 7 7 8 8 1 9 7 9 9 9 9 1 9 2
51 7 13 9 9 9 0 9 8 8 1 9 9 0 7 13 1 9 9 0 1 9 9 1 9 1 9 9 9 1 9 9 0 1 9 9 1 9 8 7 9 0 2 9 1 9 0 7 1 9 9 2
60 7 13 9 7 9 9 1 9 1 9 9 13 9 0 7 0 1 9 9 0 1 9 12 1 9 9 9 0 7 0 1 9 9 1 9 0 1 9 0 7 15 13 15 1 9 2 9 1 9 9 9 0 1 9 0 7 0 1 15 2
70 7 13 9 9 1 9 7 13 9 14 13 1 9 0 7 0 1 9 1 9 9 0 1 9 7 9 9 9 0 1 9 2 7 13 0 0 9 15 0 1 0 9 0 1 9 9 0 7 9 15 2 7 13 7 9 0 1 9 9 15 1 9 7 9 0 7 13 9 15 2
36 7 13 0 9 7 15 1 9 1 7 9 14 13 9 1 9 9 9 1 9 7 14 13 1 9 7 13 9 7 13 15 1 9 1 9 2
59 7 13 9 1 9 9 9 9 0 0 1 9 1 9 9 1 9 9 0 7 13 9 9 0 0 1 9 8 8 9 9 1 9 9 12 9 9 13 1 15 9 0 1 9 9 1 9 9 7 1 9 0 9 15 7 1 9 0 2
45 7 13 0 15 1 7 13 9 9 9 9 9 0 9 9 1 9 10 14 13 1 12 12 9 1 9 9 9 1 9 9 1 9 0 0 1 9 1 9 9 15 1 9 2 2
40 7 13 9 0 14 13 9 1 10 13 15 9 9 0 0 1 9 9 0 1 9 9 0 1 9 7 9 8 8 9 9 0 1 9 10 9 1 9 0 2
55 7 13 1 9 9 1 9 9 9 9 0 1 9 9 9 9 15 13 1 12 9 0 1 9 0 1 9 7 1 9 12 9 1 9 13 9 15 1 12 1 9 7 13 9 9 9 9 0 0 2 0 0 9 0 2
12 9 2 8 13 1 9 0 1 9 0 1 9
26 13 9 9 0 8 8 9 1 9 0 7 0 1 9 9 0 0 1 9 0 15 9 0 1 9 2
53 7 13 1 9 13 15 9 0 0 1 9 15 0 1 9 9 9 12 2 12 0 7 9 0 0 1 9 9 0 1 9 0 9 15 13 13 9 15 7 9 15 1 9 9 13 1 9 0 13 1 9 9 2
41 7 13 8 1 9 15 1 9 13 15 1 15 9 1 9 9 8 8 1 9 0 1 9 1 0 9 1 7 2 9 0 1 9 15 13 1 9 9 0 2 2
67 7 1 9 9 15 1 9 9 0 1 9 1 9 9 14 7 8 13 1 9 9 9 0 1 9 9 9 2 8 8 2 7 0 9 0 1 15 1 1 7 13 15 1 9 2 9 7 9 8 13 1 7 0 1 10 9 0 2 1 1 7 13 15 1 9 3 2
36 7 13 9 0 13 9 15 1 9 15 0 7 1 9 9 8 8 1 8 9 1 9 8 8 1 9 9 9 9 0 7 9 9 1 9 2
70 7 13 9 8 9 15 1 8 1 9 15 13 15 9 9 1 8 9 0 1 9 1 9 9 9 7 9 7 9 7 9 0 9 2 7 9 9 1 9 0 0 1 9 1 10 9 8 8 1 9 9 9 0 15 13 15 8 1 9 15 9 1 9 1 1 9 7 9 9 2
34 7 13 8 1 7 15 14 13 1 10 9 15 13 1 9 2 0 9 1 9 9 7 9 0 1 9 0 9 9 9 7 9 15 2
27 7 9 1 9 9 1 9 13 8 7 15 14 13 7 13 1 9 10 9 7 9 2 9 7 9 2 2
28 1 15 13 1 9 2 0 1 9 7 9 7 14 8 9 7 9 9 9 13 1 9 9 1 9 15 2 2
20 7 13 2 2 8 8 1 9 1 9 9 1 15 7 9 1 9 9 2 2
11 10 9 0 1 10 9 7 9 15 2 2
31 7 13 8 1 9 15 1 7 8 13 1 9 9 9 9 1 9 0 9 7 9 9 0 13 1 9 0 1 9 9 2
30 7 13 8 13 1 9 9 1 7 9 9 1 0 9 1 9 9 9 9 1 9 15 13 1 9 12 12 9 0 2
24 1 9 0 2 13 8 9 1 7 9 0 13 1 9 0 1 9 0 1 1 9 9 0 2
53 7 13 1 9 9 15 1 9 13 15 1 15 9 1 9 8 8 8 8 8 7 9 0 13 9 1 9 0 1 0 7 12 1 9 12 13 1 9 15 1 9 0 1 9 12 12 9 0 1 9 9 9 2
61 7 13 1 7 9 0 13 9 9 9 9 15 12 9 2 7 9 9 12 9 1 9 9 15 7 13 9 1 7 15 9 1 9 0 2 9 0 2 2 0 9 15 1 2 9 10 9 2 9 7 15 13 1 9 15 9 15 9 1 9 2
59 7 13 8 1 9 0 1 7 13 9 9 9 1 9 1 9 9 1 9 9 9 15 14 13 9 9 15 9 12 2 12 0 7 15 14 13 1 15 8 9 9 1 9 12 15 13 15 9 9 0 1 9 15 9 12 2 12 0 2
16 9 2 9 8 2 14 13 9 7 14 13 8 8 9 1 0
40 13 9 9 9 15 1 0 2 1 9 9 1 9 9 15 1 9 9 2 9 8 2 0 9 15 1 9 9 0 1 9 0 2 1 9 9 9 9 9 2
68 7 13 9 0 0 0 9 2 7 2 9 0 0 13 9 9 1 9 0 1 0 1 9 9 9 1 9 0 2 7 4 3 9 1 9 0 2 2 1 9 1 9 0 0 1 9 1 0 2 7 14 13 9 0 9 13 9 2 13 9 1 15 1 9 2 9 2 2
26 7 13 9 2 8 8 2 1 9 9 15 2 2 7 13 9 9 14 13 9 0 9 1 9 2 2
29 7 13 9 1 9 2 9 2 1 9 9 0 1 9 9 2 9 8 2 9 9 0 1 9 15 1 9 0 2
3 9 14 13
42 13 8 8 9 9 2 8 2 13 2 7 13 9 13 1 7 9 0 13 7 14 13 0 2 7 13 7 14 13 1 9 0 3 2 7 7 15 13 9 0 2 2
24 7 14 15 14 13 9 7 9 0 2 0 1 9 14 13 2 7 13 9 7 15 13 9 2
16 7 14 13 3 9 1 9 1 9 9 2 7 7 9 15 2
16 7 14 13 3 9 1 9 1 9 0 7 13 9 1 9 2
41 9 10 3 7 10 9 2 2 15 13 7 13 9 9 9 0 2 15 13 12 9 2 7 14 13 1 15 0 8 9 0 2 2 1 9 15 7 13 0 2 2
10 15 9 0 7 0 1 9 10 9 2
22 7 7 13 3 15 13 9 9 9 1 1 0 9 0 2 7 14 15 13 1 9 2
8 7 14 13 9 9 0 2 2
62 9 7 1 9 9 9 15 1 9 7 9 13 9 9 0 2 7 9 7 9 9 2 7 9 9 0 2 7 9 9 2 7 9 9 0 1 9 7 9 7 9 2 8 8 7 9 9 2 7 9 9 7 9 2 7 9 9 0 7 9 9 2
64 7 7 13 9 9 8 8 7 9 9 0 8 8 2 8 8 8 2 9 9 0 1 9 0 2 14 13 1 7 15 14 13 9 0 2 7 7 15 1 0 7 13 3 9 1 9 0 1 10 9 1 9 0 7 0 0 1 15 9 1 9 0 2 2
7 7 3 15 13 9 2 2
23 3 13 9 9 12 9 0 1 9 0 7 13 9 1 9 0 7 13 0 7 13 2 2
46 14 14 13 1 0 9 7 13 9 1 7 13 1 9 2 0 7 8 13 1 9 9 0 2 0 1 9 7 9 13 9 1 0 9 2 7 7 10 9 2 9 0 0 2 2 2
41 14 14 13 1 0 0 7 13 1 9 8 15 13 1 9 9 9 1 0 9 7 9 7 9 10 9 1 9 15 7 9 9 15 2 13 2 1 9 9 2 2
27 1 9 1 9 13 2 15 9 15 2 7 15 13 9 1 9 9 0 7 9 15 13 1 15 9 8 2
68 14 13 1 9 0 0 7 13 12 9 1 9 9 7 13 8 13 1 9 9 0 9 12 2 12 0 2 1 9 0 1 9 1 9 2 1 2 9 0 1 9 9 2 2 7 13 9 15 1 7 13 0 1 9 9 0 2 7 1 7 2 13 2 9 1 9 8 2
84 7 14 13 9 1 9 0 1 9 0 0 9 1 9 13 1 15 9 2 8 2 0 2 9 12 2 12 0 2 1 9 9 8 1 9 9 1 9 1 9 0 13 1 9 15 2 9 2 9 12 5 1 9 9 0 2 7 9 12 5 1 15 1 9 2 7 3 9 12 9 0 0 2 8 1 15 12 12 9 2 1 9 0 2
54 7 1 15 2 7 14 13 9 9 0 0 9 7 13 9 9 0 1 9 2 7 13 9 0 0 1 10 9 1 9 9 0 1 0 9 15 14 13 9 0 9 1 9 9 7 9 1 9 12 9 12 2 2 2
24 14 1 9 9 9 0 1 9 0 7 13 9 9 7 7 13 0 7 13 1 9 0 2 2
16 7 14 15 9 0 2 7 9 9 7 14 13 9 1 9 2
14 7 13 7 13 9 0 7 13 9 8 7 9 0 2
13 1 7 13 1 9 1 9 7 1 9 1 15 2
22 7 13 1 0 2 1 9 9 9 0 1 9 2 7 13 1 9 9 1 9 0 2
40 7 14 9 1 7 2 9 8 2 15 13 1 15 9 1 9 0 0 8 8 9 15 7 9 0 0 8 8 2 13 9 1 9 9 0 9 9 1 9 2
23 7 14 13 10 9 7 9 13 9 1 9 0 1 9 9 9 0 0 1 15 1 9 2
52 7 1 7 13 7 1 7 13 9 0 1 7 9 0 2 15 14 13 1 15 9 0 2 1 9 0 0 2 0 15 9 9 0 1 9 15 13 15 9 1 9 9 12 2 1 15 1 15 9 0 2 2
19 8 8 1 0 10 9 0 1 9 0 2 0 2 7 9 1 0 2 2
5 9 0 1 9 0
51 1 10 9 13 8 8 9 9 9 2 9 2 13 13 15 13 9 9 9 9 9 9 8 8 2 7 15 9 13 9 7 9 9 15 13 1 15 2 7 13 1 9 9 15 1 9 15 1 8 2 2
14 7 13 0 7 13 1 9 9 15 13 15 9 9 2
25 7 14 13 1 9 9 0 7 15 13 9 9 9 0 1 1 9 9 1 9 9 1 8 2 2
24 7 9 9 1 9 9 1 9 15 1 9 3 7 9 15 1 9 7 9 15 13 15 8 2
20 2 2 7 9 2 14 13 9 0 7 13 9 9 7 0 9 1 8 2 2
7 7 15 14 13 9 2 2
46 7 15 13 9 10 9 1 8 2 1 9 9 15 1 9 1 9 8 1 9 0 2 7 1 9 0 9 1 9 9 8 9 1 9 0 7 9 1 9 9 1 9 7 9 2 2
12 7 13 15 13 1 15 15 13 10 9 2 2
31 7 14 14 13 9 0 1 9 1 9 0 1 15 2 7 0 1 0 9 9 15 13 15 1 8 1 8 1 8 2 2
14 7 13 1 15 10 9 9 9 9 1 9 0 2 2
28 7 7 13 9 9 0 0 7 15 15 13 1 15 2 1 9 9 0 2 7 13 10 9 0 1 9 2 2
15 7 14 13 9 9 1 9 9 9 0 1 9 15 2 2
37 2 2 7 14 13 1 0 7 13 9 1 9 9 1 9 7 9 7 13 7 13 1 15 1 9 1 9 9 0 7 0 1 9 7 9 2 2
23 7 13 15 3 1 10 9 7 1 10 9 2 7 15 9 15 13 1 15 1 12 9 2
30 7 9 9 15 2 7 1 15 9 9 9 2 14 13 1 9 9 0 7 0 7 0 1 9 13 1 9 0 2 2
32 7 13 7 13 1 9 9 15 8 1 9 1 8 8 2 0 9 0 2 7 9 9 0 15 8 9 9 9 12 9 2 2
51 7 13 15 7 13 3 9 0 13 0 1 10 13 1 10 9 0 2 7 15 0 7 13 9 9 9 7 13 9 0 9 2 7 13 9 1 9 9 10 7 13 3 9 15 13 15 15 7 9 2 2
7 15 7 13 15 2 2 2
12 14 13 15 0 1 7 13 9 1 8 2 2
15 9 13 9 9 7 9 8 1 9 10 13 15 9 8 8
33 13 9 1 9 9 1 9 8 1 9 7 13 9 0 1 9 0 1 9 9 1 9 1 9 9 1 9 0 7 9 7 9 2
19 7 13 9 0 1 9 1 9 0 9 13 1 9 9 0 1 8 9 2
34 8 8 13 1 15 7 13 1 9 9 0 13 9 15 9 9 0 7 0 1 8 7 9 7 9 13 1 9 0 7 0 7 0 2
56 7 7 13 0 8 1 9 15 1 8 7 9 7 9 0 9 7 9 0 1 9 0 1 9 2 7 14 13 9 15 13 1 15 9 0 9 15 1 9 7 9 7 9 7 13 9 9 7 13 9 1 9 1 9 9 2
16 7 13 9 0 7 1 9 0 2 2 9 9 7 9 2 2
77 7 15 9 9 2 7 1 9 9 0 13 1 9 9 9 0 2 7 13 9 9 1 8 7 9 9 7 9 0 1 9 2 14 13 9 1 9 15 13 15 1 15 13 9 9 2 7 14 13 1 0 14 9 8 7 9 0 7 9 10 1 9 15 1 9 0 1 9 9 0 1 1 9 7 9 0 2
53 7 13 8 8 2 12 9 2 9 9 9 1 8 2 1 2 9 2 7 15 1 9 9 13 9 1 9 9 7 13 9 1 9 9 7 9 9 0 2 1 9 9 9 9 7 9 9 2 7 15 13 0 2
36 7 13 2 2 13 13 9 1 9 9 14 1 9 9 9 7 1 9 10 1 9 15 1 15 7 13 15 9 1 9 15 1 9 0 2 2
67 14 8 8 2 12 9 2 2 7 15 9 1 9 9 2 7 13 7 9 9 1 9 9 10 1 8 8 13 13 9 15 7 7 9 1 9 9 0 13 0 1 0 9 0 2 9 1 9 9 9 7 9 9 15 2 7 1 0 7 14 9 15 1 9 9 13 2
31 7 13 2 2 1 9 0 13 1 9 0 9 0 2 7 15 14 13 9 1 9 15 1 9 7 9 9 13 9 2 2
71 7 1 9 2 9 2 1 9 9 1 8 1 9 8 8 7 9 9 8 2 7 1 9 9 0 1 9 9 1 9 8 2 13 7 9 9 13 1 9 15 15 13 1 1 12 1 12 8 9 1 8 7 9 7 9 7 9 0 9 7 9 2 1 9 9 1 9 9 9 0 2
64 7 13 8 8 2 9 9 9 9 1 9 7 15 1 9 9 1 9 9 8 7 9 1 9 13 0 2 0 1 7 9 14 13 1 9 9 0 9 1 9 7 9 0 9 0 9 1 9 2 7 9 0 14 13 13 1 9 15 0 7 13 9 0 2
56 7 13 8 9 9 9 2 12 8 2 9 12 9 1 9 1 7 15 13 13 1 12 1 12 12 9 0 2 7 15 13 1 7 15 13 9 1 1 12 7 12 12 9 10 9 2 9 1 9 9 1 15 7 9 9 2
28 7 1 9 9 9 0 7 13 9 9 9 1 9 9 0 2 8 7 9 14 13 9 9 0 1 9 0 2
14 9 2 8 9 2 1 9 1 9 1 9 2 9 2
50 13 9 2 8 2 9 2 9 15 1 9 0 9 9 9 15 9 12 8 9 1 9 12 7 15 10 13 0 1 8 9 15 0 12 8 9 7 9 1 9 9 9 1 12 12 9 1 9 12 2
77 13 9 9 9 9 9 0 1 8 9 1 9 9 15 0 9 0 9 12 2 12 0 1 9 1 9 1 9 12 9 1 9 12 12 7 12 12 9 8 7 9 9 8 9 15 13 12 5 1 9 13 9 15 7 13 15 9 9 9 9 1 12 5 1 9 7 13 1 9 9 9 9 9 1 9 0 2
42 7 14 13 9 9 9 7 9 9 9 13 1 9 1 9 9 0 1 9 12 5 7 7 12 5 1 9 0 0 9 15 1 9 9 7 14 13 9 15 1 9 2
25 1 1 13 9 9 9 1 7 9 9 9 9 13 1 12 12 9 9 12 1 12 12 9 0 2
15 9 2 8 8 2 12 13 1 9 9 0 1 9 12 9
47 13 9 9 7 9 0 1 9 0 1 9 2 8 8 12 2 15 13 15 9 1 9 1 12 1 12 9 0 1 9 1 12 9 9 8 7 0 1 12 9 7 12 1 0 9 0 2
78 7 14 13 9 8 8 12 9 9 0 1 9 2 8 8 2 15 13 1 15 9 9 9 1 9 0 7 0 7 9 9 0 1 9 9 0 1 10 9 7 9 9 9 0 1 9 1 9 2 7 14 13 9 9 9 7 9 9 9 7 9 9 8 2 9 0 2 7 9 0 7 9 15 1 9 7 9 2
64 7 13 9 8 8 9 9 9 7 9 0 1 9 0 9 12 2 12 0 13 1 9 9 1 9 9 8 8 8 9 9 9 7 9 1 9 0 1 9 1 9 9 0 2 7 9 13 9 1 1 12 9 1 9 1 8 2 7 3 9 0 1 9 2
62 7 14 13 9 9 0 9 0 0 1 9 9 9 7 9 1 9 8 0 2 7 14 13 9 9 1 9 15 13 15 9 7 3 9 9 9 0 7 9 9 7 9 9 0 1 9 2 7 9 9 1 15 2 7 14 13 9 0 1 9 0 2
33 7 13 8 7 3 9 0 1 10 9 0 13 9 1 9 9 7 9 0 1 9 7 13 1 9 12 9 1 9 1 9 9 2
71 7 13 9 8 8 9 9 9 0 1 9 7 15 13 9 9 9 0 1 9 9 1 15 7 14 13 9 1 15 1 9 0 7 13 9 9 0 12 12 9 0 2 7 14 13 9 9 0 12 9 0 2 0 1 7 15 13 9 12 9 1 9 9 1 9 9 9 1 9 0 2
85 7 13 8 8 9 9 9 7 9 1 9 0 1 9 2 7 1 0 7 13 9 1 12 1 12 12 9 1 0 1 12 9 1 1 15 12 9 0 2 7 14 13 9 9 8 1 15 2 9 1 8 2 2 0 1 7 9 14 13 15 3 9 1 9 2 7 13 9 9 1 9 0 1 15 7 14 13 1 15 12 1 9 9 0 2
32 7 13 7 9 14 13 15 3 9 0 8 8 9 0 8 8 9 7 9 1 9 12 9 9 0 1 9 9 1 9 0 2
11 12 12 9 9 1 9 0 15 9 8 8
65 13 0 9 0 1 9 9 7 0 0 1 0 1 9 9 9 1 9 9 12 2 0 7 9 14 13 1 15 13 9 1 9 15 7 13 7 13 9 0 9 14 13 9 1 15 2 7 7 9 0 1 9 0 13 1 15 13 1 12 12 9 1 9 0 2
17 7 13 8 9 0 7 3 12 12 9 9 0 1 9 9 0 2
45 7 7 9 9 15 13 9 15 1 9 9 7 9 0 1 9 1 9 9 9 13 12 12 7 12 9 1 0 9 9 12 7 13 9 9 1 9 1 12 1 9 12 12 9 2
30 7 13 7 0 9 9 1 9 10 9 9 9 9 0 1 9 8 8 8 14 13 0 0 9 9 9 15 1 9 2
17 9 9 9 1 9 9 0 0 2 8 14 13 0 1 13 9 15
49 14 13 9 0 0 8 8 1 9 15 13 15 1 9 2 9 13 9 0 7 9 9 7 9 0 2 8 7 9 7 9 2 7 15 0 1 9 9 1 9 0 15 14 13 9 9 15 0 2
50 8 15 13 15 8 8 8 8 2 9 9 9 0 1 9 2 8 13 7 9 9 0 15 14 13 8 8 7 9 9 15 14 13 1 12 9 7 1 9 1 9 0 9 1 9 9 2 9 2 2
71 7 13 8 8 8 8 1 9 1 2 8 8 2 1 9 1 9 9 15 1 9 9 2 15 13 3 9 9 15 2 7 9 13 7 0 8 1 13 9 15 2 7 1 10 9 7 14 8 8 1 9 7 1 9 9 8 15 14 13 1 9 0 7 13 9 1 15 7 9 15 2
20 2 15 15 9 9 0 15 13 15 9 9 1 9 8 8 7 9 9 0 2
83 2 10 9 8 1 9 2 14 13 0 1 9 9 0 2 7 15 13 1 9 10 9 1 9 9 0 1 9 7 9 9 9 7 9 15 9 15 1 9 1 9 15 2 7 13 7 13 0 1 9 1 9 15 14 13 1 9 15 2 7 9 13 1 9 9 0 9 12 1 9 12 0 15 13 9 9 9 7 15 9 0 9 2
6 2 3 15 9 0 2
33 2 15 9 0 0 7 14 13 1 9 15 9 9 9 0 7 0 7 0 7 9 9 0 2 7 13 9 9 8 9 0 0 2
7 2 14 13 9 9 9 2
76 2 14 13 9 9 9 1 12 9 1 12 7 15 0 1 9 0 0 2 7 7 9 14 13 9 9 3 7 9 7 9 9 0 7 9 9 2 7 1 0 7 14 10 9 15 9 1 9 0 0 2 7 14 13 9 9 7 9 9 0 7 9 7 13 1 9 0 7 15 0 1 15 1 9 0 2
7 2 14 14 13 9 9 2
35 2 14 9 9 9 2 7 3 9 9 0 7 9 2 9 14 13 0 0 14 13 1 15 0 9 0 7 15 13 9 15 7 14 13 2
15 2 15 15 9 15 14 13 1 8 8 7 9 9 15 2
39 2 9 0 2 9 9 0 2 9 9 9 1 9 9 9 0 2 9 9 9 2 9 2 1 9 2 9 9 1 9 9 2 9 1 9 1 9 0 2
7 2 15 14 13 9 9 2
15 2 1 9 0 14 13 9 1 9 15 1 13 1 15 2
6 2 14 13 9 9 2
6 2 13 9 9 15 2
17 2 14 14 13 15 1 9 1 9 15 9 7 9 1 9 9 2
3 2 14 2
5 2 14 7 0 2
10 2 8 8 8 8 8 1 9 9 2
8 2 7 14 14 13 9 0 2
15 2 1 9 14 13 0 7 13 9 0 7 9 1 8 2
13 2 15 14 13 8 8 7 9 9 15 1 9 2
17 2 0 0 1 9 1 9 9 1 9 1 15 1 9 9 0 2
9 2 15 15 9 9 15 1 9 2
66 2 1 9 13 9 9 0 1 15 1 8 9 1 9 0 7 1 7 13 8 1 0 14 13 1 9 9 13 9 0 1 9 7 9 9 15 2 7 7 13 1 9 13 0 1 15 1 9 15 14 13 9 9 7 13 9 0 7 9 9 0 7 9 1 15 2
10 2 14 14 13 8 8 1 8 9 2
28 2 1 9 2 0 0 13 1 9 13 7 13 1 9 9 7 13 9 15 7 9 9 7 1 7 15 0 2
9 2 15 14 13 8 8 1 9 2
21 2 1 15 9 1 7 13 15 13 15 9 13 9 0 7 9 9 7 9 0 2
8 2 7 1 9 15 14 13 2
7 2 14 13 9 15 0 2
11 2 13 7 15 14 13 9 0 1 9 2
52 2 8 8 7 9 9 0 0 14 14 13 9 15 2 7 1 15 1 15 9 1 9 10 13 15 1 9 7 1 9 2 7 7 13 9 9 1 9 15 1 15 13 9 0 1 9 1 15 1 9 9 2
11 2 15 15 9 15 14 13 15 10 9 2
70 2 10 9 13 0 7 1 0 7 14 10 9 14 13 9 15 7 9 15 0 7 9 14 13 1 9 7 9 7 3 7 13 9 7 9 2 7 3 0 1 15 15 13 9 0 7 9 9 0 7 9 9 0 2 13 7 13 9 9 0 2 7 1 7 13 9 1 9 9 2
10 2 14 13 7 8 8 8 1 9 2
70 2 15 9 7 13 9 9 9 2 7 13 1 15 0 1 0 7 9 1 9 0 2 7 9 7 13 9 15 0 7 14 13 9 0 7 0 1 9 15 13 15 9 2 7 7 13 1 15 7 9 14 13 9 8 8 7 14 13 14 13 1 15 0 7 14 9 1 9 9 2
16 2 14 14 13 9 0 1 9 8 8 7 9 9 9 0 2
57 2 8 8 13 1 9 9 9 0 1 10 9 7 13 14 13 1 9 0 0 2 7 13 9 15 9 9 9 1 9 15 2 7 1 15 7 9 9 13 1 9 10 9 7 14 8 13 1 9 15 1 9 9 9 0 0 2
7 2 15 13 1 8 8 2
13 2 8 8 7 9 9 15 0 1 13 9 15 2
13 2 1 9 1 15 13 15 9 0 1 9 15 2
8 2 15 9 9 9 8 8 2
67 7 14 8 9 12 9 0 1 9 0 0 8 1 9 9 9 0 8 8 1 9 8 8 1 9 7 9 7 9 1 9 9 7 8 1 9 1 9 8 8 9 9 0 7 9 9 7 9 2 7 1 15 7 1 9 13 7 8 1 0 9 0 1 0 9 0 2
17 2 14 13 15 7 0 1 9 8 8 7 0 1 9 9 15 2
11 2 14 8 8 9 15 9 1 9 9 2
10 2 7 15 14 13 9 15 1 15 2
15 2 14 13 9 15 1 9 0 0 7 13 15 1 9 2
8 2 15 13 9 15 1 9 2
37 2 8 1 9 9 9 12 7 8 1 9 0 8 8 8 8 8 1 9 1 9 12 2 8 9 1 9 0 9 8 8 8 8 7 0 8 2
8 9 12 9 0 8 8 1 9
3 9 0 9
34 13 9 0 7 0 0 9 9 7 12 9 0 13 8 8 1 9 0 13 1 9 0 15 13 15 9 0 1 9 8 9 9 9 2
39 7 13 9 0 1 9 8 8 9 2 7 12 1 9 8 8 2 13 1 9 2 7 14 13 8 8 1 9 0 7 1 1 15 9 8 8 0 2 2
15 7 13 9 7 9 0 0 13 1 15 8 1 9 0 2
19 7 13 9 0 7 9 0 1 9 0 13 1 9 7 13 1 9 8 2
31 7 13 9 9 1 7 9 0 13 8 8 8 1 9 0 1 9 8 8 2 7 13 1 9 9 0 9 0 1 9 2
40 7 13 9 9 0 7 0 1 12 9 8 8 0 0 13 15 9 0 1 9 9 1 9 0 1 9 0 13 1 9 0 1 9 1 8 8 1 9 9 2
38 7 13 9 8 9 0 1 9 9 1 9 1 15 7 2 9 1 9 9 0 1 9 9 13 1 9 8 8 1 9 15 1 9 0 1 8 2 2
39 7 13 1 7 9 15 13 12 9 1 9 8 1 9 0 1 9 0 9 9 9 2 7 13 9 0 1 9 10 13 1 9 8 1 12 9 8 12 2
23 7 13 9 9 9 0 2 1 9 1 9 9 9 13 15 9 0 1 9 9 0 2 2
8 9 1 9 0 7 9 9 8
6 9 12 9 12 2 12
41 13 9 9 0 0 0 1 9 0 9 11 8 1 9 9 8 8 8 8 9 9 1 8 7 13 8 9 0 1 9 7 9 0 0 7 0 9 1 8 0 2
27 7 13 9 9 1 9 9 0 7 9 9 8 13 1 9 7 9 9 15 13 1 9 1 9 8 0 2
18 15 7 14 13 9 0 1 9 9 0 1 9 9 0 1 9 0 2
13 9 9 0 1 9 9 9 9 2 8 2 0 0
6 8 12 9 12 2 12
32 13 9 0 9 9 1 9 0 8 8 9 0 0 1 9 8 2 1 9 9 0 1 9 9 9 9 2 8 2 0 0 2
29 7 13 9 9 0 7 15 14 13 9 9 9 2 8 2 9 10 9 7 13 9 9 0 1 9 10 9 0 2
18 7 14 13 8 9 8 8 9 9 9 9 2 8 2 1 9 12 2
28 7 13 9 9 0 8 8 7 9 13 7 13 8 9 9 8 1 8 1 9 9 9 2 8 2 1 9 2
14 7 13 9 8 8 8 9 9 9 9 2 8 2 2
43 13 9 1 7 8 0 1 9 12 9 2 7 15 8 0 2 13 13 9 1 9 9 9 2 8 8 8 2 0 1 9 9 8 8 1 8 1 9 1 12 2 12 2
25 7 13 3 9 9 9 9 8 2 7 13 0 9 9 9 9 9 0 1 9 0 2 8 2 2
7 9 1 9 1 9 9 9
6 8 12 9 12 2 12
36 13 9 8 8 7 13 0 1 9 1 9 8 8 1 9 8 1 9 8 2 9 9 9 2 1 9 0 7 0 12 1 9 0 9 9 2
18 13 9 9 1 9 0 9 9 9 14 7 9 14 13 1 0 15 2
13 7 14 13 9 9 9 7 9 9 0 1 9 2
5 9 9 13 9 8
6 8 12 9 12 2 12
13 13 9 9 0 7 0 9 0 1 9 9 8 2
40 13 9 9 0 0 9 9 0 7 9 9 1 9 15 13 1 8 2 7 7 9 9 9 0 1 9 7 9 7 13 8 0 1 9 9 0 0 1 9 2
33 7 13 9 9 0 0 1 9 7 13 1 9 9 1 9 9 2 7 7 15 13 8 8 7 14 13 1 9 7 13 1 9 2
20 7 13 9 8 1 9 9 0 1 9 0 1 9 1 9 8 1 9 15 2
33 7 15 13 9 9 8 14 13 1 15 15 7 13 14 13 9 8 7 7 9 9 14 13 1 15 9 9 1 9 1 9 0 2
18 14 13 9 7 3 9 1 9 0 1 0 9 0 7 15 13 9 2
20 13 9 7 9 0 0 1 9 9 9 1 9 7 13 1 9 9 7 9 2
16 7 13 9 9 9 12 9 7 7 7 9 9 9 0 9 2
7 9 9 0 0 1 9 0
3 9 12 9
21 13 9 0 9 9 7 9 15 13 1 9 0 0 14 13 1 9 1 9 0 2
44 7 13 9 2 7 9 13 0 1 9 7 9 0 7 9 1 9 0 2 1 9 9 9 9 1 9 9 1 9 0 0 13 9 1 1 15 1 9 0 1 9 0 2 2
52 7 13 9 0 9 9 1 9 0 1 9 0 1 9 9 9 9 0 2 9 8 8 7 14 13 9 9 1 9 1 1 9 1 9 1 9 0 2 7 0 15 9 9 9 1 9 1 9 0 7 0 2
29 7 13 9 1 9 0 7 3 9 9 9 2 9 2 1 15 1 9 9 9 0 0 7 13 1 9 9 9 2
31 7 13 9 0 9 1 2 9 8 1 9 0 8 8 9 2 1 8 9 9 1 9 9 0 9 9 0 1 9 2 2
9 8 0 1 9 1 8 13 8 8
48 8 0 1 9 1 8 13 8 8 8 12 9 2 8 2 13 9 9 1 9 8 1 9 9 0 9 0 1 9 8 8 15 13 15 9 8 1 9 8 8 8 8 1 0 1 9 0 2
71 7 1 9 15 1 9 9 7 15 13 1 9 1 15 13 9 9 11 8 9 8 9 9 8 9 9 0 7 9 9 0 1 9 8 8 0 13 1 9 15 8 8 9 0 8 8 9 0 9 1 9 0 7 0 1 9 9 0 1 7 9 9 0 1 10 9 13 8 1 9 2
42 7 13 7 9 9 0 13 0 8 8 8 0 1 9 9 8 0 7 7 9 9 0 1 9 9 9 0 0 13 0 1 9 1 9 15 8 8 8 8 1 15 2
63 7 13 9 11 8 1 7 8 0 1 9 0 13 12 12 9 7 13 9 0 8 8 0 13 15 1 8 9 9 9 1 8 9 0 7 9 0 7 9 1 8 9 7 13 1 15 9 1 9 0 8 14 7 9 9 14 13 0 1 15 8 0 2
57 7 13 1 7 9 0 0 1 12 9 0 0 13 12 12 9 3 7 15 15 13 1 9 0 0 1 9 1 8 2 7 7 9 9 0 0 1 0 9 0 0 1 9 1 9 12 7 0 12 12 9 14 13 12 1 12 2
66 7 13 9 10 9 1 9 0 0 15 9 0 1 9 7 0 9 0 0 1 15 0 1 7 9 0 13 9 0 1 9 1 10 9 7 14 13 1 9 9 15 0 1 1 9 0 9 0 9 1 9 1 9 1 9 8 7 9 9 7 9 7 9 7 9 2
31 7 13 7 2 3 0 1 9 0 1 8 8 8 8 13 8 8 7 8 8 8 10 9 7 8 1 9 15 1 0 2
95 7 1 15 13 1 9 7 13 9 13 1 9 1 9 8 8 8 2 7 1 8 8 7 8 9 1 9 0 1 9 15 8 8 9 13 9 9 7 9 8 8 8 14 13 0 3 7 1 8 8 0 8 8 8 8 8 0 1 9 7 8 3 1 9 9 9 0 8 8 1 9 9 0 1 8 8 9 1 1 9 0 8 8 8 7 8 8 8 7 9 8 8 0 2 2
61 7 13 7 15 14 13 8 8 9 7 13 9 9 0 1 7 13 9 9 9 13 1 9 8 0 0 2 7 13 9 9 9 1 8 9 1 1 9 9 0 1 9 7 9 1 9 9 0 7 9 9 0 7 0 1 9 9 0 1 9 2
5 9 9 0 1 9
3 9 12 9
41 13 9 9 0 0 1 9 0 0 1 9 9 9 0 1 9 12 12 9 7 15 0 1 15 13 9 15 1 9 9 0 7 13 9 0 1 9 0 9 9 2
32 7 13 9 7 9 9 0 15 13 9 15 1 9 9 0 13 1 12 12 9 1 12 12 9 1 9 9 9 15 1 15 2
33 7 1 9 0 13 9 9 0 0 1 9 1 9 0 1 9 0 12 2 12 9 13 12 12 9 0 1 9 0 1 9 9 2
6 9 9 1 9 1 8
3 8 12 9
27 13 9 9 15 13 9 15 1 9 8 1 8 9 9 1 15 13 9 9 0 1 9 1 8 1 9 2
21 7 1 0 1 9 9 2 13 9 0 1 8 12 1 9 12 9 1 9 0 2
28 1 9 0 13 9 1 12 9 1 9 1 9 1 9 0 2 7 13 9 15 13 1 15 9 0 1 12 2
16 7 14 13 9 9 0 1 9 2 1 15 13 9 1 9 2
6 9 13 9 0 1 9
3 9 12 9
27 13 9 9 0 8 1 9 8 8 13 12 9 0 7 12 0 2 9 1 15 13 9 9 0 0 8 2
40 7 13 9 1 9 1 9 9 9 0 8 8 8 9 15 7 9 0 1 9 0 7 0 9 15 13 1 15 8 8 13 9 0 0 8 8 1 9 0 2
24 7 13 8 7 8 9 0 8 8 13 1 9 0 1 10 9 1 9 15 1 9 0 8 2
33 7 13 10 9 0 9 8 8 9 0 1 9 8 8 0 2 8 8 8 1 9 0 0 1 9 9 15 1 9 7 9 0 2
13 13 7 9 13 9 9 9 15 0 1 9 0 2
28 7 13 9 0 8 1 9 1 9 8 9 9 9 7 9 8 3 8 8 9 1 9 0 7 13 15 9 2
4 2 9 9 2
12 9 12 8 8 0 1 12 1 9 9 1 9
3 8 12 9
26 13 9 9 8 8 8 9 7 12 9 13 7 13 0 1 12 1 9 9 1 9 1 3 1 9 2
18 13 9 9 1 9 1 8 8 8 0 1 9 8 8 8 8 0 2
37 7 13 9 2 7 13 8 12 0 2 7 13 9 13 8 8 1 9 1 1 9 8 2 8 0 0 1 9 9 15 13 1 15 9 9 9 2
35 3 13 1 12 9 2 1 1 15 12 9 15 0 2 9 7 13 9 13 15 1 9 1 9 1 9 8 1 9 12 8 9 9 8 2
37 7 13 9 7 15 1 9 0 2 13 12 9 7 13 12 0 1 9 0 7 13 9 15 1 9 1 8 2 1 9 12 8 9 9 8 9 2
12 9 0 8 13 1 9 1 15 9 9 8 8
3 8 12 9
60 13 9 0 1 3 9 7 9 0 8 8 8 2 8 9 9 1 9 2 13 1 9 1 15 7 9 15 12 12 9 1 9 8 8 1 9 12 1 12 2 1 9 8 0 2 1 9 12 9 2 8 8 1 9 1 9 0 1 9 2
37 7 13 8 8 9 8 9 1 8 8 2 7 9 2 15 13 8 1 9 15 1 9 2 13 8 1 9 1 9 1 8 9 1 9 3 9 2
34 7 13 8 1 9 9 7 10 9 13 1 9 9 1 9 2 1 15 13 8 8 1 12 8 9 0 2 1 12 9 0 2 0 2
25 7 7 15 13 9 1 15 2 7 14 13 9 8 1 9 1 9 15 1 9 0 1 8 9 2
11 13 8 8 1 9 0 1 9 1 9 0
38 13 8 8 1 9 0 1 9 1 9 0 8 12 9 5 8 2 13 9 0 12 1 9 1 9 9 8 8 1 8 0 8 1 9 9 1 9 2
29 7 13 8 8 13 12 9 7 13 1 8 9 8 0 9 9 8 8 9 8 8 1 15 7 9 1 9 0 2
44 7 14 13 8 8 13 1 15 9 8 8 8 0 1 9 0 7 7 15 14 13 1 9 15 1 9 0 1 9 12 9 0 1 9 1 9 0 7 8 8 8 9 8 2
39 7 14 13 0 1 9 8 0 9 0 1 9 0 1 8 9 1 9 0 1 9 1 9 8 8 2 8 15 1 0 7 13 1 9 8 8 1 12 2
37 7 14 13 9 9 15 13 0 1 9 9 1 9 0 1 9 1 7 13 9 9 0 1 12 9 12 7 1 9 1 9 8 0 9 1 9 2
30 13 9 8 0 9 0 1 9 8 8 8 15 13 9 0 7 15 14 13 0 1 12 1 12 1 9 1 9 8 2
79 7 1 9 1 9 12 7 15 8 8 1 9 8 8 8 8 1 8 7 8 8 1 8 7 8 8 1 8 0 7 9 15 8 1 9 9 7 8 8 1 8 8 8 8 2 8 1 8 8 8 1 9 9 8 8 8 9 0 8 8 8 8 7 15 9 9 9 0 7 9 0 8 8 7 15 9 1 8 2
7 9 0 13 9 9 1 8
3 8 12 9
35 13 9 9 7 9 0 1 9 15 0 1 9 9 7 9 1 9 15 1 8 9 0 0 2 8 2 2 9 1 15 13 9 9 9 2
38 7 14 13 9 0 8 8 1 9 0 1 8 1 9 15 0 1 9 1 9 15 1 8 2 0 1 7 8 1 9 1 9 9 1 9 9 15 2
57 7 1 9 1 9 0 8 8 8 2 13 9 8 8 8 1 9 0 15 13 15 9 0 1 9 8 2 0 1 9 15 1 7 13 9 9 7 9 1 9 9 0 1 8 2 7 7 13 9 0 1 9 15 1 9 0 2
52 7 13 9 9 8 8 8 2 1 9 1 9 9 9 8 8 8 7 9 15 8 1 9 9 8 8 9 1 9 1 9 8 7 9 1 15 2 0 1 9 15 1 9 0 1 9 8 1 0 9 0 2
28 7 13 9 0 0 1 8 1 9 15 1 9 0 2 7 9 15 0 1 7 13 9 1 8 1 9 0 2
27 7 1 9 0 2 13 9 9 1 9 12 12 8 2 1 12 12 9 0 2 1 9 9 1 9 8 2
4 9 0 1 9
3 8 12 9
38 13 9 9 0 0 15 13 9 2 8 8 9 9 9 9 15 15 14 13 9 0 1 9 1 9 0 9 15 2 1 15 13 9 0 1 9 0 2
31 7 13 9 9 15 7 8 13 9 7 1 1 15 9 9 8 1 9 9 7 8 9 8 8 1 0 13 1 9 15 2
20 14 7 9 13 1 9 9 15 14 13 15 9 8 11 8 3 1 8 8 2
45 7 13 10 9 12 9 7 12 9 0 2 1 15 8 13 15 7 13 13 15 9 11 8 8 13 15 9 9 9 8 1 9 1 9 8 8 9 0 0 8 8 1 8 12 2
10 9 2 9 12 9 1 9 9 1 8
3 8 12 9
39 13 8 13 8 9 9 1 9 8 0 9 7 12 9 13 8 8 1 7 13 15 9 9 8 12 15 13 13 9 1 8 1 9 8 0 9 3 9 2
26 7 13 8 1 9 7 9 8 9 13 9 1 9 12 8 9 2 12 9 2 1 9 8 2 8 2
13 7 7 15 14 13 9 9 15 13 1 9 9 2
24 13 9 1 9 1 12 9 1 9 9 2 7 13 9 9 1 9 7 9 1 15 1 8 2
22 7 14 13 9 9 1 8 0 7 9 13 9 9 2 7 7 15 14 13 9 9 2
19 7 13 9 1 9 8 0 7 15 13 7 13 12 9 14 13 9 1 9
11 9 12 9 1 9 0 1 9 1 9 9
4 8 8 12 9
41 13 12 9 1 0 1 15 12 0 7 9 1 9 9 1 9 0 1 9 15 13 1 15 9 1 9 2 1 1 13 12 0 1 10 9 15 13 1 9 0 2
46 7 13 8 0 1 8 9 8 7 9 1 9 9 0 13 7 13 12 1 9 9 7 13 9 9 0 8 1 9 8 8 1 8 1 9 8 8 8 8 1 9 0 1 9 9 2
20 7 13 9 15 13 15 9 1 9 8 1 9 1 8 9 1 9 1 9 2
14 7 1 9 13 9 7 13 0 1 9 0 9 0 2
13 7 13 9 7 9 0 13 1 9 1 9 9 2
18 7 13 9 9 0 7 13 9 1 9 9 1 9 9 1 9 9 2
30 7 13 9 7 13 9 0 1 15 0 7 13 9 9 1 9 1 9 1 8 8 8 8 8 1 9 8 9 8 2
26 7 13 9 1 0 1 9 8 1 9 7 9 9 1 8 8 8 1 9 1 8 1 9 8 9 2
20 7 13 9 0 8 8 1 8 1 9 9 1 8 8 1 9 8 3 9 2
22 7 13 8 9 9 9 9 1 8 1 9 9 1 9 8 8 1 9 8 9 9 2
42 7 1 9 0 2 13 0 1 9 8 8 8 8 1 9 8 1 8 1 9 9 7 9 2 7 13 0 0 7 13 9 9 15 1 9 8 1 9 8 8 9 2
23 7 14 13 12 1 9 0 1 9 9 1 9 9 1 15 13 15 9 9 8 8 0 2
